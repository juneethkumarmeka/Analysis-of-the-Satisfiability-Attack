module basic_1000_10000_1500_100_levels_5xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nand U0 (N_0,In_881,In_289);
nand U1 (N_1,In_388,In_73);
and U2 (N_2,In_718,In_311);
or U3 (N_3,In_13,In_361);
and U4 (N_4,In_31,In_454);
nor U5 (N_5,In_760,In_468);
and U6 (N_6,In_800,In_834);
nor U7 (N_7,In_112,In_960);
nor U8 (N_8,In_839,In_195);
or U9 (N_9,In_652,In_461);
and U10 (N_10,In_646,In_301);
nor U11 (N_11,In_495,In_385);
nor U12 (N_12,In_169,In_623);
or U13 (N_13,In_231,In_284);
and U14 (N_14,In_151,In_903);
and U15 (N_15,In_738,In_912);
and U16 (N_16,In_191,In_547);
nor U17 (N_17,In_778,In_935);
and U18 (N_18,In_793,In_650);
nand U19 (N_19,In_210,In_619);
xor U20 (N_20,In_715,In_208);
or U21 (N_21,In_405,In_993);
or U22 (N_22,In_844,In_261);
nor U23 (N_23,In_675,In_350);
or U24 (N_24,In_882,In_494);
nor U25 (N_25,In_876,In_2);
and U26 (N_26,In_327,In_404);
xor U27 (N_27,In_434,In_355);
nand U28 (N_28,In_362,In_937);
nand U29 (N_29,In_473,In_807);
and U30 (N_30,In_310,In_471);
or U31 (N_31,In_482,In_918);
xor U32 (N_32,In_747,In_653);
nand U33 (N_33,In_886,In_833);
or U34 (N_34,In_415,In_382);
and U35 (N_35,In_459,In_896);
or U36 (N_36,In_117,In_501);
or U37 (N_37,In_865,In_828);
nor U38 (N_38,In_181,In_608);
or U39 (N_39,In_846,In_47);
or U40 (N_40,In_312,In_54);
and U41 (N_41,In_368,In_752);
or U42 (N_42,In_589,In_956);
and U43 (N_43,In_32,In_640);
and U44 (N_44,In_427,In_445);
and U45 (N_45,In_635,In_342);
and U46 (N_46,In_426,In_153);
and U47 (N_47,In_411,In_672);
xor U48 (N_48,In_814,In_82);
nand U49 (N_49,In_103,In_880);
or U50 (N_50,In_934,In_709);
and U51 (N_51,In_384,In_787);
nor U52 (N_52,In_353,In_146);
nand U53 (N_53,In_70,In_430);
nand U54 (N_54,In_546,In_509);
and U55 (N_55,In_269,In_376);
or U56 (N_56,In_543,In_618);
nor U57 (N_57,In_663,In_160);
xnor U58 (N_58,In_780,In_976);
or U59 (N_59,In_651,In_65);
nand U60 (N_60,In_120,In_945);
xnor U61 (N_61,In_830,In_741);
nor U62 (N_62,In_28,In_457);
and U63 (N_63,In_895,In_989);
and U64 (N_64,In_917,In_902);
and U65 (N_65,In_321,In_161);
xor U66 (N_66,In_818,In_176);
or U67 (N_67,In_726,In_433);
and U68 (N_68,In_229,In_308);
nand U69 (N_69,In_262,In_629);
xor U70 (N_70,In_811,In_346);
or U71 (N_71,In_343,In_140);
nand U72 (N_72,In_569,In_111);
or U73 (N_73,In_802,In_334);
nor U74 (N_74,In_21,In_467);
nand U75 (N_75,In_98,In_557);
nor U76 (N_76,In_978,In_615);
or U77 (N_77,In_227,In_237);
and U78 (N_78,In_891,In_254);
nor U79 (N_79,In_252,In_40);
or U80 (N_80,In_774,In_617);
nor U81 (N_81,In_870,In_363);
or U82 (N_82,In_916,In_720);
nor U83 (N_83,In_131,In_668);
or U84 (N_84,In_568,In_959);
or U85 (N_85,In_658,In_822);
nand U86 (N_86,In_705,In_743);
or U87 (N_87,In_123,In_590);
and U88 (N_88,In_507,In_690);
nand U89 (N_89,In_474,In_628);
or U90 (N_90,In_158,In_132);
nand U91 (N_91,In_330,In_722);
nor U92 (N_92,In_367,In_566);
nand U93 (N_93,In_729,In_483);
xnor U94 (N_94,In_148,In_128);
nand U95 (N_95,In_662,In_298);
and U96 (N_96,In_12,In_145);
nor U97 (N_97,In_186,In_126);
nor U98 (N_98,In_366,In_877);
nor U99 (N_99,In_533,In_612);
and U100 (N_100,N_61,In_719);
or U101 (N_101,In_528,In_274);
and U102 (N_102,N_77,N_95);
or U103 (N_103,In_276,In_241);
nor U104 (N_104,In_183,In_267);
nor U105 (N_105,In_104,N_86);
nor U106 (N_106,In_607,In_108);
nor U107 (N_107,In_759,In_397);
and U108 (N_108,N_84,In_998);
and U109 (N_109,In_440,N_4);
nor U110 (N_110,In_290,In_6);
and U111 (N_111,In_913,N_67);
nand U112 (N_112,In_673,In_391);
or U113 (N_113,In_990,In_666);
or U114 (N_114,In_874,In_849);
and U115 (N_115,In_323,In_523);
xor U116 (N_116,In_700,In_88);
or U117 (N_117,N_66,In_643);
xnor U118 (N_118,In_232,N_75);
nor U119 (N_119,In_531,In_41);
nor U120 (N_120,In_777,In_947);
nor U121 (N_121,N_5,N_51);
and U122 (N_122,N_0,In_857);
nand U123 (N_123,In_889,In_18);
nand U124 (N_124,N_1,In_636);
nor U125 (N_125,In_163,In_226);
or U126 (N_126,In_453,In_683);
nor U127 (N_127,In_809,In_357);
nor U128 (N_128,In_16,In_378);
or U129 (N_129,In_214,N_62);
and U130 (N_130,In_182,N_88);
and U131 (N_131,In_522,In_86);
nor U132 (N_132,In_130,In_239);
or U133 (N_133,In_105,In_565);
nor U134 (N_134,In_517,In_712);
xor U135 (N_135,In_475,In_548);
or U136 (N_136,In_905,In_399);
or U137 (N_137,In_463,In_801);
nand U138 (N_138,In_481,In_837);
nand U139 (N_139,In_806,In_604);
nor U140 (N_140,In_121,In_825);
and U141 (N_141,In_62,In_696);
nand U142 (N_142,In_894,In_413);
xnor U143 (N_143,In_34,N_68);
xnor U144 (N_144,In_782,In_33);
and U145 (N_145,In_24,N_93);
nand U146 (N_146,In_238,In_256);
nand U147 (N_147,In_742,In_178);
nor U148 (N_148,In_554,In_948);
nand U149 (N_149,In_460,In_133);
nor U150 (N_150,In_100,In_477);
and U151 (N_151,N_85,In_744);
or U152 (N_152,In_358,In_168);
nor U153 (N_153,In_584,In_717);
or U154 (N_154,In_39,In_694);
and U155 (N_155,In_570,In_975);
nor U156 (N_156,In_863,In_728);
nand U157 (N_157,In_869,In_0);
nand U158 (N_158,N_64,In_539);
nand U159 (N_159,In_724,In_671);
nor U160 (N_160,In_637,In_42);
or U161 (N_161,In_253,In_544);
nand U162 (N_162,In_841,In_390);
and U163 (N_163,In_213,In_386);
or U164 (N_164,In_419,In_952);
or U165 (N_165,In_389,In_198);
and U166 (N_166,In_138,In_446);
nand U167 (N_167,In_217,In_506);
or U168 (N_168,N_55,In_351);
nand U169 (N_169,In_771,In_188);
nand U170 (N_170,In_664,In_223);
nand U171 (N_171,In_740,In_83);
and U172 (N_172,In_502,In_278);
nor U173 (N_173,In_27,In_769);
nand U174 (N_174,In_603,In_260);
nand U175 (N_175,In_598,In_354);
and U176 (N_176,In_529,In_414);
nor U177 (N_177,In_536,In_788);
or U178 (N_178,In_964,In_450);
nor U179 (N_179,In_746,In_871);
nor U180 (N_180,In_748,In_418);
nor U181 (N_181,N_89,In_927);
nor U182 (N_182,In_957,In_470);
nand U183 (N_183,N_65,In_71);
nand U184 (N_184,In_46,N_31);
nand U185 (N_185,In_721,In_550);
or U186 (N_186,In_973,In_572);
nand U187 (N_187,In_134,In_885);
and U188 (N_188,In_375,In_94);
nand U189 (N_189,In_906,In_713);
and U190 (N_190,In_562,In_981);
nand U191 (N_191,In_551,In_630);
and U192 (N_192,In_84,N_96);
and U193 (N_193,In_703,In_19);
or U194 (N_194,N_79,In_725);
nor U195 (N_195,In_189,In_275);
or U196 (N_196,In_966,In_784);
nor U197 (N_197,N_42,In_365);
and U198 (N_198,In_320,In_63);
nand U199 (N_199,In_144,In_224);
or U200 (N_200,In_710,N_191);
nand U201 (N_201,In_85,In_369);
and U202 (N_202,In_753,In_398);
or U203 (N_203,In_974,In_72);
and U204 (N_204,In_115,In_349);
and U205 (N_205,In_90,In_395);
nand U206 (N_206,In_1,In_676);
or U207 (N_207,In_737,In_602);
nor U208 (N_208,In_949,N_17);
xor U209 (N_209,N_73,N_139);
nor U210 (N_210,In_555,In_393);
or U211 (N_211,In_215,N_9);
and U212 (N_212,N_125,In_122);
or U213 (N_213,In_707,In_597);
nand U214 (N_214,In_435,In_518);
or U215 (N_215,In_204,In_448);
xor U216 (N_216,In_986,In_45);
and U217 (N_217,N_190,In_665);
xor U218 (N_218,In_794,In_273);
nor U219 (N_219,In_827,N_80);
or U220 (N_220,In_988,N_39);
nand U221 (N_221,In_594,In_69);
and U222 (N_222,In_820,N_38);
nor U223 (N_223,In_970,In_341);
nor U224 (N_224,In_792,N_126);
nor U225 (N_225,In_401,In_36);
nand U226 (N_226,In_693,In_832);
xor U227 (N_227,In_734,In_489);
or U228 (N_228,In_35,In_466);
nor U229 (N_229,N_111,In_236);
nand U230 (N_230,In_244,In_684);
or U231 (N_231,In_864,In_883);
nand U232 (N_232,In_485,N_158);
and U233 (N_233,N_37,In_412);
nor U234 (N_234,In_867,In_135);
xor U235 (N_235,In_170,In_823);
or U236 (N_236,In_266,In_200);
nand U237 (N_237,In_255,In_3);
and U238 (N_238,In_689,In_931);
nor U239 (N_239,In_68,In_687);
and U240 (N_240,In_873,In_451);
nand U241 (N_241,N_197,In_297);
nand U242 (N_242,In_288,In_639);
nor U243 (N_243,N_109,In_862);
nor U244 (N_244,In_424,In_348);
or U245 (N_245,In_851,In_556);
nand U246 (N_246,In_534,N_110);
or U247 (N_247,In_125,In_767);
xnor U248 (N_248,In_513,In_776);
and U249 (N_249,In_152,In_541);
xnor U250 (N_250,N_167,In_464);
nor U251 (N_251,In_406,In_951);
nor U252 (N_252,In_829,N_154);
or U253 (N_253,In_439,In_516);
or U254 (N_254,In_519,In_55);
xor U255 (N_255,In_206,In_858);
and U256 (N_256,In_421,N_170);
and U257 (N_257,N_177,In_174);
nor U258 (N_258,In_370,N_143);
nand U259 (N_259,In_257,In_600);
nand U260 (N_260,N_172,In_765);
nand U261 (N_261,In_831,In_521);
nand U262 (N_262,In_129,In_296);
nand U263 (N_263,N_171,In_379);
or U264 (N_264,In_933,N_99);
or U265 (N_265,In_567,In_136);
nand U266 (N_266,In_246,In_167);
or U267 (N_267,In_842,In_797);
and U268 (N_268,N_108,In_972);
and U269 (N_269,In_968,In_591);
or U270 (N_270,N_194,In_925);
nor U271 (N_271,In_924,In_904);
nand U272 (N_272,In_585,In_372);
or U273 (N_273,N_60,N_193);
nand U274 (N_274,N_182,In_142);
or U275 (N_275,N_13,In_581);
nor U276 (N_276,In_815,In_150);
nor U277 (N_277,N_72,In_798);
nand U278 (N_278,In_22,In_808);
nand U279 (N_279,N_57,In_940);
nand U280 (N_280,In_209,In_929);
nand U281 (N_281,In_763,N_175);
or U282 (N_282,In_219,N_140);
or U283 (N_283,In_340,In_704);
nand U284 (N_284,N_132,In_279);
nand U285 (N_285,In_697,In_627);
and U286 (N_286,In_9,N_159);
and U287 (N_287,In_96,In_428);
nor U288 (N_288,In_486,In_271);
or U289 (N_289,In_243,N_50);
xor U290 (N_290,N_98,In_932);
and U291 (N_291,In_491,In_383);
or U292 (N_292,In_810,N_7);
nand U293 (N_293,N_56,In_558);
xor U294 (N_294,N_102,In_240);
nand U295 (N_295,N_169,In_272);
nor U296 (N_296,In_190,In_852);
nand U297 (N_297,N_36,N_101);
nor U298 (N_298,In_901,In_848);
nand U299 (N_299,In_282,In_364);
xnor U300 (N_300,In_80,N_92);
and U301 (N_301,In_587,N_49);
nor U302 (N_302,N_236,In_443);
and U303 (N_303,N_78,In_309);
or U304 (N_304,N_155,In_184);
xnor U305 (N_305,In_307,In_711);
or U306 (N_306,In_292,In_119);
xnor U307 (N_307,In_141,N_295);
and U308 (N_308,N_12,In_324);
and U309 (N_309,In_754,N_298);
nand U310 (N_310,In_632,N_52);
nand U311 (N_311,In_579,N_229);
nand U312 (N_312,In_884,In_772);
or U313 (N_313,In_954,In_992);
nor U314 (N_314,In_235,In_157);
nor U315 (N_315,In_766,In_498);
and U316 (N_316,In_835,N_245);
and U317 (N_317,In_840,In_775);
or U318 (N_318,In_736,In_245);
nor U319 (N_319,N_294,In_29);
or U320 (N_320,N_87,In_682);
nor U321 (N_321,In_890,N_216);
or U322 (N_322,In_611,In_4);
nor U323 (N_323,In_898,N_25);
xor U324 (N_324,In_878,N_127);
or U325 (N_325,N_181,In_124);
nor U326 (N_326,In_638,In_345);
nand U327 (N_327,N_244,In_50);
xor U328 (N_328,In_249,In_751);
and U329 (N_329,N_286,In_212);
xnor U330 (N_330,In_429,In_95);
nor U331 (N_331,N_149,In_971);
or U332 (N_332,In_270,N_43);
xnor U333 (N_333,In_165,In_394);
and U334 (N_334,In_625,In_48);
or U335 (N_335,In_53,In_511);
nor U336 (N_336,In_234,In_530);
nand U337 (N_337,In_51,In_796);
and U338 (N_338,In_432,In_113);
or U339 (N_339,N_144,In_263);
nor U340 (N_340,In_392,N_48);
or U341 (N_341,In_688,In_764);
nor U342 (N_342,In_695,In_407);
xor U343 (N_343,N_166,N_131);
or U344 (N_344,In_921,In_911);
nor U345 (N_345,N_90,In_762);
nor U346 (N_346,N_145,N_157);
nor U347 (N_347,N_271,N_100);
nand U348 (N_348,In_211,In_985);
nor U349 (N_349,In_75,N_264);
and U350 (N_350,In_164,In_425);
or U351 (N_351,N_82,In_331);
nand U352 (N_352,In_680,In_706);
xnor U353 (N_353,N_225,N_196);
or U354 (N_354,In_396,In_553);
or U355 (N_355,N_122,In_171);
xnor U356 (N_356,In_159,In_739);
nor U357 (N_357,N_185,In_866);
and U358 (N_358,In_89,In_980);
nor U359 (N_359,N_265,In_679);
or U360 (N_360,N_198,In_573);
nand U361 (N_361,N_201,In_804);
nand U362 (N_362,In_879,In_423);
and U363 (N_363,N_32,In_892);
nand U364 (N_364,In_17,In_487);
xor U365 (N_365,In_437,In_337);
nor U366 (N_366,In_549,In_175);
xnor U367 (N_367,N_287,N_234);
nor U368 (N_368,N_239,N_40);
or U369 (N_369,N_248,In_532);
nor U370 (N_370,In_381,In_561);
nor U371 (N_371,In_908,In_180);
or U372 (N_372,In_922,In_941);
and U373 (N_373,In_484,N_29);
or U374 (N_374,In_660,In_781);
nand U375 (N_375,In_854,In_93);
and U376 (N_376,N_11,In_699);
and U377 (N_377,In_76,In_930);
nor U378 (N_378,In_524,N_262);
and U379 (N_379,N_137,N_117);
or U380 (N_380,N_231,In_400);
or U381 (N_381,In_649,N_81);
nor U382 (N_382,In_610,N_156);
and U383 (N_383,In_520,In_199);
nor U384 (N_384,N_266,In_155);
or U385 (N_385,In_476,N_16);
nand U386 (N_386,In_535,In_803);
nor U387 (N_387,N_14,In_527);
and U388 (N_388,In_220,In_586);
nor U389 (N_389,In_909,In_943);
nand U390 (N_390,N_163,In_979);
nor U391 (N_391,In_860,N_176);
nand U392 (N_392,In_222,In_66);
and U393 (N_393,N_112,In_563);
nand U394 (N_394,In_387,N_97);
nand U395 (N_395,In_25,In_698);
or U396 (N_396,In_571,N_45);
xnor U397 (N_397,N_135,N_289);
and U398 (N_398,In_681,N_281);
and U399 (N_399,In_791,N_76);
xor U400 (N_400,N_189,N_369);
nor U401 (N_401,In_838,N_58);
or U402 (N_402,In_304,In_983);
xnor U403 (N_403,N_399,N_376);
nand U404 (N_404,N_6,N_272);
nor U405 (N_405,In_730,In_642);
and U406 (N_406,In_455,N_378);
or U407 (N_407,N_34,In_299);
nand U408 (N_408,In_647,In_512);
or U409 (N_409,In_773,In_295);
and U410 (N_410,In_961,In_907);
nor U411 (N_411,N_199,In_982);
or U412 (N_412,In_196,N_346);
xnor U413 (N_413,N_288,In_622);
nand U414 (N_414,In_655,In_770);
or U415 (N_415,N_284,N_382);
and U416 (N_416,N_377,In_356);
nand U417 (N_417,N_240,In_963);
or U418 (N_418,In_677,N_195);
or U419 (N_419,In_438,In_166);
or U420 (N_420,N_152,In_493);
and U421 (N_421,In_187,In_995);
nand U422 (N_422,In_23,N_116);
nor U423 (N_423,N_230,In_657);
and U424 (N_424,In_11,N_70);
nand U425 (N_425,N_304,In_325);
nor U426 (N_426,In_205,N_2);
nor U427 (N_427,N_383,In_592);
or U428 (N_428,N_308,N_279);
nand U429 (N_429,In_149,In_686);
or U430 (N_430,N_360,In_179);
nor U431 (N_431,N_41,N_277);
nand U432 (N_432,In_410,N_337);
or U433 (N_433,N_328,In_735);
and U434 (N_434,N_358,In_559);
or U435 (N_435,In_755,N_344);
nand U436 (N_436,N_254,N_71);
or U437 (N_437,In_795,In_656);
nand U438 (N_438,In_59,In_942);
or U439 (N_439,N_343,In_305);
and U440 (N_440,N_345,N_124);
xnor U441 (N_441,N_219,In_514);
or U442 (N_442,N_207,In_944);
nor U443 (N_443,In_914,In_207);
or U444 (N_444,In_708,In_286);
nor U445 (N_445,In_785,In_302);
and U446 (N_446,N_178,In_661);
nor U447 (N_447,N_379,In_251);
nor U448 (N_448,N_370,In_458);
or U449 (N_449,In_109,In_605);
nor U450 (N_450,N_119,In_230);
nor U451 (N_451,In_8,N_291);
nor U452 (N_452,In_503,N_148);
or U453 (N_453,In_44,In_380);
nand U454 (N_454,In_601,In_81);
nand U455 (N_455,N_373,N_368);
nor U456 (N_456,In_847,N_251);
or U457 (N_457,In_616,In_552);
nand U458 (N_458,N_183,N_256);
nand U459 (N_459,In_371,N_300);
or U460 (N_460,In_248,N_69);
nand U461 (N_461,N_312,In_107);
nand U462 (N_462,In_303,In_56);
nor U463 (N_463,In_172,In_875);
nand U464 (N_464,N_332,N_226);
xor U465 (N_465,In_291,N_237);
and U466 (N_466,N_363,In_283);
nand U467 (N_467,In_621,N_359);
or U468 (N_468,N_223,N_320);
or U469 (N_469,N_329,N_347);
and U470 (N_470,In_670,N_121);
or U471 (N_471,In_139,In_669);
nand U472 (N_472,N_247,N_59);
xor U473 (N_473,In_329,N_209);
nand U474 (N_474,N_250,In_10);
nor U475 (N_475,N_28,In_593);
or U476 (N_476,In_315,In_319);
nand U477 (N_477,In_888,In_654);
xnor U478 (N_478,In_580,N_255);
nor U479 (N_479,In_644,N_162);
nand U480 (N_480,N_113,N_142);
or U481 (N_481,In_318,N_187);
or U482 (N_482,In_409,In_595);
nand U483 (N_483,In_201,In_761);
or U484 (N_484,In_577,In_91);
nand U485 (N_485,In_402,N_242);
nor U486 (N_486,In_685,N_273);
and U487 (N_487,In_147,N_333);
xor U488 (N_488,N_243,In_836);
or U489 (N_489,In_64,In_15);
or U490 (N_490,N_392,N_276);
nor U491 (N_491,In_78,N_238);
and U492 (N_492,N_395,In_449);
or U493 (N_493,In_61,N_310);
nand U494 (N_494,N_348,N_263);
or U495 (N_495,N_26,In_127);
xor U496 (N_496,In_92,In_816);
nand U497 (N_497,In_648,N_387);
nor U498 (N_498,In_173,In_114);
nor U499 (N_499,N_339,N_258);
or U500 (N_500,In_408,N_114);
and U501 (N_501,N_432,N_228);
and U502 (N_502,In_545,N_361);
nor U503 (N_503,N_490,In_193);
nand U504 (N_504,N_293,N_316);
or U505 (N_505,In_900,N_365);
xor U506 (N_506,In_360,N_467);
or U507 (N_507,N_391,N_173);
and U508 (N_508,In_984,N_222);
and U509 (N_509,In_897,N_129);
and U510 (N_510,In_287,N_104);
or U511 (N_511,In_280,N_321);
xor U512 (N_512,N_331,N_317);
and U513 (N_513,N_398,N_138);
or U514 (N_514,In_162,In_259);
or U515 (N_515,N_147,N_165);
or U516 (N_516,In_991,N_478);
or U517 (N_517,In_143,In_582);
nand U518 (N_518,N_401,In_950);
and U519 (N_519,In_634,In_659);
nor U520 (N_520,In_504,In_779);
and U521 (N_521,In_118,N_53);
or U522 (N_522,N_27,N_466);
xor U523 (N_523,In_994,N_472);
nand U524 (N_524,In_861,N_210);
nor U525 (N_525,N_397,N_367);
and U526 (N_526,In_332,N_390);
nand U527 (N_527,N_128,N_355);
or U528 (N_528,In_560,N_473);
or U529 (N_529,In_843,N_349);
and U530 (N_530,N_269,N_374);
xnor U531 (N_531,N_447,In_977);
nor U532 (N_532,N_306,N_74);
nor U533 (N_533,In_633,N_402);
or U534 (N_534,N_336,N_488);
or U535 (N_535,In_317,N_8);
and U536 (N_536,N_384,N_471);
xnor U537 (N_537,N_485,N_469);
and U538 (N_538,N_318,N_307);
xnor U539 (N_539,In_939,In_859);
and U540 (N_540,In_899,N_270);
and U541 (N_541,N_380,In_420);
or U542 (N_542,N_246,N_465);
nor U543 (N_543,N_452,N_445);
nor U544 (N_544,N_285,In_37);
or U545 (N_545,N_20,In_702);
nand U546 (N_546,N_441,N_410);
nand U547 (N_547,N_440,In_202);
nand U548 (N_548,N_341,In_824);
xor U549 (N_549,In_967,In_819);
and U550 (N_550,In_745,In_60);
and U551 (N_551,N_427,In_965);
nor U552 (N_552,In_441,In_526);
and U553 (N_553,In_575,N_444);
and U554 (N_554,N_430,N_352);
nand U555 (N_555,N_151,In_328);
nand U556 (N_556,N_428,In_588);
and U557 (N_557,In_338,N_417);
or U558 (N_558,N_338,N_192);
nand U559 (N_559,In_996,In_500);
xnor U560 (N_560,In_250,In_314);
and U561 (N_561,N_409,In_641);
nor U562 (N_562,N_422,N_455);
nand U563 (N_563,In_691,N_499);
or U564 (N_564,N_44,In_915);
xor U565 (N_565,N_487,In_442);
nor U566 (N_566,N_408,In_377);
and U567 (N_567,N_400,In_77);
and U568 (N_568,In_936,N_305);
and U569 (N_569,N_406,N_448);
nor U570 (N_570,N_106,N_107);
xor U571 (N_571,N_496,In_462);
xor U572 (N_572,In_58,In_43);
or U573 (N_573,N_146,In_997);
nand U574 (N_574,In_216,N_94);
or U575 (N_575,N_443,In_101);
or U576 (N_576,N_206,N_324);
nor U577 (N_577,N_479,In_731);
and U578 (N_578,N_15,N_278);
nand U579 (N_579,N_375,N_415);
or U580 (N_580,In_316,N_454);
nand U581 (N_581,In_727,N_211);
and U582 (N_582,In_923,N_202);
or U583 (N_583,N_486,N_227);
and U584 (N_584,N_260,N_493);
or U585 (N_585,In_416,In_335);
xor U586 (N_586,In_919,N_186);
nand U587 (N_587,N_292,N_436);
nor U588 (N_588,In_480,N_217);
nand U589 (N_589,N_47,N_394);
nand U590 (N_590,In_946,N_450);
or U591 (N_591,In_756,N_351);
or U592 (N_592,In_347,In_322);
xnor U593 (N_593,N_403,N_418);
nor U594 (N_594,N_184,N_188);
nand U595 (N_595,In_456,In_510);
or U596 (N_596,N_22,In_38);
or U597 (N_597,N_389,In_540);
nand U598 (N_598,N_233,N_424);
xor U599 (N_599,N_18,In_472);
nand U600 (N_600,In_749,In_497);
or U601 (N_601,In_768,In_359);
or U602 (N_602,N_388,N_533);
xor U603 (N_603,In_7,In_478);
and U604 (N_604,In_928,N_547);
nor U605 (N_605,N_203,N_591);
nand U606 (N_606,N_435,N_290);
nor U607 (N_607,In_786,N_232);
nor U608 (N_608,In_339,In_344);
xnor U609 (N_609,N_555,N_593);
nand U610 (N_610,N_587,N_554);
and U611 (N_611,In_920,N_561);
nand U612 (N_612,N_477,N_545);
nand U613 (N_613,N_160,N_296);
and U614 (N_614,N_19,In_156);
xor U615 (N_615,In_268,In_609);
nand U616 (N_616,N_414,N_572);
and U617 (N_617,N_562,N_588);
nand U618 (N_618,In_447,N_475);
or U619 (N_619,In_624,In_614);
or U620 (N_620,N_501,N_412);
and U621 (N_621,In_106,In_576);
or U622 (N_622,N_509,In_701);
and U623 (N_623,In_293,In_496);
and U624 (N_624,N_385,N_313);
nor U625 (N_625,N_470,N_212);
nand U626 (N_626,N_489,N_595);
nand U627 (N_627,In_578,In_417);
and U628 (N_628,In_714,N_224);
nand U629 (N_629,In_542,N_557);
xor U630 (N_630,In_757,In_692);
xor U631 (N_631,N_583,In_285);
nor U632 (N_632,N_558,In_999);
or U633 (N_633,In_958,In_817);
or U634 (N_634,N_453,N_537);
nor U635 (N_635,N_449,N_353);
nor U636 (N_636,N_323,N_330);
nor U637 (N_637,N_513,N_3);
nor U638 (N_638,N_208,In_203);
and U639 (N_639,N_280,N_498);
nor U640 (N_640,N_411,N_46);
xor U641 (N_641,N_105,N_526);
xnor U642 (N_642,N_274,In_281);
or U643 (N_643,In_508,N_204);
nor U644 (N_644,N_297,N_437);
nor U645 (N_645,In_277,N_268);
and U646 (N_646,In_374,N_342);
nor U647 (N_647,N_531,N_33);
xnor U648 (N_648,In_177,In_20);
or U649 (N_649,In_750,N_421);
or U650 (N_650,In_853,In_326);
and U651 (N_651,N_275,N_568);
nor U652 (N_652,In_57,N_386);
nor U653 (N_653,N_597,In_247);
and U654 (N_654,In_910,N_516);
or U655 (N_655,N_505,N_302);
and U656 (N_656,N_393,In_228);
nor U657 (N_657,N_524,N_546);
and U658 (N_658,In_716,N_525);
xor U659 (N_659,N_54,In_233);
and U660 (N_660,N_150,In_574);
nand U661 (N_661,N_23,N_419);
or U662 (N_662,N_483,N_523);
nand U663 (N_663,N_581,In_962);
and U664 (N_664,N_404,N_21);
nor U665 (N_665,N_520,N_214);
nor U666 (N_666,N_350,In_850);
nand U667 (N_667,N_327,In_821);
xnor U668 (N_668,N_579,N_480);
xor U669 (N_669,N_476,N_503);
nand U670 (N_670,N_522,N_83);
xor U671 (N_671,In_154,N_563);
nand U672 (N_672,In_953,In_613);
nand U673 (N_673,N_511,N_24);
nor U674 (N_674,In_74,N_575);
nand U675 (N_675,N_252,N_504);
nor U676 (N_676,N_301,N_457);
nor U677 (N_677,N_314,N_259);
nor U678 (N_678,N_438,N_115);
and U679 (N_679,In_887,N_594);
nand U680 (N_680,N_538,In_789);
or U681 (N_681,In_606,N_495);
xor U682 (N_682,N_573,In_926);
or U683 (N_683,N_552,N_257);
and U684 (N_684,In_102,In_306);
nor U685 (N_685,N_407,N_442);
and U686 (N_686,N_426,N_569);
and U687 (N_687,N_543,N_420);
nor U688 (N_688,N_366,N_168);
nor U689 (N_689,In_564,N_585);
nand U690 (N_690,In_732,N_362);
nor U691 (N_691,N_439,In_790);
or U692 (N_692,In_14,N_325);
and U693 (N_693,In_242,In_97);
nor U694 (N_694,In_218,In_805);
or U695 (N_695,In_465,In_403);
nand U696 (N_696,N_534,In_258);
and U697 (N_697,N_492,In_444);
or U698 (N_698,In_645,N_434);
xnor U699 (N_699,N_213,N_123);
nor U700 (N_700,N_616,N_456);
xor U701 (N_701,In_631,N_180);
xnor U702 (N_702,N_604,N_640);
nand U703 (N_703,In_116,N_519);
nand U704 (N_704,N_689,N_215);
nand U705 (N_705,N_574,In_799);
xor U706 (N_706,N_610,N_661);
nand U707 (N_707,N_512,N_507);
or U708 (N_708,In_422,N_641);
nor U709 (N_709,N_674,N_35);
or U710 (N_710,N_607,In_492);
or U711 (N_711,N_666,In_373);
or U712 (N_712,N_571,In_723);
nor U713 (N_713,N_429,N_626);
nand U714 (N_714,N_580,N_416);
nand U715 (N_715,In_845,In_783);
and U716 (N_716,N_603,In_620);
or U717 (N_717,N_590,In_30);
xor U718 (N_718,N_664,In_110);
nor U719 (N_719,In_488,N_680);
nand U720 (N_720,N_481,N_91);
nor U721 (N_721,N_482,N_663);
and U722 (N_722,N_141,In_294);
nand U723 (N_723,In_856,N_599);
nor U724 (N_724,In_490,N_606);
xor U725 (N_725,N_565,N_577);
nand U726 (N_726,N_10,In_185);
or U727 (N_727,N_696,N_205);
or U728 (N_728,N_461,In_67);
nand U729 (N_729,In_469,N_649);
nand U730 (N_730,N_634,N_697);
or U731 (N_731,N_130,N_688);
nor U732 (N_732,N_381,In_5);
and U733 (N_733,N_576,N_174);
xnor U734 (N_734,In_79,In_192);
nand U735 (N_735,N_642,N_133);
xnor U736 (N_736,N_645,N_675);
and U737 (N_737,N_584,In_987);
nor U738 (N_738,N_589,N_518);
xor U739 (N_739,N_335,N_671);
nand U740 (N_740,N_582,N_322);
nor U741 (N_741,N_235,N_315);
nand U742 (N_742,N_659,N_530);
or U743 (N_743,N_319,N_665);
or U744 (N_744,N_502,In_479);
xor U745 (N_745,N_686,N_253);
nand U746 (N_746,N_423,N_500);
or U747 (N_747,N_463,N_508);
nor U748 (N_748,N_627,N_623);
xor U749 (N_749,N_261,N_615);
nand U750 (N_750,N_695,In_826);
nor U751 (N_751,In_758,N_532);
or U752 (N_752,N_609,N_550);
nor U753 (N_753,In_221,N_536);
xor U754 (N_754,In_893,N_458);
and U755 (N_755,N_515,N_694);
nand U756 (N_756,N_699,N_687);
xnor U757 (N_757,N_600,N_425);
or U758 (N_758,N_371,N_644);
and U759 (N_759,N_356,N_283);
and U760 (N_760,In_352,In_599);
nand U761 (N_761,N_639,In_955);
and U762 (N_762,N_654,In_667);
or U763 (N_763,N_120,N_535);
xnor U764 (N_764,N_586,N_63);
nand U765 (N_765,In_525,N_153);
nand U766 (N_766,N_354,N_542);
and U767 (N_767,N_413,N_656);
or U768 (N_768,In_225,N_396);
and U769 (N_769,N_372,N_528);
or U770 (N_770,In_52,In_499);
nor U771 (N_771,N_548,N_647);
xnor U772 (N_772,N_161,N_693);
or U773 (N_773,In_333,In_197);
nor U774 (N_774,N_431,N_491);
or U775 (N_775,N_611,In_300);
nand U776 (N_776,N_685,N_459);
nor U777 (N_777,N_340,N_357);
and U778 (N_778,N_662,N_506);
and U779 (N_779,N_698,N_241);
nand U780 (N_780,N_497,N_668);
nand U781 (N_781,N_660,N_632);
or U782 (N_782,In_87,In_969);
nand U783 (N_783,N_539,N_667);
nand U784 (N_784,N_566,In_99);
xor U785 (N_785,In_855,N_544);
nand U786 (N_786,N_136,N_670);
xor U787 (N_787,N_221,N_249);
and U788 (N_788,N_602,In_872);
xor U789 (N_789,N_484,In_813);
nand U790 (N_790,In_812,N_567);
nand U791 (N_791,N_299,N_692);
or U792 (N_792,N_179,N_433);
xnor U793 (N_793,N_510,N_631);
nor U794 (N_794,N_540,N_596);
or U795 (N_795,N_218,In_626);
or U796 (N_796,In_313,N_529);
or U797 (N_797,N_681,N_556);
nor U798 (N_798,N_633,N_514);
or U799 (N_799,N_677,N_405);
xnor U800 (N_800,N_770,N_628);
xor U801 (N_801,N_636,N_311);
and U802 (N_802,N_630,N_726);
or U803 (N_803,N_710,N_614);
and U804 (N_804,N_765,In_537);
and U805 (N_805,N_756,N_712);
nand U806 (N_806,N_725,N_732);
nand U807 (N_807,N_655,N_790);
nand U808 (N_808,N_164,N_702);
nor U809 (N_809,N_672,N_451);
nor U810 (N_810,N_768,N_624);
nand U811 (N_811,N_751,N_721);
nand U812 (N_812,N_608,N_676);
and U813 (N_813,N_762,N_780);
or U814 (N_814,N_777,N_723);
nand U815 (N_815,N_737,N_714);
and U816 (N_816,N_460,N_795);
and U817 (N_817,N_598,N_740);
nor U818 (N_818,N_700,N_334);
nor U819 (N_819,N_200,N_578);
and U820 (N_820,N_570,N_708);
nor U821 (N_821,N_564,N_755);
and U822 (N_822,In_336,N_553);
and U823 (N_823,In_583,N_786);
and U824 (N_824,N_720,N_766);
and U825 (N_825,N_669,N_303);
and U826 (N_826,N_309,N_757);
and U827 (N_827,N_783,N_787);
nor U828 (N_828,N_605,N_621);
nand U829 (N_829,N_690,N_134);
xor U830 (N_830,N_736,N_773);
and U831 (N_831,N_30,N_717);
xnor U832 (N_832,N_752,N_793);
nor U833 (N_833,N_748,N_734);
nand U834 (N_834,N_635,N_781);
nor U835 (N_835,N_638,N_684);
nand U836 (N_836,N_619,N_789);
and U837 (N_837,N_775,N_760);
and U838 (N_838,N_118,N_474);
nor U839 (N_839,N_282,N_646);
nor U840 (N_840,N_653,N_749);
and U841 (N_841,N_541,N_764);
nor U842 (N_842,N_701,In_674);
nor U843 (N_843,N_617,N_763);
xnor U844 (N_844,In_938,N_560);
and U845 (N_845,N_788,In_137);
and U846 (N_846,N_559,N_754);
nor U847 (N_847,N_724,N_678);
nor U848 (N_848,N_620,N_772);
or U849 (N_849,N_778,N_753);
nand U850 (N_850,N_742,N_730);
and U851 (N_851,N_612,N_735);
nand U852 (N_852,N_792,N_326);
nand U853 (N_853,N_728,In_431);
xnor U854 (N_854,N_791,In_596);
and U855 (N_855,N_651,In_436);
nand U856 (N_856,N_521,N_648);
xnor U857 (N_857,N_650,In_733);
nand U858 (N_858,N_746,In_49);
nand U859 (N_859,N_462,In_515);
nor U860 (N_860,In_264,N_771);
or U861 (N_861,In_868,N_711);
nand U862 (N_862,N_769,N_743);
nand U863 (N_863,In_538,N_799);
and U864 (N_864,N_704,N_682);
and U865 (N_865,N_745,N_622);
and U866 (N_866,N_652,N_798);
and U867 (N_867,N_103,N_731);
xnor U868 (N_868,N_796,N_767);
or U869 (N_869,In_452,N_679);
nor U870 (N_870,N_643,N_683);
nor U871 (N_871,N_794,N_761);
nor U872 (N_872,N_776,N_716);
nor U873 (N_873,N_551,N_727);
and U874 (N_874,N_706,N_719);
or U875 (N_875,N_707,N_779);
nand U876 (N_876,N_784,N_750);
xnor U877 (N_877,N_718,N_785);
and U878 (N_878,N_774,N_637);
nand U879 (N_879,N_364,N_618);
xnor U880 (N_880,N_592,In_26);
nand U881 (N_881,N_657,N_715);
nand U882 (N_882,N_691,N_739);
nand U883 (N_883,N_549,N_744);
and U884 (N_884,N_468,N_759);
or U885 (N_885,In_194,N_741);
nand U886 (N_886,In_678,N_601);
nand U887 (N_887,N_703,N_220);
nor U888 (N_888,N_729,N_517);
nor U889 (N_889,N_494,N_705);
and U890 (N_890,In_265,N_464);
or U891 (N_891,N_625,N_722);
or U892 (N_892,N_782,N_527);
or U893 (N_893,N_446,N_738);
or U894 (N_894,N_747,N_613);
nor U895 (N_895,N_758,N_713);
and U896 (N_896,N_797,N_629);
and U897 (N_897,N_673,In_505);
nand U898 (N_898,N_709,N_658);
nor U899 (N_899,N_267,N_733);
and U900 (N_900,N_879,N_878);
or U901 (N_901,N_820,N_876);
nor U902 (N_902,N_826,N_892);
nor U903 (N_903,N_883,N_855);
and U904 (N_904,N_866,N_801);
nor U905 (N_905,N_830,N_808);
xnor U906 (N_906,N_877,N_840);
or U907 (N_907,N_857,N_850);
nand U908 (N_908,N_839,N_895);
or U909 (N_909,N_822,N_800);
nand U910 (N_910,N_865,N_885);
and U911 (N_911,N_874,N_837);
xnor U912 (N_912,N_834,N_846);
and U913 (N_913,N_856,N_864);
nor U914 (N_914,N_827,N_852);
nand U915 (N_915,N_802,N_805);
or U916 (N_916,N_854,N_860);
nand U917 (N_917,N_858,N_881);
nor U918 (N_918,N_863,N_807);
or U919 (N_919,N_823,N_886);
or U920 (N_920,N_836,N_867);
or U921 (N_921,N_811,N_825);
xor U922 (N_922,N_831,N_803);
and U923 (N_923,N_841,N_884);
xnor U924 (N_924,N_812,N_824);
nand U925 (N_925,N_887,N_838);
or U926 (N_926,N_814,N_896);
or U927 (N_927,N_851,N_848);
nand U928 (N_928,N_875,N_816);
xor U929 (N_929,N_890,N_873);
nand U930 (N_930,N_891,N_819);
nor U931 (N_931,N_870,N_880);
xnor U932 (N_932,N_889,N_871);
nor U933 (N_933,N_832,N_845);
xnor U934 (N_934,N_868,N_847);
nor U935 (N_935,N_882,N_828);
and U936 (N_936,N_821,N_842);
nor U937 (N_937,N_869,N_898);
xnor U938 (N_938,N_859,N_844);
nand U939 (N_939,N_843,N_817);
or U940 (N_940,N_810,N_853);
nand U941 (N_941,N_893,N_861);
nor U942 (N_942,N_835,N_833);
nand U943 (N_943,N_815,N_804);
or U944 (N_944,N_806,N_829);
nor U945 (N_945,N_872,N_849);
nand U946 (N_946,N_862,N_894);
nand U947 (N_947,N_897,N_899);
nor U948 (N_948,N_809,N_813);
nor U949 (N_949,N_818,N_888);
or U950 (N_950,N_811,N_871);
nand U951 (N_951,N_890,N_888);
and U952 (N_952,N_884,N_811);
and U953 (N_953,N_864,N_861);
nor U954 (N_954,N_821,N_823);
nor U955 (N_955,N_846,N_860);
or U956 (N_956,N_890,N_891);
nor U957 (N_957,N_890,N_846);
nand U958 (N_958,N_820,N_854);
nand U959 (N_959,N_830,N_868);
nand U960 (N_960,N_897,N_837);
nor U961 (N_961,N_858,N_811);
nor U962 (N_962,N_858,N_877);
nor U963 (N_963,N_869,N_886);
and U964 (N_964,N_809,N_893);
and U965 (N_965,N_834,N_839);
nand U966 (N_966,N_829,N_833);
or U967 (N_967,N_837,N_817);
and U968 (N_968,N_818,N_852);
and U969 (N_969,N_865,N_801);
and U970 (N_970,N_892,N_851);
and U971 (N_971,N_862,N_807);
nor U972 (N_972,N_810,N_857);
or U973 (N_973,N_894,N_896);
or U974 (N_974,N_875,N_826);
nand U975 (N_975,N_813,N_826);
nor U976 (N_976,N_846,N_831);
nand U977 (N_977,N_822,N_852);
nand U978 (N_978,N_803,N_808);
nand U979 (N_979,N_887,N_803);
and U980 (N_980,N_815,N_805);
and U981 (N_981,N_836,N_838);
nand U982 (N_982,N_877,N_866);
and U983 (N_983,N_837,N_800);
nor U984 (N_984,N_879,N_848);
and U985 (N_985,N_880,N_888);
and U986 (N_986,N_836,N_896);
nand U987 (N_987,N_810,N_836);
or U988 (N_988,N_894,N_857);
or U989 (N_989,N_846,N_840);
or U990 (N_990,N_894,N_863);
and U991 (N_991,N_857,N_843);
or U992 (N_992,N_852,N_819);
nor U993 (N_993,N_849,N_836);
nor U994 (N_994,N_877,N_872);
or U995 (N_995,N_885,N_863);
or U996 (N_996,N_860,N_899);
nand U997 (N_997,N_883,N_808);
xor U998 (N_998,N_879,N_801);
and U999 (N_999,N_804,N_833);
nor U1000 (N_1000,N_965,N_941);
and U1001 (N_1001,N_959,N_942);
nand U1002 (N_1002,N_992,N_943);
and U1003 (N_1003,N_962,N_976);
and U1004 (N_1004,N_988,N_905);
and U1005 (N_1005,N_931,N_956);
and U1006 (N_1006,N_929,N_975);
or U1007 (N_1007,N_982,N_924);
xor U1008 (N_1008,N_977,N_933);
nand U1009 (N_1009,N_955,N_920);
nor U1010 (N_1010,N_967,N_910);
and U1011 (N_1011,N_961,N_949);
nand U1012 (N_1012,N_948,N_914);
or U1013 (N_1013,N_947,N_971);
nand U1014 (N_1014,N_966,N_932);
and U1015 (N_1015,N_993,N_957);
nand U1016 (N_1016,N_919,N_901);
or U1017 (N_1017,N_990,N_970);
nor U1018 (N_1018,N_918,N_907);
and U1019 (N_1019,N_954,N_936);
nand U1020 (N_1020,N_923,N_902);
and U1021 (N_1021,N_935,N_978);
nand U1022 (N_1022,N_906,N_951);
nand U1023 (N_1023,N_930,N_960);
xor U1024 (N_1024,N_927,N_984);
nor U1025 (N_1025,N_999,N_958);
xor U1026 (N_1026,N_986,N_939);
nand U1027 (N_1027,N_972,N_940);
nor U1028 (N_1028,N_994,N_925);
xnor U1029 (N_1029,N_995,N_909);
or U1030 (N_1030,N_996,N_904);
nor U1031 (N_1031,N_997,N_945);
nand U1032 (N_1032,N_974,N_968);
nor U1033 (N_1033,N_963,N_900);
nand U1034 (N_1034,N_989,N_926);
nor U1035 (N_1035,N_983,N_991);
or U1036 (N_1036,N_922,N_981);
nor U1037 (N_1037,N_937,N_987);
nor U1038 (N_1038,N_946,N_912);
nor U1039 (N_1039,N_980,N_928);
or U1040 (N_1040,N_964,N_913);
nand U1041 (N_1041,N_938,N_952);
nor U1042 (N_1042,N_903,N_979);
and U1043 (N_1043,N_915,N_998);
xor U1044 (N_1044,N_908,N_921);
nor U1045 (N_1045,N_916,N_917);
nand U1046 (N_1046,N_985,N_911);
nor U1047 (N_1047,N_973,N_969);
nand U1048 (N_1048,N_944,N_953);
nor U1049 (N_1049,N_934,N_950);
or U1050 (N_1050,N_998,N_950);
or U1051 (N_1051,N_962,N_948);
or U1052 (N_1052,N_964,N_916);
nand U1053 (N_1053,N_932,N_901);
nand U1054 (N_1054,N_962,N_969);
xnor U1055 (N_1055,N_945,N_910);
or U1056 (N_1056,N_980,N_956);
and U1057 (N_1057,N_912,N_962);
and U1058 (N_1058,N_922,N_940);
nand U1059 (N_1059,N_993,N_909);
or U1060 (N_1060,N_906,N_910);
and U1061 (N_1061,N_933,N_935);
or U1062 (N_1062,N_998,N_970);
and U1063 (N_1063,N_919,N_938);
nor U1064 (N_1064,N_908,N_966);
nor U1065 (N_1065,N_910,N_990);
and U1066 (N_1066,N_908,N_923);
and U1067 (N_1067,N_919,N_952);
nor U1068 (N_1068,N_943,N_942);
nand U1069 (N_1069,N_983,N_996);
nor U1070 (N_1070,N_990,N_974);
nor U1071 (N_1071,N_959,N_973);
nand U1072 (N_1072,N_936,N_912);
nand U1073 (N_1073,N_961,N_904);
xnor U1074 (N_1074,N_924,N_956);
and U1075 (N_1075,N_911,N_947);
nor U1076 (N_1076,N_967,N_954);
nor U1077 (N_1077,N_996,N_900);
nor U1078 (N_1078,N_902,N_907);
nor U1079 (N_1079,N_944,N_964);
or U1080 (N_1080,N_948,N_904);
and U1081 (N_1081,N_903,N_921);
nor U1082 (N_1082,N_931,N_994);
nor U1083 (N_1083,N_969,N_906);
and U1084 (N_1084,N_991,N_969);
xor U1085 (N_1085,N_918,N_962);
xnor U1086 (N_1086,N_991,N_926);
and U1087 (N_1087,N_951,N_908);
nor U1088 (N_1088,N_900,N_916);
nor U1089 (N_1089,N_960,N_972);
nor U1090 (N_1090,N_937,N_963);
and U1091 (N_1091,N_954,N_908);
nor U1092 (N_1092,N_918,N_972);
nor U1093 (N_1093,N_954,N_994);
or U1094 (N_1094,N_954,N_942);
nor U1095 (N_1095,N_902,N_946);
and U1096 (N_1096,N_962,N_944);
nor U1097 (N_1097,N_917,N_965);
xnor U1098 (N_1098,N_924,N_973);
or U1099 (N_1099,N_932,N_953);
nor U1100 (N_1100,N_1054,N_1091);
nor U1101 (N_1101,N_1044,N_1048);
nor U1102 (N_1102,N_1050,N_1058);
and U1103 (N_1103,N_1002,N_1080);
xor U1104 (N_1104,N_1038,N_1037);
and U1105 (N_1105,N_1006,N_1009);
nor U1106 (N_1106,N_1071,N_1092);
and U1107 (N_1107,N_1079,N_1028);
xnor U1108 (N_1108,N_1030,N_1046);
and U1109 (N_1109,N_1036,N_1025);
or U1110 (N_1110,N_1053,N_1077);
or U1111 (N_1111,N_1001,N_1076);
nand U1112 (N_1112,N_1020,N_1035);
nand U1113 (N_1113,N_1000,N_1089);
nor U1114 (N_1114,N_1041,N_1032);
and U1115 (N_1115,N_1017,N_1068);
xnor U1116 (N_1116,N_1051,N_1082);
nand U1117 (N_1117,N_1015,N_1087);
and U1118 (N_1118,N_1013,N_1007);
xor U1119 (N_1119,N_1052,N_1043);
or U1120 (N_1120,N_1055,N_1081);
or U1121 (N_1121,N_1060,N_1099);
and U1122 (N_1122,N_1005,N_1003);
nor U1123 (N_1123,N_1069,N_1045);
nand U1124 (N_1124,N_1011,N_1021);
nand U1125 (N_1125,N_1033,N_1084);
or U1126 (N_1126,N_1098,N_1027);
nand U1127 (N_1127,N_1040,N_1074);
and U1128 (N_1128,N_1042,N_1066);
nand U1129 (N_1129,N_1008,N_1070);
nor U1130 (N_1130,N_1023,N_1075);
and U1131 (N_1131,N_1018,N_1026);
or U1132 (N_1132,N_1039,N_1090);
xnor U1133 (N_1133,N_1093,N_1016);
and U1134 (N_1134,N_1056,N_1088);
or U1135 (N_1135,N_1067,N_1047);
and U1136 (N_1136,N_1064,N_1057);
nor U1137 (N_1137,N_1004,N_1085);
or U1138 (N_1138,N_1094,N_1029);
nand U1139 (N_1139,N_1014,N_1078);
xnor U1140 (N_1140,N_1086,N_1012);
nor U1141 (N_1141,N_1024,N_1063);
and U1142 (N_1142,N_1061,N_1083);
xnor U1143 (N_1143,N_1034,N_1059);
nor U1144 (N_1144,N_1096,N_1022);
nand U1145 (N_1145,N_1010,N_1097);
nand U1146 (N_1146,N_1031,N_1072);
nor U1147 (N_1147,N_1065,N_1095);
xor U1148 (N_1148,N_1062,N_1073);
nor U1149 (N_1149,N_1019,N_1049);
and U1150 (N_1150,N_1065,N_1040);
and U1151 (N_1151,N_1007,N_1047);
nor U1152 (N_1152,N_1022,N_1037);
nand U1153 (N_1153,N_1091,N_1051);
or U1154 (N_1154,N_1001,N_1058);
or U1155 (N_1155,N_1010,N_1095);
and U1156 (N_1156,N_1031,N_1067);
xor U1157 (N_1157,N_1086,N_1035);
nor U1158 (N_1158,N_1017,N_1028);
and U1159 (N_1159,N_1078,N_1087);
nor U1160 (N_1160,N_1017,N_1082);
nand U1161 (N_1161,N_1049,N_1034);
nor U1162 (N_1162,N_1094,N_1058);
or U1163 (N_1163,N_1060,N_1064);
nand U1164 (N_1164,N_1042,N_1012);
or U1165 (N_1165,N_1024,N_1083);
nand U1166 (N_1166,N_1092,N_1033);
and U1167 (N_1167,N_1098,N_1058);
nor U1168 (N_1168,N_1079,N_1045);
nand U1169 (N_1169,N_1094,N_1013);
nor U1170 (N_1170,N_1085,N_1042);
nor U1171 (N_1171,N_1077,N_1070);
xor U1172 (N_1172,N_1005,N_1020);
and U1173 (N_1173,N_1056,N_1086);
or U1174 (N_1174,N_1036,N_1040);
xnor U1175 (N_1175,N_1001,N_1097);
xnor U1176 (N_1176,N_1078,N_1028);
xor U1177 (N_1177,N_1070,N_1033);
and U1178 (N_1178,N_1047,N_1025);
nor U1179 (N_1179,N_1027,N_1095);
and U1180 (N_1180,N_1097,N_1044);
nor U1181 (N_1181,N_1001,N_1015);
xor U1182 (N_1182,N_1033,N_1019);
nand U1183 (N_1183,N_1023,N_1083);
nor U1184 (N_1184,N_1017,N_1062);
nor U1185 (N_1185,N_1058,N_1093);
nor U1186 (N_1186,N_1054,N_1097);
or U1187 (N_1187,N_1035,N_1037);
nand U1188 (N_1188,N_1079,N_1048);
or U1189 (N_1189,N_1079,N_1069);
xnor U1190 (N_1190,N_1007,N_1091);
and U1191 (N_1191,N_1064,N_1001);
xor U1192 (N_1192,N_1082,N_1031);
xnor U1193 (N_1193,N_1045,N_1065);
nand U1194 (N_1194,N_1068,N_1035);
nand U1195 (N_1195,N_1040,N_1066);
and U1196 (N_1196,N_1069,N_1014);
nand U1197 (N_1197,N_1065,N_1032);
nor U1198 (N_1198,N_1099,N_1010);
and U1199 (N_1199,N_1008,N_1027);
nand U1200 (N_1200,N_1148,N_1104);
nor U1201 (N_1201,N_1161,N_1173);
or U1202 (N_1202,N_1183,N_1160);
nand U1203 (N_1203,N_1129,N_1138);
and U1204 (N_1204,N_1111,N_1181);
or U1205 (N_1205,N_1170,N_1100);
and U1206 (N_1206,N_1176,N_1122);
nor U1207 (N_1207,N_1126,N_1113);
or U1208 (N_1208,N_1112,N_1182);
nor U1209 (N_1209,N_1143,N_1145);
xor U1210 (N_1210,N_1174,N_1199);
or U1211 (N_1211,N_1166,N_1190);
nand U1212 (N_1212,N_1116,N_1141);
and U1213 (N_1213,N_1168,N_1107);
xnor U1214 (N_1214,N_1191,N_1198);
and U1215 (N_1215,N_1133,N_1114);
and U1216 (N_1216,N_1178,N_1184);
nor U1217 (N_1217,N_1147,N_1149);
nand U1218 (N_1218,N_1162,N_1172);
nand U1219 (N_1219,N_1123,N_1121);
or U1220 (N_1220,N_1158,N_1137);
or U1221 (N_1221,N_1106,N_1125);
nor U1222 (N_1222,N_1177,N_1142);
nor U1223 (N_1223,N_1105,N_1128);
nor U1224 (N_1224,N_1154,N_1164);
nand U1225 (N_1225,N_1108,N_1180);
nand U1226 (N_1226,N_1130,N_1194);
nand U1227 (N_1227,N_1195,N_1192);
and U1228 (N_1228,N_1193,N_1188);
and U1229 (N_1229,N_1169,N_1151);
nor U1230 (N_1230,N_1109,N_1189);
and U1231 (N_1231,N_1159,N_1120);
or U1232 (N_1232,N_1197,N_1153);
and U1233 (N_1233,N_1175,N_1102);
and U1234 (N_1234,N_1186,N_1165);
xor U1235 (N_1235,N_1119,N_1156);
nor U1236 (N_1236,N_1101,N_1196);
nand U1237 (N_1237,N_1135,N_1167);
nand U1238 (N_1238,N_1155,N_1187);
nor U1239 (N_1239,N_1124,N_1140);
or U1240 (N_1240,N_1118,N_1171);
or U1241 (N_1241,N_1110,N_1127);
or U1242 (N_1242,N_1103,N_1157);
or U1243 (N_1243,N_1136,N_1144);
nand U1244 (N_1244,N_1146,N_1132);
and U1245 (N_1245,N_1163,N_1139);
xnor U1246 (N_1246,N_1131,N_1150);
nand U1247 (N_1247,N_1185,N_1179);
and U1248 (N_1248,N_1152,N_1134);
nor U1249 (N_1249,N_1117,N_1115);
or U1250 (N_1250,N_1154,N_1120);
and U1251 (N_1251,N_1146,N_1116);
and U1252 (N_1252,N_1195,N_1111);
nand U1253 (N_1253,N_1184,N_1164);
and U1254 (N_1254,N_1146,N_1167);
and U1255 (N_1255,N_1180,N_1113);
or U1256 (N_1256,N_1101,N_1190);
nor U1257 (N_1257,N_1136,N_1179);
xor U1258 (N_1258,N_1124,N_1130);
nand U1259 (N_1259,N_1157,N_1167);
xnor U1260 (N_1260,N_1183,N_1127);
nand U1261 (N_1261,N_1194,N_1103);
nor U1262 (N_1262,N_1151,N_1170);
or U1263 (N_1263,N_1141,N_1170);
nand U1264 (N_1264,N_1149,N_1170);
and U1265 (N_1265,N_1126,N_1112);
nor U1266 (N_1266,N_1115,N_1103);
nor U1267 (N_1267,N_1137,N_1163);
nor U1268 (N_1268,N_1173,N_1149);
and U1269 (N_1269,N_1140,N_1155);
nor U1270 (N_1270,N_1133,N_1172);
xor U1271 (N_1271,N_1148,N_1177);
nand U1272 (N_1272,N_1123,N_1186);
or U1273 (N_1273,N_1117,N_1188);
or U1274 (N_1274,N_1104,N_1115);
nor U1275 (N_1275,N_1183,N_1164);
nand U1276 (N_1276,N_1121,N_1119);
or U1277 (N_1277,N_1118,N_1123);
nand U1278 (N_1278,N_1112,N_1147);
nor U1279 (N_1279,N_1175,N_1193);
and U1280 (N_1280,N_1138,N_1161);
xor U1281 (N_1281,N_1164,N_1110);
xor U1282 (N_1282,N_1189,N_1103);
or U1283 (N_1283,N_1124,N_1138);
nor U1284 (N_1284,N_1166,N_1135);
nand U1285 (N_1285,N_1157,N_1109);
or U1286 (N_1286,N_1170,N_1153);
or U1287 (N_1287,N_1154,N_1131);
nor U1288 (N_1288,N_1133,N_1121);
or U1289 (N_1289,N_1132,N_1195);
or U1290 (N_1290,N_1160,N_1143);
or U1291 (N_1291,N_1139,N_1137);
nand U1292 (N_1292,N_1169,N_1163);
nand U1293 (N_1293,N_1154,N_1102);
nand U1294 (N_1294,N_1104,N_1121);
and U1295 (N_1295,N_1110,N_1174);
or U1296 (N_1296,N_1191,N_1152);
and U1297 (N_1297,N_1187,N_1112);
nor U1298 (N_1298,N_1167,N_1193);
nor U1299 (N_1299,N_1179,N_1120);
nand U1300 (N_1300,N_1299,N_1208);
or U1301 (N_1301,N_1298,N_1212);
nor U1302 (N_1302,N_1273,N_1266);
nand U1303 (N_1303,N_1201,N_1230);
xnor U1304 (N_1304,N_1271,N_1288);
xor U1305 (N_1305,N_1236,N_1200);
xor U1306 (N_1306,N_1275,N_1203);
and U1307 (N_1307,N_1254,N_1272);
nor U1308 (N_1308,N_1213,N_1204);
nand U1309 (N_1309,N_1209,N_1256);
nor U1310 (N_1310,N_1228,N_1297);
or U1311 (N_1311,N_1286,N_1214);
nor U1312 (N_1312,N_1211,N_1202);
or U1313 (N_1313,N_1296,N_1244);
and U1314 (N_1314,N_1278,N_1227);
and U1315 (N_1315,N_1206,N_1233);
nand U1316 (N_1316,N_1249,N_1263);
or U1317 (N_1317,N_1295,N_1223);
or U1318 (N_1318,N_1262,N_1245);
xor U1319 (N_1319,N_1205,N_1284);
nor U1320 (N_1320,N_1246,N_1225);
or U1321 (N_1321,N_1287,N_1285);
and U1322 (N_1322,N_1222,N_1290);
nor U1323 (N_1323,N_1216,N_1239);
nand U1324 (N_1324,N_1267,N_1269);
nor U1325 (N_1325,N_1232,N_1240);
nand U1326 (N_1326,N_1255,N_1221);
nor U1327 (N_1327,N_1259,N_1250);
nand U1328 (N_1328,N_1293,N_1226);
nor U1329 (N_1329,N_1294,N_1210);
nand U1330 (N_1330,N_1243,N_1291);
nand U1331 (N_1331,N_1231,N_1289);
nand U1332 (N_1332,N_1270,N_1217);
and U1333 (N_1333,N_1238,N_1215);
or U1334 (N_1334,N_1252,N_1283);
and U1335 (N_1335,N_1261,N_1251);
xnor U1336 (N_1336,N_1219,N_1260);
and U1337 (N_1337,N_1257,N_1247);
nand U1338 (N_1338,N_1253,N_1279);
xor U1339 (N_1339,N_1277,N_1218);
and U1340 (N_1340,N_1229,N_1280);
or U1341 (N_1341,N_1274,N_1237);
nand U1342 (N_1342,N_1235,N_1282);
and U1343 (N_1343,N_1264,N_1220);
or U1344 (N_1344,N_1207,N_1241);
nor U1345 (N_1345,N_1234,N_1242);
xor U1346 (N_1346,N_1281,N_1276);
xor U1347 (N_1347,N_1224,N_1292);
and U1348 (N_1348,N_1258,N_1268);
and U1349 (N_1349,N_1265,N_1248);
or U1350 (N_1350,N_1210,N_1290);
and U1351 (N_1351,N_1204,N_1262);
nor U1352 (N_1352,N_1264,N_1231);
xor U1353 (N_1353,N_1280,N_1254);
or U1354 (N_1354,N_1245,N_1285);
and U1355 (N_1355,N_1233,N_1218);
nand U1356 (N_1356,N_1279,N_1220);
and U1357 (N_1357,N_1203,N_1273);
xnor U1358 (N_1358,N_1244,N_1238);
nand U1359 (N_1359,N_1254,N_1233);
or U1360 (N_1360,N_1267,N_1255);
or U1361 (N_1361,N_1232,N_1292);
nand U1362 (N_1362,N_1221,N_1235);
nor U1363 (N_1363,N_1244,N_1222);
nor U1364 (N_1364,N_1293,N_1233);
nand U1365 (N_1365,N_1200,N_1298);
xor U1366 (N_1366,N_1242,N_1217);
xor U1367 (N_1367,N_1236,N_1271);
xor U1368 (N_1368,N_1205,N_1285);
or U1369 (N_1369,N_1275,N_1235);
or U1370 (N_1370,N_1277,N_1265);
nand U1371 (N_1371,N_1222,N_1211);
and U1372 (N_1372,N_1295,N_1241);
or U1373 (N_1373,N_1294,N_1207);
and U1374 (N_1374,N_1242,N_1238);
nor U1375 (N_1375,N_1297,N_1222);
nand U1376 (N_1376,N_1278,N_1261);
and U1377 (N_1377,N_1230,N_1270);
nand U1378 (N_1378,N_1210,N_1201);
or U1379 (N_1379,N_1251,N_1280);
nor U1380 (N_1380,N_1265,N_1263);
and U1381 (N_1381,N_1209,N_1233);
nand U1382 (N_1382,N_1234,N_1227);
nand U1383 (N_1383,N_1215,N_1219);
and U1384 (N_1384,N_1295,N_1275);
xor U1385 (N_1385,N_1243,N_1200);
nor U1386 (N_1386,N_1241,N_1238);
nand U1387 (N_1387,N_1201,N_1261);
and U1388 (N_1388,N_1232,N_1223);
nand U1389 (N_1389,N_1254,N_1246);
xor U1390 (N_1390,N_1225,N_1214);
or U1391 (N_1391,N_1203,N_1207);
nor U1392 (N_1392,N_1260,N_1299);
and U1393 (N_1393,N_1210,N_1214);
and U1394 (N_1394,N_1270,N_1288);
xnor U1395 (N_1395,N_1249,N_1234);
nand U1396 (N_1396,N_1282,N_1232);
xnor U1397 (N_1397,N_1236,N_1299);
or U1398 (N_1398,N_1252,N_1288);
nand U1399 (N_1399,N_1240,N_1203);
nand U1400 (N_1400,N_1370,N_1365);
and U1401 (N_1401,N_1385,N_1330);
and U1402 (N_1402,N_1337,N_1383);
and U1403 (N_1403,N_1345,N_1347);
or U1404 (N_1404,N_1352,N_1369);
and U1405 (N_1405,N_1314,N_1343);
or U1406 (N_1406,N_1382,N_1309);
and U1407 (N_1407,N_1357,N_1329);
and U1408 (N_1408,N_1313,N_1355);
or U1409 (N_1409,N_1324,N_1316);
or U1410 (N_1410,N_1363,N_1353);
nor U1411 (N_1411,N_1304,N_1318);
nor U1412 (N_1412,N_1361,N_1341);
nor U1413 (N_1413,N_1335,N_1381);
and U1414 (N_1414,N_1392,N_1389);
nor U1415 (N_1415,N_1350,N_1379);
and U1416 (N_1416,N_1391,N_1315);
or U1417 (N_1417,N_1398,N_1367);
xnor U1418 (N_1418,N_1322,N_1378);
and U1419 (N_1419,N_1327,N_1333);
xor U1420 (N_1420,N_1388,N_1331);
nor U1421 (N_1421,N_1377,N_1303);
and U1422 (N_1422,N_1360,N_1312);
or U1423 (N_1423,N_1339,N_1328);
or U1424 (N_1424,N_1397,N_1311);
and U1425 (N_1425,N_1334,N_1344);
and U1426 (N_1426,N_1396,N_1384);
nand U1427 (N_1427,N_1321,N_1348);
nand U1428 (N_1428,N_1342,N_1371);
and U1429 (N_1429,N_1307,N_1325);
nor U1430 (N_1430,N_1375,N_1376);
nor U1431 (N_1431,N_1351,N_1399);
and U1432 (N_1432,N_1374,N_1319);
or U1433 (N_1433,N_1394,N_1306);
or U1434 (N_1434,N_1364,N_1323);
or U1435 (N_1435,N_1301,N_1359);
xor U1436 (N_1436,N_1358,N_1349);
or U1437 (N_1437,N_1300,N_1390);
nor U1438 (N_1438,N_1387,N_1332);
nand U1439 (N_1439,N_1302,N_1373);
or U1440 (N_1440,N_1386,N_1310);
and U1441 (N_1441,N_1320,N_1308);
and U1442 (N_1442,N_1340,N_1372);
nand U1443 (N_1443,N_1368,N_1356);
xor U1444 (N_1444,N_1366,N_1336);
and U1445 (N_1445,N_1354,N_1362);
and U1446 (N_1446,N_1326,N_1317);
or U1447 (N_1447,N_1338,N_1393);
or U1448 (N_1448,N_1380,N_1305);
and U1449 (N_1449,N_1395,N_1346);
or U1450 (N_1450,N_1347,N_1358);
and U1451 (N_1451,N_1391,N_1320);
xnor U1452 (N_1452,N_1338,N_1353);
and U1453 (N_1453,N_1350,N_1339);
or U1454 (N_1454,N_1326,N_1334);
nand U1455 (N_1455,N_1375,N_1368);
and U1456 (N_1456,N_1301,N_1321);
or U1457 (N_1457,N_1394,N_1376);
nand U1458 (N_1458,N_1322,N_1314);
nand U1459 (N_1459,N_1336,N_1369);
and U1460 (N_1460,N_1354,N_1395);
nor U1461 (N_1461,N_1365,N_1378);
nand U1462 (N_1462,N_1380,N_1365);
xor U1463 (N_1463,N_1366,N_1310);
or U1464 (N_1464,N_1323,N_1371);
or U1465 (N_1465,N_1391,N_1375);
nand U1466 (N_1466,N_1381,N_1312);
nand U1467 (N_1467,N_1373,N_1377);
or U1468 (N_1468,N_1344,N_1388);
or U1469 (N_1469,N_1327,N_1377);
nand U1470 (N_1470,N_1315,N_1328);
or U1471 (N_1471,N_1349,N_1382);
xnor U1472 (N_1472,N_1307,N_1374);
and U1473 (N_1473,N_1350,N_1363);
or U1474 (N_1474,N_1379,N_1364);
nand U1475 (N_1475,N_1307,N_1327);
and U1476 (N_1476,N_1304,N_1360);
and U1477 (N_1477,N_1330,N_1335);
or U1478 (N_1478,N_1337,N_1365);
nor U1479 (N_1479,N_1300,N_1328);
nor U1480 (N_1480,N_1348,N_1352);
nor U1481 (N_1481,N_1387,N_1301);
or U1482 (N_1482,N_1347,N_1399);
nand U1483 (N_1483,N_1306,N_1314);
nor U1484 (N_1484,N_1389,N_1317);
nor U1485 (N_1485,N_1378,N_1396);
nor U1486 (N_1486,N_1392,N_1342);
and U1487 (N_1487,N_1396,N_1374);
nand U1488 (N_1488,N_1329,N_1315);
or U1489 (N_1489,N_1307,N_1399);
nand U1490 (N_1490,N_1392,N_1311);
nand U1491 (N_1491,N_1311,N_1332);
nand U1492 (N_1492,N_1302,N_1353);
and U1493 (N_1493,N_1324,N_1329);
or U1494 (N_1494,N_1338,N_1308);
xor U1495 (N_1495,N_1339,N_1320);
nor U1496 (N_1496,N_1309,N_1333);
nor U1497 (N_1497,N_1348,N_1388);
nor U1498 (N_1498,N_1365,N_1364);
or U1499 (N_1499,N_1375,N_1362);
or U1500 (N_1500,N_1400,N_1462);
or U1501 (N_1501,N_1489,N_1482);
and U1502 (N_1502,N_1414,N_1490);
nand U1503 (N_1503,N_1442,N_1427);
nand U1504 (N_1504,N_1458,N_1435);
nand U1505 (N_1505,N_1478,N_1495);
or U1506 (N_1506,N_1484,N_1421);
and U1507 (N_1507,N_1460,N_1453);
and U1508 (N_1508,N_1457,N_1447);
or U1509 (N_1509,N_1405,N_1401);
xnor U1510 (N_1510,N_1424,N_1481);
xor U1511 (N_1511,N_1467,N_1402);
nand U1512 (N_1512,N_1468,N_1451);
and U1513 (N_1513,N_1450,N_1409);
xnor U1514 (N_1514,N_1404,N_1416);
xor U1515 (N_1515,N_1423,N_1408);
or U1516 (N_1516,N_1418,N_1432);
nor U1517 (N_1517,N_1493,N_1466);
nor U1518 (N_1518,N_1443,N_1475);
nand U1519 (N_1519,N_1491,N_1441);
nand U1520 (N_1520,N_1449,N_1429);
and U1521 (N_1521,N_1469,N_1479);
or U1522 (N_1522,N_1436,N_1456);
xnor U1523 (N_1523,N_1492,N_1473);
nor U1524 (N_1524,N_1412,N_1486);
xor U1525 (N_1525,N_1415,N_1448);
nand U1526 (N_1526,N_1425,N_1485);
or U1527 (N_1527,N_1470,N_1434);
or U1528 (N_1528,N_1474,N_1422);
or U1529 (N_1529,N_1472,N_1438);
nor U1530 (N_1530,N_1444,N_1480);
or U1531 (N_1531,N_1465,N_1497);
or U1532 (N_1532,N_1496,N_1413);
and U1533 (N_1533,N_1407,N_1437);
and U1534 (N_1534,N_1476,N_1410);
and U1535 (N_1535,N_1430,N_1499);
nor U1536 (N_1536,N_1454,N_1420);
or U1537 (N_1537,N_1431,N_1455);
or U1538 (N_1538,N_1440,N_1406);
nand U1539 (N_1539,N_1403,N_1445);
and U1540 (N_1540,N_1461,N_1426);
nand U1541 (N_1541,N_1494,N_1483);
nor U1542 (N_1542,N_1459,N_1498);
xor U1543 (N_1543,N_1419,N_1446);
nor U1544 (N_1544,N_1463,N_1411);
nor U1545 (N_1545,N_1439,N_1464);
nor U1546 (N_1546,N_1477,N_1428);
and U1547 (N_1547,N_1471,N_1417);
nand U1548 (N_1548,N_1487,N_1452);
or U1549 (N_1549,N_1433,N_1488);
or U1550 (N_1550,N_1494,N_1442);
nor U1551 (N_1551,N_1481,N_1449);
nor U1552 (N_1552,N_1422,N_1446);
nor U1553 (N_1553,N_1498,N_1458);
nor U1554 (N_1554,N_1419,N_1464);
and U1555 (N_1555,N_1425,N_1495);
nor U1556 (N_1556,N_1495,N_1435);
or U1557 (N_1557,N_1445,N_1404);
xor U1558 (N_1558,N_1482,N_1439);
nor U1559 (N_1559,N_1406,N_1413);
nor U1560 (N_1560,N_1452,N_1442);
nor U1561 (N_1561,N_1448,N_1441);
xnor U1562 (N_1562,N_1432,N_1404);
nor U1563 (N_1563,N_1406,N_1466);
and U1564 (N_1564,N_1487,N_1447);
and U1565 (N_1565,N_1448,N_1489);
or U1566 (N_1566,N_1479,N_1404);
nand U1567 (N_1567,N_1484,N_1462);
and U1568 (N_1568,N_1443,N_1423);
nand U1569 (N_1569,N_1412,N_1455);
nand U1570 (N_1570,N_1439,N_1448);
or U1571 (N_1571,N_1487,N_1432);
or U1572 (N_1572,N_1451,N_1478);
nor U1573 (N_1573,N_1434,N_1412);
and U1574 (N_1574,N_1463,N_1470);
nor U1575 (N_1575,N_1420,N_1452);
or U1576 (N_1576,N_1432,N_1442);
or U1577 (N_1577,N_1428,N_1421);
or U1578 (N_1578,N_1441,N_1499);
nand U1579 (N_1579,N_1433,N_1415);
nand U1580 (N_1580,N_1402,N_1414);
nor U1581 (N_1581,N_1441,N_1428);
nand U1582 (N_1582,N_1451,N_1487);
xnor U1583 (N_1583,N_1448,N_1413);
xor U1584 (N_1584,N_1499,N_1436);
nor U1585 (N_1585,N_1430,N_1460);
nand U1586 (N_1586,N_1425,N_1451);
or U1587 (N_1587,N_1452,N_1409);
and U1588 (N_1588,N_1444,N_1468);
xor U1589 (N_1589,N_1412,N_1492);
and U1590 (N_1590,N_1430,N_1473);
and U1591 (N_1591,N_1456,N_1479);
and U1592 (N_1592,N_1436,N_1486);
or U1593 (N_1593,N_1462,N_1423);
and U1594 (N_1594,N_1466,N_1473);
nand U1595 (N_1595,N_1424,N_1405);
nand U1596 (N_1596,N_1406,N_1442);
nor U1597 (N_1597,N_1443,N_1491);
or U1598 (N_1598,N_1491,N_1439);
and U1599 (N_1599,N_1477,N_1448);
and U1600 (N_1600,N_1558,N_1573);
nand U1601 (N_1601,N_1539,N_1531);
or U1602 (N_1602,N_1567,N_1524);
nor U1603 (N_1603,N_1583,N_1564);
xnor U1604 (N_1604,N_1502,N_1571);
xnor U1605 (N_1605,N_1576,N_1520);
nand U1606 (N_1606,N_1533,N_1536);
and U1607 (N_1607,N_1590,N_1588);
nand U1608 (N_1608,N_1587,N_1563);
nand U1609 (N_1609,N_1569,N_1565);
nand U1610 (N_1610,N_1549,N_1508);
nand U1611 (N_1611,N_1530,N_1527);
and U1612 (N_1612,N_1515,N_1550);
nand U1613 (N_1613,N_1514,N_1543);
or U1614 (N_1614,N_1551,N_1513);
nand U1615 (N_1615,N_1542,N_1560);
and U1616 (N_1616,N_1526,N_1580);
nand U1617 (N_1617,N_1557,N_1541);
nor U1618 (N_1618,N_1501,N_1521);
and U1619 (N_1619,N_1538,N_1582);
xnor U1620 (N_1620,N_1599,N_1504);
nand U1621 (N_1621,N_1574,N_1503);
nor U1622 (N_1622,N_1512,N_1593);
nor U1623 (N_1623,N_1586,N_1584);
or U1624 (N_1624,N_1595,N_1554);
and U1625 (N_1625,N_1509,N_1517);
nand U1626 (N_1626,N_1547,N_1500);
or U1627 (N_1627,N_1585,N_1579);
nor U1628 (N_1628,N_1570,N_1562);
xor U1629 (N_1629,N_1535,N_1511);
nor U1630 (N_1630,N_1522,N_1540);
or U1631 (N_1631,N_1552,N_1546);
nor U1632 (N_1632,N_1548,N_1506);
nor U1633 (N_1633,N_1532,N_1516);
xor U1634 (N_1634,N_1597,N_1594);
xnor U1635 (N_1635,N_1534,N_1578);
nor U1636 (N_1636,N_1523,N_1572);
or U1637 (N_1637,N_1507,N_1589);
or U1638 (N_1638,N_1525,N_1545);
nand U1639 (N_1639,N_1559,N_1561);
nand U1640 (N_1640,N_1519,N_1592);
or U1641 (N_1641,N_1537,N_1556);
and U1642 (N_1642,N_1596,N_1518);
nand U1643 (N_1643,N_1568,N_1528);
nor U1644 (N_1644,N_1566,N_1505);
nor U1645 (N_1645,N_1529,N_1575);
or U1646 (N_1646,N_1598,N_1581);
nand U1647 (N_1647,N_1553,N_1555);
nand U1648 (N_1648,N_1577,N_1544);
or U1649 (N_1649,N_1591,N_1510);
and U1650 (N_1650,N_1500,N_1580);
or U1651 (N_1651,N_1584,N_1517);
and U1652 (N_1652,N_1571,N_1577);
or U1653 (N_1653,N_1595,N_1535);
and U1654 (N_1654,N_1579,N_1563);
or U1655 (N_1655,N_1586,N_1536);
and U1656 (N_1656,N_1547,N_1509);
nor U1657 (N_1657,N_1505,N_1540);
and U1658 (N_1658,N_1574,N_1586);
xor U1659 (N_1659,N_1535,N_1554);
nor U1660 (N_1660,N_1590,N_1535);
nand U1661 (N_1661,N_1589,N_1575);
nand U1662 (N_1662,N_1540,N_1541);
nor U1663 (N_1663,N_1548,N_1577);
or U1664 (N_1664,N_1500,N_1589);
and U1665 (N_1665,N_1502,N_1504);
nor U1666 (N_1666,N_1518,N_1544);
and U1667 (N_1667,N_1526,N_1515);
and U1668 (N_1668,N_1594,N_1543);
nand U1669 (N_1669,N_1561,N_1525);
nor U1670 (N_1670,N_1582,N_1515);
nor U1671 (N_1671,N_1523,N_1583);
nor U1672 (N_1672,N_1541,N_1510);
or U1673 (N_1673,N_1589,N_1524);
xnor U1674 (N_1674,N_1519,N_1579);
xnor U1675 (N_1675,N_1502,N_1513);
xor U1676 (N_1676,N_1596,N_1503);
nand U1677 (N_1677,N_1507,N_1516);
nand U1678 (N_1678,N_1549,N_1547);
or U1679 (N_1679,N_1558,N_1560);
or U1680 (N_1680,N_1548,N_1590);
or U1681 (N_1681,N_1577,N_1507);
and U1682 (N_1682,N_1519,N_1548);
nand U1683 (N_1683,N_1575,N_1567);
nand U1684 (N_1684,N_1557,N_1561);
or U1685 (N_1685,N_1575,N_1590);
or U1686 (N_1686,N_1549,N_1552);
or U1687 (N_1687,N_1552,N_1599);
and U1688 (N_1688,N_1521,N_1592);
nor U1689 (N_1689,N_1537,N_1573);
nand U1690 (N_1690,N_1500,N_1557);
nor U1691 (N_1691,N_1544,N_1533);
xor U1692 (N_1692,N_1571,N_1560);
nor U1693 (N_1693,N_1562,N_1561);
xnor U1694 (N_1694,N_1593,N_1562);
or U1695 (N_1695,N_1538,N_1587);
or U1696 (N_1696,N_1546,N_1512);
nand U1697 (N_1697,N_1501,N_1512);
and U1698 (N_1698,N_1501,N_1537);
nand U1699 (N_1699,N_1555,N_1576);
nor U1700 (N_1700,N_1639,N_1649);
or U1701 (N_1701,N_1619,N_1674);
nand U1702 (N_1702,N_1618,N_1627);
nor U1703 (N_1703,N_1657,N_1613);
xor U1704 (N_1704,N_1615,N_1626);
or U1705 (N_1705,N_1661,N_1641);
nand U1706 (N_1706,N_1663,N_1693);
xor U1707 (N_1707,N_1608,N_1617);
xnor U1708 (N_1708,N_1685,N_1695);
and U1709 (N_1709,N_1656,N_1659);
or U1710 (N_1710,N_1612,N_1625);
nor U1711 (N_1711,N_1600,N_1680);
or U1712 (N_1712,N_1679,N_1668);
xnor U1713 (N_1713,N_1628,N_1682);
and U1714 (N_1714,N_1690,N_1632);
or U1715 (N_1715,N_1633,N_1677);
nor U1716 (N_1716,N_1647,N_1605);
nor U1717 (N_1717,N_1609,N_1684);
and U1718 (N_1718,N_1648,N_1634);
nor U1719 (N_1719,N_1614,N_1645);
and U1720 (N_1720,N_1671,N_1692);
and U1721 (N_1721,N_1642,N_1621);
nor U1722 (N_1722,N_1638,N_1616);
nand U1723 (N_1723,N_1676,N_1603);
or U1724 (N_1724,N_1691,N_1697);
xor U1725 (N_1725,N_1678,N_1654);
nand U1726 (N_1726,N_1624,N_1629);
nand U1727 (N_1727,N_1604,N_1696);
nor U1728 (N_1728,N_1673,N_1644);
nor U1729 (N_1729,N_1653,N_1687);
nand U1730 (N_1730,N_1683,N_1620);
nand U1731 (N_1731,N_1652,N_1630);
nor U1732 (N_1732,N_1646,N_1655);
and U1733 (N_1733,N_1667,N_1640);
nor U1734 (N_1734,N_1643,N_1688);
and U1735 (N_1735,N_1675,N_1601);
xor U1736 (N_1736,N_1664,N_1636);
nand U1737 (N_1737,N_1611,N_1672);
or U1738 (N_1738,N_1622,N_1681);
nand U1739 (N_1739,N_1637,N_1651);
nor U1740 (N_1740,N_1686,N_1606);
and U1741 (N_1741,N_1602,N_1660);
nor U1742 (N_1742,N_1662,N_1669);
nor U1743 (N_1743,N_1658,N_1694);
xnor U1744 (N_1744,N_1631,N_1670);
nor U1745 (N_1745,N_1665,N_1607);
nand U1746 (N_1746,N_1698,N_1650);
xnor U1747 (N_1747,N_1689,N_1635);
nor U1748 (N_1748,N_1699,N_1610);
xor U1749 (N_1749,N_1666,N_1623);
nand U1750 (N_1750,N_1616,N_1641);
xnor U1751 (N_1751,N_1607,N_1672);
nor U1752 (N_1752,N_1622,N_1668);
nand U1753 (N_1753,N_1652,N_1601);
and U1754 (N_1754,N_1696,N_1642);
nor U1755 (N_1755,N_1666,N_1631);
and U1756 (N_1756,N_1641,N_1688);
or U1757 (N_1757,N_1600,N_1619);
nand U1758 (N_1758,N_1640,N_1682);
or U1759 (N_1759,N_1646,N_1680);
and U1760 (N_1760,N_1628,N_1630);
and U1761 (N_1761,N_1676,N_1694);
or U1762 (N_1762,N_1663,N_1680);
nor U1763 (N_1763,N_1658,N_1640);
and U1764 (N_1764,N_1677,N_1690);
or U1765 (N_1765,N_1684,N_1667);
nand U1766 (N_1766,N_1624,N_1673);
or U1767 (N_1767,N_1658,N_1634);
nor U1768 (N_1768,N_1620,N_1662);
or U1769 (N_1769,N_1664,N_1625);
and U1770 (N_1770,N_1619,N_1655);
nor U1771 (N_1771,N_1664,N_1615);
and U1772 (N_1772,N_1621,N_1643);
xnor U1773 (N_1773,N_1692,N_1652);
nand U1774 (N_1774,N_1686,N_1657);
and U1775 (N_1775,N_1615,N_1643);
nor U1776 (N_1776,N_1667,N_1658);
nand U1777 (N_1777,N_1687,N_1646);
or U1778 (N_1778,N_1697,N_1656);
nor U1779 (N_1779,N_1676,N_1670);
and U1780 (N_1780,N_1627,N_1609);
and U1781 (N_1781,N_1610,N_1636);
nand U1782 (N_1782,N_1689,N_1623);
nand U1783 (N_1783,N_1695,N_1642);
and U1784 (N_1784,N_1619,N_1680);
xnor U1785 (N_1785,N_1686,N_1610);
nand U1786 (N_1786,N_1674,N_1699);
and U1787 (N_1787,N_1664,N_1680);
xor U1788 (N_1788,N_1601,N_1687);
xor U1789 (N_1789,N_1616,N_1676);
nand U1790 (N_1790,N_1696,N_1668);
nand U1791 (N_1791,N_1641,N_1691);
nor U1792 (N_1792,N_1609,N_1648);
nor U1793 (N_1793,N_1663,N_1631);
nand U1794 (N_1794,N_1625,N_1666);
and U1795 (N_1795,N_1630,N_1672);
or U1796 (N_1796,N_1652,N_1659);
and U1797 (N_1797,N_1696,N_1603);
xnor U1798 (N_1798,N_1666,N_1656);
nand U1799 (N_1799,N_1643,N_1655);
or U1800 (N_1800,N_1736,N_1784);
nor U1801 (N_1801,N_1702,N_1787);
nor U1802 (N_1802,N_1701,N_1741);
or U1803 (N_1803,N_1754,N_1788);
and U1804 (N_1804,N_1743,N_1755);
and U1805 (N_1805,N_1762,N_1785);
nand U1806 (N_1806,N_1710,N_1720);
nand U1807 (N_1807,N_1781,N_1786);
nand U1808 (N_1808,N_1727,N_1707);
xor U1809 (N_1809,N_1732,N_1798);
or U1810 (N_1810,N_1780,N_1763);
nor U1811 (N_1811,N_1721,N_1740);
or U1812 (N_1812,N_1756,N_1723);
or U1813 (N_1813,N_1733,N_1769);
nor U1814 (N_1814,N_1717,N_1779);
xnor U1815 (N_1815,N_1709,N_1716);
nor U1816 (N_1816,N_1742,N_1796);
nor U1817 (N_1817,N_1735,N_1760);
and U1818 (N_1818,N_1767,N_1739);
and U1819 (N_1819,N_1737,N_1715);
nor U1820 (N_1820,N_1750,N_1761);
and U1821 (N_1821,N_1782,N_1766);
nand U1822 (N_1822,N_1747,N_1789);
nand U1823 (N_1823,N_1745,N_1790);
and U1824 (N_1824,N_1719,N_1793);
nor U1825 (N_1825,N_1791,N_1705);
or U1826 (N_1826,N_1783,N_1775);
nand U1827 (N_1827,N_1744,N_1752);
nand U1828 (N_1828,N_1797,N_1753);
nand U1829 (N_1829,N_1748,N_1773);
or U1830 (N_1830,N_1778,N_1731);
or U1831 (N_1831,N_1749,N_1708);
xor U1832 (N_1832,N_1795,N_1724);
nor U1833 (N_1833,N_1746,N_1777);
and U1834 (N_1834,N_1722,N_1772);
or U1835 (N_1835,N_1776,N_1712);
and U1836 (N_1836,N_1758,N_1759);
or U1837 (N_1837,N_1700,N_1726);
nand U1838 (N_1838,N_1728,N_1799);
and U1839 (N_1839,N_1770,N_1734);
and U1840 (N_1840,N_1794,N_1711);
xor U1841 (N_1841,N_1729,N_1713);
nor U1842 (N_1842,N_1751,N_1706);
and U1843 (N_1843,N_1718,N_1730);
or U1844 (N_1844,N_1738,N_1714);
nor U1845 (N_1845,N_1792,N_1725);
nand U1846 (N_1846,N_1774,N_1768);
or U1847 (N_1847,N_1703,N_1764);
nor U1848 (N_1848,N_1771,N_1757);
nor U1849 (N_1849,N_1704,N_1765);
nor U1850 (N_1850,N_1749,N_1762);
nor U1851 (N_1851,N_1724,N_1768);
and U1852 (N_1852,N_1765,N_1717);
nor U1853 (N_1853,N_1725,N_1765);
or U1854 (N_1854,N_1754,N_1705);
nor U1855 (N_1855,N_1730,N_1705);
nand U1856 (N_1856,N_1738,N_1722);
nand U1857 (N_1857,N_1712,N_1750);
and U1858 (N_1858,N_1785,N_1705);
and U1859 (N_1859,N_1739,N_1748);
nor U1860 (N_1860,N_1725,N_1772);
nor U1861 (N_1861,N_1700,N_1730);
or U1862 (N_1862,N_1727,N_1748);
nand U1863 (N_1863,N_1774,N_1786);
nand U1864 (N_1864,N_1767,N_1794);
nor U1865 (N_1865,N_1706,N_1735);
nor U1866 (N_1866,N_1720,N_1746);
or U1867 (N_1867,N_1787,N_1718);
nor U1868 (N_1868,N_1760,N_1784);
nand U1869 (N_1869,N_1769,N_1717);
xnor U1870 (N_1870,N_1728,N_1756);
and U1871 (N_1871,N_1777,N_1751);
and U1872 (N_1872,N_1762,N_1716);
or U1873 (N_1873,N_1739,N_1728);
nor U1874 (N_1874,N_1782,N_1765);
and U1875 (N_1875,N_1740,N_1750);
nand U1876 (N_1876,N_1759,N_1720);
xnor U1877 (N_1877,N_1738,N_1734);
and U1878 (N_1878,N_1704,N_1701);
nor U1879 (N_1879,N_1747,N_1717);
xnor U1880 (N_1880,N_1714,N_1794);
and U1881 (N_1881,N_1743,N_1752);
xnor U1882 (N_1882,N_1779,N_1763);
nor U1883 (N_1883,N_1710,N_1780);
or U1884 (N_1884,N_1778,N_1722);
or U1885 (N_1885,N_1710,N_1740);
nor U1886 (N_1886,N_1710,N_1742);
nand U1887 (N_1887,N_1763,N_1796);
nand U1888 (N_1888,N_1750,N_1772);
nand U1889 (N_1889,N_1768,N_1762);
nand U1890 (N_1890,N_1765,N_1747);
nand U1891 (N_1891,N_1759,N_1792);
and U1892 (N_1892,N_1777,N_1793);
nand U1893 (N_1893,N_1793,N_1715);
xor U1894 (N_1894,N_1756,N_1712);
or U1895 (N_1895,N_1780,N_1772);
xor U1896 (N_1896,N_1762,N_1729);
nand U1897 (N_1897,N_1795,N_1760);
nor U1898 (N_1898,N_1732,N_1770);
and U1899 (N_1899,N_1774,N_1716);
xnor U1900 (N_1900,N_1824,N_1859);
nand U1901 (N_1901,N_1818,N_1888);
nor U1902 (N_1902,N_1803,N_1854);
nand U1903 (N_1903,N_1850,N_1840);
nand U1904 (N_1904,N_1849,N_1842);
xor U1905 (N_1905,N_1838,N_1884);
nor U1906 (N_1906,N_1841,N_1835);
nor U1907 (N_1907,N_1866,N_1817);
nand U1908 (N_1908,N_1827,N_1876);
nor U1909 (N_1909,N_1815,N_1862);
or U1910 (N_1910,N_1800,N_1808);
nand U1911 (N_1911,N_1885,N_1845);
xnor U1912 (N_1912,N_1881,N_1847);
and U1913 (N_1913,N_1853,N_1837);
xnor U1914 (N_1914,N_1836,N_1865);
or U1915 (N_1915,N_1832,N_1891);
and U1916 (N_1916,N_1898,N_1892);
nand U1917 (N_1917,N_1863,N_1813);
or U1918 (N_1918,N_1846,N_1874);
nand U1919 (N_1919,N_1860,N_1899);
nor U1920 (N_1920,N_1896,N_1820);
nand U1921 (N_1921,N_1873,N_1858);
nor U1922 (N_1922,N_1880,N_1821);
and U1923 (N_1923,N_1822,N_1816);
nand U1924 (N_1924,N_1809,N_1844);
nand U1925 (N_1925,N_1883,N_1864);
nor U1926 (N_1926,N_1856,N_1810);
nor U1927 (N_1927,N_1807,N_1855);
nor U1928 (N_1928,N_1830,N_1806);
nand U1929 (N_1929,N_1878,N_1833);
and U1930 (N_1930,N_1831,N_1895);
and U1931 (N_1931,N_1871,N_1887);
nand U1932 (N_1932,N_1805,N_1893);
and U1933 (N_1933,N_1870,N_1889);
or U1934 (N_1934,N_1843,N_1868);
and U1935 (N_1935,N_1834,N_1801);
xnor U1936 (N_1936,N_1897,N_1890);
nand U1937 (N_1937,N_1811,N_1829);
or U1938 (N_1938,N_1879,N_1857);
nand U1939 (N_1939,N_1851,N_1826);
xor U1940 (N_1940,N_1804,N_1839);
nor U1941 (N_1941,N_1812,N_1825);
xor U1942 (N_1942,N_1869,N_1875);
nand U1943 (N_1943,N_1867,N_1823);
xor U1944 (N_1944,N_1852,N_1848);
or U1945 (N_1945,N_1814,N_1802);
or U1946 (N_1946,N_1872,N_1894);
nor U1947 (N_1947,N_1819,N_1861);
nand U1948 (N_1948,N_1877,N_1886);
or U1949 (N_1949,N_1882,N_1828);
nand U1950 (N_1950,N_1878,N_1844);
and U1951 (N_1951,N_1803,N_1851);
and U1952 (N_1952,N_1813,N_1837);
and U1953 (N_1953,N_1817,N_1828);
or U1954 (N_1954,N_1881,N_1811);
or U1955 (N_1955,N_1855,N_1890);
nor U1956 (N_1956,N_1800,N_1882);
nand U1957 (N_1957,N_1848,N_1893);
xnor U1958 (N_1958,N_1818,N_1851);
and U1959 (N_1959,N_1855,N_1819);
or U1960 (N_1960,N_1825,N_1831);
or U1961 (N_1961,N_1828,N_1841);
and U1962 (N_1962,N_1851,N_1888);
nor U1963 (N_1963,N_1898,N_1844);
nor U1964 (N_1964,N_1889,N_1830);
nor U1965 (N_1965,N_1845,N_1880);
nor U1966 (N_1966,N_1848,N_1831);
nor U1967 (N_1967,N_1885,N_1888);
xor U1968 (N_1968,N_1830,N_1841);
and U1969 (N_1969,N_1880,N_1852);
and U1970 (N_1970,N_1865,N_1852);
or U1971 (N_1971,N_1819,N_1849);
and U1972 (N_1972,N_1853,N_1818);
nor U1973 (N_1973,N_1820,N_1802);
xnor U1974 (N_1974,N_1873,N_1814);
nand U1975 (N_1975,N_1865,N_1849);
xor U1976 (N_1976,N_1823,N_1897);
nor U1977 (N_1977,N_1849,N_1870);
and U1978 (N_1978,N_1837,N_1880);
and U1979 (N_1979,N_1866,N_1894);
xnor U1980 (N_1980,N_1858,N_1854);
or U1981 (N_1981,N_1808,N_1877);
nor U1982 (N_1982,N_1867,N_1881);
nor U1983 (N_1983,N_1877,N_1873);
and U1984 (N_1984,N_1893,N_1865);
nor U1985 (N_1985,N_1880,N_1888);
or U1986 (N_1986,N_1802,N_1881);
and U1987 (N_1987,N_1849,N_1807);
xnor U1988 (N_1988,N_1847,N_1848);
nor U1989 (N_1989,N_1811,N_1841);
nor U1990 (N_1990,N_1858,N_1849);
and U1991 (N_1991,N_1863,N_1829);
nor U1992 (N_1992,N_1833,N_1847);
and U1993 (N_1993,N_1872,N_1822);
xnor U1994 (N_1994,N_1811,N_1868);
and U1995 (N_1995,N_1830,N_1839);
xnor U1996 (N_1996,N_1843,N_1813);
and U1997 (N_1997,N_1853,N_1891);
nand U1998 (N_1998,N_1878,N_1811);
or U1999 (N_1999,N_1845,N_1820);
nand U2000 (N_2000,N_1993,N_1938);
and U2001 (N_2001,N_1930,N_1990);
nor U2002 (N_2002,N_1961,N_1954);
nand U2003 (N_2003,N_1939,N_1959);
and U2004 (N_2004,N_1900,N_1980);
or U2005 (N_2005,N_1964,N_1932);
nand U2006 (N_2006,N_1913,N_1920);
nand U2007 (N_2007,N_1955,N_1902);
and U2008 (N_2008,N_1921,N_1986);
nand U2009 (N_2009,N_1916,N_1962);
xnor U2010 (N_2010,N_1994,N_1998);
nand U2011 (N_2011,N_1969,N_1935);
or U2012 (N_2012,N_1989,N_1903);
or U2013 (N_2013,N_1905,N_1950);
xor U2014 (N_2014,N_1929,N_1915);
nand U2015 (N_2015,N_1983,N_1946);
nand U2016 (N_2016,N_1909,N_1928);
xor U2017 (N_2017,N_1918,N_1901);
and U2018 (N_2018,N_1960,N_1925);
nand U2019 (N_2019,N_1988,N_1923);
nor U2020 (N_2020,N_1984,N_1976);
nand U2021 (N_2021,N_1977,N_1947);
nand U2022 (N_2022,N_1924,N_1943);
nor U2023 (N_2023,N_1934,N_1992);
and U2024 (N_2024,N_1979,N_1968);
nand U2025 (N_2025,N_1996,N_1974);
or U2026 (N_2026,N_1957,N_1963);
nor U2027 (N_2027,N_1911,N_1914);
nor U2028 (N_2028,N_1919,N_1985);
nor U2029 (N_2029,N_1978,N_1926);
xnor U2030 (N_2030,N_1970,N_1908);
and U2031 (N_2031,N_1912,N_1942);
and U2032 (N_2032,N_1966,N_1907);
or U2033 (N_2033,N_1981,N_1949);
nand U2034 (N_2034,N_1967,N_1944);
nand U2035 (N_2035,N_1975,N_1999);
or U2036 (N_2036,N_1997,N_1995);
nor U2037 (N_2037,N_1948,N_1973);
or U2038 (N_2038,N_1945,N_1956);
and U2039 (N_2039,N_1910,N_1952);
or U2040 (N_2040,N_1971,N_1931);
and U2041 (N_2041,N_1917,N_1953);
nand U2042 (N_2042,N_1987,N_1927);
or U2043 (N_2043,N_1936,N_1958);
nor U2044 (N_2044,N_1940,N_1951);
or U2045 (N_2045,N_1982,N_1991);
or U2046 (N_2046,N_1941,N_1965);
and U2047 (N_2047,N_1933,N_1904);
and U2048 (N_2048,N_1937,N_1922);
or U2049 (N_2049,N_1906,N_1972);
xnor U2050 (N_2050,N_1962,N_1914);
xnor U2051 (N_2051,N_1947,N_1907);
nor U2052 (N_2052,N_1948,N_1982);
nand U2053 (N_2053,N_1916,N_1930);
or U2054 (N_2054,N_1916,N_1988);
and U2055 (N_2055,N_1977,N_1955);
xor U2056 (N_2056,N_1901,N_1925);
nand U2057 (N_2057,N_1981,N_1956);
and U2058 (N_2058,N_1976,N_1983);
nand U2059 (N_2059,N_1981,N_1947);
xor U2060 (N_2060,N_1971,N_1935);
nor U2061 (N_2061,N_1990,N_1976);
nand U2062 (N_2062,N_1945,N_1905);
or U2063 (N_2063,N_1969,N_1981);
nor U2064 (N_2064,N_1908,N_1916);
nor U2065 (N_2065,N_1904,N_1911);
nand U2066 (N_2066,N_1930,N_1951);
nand U2067 (N_2067,N_1939,N_1946);
nor U2068 (N_2068,N_1993,N_1971);
or U2069 (N_2069,N_1956,N_1984);
xnor U2070 (N_2070,N_1903,N_1988);
and U2071 (N_2071,N_1939,N_1981);
xnor U2072 (N_2072,N_1971,N_1952);
nand U2073 (N_2073,N_1960,N_1931);
xnor U2074 (N_2074,N_1984,N_1916);
or U2075 (N_2075,N_1937,N_1935);
or U2076 (N_2076,N_1924,N_1963);
nand U2077 (N_2077,N_1936,N_1915);
and U2078 (N_2078,N_1940,N_1978);
nor U2079 (N_2079,N_1953,N_1924);
nor U2080 (N_2080,N_1914,N_1988);
nor U2081 (N_2081,N_1995,N_1991);
nor U2082 (N_2082,N_1955,N_1914);
nor U2083 (N_2083,N_1996,N_1927);
xor U2084 (N_2084,N_1931,N_1983);
xnor U2085 (N_2085,N_1909,N_1977);
or U2086 (N_2086,N_1984,N_1906);
and U2087 (N_2087,N_1980,N_1963);
nor U2088 (N_2088,N_1982,N_1972);
xor U2089 (N_2089,N_1944,N_1905);
xnor U2090 (N_2090,N_1977,N_1933);
and U2091 (N_2091,N_1997,N_1918);
or U2092 (N_2092,N_1986,N_1968);
and U2093 (N_2093,N_1948,N_1957);
nor U2094 (N_2094,N_1929,N_1912);
and U2095 (N_2095,N_1902,N_1923);
and U2096 (N_2096,N_1920,N_1969);
or U2097 (N_2097,N_1902,N_1938);
or U2098 (N_2098,N_1934,N_1965);
or U2099 (N_2099,N_1938,N_1919);
and U2100 (N_2100,N_2057,N_2061);
and U2101 (N_2101,N_2077,N_2099);
and U2102 (N_2102,N_2032,N_2037);
nor U2103 (N_2103,N_2081,N_2068);
xnor U2104 (N_2104,N_2059,N_2074);
and U2105 (N_2105,N_2097,N_2044);
xor U2106 (N_2106,N_2018,N_2058);
nand U2107 (N_2107,N_2019,N_2086);
nand U2108 (N_2108,N_2041,N_2045);
and U2109 (N_2109,N_2003,N_2043);
nand U2110 (N_2110,N_2051,N_2023);
nor U2111 (N_2111,N_2072,N_2017);
and U2112 (N_2112,N_2076,N_2080);
nand U2113 (N_2113,N_2012,N_2033);
and U2114 (N_2114,N_2079,N_2049);
and U2115 (N_2115,N_2010,N_2065);
or U2116 (N_2116,N_2093,N_2070);
nor U2117 (N_2117,N_2098,N_2024);
or U2118 (N_2118,N_2016,N_2020);
or U2119 (N_2119,N_2091,N_2052);
nor U2120 (N_2120,N_2053,N_2007);
or U2121 (N_2121,N_2083,N_2015);
nor U2122 (N_2122,N_2004,N_2002);
nor U2123 (N_2123,N_2034,N_2094);
nor U2124 (N_2124,N_2001,N_2066);
or U2125 (N_2125,N_2048,N_2089);
and U2126 (N_2126,N_2039,N_2087);
and U2127 (N_2127,N_2090,N_2055);
nand U2128 (N_2128,N_2008,N_2067);
nor U2129 (N_2129,N_2042,N_2096);
nor U2130 (N_2130,N_2028,N_2047);
nand U2131 (N_2131,N_2084,N_2062);
or U2132 (N_2132,N_2056,N_2035);
or U2133 (N_2133,N_2085,N_2046);
xor U2134 (N_2134,N_2013,N_2014);
nand U2135 (N_2135,N_2026,N_2060);
or U2136 (N_2136,N_2029,N_2000);
and U2137 (N_2137,N_2064,N_2082);
and U2138 (N_2138,N_2073,N_2036);
xnor U2139 (N_2139,N_2092,N_2040);
or U2140 (N_2140,N_2038,N_2011);
nand U2141 (N_2141,N_2069,N_2005);
or U2142 (N_2142,N_2030,N_2009);
xor U2143 (N_2143,N_2027,N_2006);
nand U2144 (N_2144,N_2050,N_2088);
or U2145 (N_2145,N_2025,N_2075);
nor U2146 (N_2146,N_2078,N_2022);
nand U2147 (N_2147,N_2071,N_2021);
nand U2148 (N_2148,N_2054,N_2031);
nand U2149 (N_2149,N_2095,N_2063);
or U2150 (N_2150,N_2053,N_2049);
nor U2151 (N_2151,N_2006,N_2072);
nand U2152 (N_2152,N_2053,N_2010);
nor U2153 (N_2153,N_2046,N_2006);
nor U2154 (N_2154,N_2050,N_2060);
and U2155 (N_2155,N_2001,N_2046);
and U2156 (N_2156,N_2008,N_2072);
nor U2157 (N_2157,N_2048,N_2054);
nand U2158 (N_2158,N_2029,N_2007);
and U2159 (N_2159,N_2069,N_2031);
nor U2160 (N_2160,N_2014,N_2046);
nand U2161 (N_2161,N_2044,N_2085);
or U2162 (N_2162,N_2056,N_2007);
and U2163 (N_2163,N_2032,N_2050);
nor U2164 (N_2164,N_2066,N_2008);
and U2165 (N_2165,N_2029,N_2017);
nand U2166 (N_2166,N_2021,N_2001);
and U2167 (N_2167,N_2069,N_2000);
and U2168 (N_2168,N_2066,N_2073);
and U2169 (N_2169,N_2048,N_2043);
or U2170 (N_2170,N_2061,N_2081);
nand U2171 (N_2171,N_2009,N_2060);
and U2172 (N_2172,N_2063,N_2046);
or U2173 (N_2173,N_2028,N_2053);
and U2174 (N_2174,N_2006,N_2034);
nand U2175 (N_2175,N_2004,N_2092);
or U2176 (N_2176,N_2032,N_2063);
and U2177 (N_2177,N_2091,N_2086);
nand U2178 (N_2178,N_2098,N_2043);
nor U2179 (N_2179,N_2090,N_2012);
nand U2180 (N_2180,N_2005,N_2020);
xnor U2181 (N_2181,N_2022,N_2073);
and U2182 (N_2182,N_2095,N_2006);
or U2183 (N_2183,N_2086,N_2017);
and U2184 (N_2184,N_2040,N_2003);
and U2185 (N_2185,N_2094,N_2028);
nor U2186 (N_2186,N_2018,N_2053);
and U2187 (N_2187,N_2036,N_2097);
and U2188 (N_2188,N_2054,N_2027);
xnor U2189 (N_2189,N_2051,N_2044);
nor U2190 (N_2190,N_2087,N_2071);
or U2191 (N_2191,N_2083,N_2001);
and U2192 (N_2192,N_2061,N_2068);
nand U2193 (N_2193,N_2066,N_2081);
and U2194 (N_2194,N_2093,N_2072);
and U2195 (N_2195,N_2057,N_2092);
or U2196 (N_2196,N_2067,N_2025);
nor U2197 (N_2197,N_2078,N_2049);
xnor U2198 (N_2198,N_2006,N_2084);
nor U2199 (N_2199,N_2076,N_2007);
nor U2200 (N_2200,N_2114,N_2180);
nor U2201 (N_2201,N_2148,N_2199);
nand U2202 (N_2202,N_2176,N_2166);
nand U2203 (N_2203,N_2163,N_2121);
nor U2204 (N_2204,N_2184,N_2137);
nor U2205 (N_2205,N_2157,N_2123);
nor U2206 (N_2206,N_2143,N_2187);
or U2207 (N_2207,N_2146,N_2191);
or U2208 (N_2208,N_2102,N_2153);
and U2209 (N_2209,N_2150,N_2134);
nor U2210 (N_2210,N_2152,N_2129);
nand U2211 (N_2211,N_2155,N_2109);
or U2212 (N_2212,N_2124,N_2169);
and U2213 (N_2213,N_2179,N_2131);
nand U2214 (N_2214,N_2172,N_2167);
nor U2215 (N_2215,N_2151,N_2162);
and U2216 (N_2216,N_2110,N_2108);
nand U2217 (N_2217,N_2107,N_2178);
or U2218 (N_2218,N_2156,N_2103);
and U2219 (N_2219,N_2173,N_2174);
or U2220 (N_2220,N_2115,N_2100);
and U2221 (N_2221,N_2111,N_2125);
nor U2222 (N_2222,N_2168,N_2101);
and U2223 (N_2223,N_2164,N_2112);
nor U2224 (N_2224,N_2127,N_2133);
and U2225 (N_2225,N_2198,N_2185);
nor U2226 (N_2226,N_2106,N_2175);
or U2227 (N_2227,N_2141,N_2117);
nor U2228 (N_2228,N_2139,N_2189);
nor U2229 (N_2229,N_2188,N_2116);
or U2230 (N_2230,N_2149,N_2195);
and U2231 (N_2231,N_2140,N_2138);
and U2232 (N_2232,N_2122,N_2160);
or U2233 (N_2233,N_2171,N_2130);
nand U2234 (N_2234,N_2170,N_2158);
nor U2235 (N_2235,N_2192,N_2136);
nand U2236 (N_2236,N_2193,N_2120);
xnor U2237 (N_2237,N_2132,N_2119);
and U2238 (N_2238,N_2135,N_2154);
nand U2239 (N_2239,N_2104,N_2147);
xnor U2240 (N_2240,N_2177,N_2118);
or U2241 (N_2241,N_2142,N_2105);
or U2242 (N_2242,N_2159,N_2190);
and U2243 (N_2243,N_2183,N_2197);
and U2244 (N_2244,N_2181,N_2126);
or U2245 (N_2245,N_2145,N_2194);
nand U2246 (N_2246,N_2165,N_2196);
or U2247 (N_2247,N_2186,N_2161);
and U2248 (N_2248,N_2182,N_2144);
or U2249 (N_2249,N_2128,N_2113);
nand U2250 (N_2250,N_2162,N_2166);
nor U2251 (N_2251,N_2123,N_2199);
nor U2252 (N_2252,N_2112,N_2131);
nor U2253 (N_2253,N_2189,N_2130);
or U2254 (N_2254,N_2193,N_2164);
nand U2255 (N_2255,N_2188,N_2131);
nor U2256 (N_2256,N_2199,N_2164);
nor U2257 (N_2257,N_2103,N_2163);
and U2258 (N_2258,N_2109,N_2193);
or U2259 (N_2259,N_2133,N_2195);
and U2260 (N_2260,N_2148,N_2160);
xnor U2261 (N_2261,N_2142,N_2187);
nand U2262 (N_2262,N_2189,N_2137);
and U2263 (N_2263,N_2149,N_2165);
or U2264 (N_2264,N_2166,N_2106);
nand U2265 (N_2265,N_2168,N_2165);
and U2266 (N_2266,N_2104,N_2131);
nand U2267 (N_2267,N_2122,N_2123);
and U2268 (N_2268,N_2192,N_2133);
nand U2269 (N_2269,N_2153,N_2104);
and U2270 (N_2270,N_2160,N_2107);
nor U2271 (N_2271,N_2129,N_2133);
nor U2272 (N_2272,N_2146,N_2117);
xnor U2273 (N_2273,N_2150,N_2140);
or U2274 (N_2274,N_2100,N_2127);
nor U2275 (N_2275,N_2100,N_2181);
nor U2276 (N_2276,N_2172,N_2155);
or U2277 (N_2277,N_2133,N_2140);
nand U2278 (N_2278,N_2173,N_2117);
and U2279 (N_2279,N_2157,N_2144);
and U2280 (N_2280,N_2109,N_2163);
and U2281 (N_2281,N_2155,N_2178);
nand U2282 (N_2282,N_2192,N_2149);
nand U2283 (N_2283,N_2190,N_2145);
or U2284 (N_2284,N_2172,N_2146);
nand U2285 (N_2285,N_2102,N_2185);
nor U2286 (N_2286,N_2113,N_2167);
nor U2287 (N_2287,N_2134,N_2107);
nor U2288 (N_2288,N_2142,N_2160);
nand U2289 (N_2289,N_2152,N_2145);
xor U2290 (N_2290,N_2134,N_2157);
nand U2291 (N_2291,N_2151,N_2137);
xnor U2292 (N_2292,N_2138,N_2102);
nor U2293 (N_2293,N_2174,N_2181);
nand U2294 (N_2294,N_2197,N_2166);
or U2295 (N_2295,N_2162,N_2126);
nand U2296 (N_2296,N_2199,N_2165);
and U2297 (N_2297,N_2176,N_2153);
nand U2298 (N_2298,N_2105,N_2123);
nand U2299 (N_2299,N_2115,N_2185);
xor U2300 (N_2300,N_2297,N_2211);
xnor U2301 (N_2301,N_2281,N_2229);
and U2302 (N_2302,N_2215,N_2238);
nand U2303 (N_2303,N_2254,N_2296);
nand U2304 (N_2304,N_2280,N_2240);
nor U2305 (N_2305,N_2214,N_2282);
and U2306 (N_2306,N_2201,N_2255);
xnor U2307 (N_2307,N_2250,N_2248);
or U2308 (N_2308,N_2251,N_2206);
and U2309 (N_2309,N_2217,N_2290);
nor U2310 (N_2310,N_2204,N_2253);
or U2311 (N_2311,N_2295,N_2224);
and U2312 (N_2312,N_2291,N_2221);
nand U2313 (N_2313,N_2261,N_2269);
and U2314 (N_2314,N_2228,N_2230);
and U2315 (N_2315,N_2278,N_2267);
and U2316 (N_2316,N_2239,N_2292);
nand U2317 (N_2317,N_2213,N_2294);
nand U2318 (N_2318,N_2232,N_2271);
nor U2319 (N_2319,N_2283,N_2209);
nand U2320 (N_2320,N_2262,N_2244);
or U2321 (N_2321,N_2298,N_2243);
nand U2322 (N_2322,N_2222,N_2279);
nor U2323 (N_2323,N_2235,N_2287);
nand U2324 (N_2324,N_2207,N_2225);
and U2325 (N_2325,N_2219,N_2299);
and U2326 (N_2326,N_2241,N_2263);
or U2327 (N_2327,N_2202,N_2285);
or U2328 (N_2328,N_2276,N_2245);
nor U2329 (N_2329,N_2210,N_2272);
or U2330 (N_2330,N_2275,N_2226);
nor U2331 (N_2331,N_2247,N_2212);
and U2332 (N_2332,N_2268,N_2258);
nor U2333 (N_2333,N_2227,N_2256);
nor U2334 (N_2334,N_2289,N_2265);
or U2335 (N_2335,N_2237,N_2249);
and U2336 (N_2336,N_2284,N_2231);
nor U2337 (N_2337,N_2270,N_2260);
and U2338 (N_2338,N_2233,N_2259);
or U2339 (N_2339,N_2218,N_2257);
or U2340 (N_2340,N_2252,N_2277);
nand U2341 (N_2341,N_2234,N_2208);
or U2342 (N_2342,N_2236,N_2216);
nor U2343 (N_2343,N_2203,N_2264);
and U2344 (N_2344,N_2246,N_2286);
or U2345 (N_2345,N_2205,N_2200);
or U2346 (N_2346,N_2242,N_2274);
or U2347 (N_2347,N_2273,N_2220);
and U2348 (N_2348,N_2288,N_2266);
nor U2349 (N_2349,N_2223,N_2293);
nor U2350 (N_2350,N_2270,N_2247);
nor U2351 (N_2351,N_2215,N_2229);
xnor U2352 (N_2352,N_2277,N_2273);
nor U2353 (N_2353,N_2257,N_2222);
or U2354 (N_2354,N_2209,N_2233);
or U2355 (N_2355,N_2237,N_2201);
and U2356 (N_2356,N_2200,N_2234);
nand U2357 (N_2357,N_2219,N_2248);
nand U2358 (N_2358,N_2247,N_2228);
nor U2359 (N_2359,N_2296,N_2284);
nor U2360 (N_2360,N_2269,N_2234);
and U2361 (N_2361,N_2286,N_2276);
or U2362 (N_2362,N_2248,N_2227);
nand U2363 (N_2363,N_2234,N_2264);
and U2364 (N_2364,N_2200,N_2288);
and U2365 (N_2365,N_2265,N_2232);
nand U2366 (N_2366,N_2294,N_2244);
nand U2367 (N_2367,N_2223,N_2292);
nand U2368 (N_2368,N_2251,N_2212);
nor U2369 (N_2369,N_2292,N_2295);
and U2370 (N_2370,N_2234,N_2282);
and U2371 (N_2371,N_2232,N_2297);
and U2372 (N_2372,N_2293,N_2249);
or U2373 (N_2373,N_2200,N_2287);
xnor U2374 (N_2374,N_2270,N_2213);
or U2375 (N_2375,N_2205,N_2273);
or U2376 (N_2376,N_2259,N_2208);
nand U2377 (N_2377,N_2276,N_2242);
nand U2378 (N_2378,N_2219,N_2202);
or U2379 (N_2379,N_2215,N_2222);
or U2380 (N_2380,N_2255,N_2248);
or U2381 (N_2381,N_2229,N_2279);
and U2382 (N_2382,N_2264,N_2274);
nor U2383 (N_2383,N_2244,N_2248);
xnor U2384 (N_2384,N_2292,N_2250);
nor U2385 (N_2385,N_2241,N_2249);
nor U2386 (N_2386,N_2297,N_2204);
nor U2387 (N_2387,N_2260,N_2266);
nand U2388 (N_2388,N_2270,N_2274);
and U2389 (N_2389,N_2229,N_2205);
nand U2390 (N_2390,N_2267,N_2241);
nand U2391 (N_2391,N_2224,N_2201);
nand U2392 (N_2392,N_2287,N_2282);
or U2393 (N_2393,N_2237,N_2215);
nand U2394 (N_2394,N_2258,N_2273);
nor U2395 (N_2395,N_2200,N_2259);
nand U2396 (N_2396,N_2224,N_2267);
and U2397 (N_2397,N_2274,N_2200);
nand U2398 (N_2398,N_2261,N_2295);
and U2399 (N_2399,N_2254,N_2278);
and U2400 (N_2400,N_2361,N_2374);
nor U2401 (N_2401,N_2331,N_2345);
nand U2402 (N_2402,N_2307,N_2390);
nor U2403 (N_2403,N_2311,N_2308);
nor U2404 (N_2404,N_2342,N_2366);
and U2405 (N_2405,N_2339,N_2363);
and U2406 (N_2406,N_2322,N_2320);
or U2407 (N_2407,N_2337,N_2319);
nor U2408 (N_2408,N_2351,N_2312);
xnor U2409 (N_2409,N_2383,N_2303);
or U2410 (N_2410,N_2326,N_2385);
or U2411 (N_2411,N_2382,N_2356);
and U2412 (N_2412,N_2340,N_2394);
and U2413 (N_2413,N_2358,N_2341);
and U2414 (N_2414,N_2355,N_2344);
and U2415 (N_2415,N_2372,N_2349);
nand U2416 (N_2416,N_2364,N_2397);
nor U2417 (N_2417,N_2368,N_2388);
and U2418 (N_2418,N_2353,N_2310);
xnor U2419 (N_2419,N_2317,N_2362);
nor U2420 (N_2420,N_2314,N_2332);
or U2421 (N_2421,N_2305,N_2348);
nor U2422 (N_2422,N_2334,N_2371);
and U2423 (N_2423,N_2313,N_2395);
nor U2424 (N_2424,N_2323,N_2376);
and U2425 (N_2425,N_2398,N_2389);
or U2426 (N_2426,N_2352,N_2346);
or U2427 (N_2427,N_2391,N_2301);
and U2428 (N_2428,N_2359,N_2316);
and U2429 (N_2429,N_2321,N_2399);
or U2430 (N_2430,N_2318,N_2375);
nand U2431 (N_2431,N_2328,N_2360);
and U2432 (N_2432,N_2327,N_2336);
nand U2433 (N_2433,N_2350,N_2300);
and U2434 (N_2434,N_2325,N_2302);
nor U2435 (N_2435,N_2330,N_2338);
or U2436 (N_2436,N_2333,N_2324);
nor U2437 (N_2437,N_2315,N_2306);
or U2438 (N_2438,N_2393,N_2354);
and U2439 (N_2439,N_2387,N_2335);
and U2440 (N_2440,N_2370,N_2309);
xor U2441 (N_2441,N_2367,N_2396);
nand U2442 (N_2442,N_2365,N_2392);
xor U2443 (N_2443,N_2381,N_2380);
and U2444 (N_2444,N_2386,N_2304);
nor U2445 (N_2445,N_2384,N_2329);
xnor U2446 (N_2446,N_2347,N_2377);
nor U2447 (N_2447,N_2343,N_2369);
and U2448 (N_2448,N_2373,N_2357);
nand U2449 (N_2449,N_2379,N_2378);
or U2450 (N_2450,N_2310,N_2394);
or U2451 (N_2451,N_2387,N_2311);
and U2452 (N_2452,N_2388,N_2336);
nand U2453 (N_2453,N_2317,N_2347);
nor U2454 (N_2454,N_2318,N_2377);
nor U2455 (N_2455,N_2314,N_2396);
and U2456 (N_2456,N_2315,N_2319);
nand U2457 (N_2457,N_2372,N_2320);
nand U2458 (N_2458,N_2371,N_2367);
or U2459 (N_2459,N_2382,N_2371);
xnor U2460 (N_2460,N_2371,N_2325);
nor U2461 (N_2461,N_2386,N_2381);
nor U2462 (N_2462,N_2319,N_2386);
or U2463 (N_2463,N_2389,N_2372);
xor U2464 (N_2464,N_2343,N_2386);
nor U2465 (N_2465,N_2368,N_2338);
nor U2466 (N_2466,N_2327,N_2342);
nand U2467 (N_2467,N_2374,N_2363);
or U2468 (N_2468,N_2365,N_2303);
xor U2469 (N_2469,N_2353,N_2360);
nor U2470 (N_2470,N_2384,N_2314);
and U2471 (N_2471,N_2348,N_2318);
nand U2472 (N_2472,N_2317,N_2321);
xnor U2473 (N_2473,N_2312,N_2336);
nand U2474 (N_2474,N_2376,N_2349);
nor U2475 (N_2475,N_2319,N_2335);
nand U2476 (N_2476,N_2308,N_2361);
and U2477 (N_2477,N_2345,N_2359);
or U2478 (N_2478,N_2308,N_2309);
or U2479 (N_2479,N_2337,N_2338);
or U2480 (N_2480,N_2377,N_2395);
nand U2481 (N_2481,N_2348,N_2391);
or U2482 (N_2482,N_2372,N_2318);
and U2483 (N_2483,N_2377,N_2328);
nand U2484 (N_2484,N_2334,N_2374);
nor U2485 (N_2485,N_2380,N_2384);
or U2486 (N_2486,N_2396,N_2347);
nor U2487 (N_2487,N_2364,N_2357);
or U2488 (N_2488,N_2307,N_2319);
nand U2489 (N_2489,N_2359,N_2342);
and U2490 (N_2490,N_2334,N_2338);
nand U2491 (N_2491,N_2394,N_2354);
xnor U2492 (N_2492,N_2318,N_2330);
nand U2493 (N_2493,N_2374,N_2308);
nor U2494 (N_2494,N_2333,N_2347);
or U2495 (N_2495,N_2332,N_2383);
nor U2496 (N_2496,N_2347,N_2341);
and U2497 (N_2497,N_2353,N_2339);
or U2498 (N_2498,N_2332,N_2392);
or U2499 (N_2499,N_2358,N_2380);
and U2500 (N_2500,N_2481,N_2483);
xor U2501 (N_2501,N_2407,N_2419);
nor U2502 (N_2502,N_2441,N_2404);
or U2503 (N_2503,N_2431,N_2424);
xor U2504 (N_2504,N_2405,N_2468);
xor U2505 (N_2505,N_2463,N_2421);
or U2506 (N_2506,N_2418,N_2489);
and U2507 (N_2507,N_2408,N_2477);
nand U2508 (N_2508,N_2471,N_2479);
and U2509 (N_2509,N_2432,N_2485);
and U2510 (N_2510,N_2449,N_2437);
and U2511 (N_2511,N_2497,N_2434);
and U2512 (N_2512,N_2425,N_2484);
and U2513 (N_2513,N_2415,N_2448);
nand U2514 (N_2514,N_2402,N_2487);
and U2515 (N_2515,N_2416,N_2410);
or U2516 (N_2516,N_2457,N_2451);
nand U2517 (N_2517,N_2495,N_2429);
and U2518 (N_2518,N_2488,N_2423);
and U2519 (N_2519,N_2470,N_2450);
and U2520 (N_2520,N_2406,N_2465);
xnor U2521 (N_2521,N_2435,N_2433);
xnor U2522 (N_2522,N_2454,N_2460);
nor U2523 (N_2523,N_2440,N_2459);
xor U2524 (N_2524,N_2486,N_2494);
and U2525 (N_2525,N_2469,N_2438);
or U2526 (N_2526,N_2475,N_2401);
and U2527 (N_2527,N_2420,N_2467);
nor U2528 (N_2528,N_2473,N_2456);
and U2529 (N_2529,N_2409,N_2400);
xor U2530 (N_2530,N_2492,N_2474);
nand U2531 (N_2531,N_2462,N_2453);
nor U2532 (N_2532,N_2427,N_2452);
nor U2533 (N_2533,N_2458,N_2478);
and U2534 (N_2534,N_2455,N_2490);
and U2535 (N_2535,N_2466,N_2439);
nand U2536 (N_2536,N_2428,N_2443);
and U2537 (N_2537,N_2417,N_2413);
nor U2538 (N_2538,N_2426,N_2464);
nand U2539 (N_2539,N_2499,N_2491);
nor U2540 (N_2540,N_2422,N_2480);
nand U2541 (N_2541,N_2442,N_2482);
or U2542 (N_2542,N_2436,N_2496);
nand U2543 (N_2543,N_2447,N_2476);
and U2544 (N_2544,N_2430,N_2461);
or U2545 (N_2545,N_2414,N_2472);
or U2546 (N_2546,N_2445,N_2498);
nand U2547 (N_2547,N_2411,N_2493);
and U2548 (N_2548,N_2403,N_2444);
and U2549 (N_2549,N_2446,N_2412);
or U2550 (N_2550,N_2481,N_2469);
nor U2551 (N_2551,N_2410,N_2474);
and U2552 (N_2552,N_2459,N_2426);
nor U2553 (N_2553,N_2410,N_2413);
nand U2554 (N_2554,N_2407,N_2497);
nor U2555 (N_2555,N_2429,N_2472);
and U2556 (N_2556,N_2485,N_2466);
nand U2557 (N_2557,N_2496,N_2417);
nor U2558 (N_2558,N_2474,N_2434);
nor U2559 (N_2559,N_2481,N_2407);
and U2560 (N_2560,N_2493,N_2485);
nand U2561 (N_2561,N_2430,N_2415);
nor U2562 (N_2562,N_2424,N_2447);
nand U2563 (N_2563,N_2462,N_2444);
nor U2564 (N_2564,N_2436,N_2405);
xor U2565 (N_2565,N_2462,N_2450);
nand U2566 (N_2566,N_2487,N_2480);
nor U2567 (N_2567,N_2424,N_2446);
nor U2568 (N_2568,N_2440,N_2407);
xor U2569 (N_2569,N_2426,N_2429);
nor U2570 (N_2570,N_2416,N_2456);
nor U2571 (N_2571,N_2471,N_2429);
nor U2572 (N_2572,N_2433,N_2440);
nor U2573 (N_2573,N_2412,N_2450);
or U2574 (N_2574,N_2458,N_2493);
or U2575 (N_2575,N_2419,N_2463);
xor U2576 (N_2576,N_2421,N_2432);
and U2577 (N_2577,N_2452,N_2450);
nand U2578 (N_2578,N_2422,N_2408);
xnor U2579 (N_2579,N_2436,N_2464);
or U2580 (N_2580,N_2496,N_2470);
nor U2581 (N_2581,N_2497,N_2465);
or U2582 (N_2582,N_2483,N_2443);
and U2583 (N_2583,N_2401,N_2402);
nand U2584 (N_2584,N_2467,N_2427);
and U2585 (N_2585,N_2477,N_2436);
nor U2586 (N_2586,N_2447,N_2415);
nor U2587 (N_2587,N_2423,N_2462);
or U2588 (N_2588,N_2444,N_2472);
xnor U2589 (N_2589,N_2485,N_2486);
and U2590 (N_2590,N_2447,N_2440);
nand U2591 (N_2591,N_2419,N_2467);
nor U2592 (N_2592,N_2400,N_2453);
or U2593 (N_2593,N_2431,N_2450);
or U2594 (N_2594,N_2420,N_2469);
or U2595 (N_2595,N_2485,N_2469);
nand U2596 (N_2596,N_2403,N_2417);
xor U2597 (N_2597,N_2419,N_2461);
nand U2598 (N_2598,N_2411,N_2498);
nand U2599 (N_2599,N_2452,N_2472);
or U2600 (N_2600,N_2572,N_2547);
nand U2601 (N_2601,N_2581,N_2577);
and U2602 (N_2602,N_2576,N_2511);
and U2603 (N_2603,N_2554,N_2550);
nor U2604 (N_2604,N_2525,N_2557);
and U2605 (N_2605,N_2519,N_2549);
nand U2606 (N_2606,N_2575,N_2535);
or U2607 (N_2607,N_2558,N_2500);
nand U2608 (N_2608,N_2521,N_2561);
nand U2609 (N_2609,N_2545,N_2586);
nand U2610 (N_2610,N_2582,N_2593);
or U2611 (N_2611,N_2506,N_2569);
nand U2612 (N_2612,N_2513,N_2508);
xnor U2613 (N_2613,N_2505,N_2515);
xnor U2614 (N_2614,N_2542,N_2523);
or U2615 (N_2615,N_2592,N_2534);
or U2616 (N_2616,N_2579,N_2590);
and U2617 (N_2617,N_2585,N_2531);
and U2618 (N_2618,N_2552,N_2502);
and U2619 (N_2619,N_2539,N_2504);
xor U2620 (N_2620,N_2571,N_2530);
nand U2621 (N_2621,N_2587,N_2536);
xnor U2622 (N_2622,N_2599,N_2598);
nor U2623 (N_2623,N_2516,N_2520);
nor U2624 (N_2624,N_2533,N_2594);
xor U2625 (N_2625,N_2589,N_2565);
xor U2626 (N_2626,N_2597,N_2596);
nor U2627 (N_2627,N_2566,N_2564);
and U2628 (N_2628,N_2563,N_2560);
or U2629 (N_2629,N_2507,N_2538);
nand U2630 (N_2630,N_2518,N_2527);
nor U2631 (N_2631,N_2546,N_2532);
nand U2632 (N_2632,N_2529,N_2559);
xnor U2633 (N_2633,N_2562,N_2583);
nand U2634 (N_2634,N_2573,N_2540);
or U2635 (N_2635,N_2556,N_2501);
xnor U2636 (N_2636,N_2568,N_2514);
nor U2637 (N_2637,N_2512,N_2509);
nand U2638 (N_2638,N_2510,N_2524);
or U2639 (N_2639,N_2541,N_2551);
xnor U2640 (N_2640,N_2548,N_2574);
and U2641 (N_2641,N_2567,N_2526);
nor U2642 (N_2642,N_2544,N_2517);
xnor U2643 (N_2643,N_2528,N_2537);
nand U2644 (N_2644,N_2591,N_2555);
or U2645 (N_2645,N_2522,N_2553);
nor U2646 (N_2646,N_2503,N_2580);
nor U2647 (N_2647,N_2570,N_2588);
nor U2648 (N_2648,N_2595,N_2584);
nand U2649 (N_2649,N_2543,N_2578);
nor U2650 (N_2650,N_2517,N_2550);
and U2651 (N_2651,N_2543,N_2537);
or U2652 (N_2652,N_2581,N_2592);
and U2653 (N_2653,N_2580,N_2568);
nor U2654 (N_2654,N_2594,N_2548);
nand U2655 (N_2655,N_2590,N_2527);
nand U2656 (N_2656,N_2590,N_2503);
nor U2657 (N_2657,N_2510,N_2599);
xor U2658 (N_2658,N_2597,N_2561);
xnor U2659 (N_2659,N_2597,N_2502);
or U2660 (N_2660,N_2524,N_2592);
and U2661 (N_2661,N_2563,N_2522);
nand U2662 (N_2662,N_2543,N_2576);
nand U2663 (N_2663,N_2579,N_2566);
and U2664 (N_2664,N_2567,N_2507);
or U2665 (N_2665,N_2500,N_2515);
or U2666 (N_2666,N_2549,N_2583);
or U2667 (N_2667,N_2513,N_2533);
nand U2668 (N_2668,N_2530,N_2573);
nand U2669 (N_2669,N_2552,N_2590);
nand U2670 (N_2670,N_2590,N_2532);
and U2671 (N_2671,N_2512,N_2551);
or U2672 (N_2672,N_2544,N_2597);
or U2673 (N_2673,N_2510,N_2534);
nand U2674 (N_2674,N_2544,N_2563);
and U2675 (N_2675,N_2515,N_2576);
or U2676 (N_2676,N_2502,N_2572);
nor U2677 (N_2677,N_2598,N_2519);
nor U2678 (N_2678,N_2526,N_2517);
and U2679 (N_2679,N_2594,N_2514);
nand U2680 (N_2680,N_2522,N_2535);
nor U2681 (N_2681,N_2522,N_2508);
and U2682 (N_2682,N_2592,N_2532);
and U2683 (N_2683,N_2531,N_2507);
nor U2684 (N_2684,N_2528,N_2564);
nand U2685 (N_2685,N_2516,N_2530);
nand U2686 (N_2686,N_2562,N_2596);
and U2687 (N_2687,N_2547,N_2567);
or U2688 (N_2688,N_2592,N_2529);
or U2689 (N_2689,N_2597,N_2563);
or U2690 (N_2690,N_2566,N_2549);
and U2691 (N_2691,N_2595,N_2507);
nand U2692 (N_2692,N_2566,N_2512);
and U2693 (N_2693,N_2536,N_2590);
nor U2694 (N_2694,N_2590,N_2558);
nand U2695 (N_2695,N_2544,N_2511);
nand U2696 (N_2696,N_2560,N_2541);
or U2697 (N_2697,N_2549,N_2514);
nor U2698 (N_2698,N_2555,N_2519);
or U2699 (N_2699,N_2524,N_2565);
nand U2700 (N_2700,N_2694,N_2693);
nor U2701 (N_2701,N_2631,N_2646);
nand U2702 (N_2702,N_2658,N_2696);
nor U2703 (N_2703,N_2605,N_2692);
nor U2704 (N_2704,N_2688,N_2624);
nand U2705 (N_2705,N_2687,N_2648);
nand U2706 (N_2706,N_2675,N_2616);
nand U2707 (N_2707,N_2666,N_2604);
and U2708 (N_2708,N_2637,N_2671);
nor U2709 (N_2709,N_2654,N_2652);
nor U2710 (N_2710,N_2651,N_2614);
nand U2711 (N_2711,N_2649,N_2657);
and U2712 (N_2712,N_2613,N_2620);
nor U2713 (N_2713,N_2639,N_2626);
nand U2714 (N_2714,N_2655,N_2608);
and U2715 (N_2715,N_2683,N_2674);
and U2716 (N_2716,N_2698,N_2603);
or U2717 (N_2717,N_2630,N_2664);
or U2718 (N_2718,N_2650,N_2686);
nor U2719 (N_2719,N_2677,N_2622);
and U2720 (N_2720,N_2660,N_2665);
and U2721 (N_2721,N_2629,N_2645);
nor U2722 (N_2722,N_2647,N_2625);
or U2723 (N_2723,N_2640,N_2627);
or U2724 (N_2724,N_2610,N_2667);
or U2725 (N_2725,N_2634,N_2697);
nor U2726 (N_2726,N_2632,N_2691);
and U2727 (N_2727,N_2621,N_2602);
or U2728 (N_2728,N_2609,N_2685);
or U2729 (N_2729,N_2661,N_2606);
and U2730 (N_2730,N_2607,N_2600);
nand U2731 (N_2731,N_2653,N_2695);
and U2732 (N_2732,N_2662,N_2680);
and U2733 (N_2733,N_2628,N_2643);
nor U2734 (N_2734,N_2681,N_2659);
or U2735 (N_2735,N_2617,N_2670);
xnor U2736 (N_2736,N_2684,N_2668);
nand U2737 (N_2737,N_2669,N_2663);
and U2738 (N_2738,N_2612,N_2689);
xor U2739 (N_2739,N_2638,N_2618);
nand U2740 (N_2740,N_2679,N_2636);
nor U2741 (N_2741,N_2642,N_2656);
or U2742 (N_2742,N_2641,N_2635);
nor U2743 (N_2743,N_2633,N_2699);
and U2744 (N_2744,N_2644,N_2623);
and U2745 (N_2745,N_2676,N_2673);
or U2746 (N_2746,N_2611,N_2678);
xnor U2747 (N_2747,N_2690,N_2619);
nor U2748 (N_2748,N_2682,N_2601);
nor U2749 (N_2749,N_2615,N_2672);
nand U2750 (N_2750,N_2665,N_2641);
nand U2751 (N_2751,N_2604,N_2659);
xor U2752 (N_2752,N_2660,N_2671);
and U2753 (N_2753,N_2639,N_2696);
nand U2754 (N_2754,N_2692,N_2662);
or U2755 (N_2755,N_2662,N_2689);
nor U2756 (N_2756,N_2677,N_2656);
xor U2757 (N_2757,N_2666,N_2646);
or U2758 (N_2758,N_2654,N_2625);
or U2759 (N_2759,N_2649,N_2670);
and U2760 (N_2760,N_2661,N_2637);
and U2761 (N_2761,N_2695,N_2671);
nand U2762 (N_2762,N_2668,N_2648);
nor U2763 (N_2763,N_2663,N_2659);
nand U2764 (N_2764,N_2660,N_2677);
xor U2765 (N_2765,N_2657,N_2671);
and U2766 (N_2766,N_2675,N_2662);
nor U2767 (N_2767,N_2664,N_2654);
or U2768 (N_2768,N_2606,N_2626);
nand U2769 (N_2769,N_2694,N_2685);
or U2770 (N_2770,N_2614,N_2641);
nand U2771 (N_2771,N_2619,N_2692);
nand U2772 (N_2772,N_2618,N_2671);
nor U2773 (N_2773,N_2664,N_2626);
xor U2774 (N_2774,N_2649,N_2655);
or U2775 (N_2775,N_2673,N_2670);
xor U2776 (N_2776,N_2659,N_2635);
nor U2777 (N_2777,N_2662,N_2695);
xnor U2778 (N_2778,N_2605,N_2609);
nor U2779 (N_2779,N_2657,N_2680);
nor U2780 (N_2780,N_2683,N_2610);
or U2781 (N_2781,N_2636,N_2622);
or U2782 (N_2782,N_2636,N_2662);
xor U2783 (N_2783,N_2621,N_2600);
nor U2784 (N_2784,N_2663,N_2630);
or U2785 (N_2785,N_2640,N_2691);
nand U2786 (N_2786,N_2601,N_2657);
or U2787 (N_2787,N_2660,N_2679);
and U2788 (N_2788,N_2635,N_2616);
or U2789 (N_2789,N_2623,N_2617);
and U2790 (N_2790,N_2670,N_2652);
nand U2791 (N_2791,N_2689,N_2656);
or U2792 (N_2792,N_2655,N_2621);
nor U2793 (N_2793,N_2632,N_2683);
xor U2794 (N_2794,N_2644,N_2665);
nor U2795 (N_2795,N_2657,N_2687);
nand U2796 (N_2796,N_2667,N_2647);
or U2797 (N_2797,N_2653,N_2692);
xor U2798 (N_2798,N_2622,N_2637);
nor U2799 (N_2799,N_2659,N_2674);
xor U2800 (N_2800,N_2742,N_2700);
nor U2801 (N_2801,N_2797,N_2720);
xnor U2802 (N_2802,N_2783,N_2778);
nand U2803 (N_2803,N_2728,N_2754);
and U2804 (N_2804,N_2788,N_2708);
nor U2805 (N_2805,N_2758,N_2761);
nand U2806 (N_2806,N_2701,N_2771);
nand U2807 (N_2807,N_2751,N_2795);
and U2808 (N_2808,N_2787,N_2765);
or U2809 (N_2809,N_2769,N_2743);
or U2810 (N_2810,N_2781,N_2791);
nand U2811 (N_2811,N_2774,N_2779);
and U2812 (N_2812,N_2723,N_2713);
and U2813 (N_2813,N_2711,N_2757);
and U2814 (N_2814,N_2741,N_2702);
nor U2815 (N_2815,N_2799,N_2782);
and U2816 (N_2816,N_2746,N_2772);
nor U2817 (N_2817,N_2704,N_2748);
nor U2818 (N_2818,N_2775,N_2730);
or U2819 (N_2819,N_2726,N_2764);
nand U2820 (N_2820,N_2763,N_2747);
or U2821 (N_2821,N_2712,N_2721);
nor U2822 (N_2822,N_2759,N_2738);
nand U2823 (N_2823,N_2784,N_2744);
nor U2824 (N_2824,N_2715,N_2770);
nand U2825 (N_2825,N_2798,N_2718);
or U2826 (N_2826,N_2729,N_2756);
nand U2827 (N_2827,N_2705,N_2727);
and U2828 (N_2828,N_2755,N_2722);
or U2829 (N_2829,N_2709,N_2749);
xor U2830 (N_2830,N_2714,N_2719);
nand U2831 (N_2831,N_2716,N_2768);
and U2832 (N_2832,N_2777,N_2734);
xnor U2833 (N_2833,N_2737,N_2796);
or U2834 (N_2834,N_2739,N_2732);
and U2835 (N_2835,N_2703,N_2762);
and U2836 (N_2836,N_2717,N_2706);
nand U2837 (N_2837,N_2773,N_2767);
and U2838 (N_2838,N_2750,N_2760);
nand U2839 (N_2839,N_2780,N_2710);
or U2840 (N_2840,N_2794,N_2766);
nor U2841 (N_2841,N_2785,N_2753);
nand U2842 (N_2842,N_2725,N_2745);
xnor U2843 (N_2843,N_2740,N_2736);
or U2844 (N_2844,N_2735,N_2786);
nor U2845 (N_2845,N_2731,N_2793);
nand U2846 (N_2846,N_2724,N_2752);
nand U2847 (N_2847,N_2707,N_2733);
and U2848 (N_2848,N_2792,N_2776);
xor U2849 (N_2849,N_2790,N_2789);
or U2850 (N_2850,N_2787,N_2715);
and U2851 (N_2851,N_2718,N_2738);
or U2852 (N_2852,N_2727,N_2723);
nand U2853 (N_2853,N_2793,N_2790);
or U2854 (N_2854,N_2719,N_2761);
or U2855 (N_2855,N_2796,N_2795);
and U2856 (N_2856,N_2798,N_2744);
and U2857 (N_2857,N_2760,N_2759);
xor U2858 (N_2858,N_2784,N_2754);
nor U2859 (N_2859,N_2726,N_2722);
or U2860 (N_2860,N_2721,N_2716);
xor U2861 (N_2861,N_2735,N_2764);
nor U2862 (N_2862,N_2733,N_2734);
and U2863 (N_2863,N_2751,N_2774);
nand U2864 (N_2864,N_2780,N_2756);
nand U2865 (N_2865,N_2712,N_2757);
nand U2866 (N_2866,N_2758,N_2780);
or U2867 (N_2867,N_2715,N_2754);
and U2868 (N_2868,N_2788,N_2717);
and U2869 (N_2869,N_2766,N_2757);
nand U2870 (N_2870,N_2723,N_2799);
nor U2871 (N_2871,N_2783,N_2791);
and U2872 (N_2872,N_2704,N_2772);
nor U2873 (N_2873,N_2777,N_2720);
nor U2874 (N_2874,N_2776,N_2794);
and U2875 (N_2875,N_2787,N_2753);
or U2876 (N_2876,N_2798,N_2739);
or U2877 (N_2877,N_2760,N_2731);
nand U2878 (N_2878,N_2735,N_2754);
or U2879 (N_2879,N_2729,N_2750);
or U2880 (N_2880,N_2720,N_2760);
nand U2881 (N_2881,N_2796,N_2759);
and U2882 (N_2882,N_2766,N_2770);
and U2883 (N_2883,N_2751,N_2771);
or U2884 (N_2884,N_2794,N_2737);
xor U2885 (N_2885,N_2794,N_2791);
nand U2886 (N_2886,N_2779,N_2754);
nand U2887 (N_2887,N_2703,N_2741);
and U2888 (N_2888,N_2795,N_2757);
nor U2889 (N_2889,N_2754,N_2722);
nor U2890 (N_2890,N_2730,N_2703);
nor U2891 (N_2891,N_2767,N_2725);
nor U2892 (N_2892,N_2793,N_2740);
and U2893 (N_2893,N_2731,N_2745);
nand U2894 (N_2894,N_2778,N_2749);
xor U2895 (N_2895,N_2765,N_2742);
nand U2896 (N_2896,N_2773,N_2722);
nor U2897 (N_2897,N_2743,N_2794);
nor U2898 (N_2898,N_2727,N_2700);
nand U2899 (N_2899,N_2719,N_2770);
nor U2900 (N_2900,N_2885,N_2874);
nor U2901 (N_2901,N_2832,N_2890);
and U2902 (N_2902,N_2809,N_2863);
nand U2903 (N_2903,N_2829,N_2826);
nor U2904 (N_2904,N_2873,N_2811);
and U2905 (N_2905,N_2896,N_2815);
or U2906 (N_2906,N_2879,N_2833);
or U2907 (N_2907,N_2869,N_2837);
nor U2908 (N_2908,N_2802,N_2824);
nand U2909 (N_2909,N_2816,N_2857);
nor U2910 (N_2910,N_2871,N_2821);
nand U2911 (N_2911,N_2839,N_2855);
nor U2912 (N_2912,N_2868,N_2875);
or U2913 (N_2913,N_2860,N_2813);
or U2914 (N_2914,N_2856,N_2817);
nor U2915 (N_2915,N_2814,N_2853);
nor U2916 (N_2916,N_2846,N_2889);
nand U2917 (N_2917,N_2897,N_2835);
nand U2918 (N_2918,N_2831,N_2820);
or U2919 (N_2919,N_2844,N_2877);
nand U2920 (N_2920,N_2800,N_2812);
nand U2921 (N_2921,N_2838,N_2825);
and U2922 (N_2922,N_2881,N_2852);
or U2923 (N_2923,N_2888,N_2851);
or U2924 (N_2924,N_2867,N_2861);
nor U2925 (N_2925,N_2858,N_2805);
and U2926 (N_2926,N_2834,N_2878);
nand U2927 (N_2927,N_2893,N_2840);
nand U2928 (N_2928,N_2848,N_2827);
or U2929 (N_2929,N_2849,N_2842);
nor U2930 (N_2930,N_2859,N_2872);
or U2931 (N_2931,N_2882,N_2818);
and U2932 (N_2932,N_2836,N_2822);
nand U2933 (N_2933,N_2801,N_2854);
and U2934 (N_2934,N_2843,N_2864);
nor U2935 (N_2935,N_2883,N_2804);
xor U2936 (N_2936,N_2887,N_2891);
or U2937 (N_2937,N_2819,N_2870);
and U2938 (N_2938,N_2865,N_2862);
nand U2939 (N_2939,N_2828,N_2806);
and U2940 (N_2940,N_2847,N_2880);
nand U2941 (N_2941,N_2886,N_2823);
nor U2942 (N_2942,N_2895,N_2884);
nand U2943 (N_2943,N_2807,N_2898);
or U2944 (N_2944,N_2894,N_2866);
or U2945 (N_2945,N_2810,N_2876);
and U2946 (N_2946,N_2841,N_2850);
nor U2947 (N_2947,N_2803,N_2892);
nor U2948 (N_2948,N_2808,N_2899);
nand U2949 (N_2949,N_2830,N_2845);
and U2950 (N_2950,N_2848,N_2837);
nand U2951 (N_2951,N_2865,N_2858);
nor U2952 (N_2952,N_2815,N_2832);
and U2953 (N_2953,N_2853,N_2830);
nor U2954 (N_2954,N_2827,N_2885);
or U2955 (N_2955,N_2883,N_2871);
nand U2956 (N_2956,N_2895,N_2813);
nor U2957 (N_2957,N_2850,N_2801);
nand U2958 (N_2958,N_2887,N_2880);
nand U2959 (N_2959,N_2840,N_2877);
or U2960 (N_2960,N_2807,N_2822);
nor U2961 (N_2961,N_2830,N_2841);
or U2962 (N_2962,N_2849,N_2875);
nand U2963 (N_2963,N_2813,N_2840);
and U2964 (N_2964,N_2828,N_2808);
nor U2965 (N_2965,N_2826,N_2864);
nor U2966 (N_2966,N_2843,N_2831);
nor U2967 (N_2967,N_2849,N_2856);
and U2968 (N_2968,N_2810,N_2878);
or U2969 (N_2969,N_2859,N_2877);
nor U2970 (N_2970,N_2808,N_2842);
nand U2971 (N_2971,N_2898,N_2825);
xor U2972 (N_2972,N_2898,N_2869);
and U2973 (N_2973,N_2842,N_2823);
or U2974 (N_2974,N_2880,N_2843);
nor U2975 (N_2975,N_2836,N_2860);
nor U2976 (N_2976,N_2829,N_2893);
and U2977 (N_2977,N_2847,N_2894);
and U2978 (N_2978,N_2872,N_2880);
nor U2979 (N_2979,N_2841,N_2865);
and U2980 (N_2980,N_2843,N_2821);
and U2981 (N_2981,N_2815,N_2879);
nand U2982 (N_2982,N_2839,N_2878);
nand U2983 (N_2983,N_2835,N_2858);
nand U2984 (N_2984,N_2860,N_2892);
or U2985 (N_2985,N_2867,N_2884);
or U2986 (N_2986,N_2817,N_2809);
or U2987 (N_2987,N_2828,N_2894);
or U2988 (N_2988,N_2824,N_2899);
and U2989 (N_2989,N_2875,N_2822);
nand U2990 (N_2990,N_2891,N_2808);
or U2991 (N_2991,N_2870,N_2874);
nand U2992 (N_2992,N_2872,N_2861);
or U2993 (N_2993,N_2885,N_2849);
and U2994 (N_2994,N_2838,N_2856);
or U2995 (N_2995,N_2867,N_2808);
nor U2996 (N_2996,N_2842,N_2834);
xnor U2997 (N_2997,N_2813,N_2854);
xnor U2998 (N_2998,N_2899,N_2877);
nand U2999 (N_2999,N_2846,N_2803);
xor U3000 (N_3000,N_2987,N_2924);
nor U3001 (N_3001,N_2991,N_2938);
nand U3002 (N_3002,N_2929,N_2914);
or U3003 (N_3003,N_2901,N_2954);
xnor U3004 (N_3004,N_2998,N_2916);
or U3005 (N_3005,N_2968,N_2970);
or U3006 (N_3006,N_2956,N_2967);
or U3007 (N_3007,N_2941,N_2911);
nor U3008 (N_3008,N_2995,N_2993);
or U3009 (N_3009,N_2958,N_2978);
or U3010 (N_3010,N_2955,N_2928);
and U3011 (N_3011,N_2962,N_2939);
nand U3012 (N_3012,N_2944,N_2990);
nand U3013 (N_3013,N_2900,N_2980);
nor U3014 (N_3014,N_2930,N_2981);
and U3015 (N_3015,N_2971,N_2952);
and U3016 (N_3016,N_2948,N_2963);
or U3017 (N_3017,N_2909,N_2918);
or U3018 (N_3018,N_2917,N_2965);
xnor U3019 (N_3019,N_2947,N_2932);
or U3020 (N_3020,N_2996,N_2985);
nor U3021 (N_3021,N_2988,N_2935);
and U3022 (N_3022,N_2982,N_2910);
and U3023 (N_3023,N_2975,N_2979);
or U3024 (N_3024,N_2950,N_2926);
and U3025 (N_3025,N_2961,N_2994);
nand U3026 (N_3026,N_2920,N_2977);
nor U3027 (N_3027,N_2942,N_2915);
nand U3028 (N_3028,N_2986,N_2933);
or U3029 (N_3029,N_2960,N_2943);
nand U3030 (N_3030,N_2922,N_2984);
nand U3031 (N_3031,N_2903,N_2964);
or U3032 (N_3032,N_2905,N_2953);
xor U3033 (N_3033,N_2999,N_2936);
or U3034 (N_3034,N_2937,N_2966);
or U3035 (N_3035,N_2921,N_2983);
nand U3036 (N_3036,N_2908,N_2989);
nor U3037 (N_3037,N_2913,N_2904);
or U3038 (N_3038,N_2927,N_2912);
and U3039 (N_3039,N_2949,N_2976);
xnor U3040 (N_3040,N_2946,N_2951);
and U3041 (N_3041,N_2972,N_2934);
nand U3042 (N_3042,N_2973,N_2940);
or U3043 (N_3043,N_2945,N_2957);
or U3044 (N_3044,N_2907,N_2959);
or U3045 (N_3045,N_2931,N_2923);
nand U3046 (N_3046,N_2992,N_2906);
and U3047 (N_3047,N_2902,N_2925);
nand U3048 (N_3048,N_2969,N_2997);
or U3049 (N_3049,N_2974,N_2919);
nor U3050 (N_3050,N_2913,N_2951);
nor U3051 (N_3051,N_2988,N_2998);
and U3052 (N_3052,N_2972,N_2924);
or U3053 (N_3053,N_2964,N_2994);
and U3054 (N_3054,N_2918,N_2995);
or U3055 (N_3055,N_2978,N_2936);
and U3056 (N_3056,N_2948,N_2999);
xnor U3057 (N_3057,N_2902,N_2992);
and U3058 (N_3058,N_2988,N_2915);
and U3059 (N_3059,N_2935,N_2989);
nand U3060 (N_3060,N_2973,N_2996);
nand U3061 (N_3061,N_2992,N_2929);
and U3062 (N_3062,N_2993,N_2955);
nor U3063 (N_3063,N_2949,N_2979);
and U3064 (N_3064,N_2945,N_2906);
nand U3065 (N_3065,N_2973,N_2937);
nand U3066 (N_3066,N_2980,N_2903);
nand U3067 (N_3067,N_2938,N_2906);
nand U3068 (N_3068,N_2925,N_2998);
nand U3069 (N_3069,N_2905,N_2902);
nor U3070 (N_3070,N_2931,N_2916);
nor U3071 (N_3071,N_2966,N_2952);
nand U3072 (N_3072,N_2910,N_2932);
and U3073 (N_3073,N_2924,N_2913);
nand U3074 (N_3074,N_2914,N_2955);
nand U3075 (N_3075,N_2968,N_2995);
nand U3076 (N_3076,N_2920,N_2928);
nand U3077 (N_3077,N_2951,N_2911);
nor U3078 (N_3078,N_2980,N_2963);
and U3079 (N_3079,N_2941,N_2915);
xor U3080 (N_3080,N_2991,N_2971);
nand U3081 (N_3081,N_2994,N_2957);
nand U3082 (N_3082,N_2976,N_2925);
xnor U3083 (N_3083,N_2964,N_2908);
or U3084 (N_3084,N_2961,N_2974);
or U3085 (N_3085,N_2973,N_2960);
xnor U3086 (N_3086,N_2907,N_2979);
nor U3087 (N_3087,N_2971,N_2978);
and U3088 (N_3088,N_2957,N_2908);
and U3089 (N_3089,N_2924,N_2937);
or U3090 (N_3090,N_2925,N_2907);
and U3091 (N_3091,N_2907,N_2968);
and U3092 (N_3092,N_2998,N_2983);
nand U3093 (N_3093,N_2985,N_2998);
nand U3094 (N_3094,N_2955,N_2989);
and U3095 (N_3095,N_2908,N_2969);
nor U3096 (N_3096,N_2993,N_2969);
nand U3097 (N_3097,N_2941,N_2919);
or U3098 (N_3098,N_2909,N_2980);
nand U3099 (N_3099,N_2911,N_2916);
nor U3100 (N_3100,N_3019,N_3026);
or U3101 (N_3101,N_3044,N_3034);
nor U3102 (N_3102,N_3081,N_3071);
nor U3103 (N_3103,N_3067,N_3089);
nand U3104 (N_3104,N_3069,N_3090);
and U3105 (N_3105,N_3094,N_3014);
nor U3106 (N_3106,N_3084,N_3011);
or U3107 (N_3107,N_3021,N_3099);
nor U3108 (N_3108,N_3045,N_3027);
nor U3109 (N_3109,N_3066,N_3055);
nand U3110 (N_3110,N_3073,N_3062);
xor U3111 (N_3111,N_3018,N_3063);
and U3112 (N_3112,N_3036,N_3048);
nor U3113 (N_3113,N_3086,N_3038);
and U3114 (N_3114,N_3007,N_3041);
nor U3115 (N_3115,N_3075,N_3097);
or U3116 (N_3116,N_3060,N_3005);
nor U3117 (N_3117,N_3050,N_3072);
and U3118 (N_3118,N_3095,N_3098);
and U3119 (N_3119,N_3083,N_3059);
nand U3120 (N_3120,N_3043,N_3047);
or U3121 (N_3121,N_3056,N_3017);
nor U3122 (N_3122,N_3054,N_3016);
and U3123 (N_3123,N_3057,N_3096);
or U3124 (N_3124,N_3042,N_3035);
or U3125 (N_3125,N_3046,N_3087);
nand U3126 (N_3126,N_3093,N_3092);
xnor U3127 (N_3127,N_3085,N_3000);
nor U3128 (N_3128,N_3082,N_3061);
xnor U3129 (N_3129,N_3070,N_3010);
xnor U3130 (N_3130,N_3032,N_3004);
nand U3131 (N_3131,N_3052,N_3088);
nor U3132 (N_3132,N_3040,N_3080);
xnor U3133 (N_3133,N_3015,N_3020);
nor U3134 (N_3134,N_3076,N_3091);
or U3135 (N_3135,N_3065,N_3058);
or U3136 (N_3136,N_3074,N_3078);
nor U3137 (N_3137,N_3029,N_3008);
and U3138 (N_3138,N_3079,N_3006);
and U3139 (N_3139,N_3030,N_3053);
nor U3140 (N_3140,N_3024,N_3039);
nor U3141 (N_3141,N_3028,N_3064);
or U3142 (N_3142,N_3033,N_3003);
nand U3143 (N_3143,N_3077,N_3051);
or U3144 (N_3144,N_3049,N_3023);
or U3145 (N_3145,N_3012,N_3068);
or U3146 (N_3146,N_3009,N_3025);
and U3147 (N_3147,N_3013,N_3002);
and U3148 (N_3148,N_3001,N_3037);
nor U3149 (N_3149,N_3022,N_3031);
nand U3150 (N_3150,N_3061,N_3087);
nor U3151 (N_3151,N_3004,N_3030);
and U3152 (N_3152,N_3089,N_3049);
nand U3153 (N_3153,N_3007,N_3076);
nor U3154 (N_3154,N_3024,N_3072);
nand U3155 (N_3155,N_3025,N_3018);
and U3156 (N_3156,N_3038,N_3012);
or U3157 (N_3157,N_3010,N_3049);
xor U3158 (N_3158,N_3084,N_3043);
nor U3159 (N_3159,N_3015,N_3024);
nand U3160 (N_3160,N_3070,N_3028);
nand U3161 (N_3161,N_3094,N_3086);
nand U3162 (N_3162,N_3029,N_3094);
nand U3163 (N_3163,N_3012,N_3048);
nand U3164 (N_3164,N_3018,N_3087);
nand U3165 (N_3165,N_3005,N_3090);
or U3166 (N_3166,N_3024,N_3041);
nor U3167 (N_3167,N_3072,N_3040);
or U3168 (N_3168,N_3087,N_3058);
nand U3169 (N_3169,N_3089,N_3094);
and U3170 (N_3170,N_3043,N_3044);
nand U3171 (N_3171,N_3076,N_3070);
and U3172 (N_3172,N_3051,N_3025);
or U3173 (N_3173,N_3085,N_3093);
nand U3174 (N_3174,N_3014,N_3077);
nor U3175 (N_3175,N_3012,N_3036);
or U3176 (N_3176,N_3073,N_3075);
xnor U3177 (N_3177,N_3031,N_3024);
nand U3178 (N_3178,N_3095,N_3020);
and U3179 (N_3179,N_3069,N_3006);
or U3180 (N_3180,N_3088,N_3075);
or U3181 (N_3181,N_3032,N_3042);
or U3182 (N_3182,N_3009,N_3028);
xor U3183 (N_3183,N_3060,N_3010);
and U3184 (N_3184,N_3093,N_3029);
nand U3185 (N_3185,N_3093,N_3065);
nand U3186 (N_3186,N_3011,N_3059);
or U3187 (N_3187,N_3042,N_3023);
nand U3188 (N_3188,N_3022,N_3035);
or U3189 (N_3189,N_3031,N_3026);
nand U3190 (N_3190,N_3068,N_3031);
nor U3191 (N_3191,N_3044,N_3054);
or U3192 (N_3192,N_3099,N_3028);
and U3193 (N_3193,N_3062,N_3063);
xnor U3194 (N_3194,N_3043,N_3096);
xor U3195 (N_3195,N_3084,N_3047);
nand U3196 (N_3196,N_3010,N_3021);
and U3197 (N_3197,N_3012,N_3049);
and U3198 (N_3198,N_3013,N_3035);
nand U3199 (N_3199,N_3053,N_3084);
and U3200 (N_3200,N_3196,N_3174);
nand U3201 (N_3201,N_3145,N_3157);
nor U3202 (N_3202,N_3118,N_3112);
or U3203 (N_3203,N_3189,N_3137);
nand U3204 (N_3204,N_3142,N_3123);
nor U3205 (N_3205,N_3114,N_3194);
and U3206 (N_3206,N_3152,N_3104);
xor U3207 (N_3207,N_3120,N_3165);
and U3208 (N_3208,N_3163,N_3166);
nor U3209 (N_3209,N_3159,N_3143);
nor U3210 (N_3210,N_3138,N_3121);
xnor U3211 (N_3211,N_3124,N_3140);
and U3212 (N_3212,N_3126,N_3117);
nand U3213 (N_3213,N_3115,N_3182);
nor U3214 (N_3214,N_3141,N_3100);
nand U3215 (N_3215,N_3193,N_3156);
or U3216 (N_3216,N_3135,N_3186);
nand U3217 (N_3217,N_3158,N_3187);
and U3218 (N_3218,N_3128,N_3134);
or U3219 (N_3219,N_3151,N_3192);
nand U3220 (N_3220,N_3122,N_3136);
nand U3221 (N_3221,N_3102,N_3129);
or U3222 (N_3222,N_3103,N_3171);
nand U3223 (N_3223,N_3149,N_3148);
nor U3224 (N_3224,N_3133,N_3116);
and U3225 (N_3225,N_3132,N_3175);
nand U3226 (N_3226,N_3125,N_3176);
or U3227 (N_3227,N_3107,N_3153);
xnor U3228 (N_3228,N_3188,N_3190);
and U3229 (N_3229,N_3110,N_3184);
or U3230 (N_3230,N_3183,N_3147);
and U3231 (N_3231,N_3106,N_3150);
or U3232 (N_3232,N_3169,N_3162);
and U3233 (N_3233,N_3179,N_3154);
nor U3234 (N_3234,N_3178,N_3195);
nor U3235 (N_3235,N_3164,N_3173);
or U3236 (N_3236,N_3198,N_3105);
nand U3237 (N_3237,N_3130,N_3139);
nor U3238 (N_3238,N_3101,N_3197);
nand U3239 (N_3239,N_3167,N_3160);
or U3240 (N_3240,N_3170,N_3113);
nand U3241 (N_3241,N_3127,N_3199);
and U3242 (N_3242,N_3181,N_3131);
nor U3243 (N_3243,N_3146,N_3109);
nand U3244 (N_3244,N_3108,N_3119);
or U3245 (N_3245,N_3155,N_3161);
and U3246 (N_3246,N_3168,N_3185);
nand U3247 (N_3247,N_3144,N_3191);
or U3248 (N_3248,N_3172,N_3177);
nand U3249 (N_3249,N_3111,N_3180);
or U3250 (N_3250,N_3157,N_3196);
and U3251 (N_3251,N_3167,N_3109);
xnor U3252 (N_3252,N_3157,N_3106);
nor U3253 (N_3253,N_3135,N_3196);
nor U3254 (N_3254,N_3136,N_3137);
nand U3255 (N_3255,N_3128,N_3127);
and U3256 (N_3256,N_3178,N_3184);
xnor U3257 (N_3257,N_3155,N_3178);
or U3258 (N_3258,N_3190,N_3158);
or U3259 (N_3259,N_3110,N_3113);
nand U3260 (N_3260,N_3101,N_3100);
nor U3261 (N_3261,N_3182,N_3107);
and U3262 (N_3262,N_3193,N_3126);
or U3263 (N_3263,N_3181,N_3108);
nand U3264 (N_3264,N_3134,N_3149);
and U3265 (N_3265,N_3139,N_3182);
nand U3266 (N_3266,N_3147,N_3154);
nor U3267 (N_3267,N_3173,N_3163);
nand U3268 (N_3268,N_3173,N_3174);
or U3269 (N_3269,N_3197,N_3131);
nand U3270 (N_3270,N_3175,N_3149);
or U3271 (N_3271,N_3166,N_3154);
or U3272 (N_3272,N_3153,N_3139);
nand U3273 (N_3273,N_3131,N_3183);
nand U3274 (N_3274,N_3125,N_3177);
nor U3275 (N_3275,N_3120,N_3136);
nor U3276 (N_3276,N_3103,N_3131);
and U3277 (N_3277,N_3162,N_3197);
xor U3278 (N_3278,N_3148,N_3128);
nor U3279 (N_3279,N_3175,N_3127);
nor U3280 (N_3280,N_3199,N_3172);
or U3281 (N_3281,N_3190,N_3199);
nor U3282 (N_3282,N_3158,N_3197);
and U3283 (N_3283,N_3120,N_3127);
and U3284 (N_3284,N_3152,N_3159);
nor U3285 (N_3285,N_3127,N_3197);
or U3286 (N_3286,N_3144,N_3161);
and U3287 (N_3287,N_3165,N_3134);
nand U3288 (N_3288,N_3139,N_3155);
or U3289 (N_3289,N_3175,N_3129);
nor U3290 (N_3290,N_3172,N_3118);
xor U3291 (N_3291,N_3119,N_3174);
nand U3292 (N_3292,N_3101,N_3121);
nor U3293 (N_3293,N_3194,N_3195);
or U3294 (N_3294,N_3156,N_3154);
nand U3295 (N_3295,N_3102,N_3163);
nor U3296 (N_3296,N_3125,N_3137);
or U3297 (N_3297,N_3184,N_3137);
xor U3298 (N_3298,N_3135,N_3140);
nand U3299 (N_3299,N_3154,N_3130);
and U3300 (N_3300,N_3223,N_3220);
and U3301 (N_3301,N_3215,N_3271);
xor U3302 (N_3302,N_3221,N_3237);
and U3303 (N_3303,N_3277,N_3236);
nor U3304 (N_3304,N_3234,N_3243);
or U3305 (N_3305,N_3268,N_3206);
or U3306 (N_3306,N_3257,N_3227);
and U3307 (N_3307,N_3245,N_3289);
nand U3308 (N_3308,N_3274,N_3238);
nand U3309 (N_3309,N_3283,N_3228);
nand U3310 (N_3310,N_3284,N_3280);
and U3311 (N_3311,N_3248,N_3203);
and U3312 (N_3312,N_3265,N_3230);
nor U3313 (N_3313,N_3211,N_3252);
xor U3314 (N_3314,N_3273,N_3299);
and U3315 (N_3315,N_3270,N_3249);
nand U3316 (N_3316,N_3276,N_3225);
nand U3317 (N_3317,N_3294,N_3285);
or U3318 (N_3318,N_3207,N_3290);
nor U3319 (N_3319,N_3247,N_3250);
or U3320 (N_3320,N_3232,N_3200);
nor U3321 (N_3321,N_3264,N_3214);
and U3322 (N_3322,N_3224,N_3278);
nor U3323 (N_3323,N_3288,N_3239);
xor U3324 (N_3324,N_3205,N_3260);
nor U3325 (N_3325,N_3254,N_3235);
nand U3326 (N_3326,N_3287,N_3229);
nand U3327 (N_3327,N_3209,N_3253);
nand U3328 (N_3328,N_3233,N_3275);
and U3329 (N_3329,N_3202,N_3258);
nor U3330 (N_3330,N_3246,N_3231);
or U3331 (N_3331,N_3222,N_3216);
and U3332 (N_3332,N_3298,N_3259);
and U3333 (N_3333,N_3262,N_3219);
and U3334 (N_3334,N_3267,N_3217);
or U3335 (N_3335,N_3201,N_3266);
xnor U3336 (N_3336,N_3244,N_3208);
or U3337 (N_3337,N_3293,N_3292);
and U3338 (N_3338,N_3272,N_3255);
nand U3339 (N_3339,N_3213,N_3240);
nor U3340 (N_3340,N_3269,N_3204);
xor U3341 (N_3341,N_3281,N_3286);
or U3342 (N_3342,N_3212,N_3296);
and U3343 (N_3343,N_3282,N_3251);
nand U3344 (N_3344,N_3261,N_3241);
or U3345 (N_3345,N_3218,N_3297);
or U3346 (N_3346,N_3210,N_3242);
nor U3347 (N_3347,N_3226,N_3279);
or U3348 (N_3348,N_3291,N_3263);
or U3349 (N_3349,N_3295,N_3256);
and U3350 (N_3350,N_3291,N_3233);
nor U3351 (N_3351,N_3216,N_3277);
and U3352 (N_3352,N_3280,N_3292);
nand U3353 (N_3353,N_3273,N_3275);
nor U3354 (N_3354,N_3215,N_3245);
nand U3355 (N_3355,N_3254,N_3225);
or U3356 (N_3356,N_3230,N_3258);
nand U3357 (N_3357,N_3273,N_3232);
xnor U3358 (N_3358,N_3272,N_3277);
nand U3359 (N_3359,N_3240,N_3231);
nand U3360 (N_3360,N_3291,N_3253);
nor U3361 (N_3361,N_3249,N_3285);
nand U3362 (N_3362,N_3277,N_3263);
nand U3363 (N_3363,N_3252,N_3203);
nand U3364 (N_3364,N_3226,N_3222);
xnor U3365 (N_3365,N_3258,N_3250);
or U3366 (N_3366,N_3295,N_3206);
or U3367 (N_3367,N_3278,N_3254);
and U3368 (N_3368,N_3274,N_3230);
and U3369 (N_3369,N_3287,N_3256);
or U3370 (N_3370,N_3204,N_3209);
and U3371 (N_3371,N_3257,N_3279);
nor U3372 (N_3372,N_3291,N_3220);
nor U3373 (N_3373,N_3236,N_3256);
or U3374 (N_3374,N_3292,N_3203);
and U3375 (N_3375,N_3220,N_3240);
nand U3376 (N_3376,N_3287,N_3266);
nand U3377 (N_3377,N_3294,N_3206);
nor U3378 (N_3378,N_3253,N_3251);
nor U3379 (N_3379,N_3297,N_3223);
or U3380 (N_3380,N_3261,N_3285);
nand U3381 (N_3381,N_3209,N_3210);
nor U3382 (N_3382,N_3281,N_3204);
nor U3383 (N_3383,N_3247,N_3297);
or U3384 (N_3384,N_3267,N_3277);
and U3385 (N_3385,N_3262,N_3232);
nor U3386 (N_3386,N_3226,N_3228);
or U3387 (N_3387,N_3291,N_3243);
and U3388 (N_3388,N_3264,N_3260);
and U3389 (N_3389,N_3211,N_3209);
and U3390 (N_3390,N_3296,N_3217);
xor U3391 (N_3391,N_3260,N_3237);
nor U3392 (N_3392,N_3205,N_3289);
and U3393 (N_3393,N_3247,N_3276);
nand U3394 (N_3394,N_3219,N_3298);
nor U3395 (N_3395,N_3251,N_3211);
nor U3396 (N_3396,N_3239,N_3231);
nand U3397 (N_3397,N_3210,N_3230);
xor U3398 (N_3398,N_3253,N_3206);
or U3399 (N_3399,N_3215,N_3233);
nor U3400 (N_3400,N_3396,N_3344);
nor U3401 (N_3401,N_3307,N_3389);
xor U3402 (N_3402,N_3328,N_3358);
and U3403 (N_3403,N_3385,N_3354);
nand U3404 (N_3404,N_3330,N_3313);
nor U3405 (N_3405,N_3382,N_3336);
or U3406 (N_3406,N_3342,N_3341);
nor U3407 (N_3407,N_3349,N_3376);
nor U3408 (N_3408,N_3332,N_3317);
or U3409 (N_3409,N_3318,N_3325);
nor U3410 (N_3410,N_3390,N_3378);
nand U3411 (N_3411,N_3365,N_3361);
nand U3412 (N_3412,N_3345,N_3329);
nor U3413 (N_3413,N_3327,N_3340);
nor U3414 (N_3414,N_3305,N_3374);
and U3415 (N_3415,N_3322,N_3360);
and U3416 (N_3416,N_3366,N_3356);
nand U3417 (N_3417,N_3309,N_3363);
nor U3418 (N_3418,N_3352,N_3310);
nand U3419 (N_3419,N_3324,N_3381);
xnor U3420 (N_3420,N_3370,N_3302);
and U3421 (N_3421,N_3368,N_3306);
or U3422 (N_3422,N_3399,N_3393);
nor U3423 (N_3423,N_3312,N_3321);
nor U3424 (N_3424,N_3364,N_3371);
nand U3425 (N_3425,N_3369,N_3347);
and U3426 (N_3426,N_3362,N_3333);
nor U3427 (N_3427,N_3398,N_3343);
nand U3428 (N_3428,N_3377,N_3335);
or U3429 (N_3429,N_3392,N_3346);
xnor U3430 (N_3430,N_3394,N_3380);
and U3431 (N_3431,N_3315,N_3334);
nand U3432 (N_3432,N_3331,N_3373);
or U3433 (N_3433,N_3301,N_3372);
nor U3434 (N_3434,N_3311,N_3386);
nand U3435 (N_3435,N_3339,N_3359);
nor U3436 (N_3436,N_3303,N_3397);
nand U3437 (N_3437,N_3391,N_3338);
nor U3438 (N_3438,N_3384,N_3379);
xor U3439 (N_3439,N_3351,N_3326);
nor U3440 (N_3440,N_3304,N_3316);
nand U3441 (N_3441,N_3357,N_3383);
nand U3442 (N_3442,N_3348,N_3375);
and U3443 (N_3443,N_3319,N_3387);
nand U3444 (N_3444,N_3323,N_3320);
nand U3445 (N_3445,N_3395,N_3308);
nor U3446 (N_3446,N_3314,N_3350);
nor U3447 (N_3447,N_3337,N_3353);
nand U3448 (N_3448,N_3388,N_3367);
and U3449 (N_3449,N_3355,N_3300);
nand U3450 (N_3450,N_3383,N_3345);
nand U3451 (N_3451,N_3345,N_3393);
nand U3452 (N_3452,N_3339,N_3302);
nor U3453 (N_3453,N_3320,N_3306);
nor U3454 (N_3454,N_3387,N_3363);
and U3455 (N_3455,N_3379,N_3382);
or U3456 (N_3456,N_3339,N_3384);
nand U3457 (N_3457,N_3385,N_3328);
nand U3458 (N_3458,N_3321,N_3318);
and U3459 (N_3459,N_3341,N_3399);
or U3460 (N_3460,N_3345,N_3369);
xor U3461 (N_3461,N_3319,N_3361);
nor U3462 (N_3462,N_3376,N_3304);
nand U3463 (N_3463,N_3310,N_3302);
and U3464 (N_3464,N_3352,N_3306);
nor U3465 (N_3465,N_3345,N_3332);
xnor U3466 (N_3466,N_3364,N_3369);
nand U3467 (N_3467,N_3380,N_3349);
nor U3468 (N_3468,N_3388,N_3337);
and U3469 (N_3469,N_3362,N_3343);
nor U3470 (N_3470,N_3344,N_3379);
nor U3471 (N_3471,N_3305,N_3316);
and U3472 (N_3472,N_3392,N_3330);
xor U3473 (N_3473,N_3307,N_3344);
or U3474 (N_3474,N_3333,N_3360);
or U3475 (N_3475,N_3335,N_3336);
nor U3476 (N_3476,N_3317,N_3323);
nor U3477 (N_3477,N_3390,N_3343);
or U3478 (N_3478,N_3314,N_3384);
nand U3479 (N_3479,N_3380,N_3347);
or U3480 (N_3480,N_3328,N_3355);
nand U3481 (N_3481,N_3334,N_3391);
nor U3482 (N_3482,N_3330,N_3364);
nand U3483 (N_3483,N_3350,N_3317);
nand U3484 (N_3484,N_3307,N_3327);
or U3485 (N_3485,N_3300,N_3317);
xnor U3486 (N_3486,N_3367,N_3345);
or U3487 (N_3487,N_3399,N_3378);
xor U3488 (N_3488,N_3336,N_3314);
nor U3489 (N_3489,N_3359,N_3352);
nor U3490 (N_3490,N_3357,N_3329);
and U3491 (N_3491,N_3328,N_3387);
or U3492 (N_3492,N_3367,N_3369);
nor U3493 (N_3493,N_3337,N_3356);
nor U3494 (N_3494,N_3341,N_3334);
xor U3495 (N_3495,N_3392,N_3321);
xor U3496 (N_3496,N_3331,N_3302);
and U3497 (N_3497,N_3330,N_3368);
nor U3498 (N_3498,N_3321,N_3355);
nand U3499 (N_3499,N_3371,N_3333);
or U3500 (N_3500,N_3405,N_3437);
nand U3501 (N_3501,N_3498,N_3486);
and U3502 (N_3502,N_3474,N_3427);
nor U3503 (N_3503,N_3432,N_3431);
nor U3504 (N_3504,N_3447,N_3455);
xnor U3505 (N_3505,N_3414,N_3457);
or U3506 (N_3506,N_3407,N_3442);
and U3507 (N_3507,N_3422,N_3409);
or U3508 (N_3508,N_3492,N_3443);
nand U3509 (N_3509,N_3456,N_3448);
nand U3510 (N_3510,N_3461,N_3458);
nor U3511 (N_3511,N_3404,N_3425);
or U3512 (N_3512,N_3468,N_3454);
and U3513 (N_3513,N_3487,N_3491);
nor U3514 (N_3514,N_3403,N_3412);
xnor U3515 (N_3515,N_3430,N_3482);
or U3516 (N_3516,N_3444,N_3459);
and U3517 (N_3517,N_3421,N_3424);
and U3518 (N_3518,N_3433,N_3472);
xor U3519 (N_3519,N_3466,N_3411);
nand U3520 (N_3520,N_3480,N_3462);
and U3521 (N_3521,N_3453,N_3475);
or U3522 (N_3522,N_3493,N_3495);
and U3523 (N_3523,N_3467,N_3406);
nand U3524 (N_3524,N_3452,N_3441);
xor U3525 (N_3525,N_3479,N_3499);
and U3526 (N_3526,N_3477,N_3496);
and U3527 (N_3527,N_3402,N_3439);
and U3528 (N_3528,N_3428,N_3445);
and U3529 (N_3529,N_3484,N_3446);
nand U3530 (N_3530,N_3469,N_3408);
or U3531 (N_3531,N_3436,N_3470);
or U3532 (N_3532,N_3490,N_3451);
nor U3533 (N_3533,N_3464,N_3418);
nor U3534 (N_3534,N_3460,N_3473);
nor U3535 (N_3535,N_3438,N_3400);
nand U3536 (N_3536,N_3434,N_3440);
nand U3537 (N_3537,N_3450,N_3419);
or U3538 (N_3538,N_3485,N_3413);
or U3539 (N_3539,N_3478,N_3415);
and U3540 (N_3540,N_3483,N_3423);
and U3541 (N_3541,N_3481,N_3435);
xnor U3542 (N_3542,N_3476,N_3497);
xnor U3543 (N_3543,N_3426,N_3417);
or U3544 (N_3544,N_3429,N_3463);
xor U3545 (N_3545,N_3449,N_3410);
xnor U3546 (N_3546,N_3416,N_3471);
xor U3547 (N_3547,N_3420,N_3494);
and U3548 (N_3548,N_3489,N_3465);
nand U3549 (N_3549,N_3488,N_3401);
nor U3550 (N_3550,N_3423,N_3470);
nand U3551 (N_3551,N_3487,N_3401);
or U3552 (N_3552,N_3497,N_3467);
and U3553 (N_3553,N_3408,N_3477);
nand U3554 (N_3554,N_3416,N_3445);
or U3555 (N_3555,N_3409,N_3431);
nand U3556 (N_3556,N_3409,N_3491);
or U3557 (N_3557,N_3496,N_3414);
nand U3558 (N_3558,N_3484,N_3408);
and U3559 (N_3559,N_3452,N_3494);
and U3560 (N_3560,N_3497,N_3477);
and U3561 (N_3561,N_3494,N_3402);
or U3562 (N_3562,N_3461,N_3488);
nor U3563 (N_3563,N_3436,N_3421);
and U3564 (N_3564,N_3469,N_3409);
nand U3565 (N_3565,N_3458,N_3481);
or U3566 (N_3566,N_3463,N_3436);
xor U3567 (N_3567,N_3411,N_3420);
and U3568 (N_3568,N_3477,N_3468);
xnor U3569 (N_3569,N_3408,N_3446);
nand U3570 (N_3570,N_3457,N_3406);
nor U3571 (N_3571,N_3494,N_3438);
or U3572 (N_3572,N_3472,N_3490);
nor U3573 (N_3573,N_3489,N_3486);
nor U3574 (N_3574,N_3453,N_3421);
and U3575 (N_3575,N_3436,N_3492);
xnor U3576 (N_3576,N_3448,N_3466);
or U3577 (N_3577,N_3499,N_3431);
or U3578 (N_3578,N_3475,N_3422);
and U3579 (N_3579,N_3455,N_3427);
nand U3580 (N_3580,N_3403,N_3489);
and U3581 (N_3581,N_3436,N_3403);
xnor U3582 (N_3582,N_3496,N_3422);
nor U3583 (N_3583,N_3471,N_3486);
xor U3584 (N_3584,N_3490,N_3457);
nor U3585 (N_3585,N_3486,N_3455);
nor U3586 (N_3586,N_3456,N_3481);
xnor U3587 (N_3587,N_3428,N_3466);
nor U3588 (N_3588,N_3445,N_3405);
or U3589 (N_3589,N_3471,N_3431);
nand U3590 (N_3590,N_3431,N_3472);
nand U3591 (N_3591,N_3470,N_3469);
nor U3592 (N_3592,N_3471,N_3458);
xor U3593 (N_3593,N_3462,N_3423);
and U3594 (N_3594,N_3460,N_3461);
or U3595 (N_3595,N_3471,N_3403);
nand U3596 (N_3596,N_3408,N_3461);
nor U3597 (N_3597,N_3474,N_3467);
and U3598 (N_3598,N_3499,N_3423);
xnor U3599 (N_3599,N_3426,N_3457);
nor U3600 (N_3600,N_3576,N_3579);
nand U3601 (N_3601,N_3531,N_3547);
nor U3602 (N_3602,N_3538,N_3566);
or U3603 (N_3603,N_3511,N_3528);
nand U3604 (N_3604,N_3548,N_3508);
nand U3605 (N_3605,N_3561,N_3556);
or U3606 (N_3606,N_3559,N_3587);
nor U3607 (N_3607,N_3560,N_3570);
nor U3608 (N_3608,N_3518,N_3504);
nor U3609 (N_3609,N_3529,N_3539);
nor U3610 (N_3610,N_3537,N_3563);
or U3611 (N_3611,N_3581,N_3567);
and U3612 (N_3612,N_3526,N_3507);
nor U3613 (N_3613,N_3501,N_3588);
nand U3614 (N_3614,N_3525,N_3589);
nand U3615 (N_3615,N_3586,N_3549);
or U3616 (N_3616,N_3564,N_3505);
nand U3617 (N_3617,N_3598,N_3592);
and U3618 (N_3618,N_3568,N_3558);
nor U3619 (N_3619,N_3574,N_3562);
and U3620 (N_3620,N_3516,N_3542);
and U3621 (N_3621,N_3512,N_3506);
nand U3622 (N_3622,N_3555,N_3543);
or U3623 (N_3623,N_3521,N_3580);
and U3624 (N_3624,N_3534,N_3551);
nand U3625 (N_3625,N_3522,N_3535);
xor U3626 (N_3626,N_3597,N_3500);
and U3627 (N_3627,N_3540,N_3583);
nor U3628 (N_3628,N_3554,N_3523);
nand U3629 (N_3629,N_3596,N_3572);
nor U3630 (N_3630,N_3577,N_3546);
nor U3631 (N_3631,N_3599,N_3502);
and U3632 (N_3632,N_3536,N_3524);
nand U3633 (N_3633,N_3544,N_3552);
nor U3634 (N_3634,N_3532,N_3513);
and U3635 (N_3635,N_3578,N_3514);
or U3636 (N_3636,N_3520,N_3575);
nor U3637 (N_3637,N_3533,N_3550);
and U3638 (N_3638,N_3595,N_3503);
nand U3639 (N_3639,N_3557,N_3519);
nor U3640 (N_3640,N_3541,N_3585);
nand U3641 (N_3641,N_3584,N_3545);
nor U3642 (N_3642,N_3530,N_3515);
nor U3643 (N_3643,N_3594,N_3553);
or U3644 (N_3644,N_3510,N_3573);
xnor U3645 (N_3645,N_3565,N_3509);
and U3646 (N_3646,N_3593,N_3527);
nor U3647 (N_3647,N_3582,N_3591);
or U3648 (N_3648,N_3571,N_3569);
nor U3649 (N_3649,N_3590,N_3517);
nor U3650 (N_3650,N_3517,N_3521);
or U3651 (N_3651,N_3568,N_3556);
and U3652 (N_3652,N_3556,N_3513);
nand U3653 (N_3653,N_3528,N_3512);
nand U3654 (N_3654,N_3569,N_3511);
nand U3655 (N_3655,N_3510,N_3506);
or U3656 (N_3656,N_3590,N_3586);
nor U3657 (N_3657,N_3513,N_3500);
nor U3658 (N_3658,N_3556,N_3519);
and U3659 (N_3659,N_3531,N_3563);
or U3660 (N_3660,N_3509,N_3503);
or U3661 (N_3661,N_3557,N_3522);
xnor U3662 (N_3662,N_3534,N_3548);
nand U3663 (N_3663,N_3596,N_3578);
and U3664 (N_3664,N_3538,N_3505);
and U3665 (N_3665,N_3563,N_3500);
or U3666 (N_3666,N_3590,N_3595);
and U3667 (N_3667,N_3564,N_3526);
or U3668 (N_3668,N_3571,N_3500);
or U3669 (N_3669,N_3539,N_3570);
nand U3670 (N_3670,N_3551,N_3595);
nor U3671 (N_3671,N_3572,N_3516);
nand U3672 (N_3672,N_3500,N_3530);
nor U3673 (N_3673,N_3558,N_3513);
and U3674 (N_3674,N_3542,N_3505);
or U3675 (N_3675,N_3562,N_3500);
and U3676 (N_3676,N_3568,N_3587);
nand U3677 (N_3677,N_3527,N_3557);
nor U3678 (N_3678,N_3510,N_3549);
and U3679 (N_3679,N_3561,N_3574);
nand U3680 (N_3680,N_3520,N_3557);
and U3681 (N_3681,N_3516,N_3579);
nor U3682 (N_3682,N_3542,N_3536);
nand U3683 (N_3683,N_3599,N_3523);
nand U3684 (N_3684,N_3583,N_3542);
nand U3685 (N_3685,N_3581,N_3520);
nand U3686 (N_3686,N_3572,N_3552);
or U3687 (N_3687,N_3516,N_3550);
and U3688 (N_3688,N_3515,N_3532);
nor U3689 (N_3689,N_3541,N_3531);
nand U3690 (N_3690,N_3517,N_3561);
nor U3691 (N_3691,N_3544,N_3514);
and U3692 (N_3692,N_3578,N_3552);
and U3693 (N_3693,N_3579,N_3545);
nor U3694 (N_3694,N_3526,N_3506);
and U3695 (N_3695,N_3574,N_3575);
nand U3696 (N_3696,N_3545,N_3519);
nand U3697 (N_3697,N_3585,N_3502);
and U3698 (N_3698,N_3530,N_3540);
or U3699 (N_3699,N_3568,N_3549);
and U3700 (N_3700,N_3601,N_3692);
nor U3701 (N_3701,N_3629,N_3696);
or U3702 (N_3702,N_3603,N_3663);
nor U3703 (N_3703,N_3690,N_3619);
or U3704 (N_3704,N_3666,N_3693);
and U3705 (N_3705,N_3644,N_3625);
nand U3706 (N_3706,N_3686,N_3639);
nor U3707 (N_3707,N_3646,N_3679);
xor U3708 (N_3708,N_3650,N_3635);
nor U3709 (N_3709,N_3617,N_3614);
nand U3710 (N_3710,N_3685,N_3630);
or U3711 (N_3711,N_3682,N_3645);
and U3712 (N_3712,N_3678,N_3660);
or U3713 (N_3713,N_3640,N_3615);
nand U3714 (N_3714,N_3602,N_3609);
nand U3715 (N_3715,N_3659,N_3622);
and U3716 (N_3716,N_3699,N_3676);
xnor U3717 (N_3717,N_3626,N_3611);
or U3718 (N_3718,N_3612,N_3616);
and U3719 (N_3719,N_3687,N_3671);
nor U3720 (N_3720,N_3642,N_3621);
nor U3721 (N_3721,N_3655,N_3653);
nand U3722 (N_3722,N_3641,N_3689);
and U3723 (N_3723,N_3667,N_3652);
nor U3724 (N_3724,N_3684,N_3634);
nor U3725 (N_3725,N_3680,N_3638);
nor U3726 (N_3726,N_3688,N_3698);
nand U3727 (N_3727,N_3632,N_3669);
or U3728 (N_3728,N_3600,N_3604);
or U3729 (N_3729,N_3610,N_3647);
nor U3730 (N_3730,N_3683,N_3636);
xor U3731 (N_3731,N_3651,N_3658);
and U3732 (N_3732,N_3670,N_3605);
or U3733 (N_3733,N_3627,N_3620);
and U3734 (N_3734,N_3668,N_3695);
xnor U3735 (N_3735,N_3674,N_3633);
or U3736 (N_3736,N_3656,N_3694);
nand U3737 (N_3737,N_3665,N_3662);
nor U3738 (N_3738,N_3628,N_3637);
or U3739 (N_3739,N_3661,N_3697);
or U3740 (N_3740,N_3681,N_3664);
or U3741 (N_3741,N_3649,N_3657);
xor U3742 (N_3742,N_3654,N_3673);
nand U3743 (N_3743,N_3648,N_3608);
nor U3744 (N_3744,N_3631,N_3675);
nand U3745 (N_3745,N_3618,N_3623);
or U3746 (N_3746,N_3677,N_3691);
nor U3747 (N_3747,N_3607,N_3672);
nor U3748 (N_3748,N_3643,N_3613);
or U3749 (N_3749,N_3606,N_3624);
and U3750 (N_3750,N_3690,N_3695);
or U3751 (N_3751,N_3612,N_3602);
and U3752 (N_3752,N_3608,N_3669);
or U3753 (N_3753,N_3668,N_3680);
or U3754 (N_3754,N_3649,N_3687);
nand U3755 (N_3755,N_3697,N_3674);
and U3756 (N_3756,N_3695,N_3672);
xor U3757 (N_3757,N_3621,N_3638);
and U3758 (N_3758,N_3690,N_3605);
or U3759 (N_3759,N_3678,N_3600);
xor U3760 (N_3760,N_3675,N_3643);
xnor U3761 (N_3761,N_3606,N_3601);
nor U3762 (N_3762,N_3667,N_3644);
xnor U3763 (N_3763,N_3622,N_3608);
nand U3764 (N_3764,N_3666,N_3607);
xor U3765 (N_3765,N_3665,N_3691);
nor U3766 (N_3766,N_3698,N_3646);
and U3767 (N_3767,N_3607,N_3699);
and U3768 (N_3768,N_3664,N_3643);
nand U3769 (N_3769,N_3610,N_3654);
or U3770 (N_3770,N_3612,N_3637);
and U3771 (N_3771,N_3632,N_3607);
and U3772 (N_3772,N_3647,N_3681);
nand U3773 (N_3773,N_3670,N_3600);
nand U3774 (N_3774,N_3696,N_3686);
and U3775 (N_3775,N_3688,N_3683);
and U3776 (N_3776,N_3637,N_3608);
nor U3777 (N_3777,N_3662,N_3657);
nor U3778 (N_3778,N_3689,N_3615);
and U3779 (N_3779,N_3601,N_3634);
or U3780 (N_3780,N_3658,N_3640);
nor U3781 (N_3781,N_3615,N_3675);
nor U3782 (N_3782,N_3655,N_3679);
nand U3783 (N_3783,N_3639,N_3668);
and U3784 (N_3784,N_3653,N_3682);
nor U3785 (N_3785,N_3677,N_3652);
or U3786 (N_3786,N_3671,N_3626);
and U3787 (N_3787,N_3609,N_3699);
xnor U3788 (N_3788,N_3683,N_3637);
and U3789 (N_3789,N_3664,N_3665);
nand U3790 (N_3790,N_3630,N_3635);
and U3791 (N_3791,N_3615,N_3695);
and U3792 (N_3792,N_3624,N_3691);
nand U3793 (N_3793,N_3615,N_3610);
nor U3794 (N_3794,N_3683,N_3690);
xor U3795 (N_3795,N_3694,N_3616);
nand U3796 (N_3796,N_3619,N_3660);
xnor U3797 (N_3797,N_3662,N_3652);
nand U3798 (N_3798,N_3665,N_3685);
nor U3799 (N_3799,N_3643,N_3603);
nand U3800 (N_3800,N_3732,N_3751);
xor U3801 (N_3801,N_3725,N_3737);
or U3802 (N_3802,N_3704,N_3774);
nand U3803 (N_3803,N_3759,N_3717);
nand U3804 (N_3804,N_3753,N_3784);
nor U3805 (N_3805,N_3734,N_3716);
nand U3806 (N_3806,N_3785,N_3703);
and U3807 (N_3807,N_3798,N_3792);
nor U3808 (N_3808,N_3773,N_3711);
and U3809 (N_3809,N_3793,N_3768);
nor U3810 (N_3810,N_3743,N_3763);
and U3811 (N_3811,N_3740,N_3714);
or U3812 (N_3812,N_3718,N_3720);
or U3813 (N_3813,N_3735,N_3701);
nand U3814 (N_3814,N_3777,N_3754);
and U3815 (N_3815,N_3772,N_3721);
nand U3816 (N_3816,N_3702,N_3788);
xnor U3817 (N_3817,N_3797,N_3766);
or U3818 (N_3818,N_3700,N_3762);
or U3819 (N_3819,N_3731,N_3713);
xor U3820 (N_3820,N_3765,N_3769);
nand U3821 (N_3821,N_3715,N_3787);
xor U3822 (N_3822,N_3757,N_3761);
nand U3823 (N_3823,N_3747,N_3707);
nor U3824 (N_3824,N_3723,N_3730);
nor U3825 (N_3825,N_3775,N_3745);
or U3826 (N_3826,N_3764,N_3779);
nor U3827 (N_3827,N_3750,N_3780);
and U3828 (N_3828,N_3771,N_3719);
or U3829 (N_3829,N_3708,N_3712);
or U3830 (N_3830,N_3739,N_3755);
xnor U3831 (N_3831,N_3749,N_3795);
nor U3832 (N_3832,N_3786,N_3776);
xnor U3833 (N_3833,N_3783,N_3778);
or U3834 (N_3834,N_3741,N_3724);
and U3835 (N_3835,N_3733,N_3729);
nor U3836 (N_3836,N_3727,N_3790);
nand U3837 (N_3837,N_3742,N_3706);
and U3838 (N_3838,N_3736,N_3726);
nor U3839 (N_3839,N_3760,N_3710);
or U3840 (N_3840,N_3799,N_3748);
and U3841 (N_3841,N_3781,N_3709);
or U3842 (N_3842,N_3738,N_3746);
and U3843 (N_3843,N_3752,N_3789);
xnor U3844 (N_3844,N_3770,N_3744);
or U3845 (N_3845,N_3728,N_3796);
xor U3846 (N_3846,N_3722,N_3782);
nand U3847 (N_3847,N_3756,N_3758);
nand U3848 (N_3848,N_3794,N_3791);
and U3849 (N_3849,N_3767,N_3705);
and U3850 (N_3850,N_3727,N_3754);
or U3851 (N_3851,N_3711,N_3729);
or U3852 (N_3852,N_3704,N_3794);
nand U3853 (N_3853,N_3736,N_3776);
and U3854 (N_3854,N_3719,N_3752);
nand U3855 (N_3855,N_3797,N_3742);
and U3856 (N_3856,N_3788,N_3781);
and U3857 (N_3857,N_3718,N_3787);
xor U3858 (N_3858,N_3772,N_3791);
nand U3859 (N_3859,N_3701,N_3758);
nor U3860 (N_3860,N_3796,N_3731);
nand U3861 (N_3861,N_3751,N_3731);
nor U3862 (N_3862,N_3767,N_3791);
and U3863 (N_3863,N_3768,N_3720);
nor U3864 (N_3864,N_3729,N_3707);
and U3865 (N_3865,N_3786,N_3714);
and U3866 (N_3866,N_3740,N_3780);
xor U3867 (N_3867,N_3708,N_3734);
and U3868 (N_3868,N_3766,N_3743);
and U3869 (N_3869,N_3774,N_3763);
nand U3870 (N_3870,N_3739,N_3762);
and U3871 (N_3871,N_3776,N_3717);
or U3872 (N_3872,N_3748,N_3776);
nor U3873 (N_3873,N_3723,N_3777);
or U3874 (N_3874,N_3711,N_3795);
nor U3875 (N_3875,N_3750,N_3792);
and U3876 (N_3876,N_3761,N_3738);
nor U3877 (N_3877,N_3761,N_3781);
or U3878 (N_3878,N_3771,N_3791);
and U3879 (N_3879,N_3717,N_3785);
nand U3880 (N_3880,N_3749,N_3757);
nor U3881 (N_3881,N_3750,N_3784);
and U3882 (N_3882,N_3751,N_3776);
or U3883 (N_3883,N_3723,N_3785);
xor U3884 (N_3884,N_3773,N_3736);
or U3885 (N_3885,N_3729,N_3725);
and U3886 (N_3886,N_3746,N_3752);
and U3887 (N_3887,N_3762,N_3794);
nor U3888 (N_3888,N_3762,N_3745);
xnor U3889 (N_3889,N_3708,N_3709);
and U3890 (N_3890,N_3742,N_3788);
or U3891 (N_3891,N_3727,N_3775);
nand U3892 (N_3892,N_3723,N_3778);
nand U3893 (N_3893,N_3720,N_3799);
or U3894 (N_3894,N_3720,N_3760);
and U3895 (N_3895,N_3717,N_3732);
nand U3896 (N_3896,N_3780,N_3795);
nand U3897 (N_3897,N_3757,N_3737);
and U3898 (N_3898,N_3712,N_3755);
and U3899 (N_3899,N_3740,N_3760);
and U3900 (N_3900,N_3825,N_3894);
and U3901 (N_3901,N_3892,N_3861);
xor U3902 (N_3902,N_3805,N_3829);
nand U3903 (N_3903,N_3804,N_3899);
xor U3904 (N_3904,N_3814,N_3832);
or U3905 (N_3905,N_3890,N_3860);
or U3906 (N_3906,N_3809,N_3867);
xnor U3907 (N_3907,N_3803,N_3807);
and U3908 (N_3908,N_3883,N_3834);
nand U3909 (N_3909,N_3877,N_3823);
and U3910 (N_3910,N_3887,N_3884);
nand U3911 (N_3911,N_3872,N_3839);
nor U3912 (N_3912,N_3878,N_3830);
or U3913 (N_3913,N_3857,N_3876);
or U3914 (N_3914,N_3855,N_3879);
and U3915 (N_3915,N_3808,N_3874);
or U3916 (N_3916,N_3816,N_3800);
or U3917 (N_3917,N_3858,N_3862);
nand U3918 (N_3918,N_3806,N_3838);
xor U3919 (N_3919,N_3870,N_3851);
or U3920 (N_3920,N_3801,N_3813);
nor U3921 (N_3921,N_3875,N_3835);
or U3922 (N_3922,N_3827,N_3895);
and U3923 (N_3923,N_3869,N_3837);
or U3924 (N_3924,N_3882,N_3811);
and U3925 (N_3925,N_3856,N_3889);
and U3926 (N_3926,N_3810,N_3886);
or U3927 (N_3927,N_3819,N_3897);
nand U3928 (N_3928,N_3844,N_3843);
or U3929 (N_3929,N_3893,N_3896);
nor U3930 (N_3930,N_3802,N_3868);
nor U3931 (N_3931,N_3847,N_3865);
or U3932 (N_3932,N_3812,N_3871);
or U3933 (N_3933,N_3820,N_3888);
nand U3934 (N_3934,N_3898,N_3822);
and U3935 (N_3935,N_3840,N_3831);
or U3936 (N_3936,N_3815,N_3845);
nand U3937 (N_3937,N_3853,N_3891);
or U3938 (N_3938,N_3852,N_3866);
or U3939 (N_3939,N_3850,N_3846);
nand U3940 (N_3940,N_3836,N_3854);
nand U3941 (N_3941,N_3881,N_3817);
or U3942 (N_3942,N_3864,N_3826);
xor U3943 (N_3943,N_3818,N_3821);
nor U3944 (N_3944,N_3880,N_3833);
and U3945 (N_3945,N_3859,N_3885);
or U3946 (N_3946,N_3841,N_3863);
xnor U3947 (N_3947,N_3849,N_3824);
nand U3948 (N_3948,N_3848,N_3828);
and U3949 (N_3949,N_3842,N_3873);
and U3950 (N_3950,N_3810,N_3802);
and U3951 (N_3951,N_3801,N_3826);
and U3952 (N_3952,N_3892,N_3811);
nand U3953 (N_3953,N_3854,N_3803);
and U3954 (N_3954,N_3803,N_3839);
and U3955 (N_3955,N_3846,N_3890);
xnor U3956 (N_3956,N_3839,N_3876);
nand U3957 (N_3957,N_3898,N_3870);
or U3958 (N_3958,N_3835,N_3812);
and U3959 (N_3959,N_3866,N_3887);
nor U3960 (N_3960,N_3821,N_3857);
nand U3961 (N_3961,N_3870,N_3869);
nand U3962 (N_3962,N_3832,N_3820);
and U3963 (N_3963,N_3899,N_3818);
and U3964 (N_3964,N_3839,N_3810);
nand U3965 (N_3965,N_3848,N_3844);
or U3966 (N_3966,N_3811,N_3881);
or U3967 (N_3967,N_3847,N_3886);
and U3968 (N_3968,N_3814,N_3863);
nor U3969 (N_3969,N_3822,N_3843);
or U3970 (N_3970,N_3852,N_3818);
and U3971 (N_3971,N_3825,N_3861);
or U3972 (N_3972,N_3831,N_3815);
nor U3973 (N_3973,N_3823,N_3825);
nand U3974 (N_3974,N_3857,N_3818);
and U3975 (N_3975,N_3845,N_3807);
or U3976 (N_3976,N_3879,N_3887);
nor U3977 (N_3977,N_3869,N_3881);
or U3978 (N_3978,N_3840,N_3898);
or U3979 (N_3979,N_3844,N_3806);
nor U3980 (N_3980,N_3861,N_3838);
or U3981 (N_3981,N_3827,N_3851);
nand U3982 (N_3982,N_3828,N_3880);
or U3983 (N_3983,N_3876,N_3885);
or U3984 (N_3984,N_3886,N_3877);
and U3985 (N_3985,N_3852,N_3804);
nor U3986 (N_3986,N_3832,N_3872);
xor U3987 (N_3987,N_3855,N_3821);
xor U3988 (N_3988,N_3861,N_3818);
nor U3989 (N_3989,N_3867,N_3839);
xnor U3990 (N_3990,N_3853,N_3807);
nand U3991 (N_3991,N_3854,N_3896);
nor U3992 (N_3992,N_3824,N_3822);
nand U3993 (N_3993,N_3871,N_3890);
and U3994 (N_3994,N_3821,N_3810);
and U3995 (N_3995,N_3838,N_3840);
xnor U3996 (N_3996,N_3850,N_3866);
nor U3997 (N_3997,N_3823,N_3889);
nor U3998 (N_3998,N_3882,N_3836);
nand U3999 (N_3999,N_3816,N_3851);
nand U4000 (N_4000,N_3993,N_3938);
or U4001 (N_4001,N_3943,N_3963);
or U4002 (N_4002,N_3957,N_3948);
or U4003 (N_4003,N_3934,N_3964);
nand U4004 (N_4004,N_3940,N_3924);
or U4005 (N_4005,N_3992,N_3962);
or U4006 (N_4006,N_3945,N_3904);
and U4007 (N_4007,N_3985,N_3961);
nor U4008 (N_4008,N_3929,N_3920);
nor U4009 (N_4009,N_3944,N_3967);
nand U4010 (N_4010,N_3995,N_3950);
or U4011 (N_4011,N_3931,N_3956);
or U4012 (N_4012,N_3901,N_3921);
nor U4013 (N_4013,N_3973,N_3927);
nor U4014 (N_4014,N_3959,N_3988);
or U4015 (N_4015,N_3926,N_3905);
nor U4016 (N_4016,N_3968,N_3946);
nor U4017 (N_4017,N_3928,N_3994);
or U4018 (N_4018,N_3980,N_3936);
nand U4019 (N_4019,N_3941,N_3979);
nand U4020 (N_4020,N_3977,N_3982);
nand U4021 (N_4021,N_3999,N_3912);
and U4022 (N_4022,N_3908,N_3939);
nor U4023 (N_4023,N_3965,N_3933);
nor U4024 (N_4024,N_3917,N_3906);
and U4025 (N_4025,N_3997,N_3996);
xor U4026 (N_4026,N_3932,N_3969);
or U4027 (N_4027,N_3974,N_3998);
nand U4028 (N_4028,N_3970,N_3925);
and U4029 (N_4029,N_3910,N_3989);
or U4030 (N_4030,N_3990,N_3955);
nand U4031 (N_4031,N_3986,N_3958);
nor U4032 (N_4032,N_3942,N_3952);
and U4033 (N_4033,N_3915,N_3902);
and U4034 (N_4034,N_3975,N_3923);
nor U4035 (N_4035,N_3900,N_3971);
and U4036 (N_4036,N_3951,N_3913);
nand U4037 (N_4037,N_3978,N_3907);
or U4038 (N_4038,N_3914,N_3937);
nand U4039 (N_4039,N_3903,N_3953);
nor U4040 (N_4040,N_3981,N_3991);
and U4041 (N_4041,N_3930,N_3983);
and U4042 (N_4042,N_3987,N_3935);
and U4043 (N_4043,N_3918,N_3919);
or U4044 (N_4044,N_3972,N_3954);
and U4045 (N_4045,N_3984,N_3922);
or U4046 (N_4046,N_3976,N_3949);
nand U4047 (N_4047,N_3916,N_3947);
nand U4048 (N_4048,N_3966,N_3909);
nand U4049 (N_4049,N_3960,N_3911);
xor U4050 (N_4050,N_3986,N_3999);
nand U4051 (N_4051,N_3959,N_3917);
nand U4052 (N_4052,N_3961,N_3997);
xnor U4053 (N_4053,N_3928,N_3952);
or U4054 (N_4054,N_3957,N_3932);
and U4055 (N_4055,N_3981,N_3949);
nand U4056 (N_4056,N_3994,N_3915);
nand U4057 (N_4057,N_3929,N_3982);
or U4058 (N_4058,N_3955,N_3998);
or U4059 (N_4059,N_3973,N_3996);
or U4060 (N_4060,N_3986,N_3941);
nand U4061 (N_4061,N_3976,N_3974);
nand U4062 (N_4062,N_3989,N_3968);
xor U4063 (N_4063,N_3924,N_3964);
or U4064 (N_4064,N_3971,N_3967);
nor U4065 (N_4065,N_3936,N_3918);
xnor U4066 (N_4066,N_3992,N_3941);
nand U4067 (N_4067,N_3910,N_3948);
and U4068 (N_4068,N_3901,N_3905);
and U4069 (N_4069,N_3938,N_3948);
xor U4070 (N_4070,N_3989,N_3973);
or U4071 (N_4071,N_3923,N_3928);
nand U4072 (N_4072,N_3984,N_3919);
nor U4073 (N_4073,N_3908,N_3900);
nor U4074 (N_4074,N_3952,N_3968);
nor U4075 (N_4075,N_3935,N_3952);
nand U4076 (N_4076,N_3972,N_3915);
nor U4077 (N_4077,N_3933,N_3938);
nor U4078 (N_4078,N_3949,N_3980);
xnor U4079 (N_4079,N_3953,N_3927);
nor U4080 (N_4080,N_3991,N_3975);
nor U4081 (N_4081,N_3932,N_3909);
and U4082 (N_4082,N_3911,N_3901);
nor U4083 (N_4083,N_3997,N_3953);
nor U4084 (N_4084,N_3914,N_3941);
nand U4085 (N_4085,N_3954,N_3927);
nand U4086 (N_4086,N_3975,N_3996);
nand U4087 (N_4087,N_3915,N_3923);
nand U4088 (N_4088,N_3964,N_3925);
or U4089 (N_4089,N_3960,N_3984);
and U4090 (N_4090,N_3999,N_3981);
nand U4091 (N_4091,N_3949,N_3909);
nor U4092 (N_4092,N_3920,N_3939);
nand U4093 (N_4093,N_3962,N_3917);
and U4094 (N_4094,N_3918,N_3954);
nand U4095 (N_4095,N_3928,N_3916);
and U4096 (N_4096,N_3954,N_3977);
and U4097 (N_4097,N_3983,N_3918);
and U4098 (N_4098,N_3970,N_3951);
xnor U4099 (N_4099,N_3941,N_3933);
nor U4100 (N_4100,N_4031,N_4090);
nand U4101 (N_4101,N_4034,N_4033);
or U4102 (N_4102,N_4015,N_4027);
nand U4103 (N_4103,N_4045,N_4057);
and U4104 (N_4104,N_4020,N_4092);
nor U4105 (N_4105,N_4017,N_4066);
xnor U4106 (N_4106,N_4003,N_4049);
nor U4107 (N_4107,N_4052,N_4075);
nor U4108 (N_4108,N_4094,N_4098);
and U4109 (N_4109,N_4018,N_4064);
or U4110 (N_4110,N_4035,N_4029);
nor U4111 (N_4111,N_4096,N_4089);
nand U4112 (N_4112,N_4056,N_4065);
nand U4113 (N_4113,N_4051,N_4070);
nand U4114 (N_4114,N_4022,N_4059);
and U4115 (N_4115,N_4000,N_4080);
nand U4116 (N_4116,N_4006,N_4001);
nor U4117 (N_4117,N_4041,N_4055);
nor U4118 (N_4118,N_4014,N_4009);
nor U4119 (N_4119,N_4082,N_4058);
nor U4120 (N_4120,N_4093,N_4077);
xnor U4121 (N_4121,N_4071,N_4043);
nor U4122 (N_4122,N_4028,N_4091);
or U4123 (N_4123,N_4078,N_4030);
nand U4124 (N_4124,N_4004,N_4061);
xnor U4125 (N_4125,N_4087,N_4074);
nand U4126 (N_4126,N_4069,N_4016);
nor U4127 (N_4127,N_4086,N_4042);
and U4128 (N_4128,N_4005,N_4054);
nor U4129 (N_4129,N_4036,N_4010);
nor U4130 (N_4130,N_4079,N_4012);
nor U4131 (N_4131,N_4060,N_4047);
and U4132 (N_4132,N_4068,N_4099);
nor U4133 (N_4133,N_4038,N_4050);
and U4134 (N_4134,N_4083,N_4067);
and U4135 (N_4135,N_4025,N_4019);
nand U4136 (N_4136,N_4076,N_4008);
nor U4137 (N_4137,N_4088,N_4026);
nor U4138 (N_4138,N_4039,N_4081);
and U4139 (N_4139,N_4023,N_4046);
nand U4140 (N_4140,N_4063,N_4073);
or U4141 (N_4141,N_4024,N_4021);
and U4142 (N_4142,N_4007,N_4084);
or U4143 (N_4143,N_4053,N_4072);
nand U4144 (N_4144,N_4037,N_4044);
or U4145 (N_4145,N_4032,N_4048);
and U4146 (N_4146,N_4097,N_4040);
and U4147 (N_4147,N_4062,N_4002);
nor U4148 (N_4148,N_4085,N_4011);
nand U4149 (N_4149,N_4013,N_4095);
nor U4150 (N_4150,N_4045,N_4033);
or U4151 (N_4151,N_4096,N_4049);
nand U4152 (N_4152,N_4043,N_4087);
and U4153 (N_4153,N_4099,N_4055);
xnor U4154 (N_4154,N_4084,N_4041);
and U4155 (N_4155,N_4002,N_4047);
nor U4156 (N_4156,N_4050,N_4058);
or U4157 (N_4157,N_4012,N_4051);
or U4158 (N_4158,N_4097,N_4079);
nand U4159 (N_4159,N_4097,N_4010);
nand U4160 (N_4160,N_4034,N_4072);
nand U4161 (N_4161,N_4057,N_4020);
nand U4162 (N_4162,N_4074,N_4011);
or U4163 (N_4163,N_4030,N_4033);
nand U4164 (N_4164,N_4058,N_4089);
and U4165 (N_4165,N_4098,N_4030);
and U4166 (N_4166,N_4048,N_4009);
nor U4167 (N_4167,N_4077,N_4021);
nand U4168 (N_4168,N_4044,N_4009);
xor U4169 (N_4169,N_4016,N_4079);
nor U4170 (N_4170,N_4059,N_4097);
xor U4171 (N_4171,N_4016,N_4045);
or U4172 (N_4172,N_4086,N_4097);
nand U4173 (N_4173,N_4034,N_4064);
and U4174 (N_4174,N_4027,N_4032);
nor U4175 (N_4175,N_4021,N_4045);
and U4176 (N_4176,N_4001,N_4021);
xnor U4177 (N_4177,N_4091,N_4097);
nor U4178 (N_4178,N_4057,N_4076);
and U4179 (N_4179,N_4008,N_4039);
and U4180 (N_4180,N_4029,N_4025);
nand U4181 (N_4181,N_4088,N_4047);
nand U4182 (N_4182,N_4079,N_4017);
or U4183 (N_4183,N_4067,N_4095);
or U4184 (N_4184,N_4070,N_4031);
nand U4185 (N_4185,N_4025,N_4018);
nand U4186 (N_4186,N_4045,N_4066);
xor U4187 (N_4187,N_4061,N_4063);
nor U4188 (N_4188,N_4004,N_4024);
nand U4189 (N_4189,N_4076,N_4027);
or U4190 (N_4190,N_4072,N_4061);
or U4191 (N_4191,N_4057,N_4093);
and U4192 (N_4192,N_4019,N_4028);
and U4193 (N_4193,N_4020,N_4053);
nor U4194 (N_4194,N_4060,N_4042);
nor U4195 (N_4195,N_4076,N_4043);
or U4196 (N_4196,N_4087,N_4067);
nor U4197 (N_4197,N_4091,N_4083);
nand U4198 (N_4198,N_4081,N_4052);
or U4199 (N_4199,N_4002,N_4086);
or U4200 (N_4200,N_4199,N_4195);
or U4201 (N_4201,N_4167,N_4134);
nor U4202 (N_4202,N_4100,N_4156);
nand U4203 (N_4203,N_4107,N_4111);
xor U4204 (N_4204,N_4154,N_4109);
nor U4205 (N_4205,N_4191,N_4184);
and U4206 (N_4206,N_4139,N_4135);
nor U4207 (N_4207,N_4143,N_4130);
nand U4208 (N_4208,N_4123,N_4157);
nand U4209 (N_4209,N_4128,N_4122);
xor U4210 (N_4210,N_4155,N_4147);
and U4211 (N_4211,N_4161,N_4106);
or U4212 (N_4212,N_4102,N_4112);
xnor U4213 (N_4213,N_4133,N_4163);
nand U4214 (N_4214,N_4182,N_4117);
and U4215 (N_4215,N_4183,N_4185);
nand U4216 (N_4216,N_4108,N_4137);
nor U4217 (N_4217,N_4170,N_4110);
or U4218 (N_4218,N_4101,N_4190);
nand U4219 (N_4219,N_4150,N_4164);
and U4220 (N_4220,N_4198,N_4169);
and U4221 (N_4221,N_4151,N_4196);
nor U4222 (N_4222,N_4126,N_4166);
and U4223 (N_4223,N_4132,N_4116);
and U4224 (N_4224,N_4175,N_4189);
xor U4225 (N_4225,N_4168,N_4146);
and U4226 (N_4226,N_4193,N_4121);
or U4227 (N_4227,N_4173,N_4174);
or U4228 (N_4228,N_4152,N_4165);
xnor U4229 (N_4229,N_4188,N_4142);
or U4230 (N_4230,N_4172,N_4124);
xnor U4231 (N_4231,N_4158,N_4118);
nor U4232 (N_4232,N_4127,N_4171);
nand U4233 (N_4233,N_4138,N_4114);
xnor U4234 (N_4234,N_4197,N_4160);
nand U4235 (N_4235,N_4179,N_4145);
nand U4236 (N_4236,N_4105,N_4176);
and U4237 (N_4237,N_4148,N_4192);
or U4238 (N_4238,N_4125,N_4194);
nor U4239 (N_4239,N_4113,N_4141);
nor U4240 (N_4240,N_4120,N_4149);
nor U4241 (N_4241,N_4177,N_4115);
or U4242 (N_4242,N_4186,N_4103);
or U4243 (N_4243,N_4153,N_4136);
and U4244 (N_4244,N_4162,N_4104);
xnor U4245 (N_4245,N_4119,N_4144);
or U4246 (N_4246,N_4131,N_4129);
nor U4247 (N_4247,N_4159,N_4187);
nand U4248 (N_4248,N_4178,N_4180);
xor U4249 (N_4249,N_4181,N_4140);
and U4250 (N_4250,N_4142,N_4128);
xor U4251 (N_4251,N_4189,N_4121);
nor U4252 (N_4252,N_4185,N_4140);
nand U4253 (N_4253,N_4135,N_4103);
nand U4254 (N_4254,N_4148,N_4197);
and U4255 (N_4255,N_4183,N_4192);
and U4256 (N_4256,N_4156,N_4141);
and U4257 (N_4257,N_4145,N_4146);
and U4258 (N_4258,N_4133,N_4192);
nor U4259 (N_4259,N_4101,N_4149);
or U4260 (N_4260,N_4182,N_4161);
or U4261 (N_4261,N_4175,N_4122);
and U4262 (N_4262,N_4199,N_4133);
xnor U4263 (N_4263,N_4142,N_4190);
nor U4264 (N_4264,N_4179,N_4103);
nor U4265 (N_4265,N_4138,N_4136);
nand U4266 (N_4266,N_4167,N_4124);
and U4267 (N_4267,N_4122,N_4126);
and U4268 (N_4268,N_4129,N_4166);
or U4269 (N_4269,N_4105,N_4157);
nand U4270 (N_4270,N_4152,N_4186);
xnor U4271 (N_4271,N_4108,N_4162);
and U4272 (N_4272,N_4159,N_4162);
or U4273 (N_4273,N_4111,N_4178);
and U4274 (N_4274,N_4169,N_4159);
nand U4275 (N_4275,N_4120,N_4155);
or U4276 (N_4276,N_4175,N_4132);
and U4277 (N_4277,N_4184,N_4189);
nand U4278 (N_4278,N_4156,N_4159);
nor U4279 (N_4279,N_4175,N_4147);
xnor U4280 (N_4280,N_4117,N_4141);
and U4281 (N_4281,N_4129,N_4105);
or U4282 (N_4282,N_4184,N_4105);
xnor U4283 (N_4283,N_4189,N_4130);
nand U4284 (N_4284,N_4137,N_4105);
nor U4285 (N_4285,N_4130,N_4113);
nor U4286 (N_4286,N_4184,N_4148);
nand U4287 (N_4287,N_4102,N_4127);
and U4288 (N_4288,N_4119,N_4190);
or U4289 (N_4289,N_4108,N_4112);
xnor U4290 (N_4290,N_4155,N_4196);
nor U4291 (N_4291,N_4122,N_4168);
nand U4292 (N_4292,N_4135,N_4104);
or U4293 (N_4293,N_4151,N_4173);
and U4294 (N_4294,N_4127,N_4196);
and U4295 (N_4295,N_4140,N_4126);
or U4296 (N_4296,N_4166,N_4122);
nand U4297 (N_4297,N_4133,N_4174);
xor U4298 (N_4298,N_4166,N_4106);
xnor U4299 (N_4299,N_4159,N_4185);
nor U4300 (N_4300,N_4245,N_4221);
nor U4301 (N_4301,N_4213,N_4295);
and U4302 (N_4302,N_4210,N_4226);
nor U4303 (N_4303,N_4260,N_4218);
nand U4304 (N_4304,N_4264,N_4228);
or U4305 (N_4305,N_4238,N_4263);
nand U4306 (N_4306,N_4256,N_4271);
and U4307 (N_4307,N_4244,N_4243);
xor U4308 (N_4308,N_4273,N_4266);
and U4309 (N_4309,N_4223,N_4270);
nand U4310 (N_4310,N_4209,N_4251);
nor U4311 (N_4311,N_4235,N_4233);
and U4312 (N_4312,N_4275,N_4222);
nor U4313 (N_4313,N_4202,N_4237);
or U4314 (N_4314,N_4211,N_4299);
and U4315 (N_4315,N_4239,N_4288);
and U4316 (N_4316,N_4284,N_4296);
nand U4317 (N_4317,N_4293,N_4272);
xnor U4318 (N_4318,N_4246,N_4280);
and U4319 (N_4319,N_4200,N_4217);
and U4320 (N_4320,N_4206,N_4247);
nand U4321 (N_4321,N_4208,N_4279);
nand U4322 (N_4322,N_4281,N_4220);
nand U4323 (N_4323,N_4276,N_4240);
and U4324 (N_4324,N_4250,N_4259);
nor U4325 (N_4325,N_4249,N_4292);
and U4326 (N_4326,N_4278,N_4229);
or U4327 (N_4327,N_4262,N_4214);
or U4328 (N_4328,N_4212,N_4285);
or U4329 (N_4329,N_4289,N_4231);
nor U4330 (N_4330,N_4267,N_4290);
or U4331 (N_4331,N_4282,N_4242);
nand U4332 (N_4332,N_4287,N_4207);
xnor U4333 (N_4333,N_4286,N_4274);
nor U4334 (N_4334,N_4234,N_4261);
or U4335 (N_4335,N_4241,N_4201);
or U4336 (N_4336,N_4204,N_4291);
or U4337 (N_4337,N_4283,N_4248);
nor U4338 (N_4338,N_4227,N_4236);
or U4339 (N_4339,N_4265,N_4203);
and U4340 (N_4340,N_4297,N_4224);
nand U4341 (N_4341,N_4294,N_4219);
or U4342 (N_4342,N_4254,N_4277);
or U4343 (N_4343,N_4232,N_4253);
nor U4344 (N_4344,N_4225,N_4215);
nor U4345 (N_4345,N_4269,N_4258);
nor U4346 (N_4346,N_4268,N_4257);
nand U4347 (N_4347,N_4216,N_4252);
nand U4348 (N_4348,N_4205,N_4298);
nand U4349 (N_4349,N_4255,N_4230);
nand U4350 (N_4350,N_4286,N_4280);
nor U4351 (N_4351,N_4253,N_4246);
and U4352 (N_4352,N_4274,N_4202);
nand U4353 (N_4353,N_4216,N_4283);
nand U4354 (N_4354,N_4250,N_4289);
nand U4355 (N_4355,N_4296,N_4289);
and U4356 (N_4356,N_4262,N_4290);
nand U4357 (N_4357,N_4203,N_4229);
or U4358 (N_4358,N_4254,N_4260);
and U4359 (N_4359,N_4207,N_4263);
nor U4360 (N_4360,N_4202,N_4230);
or U4361 (N_4361,N_4246,N_4214);
and U4362 (N_4362,N_4226,N_4214);
and U4363 (N_4363,N_4272,N_4240);
nand U4364 (N_4364,N_4286,N_4201);
nand U4365 (N_4365,N_4232,N_4285);
nand U4366 (N_4366,N_4200,N_4226);
and U4367 (N_4367,N_4256,N_4279);
nand U4368 (N_4368,N_4279,N_4271);
and U4369 (N_4369,N_4246,N_4262);
xor U4370 (N_4370,N_4264,N_4248);
and U4371 (N_4371,N_4293,N_4294);
nand U4372 (N_4372,N_4216,N_4241);
nor U4373 (N_4373,N_4289,N_4265);
xnor U4374 (N_4374,N_4296,N_4273);
nor U4375 (N_4375,N_4255,N_4275);
and U4376 (N_4376,N_4217,N_4281);
or U4377 (N_4377,N_4285,N_4257);
nand U4378 (N_4378,N_4296,N_4206);
nand U4379 (N_4379,N_4226,N_4259);
or U4380 (N_4380,N_4208,N_4281);
xor U4381 (N_4381,N_4249,N_4205);
and U4382 (N_4382,N_4201,N_4225);
and U4383 (N_4383,N_4249,N_4220);
and U4384 (N_4384,N_4201,N_4267);
and U4385 (N_4385,N_4229,N_4288);
or U4386 (N_4386,N_4201,N_4207);
nand U4387 (N_4387,N_4262,N_4259);
or U4388 (N_4388,N_4211,N_4284);
and U4389 (N_4389,N_4243,N_4234);
and U4390 (N_4390,N_4260,N_4208);
and U4391 (N_4391,N_4208,N_4225);
or U4392 (N_4392,N_4291,N_4299);
nor U4393 (N_4393,N_4241,N_4234);
nor U4394 (N_4394,N_4280,N_4249);
nand U4395 (N_4395,N_4242,N_4209);
nand U4396 (N_4396,N_4253,N_4224);
xor U4397 (N_4397,N_4263,N_4224);
and U4398 (N_4398,N_4271,N_4200);
and U4399 (N_4399,N_4245,N_4200);
nor U4400 (N_4400,N_4307,N_4381);
and U4401 (N_4401,N_4352,N_4384);
nor U4402 (N_4402,N_4301,N_4375);
and U4403 (N_4403,N_4365,N_4318);
nor U4404 (N_4404,N_4396,N_4321);
nor U4405 (N_4405,N_4336,N_4303);
and U4406 (N_4406,N_4387,N_4322);
xnor U4407 (N_4407,N_4376,N_4379);
and U4408 (N_4408,N_4347,N_4357);
or U4409 (N_4409,N_4385,N_4345);
and U4410 (N_4410,N_4350,N_4325);
nor U4411 (N_4411,N_4320,N_4348);
or U4412 (N_4412,N_4340,N_4392);
nor U4413 (N_4413,N_4333,N_4383);
and U4414 (N_4414,N_4369,N_4351);
nand U4415 (N_4415,N_4316,N_4304);
and U4416 (N_4416,N_4367,N_4344);
or U4417 (N_4417,N_4308,N_4310);
or U4418 (N_4418,N_4326,N_4373);
and U4419 (N_4419,N_4389,N_4338);
or U4420 (N_4420,N_4328,N_4354);
nor U4421 (N_4421,N_4315,N_4323);
or U4422 (N_4422,N_4331,N_4368);
xor U4423 (N_4423,N_4332,N_4370);
xor U4424 (N_4424,N_4341,N_4349);
and U4425 (N_4425,N_4339,N_4362);
or U4426 (N_4426,N_4342,N_4363);
nor U4427 (N_4427,N_4371,N_4399);
nor U4428 (N_4428,N_4395,N_4397);
xor U4429 (N_4429,N_4393,N_4334);
xor U4430 (N_4430,N_4305,N_4317);
nand U4431 (N_4431,N_4327,N_4335);
nand U4432 (N_4432,N_4309,N_4378);
nand U4433 (N_4433,N_4374,N_4302);
and U4434 (N_4434,N_4300,N_4382);
or U4435 (N_4435,N_4319,N_4390);
xor U4436 (N_4436,N_4306,N_4386);
or U4437 (N_4437,N_4329,N_4356);
nor U4438 (N_4438,N_4355,N_4311);
or U4439 (N_4439,N_4314,N_4388);
xor U4440 (N_4440,N_4359,N_4391);
nor U4441 (N_4441,N_4394,N_4377);
nand U4442 (N_4442,N_4346,N_4330);
nor U4443 (N_4443,N_4372,N_4358);
or U4444 (N_4444,N_4398,N_4380);
nor U4445 (N_4445,N_4313,N_4364);
xor U4446 (N_4446,N_4360,N_4343);
xor U4447 (N_4447,N_4353,N_4337);
and U4448 (N_4448,N_4361,N_4366);
nor U4449 (N_4449,N_4324,N_4312);
xor U4450 (N_4450,N_4325,N_4391);
and U4451 (N_4451,N_4336,N_4347);
or U4452 (N_4452,N_4300,N_4351);
and U4453 (N_4453,N_4366,N_4387);
or U4454 (N_4454,N_4370,N_4337);
and U4455 (N_4455,N_4367,N_4390);
nor U4456 (N_4456,N_4382,N_4350);
or U4457 (N_4457,N_4311,N_4304);
and U4458 (N_4458,N_4356,N_4314);
and U4459 (N_4459,N_4324,N_4333);
xor U4460 (N_4460,N_4369,N_4307);
nand U4461 (N_4461,N_4374,N_4323);
or U4462 (N_4462,N_4376,N_4307);
nand U4463 (N_4463,N_4377,N_4308);
nand U4464 (N_4464,N_4351,N_4340);
or U4465 (N_4465,N_4357,N_4325);
and U4466 (N_4466,N_4389,N_4336);
and U4467 (N_4467,N_4397,N_4349);
nand U4468 (N_4468,N_4322,N_4394);
and U4469 (N_4469,N_4315,N_4327);
nand U4470 (N_4470,N_4397,N_4380);
xnor U4471 (N_4471,N_4335,N_4383);
or U4472 (N_4472,N_4352,N_4327);
nand U4473 (N_4473,N_4370,N_4316);
xnor U4474 (N_4474,N_4387,N_4368);
nand U4475 (N_4475,N_4369,N_4352);
or U4476 (N_4476,N_4319,N_4323);
nor U4477 (N_4477,N_4308,N_4319);
nor U4478 (N_4478,N_4334,N_4351);
nand U4479 (N_4479,N_4331,N_4303);
nand U4480 (N_4480,N_4301,N_4377);
nor U4481 (N_4481,N_4381,N_4303);
xnor U4482 (N_4482,N_4342,N_4348);
nor U4483 (N_4483,N_4397,N_4338);
and U4484 (N_4484,N_4353,N_4329);
or U4485 (N_4485,N_4330,N_4377);
and U4486 (N_4486,N_4377,N_4390);
nand U4487 (N_4487,N_4379,N_4322);
xnor U4488 (N_4488,N_4385,N_4369);
or U4489 (N_4489,N_4347,N_4321);
and U4490 (N_4490,N_4377,N_4337);
nand U4491 (N_4491,N_4329,N_4380);
nor U4492 (N_4492,N_4359,N_4357);
nor U4493 (N_4493,N_4391,N_4356);
nand U4494 (N_4494,N_4337,N_4323);
nand U4495 (N_4495,N_4384,N_4305);
nand U4496 (N_4496,N_4310,N_4330);
nor U4497 (N_4497,N_4389,N_4323);
xor U4498 (N_4498,N_4375,N_4392);
nand U4499 (N_4499,N_4313,N_4355);
xnor U4500 (N_4500,N_4455,N_4418);
or U4501 (N_4501,N_4431,N_4489);
nor U4502 (N_4502,N_4433,N_4417);
or U4503 (N_4503,N_4481,N_4478);
nand U4504 (N_4504,N_4479,N_4416);
and U4505 (N_4505,N_4421,N_4487);
and U4506 (N_4506,N_4465,N_4493);
nand U4507 (N_4507,N_4406,N_4486);
and U4508 (N_4508,N_4452,N_4471);
or U4509 (N_4509,N_4469,N_4461);
and U4510 (N_4510,N_4442,N_4467);
and U4511 (N_4511,N_4496,N_4420);
nand U4512 (N_4512,N_4498,N_4474);
xor U4513 (N_4513,N_4429,N_4483);
and U4514 (N_4514,N_4482,N_4468);
nor U4515 (N_4515,N_4404,N_4475);
nand U4516 (N_4516,N_4435,N_4466);
nand U4517 (N_4517,N_4462,N_4427);
and U4518 (N_4518,N_4400,N_4432);
nor U4519 (N_4519,N_4444,N_4436);
nor U4520 (N_4520,N_4495,N_4440);
nor U4521 (N_4521,N_4454,N_4439);
nand U4522 (N_4522,N_4409,N_4443);
nand U4523 (N_4523,N_4476,N_4470);
nand U4524 (N_4524,N_4428,N_4456);
nor U4525 (N_4525,N_4480,N_4463);
xor U4526 (N_4526,N_4494,N_4407);
and U4527 (N_4527,N_4419,N_4472);
nand U4528 (N_4528,N_4445,N_4424);
nor U4529 (N_4529,N_4459,N_4437);
or U4530 (N_4530,N_4405,N_4492);
xor U4531 (N_4531,N_4447,N_4422);
nor U4532 (N_4532,N_4453,N_4488);
and U4533 (N_4533,N_4425,N_4460);
or U4534 (N_4534,N_4402,N_4412);
nand U4535 (N_4535,N_4423,N_4490);
nand U4536 (N_4536,N_4401,N_4410);
nand U4537 (N_4537,N_4411,N_4438);
nand U4538 (N_4538,N_4414,N_4497);
nand U4539 (N_4539,N_4485,N_4451);
and U4540 (N_4540,N_4426,N_4464);
nand U4541 (N_4541,N_4408,N_4477);
nand U4542 (N_4542,N_4499,N_4458);
nor U4543 (N_4543,N_4430,N_4415);
or U4544 (N_4544,N_4484,N_4413);
or U4545 (N_4545,N_4448,N_4450);
nor U4546 (N_4546,N_4457,N_4473);
nand U4547 (N_4547,N_4434,N_4449);
or U4548 (N_4548,N_4491,N_4403);
and U4549 (N_4549,N_4441,N_4446);
nand U4550 (N_4550,N_4442,N_4498);
nor U4551 (N_4551,N_4419,N_4482);
nand U4552 (N_4552,N_4428,N_4409);
and U4553 (N_4553,N_4472,N_4414);
nand U4554 (N_4554,N_4474,N_4447);
or U4555 (N_4555,N_4487,N_4430);
xor U4556 (N_4556,N_4406,N_4430);
nor U4557 (N_4557,N_4470,N_4409);
or U4558 (N_4558,N_4465,N_4415);
nand U4559 (N_4559,N_4483,N_4490);
and U4560 (N_4560,N_4480,N_4420);
xor U4561 (N_4561,N_4407,N_4449);
nor U4562 (N_4562,N_4410,N_4462);
nand U4563 (N_4563,N_4483,N_4423);
nor U4564 (N_4564,N_4472,N_4420);
and U4565 (N_4565,N_4450,N_4441);
and U4566 (N_4566,N_4432,N_4461);
nor U4567 (N_4567,N_4418,N_4440);
or U4568 (N_4568,N_4472,N_4490);
nor U4569 (N_4569,N_4492,N_4425);
nor U4570 (N_4570,N_4461,N_4456);
and U4571 (N_4571,N_4426,N_4438);
xor U4572 (N_4572,N_4415,N_4406);
and U4573 (N_4573,N_4450,N_4493);
and U4574 (N_4574,N_4425,N_4475);
and U4575 (N_4575,N_4412,N_4471);
or U4576 (N_4576,N_4417,N_4412);
and U4577 (N_4577,N_4494,N_4433);
nor U4578 (N_4578,N_4402,N_4448);
and U4579 (N_4579,N_4463,N_4440);
or U4580 (N_4580,N_4496,N_4450);
and U4581 (N_4581,N_4485,N_4438);
and U4582 (N_4582,N_4459,N_4486);
nor U4583 (N_4583,N_4479,N_4467);
and U4584 (N_4584,N_4454,N_4428);
xnor U4585 (N_4585,N_4419,N_4415);
nor U4586 (N_4586,N_4440,N_4434);
and U4587 (N_4587,N_4457,N_4455);
nor U4588 (N_4588,N_4431,N_4443);
and U4589 (N_4589,N_4461,N_4489);
and U4590 (N_4590,N_4438,N_4403);
or U4591 (N_4591,N_4406,N_4492);
and U4592 (N_4592,N_4434,N_4439);
nor U4593 (N_4593,N_4483,N_4458);
nand U4594 (N_4594,N_4474,N_4413);
nor U4595 (N_4595,N_4461,N_4483);
and U4596 (N_4596,N_4448,N_4445);
nor U4597 (N_4597,N_4454,N_4496);
xor U4598 (N_4598,N_4448,N_4440);
and U4599 (N_4599,N_4493,N_4454);
nand U4600 (N_4600,N_4505,N_4514);
nand U4601 (N_4601,N_4571,N_4578);
nand U4602 (N_4602,N_4573,N_4534);
nor U4603 (N_4603,N_4548,N_4563);
nand U4604 (N_4604,N_4598,N_4524);
nor U4605 (N_4605,N_4575,N_4512);
nor U4606 (N_4606,N_4545,N_4549);
or U4607 (N_4607,N_4579,N_4509);
nor U4608 (N_4608,N_4569,N_4517);
nor U4609 (N_4609,N_4551,N_4580);
and U4610 (N_4610,N_4538,N_4594);
xnor U4611 (N_4611,N_4555,N_4504);
nor U4612 (N_4612,N_4539,N_4570);
nand U4613 (N_4613,N_4596,N_4576);
nor U4614 (N_4614,N_4567,N_4523);
and U4615 (N_4615,N_4595,N_4581);
nand U4616 (N_4616,N_4584,N_4521);
nor U4617 (N_4617,N_4529,N_4593);
nand U4618 (N_4618,N_4564,N_4518);
nor U4619 (N_4619,N_4519,N_4585);
and U4620 (N_4620,N_4520,N_4516);
nor U4621 (N_4621,N_4515,N_4531);
or U4622 (N_4622,N_4507,N_4550);
or U4623 (N_4623,N_4542,N_4508);
nand U4624 (N_4624,N_4566,N_4546);
nand U4625 (N_4625,N_4556,N_4528);
nand U4626 (N_4626,N_4536,N_4583);
or U4627 (N_4627,N_4582,N_4527);
nand U4628 (N_4628,N_4553,N_4503);
nand U4629 (N_4629,N_4590,N_4561);
xor U4630 (N_4630,N_4513,N_4589);
or U4631 (N_4631,N_4547,N_4537);
or U4632 (N_4632,N_4543,N_4502);
nand U4633 (N_4633,N_4558,N_4560);
nand U4634 (N_4634,N_4535,N_4500);
nor U4635 (N_4635,N_4510,N_4540);
and U4636 (N_4636,N_4591,N_4559);
nand U4637 (N_4637,N_4532,N_4599);
or U4638 (N_4638,N_4588,N_4574);
nor U4639 (N_4639,N_4541,N_4587);
xor U4640 (N_4640,N_4530,N_4557);
or U4641 (N_4641,N_4565,N_4525);
and U4642 (N_4642,N_4552,N_4506);
and U4643 (N_4643,N_4554,N_4577);
or U4644 (N_4644,N_4572,N_4568);
nand U4645 (N_4645,N_4511,N_4562);
nand U4646 (N_4646,N_4501,N_4544);
or U4647 (N_4647,N_4533,N_4522);
and U4648 (N_4648,N_4586,N_4597);
xor U4649 (N_4649,N_4526,N_4592);
nand U4650 (N_4650,N_4518,N_4587);
xnor U4651 (N_4651,N_4530,N_4548);
nand U4652 (N_4652,N_4503,N_4551);
nor U4653 (N_4653,N_4581,N_4534);
nand U4654 (N_4654,N_4565,N_4521);
nand U4655 (N_4655,N_4546,N_4589);
or U4656 (N_4656,N_4530,N_4585);
nor U4657 (N_4657,N_4586,N_4519);
nand U4658 (N_4658,N_4503,N_4561);
nor U4659 (N_4659,N_4585,N_4538);
nand U4660 (N_4660,N_4538,N_4542);
and U4661 (N_4661,N_4584,N_4585);
and U4662 (N_4662,N_4538,N_4565);
nor U4663 (N_4663,N_4548,N_4503);
xor U4664 (N_4664,N_4520,N_4551);
and U4665 (N_4665,N_4577,N_4502);
or U4666 (N_4666,N_4557,N_4518);
nor U4667 (N_4667,N_4576,N_4511);
and U4668 (N_4668,N_4579,N_4522);
nor U4669 (N_4669,N_4586,N_4525);
or U4670 (N_4670,N_4553,N_4596);
xnor U4671 (N_4671,N_4508,N_4526);
nand U4672 (N_4672,N_4530,N_4599);
and U4673 (N_4673,N_4533,N_4520);
nor U4674 (N_4674,N_4588,N_4522);
and U4675 (N_4675,N_4540,N_4511);
nor U4676 (N_4676,N_4513,N_4564);
and U4677 (N_4677,N_4565,N_4540);
or U4678 (N_4678,N_4598,N_4526);
and U4679 (N_4679,N_4523,N_4580);
or U4680 (N_4680,N_4538,N_4597);
nor U4681 (N_4681,N_4595,N_4574);
nor U4682 (N_4682,N_4537,N_4523);
and U4683 (N_4683,N_4592,N_4547);
or U4684 (N_4684,N_4526,N_4563);
and U4685 (N_4685,N_4582,N_4523);
xnor U4686 (N_4686,N_4547,N_4584);
or U4687 (N_4687,N_4564,N_4583);
nand U4688 (N_4688,N_4501,N_4586);
nand U4689 (N_4689,N_4505,N_4580);
or U4690 (N_4690,N_4536,N_4501);
or U4691 (N_4691,N_4595,N_4539);
nand U4692 (N_4692,N_4502,N_4575);
xor U4693 (N_4693,N_4528,N_4584);
xor U4694 (N_4694,N_4507,N_4538);
nor U4695 (N_4695,N_4574,N_4583);
nand U4696 (N_4696,N_4586,N_4555);
nor U4697 (N_4697,N_4514,N_4504);
nand U4698 (N_4698,N_4554,N_4532);
nand U4699 (N_4699,N_4527,N_4504);
or U4700 (N_4700,N_4676,N_4647);
nand U4701 (N_4701,N_4654,N_4608);
or U4702 (N_4702,N_4661,N_4697);
and U4703 (N_4703,N_4609,N_4681);
xor U4704 (N_4704,N_4600,N_4639);
nor U4705 (N_4705,N_4698,N_4638);
nor U4706 (N_4706,N_4607,N_4664);
or U4707 (N_4707,N_4651,N_4688);
nor U4708 (N_4708,N_4689,N_4628);
nand U4709 (N_4709,N_4640,N_4643);
or U4710 (N_4710,N_4632,N_4690);
nand U4711 (N_4711,N_4668,N_4614);
or U4712 (N_4712,N_4653,N_4613);
nand U4713 (N_4713,N_4626,N_4660);
or U4714 (N_4714,N_4627,N_4618);
or U4715 (N_4715,N_4629,N_4602);
or U4716 (N_4716,N_4683,N_4657);
or U4717 (N_4717,N_4642,N_4658);
nor U4718 (N_4718,N_4666,N_4695);
or U4719 (N_4719,N_4636,N_4691);
and U4720 (N_4720,N_4696,N_4617);
and U4721 (N_4721,N_4693,N_4685);
nor U4722 (N_4722,N_4645,N_4623);
and U4723 (N_4723,N_4699,N_4601);
and U4724 (N_4724,N_4652,N_4615);
xnor U4725 (N_4725,N_4631,N_4678);
nand U4726 (N_4726,N_4692,N_4605);
nand U4727 (N_4727,N_4619,N_4659);
nand U4728 (N_4728,N_4646,N_4633);
or U4729 (N_4729,N_4663,N_4606);
nand U4730 (N_4730,N_4649,N_4644);
nor U4731 (N_4731,N_4684,N_4622);
nand U4732 (N_4732,N_4662,N_4612);
or U4733 (N_4733,N_4641,N_4637);
xnor U4734 (N_4734,N_4635,N_4621);
or U4735 (N_4735,N_4620,N_4669);
nand U4736 (N_4736,N_4687,N_4648);
and U4737 (N_4737,N_4650,N_4665);
nor U4738 (N_4738,N_4634,N_4694);
nand U4739 (N_4739,N_4667,N_4671);
nor U4740 (N_4740,N_4686,N_4625);
nand U4741 (N_4741,N_4656,N_4655);
xnor U4742 (N_4742,N_4672,N_4616);
nand U4743 (N_4743,N_4604,N_4630);
nand U4744 (N_4744,N_4675,N_4682);
and U4745 (N_4745,N_4610,N_4679);
xnor U4746 (N_4746,N_4674,N_4603);
xor U4747 (N_4747,N_4677,N_4680);
nand U4748 (N_4748,N_4624,N_4670);
xor U4749 (N_4749,N_4673,N_4611);
xor U4750 (N_4750,N_4632,N_4682);
and U4751 (N_4751,N_4667,N_4676);
xnor U4752 (N_4752,N_4693,N_4676);
or U4753 (N_4753,N_4647,N_4635);
nand U4754 (N_4754,N_4686,N_4698);
and U4755 (N_4755,N_4679,N_4699);
nor U4756 (N_4756,N_4678,N_4684);
nor U4757 (N_4757,N_4676,N_4672);
nor U4758 (N_4758,N_4621,N_4646);
or U4759 (N_4759,N_4617,N_4669);
nand U4760 (N_4760,N_4698,N_4609);
nor U4761 (N_4761,N_4628,N_4618);
and U4762 (N_4762,N_4681,N_4626);
xor U4763 (N_4763,N_4632,N_4644);
nor U4764 (N_4764,N_4609,N_4672);
and U4765 (N_4765,N_4623,N_4606);
or U4766 (N_4766,N_4661,N_4683);
or U4767 (N_4767,N_4682,N_4693);
nand U4768 (N_4768,N_4669,N_4642);
nor U4769 (N_4769,N_4687,N_4684);
or U4770 (N_4770,N_4648,N_4660);
nand U4771 (N_4771,N_4667,N_4648);
nand U4772 (N_4772,N_4621,N_4676);
nor U4773 (N_4773,N_4646,N_4658);
and U4774 (N_4774,N_4655,N_4668);
xor U4775 (N_4775,N_4672,N_4606);
nand U4776 (N_4776,N_4626,N_4661);
or U4777 (N_4777,N_4635,N_4633);
or U4778 (N_4778,N_4669,N_4686);
and U4779 (N_4779,N_4674,N_4627);
nor U4780 (N_4780,N_4636,N_4689);
nand U4781 (N_4781,N_4627,N_4614);
nand U4782 (N_4782,N_4663,N_4640);
and U4783 (N_4783,N_4671,N_4683);
and U4784 (N_4784,N_4672,N_4607);
nor U4785 (N_4785,N_4603,N_4606);
nor U4786 (N_4786,N_4624,N_4699);
or U4787 (N_4787,N_4676,N_4687);
and U4788 (N_4788,N_4634,N_4606);
or U4789 (N_4789,N_4672,N_4602);
nor U4790 (N_4790,N_4619,N_4692);
and U4791 (N_4791,N_4620,N_4665);
nor U4792 (N_4792,N_4669,N_4687);
nand U4793 (N_4793,N_4671,N_4675);
or U4794 (N_4794,N_4673,N_4656);
nand U4795 (N_4795,N_4687,N_4606);
nand U4796 (N_4796,N_4631,N_4661);
and U4797 (N_4797,N_4662,N_4614);
nor U4798 (N_4798,N_4661,N_4673);
nand U4799 (N_4799,N_4671,N_4635);
or U4800 (N_4800,N_4799,N_4736);
nor U4801 (N_4801,N_4730,N_4741);
or U4802 (N_4802,N_4781,N_4709);
or U4803 (N_4803,N_4748,N_4740);
nand U4804 (N_4804,N_4758,N_4732);
or U4805 (N_4805,N_4771,N_4765);
nor U4806 (N_4806,N_4782,N_4718);
and U4807 (N_4807,N_4723,N_4789);
and U4808 (N_4808,N_4791,N_4752);
or U4809 (N_4809,N_4735,N_4762);
nand U4810 (N_4810,N_4753,N_4727);
and U4811 (N_4811,N_4760,N_4792);
or U4812 (N_4812,N_4761,N_4734);
xnor U4813 (N_4813,N_4744,N_4783);
nand U4814 (N_4814,N_4745,N_4726);
and U4815 (N_4815,N_4721,N_4788);
and U4816 (N_4816,N_4764,N_4767);
or U4817 (N_4817,N_4712,N_4777);
and U4818 (N_4818,N_4702,N_4706);
nand U4819 (N_4819,N_4776,N_4763);
nand U4820 (N_4820,N_4707,N_4793);
xnor U4821 (N_4821,N_4739,N_4780);
nand U4822 (N_4822,N_4756,N_4749);
and U4823 (N_4823,N_4785,N_4773);
nand U4824 (N_4824,N_4779,N_4701);
nand U4825 (N_4825,N_4746,N_4733);
and U4826 (N_4826,N_4742,N_4757);
and U4827 (N_4827,N_4769,N_4750);
nor U4828 (N_4828,N_4724,N_4704);
xor U4829 (N_4829,N_4705,N_4775);
or U4830 (N_4830,N_4798,N_4738);
or U4831 (N_4831,N_4755,N_4796);
or U4832 (N_4832,N_4794,N_4784);
nand U4833 (N_4833,N_4731,N_4703);
nor U4834 (N_4834,N_4720,N_4747);
or U4835 (N_4835,N_4722,N_4719);
or U4836 (N_4836,N_4795,N_4708);
nor U4837 (N_4837,N_4797,N_4711);
xor U4838 (N_4838,N_4759,N_4714);
nand U4839 (N_4839,N_4710,N_4790);
nand U4840 (N_4840,N_4766,N_4754);
nor U4841 (N_4841,N_4770,N_4743);
nand U4842 (N_4842,N_4717,N_4787);
or U4843 (N_4843,N_4768,N_4728);
and U4844 (N_4844,N_4737,N_4774);
nand U4845 (N_4845,N_4729,N_4778);
nor U4846 (N_4846,N_4725,N_4751);
nor U4847 (N_4847,N_4700,N_4772);
and U4848 (N_4848,N_4715,N_4716);
nor U4849 (N_4849,N_4713,N_4786);
or U4850 (N_4850,N_4715,N_4788);
xnor U4851 (N_4851,N_4795,N_4710);
nor U4852 (N_4852,N_4709,N_4732);
nor U4853 (N_4853,N_4749,N_4784);
nor U4854 (N_4854,N_4750,N_4784);
and U4855 (N_4855,N_4798,N_4792);
xnor U4856 (N_4856,N_4750,N_4782);
nand U4857 (N_4857,N_4777,N_4771);
xnor U4858 (N_4858,N_4759,N_4710);
nor U4859 (N_4859,N_4704,N_4740);
nand U4860 (N_4860,N_4751,N_4785);
and U4861 (N_4861,N_4725,N_4745);
and U4862 (N_4862,N_4703,N_4754);
and U4863 (N_4863,N_4781,N_4721);
nor U4864 (N_4864,N_4736,N_4796);
and U4865 (N_4865,N_4727,N_4751);
and U4866 (N_4866,N_4765,N_4733);
or U4867 (N_4867,N_4750,N_4788);
or U4868 (N_4868,N_4711,N_4737);
and U4869 (N_4869,N_4755,N_4769);
nand U4870 (N_4870,N_4759,N_4708);
nand U4871 (N_4871,N_4765,N_4792);
nor U4872 (N_4872,N_4785,N_4722);
nor U4873 (N_4873,N_4733,N_4776);
nand U4874 (N_4874,N_4760,N_4787);
nand U4875 (N_4875,N_4789,N_4702);
nand U4876 (N_4876,N_4743,N_4710);
and U4877 (N_4877,N_4742,N_4728);
or U4878 (N_4878,N_4776,N_4781);
and U4879 (N_4879,N_4741,N_4705);
nand U4880 (N_4880,N_4787,N_4763);
or U4881 (N_4881,N_4731,N_4755);
or U4882 (N_4882,N_4744,N_4773);
or U4883 (N_4883,N_4756,N_4718);
nor U4884 (N_4884,N_4752,N_4754);
nor U4885 (N_4885,N_4761,N_4744);
or U4886 (N_4886,N_4744,N_4780);
or U4887 (N_4887,N_4756,N_4710);
and U4888 (N_4888,N_4746,N_4710);
or U4889 (N_4889,N_4728,N_4705);
nor U4890 (N_4890,N_4723,N_4790);
nor U4891 (N_4891,N_4726,N_4780);
or U4892 (N_4892,N_4750,N_4753);
and U4893 (N_4893,N_4729,N_4779);
nor U4894 (N_4894,N_4775,N_4759);
nand U4895 (N_4895,N_4702,N_4766);
and U4896 (N_4896,N_4771,N_4793);
nand U4897 (N_4897,N_4791,N_4744);
or U4898 (N_4898,N_4774,N_4773);
nand U4899 (N_4899,N_4752,N_4771);
or U4900 (N_4900,N_4845,N_4856);
or U4901 (N_4901,N_4825,N_4861);
nor U4902 (N_4902,N_4854,N_4817);
nand U4903 (N_4903,N_4853,N_4842);
nor U4904 (N_4904,N_4829,N_4808);
nor U4905 (N_4905,N_4877,N_4879);
or U4906 (N_4906,N_4850,N_4863);
nor U4907 (N_4907,N_4883,N_4858);
and U4908 (N_4908,N_4897,N_4843);
or U4909 (N_4909,N_4881,N_4831);
or U4910 (N_4910,N_4888,N_4822);
xnor U4911 (N_4911,N_4847,N_4837);
nor U4912 (N_4912,N_4840,N_4846);
nor U4913 (N_4913,N_4813,N_4809);
nand U4914 (N_4914,N_4836,N_4864);
nand U4915 (N_4915,N_4814,N_4884);
nand U4916 (N_4916,N_4844,N_4875);
and U4917 (N_4917,N_4886,N_4895);
nor U4918 (N_4918,N_4832,N_4835);
nand U4919 (N_4919,N_4824,N_4859);
xor U4920 (N_4920,N_4880,N_4876);
nand U4921 (N_4921,N_4872,N_4834);
nor U4922 (N_4922,N_4860,N_4801);
xor U4923 (N_4923,N_4870,N_4849);
or U4924 (N_4924,N_4894,N_4818);
nand U4925 (N_4925,N_4841,N_4819);
and U4926 (N_4926,N_4828,N_4807);
nand U4927 (N_4927,N_4890,N_4857);
nor U4928 (N_4928,N_4804,N_4803);
or U4929 (N_4929,N_4805,N_4852);
and U4930 (N_4930,N_4891,N_4893);
or U4931 (N_4931,N_4867,N_4810);
xor U4932 (N_4932,N_4869,N_4878);
or U4933 (N_4933,N_4800,N_4868);
nand U4934 (N_4934,N_4865,N_4815);
nand U4935 (N_4935,N_4823,N_4855);
and U4936 (N_4936,N_4887,N_4838);
nor U4937 (N_4937,N_4820,N_4892);
xnor U4938 (N_4938,N_4816,N_4811);
and U4939 (N_4939,N_4848,N_4871);
or U4940 (N_4940,N_4874,N_4898);
nand U4941 (N_4941,N_4821,N_4833);
or U4942 (N_4942,N_4839,N_4899);
nor U4943 (N_4943,N_4826,N_4806);
nand U4944 (N_4944,N_4885,N_4830);
and U4945 (N_4945,N_4873,N_4812);
and U4946 (N_4946,N_4862,N_4896);
or U4947 (N_4947,N_4827,N_4851);
or U4948 (N_4948,N_4882,N_4802);
and U4949 (N_4949,N_4889,N_4866);
or U4950 (N_4950,N_4882,N_4883);
or U4951 (N_4951,N_4849,N_4899);
or U4952 (N_4952,N_4831,N_4852);
or U4953 (N_4953,N_4815,N_4805);
and U4954 (N_4954,N_4833,N_4855);
and U4955 (N_4955,N_4859,N_4847);
or U4956 (N_4956,N_4841,N_4816);
and U4957 (N_4957,N_4804,N_4844);
nor U4958 (N_4958,N_4814,N_4832);
and U4959 (N_4959,N_4821,N_4823);
xor U4960 (N_4960,N_4811,N_4807);
nor U4961 (N_4961,N_4872,N_4862);
nor U4962 (N_4962,N_4842,N_4846);
nor U4963 (N_4963,N_4880,N_4871);
nand U4964 (N_4964,N_4890,N_4847);
xor U4965 (N_4965,N_4890,N_4867);
or U4966 (N_4966,N_4814,N_4823);
or U4967 (N_4967,N_4848,N_4868);
or U4968 (N_4968,N_4812,N_4882);
nor U4969 (N_4969,N_4803,N_4835);
nor U4970 (N_4970,N_4812,N_4897);
and U4971 (N_4971,N_4872,N_4857);
nand U4972 (N_4972,N_4837,N_4845);
and U4973 (N_4973,N_4853,N_4823);
or U4974 (N_4974,N_4824,N_4812);
nor U4975 (N_4975,N_4854,N_4860);
nand U4976 (N_4976,N_4812,N_4886);
and U4977 (N_4977,N_4878,N_4870);
and U4978 (N_4978,N_4897,N_4888);
nor U4979 (N_4979,N_4896,N_4858);
nand U4980 (N_4980,N_4898,N_4806);
or U4981 (N_4981,N_4846,N_4893);
nor U4982 (N_4982,N_4858,N_4832);
nor U4983 (N_4983,N_4895,N_4884);
or U4984 (N_4984,N_4805,N_4894);
nand U4985 (N_4985,N_4873,N_4830);
nand U4986 (N_4986,N_4808,N_4813);
nor U4987 (N_4987,N_4893,N_4802);
or U4988 (N_4988,N_4866,N_4860);
nor U4989 (N_4989,N_4812,N_4828);
or U4990 (N_4990,N_4805,N_4825);
nand U4991 (N_4991,N_4824,N_4845);
nand U4992 (N_4992,N_4852,N_4882);
xnor U4993 (N_4993,N_4840,N_4895);
and U4994 (N_4994,N_4861,N_4883);
and U4995 (N_4995,N_4870,N_4895);
nor U4996 (N_4996,N_4850,N_4893);
xor U4997 (N_4997,N_4817,N_4849);
nand U4998 (N_4998,N_4856,N_4867);
and U4999 (N_4999,N_4804,N_4807);
nand U5000 (N_5000,N_4928,N_4966);
or U5001 (N_5001,N_4985,N_4961);
xnor U5002 (N_5002,N_4965,N_4973);
and U5003 (N_5003,N_4907,N_4934);
nand U5004 (N_5004,N_4901,N_4984);
or U5005 (N_5005,N_4914,N_4975);
xor U5006 (N_5006,N_4991,N_4938);
or U5007 (N_5007,N_4983,N_4996);
or U5008 (N_5008,N_4923,N_4962);
and U5009 (N_5009,N_4908,N_4954);
nor U5010 (N_5010,N_4902,N_4955);
and U5011 (N_5011,N_4950,N_4968);
or U5012 (N_5012,N_4913,N_4929);
nand U5013 (N_5013,N_4967,N_4932);
nand U5014 (N_5014,N_4953,N_4919);
or U5015 (N_5015,N_4921,N_4992);
nor U5016 (N_5016,N_4974,N_4942);
or U5017 (N_5017,N_4920,N_4916);
xor U5018 (N_5018,N_4910,N_4944);
and U5019 (N_5019,N_4939,N_4937);
or U5020 (N_5020,N_4918,N_4960);
or U5021 (N_5021,N_4997,N_4911);
nor U5022 (N_5022,N_4957,N_4917);
nand U5023 (N_5023,N_4906,N_4982);
or U5024 (N_5024,N_4976,N_4930);
xnor U5025 (N_5025,N_4980,N_4989);
nand U5026 (N_5026,N_4999,N_4926);
xnor U5027 (N_5027,N_4998,N_4900);
and U5028 (N_5028,N_4943,N_4963);
and U5029 (N_5029,N_4958,N_4922);
and U5030 (N_5030,N_4935,N_4993);
xnor U5031 (N_5031,N_4940,N_4990);
xor U5032 (N_5032,N_4915,N_4948);
or U5033 (N_5033,N_4972,N_4970);
and U5034 (N_5034,N_4969,N_4925);
and U5035 (N_5035,N_4956,N_4947);
nor U5036 (N_5036,N_4994,N_4981);
xnor U5037 (N_5037,N_4959,N_4995);
and U5038 (N_5038,N_4931,N_4912);
and U5039 (N_5039,N_4909,N_4905);
nand U5040 (N_5040,N_4946,N_4951);
or U5041 (N_5041,N_4986,N_4936);
nand U5042 (N_5042,N_4927,N_4979);
or U5043 (N_5043,N_4941,N_4952);
xnor U5044 (N_5044,N_4903,N_4904);
and U5045 (N_5045,N_4949,N_4987);
and U5046 (N_5046,N_4964,N_4978);
or U5047 (N_5047,N_4945,N_4988);
nand U5048 (N_5048,N_4924,N_4933);
nor U5049 (N_5049,N_4977,N_4971);
nand U5050 (N_5050,N_4973,N_4919);
and U5051 (N_5051,N_4921,N_4999);
nor U5052 (N_5052,N_4941,N_4919);
nor U5053 (N_5053,N_4900,N_4988);
nand U5054 (N_5054,N_4978,N_4930);
or U5055 (N_5055,N_4934,N_4947);
nor U5056 (N_5056,N_4976,N_4989);
nor U5057 (N_5057,N_4986,N_4923);
nand U5058 (N_5058,N_4931,N_4989);
or U5059 (N_5059,N_4962,N_4902);
nor U5060 (N_5060,N_4993,N_4905);
or U5061 (N_5061,N_4965,N_4932);
nor U5062 (N_5062,N_4935,N_4948);
nor U5063 (N_5063,N_4934,N_4908);
or U5064 (N_5064,N_4929,N_4968);
and U5065 (N_5065,N_4979,N_4991);
nor U5066 (N_5066,N_4945,N_4937);
nor U5067 (N_5067,N_4983,N_4989);
nor U5068 (N_5068,N_4916,N_4959);
xor U5069 (N_5069,N_4933,N_4995);
nor U5070 (N_5070,N_4981,N_4928);
nor U5071 (N_5071,N_4934,N_4971);
and U5072 (N_5072,N_4957,N_4937);
nand U5073 (N_5073,N_4997,N_4906);
and U5074 (N_5074,N_4917,N_4928);
xnor U5075 (N_5075,N_4948,N_4964);
and U5076 (N_5076,N_4919,N_4990);
nor U5077 (N_5077,N_4919,N_4969);
nor U5078 (N_5078,N_4921,N_4956);
or U5079 (N_5079,N_4984,N_4922);
or U5080 (N_5080,N_4932,N_4959);
nand U5081 (N_5081,N_4953,N_4971);
or U5082 (N_5082,N_4956,N_4953);
nor U5083 (N_5083,N_4918,N_4958);
nor U5084 (N_5084,N_4931,N_4958);
and U5085 (N_5085,N_4974,N_4921);
nor U5086 (N_5086,N_4985,N_4973);
and U5087 (N_5087,N_4929,N_4902);
nand U5088 (N_5088,N_4914,N_4969);
xor U5089 (N_5089,N_4959,N_4953);
and U5090 (N_5090,N_4918,N_4920);
or U5091 (N_5091,N_4932,N_4968);
nand U5092 (N_5092,N_4916,N_4918);
or U5093 (N_5093,N_4931,N_4945);
or U5094 (N_5094,N_4998,N_4916);
or U5095 (N_5095,N_4930,N_4966);
nor U5096 (N_5096,N_4946,N_4950);
nor U5097 (N_5097,N_4925,N_4915);
or U5098 (N_5098,N_4979,N_4997);
nand U5099 (N_5099,N_4965,N_4915);
and U5100 (N_5100,N_5013,N_5029);
and U5101 (N_5101,N_5090,N_5088);
or U5102 (N_5102,N_5073,N_5066);
or U5103 (N_5103,N_5007,N_5052);
nand U5104 (N_5104,N_5093,N_5087);
and U5105 (N_5105,N_5060,N_5036);
or U5106 (N_5106,N_5047,N_5082);
xnor U5107 (N_5107,N_5034,N_5035);
nand U5108 (N_5108,N_5018,N_5065);
nand U5109 (N_5109,N_5039,N_5080);
nor U5110 (N_5110,N_5075,N_5097);
xnor U5111 (N_5111,N_5048,N_5068);
and U5112 (N_5112,N_5085,N_5062);
nor U5113 (N_5113,N_5050,N_5030);
nand U5114 (N_5114,N_5053,N_5067);
or U5115 (N_5115,N_5045,N_5072);
nor U5116 (N_5116,N_5070,N_5061);
or U5117 (N_5117,N_5023,N_5041);
and U5118 (N_5118,N_5042,N_5046);
xor U5119 (N_5119,N_5057,N_5074);
and U5120 (N_5120,N_5028,N_5038);
or U5121 (N_5121,N_5021,N_5032);
and U5122 (N_5122,N_5076,N_5006);
or U5123 (N_5123,N_5025,N_5010);
and U5124 (N_5124,N_5033,N_5044);
nand U5125 (N_5125,N_5043,N_5058);
nand U5126 (N_5126,N_5089,N_5055);
nor U5127 (N_5127,N_5022,N_5009);
and U5128 (N_5128,N_5083,N_5064);
nor U5129 (N_5129,N_5069,N_5000);
nand U5130 (N_5130,N_5096,N_5081);
nand U5131 (N_5131,N_5011,N_5098);
nand U5132 (N_5132,N_5063,N_5020);
and U5133 (N_5133,N_5084,N_5024);
nand U5134 (N_5134,N_5015,N_5078);
xnor U5135 (N_5135,N_5040,N_5086);
and U5136 (N_5136,N_5091,N_5017);
and U5137 (N_5137,N_5005,N_5008);
or U5138 (N_5138,N_5079,N_5016);
and U5139 (N_5139,N_5031,N_5014);
nor U5140 (N_5140,N_5003,N_5037);
nor U5141 (N_5141,N_5051,N_5077);
and U5142 (N_5142,N_5004,N_5099);
or U5143 (N_5143,N_5071,N_5092);
nor U5144 (N_5144,N_5002,N_5054);
xnor U5145 (N_5145,N_5049,N_5027);
nand U5146 (N_5146,N_5056,N_5059);
or U5147 (N_5147,N_5026,N_5012);
and U5148 (N_5148,N_5019,N_5095);
nand U5149 (N_5149,N_5001,N_5094);
and U5150 (N_5150,N_5011,N_5038);
nand U5151 (N_5151,N_5013,N_5082);
nor U5152 (N_5152,N_5063,N_5053);
or U5153 (N_5153,N_5045,N_5046);
and U5154 (N_5154,N_5012,N_5054);
and U5155 (N_5155,N_5065,N_5009);
nor U5156 (N_5156,N_5021,N_5074);
and U5157 (N_5157,N_5062,N_5064);
or U5158 (N_5158,N_5047,N_5033);
nor U5159 (N_5159,N_5031,N_5095);
and U5160 (N_5160,N_5081,N_5076);
xnor U5161 (N_5161,N_5063,N_5099);
and U5162 (N_5162,N_5072,N_5005);
xor U5163 (N_5163,N_5075,N_5025);
nand U5164 (N_5164,N_5096,N_5003);
and U5165 (N_5165,N_5009,N_5030);
or U5166 (N_5166,N_5004,N_5054);
or U5167 (N_5167,N_5043,N_5088);
and U5168 (N_5168,N_5023,N_5001);
nor U5169 (N_5169,N_5011,N_5025);
and U5170 (N_5170,N_5075,N_5063);
and U5171 (N_5171,N_5029,N_5043);
nor U5172 (N_5172,N_5098,N_5042);
or U5173 (N_5173,N_5041,N_5003);
or U5174 (N_5174,N_5054,N_5078);
and U5175 (N_5175,N_5036,N_5095);
or U5176 (N_5176,N_5010,N_5089);
nand U5177 (N_5177,N_5018,N_5009);
or U5178 (N_5178,N_5094,N_5046);
or U5179 (N_5179,N_5089,N_5086);
xnor U5180 (N_5180,N_5079,N_5037);
and U5181 (N_5181,N_5037,N_5090);
nand U5182 (N_5182,N_5015,N_5067);
nand U5183 (N_5183,N_5050,N_5058);
nand U5184 (N_5184,N_5066,N_5058);
nand U5185 (N_5185,N_5053,N_5017);
nor U5186 (N_5186,N_5088,N_5002);
or U5187 (N_5187,N_5077,N_5023);
and U5188 (N_5188,N_5027,N_5052);
nor U5189 (N_5189,N_5094,N_5020);
nand U5190 (N_5190,N_5072,N_5095);
nor U5191 (N_5191,N_5092,N_5096);
nor U5192 (N_5192,N_5030,N_5014);
xor U5193 (N_5193,N_5032,N_5085);
nand U5194 (N_5194,N_5046,N_5085);
nor U5195 (N_5195,N_5003,N_5027);
and U5196 (N_5196,N_5046,N_5096);
nand U5197 (N_5197,N_5001,N_5078);
and U5198 (N_5198,N_5081,N_5018);
nor U5199 (N_5199,N_5032,N_5055);
or U5200 (N_5200,N_5106,N_5130);
and U5201 (N_5201,N_5169,N_5197);
and U5202 (N_5202,N_5105,N_5167);
nand U5203 (N_5203,N_5175,N_5166);
nor U5204 (N_5204,N_5193,N_5156);
or U5205 (N_5205,N_5145,N_5126);
nor U5206 (N_5206,N_5109,N_5153);
and U5207 (N_5207,N_5194,N_5144);
nand U5208 (N_5208,N_5143,N_5186);
nor U5209 (N_5209,N_5136,N_5137);
and U5210 (N_5210,N_5168,N_5110);
or U5211 (N_5211,N_5149,N_5170);
nor U5212 (N_5212,N_5178,N_5114);
and U5213 (N_5213,N_5101,N_5176);
xnor U5214 (N_5214,N_5177,N_5117);
nor U5215 (N_5215,N_5115,N_5134);
or U5216 (N_5216,N_5171,N_5133);
nand U5217 (N_5217,N_5154,N_5174);
nor U5218 (N_5218,N_5199,N_5112);
or U5219 (N_5219,N_5128,N_5108);
and U5220 (N_5220,N_5119,N_5187);
and U5221 (N_5221,N_5165,N_5102);
nand U5222 (N_5222,N_5161,N_5122);
nor U5223 (N_5223,N_5118,N_5127);
xor U5224 (N_5224,N_5140,N_5159);
or U5225 (N_5225,N_5121,N_5173);
and U5226 (N_5226,N_5190,N_5185);
or U5227 (N_5227,N_5198,N_5129);
or U5228 (N_5228,N_5107,N_5103);
nand U5229 (N_5229,N_5151,N_5124);
and U5230 (N_5230,N_5164,N_5131);
and U5231 (N_5231,N_5111,N_5120);
xor U5232 (N_5232,N_5148,N_5142);
nor U5233 (N_5233,N_5162,N_5160);
nand U5234 (N_5234,N_5192,N_5195);
nand U5235 (N_5235,N_5100,N_5141);
xor U5236 (N_5236,N_5155,N_5181);
nor U5237 (N_5237,N_5183,N_5116);
or U5238 (N_5238,N_5157,N_5132);
and U5239 (N_5239,N_5135,N_5189);
nand U5240 (N_5240,N_5180,N_5158);
or U5241 (N_5241,N_5182,N_5191);
nand U5242 (N_5242,N_5184,N_5179);
nand U5243 (N_5243,N_5104,N_5123);
nor U5244 (N_5244,N_5147,N_5172);
nor U5245 (N_5245,N_5163,N_5188);
or U5246 (N_5246,N_5113,N_5139);
nand U5247 (N_5247,N_5146,N_5125);
nand U5248 (N_5248,N_5150,N_5196);
nand U5249 (N_5249,N_5138,N_5152);
nand U5250 (N_5250,N_5165,N_5132);
and U5251 (N_5251,N_5140,N_5160);
or U5252 (N_5252,N_5176,N_5110);
nor U5253 (N_5253,N_5150,N_5184);
nor U5254 (N_5254,N_5133,N_5122);
or U5255 (N_5255,N_5197,N_5147);
nand U5256 (N_5256,N_5155,N_5129);
nand U5257 (N_5257,N_5164,N_5178);
and U5258 (N_5258,N_5193,N_5174);
nand U5259 (N_5259,N_5159,N_5146);
and U5260 (N_5260,N_5151,N_5153);
xnor U5261 (N_5261,N_5182,N_5188);
and U5262 (N_5262,N_5173,N_5186);
nand U5263 (N_5263,N_5173,N_5179);
nor U5264 (N_5264,N_5187,N_5151);
and U5265 (N_5265,N_5190,N_5171);
and U5266 (N_5266,N_5159,N_5124);
or U5267 (N_5267,N_5121,N_5158);
or U5268 (N_5268,N_5142,N_5106);
and U5269 (N_5269,N_5116,N_5150);
and U5270 (N_5270,N_5194,N_5185);
and U5271 (N_5271,N_5158,N_5177);
or U5272 (N_5272,N_5133,N_5182);
nor U5273 (N_5273,N_5147,N_5164);
nor U5274 (N_5274,N_5112,N_5119);
xor U5275 (N_5275,N_5131,N_5110);
or U5276 (N_5276,N_5134,N_5188);
nand U5277 (N_5277,N_5193,N_5166);
nor U5278 (N_5278,N_5150,N_5129);
or U5279 (N_5279,N_5137,N_5185);
and U5280 (N_5280,N_5140,N_5128);
or U5281 (N_5281,N_5195,N_5184);
and U5282 (N_5282,N_5155,N_5198);
nand U5283 (N_5283,N_5130,N_5119);
nand U5284 (N_5284,N_5174,N_5115);
nor U5285 (N_5285,N_5170,N_5142);
nor U5286 (N_5286,N_5150,N_5139);
xor U5287 (N_5287,N_5162,N_5174);
nor U5288 (N_5288,N_5113,N_5114);
nand U5289 (N_5289,N_5148,N_5182);
or U5290 (N_5290,N_5100,N_5186);
nand U5291 (N_5291,N_5197,N_5125);
or U5292 (N_5292,N_5115,N_5184);
or U5293 (N_5293,N_5149,N_5115);
nor U5294 (N_5294,N_5177,N_5108);
and U5295 (N_5295,N_5169,N_5189);
nand U5296 (N_5296,N_5137,N_5182);
and U5297 (N_5297,N_5124,N_5148);
nor U5298 (N_5298,N_5126,N_5153);
nor U5299 (N_5299,N_5140,N_5192);
and U5300 (N_5300,N_5273,N_5270);
nand U5301 (N_5301,N_5254,N_5292);
and U5302 (N_5302,N_5243,N_5255);
nand U5303 (N_5303,N_5281,N_5221);
nor U5304 (N_5304,N_5204,N_5286);
or U5305 (N_5305,N_5282,N_5252);
nor U5306 (N_5306,N_5213,N_5232);
or U5307 (N_5307,N_5265,N_5290);
and U5308 (N_5308,N_5271,N_5212);
and U5309 (N_5309,N_5247,N_5256);
or U5310 (N_5310,N_5264,N_5283);
nand U5311 (N_5311,N_5298,N_5285);
or U5312 (N_5312,N_5246,N_5279);
and U5313 (N_5313,N_5280,N_5262);
and U5314 (N_5314,N_5234,N_5228);
and U5315 (N_5315,N_5261,N_5244);
nor U5316 (N_5316,N_5245,N_5297);
and U5317 (N_5317,N_5250,N_5291);
nor U5318 (N_5318,N_5293,N_5288);
nand U5319 (N_5319,N_5249,N_5241);
and U5320 (N_5320,N_5203,N_5269);
and U5321 (N_5321,N_5253,N_5216);
nand U5322 (N_5322,N_5251,N_5207);
nand U5323 (N_5323,N_5294,N_5258);
and U5324 (N_5324,N_5233,N_5259);
xor U5325 (N_5325,N_5202,N_5235);
nor U5326 (N_5326,N_5278,N_5225);
nand U5327 (N_5327,N_5231,N_5260);
or U5328 (N_5328,N_5200,N_5263);
nor U5329 (N_5329,N_5248,N_5287);
nor U5330 (N_5330,N_5284,N_5211);
nor U5331 (N_5331,N_5274,N_5296);
or U5332 (N_5332,N_5242,N_5209);
nand U5333 (N_5333,N_5238,N_5257);
nor U5334 (N_5334,N_5205,N_5227);
nor U5335 (N_5335,N_5220,N_5240);
nor U5336 (N_5336,N_5295,N_5236);
or U5337 (N_5337,N_5266,N_5223);
or U5338 (N_5338,N_5222,N_5208);
xnor U5339 (N_5339,N_5201,N_5224);
and U5340 (N_5340,N_5277,N_5226);
and U5341 (N_5341,N_5229,N_5206);
nor U5342 (N_5342,N_5299,N_5267);
and U5343 (N_5343,N_5210,N_5217);
nor U5344 (N_5344,N_5275,N_5289);
and U5345 (N_5345,N_5215,N_5214);
or U5346 (N_5346,N_5239,N_5272);
and U5347 (N_5347,N_5237,N_5276);
xnor U5348 (N_5348,N_5230,N_5218);
and U5349 (N_5349,N_5268,N_5219);
nor U5350 (N_5350,N_5207,N_5289);
and U5351 (N_5351,N_5204,N_5222);
and U5352 (N_5352,N_5200,N_5216);
and U5353 (N_5353,N_5243,N_5269);
and U5354 (N_5354,N_5278,N_5292);
and U5355 (N_5355,N_5222,N_5230);
and U5356 (N_5356,N_5280,N_5248);
or U5357 (N_5357,N_5231,N_5213);
nor U5358 (N_5358,N_5223,N_5216);
nand U5359 (N_5359,N_5210,N_5222);
nand U5360 (N_5360,N_5200,N_5220);
and U5361 (N_5361,N_5221,N_5239);
nand U5362 (N_5362,N_5298,N_5206);
or U5363 (N_5363,N_5268,N_5258);
or U5364 (N_5364,N_5286,N_5209);
or U5365 (N_5365,N_5279,N_5245);
nor U5366 (N_5366,N_5271,N_5229);
or U5367 (N_5367,N_5225,N_5290);
and U5368 (N_5368,N_5284,N_5261);
or U5369 (N_5369,N_5216,N_5298);
nor U5370 (N_5370,N_5219,N_5261);
or U5371 (N_5371,N_5236,N_5205);
xor U5372 (N_5372,N_5299,N_5273);
or U5373 (N_5373,N_5207,N_5296);
and U5374 (N_5374,N_5219,N_5254);
nand U5375 (N_5375,N_5276,N_5214);
nand U5376 (N_5376,N_5287,N_5265);
or U5377 (N_5377,N_5254,N_5267);
or U5378 (N_5378,N_5270,N_5215);
nand U5379 (N_5379,N_5228,N_5293);
or U5380 (N_5380,N_5223,N_5258);
and U5381 (N_5381,N_5225,N_5279);
and U5382 (N_5382,N_5239,N_5275);
and U5383 (N_5383,N_5219,N_5294);
or U5384 (N_5384,N_5233,N_5270);
and U5385 (N_5385,N_5229,N_5214);
nor U5386 (N_5386,N_5222,N_5252);
nand U5387 (N_5387,N_5280,N_5252);
or U5388 (N_5388,N_5278,N_5261);
nor U5389 (N_5389,N_5271,N_5276);
and U5390 (N_5390,N_5255,N_5295);
and U5391 (N_5391,N_5248,N_5216);
xor U5392 (N_5392,N_5220,N_5273);
and U5393 (N_5393,N_5222,N_5216);
nor U5394 (N_5394,N_5212,N_5259);
or U5395 (N_5395,N_5221,N_5242);
nand U5396 (N_5396,N_5285,N_5219);
nor U5397 (N_5397,N_5234,N_5229);
nand U5398 (N_5398,N_5297,N_5207);
and U5399 (N_5399,N_5219,N_5288);
and U5400 (N_5400,N_5371,N_5372);
xnor U5401 (N_5401,N_5302,N_5312);
nor U5402 (N_5402,N_5326,N_5380);
nand U5403 (N_5403,N_5313,N_5398);
or U5404 (N_5404,N_5325,N_5386);
nor U5405 (N_5405,N_5387,N_5365);
nor U5406 (N_5406,N_5314,N_5394);
nor U5407 (N_5407,N_5392,N_5355);
nand U5408 (N_5408,N_5342,N_5321);
and U5409 (N_5409,N_5337,N_5328);
xnor U5410 (N_5410,N_5399,N_5327);
or U5411 (N_5411,N_5360,N_5315);
nor U5412 (N_5412,N_5362,N_5332);
nand U5413 (N_5413,N_5357,N_5384);
and U5414 (N_5414,N_5334,N_5350);
or U5415 (N_5415,N_5366,N_5309);
or U5416 (N_5416,N_5329,N_5338);
and U5417 (N_5417,N_5318,N_5367);
or U5418 (N_5418,N_5359,N_5349);
and U5419 (N_5419,N_5310,N_5381);
and U5420 (N_5420,N_5391,N_5396);
or U5421 (N_5421,N_5333,N_5375);
xor U5422 (N_5422,N_5351,N_5356);
or U5423 (N_5423,N_5388,N_5378);
nand U5424 (N_5424,N_5361,N_5300);
and U5425 (N_5425,N_5305,N_5363);
nand U5426 (N_5426,N_5304,N_5323);
and U5427 (N_5427,N_5330,N_5320);
or U5428 (N_5428,N_5340,N_5335);
and U5429 (N_5429,N_5390,N_5341);
nand U5430 (N_5430,N_5358,N_5368);
nand U5431 (N_5431,N_5395,N_5370);
and U5432 (N_5432,N_5379,N_5397);
nand U5433 (N_5433,N_5343,N_5383);
nor U5434 (N_5434,N_5364,N_5345);
or U5435 (N_5435,N_5347,N_5308);
and U5436 (N_5436,N_5348,N_5382);
or U5437 (N_5437,N_5306,N_5373);
and U5438 (N_5438,N_5322,N_5353);
xnor U5439 (N_5439,N_5393,N_5352);
xnor U5440 (N_5440,N_5377,N_5331);
nor U5441 (N_5441,N_5339,N_5303);
and U5442 (N_5442,N_5385,N_5346);
nor U5443 (N_5443,N_5319,N_5324);
nor U5444 (N_5444,N_5389,N_5344);
nor U5445 (N_5445,N_5369,N_5311);
nand U5446 (N_5446,N_5354,N_5336);
or U5447 (N_5447,N_5316,N_5376);
nand U5448 (N_5448,N_5374,N_5307);
and U5449 (N_5449,N_5317,N_5301);
nand U5450 (N_5450,N_5392,N_5326);
and U5451 (N_5451,N_5349,N_5384);
or U5452 (N_5452,N_5310,N_5369);
and U5453 (N_5453,N_5300,N_5394);
or U5454 (N_5454,N_5354,N_5377);
nor U5455 (N_5455,N_5378,N_5344);
nor U5456 (N_5456,N_5348,N_5347);
nor U5457 (N_5457,N_5343,N_5326);
and U5458 (N_5458,N_5391,N_5386);
or U5459 (N_5459,N_5317,N_5314);
xnor U5460 (N_5460,N_5375,N_5376);
nand U5461 (N_5461,N_5366,N_5369);
nor U5462 (N_5462,N_5334,N_5352);
nand U5463 (N_5463,N_5303,N_5341);
nand U5464 (N_5464,N_5300,N_5318);
and U5465 (N_5465,N_5326,N_5319);
or U5466 (N_5466,N_5309,N_5347);
nor U5467 (N_5467,N_5386,N_5336);
nor U5468 (N_5468,N_5302,N_5353);
and U5469 (N_5469,N_5366,N_5315);
and U5470 (N_5470,N_5344,N_5326);
nand U5471 (N_5471,N_5324,N_5339);
or U5472 (N_5472,N_5394,N_5335);
and U5473 (N_5473,N_5336,N_5321);
nor U5474 (N_5474,N_5356,N_5361);
xnor U5475 (N_5475,N_5338,N_5387);
and U5476 (N_5476,N_5378,N_5305);
and U5477 (N_5477,N_5311,N_5334);
nor U5478 (N_5478,N_5346,N_5353);
or U5479 (N_5479,N_5398,N_5340);
nor U5480 (N_5480,N_5361,N_5326);
nand U5481 (N_5481,N_5370,N_5329);
and U5482 (N_5482,N_5397,N_5344);
nor U5483 (N_5483,N_5360,N_5324);
nand U5484 (N_5484,N_5375,N_5322);
nand U5485 (N_5485,N_5356,N_5329);
or U5486 (N_5486,N_5379,N_5332);
or U5487 (N_5487,N_5350,N_5347);
or U5488 (N_5488,N_5357,N_5351);
and U5489 (N_5489,N_5333,N_5376);
xnor U5490 (N_5490,N_5361,N_5357);
or U5491 (N_5491,N_5335,N_5314);
xnor U5492 (N_5492,N_5331,N_5395);
nor U5493 (N_5493,N_5380,N_5395);
nand U5494 (N_5494,N_5323,N_5322);
nand U5495 (N_5495,N_5315,N_5300);
nand U5496 (N_5496,N_5393,N_5381);
xnor U5497 (N_5497,N_5312,N_5329);
nor U5498 (N_5498,N_5346,N_5382);
nor U5499 (N_5499,N_5379,N_5392);
xnor U5500 (N_5500,N_5473,N_5448);
nor U5501 (N_5501,N_5457,N_5442);
and U5502 (N_5502,N_5495,N_5430);
or U5503 (N_5503,N_5431,N_5459);
nor U5504 (N_5504,N_5477,N_5452);
nor U5505 (N_5505,N_5446,N_5410);
xor U5506 (N_5506,N_5419,N_5440);
and U5507 (N_5507,N_5449,N_5428);
xnor U5508 (N_5508,N_5417,N_5484);
and U5509 (N_5509,N_5456,N_5407);
nand U5510 (N_5510,N_5409,N_5438);
nand U5511 (N_5511,N_5422,N_5474);
or U5512 (N_5512,N_5489,N_5445);
nor U5513 (N_5513,N_5411,N_5492);
nor U5514 (N_5514,N_5403,N_5404);
and U5515 (N_5515,N_5466,N_5468);
nand U5516 (N_5516,N_5485,N_5471);
nand U5517 (N_5517,N_5488,N_5481);
or U5518 (N_5518,N_5415,N_5453);
or U5519 (N_5519,N_5491,N_5494);
nand U5520 (N_5520,N_5434,N_5454);
nor U5521 (N_5521,N_5482,N_5406);
or U5522 (N_5522,N_5435,N_5443);
nor U5523 (N_5523,N_5401,N_5498);
and U5524 (N_5524,N_5447,N_5450);
or U5525 (N_5525,N_5424,N_5496);
nand U5526 (N_5526,N_5432,N_5423);
nor U5527 (N_5527,N_5475,N_5437);
or U5528 (N_5528,N_5467,N_5478);
and U5529 (N_5529,N_5408,N_5433);
and U5530 (N_5530,N_5497,N_5421);
and U5531 (N_5531,N_5426,N_5476);
nor U5532 (N_5532,N_5402,N_5487);
nor U5533 (N_5533,N_5479,N_5465);
nand U5534 (N_5534,N_5483,N_5472);
or U5535 (N_5535,N_5400,N_5486);
and U5536 (N_5536,N_5420,N_5441);
xnor U5537 (N_5537,N_5416,N_5436);
and U5538 (N_5538,N_5460,N_5490);
nand U5539 (N_5539,N_5464,N_5451);
nor U5540 (N_5540,N_5429,N_5462);
or U5541 (N_5541,N_5439,N_5461);
xnor U5542 (N_5542,N_5427,N_5444);
and U5543 (N_5543,N_5425,N_5463);
nor U5544 (N_5544,N_5455,N_5418);
and U5545 (N_5545,N_5499,N_5413);
xor U5546 (N_5546,N_5480,N_5458);
nand U5547 (N_5547,N_5470,N_5405);
nand U5548 (N_5548,N_5414,N_5469);
xor U5549 (N_5549,N_5412,N_5493);
and U5550 (N_5550,N_5487,N_5489);
nand U5551 (N_5551,N_5491,N_5477);
nand U5552 (N_5552,N_5419,N_5470);
and U5553 (N_5553,N_5483,N_5445);
and U5554 (N_5554,N_5453,N_5438);
and U5555 (N_5555,N_5467,N_5450);
or U5556 (N_5556,N_5490,N_5416);
nand U5557 (N_5557,N_5410,N_5422);
and U5558 (N_5558,N_5488,N_5446);
nor U5559 (N_5559,N_5493,N_5474);
nand U5560 (N_5560,N_5450,N_5474);
nand U5561 (N_5561,N_5473,N_5403);
and U5562 (N_5562,N_5487,N_5438);
and U5563 (N_5563,N_5433,N_5402);
nand U5564 (N_5564,N_5446,N_5493);
xnor U5565 (N_5565,N_5444,N_5441);
or U5566 (N_5566,N_5421,N_5498);
or U5567 (N_5567,N_5423,N_5465);
nand U5568 (N_5568,N_5496,N_5465);
and U5569 (N_5569,N_5448,N_5414);
xor U5570 (N_5570,N_5449,N_5408);
xor U5571 (N_5571,N_5486,N_5420);
nor U5572 (N_5572,N_5441,N_5424);
nand U5573 (N_5573,N_5410,N_5412);
nor U5574 (N_5574,N_5464,N_5480);
or U5575 (N_5575,N_5433,N_5406);
nand U5576 (N_5576,N_5441,N_5466);
nand U5577 (N_5577,N_5481,N_5498);
or U5578 (N_5578,N_5470,N_5437);
or U5579 (N_5579,N_5451,N_5420);
xnor U5580 (N_5580,N_5475,N_5426);
or U5581 (N_5581,N_5463,N_5431);
and U5582 (N_5582,N_5494,N_5407);
and U5583 (N_5583,N_5417,N_5406);
or U5584 (N_5584,N_5451,N_5462);
nand U5585 (N_5585,N_5451,N_5457);
nor U5586 (N_5586,N_5451,N_5428);
and U5587 (N_5587,N_5405,N_5463);
or U5588 (N_5588,N_5473,N_5487);
nand U5589 (N_5589,N_5498,N_5431);
nor U5590 (N_5590,N_5459,N_5442);
or U5591 (N_5591,N_5410,N_5423);
or U5592 (N_5592,N_5415,N_5428);
and U5593 (N_5593,N_5480,N_5475);
or U5594 (N_5594,N_5441,N_5464);
or U5595 (N_5595,N_5437,N_5407);
xor U5596 (N_5596,N_5499,N_5489);
xnor U5597 (N_5597,N_5402,N_5457);
and U5598 (N_5598,N_5407,N_5480);
nor U5599 (N_5599,N_5460,N_5499);
nand U5600 (N_5600,N_5568,N_5584);
xor U5601 (N_5601,N_5588,N_5523);
or U5602 (N_5602,N_5576,N_5507);
nand U5603 (N_5603,N_5549,N_5522);
or U5604 (N_5604,N_5515,N_5506);
nand U5605 (N_5605,N_5579,N_5575);
xnor U5606 (N_5606,N_5535,N_5578);
xnor U5607 (N_5607,N_5577,N_5503);
or U5608 (N_5608,N_5580,N_5542);
or U5609 (N_5609,N_5598,N_5557);
and U5610 (N_5610,N_5555,N_5534);
nand U5611 (N_5611,N_5596,N_5539);
xnor U5612 (N_5612,N_5513,N_5536);
xor U5613 (N_5613,N_5569,N_5512);
and U5614 (N_5614,N_5520,N_5566);
xor U5615 (N_5615,N_5543,N_5532);
nand U5616 (N_5616,N_5529,N_5531);
nand U5617 (N_5617,N_5551,N_5519);
xor U5618 (N_5618,N_5563,N_5502);
and U5619 (N_5619,N_5501,N_5504);
nand U5620 (N_5620,N_5525,N_5537);
nor U5621 (N_5621,N_5517,N_5527);
or U5622 (N_5622,N_5565,N_5589);
xor U5623 (N_5623,N_5516,N_5571);
nand U5624 (N_5624,N_5554,N_5528);
nor U5625 (N_5625,N_5594,N_5590);
nor U5626 (N_5626,N_5581,N_5548);
nand U5627 (N_5627,N_5544,N_5573);
nand U5628 (N_5628,N_5509,N_5591);
nand U5629 (N_5629,N_5592,N_5559);
nand U5630 (N_5630,N_5505,N_5541);
nand U5631 (N_5631,N_5524,N_5599);
and U5632 (N_5632,N_5582,N_5526);
or U5633 (N_5633,N_5538,N_5545);
nor U5634 (N_5634,N_5560,N_5500);
and U5635 (N_5635,N_5595,N_5561);
xor U5636 (N_5636,N_5593,N_5514);
or U5637 (N_5637,N_5540,N_5546);
and U5638 (N_5638,N_5558,N_5562);
and U5639 (N_5639,N_5552,N_5556);
nor U5640 (N_5640,N_5518,N_5587);
nor U5641 (N_5641,N_5521,N_5586);
and U5642 (N_5642,N_5533,N_5553);
or U5643 (N_5643,N_5508,N_5564);
or U5644 (N_5644,N_5547,N_5510);
xnor U5645 (N_5645,N_5530,N_5567);
and U5646 (N_5646,N_5511,N_5583);
nor U5647 (N_5647,N_5597,N_5570);
or U5648 (N_5648,N_5550,N_5585);
xnor U5649 (N_5649,N_5574,N_5572);
xor U5650 (N_5650,N_5595,N_5576);
or U5651 (N_5651,N_5572,N_5599);
and U5652 (N_5652,N_5523,N_5514);
or U5653 (N_5653,N_5578,N_5559);
nand U5654 (N_5654,N_5578,N_5539);
nand U5655 (N_5655,N_5552,N_5555);
or U5656 (N_5656,N_5551,N_5547);
xor U5657 (N_5657,N_5507,N_5595);
and U5658 (N_5658,N_5589,N_5530);
nand U5659 (N_5659,N_5543,N_5571);
or U5660 (N_5660,N_5536,N_5546);
nor U5661 (N_5661,N_5526,N_5591);
nor U5662 (N_5662,N_5589,N_5531);
or U5663 (N_5663,N_5529,N_5586);
nor U5664 (N_5664,N_5510,N_5515);
and U5665 (N_5665,N_5546,N_5545);
or U5666 (N_5666,N_5548,N_5585);
nand U5667 (N_5667,N_5557,N_5581);
and U5668 (N_5668,N_5578,N_5541);
and U5669 (N_5669,N_5503,N_5588);
nand U5670 (N_5670,N_5569,N_5576);
and U5671 (N_5671,N_5597,N_5591);
and U5672 (N_5672,N_5597,N_5558);
and U5673 (N_5673,N_5517,N_5574);
or U5674 (N_5674,N_5566,N_5569);
nand U5675 (N_5675,N_5507,N_5599);
xnor U5676 (N_5676,N_5576,N_5536);
nand U5677 (N_5677,N_5522,N_5518);
or U5678 (N_5678,N_5547,N_5589);
nor U5679 (N_5679,N_5522,N_5588);
xor U5680 (N_5680,N_5561,N_5566);
nor U5681 (N_5681,N_5527,N_5562);
and U5682 (N_5682,N_5567,N_5566);
and U5683 (N_5683,N_5598,N_5571);
or U5684 (N_5684,N_5519,N_5532);
or U5685 (N_5685,N_5543,N_5554);
nand U5686 (N_5686,N_5543,N_5531);
and U5687 (N_5687,N_5573,N_5583);
nand U5688 (N_5688,N_5508,N_5546);
nand U5689 (N_5689,N_5503,N_5523);
xor U5690 (N_5690,N_5591,N_5568);
nor U5691 (N_5691,N_5527,N_5578);
and U5692 (N_5692,N_5521,N_5520);
nor U5693 (N_5693,N_5519,N_5527);
or U5694 (N_5694,N_5534,N_5505);
xnor U5695 (N_5695,N_5560,N_5596);
xor U5696 (N_5696,N_5525,N_5510);
xnor U5697 (N_5697,N_5541,N_5506);
and U5698 (N_5698,N_5508,N_5584);
or U5699 (N_5699,N_5511,N_5571);
and U5700 (N_5700,N_5658,N_5656);
or U5701 (N_5701,N_5602,N_5623);
xor U5702 (N_5702,N_5606,N_5680);
and U5703 (N_5703,N_5644,N_5666);
and U5704 (N_5704,N_5635,N_5693);
nor U5705 (N_5705,N_5692,N_5636);
nand U5706 (N_5706,N_5682,N_5672);
nand U5707 (N_5707,N_5673,N_5696);
nor U5708 (N_5708,N_5657,N_5649);
or U5709 (N_5709,N_5664,N_5608);
nor U5710 (N_5710,N_5683,N_5605);
and U5711 (N_5711,N_5618,N_5652);
or U5712 (N_5712,N_5642,N_5612);
or U5713 (N_5713,N_5669,N_5622);
or U5714 (N_5714,N_5629,N_5681);
or U5715 (N_5715,N_5613,N_5600);
nand U5716 (N_5716,N_5616,N_5655);
nor U5717 (N_5717,N_5684,N_5625);
nand U5718 (N_5718,N_5626,N_5617);
nand U5719 (N_5719,N_5651,N_5695);
and U5720 (N_5720,N_5671,N_5633);
nor U5721 (N_5721,N_5674,N_5687);
and U5722 (N_5722,N_5638,N_5637);
nor U5723 (N_5723,N_5676,N_5641);
nor U5724 (N_5724,N_5694,N_5661);
nor U5725 (N_5725,N_5662,N_5610);
and U5726 (N_5726,N_5667,N_5631);
nor U5727 (N_5727,N_5632,N_5688);
xnor U5728 (N_5728,N_5691,N_5677);
nor U5729 (N_5729,N_5686,N_5670);
nand U5730 (N_5730,N_5690,N_5659);
nand U5731 (N_5731,N_5699,N_5627);
xor U5732 (N_5732,N_5648,N_5653);
and U5733 (N_5733,N_5685,N_5615);
xor U5734 (N_5734,N_5634,N_5650);
xor U5735 (N_5735,N_5609,N_5665);
nor U5736 (N_5736,N_5620,N_5645);
and U5737 (N_5737,N_5679,N_5630);
or U5738 (N_5738,N_5639,N_5624);
nand U5739 (N_5739,N_5647,N_5654);
nor U5740 (N_5740,N_5628,N_5663);
or U5741 (N_5741,N_5611,N_5619);
nor U5742 (N_5742,N_5614,N_5678);
and U5743 (N_5743,N_5646,N_5607);
nor U5744 (N_5744,N_5660,N_5668);
and U5745 (N_5745,N_5698,N_5601);
nand U5746 (N_5746,N_5643,N_5604);
and U5747 (N_5747,N_5689,N_5697);
nor U5748 (N_5748,N_5621,N_5640);
nand U5749 (N_5749,N_5675,N_5603);
and U5750 (N_5750,N_5602,N_5615);
and U5751 (N_5751,N_5687,N_5647);
or U5752 (N_5752,N_5647,N_5664);
and U5753 (N_5753,N_5685,N_5671);
nor U5754 (N_5754,N_5690,N_5619);
nor U5755 (N_5755,N_5643,N_5601);
nand U5756 (N_5756,N_5672,N_5613);
nand U5757 (N_5757,N_5621,N_5649);
or U5758 (N_5758,N_5676,N_5686);
or U5759 (N_5759,N_5616,N_5603);
nand U5760 (N_5760,N_5655,N_5626);
and U5761 (N_5761,N_5652,N_5687);
xor U5762 (N_5762,N_5645,N_5684);
xnor U5763 (N_5763,N_5667,N_5625);
or U5764 (N_5764,N_5618,N_5601);
or U5765 (N_5765,N_5617,N_5629);
or U5766 (N_5766,N_5640,N_5668);
or U5767 (N_5767,N_5665,N_5657);
or U5768 (N_5768,N_5613,N_5656);
and U5769 (N_5769,N_5671,N_5657);
and U5770 (N_5770,N_5652,N_5643);
and U5771 (N_5771,N_5689,N_5643);
nand U5772 (N_5772,N_5643,N_5685);
or U5773 (N_5773,N_5630,N_5611);
nor U5774 (N_5774,N_5601,N_5678);
or U5775 (N_5775,N_5627,N_5648);
and U5776 (N_5776,N_5653,N_5685);
xor U5777 (N_5777,N_5680,N_5602);
nor U5778 (N_5778,N_5600,N_5620);
or U5779 (N_5779,N_5689,N_5692);
or U5780 (N_5780,N_5680,N_5648);
and U5781 (N_5781,N_5617,N_5667);
nand U5782 (N_5782,N_5652,N_5635);
and U5783 (N_5783,N_5678,N_5634);
and U5784 (N_5784,N_5639,N_5601);
nor U5785 (N_5785,N_5611,N_5643);
or U5786 (N_5786,N_5628,N_5639);
and U5787 (N_5787,N_5606,N_5683);
and U5788 (N_5788,N_5637,N_5604);
nand U5789 (N_5789,N_5635,N_5604);
nand U5790 (N_5790,N_5600,N_5684);
nor U5791 (N_5791,N_5637,N_5694);
xnor U5792 (N_5792,N_5637,N_5662);
and U5793 (N_5793,N_5678,N_5635);
nor U5794 (N_5794,N_5653,N_5644);
and U5795 (N_5795,N_5647,N_5631);
and U5796 (N_5796,N_5695,N_5653);
and U5797 (N_5797,N_5673,N_5672);
nand U5798 (N_5798,N_5673,N_5654);
xor U5799 (N_5799,N_5654,N_5622);
and U5800 (N_5800,N_5727,N_5720);
or U5801 (N_5801,N_5776,N_5704);
nor U5802 (N_5802,N_5778,N_5761);
and U5803 (N_5803,N_5702,N_5754);
or U5804 (N_5804,N_5707,N_5743);
and U5805 (N_5805,N_5755,N_5701);
nand U5806 (N_5806,N_5722,N_5758);
xor U5807 (N_5807,N_5737,N_5738);
nand U5808 (N_5808,N_5762,N_5712);
or U5809 (N_5809,N_5732,N_5751);
or U5810 (N_5810,N_5765,N_5793);
and U5811 (N_5811,N_5724,N_5796);
nor U5812 (N_5812,N_5794,N_5708);
and U5813 (N_5813,N_5786,N_5757);
or U5814 (N_5814,N_5716,N_5760);
or U5815 (N_5815,N_5753,N_5798);
nand U5816 (N_5816,N_5723,N_5779);
nand U5817 (N_5817,N_5739,N_5797);
nand U5818 (N_5818,N_5766,N_5767);
nor U5819 (N_5819,N_5717,N_5714);
nand U5820 (N_5820,N_5773,N_5742);
nor U5821 (N_5821,N_5740,N_5782);
xnor U5822 (N_5822,N_5731,N_5700);
or U5823 (N_5823,N_5777,N_5772);
nor U5824 (N_5824,N_5735,N_5728);
nand U5825 (N_5825,N_5703,N_5750);
and U5826 (N_5826,N_5706,N_5715);
or U5827 (N_5827,N_5780,N_5736);
nand U5828 (N_5828,N_5729,N_5792);
or U5829 (N_5829,N_5734,N_5771);
nand U5830 (N_5830,N_5787,N_5788);
or U5831 (N_5831,N_5774,N_5745);
and U5832 (N_5832,N_5713,N_5781);
or U5833 (N_5833,N_5783,N_5770);
nand U5834 (N_5834,N_5752,N_5763);
xnor U5835 (N_5835,N_5759,N_5799);
nor U5836 (N_5836,N_5764,N_5709);
nand U5837 (N_5837,N_5790,N_5784);
nor U5838 (N_5838,N_5705,N_5730);
or U5839 (N_5839,N_5718,N_5725);
nor U5840 (N_5840,N_5775,N_5710);
or U5841 (N_5841,N_5748,N_5719);
and U5842 (N_5842,N_5795,N_5744);
nand U5843 (N_5843,N_5747,N_5791);
or U5844 (N_5844,N_5756,N_5726);
or U5845 (N_5845,N_5741,N_5789);
and U5846 (N_5846,N_5711,N_5769);
xnor U5847 (N_5847,N_5721,N_5733);
nand U5848 (N_5848,N_5746,N_5749);
and U5849 (N_5849,N_5768,N_5785);
nand U5850 (N_5850,N_5747,N_5752);
nor U5851 (N_5851,N_5756,N_5794);
nand U5852 (N_5852,N_5719,N_5741);
nor U5853 (N_5853,N_5757,N_5733);
xor U5854 (N_5854,N_5721,N_5738);
nand U5855 (N_5855,N_5759,N_5724);
nand U5856 (N_5856,N_5780,N_5739);
or U5857 (N_5857,N_5704,N_5749);
xor U5858 (N_5858,N_5707,N_5789);
nand U5859 (N_5859,N_5771,N_5784);
and U5860 (N_5860,N_5717,N_5776);
or U5861 (N_5861,N_5719,N_5749);
nor U5862 (N_5862,N_5732,N_5774);
and U5863 (N_5863,N_5730,N_5707);
or U5864 (N_5864,N_5751,N_5737);
nor U5865 (N_5865,N_5769,N_5780);
nor U5866 (N_5866,N_5758,N_5709);
and U5867 (N_5867,N_5785,N_5775);
or U5868 (N_5868,N_5772,N_5756);
nand U5869 (N_5869,N_5713,N_5759);
nor U5870 (N_5870,N_5777,N_5723);
nor U5871 (N_5871,N_5761,N_5770);
and U5872 (N_5872,N_5766,N_5771);
or U5873 (N_5873,N_5735,N_5760);
or U5874 (N_5874,N_5797,N_5751);
and U5875 (N_5875,N_5759,N_5726);
xor U5876 (N_5876,N_5795,N_5785);
and U5877 (N_5877,N_5730,N_5716);
and U5878 (N_5878,N_5769,N_5708);
or U5879 (N_5879,N_5757,N_5797);
or U5880 (N_5880,N_5763,N_5743);
or U5881 (N_5881,N_5776,N_5768);
nor U5882 (N_5882,N_5709,N_5791);
nor U5883 (N_5883,N_5709,N_5701);
nor U5884 (N_5884,N_5752,N_5703);
or U5885 (N_5885,N_5754,N_5735);
or U5886 (N_5886,N_5747,N_5731);
nand U5887 (N_5887,N_5757,N_5784);
or U5888 (N_5888,N_5706,N_5734);
nor U5889 (N_5889,N_5788,N_5727);
or U5890 (N_5890,N_5761,N_5701);
nand U5891 (N_5891,N_5799,N_5780);
xnor U5892 (N_5892,N_5714,N_5785);
or U5893 (N_5893,N_5724,N_5761);
or U5894 (N_5894,N_5789,N_5732);
nor U5895 (N_5895,N_5740,N_5783);
nand U5896 (N_5896,N_5794,N_5764);
nand U5897 (N_5897,N_5737,N_5741);
or U5898 (N_5898,N_5795,N_5724);
nand U5899 (N_5899,N_5732,N_5785);
or U5900 (N_5900,N_5886,N_5899);
nand U5901 (N_5901,N_5871,N_5861);
or U5902 (N_5902,N_5832,N_5888);
nand U5903 (N_5903,N_5838,N_5821);
or U5904 (N_5904,N_5874,N_5810);
and U5905 (N_5905,N_5815,N_5820);
nand U5906 (N_5906,N_5893,N_5822);
and U5907 (N_5907,N_5812,N_5840);
xnor U5908 (N_5908,N_5885,N_5864);
nor U5909 (N_5909,N_5870,N_5826);
nand U5910 (N_5910,N_5839,N_5866);
xor U5911 (N_5911,N_5828,N_5860);
nor U5912 (N_5912,N_5887,N_5804);
and U5913 (N_5913,N_5849,N_5836);
nand U5914 (N_5914,N_5805,N_5831);
nand U5915 (N_5915,N_5894,N_5825);
and U5916 (N_5916,N_5813,N_5800);
and U5917 (N_5917,N_5803,N_5869);
and U5918 (N_5918,N_5881,N_5848);
or U5919 (N_5919,N_5867,N_5806);
or U5920 (N_5920,N_5814,N_5837);
and U5921 (N_5921,N_5817,N_5880);
or U5922 (N_5922,N_5863,N_5823);
and U5923 (N_5923,N_5842,N_5873);
nor U5924 (N_5924,N_5895,N_5850);
nor U5925 (N_5925,N_5879,N_5816);
and U5926 (N_5926,N_5856,N_5876);
or U5927 (N_5927,N_5896,N_5851);
nand U5928 (N_5928,N_5834,N_5875);
nor U5929 (N_5929,N_5808,N_5854);
and U5930 (N_5930,N_5890,N_5855);
and U5931 (N_5931,N_5882,N_5807);
nand U5932 (N_5932,N_5884,N_5819);
or U5933 (N_5933,N_5830,N_5847);
and U5934 (N_5934,N_5868,N_5862);
nand U5935 (N_5935,N_5827,N_5889);
or U5936 (N_5936,N_5898,N_5844);
nand U5937 (N_5937,N_5853,N_5883);
or U5938 (N_5938,N_5811,N_5801);
or U5939 (N_5939,N_5835,N_5843);
xor U5940 (N_5940,N_5833,N_5892);
nand U5941 (N_5941,N_5845,N_5877);
or U5942 (N_5942,N_5802,N_5846);
xnor U5943 (N_5943,N_5865,N_5872);
nand U5944 (N_5944,N_5857,N_5809);
nor U5945 (N_5945,N_5818,N_5824);
nand U5946 (N_5946,N_5841,N_5829);
nor U5947 (N_5947,N_5891,N_5897);
and U5948 (N_5948,N_5858,N_5859);
nand U5949 (N_5949,N_5878,N_5852);
nor U5950 (N_5950,N_5819,N_5837);
or U5951 (N_5951,N_5868,N_5855);
nor U5952 (N_5952,N_5829,N_5899);
nand U5953 (N_5953,N_5874,N_5892);
nand U5954 (N_5954,N_5855,N_5882);
nor U5955 (N_5955,N_5849,N_5880);
nor U5956 (N_5956,N_5885,N_5842);
and U5957 (N_5957,N_5885,N_5865);
or U5958 (N_5958,N_5880,N_5848);
nand U5959 (N_5959,N_5855,N_5822);
nor U5960 (N_5960,N_5835,N_5849);
or U5961 (N_5961,N_5854,N_5800);
xnor U5962 (N_5962,N_5831,N_5891);
or U5963 (N_5963,N_5868,N_5874);
or U5964 (N_5964,N_5895,N_5854);
xor U5965 (N_5965,N_5883,N_5863);
and U5966 (N_5966,N_5885,N_5835);
nor U5967 (N_5967,N_5811,N_5888);
xnor U5968 (N_5968,N_5886,N_5887);
nand U5969 (N_5969,N_5835,N_5898);
or U5970 (N_5970,N_5868,N_5813);
nor U5971 (N_5971,N_5868,N_5809);
and U5972 (N_5972,N_5810,N_5886);
and U5973 (N_5973,N_5852,N_5831);
nand U5974 (N_5974,N_5861,N_5827);
or U5975 (N_5975,N_5885,N_5804);
nor U5976 (N_5976,N_5883,N_5864);
xnor U5977 (N_5977,N_5851,N_5857);
nor U5978 (N_5978,N_5844,N_5881);
or U5979 (N_5979,N_5875,N_5841);
or U5980 (N_5980,N_5884,N_5878);
nor U5981 (N_5981,N_5888,N_5834);
nor U5982 (N_5982,N_5893,N_5829);
and U5983 (N_5983,N_5820,N_5853);
or U5984 (N_5984,N_5855,N_5823);
nor U5985 (N_5985,N_5814,N_5825);
or U5986 (N_5986,N_5812,N_5813);
nor U5987 (N_5987,N_5842,N_5809);
nand U5988 (N_5988,N_5897,N_5806);
xnor U5989 (N_5989,N_5853,N_5841);
nand U5990 (N_5990,N_5884,N_5868);
or U5991 (N_5991,N_5898,N_5897);
and U5992 (N_5992,N_5853,N_5891);
and U5993 (N_5993,N_5805,N_5863);
or U5994 (N_5994,N_5815,N_5840);
or U5995 (N_5995,N_5826,N_5865);
nor U5996 (N_5996,N_5853,N_5866);
and U5997 (N_5997,N_5815,N_5894);
nand U5998 (N_5998,N_5899,N_5865);
or U5999 (N_5999,N_5832,N_5833);
and U6000 (N_6000,N_5941,N_5950);
nor U6001 (N_6001,N_5968,N_5944);
xnor U6002 (N_6002,N_5978,N_5981);
nor U6003 (N_6003,N_5923,N_5984);
nand U6004 (N_6004,N_5952,N_5917);
or U6005 (N_6005,N_5908,N_5966);
or U6006 (N_6006,N_5976,N_5913);
nor U6007 (N_6007,N_5988,N_5906);
and U6008 (N_6008,N_5982,N_5971);
nand U6009 (N_6009,N_5947,N_5965);
nor U6010 (N_6010,N_5929,N_5959);
nor U6011 (N_6011,N_5951,N_5905);
and U6012 (N_6012,N_5922,N_5914);
nor U6013 (N_6013,N_5933,N_5928);
and U6014 (N_6014,N_5920,N_5937);
nand U6015 (N_6015,N_5915,N_5919);
nor U6016 (N_6016,N_5991,N_5935);
or U6017 (N_6017,N_5942,N_5975);
nor U6018 (N_6018,N_5945,N_5980);
nand U6019 (N_6019,N_5996,N_5961);
or U6020 (N_6020,N_5967,N_5946);
nand U6021 (N_6021,N_5958,N_5932);
nand U6022 (N_6022,N_5902,N_5964);
nor U6023 (N_6023,N_5960,N_5910);
nand U6024 (N_6024,N_5948,N_5977);
xnor U6025 (N_6025,N_5916,N_5953);
nor U6026 (N_6026,N_5992,N_5911);
or U6027 (N_6027,N_5912,N_5985);
nand U6028 (N_6028,N_5990,N_5927);
nor U6029 (N_6029,N_5999,N_5957);
and U6030 (N_6030,N_5903,N_5970);
or U6031 (N_6031,N_5936,N_5997);
or U6032 (N_6032,N_5921,N_5938);
nand U6033 (N_6033,N_5973,N_5986);
and U6034 (N_6034,N_5979,N_5924);
xnor U6035 (N_6035,N_5974,N_5925);
nor U6036 (N_6036,N_5901,N_5949);
and U6037 (N_6037,N_5962,N_5907);
xor U6038 (N_6038,N_5995,N_5900);
or U6039 (N_6039,N_5994,N_5989);
nand U6040 (N_6040,N_5955,N_5931);
nand U6041 (N_6041,N_5987,N_5943);
nor U6042 (N_6042,N_5954,N_5993);
nand U6043 (N_6043,N_5939,N_5930);
nor U6044 (N_6044,N_5904,N_5934);
nor U6045 (N_6045,N_5909,N_5969);
and U6046 (N_6046,N_5918,N_5926);
xor U6047 (N_6047,N_5972,N_5983);
xor U6048 (N_6048,N_5940,N_5956);
xor U6049 (N_6049,N_5963,N_5998);
and U6050 (N_6050,N_5938,N_5992);
or U6051 (N_6051,N_5905,N_5971);
xor U6052 (N_6052,N_5954,N_5926);
and U6053 (N_6053,N_5995,N_5956);
nor U6054 (N_6054,N_5954,N_5985);
xnor U6055 (N_6055,N_5905,N_5940);
nand U6056 (N_6056,N_5976,N_5961);
xor U6057 (N_6057,N_5942,N_5958);
and U6058 (N_6058,N_5983,N_5968);
and U6059 (N_6059,N_5951,N_5964);
xor U6060 (N_6060,N_5957,N_5910);
nor U6061 (N_6061,N_5928,N_5944);
nand U6062 (N_6062,N_5958,N_5914);
nor U6063 (N_6063,N_5958,N_5948);
nor U6064 (N_6064,N_5964,N_5990);
xnor U6065 (N_6065,N_5995,N_5922);
or U6066 (N_6066,N_5962,N_5985);
or U6067 (N_6067,N_5997,N_5952);
nor U6068 (N_6068,N_5905,N_5987);
or U6069 (N_6069,N_5991,N_5968);
or U6070 (N_6070,N_5941,N_5907);
and U6071 (N_6071,N_5959,N_5915);
or U6072 (N_6072,N_5967,N_5994);
nand U6073 (N_6073,N_5972,N_5982);
nor U6074 (N_6074,N_5957,N_5911);
and U6075 (N_6075,N_5940,N_5992);
nand U6076 (N_6076,N_5985,N_5935);
nor U6077 (N_6077,N_5901,N_5986);
nand U6078 (N_6078,N_5962,N_5952);
nand U6079 (N_6079,N_5998,N_5924);
and U6080 (N_6080,N_5959,N_5946);
nor U6081 (N_6081,N_5909,N_5995);
or U6082 (N_6082,N_5992,N_5994);
nor U6083 (N_6083,N_5947,N_5914);
nor U6084 (N_6084,N_5910,N_5903);
xnor U6085 (N_6085,N_5967,N_5972);
nor U6086 (N_6086,N_5989,N_5976);
and U6087 (N_6087,N_5985,N_5965);
or U6088 (N_6088,N_5977,N_5992);
nor U6089 (N_6089,N_5928,N_5965);
nand U6090 (N_6090,N_5913,N_5910);
and U6091 (N_6091,N_5997,N_5989);
xnor U6092 (N_6092,N_5948,N_5952);
and U6093 (N_6093,N_5991,N_5990);
and U6094 (N_6094,N_5927,N_5952);
nand U6095 (N_6095,N_5943,N_5921);
nand U6096 (N_6096,N_5974,N_5932);
and U6097 (N_6097,N_5934,N_5910);
or U6098 (N_6098,N_5914,N_5935);
or U6099 (N_6099,N_5908,N_5984);
nor U6100 (N_6100,N_6001,N_6011);
or U6101 (N_6101,N_6034,N_6095);
nor U6102 (N_6102,N_6022,N_6039);
or U6103 (N_6103,N_6042,N_6007);
nor U6104 (N_6104,N_6056,N_6040);
and U6105 (N_6105,N_6072,N_6093);
and U6106 (N_6106,N_6053,N_6012);
nand U6107 (N_6107,N_6018,N_6008);
xnor U6108 (N_6108,N_6021,N_6009);
or U6109 (N_6109,N_6047,N_6055);
xnor U6110 (N_6110,N_6028,N_6010);
nand U6111 (N_6111,N_6014,N_6019);
or U6112 (N_6112,N_6045,N_6086);
xor U6113 (N_6113,N_6067,N_6080);
nand U6114 (N_6114,N_6091,N_6025);
nand U6115 (N_6115,N_6063,N_6015);
and U6116 (N_6116,N_6030,N_6006);
and U6117 (N_6117,N_6016,N_6046);
nand U6118 (N_6118,N_6043,N_6033);
nand U6119 (N_6119,N_6004,N_6085);
nand U6120 (N_6120,N_6069,N_6092);
or U6121 (N_6121,N_6079,N_6081);
or U6122 (N_6122,N_6057,N_6099);
and U6123 (N_6123,N_6089,N_6027);
nor U6124 (N_6124,N_6097,N_6084);
nor U6125 (N_6125,N_6082,N_6071);
or U6126 (N_6126,N_6044,N_6017);
nor U6127 (N_6127,N_6098,N_6029);
nor U6128 (N_6128,N_6078,N_6074);
and U6129 (N_6129,N_6096,N_6094);
and U6130 (N_6130,N_6041,N_6061);
or U6131 (N_6131,N_6038,N_6005);
and U6132 (N_6132,N_6003,N_6060);
and U6133 (N_6133,N_6050,N_6020);
nand U6134 (N_6134,N_6023,N_6077);
xor U6135 (N_6135,N_6064,N_6088);
and U6136 (N_6136,N_6037,N_6070);
and U6137 (N_6137,N_6076,N_6052);
nor U6138 (N_6138,N_6051,N_6059);
and U6139 (N_6139,N_6087,N_6090);
or U6140 (N_6140,N_6073,N_6002);
nand U6141 (N_6141,N_6066,N_6035);
and U6142 (N_6142,N_6062,N_6024);
nor U6143 (N_6143,N_6068,N_6049);
nor U6144 (N_6144,N_6048,N_6054);
nand U6145 (N_6145,N_6065,N_6036);
and U6146 (N_6146,N_6013,N_6032);
nor U6147 (N_6147,N_6026,N_6083);
nand U6148 (N_6148,N_6000,N_6031);
and U6149 (N_6149,N_6058,N_6075);
nand U6150 (N_6150,N_6019,N_6026);
and U6151 (N_6151,N_6032,N_6002);
nor U6152 (N_6152,N_6061,N_6034);
nand U6153 (N_6153,N_6012,N_6038);
and U6154 (N_6154,N_6068,N_6083);
nor U6155 (N_6155,N_6021,N_6047);
nor U6156 (N_6156,N_6070,N_6067);
nand U6157 (N_6157,N_6030,N_6043);
nand U6158 (N_6158,N_6067,N_6082);
and U6159 (N_6159,N_6012,N_6098);
xnor U6160 (N_6160,N_6041,N_6001);
or U6161 (N_6161,N_6000,N_6005);
nor U6162 (N_6162,N_6054,N_6034);
nand U6163 (N_6163,N_6024,N_6034);
nor U6164 (N_6164,N_6059,N_6003);
or U6165 (N_6165,N_6086,N_6054);
and U6166 (N_6166,N_6085,N_6002);
nand U6167 (N_6167,N_6019,N_6007);
nor U6168 (N_6168,N_6035,N_6063);
and U6169 (N_6169,N_6023,N_6034);
nor U6170 (N_6170,N_6064,N_6092);
nand U6171 (N_6171,N_6043,N_6056);
nand U6172 (N_6172,N_6063,N_6096);
or U6173 (N_6173,N_6098,N_6062);
nor U6174 (N_6174,N_6035,N_6056);
or U6175 (N_6175,N_6043,N_6031);
nand U6176 (N_6176,N_6010,N_6093);
nor U6177 (N_6177,N_6054,N_6060);
nor U6178 (N_6178,N_6045,N_6028);
nand U6179 (N_6179,N_6046,N_6082);
or U6180 (N_6180,N_6042,N_6079);
xnor U6181 (N_6181,N_6099,N_6013);
nand U6182 (N_6182,N_6064,N_6021);
nor U6183 (N_6183,N_6009,N_6026);
nand U6184 (N_6184,N_6095,N_6005);
nand U6185 (N_6185,N_6006,N_6073);
or U6186 (N_6186,N_6006,N_6032);
or U6187 (N_6187,N_6056,N_6054);
or U6188 (N_6188,N_6065,N_6004);
or U6189 (N_6189,N_6056,N_6027);
nor U6190 (N_6190,N_6081,N_6028);
or U6191 (N_6191,N_6020,N_6098);
or U6192 (N_6192,N_6040,N_6039);
nand U6193 (N_6193,N_6041,N_6076);
nor U6194 (N_6194,N_6092,N_6001);
and U6195 (N_6195,N_6092,N_6082);
or U6196 (N_6196,N_6057,N_6024);
and U6197 (N_6197,N_6086,N_6075);
nand U6198 (N_6198,N_6050,N_6038);
or U6199 (N_6199,N_6038,N_6070);
xor U6200 (N_6200,N_6116,N_6184);
nor U6201 (N_6201,N_6182,N_6123);
nor U6202 (N_6202,N_6100,N_6103);
nor U6203 (N_6203,N_6136,N_6124);
nor U6204 (N_6204,N_6126,N_6185);
or U6205 (N_6205,N_6158,N_6189);
nor U6206 (N_6206,N_6161,N_6131);
nor U6207 (N_6207,N_6178,N_6176);
and U6208 (N_6208,N_6191,N_6110);
and U6209 (N_6209,N_6127,N_6135);
and U6210 (N_6210,N_6198,N_6190);
nand U6211 (N_6211,N_6105,N_6199);
xor U6212 (N_6212,N_6129,N_6119);
nand U6213 (N_6213,N_6114,N_6192);
nor U6214 (N_6214,N_6106,N_6156);
nand U6215 (N_6215,N_6164,N_6170);
and U6216 (N_6216,N_6138,N_6115);
nor U6217 (N_6217,N_6187,N_6162);
nor U6218 (N_6218,N_6142,N_6153);
nor U6219 (N_6219,N_6148,N_6188);
nand U6220 (N_6220,N_6167,N_6137);
or U6221 (N_6221,N_6173,N_6165);
and U6222 (N_6222,N_6108,N_6125);
nor U6223 (N_6223,N_6134,N_6147);
or U6224 (N_6224,N_6171,N_6195);
xnor U6225 (N_6225,N_6139,N_6120);
or U6226 (N_6226,N_6193,N_6163);
nor U6227 (N_6227,N_6104,N_6102);
nand U6228 (N_6228,N_6183,N_6101);
or U6229 (N_6229,N_6196,N_6133);
xnor U6230 (N_6230,N_6118,N_6112);
and U6231 (N_6231,N_6157,N_6155);
nand U6232 (N_6232,N_6122,N_6111);
nor U6233 (N_6233,N_6169,N_6179);
nand U6234 (N_6234,N_6194,N_6107);
nand U6235 (N_6235,N_6175,N_6128);
xnor U6236 (N_6236,N_6121,N_6151);
nand U6237 (N_6237,N_6168,N_6186);
nor U6238 (N_6238,N_6143,N_6150);
and U6239 (N_6239,N_6160,N_6166);
nand U6240 (N_6240,N_6159,N_6130);
nor U6241 (N_6241,N_6132,N_6141);
xor U6242 (N_6242,N_6152,N_6181);
nand U6243 (N_6243,N_6144,N_6177);
or U6244 (N_6244,N_6174,N_6117);
nor U6245 (N_6245,N_6197,N_6140);
and U6246 (N_6246,N_6146,N_6172);
or U6247 (N_6247,N_6109,N_6180);
xor U6248 (N_6248,N_6149,N_6113);
xor U6249 (N_6249,N_6145,N_6154);
and U6250 (N_6250,N_6110,N_6187);
nand U6251 (N_6251,N_6140,N_6101);
and U6252 (N_6252,N_6125,N_6127);
and U6253 (N_6253,N_6113,N_6137);
or U6254 (N_6254,N_6194,N_6198);
and U6255 (N_6255,N_6115,N_6132);
nand U6256 (N_6256,N_6133,N_6103);
nor U6257 (N_6257,N_6144,N_6169);
nor U6258 (N_6258,N_6199,N_6130);
or U6259 (N_6259,N_6183,N_6102);
and U6260 (N_6260,N_6186,N_6175);
nor U6261 (N_6261,N_6158,N_6106);
and U6262 (N_6262,N_6199,N_6193);
or U6263 (N_6263,N_6147,N_6158);
or U6264 (N_6264,N_6120,N_6163);
nor U6265 (N_6265,N_6129,N_6171);
or U6266 (N_6266,N_6154,N_6132);
or U6267 (N_6267,N_6124,N_6110);
or U6268 (N_6268,N_6148,N_6144);
nor U6269 (N_6269,N_6168,N_6167);
or U6270 (N_6270,N_6194,N_6181);
and U6271 (N_6271,N_6137,N_6189);
nand U6272 (N_6272,N_6145,N_6196);
or U6273 (N_6273,N_6144,N_6182);
nor U6274 (N_6274,N_6153,N_6156);
xor U6275 (N_6275,N_6130,N_6110);
xnor U6276 (N_6276,N_6186,N_6177);
nor U6277 (N_6277,N_6166,N_6111);
xor U6278 (N_6278,N_6183,N_6116);
and U6279 (N_6279,N_6177,N_6161);
or U6280 (N_6280,N_6112,N_6101);
or U6281 (N_6281,N_6174,N_6176);
nand U6282 (N_6282,N_6170,N_6106);
xnor U6283 (N_6283,N_6142,N_6185);
nand U6284 (N_6284,N_6175,N_6152);
and U6285 (N_6285,N_6109,N_6113);
nand U6286 (N_6286,N_6130,N_6139);
and U6287 (N_6287,N_6141,N_6114);
or U6288 (N_6288,N_6145,N_6185);
nand U6289 (N_6289,N_6194,N_6100);
and U6290 (N_6290,N_6147,N_6116);
nand U6291 (N_6291,N_6177,N_6129);
nand U6292 (N_6292,N_6115,N_6158);
and U6293 (N_6293,N_6192,N_6193);
nor U6294 (N_6294,N_6177,N_6189);
nor U6295 (N_6295,N_6195,N_6181);
or U6296 (N_6296,N_6191,N_6159);
nor U6297 (N_6297,N_6165,N_6109);
or U6298 (N_6298,N_6188,N_6130);
xnor U6299 (N_6299,N_6121,N_6191);
or U6300 (N_6300,N_6269,N_6277);
or U6301 (N_6301,N_6224,N_6268);
xor U6302 (N_6302,N_6209,N_6204);
or U6303 (N_6303,N_6203,N_6258);
and U6304 (N_6304,N_6267,N_6275);
or U6305 (N_6305,N_6281,N_6295);
nand U6306 (N_6306,N_6208,N_6256);
nand U6307 (N_6307,N_6261,N_6244);
and U6308 (N_6308,N_6255,N_6252);
and U6309 (N_6309,N_6290,N_6214);
and U6310 (N_6310,N_6202,N_6232);
and U6311 (N_6311,N_6279,N_6219);
nor U6312 (N_6312,N_6207,N_6238);
nand U6313 (N_6313,N_6286,N_6270);
or U6314 (N_6314,N_6220,N_6212);
nand U6315 (N_6315,N_6240,N_6278);
or U6316 (N_6316,N_6205,N_6235);
nor U6317 (N_6317,N_6284,N_6210);
or U6318 (N_6318,N_6222,N_6274);
or U6319 (N_6319,N_6213,N_6236);
nor U6320 (N_6320,N_6216,N_6226);
nand U6321 (N_6321,N_6296,N_6289);
nand U6322 (N_6322,N_6294,N_6237);
or U6323 (N_6323,N_6234,N_6266);
nor U6324 (N_6324,N_6283,N_6221);
nand U6325 (N_6325,N_6271,N_6265);
nor U6326 (N_6326,N_6227,N_6282);
or U6327 (N_6327,N_6239,N_6262);
or U6328 (N_6328,N_6251,N_6280);
or U6329 (N_6329,N_6217,N_6287);
nor U6330 (N_6330,N_6242,N_6245);
and U6331 (N_6331,N_6292,N_6285);
and U6332 (N_6332,N_6250,N_6288);
nand U6333 (N_6333,N_6206,N_6247);
nor U6334 (N_6334,N_6228,N_6230);
and U6335 (N_6335,N_6259,N_6218);
or U6336 (N_6336,N_6297,N_6241);
or U6337 (N_6337,N_6254,N_6263);
nor U6338 (N_6338,N_6273,N_6225);
or U6339 (N_6339,N_6249,N_6243);
and U6340 (N_6340,N_6211,N_6231);
nor U6341 (N_6341,N_6233,N_6298);
nand U6342 (N_6342,N_6215,N_6246);
nor U6343 (N_6343,N_6223,N_6257);
and U6344 (N_6344,N_6291,N_6264);
nor U6345 (N_6345,N_6276,N_6201);
nand U6346 (N_6346,N_6248,N_6260);
nand U6347 (N_6347,N_6200,N_6253);
nand U6348 (N_6348,N_6293,N_6272);
and U6349 (N_6349,N_6299,N_6229);
nor U6350 (N_6350,N_6210,N_6229);
and U6351 (N_6351,N_6204,N_6288);
nand U6352 (N_6352,N_6211,N_6207);
or U6353 (N_6353,N_6219,N_6280);
nor U6354 (N_6354,N_6273,N_6242);
and U6355 (N_6355,N_6289,N_6227);
nor U6356 (N_6356,N_6281,N_6215);
nand U6357 (N_6357,N_6287,N_6279);
nor U6358 (N_6358,N_6207,N_6223);
and U6359 (N_6359,N_6238,N_6223);
or U6360 (N_6360,N_6200,N_6217);
nor U6361 (N_6361,N_6283,N_6279);
or U6362 (N_6362,N_6243,N_6205);
or U6363 (N_6363,N_6210,N_6257);
and U6364 (N_6364,N_6210,N_6248);
nand U6365 (N_6365,N_6239,N_6291);
xor U6366 (N_6366,N_6267,N_6295);
nor U6367 (N_6367,N_6207,N_6270);
and U6368 (N_6368,N_6209,N_6268);
nand U6369 (N_6369,N_6250,N_6208);
nor U6370 (N_6370,N_6268,N_6293);
and U6371 (N_6371,N_6231,N_6225);
xor U6372 (N_6372,N_6288,N_6255);
or U6373 (N_6373,N_6290,N_6263);
or U6374 (N_6374,N_6292,N_6274);
nor U6375 (N_6375,N_6269,N_6245);
and U6376 (N_6376,N_6268,N_6246);
and U6377 (N_6377,N_6274,N_6229);
or U6378 (N_6378,N_6234,N_6281);
nand U6379 (N_6379,N_6283,N_6276);
and U6380 (N_6380,N_6292,N_6235);
or U6381 (N_6381,N_6280,N_6239);
or U6382 (N_6382,N_6249,N_6268);
nand U6383 (N_6383,N_6216,N_6282);
xnor U6384 (N_6384,N_6284,N_6222);
and U6385 (N_6385,N_6267,N_6293);
nor U6386 (N_6386,N_6250,N_6286);
or U6387 (N_6387,N_6252,N_6291);
and U6388 (N_6388,N_6201,N_6274);
nand U6389 (N_6389,N_6262,N_6212);
nor U6390 (N_6390,N_6239,N_6256);
xor U6391 (N_6391,N_6289,N_6213);
nor U6392 (N_6392,N_6271,N_6238);
nand U6393 (N_6393,N_6288,N_6223);
xor U6394 (N_6394,N_6220,N_6267);
and U6395 (N_6395,N_6280,N_6291);
and U6396 (N_6396,N_6283,N_6215);
xor U6397 (N_6397,N_6234,N_6227);
nor U6398 (N_6398,N_6226,N_6282);
or U6399 (N_6399,N_6206,N_6222);
nor U6400 (N_6400,N_6368,N_6387);
nor U6401 (N_6401,N_6351,N_6373);
nand U6402 (N_6402,N_6301,N_6356);
nand U6403 (N_6403,N_6398,N_6384);
and U6404 (N_6404,N_6348,N_6334);
and U6405 (N_6405,N_6338,N_6365);
or U6406 (N_6406,N_6374,N_6382);
xnor U6407 (N_6407,N_6347,N_6320);
and U6408 (N_6408,N_6300,N_6326);
or U6409 (N_6409,N_6325,N_6367);
and U6410 (N_6410,N_6360,N_6375);
nor U6411 (N_6411,N_6371,N_6319);
nor U6412 (N_6412,N_6395,N_6303);
or U6413 (N_6413,N_6317,N_6341);
nor U6414 (N_6414,N_6396,N_6315);
nor U6415 (N_6415,N_6345,N_6344);
nand U6416 (N_6416,N_6324,N_6391);
or U6417 (N_6417,N_6380,N_6363);
nor U6418 (N_6418,N_6333,N_6392);
and U6419 (N_6419,N_6305,N_6352);
nor U6420 (N_6420,N_6331,N_6349);
nand U6421 (N_6421,N_6307,N_6308);
or U6422 (N_6422,N_6362,N_6327);
nand U6423 (N_6423,N_6381,N_6383);
or U6424 (N_6424,N_6311,N_6309);
and U6425 (N_6425,N_6377,N_6323);
or U6426 (N_6426,N_6353,N_6337);
or U6427 (N_6427,N_6310,N_6394);
xor U6428 (N_6428,N_6390,N_6379);
nor U6429 (N_6429,N_6386,N_6372);
nor U6430 (N_6430,N_6350,N_6335);
nor U6431 (N_6431,N_6306,N_6366);
nand U6432 (N_6432,N_6312,N_6378);
xor U6433 (N_6433,N_6355,N_6321);
nand U6434 (N_6434,N_6358,N_6364);
xnor U6435 (N_6435,N_6314,N_6330);
or U6436 (N_6436,N_6343,N_6332);
nor U6437 (N_6437,N_6385,N_6361);
nand U6438 (N_6438,N_6316,N_6342);
and U6439 (N_6439,N_6389,N_6357);
and U6440 (N_6440,N_6318,N_6328);
nor U6441 (N_6441,N_6313,N_6322);
and U6442 (N_6442,N_6302,N_6354);
nor U6443 (N_6443,N_6397,N_6393);
xor U6444 (N_6444,N_6359,N_6340);
nand U6445 (N_6445,N_6388,N_6336);
nor U6446 (N_6446,N_6376,N_6369);
or U6447 (N_6447,N_6339,N_6370);
nand U6448 (N_6448,N_6399,N_6346);
or U6449 (N_6449,N_6304,N_6329);
or U6450 (N_6450,N_6395,N_6347);
or U6451 (N_6451,N_6314,N_6385);
nor U6452 (N_6452,N_6364,N_6346);
nor U6453 (N_6453,N_6372,N_6353);
nor U6454 (N_6454,N_6399,N_6312);
nor U6455 (N_6455,N_6369,N_6340);
and U6456 (N_6456,N_6350,N_6324);
and U6457 (N_6457,N_6312,N_6340);
xnor U6458 (N_6458,N_6338,N_6343);
and U6459 (N_6459,N_6365,N_6393);
or U6460 (N_6460,N_6363,N_6308);
nor U6461 (N_6461,N_6357,N_6330);
nor U6462 (N_6462,N_6371,N_6368);
nand U6463 (N_6463,N_6346,N_6353);
xor U6464 (N_6464,N_6363,N_6391);
xor U6465 (N_6465,N_6391,N_6384);
nand U6466 (N_6466,N_6365,N_6384);
nand U6467 (N_6467,N_6398,N_6333);
and U6468 (N_6468,N_6319,N_6358);
or U6469 (N_6469,N_6383,N_6386);
nor U6470 (N_6470,N_6309,N_6317);
nand U6471 (N_6471,N_6396,N_6369);
nor U6472 (N_6472,N_6357,N_6351);
and U6473 (N_6473,N_6329,N_6363);
and U6474 (N_6474,N_6325,N_6365);
nor U6475 (N_6475,N_6320,N_6394);
nor U6476 (N_6476,N_6347,N_6373);
or U6477 (N_6477,N_6340,N_6338);
and U6478 (N_6478,N_6318,N_6332);
and U6479 (N_6479,N_6366,N_6344);
nand U6480 (N_6480,N_6382,N_6356);
nor U6481 (N_6481,N_6376,N_6372);
and U6482 (N_6482,N_6309,N_6349);
or U6483 (N_6483,N_6324,N_6364);
or U6484 (N_6484,N_6309,N_6399);
xor U6485 (N_6485,N_6364,N_6383);
or U6486 (N_6486,N_6327,N_6304);
nor U6487 (N_6487,N_6305,N_6362);
nand U6488 (N_6488,N_6386,N_6333);
nor U6489 (N_6489,N_6304,N_6376);
nand U6490 (N_6490,N_6346,N_6308);
nor U6491 (N_6491,N_6314,N_6383);
xor U6492 (N_6492,N_6356,N_6384);
and U6493 (N_6493,N_6322,N_6346);
or U6494 (N_6494,N_6318,N_6317);
nand U6495 (N_6495,N_6388,N_6318);
nand U6496 (N_6496,N_6335,N_6334);
xnor U6497 (N_6497,N_6393,N_6387);
nor U6498 (N_6498,N_6340,N_6343);
or U6499 (N_6499,N_6348,N_6316);
nand U6500 (N_6500,N_6451,N_6468);
xnor U6501 (N_6501,N_6440,N_6484);
nor U6502 (N_6502,N_6473,N_6401);
and U6503 (N_6503,N_6433,N_6487);
nor U6504 (N_6504,N_6492,N_6431);
and U6505 (N_6505,N_6467,N_6491);
and U6506 (N_6506,N_6407,N_6488);
nand U6507 (N_6507,N_6432,N_6489);
or U6508 (N_6508,N_6434,N_6441);
nor U6509 (N_6509,N_6445,N_6465);
nand U6510 (N_6510,N_6459,N_6429);
or U6511 (N_6511,N_6411,N_6493);
nor U6512 (N_6512,N_6405,N_6454);
nand U6513 (N_6513,N_6442,N_6475);
nand U6514 (N_6514,N_6412,N_6406);
and U6515 (N_6515,N_6486,N_6477);
xnor U6516 (N_6516,N_6427,N_6483);
xor U6517 (N_6517,N_6472,N_6474);
nor U6518 (N_6518,N_6490,N_6455);
and U6519 (N_6519,N_6423,N_6419);
xor U6520 (N_6520,N_6485,N_6424);
nand U6521 (N_6521,N_6404,N_6400);
and U6522 (N_6522,N_6415,N_6437);
nand U6523 (N_6523,N_6476,N_6478);
xnor U6524 (N_6524,N_6402,N_6439);
and U6525 (N_6525,N_6458,N_6418);
xnor U6526 (N_6526,N_6425,N_6479);
xor U6527 (N_6527,N_6456,N_6460);
and U6528 (N_6528,N_6417,N_6403);
and U6529 (N_6529,N_6462,N_6422);
or U6530 (N_6530,N_6446,N_6471);
xor U6531 (N_6531,N_6482,N_6428);
or U6532 (N_6532,N_6470,N_6447);
and U6533 (N_6533,N_6448,N_6453);
nor U6534 (N_6534,N_6452,N_6466);
nand U6535 (N_6535,N_6481,N_6410);
nand U6536 (N_6536,N_6457,N_6464);
and U6537 (N_6537,N_6414,N_6495);
and U6538 (N_6538,N_6469,N_6444);
or U6539 (N_6539,N_6436,N_6430);
nor U6540 (N_6540,N_6450,N_6413);
nor U6541 (N_6541,N_6426,N_6480);
nor U6542 (N_6542,N_6420,N_6438);
nor U6543 (N_6543,N_6498,N_6499);
or U6544 (N_6544,N_6497,N_6463);
nand U6545 (N_6545,N_6494,N_6421);
nand U6546 (N_6546,N_6408,N_6416);
or U6547 (N_6547,N_6435,N_6496);
and U6548 (N_6548,N_6409,N_6449);
and U6549 (N_6549,N_6461,N_6443);
and U6550 (N_6550,N_6486,N_6460);
or U6551 (N_6551,N_6478,N_6441);
nor U6552 (N_6552,N_6440,N_6496);
or U6553 (N_6553,N_6494,N_6400);
or U6554 (N_6554,N_6482,N_6487);
or U6555 (N_6555,N_6442,N_6496);
nand U6556 (N_6556,N_6457,N_6417);
or U6557 (N_6557,N_6418,N_6470);
nor U6558 (N_6558,N_6434,N_6404);
and U6559 (N_6559,N_6478,N_6425);
xor U6560 (N_6560,N_6441,N_6460);
nand U6561 (N_6561,N_6411,N_6444);
xnor U6562 (N_6562,N_6452,N_6469);
and U6563 (N_6563,N_6434,N_6485);
or U6564 (N_6564,N_6425,N_6470);
nand U6565 (N_6565,N_6484,N_6498);
nor U6566 (N_6566,N_6494,N_6450);
nor U6567 (N_6567,N_6489,N_6463);
or U6568 (N_6568,N_6426,N_6465);
nand U6569 (N_6569,N_6465,N_6456);
or U6570 (N_6570,N_6482,N_6496);
nor U6571 (N_6571,N_6498,N_6410);
nor U6572 (N_6572,N_6420,N_6460);
nand U6573 (N_6573,N_6476,N_6464);
nor U6574 (N_6574,N_6401,N_6435);
nand U6575 (N_6575,N_6436,N_6426);
nor U6576 (N_6576,N_6459,N_6483);
and U6577 (N_6577,N_6444,N_6421);
or U6578 (N_6578,N_6466,N_6410);
and U6579 (N_6579,N_6495,N_6486);
and U6580 (N_6580,N_6405,N_6440);
and U6581 (N_6581,N_6400,N_6453);
or U6582 (N_6582,N_6449,N_6473);
nor U6583 (N_6583,N_6491,N_6438);
nand U6584 (N_6584,N_6458,N_6492);
or U6585 (N_6585,N_6476,N_6441);
or U6586 (N_6586,N_6494,N_6438);
nand U6587 (N_6587,N_6461,N_6499);
and U6588 (N_6588,N_6427,N_6464);
nand U6589 (N_6589,N_6445,N_6455);
or U6590 (N_6590,N_6457,N_6435);
nand U6591 (N_6591,N_6499,N_6400);
nand U6592 (N_6592,N_6438,N_6483);
nand U6593 (N_6593,N_6498,N_6414);
nor U6594 (N_6594,N_6484,N_6453);
nor U6595 (N_6595,N_6491,N_6487);
nand U6596 (N_6596,N_6439,N_6469);
or U6597 (N_6597,N_6446,N_6490);
nor U6598 (N_6598,N_6478,N_6455);
nand U6599 (N_6599,N_6492,N_6406);
or U6600 (N_6600,N_6594,N_6596);
or U6601 (N_6601,N_6535,N_6509);
or U6602 (N_6602,N_6554,N_6531);
nor U6603 (N_6603,N_6567,N_6542);
or U6604 (N_6604,N_6519,N_6558);
nand U6605 (N_6605,N_6577,N_6588);
nor U6606 (N_6606,N_6552,N_6510);
nand U6607 (N_6607,N_6502,N_6562);
or U6608 (N_6608,N_6533,N_6561);
xor U6609 (N_6609,N_6526,N_6565);
xnor U6610 (N_6610,N_6597,N_6575);
and U6611 (N_6611,N_6549,N_6546);
nand U6612 (N_6612,N_6574,N_6581);
or U6613 (N_6613,N_6569,N_6557);
or U6614 (N_6614,N_6541,N_6590);
nand U6615 (N_6615,N_6548,N_6578);
xor U6616 (N_6616,N_6570,N_6550);
nand U6617 (N_6617,N_6544,N_6523);
or U6618 (N_6618,N_6527,N_6504);
xor U6619 (N_6619,N_6508,N_6589);
nand U6620 (N_6620,N_6572,N_6586);
nor U6621 (N_6621,N_6566,N_6556);
and U6622 (N_6622,N_6571,N_6505);
nor U6623 (N_6623,N_6585,N_6584);
nor U6624 (N_6624,N_6559,N_6540);
and U6625 (N_6625,N_6551,N_6507);
nor U6626 (N_6626,N_6516,N_6555);
nor U6627 (N_6627,N_6532,N_6587);
and U6628 (N_6628,N_6529,N_6511);
nor U6629 (N_6629,N_6525,N_6560);
nand U6630 (N_6630,N_6543,N_6564);
nand U6631 (N_6631,N_6583,N_6545);
and U6632 (N_6632,N_6517,N_6518);
nand U6633 (N_6633,N_6563,N_6591);
and U6634 (N_6634,N_6528,N_6568);
nor U6635 (N_6635,N_6582,N_6599);
or U6636 (N_6636,N_6538,N_6547);
or U6637 (N_6637,N_6520,N_6513);
and U6638 (N_6638,N_6576,N_6592);
and U6639 (N_6639,N_6514,N_6500);
nor U6640 (N_6640,N_6595,N_6553);
or U6641 (N_6641,N_6580,N_6573);
nor U6642 (N_6642,N_6579,N_6522);
nor U6643 (N_6643,N_6593,N_6598);
and U6644 (N_6644,N_6536,N_6501);
and U6645 (N_6645,N_6503,N_6512);
nand U6646 (N_6646,N_6530,N_6515);
nand U6647 (N_6647,N_6537,N_6521);
or U6648 (N_6648,N_6534,N_6524);
and U6649 (N_6649,N_6539,N_6506);
and U6650 (N_6650,N_6549,N_6583);
or U6651 (N_6651,N_6562,N_6561);
and U6652 (N_6652,N_6507,N_6554);
or U6653 (N_6653,N_6562,N_6560);
xor U6654 (N_6654,N_6585,N_6567);
nand U6655 (N_6655,N_6581,N_6568);
nand U6656 (N_6656,N_6542,N_6582);
nor U6657 (N_6657,N_6525,N_6516);
or U6658 (N_6658,N_6522,N_6574);
nor U6659 (N_6659,N_6569,N_6538);
nand U6660 (N_6660,N_6586,N_6570);
nand U6661 (N_6661,N_6561,N_6567);
nor U6662 (N_6662,N_6500,N_6587);
nand U6663 (N_6663,N_6539,N_6571);
nand U6664 (N_6664,N_6501,N_6599);
and U6665 (N_6665,N_6511,N_6559);
or U6666 (N_6666,N_6524,N_6531);
and U6667 (N_6667,N_6530,N_6588);
nor U6668 (N_6668,N_6527,N_6503);
xnor U6669 (N_6669,N_6504,N_6574);
nor U6670 (N_6670,N_6528,N_6579);
or U6671 (N_6671,N_6567,N_6528);
nor U6672 (N_6672,N_6573,N_6561);
nor U6673 (N_6673,N_6540,N_6554);
or U6674 (N_6674,N_6529,N_6540);
nand U6675 (N_6675,N_6537,N_6592);
nor U6676 (N_6676,N_6597,N_6508);
nand U6677 (N_6677,N_6551,N_6540);
or U6678 (N_6678,N_6508,N_6599);
nor U6679 (N_6679,N_6510,N_6597);
nand U6680 (N_6680,N_6506,N_6528);
or U6681 (N_6681,N_6572,N_6522);
or U6682 (N_6682,N_6584,N_6572);
nor U6683 (N_6683,N_6524,N_6580);
nand U6684 (N_6684,N_6519,N_6537);
nand U6685 (N_6685,N_6580,N_6596);
nand U6686 (N_6686,N_6501,N_6557);
nor U6687 (N_6687,N_6524,N_6558);
nand U6688 (N_6688,N_6571,N_6568);
and U6689 (N_6689,N_6592,N_6538);
nor U6690 (N_6690,N_6537,N_6570);
or U6691 (N_6691,N_6509,N_6507);
or U6692 (N_6692,N_6594,N_6571);
nor U6693 (N_6693,N_6562,N_6518);
nand U6694 (N_6694,N_6531,N_6582);
nor U6695 (N_6695,N_6580,N_6522);
and U6696 (N_6696,N_6568,N_6541);
and U6697 (N_6697,N_6504,N_6557);
or U6698 (N_6698,N_6539,N_6563);
or U6699 (N_6699,N_6564,N_6595);
or U6700 (N_6700,N_6601,N_6676);
and U6701 (N_6701,N_6684,N_6696);
nor U6702 (N_6702,N_6609,N_6620);
nand U6703 (N_6703,N_6673,N_6607);
and U6704 (N_6704,N_6685,N_6675);
and U6705 (N_6705,N_6648,N_6625);
and U6706 (N_6706,N_6666,N_6699);
nand U6707 (N_6707,N_6682,N_6650);
and U6708 (N_6708,N_6612,N_6653);
nand U6709 (N_6709,N_6678,N_6626);
or U6710 (N_6710,N_6674,N_6665);
nand U6711 (N_6711,N_6640,N_6667);
and U6712 (N_6712,N_6634,N_6656);
or U6713 (N_6713,N_6631,N_6693);
and U6714 (N_6714,N_6659,N_6668);
and U6715 (N_6715,N_6679,N_6641);
or U6716 (N_6716,N_6604,N_6611);
nand U6717 (N_6717,N_6617,N_6613);
nor U6718 (N_6718,N_6654,N_6651);
nand U6719 (N_6719,N_6647,N_6600);
and U6720 (N_6720,N_6662,N_6681);
and U6721 (N_6721,N_6677,N_6695);
and U6722 (N_6722,N_6687,N_6622);
nand U6723 (N_6723,N_6646,N_6670);
nand U6724 (N_6724,N_6649,N_6642);
and U6725 (N_6725,N_6697,N_6618);
nor U6726 (N_6726,N_6637,N_6616);
or U6727 (N_6727,N_6610,N_6664);
nand U6728 (N_6728,N_6680,N_6606);
or U6729 (N_6729,N_6658,N_6657);
or U6730 (N_6730,N_6619,N_6688);
xnor U6731 (N_6731,N_6615,N_6660);
nor U6732 (N_6732,N_6692,N_6672);
nor U6733 (N_6733,N_6603,N_6661);
nand U6734 (N_6734,N_6624,N_6623);
nand U6735 (N_6735,N_6671,N_6636);
nor U6736 (N_6736,N_6663,N_6605);
nor U6737 (N_6737,N_6608,N_6645);
nand U6738 (N_6738,N_6669,N_6627);
nand U6739 (N_6739,N_6633,N_6630);
and U6740 (N_6740,N_6629,N_6694);
and U6741 (N_6741,N_6632,N_6683);
and U6742 (N_6742,N_6655,N_6652);
or U6743 (N_6743,N_6639,N_6638);
or U6744 (N_6744,N_6628,N_6644);
nand U6745 (N_6745,N_6621,N_6614);
nand U6746 (N_6746,N_6691,N_6689);
nor U6747 (N_6747,N_6635,N_6690);
nor U6748 (N_6748,N_6686,N_6602);
or U6749 (N_6749,N_6643,N_6698);
nor U6750 (N_6750,N_6604,N_6640);
and U6751 (N_6751,N_6628,N_6600);
nor U6752 (N_6752,N_6663,N_6611);
or U6753 (N_6753,N_6638,N_6667);
xnor U6754 (N_6754,N_6684,N_6687);
nand U6755 (N_6755,N_6650,N_6634);
nand U6756 (N_6756,N_6675,N_6689);
and U6757 (N_6757,N_6603,N_6645);
nand U6758 (N_6758,N_6668,N_6631);
nand U6759 (N_6759,N_6674,N_6692);
nor U6760 (N_6760,N_6675,N_6668);
and U6761 (N_6761,N_6642,N_6632);
and U6762 (N_6762,N_6633,N_6607);
nand U6763 (N_6763,N_6643,N_6657);
or U6764 (N_6764,N_6636,N_6687);
xnor U6765 (N_6765,N_6677,N_6658);
xor U6766 (N_6766,N_6630,N_6657);
nor U6767 (N_6767,N_6600,N_6694);
or U6768 (N_6768,N_6628,N_6656);
and U6769 (N_6769,N_6630,N_6648);
nand U6770 (N_6770,N_6642,N_6689);
nor U6771 (N_6771,N_6621,N_6623);
and U6772 (N_6772,N_6636,N_6600);
and U6773 (N_6773,N_6664,N_6611);
nand U6774 (N_6774,N_6667,N_6669);
or U6775 (N_6775,N_6623,N_6603);
nand U6776 (N_6776,N_6664,N_6651);
nor U6777 (N_6777,N_6616,N_6663);
nor U6778 (N_6778,N_6655,N_6605);
or U6779 (N_6779,N_6654,N_6645);
or U6780 (N_6780,N_6623,N_6629);
nor U6781 (N_6781,N_6687,N_6631);
xnor U6782 (N_6782,N_6645,N_6613);
and U6783 (N_6783,N_6663,N_6627);
nor U6784 (N_6784,N_6631,N_6637);
nand U6785 (N_6785,N_6667,N_6652);
or U6786 (N_6786,N_6616,N_6666);
nand U6787 (N_6787,N_6673,N_6682);
and U6788 (N_6788,N_6604,N_6610);
nor U6789 (N_6789,N_6606,N_6689);
xor U6790 (N_6790,N_6638,N_6656);
and U6791 (N_6791,N_6645,N_6667);
nand U6792 (N_6792,N_6615,N_6604);
or U6793 (N_6793,N_6602,N_6619);
nor U6794 (N_6794,N_6676,N_6625);
and U6795 (N_6795,N_6625,N_6634);
nor U6796 (N_6796,N_6608,N_6626);
nor U6797 (N_6797,N_6698,N_6603);
or U6798 (N_6798,N_6612,N_6605);
or U6799 (N_6799,N_6664,N_6646);
nor U6800 (N_6800,N_6704,N_6716);
nor U6801 (N_6801,N_6703,N_6735);
or U6802 (N_6802,N_6762,N_6709);
and U6803 (N_6803,N_6784,N_6740);
nand U6804 (N_6804,N_6751,N_6700);
and U6805 (N_6805,N_6705,N_6742);
nand U6806 (N_6806,N_6774,N_6790);
or U6807 (N_6807,N_6749,N_6739);
and U6808 (N_6808,N_6721,N_6778);
or U6809 (N_6809,N_6767,N_6781);
or U6810 (N_6810,N_6711,N_6769);
or U6811 (N_6811,N_6741,N_6791);
and U6812 (N_6812,N_6702,N_6776);
nand U6813 (N_6813,N_6792,N_6730);
nor U6814 (N_6814,N_6787,N_6731);
nand U6815 (N_6815,N_6725,N_6763);
and U6816 (N_6816,N_6772,N_6723);
nor U6817 (N_6817,N_6732,N_6783);
nand U6818 (N_6818,N_6759,N_6768);
nand U6819 (N_6819,N_6770,N_6715);
and U6820 (N_6820,N_6718,N_6757);
nor U6821 (N_6821,N_6746,N_6799);
nand U6822 (N_6822,N_6708,N_6727);
and U6823 (N_6823,N_6728,N_6745);
xor U6824 (N_6824,N_6760,N_6707);
nand U6825 (N_6825,N_6722,N_6737);
and U6826 (N_6826,N_6710,N_6750);
nand U6827 (N_6827,N_6797,N_6753);
and U6828 (N_6828,N_6766,N_6782);
or U6829 (N_6829,N_6761,N_6758);
and U6830 (N_6830,N_6795,N_6771);
nand U6831 (N_6831,N_6748,N_6777);
and U6832 (N_6832,N_6743,N_6733);
or U6833 (N_6833,N_6714,N_6764);
or U6834 (N_6834,N_6765,N_6747);
xnor U6835 (N_6835,N_6793,N_6779);
nand U6836 (N_6836,N_6726,N_6736);
nand U6837 (N_6837,N_6796,N_6701);
nand U6838 (N_6838,N_6755,N_6754);
nand U6839 (N_6839,N_6752,N_6734);
nor U6840 (N_6840,N_6744,N_6786);
nor U6841 (N_6841,N_6738,N_6788);
and U6842 (N_6842,N_6720,N_6712);
nor U6843 (N_6843,N_6794,N_6785);
or U6844 (N_6844,N_6706,N_6789);
or U6845 (N_6845,N_6713,N_6775);
nand U6846 (N_6846,N_6756,N_6717);
or U6847 (N_6847,N_6719,N_6773);
or U6848 (N_6848,N_6798,N_6729);
nor U6849 (N_6849,N_6724,N_6780);
nor U6850 (N_6850,N_6798,N_6748);
and U6851 (N_6851,N_6715,N_6765);
nand U6852 (N_6852,N_6776,N_6758);
nand U6853 (N_6853,N_6758,N_6717);
nor U6854 (N_6854,N_6729,N_6718);
nand U6855 (N_6855,N_6764,N_6751);
nor U6856 (N_6856,N_6758,N_6714);
and U6857 (N_6857,N_6787,N_6770);
nor U6858 (N_6858,N_6779,N_6700);
and U6859 (N_6859,N_6701,N_6745);
and U6860 (N_6860,N_6757,N_6700);
or U6861 (N_6861,N_6705,N_6779);
or U6862 (N_6862,N_6717,N_6749);
nor U6863 (N_6863,N_6785,N_6773);
or U6864 (N_6864,N_6788,N_6772);
nand U6865 (N_6865,N_6760,N_6799);
or U6866 (N_6866,N_6763,N_6709);
or U6867 (N_6867,N_6708,N_6760);
or U6868 (N_6868,N_6743,N_6748);
and U6869 (N_6869,N_6764,N_6740);
and U6870 (N_6870,N_6743,N_6789);
nand U6871 (N_6871,N_6723,N_6749);
nor U6872 (N_6872,N_6791,N_6780);
and U6873 (N_6873,N_6774,N_6735);
or U6874 (N_6874,N_6754,N_6785);
nor U6875 (N_6875,N_6742,N_6700);
xnor U6876 (N_6876,N_6767,N_6753);
nor U6877 (N_6877,N_6744,N_6799);
nor U6878 (N_6878,N_6737,N_6713);
nor U6879 (N_6879,N_6787,N_6794);
nor U6880 (N_6880,N_6782,N_6775);
nand U6881 (N_6881,N_6786,N_6727);
nand U6882 (N_6882,N_6700,N_6738);
nand U6883 (N_6883,N_6735,N_6795);
nand U6884 (N_6884,N_6791,N_6700);
xnor U6885 (N_6885,N_6751,N_6727);
nor U6886 (N_6886,N_6796,N_6711);
nor U6887 (N_6887,N_6794,N_6710);
nor U6888 (N_6888,N_6772,N_6774);
and U6889 (N_6889,N_6761,N_6714);
nor U6890 (N_6890,N_6762,N_6798);
xor U6891 (N_6891,N_6767,N_6730);
nand U6892 (N_6892,N_6779,N_6710);
and U6893 (N_6893,N_6731,N_6754);
or U6894 (N_6894,N_6726,N_6785);
nand U6895 (N_6895,N_6743,N_6700);
and U6896 (N_6896,N_6782,N_6701);
and U6897 (N_6897,N_6704,N_6792);
nor U6898 (N_6898,N_6702,N_6772);
xor U6899 (N_6899,N_6709,N_6798);
xor U6900 (N_6900,N_6812,N_6809);
and U6901 (N_6901,N_6843,N_6864);
nor U6902 (N_6902,N_6879,N_6854);
nand U6903 (N_6903,N_6826,N_6827);
nand U6904 (N_6904,N_6883,N_6841);
and U6905 (N_6905,N_6867,N_6859);
and U6906 (N_6906,N_6886,N_6866);
nand U6907 (N_6907,N_6865,N_6823);
nor U6908 (N_6908,N_6821,N_6846);
nor U6909 (N_6909,N_6804,N_6882);
xnor U6910 (N_6910,N_6825,N_6892);
nand U6911 (N_6911,N_6813,N_6822);
nand U6912 (N_6912,N_6818,N_6811);
nand U6913 (N_6913,N_6840,N_6885);
or U6914 (N_6914,N_6808,N_6848);
nor U6915 (N_6915,N_6838,N_6837);
nor U6916 (N_6916,N_6836,N_6876);
or U6917 (N_6917,N_6881,N_6862);
nand U6918 (N_6918,N_6860,N_6807);
or U6919 (N_6919,N_6891,N_6829);
and U6920 (N_6920,N_6894,N_6802);
and U6921 (N_6921,N_6828,N_6889);
nand U6922 (N_6922,N_6897,N_6877);
nand U6923 (N_6923,N_6888,N_6814);
nand U6924 (N_6924,N_6805,N_6853);
nand U6925 (N_6925,N_6815,N_6839);
xnor U6926 (N_6926,N_6852,N_6842);
nor U6927 (N_6927,N_6816,N_6884);
nand U6928 (N_6928,N_6851,N_6820);
and U6929 (N_6929,N_6834,N_6874);
or U6930 (N_6930,N_6806,N_6855);
nand U6931 (N_6931,N_6810,N_6847);
xor U6932 (N_6932,N_6872,N_6857);
and U6933 (N_6933,N_6870,N_6833);
xor U6934 (N_6934,N_6896,N_6869);
nor U6935 (N_6935,N_6845,N_6875);
nand U6936 (N_6936,N_6873,N_6868);
xor U6937 (N_6937,N_6858,N_6850);
nand U6938 (N_6938,N_6880,N_6844);
or U6939 (N_6939,N_6893,N_6878);
nand U6940 (N_6940,N_6856,N_6832);
nor U6941 (N_6941,N_6887,N_6899);
and U6942 (N_6942,N_6861,N_6824);
nand U6943 (N_6943,N_6817,N_6830);
nor U6944 (N_6944,N_6898,N_6871);
nor U6945 (N_6945,N_6895,N_6800);
nand U6946 (N_6946,N_6863,N_6819);
nand U6947 (N_6947,N_6831,N_6801);
xnor U6948 (N_6948,N_6890,N_6849);
xor U6949 (N_6949,N_6835,N_6803);
nand U6950 (N_6950,N_6826,N_6807);
nor U6951 (N_6951,N_6829,N_6851);
nand U6952 (N_6952,N_6843,N_6873);
nand U6953 (N_6953,N_6864,N_6816);
or U6954 (N_6954,N_6834,N_6870);
or U6955 (N_6955,N_6829,N_6821);
nand U6956 (N_6956,N_6873,N_6871);
and U6957 (N_6957,N_6826,N_6896);
nor U6958 (N_6958,N_6890,N_6888);
xnor U6959 (N_6959,N_6872,N_6807);
xor U6960 (N_6960,N_6869,N_6879);
and U6961 (N_6961,N_6809,N_6858);
and U6962 (N_6962,N_6851,N_6874);
or U6963 (N_6963,N_6852,N_6885);
nand U6964 (N_6964,N_6860,N_6819);
or U6965 (N_6965,N_6889,N_6899);
nand U6966 (N_6966,N_6856,N_6869);
or U6967 (N_6967,N_6808,N_6836);
and U6968 (N_6968,N_6892,N_6817);
xnor U6969 (N_6969,N_6848,N_6836);
and U6970 (N_6970,N_6847,N_6879);
nor U6971 (N_6971,N_6826,N_6888);
and U6972 (N_6972,N_6874,N_6815);
and U6973 (N_6973,N_6890,N_6837);
nand U6974 (N_6974,N_6878,N_6865);
nand U6975 (N_6975,N_6898,N_6861);
nor U6976 (N_6976,N_6818,N_6844);
and U6977 (N_6977,N_6878,N_6839);
nand U6978 (N_6978,N_6806,N_6876);
and U6979 (N_6979,N_6894,N_6812);
nand U6980 (N_6980,N_6881,N_6827);
and U6981 (N_6981,N_6858,N_6836);
xnor U6982 (N_6982,N_6854,N_6866);
and U6983 (N_6983,N_6843,N_6889);
or U6984 (N_6984,N_6851,N_6831);
and U6985 (N_6985,N_6861,N_6846);
and U6986 (N_6986,N_6856,N_6824);
and U6987 (N_6987,N_6808,N_6866);
xor U6988 (N_6988,N_6820,N_6818);
nor U6989 (N_6989,N_6886,N_6815);
nor U6990 (N_6990,N_6839,N_6887);
or U6991 (N_6991,N_6856,N_6884);
nand U6992 (N_6992,N_6848,N_6822);
nand U6993 (N_6993,N_6867,N_6898);
or U6994 (N_6994,N_6892,N_6844);
nor U6995 (N_6995,N_6871,N_6860);
nand U6996 (N_6996,N_6848,N_6865);
xor U6997 (N_6997,N_6865,N_6838);
and U6998 (N_6998,N_6825,N_6852);
nand U6999 (N_6999,N_6813,N_6829);
xor U7000 (N_7000,N_6944,N_6928);
nor U7001 (N_7001,N_6988,N_6934);
and U7002 (N_7002,N_6943,N_6941);
nor U7003 (N_7003,N_6964,N_6965);
and U7004 (N_7004,N_6926,N_6915);
xor U7005 (N_7005,N_6962,N_6942);
nor U7006 (N_7006,N_6956,N_6925);
and U7007 (N_7007,N_6980,N_6911);
and U7008 (N_7008,N_6952,N_6985);
xnor U7009 (N_7009,N_6916,N_6951);
nand U7010 (N_7010,N_6927,N_6969);
nand U7011 (N_7011,N_6905,N_6932);
and U7012 (N_7012,N_6975,N_6963);
nand U7013 (N_7013,N_6960,N_6938);
and U7014 (N_7014,N_6961,N_6993);
xor U7015 (N_7015,N_6953,N_6968);
nand U7016 (N_7016,N_6977,N_6999);
nor U7017 (N_7017,N_6936,N_6971);
xnor U7018 (N_7018,N_6990,N_6918);
nor U7019 (N_7019,N_6973,N_6970);
and U7020 (N_7020,N_6907,N_6998);
and U7021 (N_7021,N_6919,N_6981);
nor U7022 (N_7022,N_6913,N_6921);
and U7023 (N_7023,N_6939,N_6955);
nand U7024 (N_7024,N_6974,N_6914);
or U7025 (N_7025,N_6930,N_6959);
nand U7026 (N_7026,N_6997,N_6978);
and U7027 (N_7027,N_6992,N_6991);
or U7028 (N_7028,N_6994,N_6924);
nor U7029 (N_7029,N_6979,N_6940);
nor U7030 (N_7030,N_6917,N_6945);
nor U7031 (N_7031,N_6984,N_6937);
nand U7032 (N_7032,N_6947,N_6904);
nor U7033 (N_7033,N_6972,N_6908);
nand U7034 (N_7034,N_6967,N_6900);
xnor U7035 (N_7035,N_6986,N_6949);
or U7036 (N_7036,N_6912,N_6950);
or U7037 (N_7037,N_6920,N_6989);
nor U7038 (N_7038,N_6954,N_6966);
xnor U7039 (N_7039,N_6983,N_6929);
xor U7040 (N_7040,N_6996,N_6948);
nor U7041 (N_7041,N_6906,N_6931);
and U7042 (N_7042,N_6946,N_6910);
nor U7043 (N_7043,N_6901,N_6982);
and U7044 (N_7044,N_6903,N_6923);
and U7045 (N_7045,N_6935,N_6933);
nand U7046 (N_7046,N_6957,N_6909);
or U7047 (N_7047,N_6987,N_6902);
xnor U7048 (N_7048,N_6922,N_6995);
nand U7049 (N_7049,N_6958,N_6976);
nand U7050 (N_7050,N_6963,N_6950);
and U7051 (N_7051,N_6987,N_6924);
xor U7052 (N_7052,N_6988,N_6994);
and U7053 (N_7053,N_6965,N_6950);
or U7054 (N_7054,N_6913,N_6982);
nand U7055 (N_7055,N_6910,N_6936);
nand U7056 (N_7056,N_6911,N_6903);
nand U7057 (N_7057,N_6911,N_6917);
nor U7058 (N_7058,N_6954,N_6926);
or U7059 (N_7059,N_6989,N_6945);
nand U7060 (N_7060,N_6910,N_6956);
and U7061 (N_7061,N_6994,N_6928);
xor U7062 (N_7062,N_6918,N_6910);
or U7063 (N_7063,N_6954,N_6992);
nand U7064 (N_7064,N_6938,N_6980);
nor U7065 (N_7065,N_6934,N_6987);
or U7066 (N_7066,N_6948,N_6960);
nand U7067 (N_7067,N_6966,N_6995);
and U7068 (N_7068,N_6926,N_6922);
nand U7069 (N_7069,N_6906,N_6979);
xor U7070 (N_7070,N_6941,N_6953);
and U7071 (N_7071,N_6907,N_6984);
nor U7072 (N_7072,N_6995,N_6986);
nor U7073 (N_7073,N_6917,N_6916);
nor U7074 (N_7074,N_6946,N_6906);
or U7075 (N_7075,N_6997,N_6974);
nand U7076 (N_7076,N_6914,N_6948);
nand U7077 (N_7077,N_6995,N_6921);
or U7078 (N_7078,N_6993,N_6912);
or U7079 (N_7079,N_6919,N_6946);
and U7080 (N_7080,N_6952,N_6965);
or U7081 (N_7081,N_6902,N_6969);
nand U7082 (N_7082,N_6946,N_6968);
nor U7083 (N_7083,N_6999,N_6921);
or U7084 (N_7084,N_6999,N_6987);
nand U7085 (N_7085,N_6999,N_6971);
nor U7086 (N_7086,N_6916,N_6952);
or U7087 (N_7087,N_6900,N_6942);
or U7088 (N_7088,N_6923,N_6906);
nor U7089 (N_7089,N_6904,N_6979);
or U7090 (N_7090,N_6913,N_6974);
or U7091 (N_7091,N_6968,N_6983);
and U7092 (N_7092,N_6952,N_6987);
nand U7093 (N_7093,N_6974,N_6980);
xor U7094 (N_7094,N_6904,N_6921);
nor U7095 (N_7095,N_6951,N_6952);
nand U7096 (N_7096,N_6950,N_6910);
or U7097 (N_7097,N_6918,N_6911);
or U7098 (N_7098,N_6947,N_6934);
or U7099 (N_7099,N_6961,N_6925);
or U7100 (N_7100,N_7068,N_7088);
nand U7101 (N_7101,N_7075,N_7096);
nand U7102 (N_7102,N_7072,N_7024);
and U7103 (N_7103,N_7042,N_7039);
or U7104 (N_7104,N_7025,N_7090);
and U7105 (N_7105,N_7078,N_7029);
or U7106 (N_7106,N_7002,N_7070);
nor U7107 (N_7107,N_7067,N_7058);
and U7108 (N_7108,N_7097,N_7069);
nor U7109 (N_7109,N_7092,N_7099);
and U7110 (N_7110,N_7044,N_7041);
or U7111 (N_7111,N_7031,N_7045);
nand U7112 (N_7112,N_7089,N_7001);
nand U7113 (N_7113,N_7063,N_7038);
nand U7114 (N_7114,N_7053,N_7060);
nand U7115 (N_7115,N_7030,N_7013);
xor U7116 (N_7116,N_7021,N_7037);
xnor U7117 (N_7117,N_7065,N_7057);
and U7118 (N_7118,N_7005,N_7085);
or U7119 (N_7119,N_7054,N_7056);
xnor U7120 (N_7120,N_7074,N_7084);
or U7121 (N_7121,N_7083,N_7043);
nand U7122 (N_7122,N_7079,N_7094);
xor U7123 (N_7123,N_7007,N_7027);
nor U7124 (N_7124,N_7009,N_7049);
nor U7125 (N_7125,N_7026,N_7014);
xnor U7126 (N_7126,N_7040,N_7073);
nand U7127 (N_7127,N_7003,N_7036);
nor U7128 (N_7128,N_7066,N_7091);
xor U7129 (N_7129,N_7046,N_7076);
nor U7130 (N_7130,N_7004,N_7052);
and U7131 (N_7131,N_7047,N_7062);
nand U7132 (N_7132,N_7087,N_7051);
and U7133 (N_7133,N_7019,N_7082);
nor U7134 (N_7134,N_7035,N_7080);
nand U7135 (N_7135,N_7020,N_7008);
nand U7136 (N_7136,N_7016,N_7050);
xor U7137 (N_7137,N_7086,N_7010);
nor U7138 (N_7138,N_7028,N_7022);
and U7139 (N_7139,N_7055,N_7006);
nor U7140 (N_7140,N_7033,N_7093);
nand U7141 (N_7141,N_7011,N_7000);
nand U7142 (N_7142,N_7064,N_7077);
nand U7143 (N_7143,N_7018,N_7098);
nor U7144 (N_7144,N_7071,N_7048);
and U7145 (N_7145,N_7017,N_7061);
nor U7146 (N_7146,N_7095,N_7034);
or U7147 (N_7147,N_7023,N_7081);
nor U7148 (N_7148,N_7032,N_7015);
nor U7149 (N_7149,N_7059,N_7012);
nand U7150 (N_7150,N_7089,N_7087);
and U7151 (N_7151,N_7021,N_7051);
nor U7152 (N_7152,N_7036,N_7039);
and U7153 (N_7153,N_7041,N_7080);
nand U7154 (N_7154,N_7028,N_7085);
nor U7155 (N_7155,N_7061,N_7035);
or U7156 (N_7156,N_7063,N_7045);
or U7157 (N_7157,N_7074,N_7010);
nand U7158 (N_7158,N_7071,N_7095);
nor U7159 (N_7159,N_7042,N_7050);
xnor U7160 (N_7160,N_7049,N_7099);
nand U7161 (N_7161,N_7074,N_7012);
or U7162 (N_7162,N_7036,N_7069);
and U7163 (N_7163,N_7065,N_7090);
nor U7164 (N_7164,N_7049,N_7067);
and U7165 (N_7165,N_7017,N_7089);
and U7166 (N_7166,N_7076,N_7098);
or U7167 (N_7167,N_7027,N_7030);
xor U7168 (N_7168,N_7079,N_7040);
or U7169 (N_7169,N_7064,N_7038);
nand U7170 (N_7170,N_7010,N_7081);
and U7171 (N_7171,N_7030,N_7063);
or U7172 (N_7172,N_7064,N_7091);
nor U7173 (N_7173,N_7083,N_7015);
nand U7174 (N_7174,N_7074,N_7054);
or U7175 (N_7175,N_7033,N_7068);
and U7176 (N_7176,N_7007,N_7046);
or U7177 (N_7177,N_7077,N_7016);
nand U7178 (N_7178,N_7072,N_7003);
nor U7179 (N_7179,N_7006,N_7031);
nand U7180 (N_7180,N_7022,N_7020);
nand U7181 (N_7181,N_7016,N_7090);
xor U7182 (N_7182,N_7097,N_7052);
nor U7183 (N_7183,N_7033,N_7049);
nor U7184 (N_7184,N_7006,N_7094);
nor U7185 (N_7185,N_7084,N_7064);
xnor U7186 (N_7186,N_7091,N_7032);
nor U7187 (N_7187,N_7033,N_7014);
nand U7188 (N_7188,N_7011,N_7040);
xnor U7189 (N_7189,N_7010,N_7007);
and U7190 (N_7190,N_7009,N_7018);
and U7191 (N_7191,N_7037,N_7016);
and U7192 (N_7192,N_7033,N_7036);
nand U7193 (N_7193,N_7057,N_7008);
and U7194 (N_7194,N_7098,N_7023);
nand U7195 (N_7195,N_7001,N_7045);
nor U7196 (N_7196,N_7097,N_7037);
and U7197 (N_7197,N_7010,N_7055);
and U7198 (N_7198,N_7018,N_7097);
and U7199 (N_7199,N_7062,N_7034);
or U7200 (N_7200,N_7197,N_7158);
nand U7201 (N_7201,N_7122,N_7142);
and U7202 (N_7202,N_7192,N_7171);
and U7203 (N_7203,N_7139,N_7130);
nand U7204 (N_7204,N_7180,N_7153);
and U7205 (N_7205,N_7103,N_7133);
and U7206 (N_7206,N_7157,N_7131);
and U7207 (N_7207,N_7116,N_7175);
or U7208 (N_7208,N_7163,N_7169);
nor U7209 (N_7209,N_7114,N_7143);
nand U7210 (N_7210,N_7132,N_7117);
or U7211 (N_7211,N_7199,N_7161);
and U7212 (N_7212,N_7172,N_7145);
nor U7213 (N_7213,N_7155,N_7140);
or U7214 (N_7214,N_7174,N_7127);
nand U7215 (N_7215,N_7107,N_7150);
nor U7216 (N_7216,N_7193,N_7147);
nand U7217 (N_7217,N_7151,N_7101);
nand U7218 (N_7218,N_7144,N_7166);
nand U7219 (N_7219,N_7181,N_7198);
nor U7220 (N_7220,N_7136,N_7164);
nand U7221 (N_7221,N_7120,N_7141);
nand U7222 (N_7222,N_7191,N_7173);
xnor U7223 (N_7223,N_7188,N_7146);
nor U7224 (N_7224,N_7184,N_7168);
or U7225 (N_7225,N_7121,N_7100);
nor U7226 (N_7226,N_7167,N_7135);
and U7227 (N_7227,N_7152,N_7119);
or U7228 (N_7228,N_7104,N_7126);
or U7229 (N_7229,N_7115,N_7148);
or U7230 (N_7230,N_7176,N_7178);
xnor U7231 (N_7231,N_7128,N_7125);
or U7232 (N_7232,N_7190,N_7154);
nand U7233 (N_7233,N_7156,N_7129);
xnor U7234 (N_7234,N_7102,N_7165);
nand U7235 (N_7235,N_7113,N_7179);
nor U7236 (N_7236,N_7124,N_7106);
nand U7237 (N_7237,N_7137,N_7118);
and U7238 (N_7238,N_7112,N_7177);
or U7239 (N_7239,N_7111,N_7182);
xor U7240 (N_7240,N_7134,N_7195);
xor U7241 (N_7241,N_7109,N_7162);
nand U7242 (N_7242,N_7149,N_7196);
nor U7243 (N_7243,N_7138,N_7159);
nand U7244 (N_7244,N_7189,N_7185);
nor U7245 (N_7245,N_7160,N_7186);
and U7246 (N_7246,N_7105,N_7187);
and U7247 (N_7247,N_7183,N_7108);
nand U7248 (N_7248,N_7110,N_7123);
nor U7249 (N_7249,N_7194,N_7170);
xnor U7250 (N_7250,N_7163,N_7103);
or U7251 (N_7251,N_7105,N_7179);
nor U7252 (N_7252,N_7164,N_7133);
xor U7253 (N_7253,N_7182,N_7127);
or U7254 (N_7254,N_7122,N_7194);
or U7255 (N_7255,N_7159,N_7105);
and U7256 (N_7256,N_7141,N_7177);
nand U7257 (N_7257,N_7135,N_7132);
xor U7258 (N_7258,N_7178,N_7107);
nand U7259 (N_7259,N_7120,N_7197);
and U7260 (N_7260,N_7151,N_7110);
or U7261 (N_7261,N_7199,N_7176);
and U7262 (N_7262,N_7164,N_7191);
nor U7263 (N_7263,N_7160,N_7122);
xnor U7264 (N_7264,N_7139,N_7141);
or U7265 (N_7265,N_7155,N_7146);
and U7266 (N_7266,N_7136,N_7112);
nor U7267 (N_7267,N_7167,N_7119);
nor U7268 (N_7268,N_7155,N_7118);
nand U7269 (N_7269,N_7109,N_7197);
nor U7270 (N_7270,N_7144,N_7101);
or U7271 (N_7271,N_7148,N_7120);
or U7272 (N_7272,N_7113,N_7123);
xnor U7273 (N_7273,N_7167,N_7185);
or U7274 (N_7274,N_7181,N_7147);
or U7275 (N_7275,N_7177,N_7106);
nand U7276 (N_7276,N_7117,N_7108);
nand U7277 (N_7277,N_7134,N_7158);
nand U7278 (N_7278,N_7137,N_7182);
nand U7279 (N_7279,N_7109,N_7102);
nor U7280 (N_7280,N_7111,N_7132);
nand U7281 (N_7281,N_7174,N_7175);
nand U7282 (N_7282,N_7197,N_7198);
or U7283 (N_7283,N_7193,N_7156);
nand U7284 (N_7284,N_7100,N_7159);
nor U7285 (N_7285,N_7186,N_7118);
or U7286 (N_7286,N_7197,N_7106);
nor U7287 (N_7287,N_7112,N_7197);
xnor U7288 (N_7288,N_7159,N_7175);
nor U7289 (N_7289,N_7105,N_7101);
nor U7290 (N_7290,N_7123,N_7193);
nand U7291 (N_7291,N_7129,N_7120);
nand U7292 (N_7292,N_7157,N_7133);
nor U7293 (N_7293,N_7135,N_7160);
nand U7294 (N_7294,N_7107,N_7180);
or U7295 (N_7295,N_7187,N_7109);
and U7296 (N_7296,N_7123,N_7150);
and U7297 (N_7297,N_7107,N_7147);
nand U7298 (N_7298,N_7154,N_7105);
xor U7299 (N_7299,N_7166,N_7113);
nor U7300 (N_7300,N_7216,N_7249);
xor U7301 (N_7301,N_7287,N_7232);
or U7302 (N_7302,N_7271,N_7227);
nor U7303 (N_7303,N_7291,N_7261);
nor U7304 (N_7304,N_7234,N_7274);
and U7305 (N_7305,N_7236,N_7209);
nand U7306 (N_7306,N_7282,N_7260);
nor U7307 (N_7307,N_7241,N_7247);
or U7308 (N_7308,N_7206,N_7252);
nand U7309 (N_7309,N_7270,N_7267);
nor U7310 (N_7310,N_7245,N_7259);
or U7311 (N_7311,N_7200,N_7279);
or U7312 (N_7312,N_7207,N_7263);
nand U7313 (N_7313,N_7254,N_7215);
or U7314 (N_7314,N_7225,N_7242);
nand U7315 (N_7315,N_7257,N_7201);
or U7316 (N_7316,N_7204,N_7275);
nand U7317 (N_7317,N_7202,N_7219);
nand U7318 (N_7318,N_7285,N_7273);
xnor U7319 (N_7319,N_7238,N_7233);
nand U7320 (N_7320,N_7217,N_7296);
nor U7321 (N_7321,N_7251,N_7290);
nor U7322 (N_7322,N_7281,N_7210);
or U7323 (N_7323,N_7226,N_7214);
and U7324 (N_7324,N_7293,N_7221);
xnor U7325 (N_7325,N_7212,N_7294);
nor U7326 (N_7326,N_7235,N_7246);
and U7327 (N_7327,N_7278,N_7292);
nand U7328 (N_7328,N_7262,N_7298);
or U7329 (N_7329,N_7228,N_7272);
nand U7330 (N_7330,N_7237,N_7256);
xnor U7331 (N_7331,N_7243,N_7222);
or U7332 (N_7332,N_7203,N_7269);
nand U7333 (N_7333,N_7248,N_7299);
xor U7334 (N_7334,N_7218,N_7213);
or U7335 (N_7335,N_7289,N_7244);
nand U7336 (N_7336,N_7240,N_7205);
nand U7337 (N_7337,N_7224,N_7265);
nand U7338 (N_7338,N_7220,N_7258);
or U7339 (N_7339,N_7211,N_7231);
and U7340 (N_7340,N_7295,N_7288);
and U7341 (N_7341,N_7297,N_7283);
xor U7342 (N_7342,N_7250,N_7264);
and U7343 (N_7343,N_7255,N_7208);
nand U7344 (N_7344,N_7229,N_7239);
nor U7345 (N_7345,N_7284,N_7223);
nand U7346 (N_7346,N_7268,N_7280);
nand U7347 (N_7347,N_7266,N_7230);
or U7348 (N_7348,N_7286,N_7276);
and U7349 (N_7349,N_7277,N_7253);
nand U7350 (N_7350,N_7289,N_7209);
or U7351 (N_7351,N_7287,N_7206);
and U7352 (N_7352,N_7238,N_7257);
xor U7353 (N_7353,N_7258,N_7200);
nand U7354 (N_7354,N_7227,N_7225);
nor U7355 (N_7355,N_7255,N_7263);
nor U7356 (N_7356,N_7205,N_7255);
nand U7357 (N_7357,N_7268,N_7227);
and U7358 (N_7358,N_7261,N_7208);
nor U7359 (N_7359,N_7273,N_7206);
nand U7360 (N_7360,N_7233,N_7275);
nand U7361 (N_7361,N_7270,N_7209);
or U7362 (N_7362,N_7258,N_7223);
and U7363 (N_7363,N_7236,N_7217);
and U7364 (N_7364,N_7294,N_7283);
and U7365 (N_7365,N_7294,N_7221);
or U7366 (N_7366,N_7226,N_7267);
nor U7367 (N_7367,N_7260,N_7209);
nand U7368 (N_7368,N_7252,N_7222);
and U7369 (N_7369,N_7236,N_7273);
xnor U7370 (N_7370,N_7209,N_7266);
or U7371 (N_7371,N_7200,N_7277);
and U7372 (N_7372,N_7242,N_7272);
and U7373 (N_7373,N_7276,N_7221);
or U7374 (N_7374,N_7203,N_7268);
and U7375 (N_7375,N_7256,N_7253);
and U7376 (N_7376,N_7281,N_7230);
or U7377 (N_7377,N_7222,N_7296);
or U7378 (N_7378,N_7297,N_7247);
nand U7379 (N_7379,N_7231,N_7268);
nor U7380 (N_7380,N_7282,N_7228);
nand U7381 (N_7381,N_7215,N_7247);
nand U7382 (N_7382,N_7245,N_7217);
and U7383 (N_7383,N_7255,N_7287);
nand U7384 (N_7384,N_7293,N_7288);
and U7385 (N_7385,N_7245,N_7263);
or U7386 (N_7386,N_7294,N_7211);
nand U7387 (N_7387,N_7262,N_7282);
or U7388 (N_7388,N_7223,N_7209);
and U7389 (N_7389,N_7209,N_7227);
nand U7390 (N_7390,N_7275,N_7272);
nor U7391 (N_7391,N_7214,N_7207);
and U7392 (N_7392,N_7226,N_7255);
or U7393 (N_7393,N_7288,N_7255);
or U7394 (N_7394,N_7279,N_7245);
or U7395 (N_7395,N_7213,N_7254);
nor U7396 (N_7396,N_7238,N_7205);
or U7397 (N_7397,N_7200,N_7283);
nor U7398 (N_7398,N_7281,N_7255);
and U7399 (N_7399,N_7297,N_7294);
or U7400 (N_7400,N_7383,N_7308);
nand U7401 (N_7401,N_7397,N_7375);
nand U7402 (N_7402,N_7365,N_7362);
and U7403 (N_7403,N_7391,N_7395);
and U7404 (N_7404,N_7368,N_7357);
or U7405 (N_7405,N_7367,N_7355);
and U7406 (N_7406,N_7312,N_7333);
and U7407 (N_7407,N_7381,N_7344);
or U7408 (N_7408,N_7346,N_7348);
nor U7409 (N_7409,N_7345,N_7329);
nor U7410 (N_7410,N_7351,N_7306);
or U7411 (N_7411,N_7324,N_7311);
and U7412 (N_7412,N_7317,N_7307);
and U7413 (N_7413,N_7380,N_7379);
nand U7414 (N_7414,N_7332,N_7376);
or U7415 (N_7415,N_7334,N_7382);
and U7416 (N_7416,N_7315,N_7390);
or U7417 (N_7417,N_7342,N_7356);
or U7418 (N_7418,N_7321,N_7335);
nor U7419 (N_7419,N_7310,N_7386);
or U7420 (N_7420,N_7349,N_7314);
xor U7421 (N_7421,N_7331,N_7385);
or U7422 (N_7422,N_7302,N_7353);
and U7423 (N_7423,N_7341,N_7374);
xor U7424 (N_7424,N_7325,N_7303);
xnor U7425 (N_7425,N_7350,N_7352);
nand U7426 (N_7426,N_7316,N_7394);
nor U7427 (N_7427,N_7328,N_7388);
nand U7428 (N_7428,N_7322,N_7389);
nand U7429 (N_7429,N_7326,N_7392);
nor U7430 (N_7430,N_7370,N_7359);
and U7431 (N_7431,N_7301,N_7347);
and U7432 (N_7432,N_7399,N_7323);
and U7433 (N_7433,N_7377,N_7300);
nor U7434 (N_7434,N_7336,N_7327);
xnor U7435 (N_7435,N_7398,N_7369);
nand U7436 (N_7436,N_7318,N_7358);
xor U7437 (N_7437,N_7372,N_7313);
xor U7438 (N_7438,N_7396,N_7384);
or U7439 (N_7439,N_7364,N_7393);
and U7440 (N_7440,N_7373,N_7387);
xnor U7441 (N_7441,N_7363,N_7354);
or U7442 (N_7442,N_7305,N_7309);
and U7443 (N_7443,N_7371,N_7366);
xnor U7444 (N_7444,N_7320,N_7340);
xnor U7445 (N_7445,N_7330,N_7361);
nand U7446 (N_7446,N_7378,N_7339);
nand U7447 (N_7447,N_7319,N_7343);
nor U7448 (N_7448,N_7337,N_7304);
or U7449 (N_7449,N_7338,N_7360);
and U7450 (N_7450,N_7359,N_7399);
and U7451 (N_7451,N_7373,N_7336);
or U7452 (N_7452,N_7331,N_7391);
or U7453 (N_7453,N_7300,N_7358);
and U7454 (N_7454,N_7336,N_7332);
nor U7455 (N_7455,N_7334,N_7396);
and U7456 (N_7456,N_7365,N_7357);
xor U7457 (N_7457,N_7395,N_7302);
xor U7458 (N_7458,N_7376,N_7314);
or U7459 (N_7459,N_7304,N_7387);
or U7460 (N_7460,N_7311,N_7359);
and U7461 (N_7461,N_7336,N_7380);
or U7462 (N_7462,N_7389,N_7381);
xor U7463 (N_7463,N_7313,N_7356);
or U7464 (N_7464,N_7347,N_7323);
nor U7465 (N_7465,N_7370,N_7390);
nand U7466 (N_7466,N_7385,N_7370);
nor U7467 (N_7467,N_7310,N_7341);
nor U7468 (N_7468,N_7327,N_7334);
and U7469 (N_7469,N_7374,N_7377);
nand U7470 (N_7470,N_7337,N_7366);
nor U7471 (N_7471,N_7389,N_7351);
nor U7472 (N_7472,N_7399,N_7369);
nand U7473 (N_7473,N_7383,N_7376);
nor U7474 (N_7474,N_7379,N_7349);
or U7475 (N_7475,N_7329,N_7323);
nor U7476 (N_7476,N_7346,N_7304);
nor U7477 (N_7477,N_7383,N_7320);
nand U7478 (N_7478,N_7362,N_7390);
and U7479 (N_7479,N_7338,N_7355);
or U7480 (N_7480,N_7319,N_7323);
and U7481 (N_7481,N_7351,N_7399);
and U7482 (N_7482,N_7376,N_7344);
nand U7483 (N_7483,N_7328,N_7335);
nand U7484 (N_7484,N_7342,N_7382);
nand U7485 (N_7485,N_7344,N_7306);
and U7486 (N_7486,N_7332,N_7364);
xnor U7487 (N_7487,N_7361,N_7353);
or U7488 (N_7488,N_7353,N_7301);
nand U7489 (N_7489,N_7393,N_7338);
xor U7490 (N_7490,N_7375,N_7383);
xnor U7491 (N_7491,N_7349,N_7325);
nand U7492 (N_7492,N_7300,N_7387);
and U7493 (N_7493,N_7389,N_7345);
nand U7494 (N_7494,N_7345,N_7356);
xor U7495 (N_7495,N_7369,N_7325);
nand U7496 (N_7496,N_7331,N_7395);
nor U7497 (N_7497,N_7319,N_7302);
nand U7498 (N_7498,N_7373,N_7304);
and U7499 (N_7499,N_7320,N_7301);
and U7500 (N_7500,N_7409,N_7419);
nand U7501 (N_7501,N_7432,N_7455);
and U7502 (N_7502,N_7422,N_7447);
nor U7503 (N_7503,N_7457,N_7407);
and U7504 (N_7504,N_7414,N_7489);
nand U7505 (N_7505,N_7458,N_7465);
or U7506 (N_7506,N_7430,N_7429);
nor U7507 (N_7507,N_7497,N_7482);
xnor U7508 (N_7508,N_7402,N_7463);
and U7509 (N_7509,N_7441,N_7498);
nand U7510 (N_7510,N_7464,N_7484);
and U7511 (N_7511,N_7480,N_7462);
or U7512 (N_7512,N_7454,N_7485);
xnor U7513 (N_7513,N_7493,N_7475);
or U7514 (N_7514,N_7445,N_7421);
or U7515 (N_7515,N_7477,N_7452);
xor U7516 (N_7516,N_7486,N_7490);
xnor U7517 (N_7517,N_7424,N_7471);
and U7518 (N_7518,N_7438,N_7496);
and U7519 (N_7519,N_7467,N_7418);
nor U7520 (N_7520,N_7433,N_7423);
nand U7521 (N_7521,N_7405,N_7406);
nor U7522 (N_7522,N_7479,N_7468);
or U7523 (N_7523,N_7470,N_7488);
nor U7524 (N_7524,N_7437,N_7495);
nand U7525 (N_7525,N_7416,N_7446);
nand U7526 (N_7526,N_7449,N_7434);
nor U7527 (N_7527,N_7448,N_7400);
nor U7528 (N_7528,N_7426,N_7499);
xnor U7529 (N_7529,N_7473,N_7492);
or U7530 (N_7530,N_7415,N_7478);
and U7531 (N_7531,N_7403,N_7476);
and U7532 (N_7532,N_7487,N_7451);
nor U7533 (N_7533,N_7491,N_7401);
nand U7534 (N_7534,N_7412,N_7481);
nand U7535 (N_7535,N_7453,N_7413);
nand U7536 (N_7536,N_7450,N_7428);
xnor U7537 (N_7537,N_7436,N_7474);
nand U7538 (N_7538,N_7461,N_7460);
or U7539 (N_7539,N_7410,N_7472);
nand U7540 (N_7540,N_7411,N_7431);
nor U7541 (N_7541,N_7443,N_7417);
or U7542 (N_7542,N_7404,N_7439);
nand U7543 (N_7543,N_7483,N_7459);
nand U7544 (N_7544,N_7420,N_7408);
nor U7545 (N_7545,N_7466,N_7469);
nand U7546 (N_7546,N_7435,N_7425);
or U7547 (N_7547,N_7456,N_7427);
and U7548 (N_7548,N_7494,N_7440);
nand U7549 (N_7549,N_7442,N_7444);
and U7550 (N_7550,N_7409,N_7478);
nand U7551 (N_7551,N_7428,N_7457);
or U7552 (N_7552,N_7463,N_7481);
nand U7553 (N_7553,N_7488,N_7455);
nand U7554 (N_7554,N_7446,N_7466);
nor U7555 (N_7555,N_7471,N_7473);
or U7556 (N_7556,N_7408,N_7406);
or U7557 (N_7557,N_7448,N_7425);
and U7558 (N_7558,N_7419,N_7486);
nand U7559 (N_7559,N_7445,N_7457);
nand U7560 (N_7560,N_7481,N_7417);
nand U7561 (N_7561,N_7405,N_7411);
nor U7562 (N_7562,N_7430,N_7425);
nor U7563 (N_7563,N_7410,N_7430);
or U7564 (N_7564,N_7439,N_7424);
and U7565 (N_7565,N_7474,N_7428);
nor U7566 (N_7566,N_7428,N_7407);
and U7567 (N_7567,N_7461,N_7434);
or U7568 (N_7568,N_7426,N_7470);
nand U7569 (N_7569,N_7457,N_7491);
nor U7570 (N_7570,N_7488,N_7493);
nand U7571 (N_7571,N_7460,N_7423);
nand U7572 (N_7572,N_7442,N_7472);
nor U7573 (N_7573,N_7471,N_7439);
nor U7574 (N_7574,N_7408,N_7497);
and U7575 (N_7575,N_7419,N_7413);
and U7576 (N_7576,N_7405,N_7449);
nand U7577 (N_7577,N_7469,N_7433);
and U7578 (N_7578,N_7429,N_7483);
nand U7579 (N_7579,N_7482,N_7406);
xor U7580 (N_7580,N_7483,N_7437);
nand U7581 (N_7581,N_7454,N_7416);
or U7582 (N_7582,N_7414,N_7437);
nand U7583 (N_7583,N_7451,N_7480);
and U7584 (N_7584,N_7488,N_7418);
or U7585 (N_7585,N_7473,N_7479);
xor U7586 (N_7586,N_7406,N_7444);
nor U7587 (N_7587,N_7410,N_7438);
nor U7588 (N_7588,N_7401,N_7459);
nor U7589 (N_7589,N_7412,N_7432);
nor U7590 (N_7590,N_7429,N_7493);
or U7591 (N_7591,N_7475,N_7489);
nor U7592 (N_7592,N_7451,N_7464);
or U7593 (N_7593,N_7492,N_7413);
nor U7594 (N_7594,N_7430,N_7473);
nor U7595 (N_7595,N_7492,N_7439);
and U7596 (N_7596,N_7422,N_7418);
nand U7597 (N_7597,N_7471,N_7435);
nor U7598 (N_7598,N_7433,N_7439);
xor U7599 (N_7599,N_7440,N_7463);
xnor U7600 (N_7600,N_7544,N_7516);
nor U7601 (N_7601,N_7535,N_7596);
or U7602 (N_7602,N_7501,N_7594);
and U7603 (N_7603,N_7588,N_7570);
and U7604 (N_7604,N_7574,N_7587);
or U7605 (N_7605,N_7532,N_7531);
and U7606 (N_7606,N_7565,N_7549);
or U7607 (N_7607,N_7595,N_7599);
nand U7608 (N_7608,N_7541,N_7509);
and U7609 (N_7609,N_7542,N_7507);
nor U7610 (N_7610,N_7543,N_7579);
nand U7611 (N_7611,N_7548,N_7521);
nand U7612 (N_7612,N_7520,N_7527);
and U7613 (N_7613,N_7503,N_7502);
nor U7614 (N_7614,N_7590,N_7589);
nand U7615 (N_7615,N_7586,N_7552);
nand U7616 (N_7616,N_7554,N_7575);
nor U7617 (N_7617,N_7564,N_7517);
xnor U7618 (N_7618,N_7505,N_7577);
or U7619 (N_7619,N_7513,N_7539);
or U7620 (N_7620,N_7555,N_7510);
nor U7621 (N_7621,N_7545,N_7567);
xor U7622 (N_7622,N_7523,N_7562);
xnor U7623 (N_7623,N_7593,N_7504);
and U7624 (N_7624,N_7512,N_7511);
and U7625 (N_7625,N_7530,N_7569);
nand U7626 (N_7626,N_7572,N_7525);
or U7627 (N_7627,N_7550,N_7578);
or U7628 (N_7628,N_7561,N_7529);
nor U7629 (N_7629,N_7566,N_7592);
and U7630 (N_7630,N_7524,N_7568);
nor U7631 (N_7631,N_7580,N_7500);
nand U7632 (N_7632,N_7519,N_7522);
or U7633 (N_7633,N_7560,N_7581);
nor U7634 (N_7634,N_7556,N_7576);
and U7635 (N_7635,N_7508,N_7585);
and U7636 (N_7636,N_7518,N_7598);
and U7637 (N_7637,N_7558,N_7536);
and U7638 (N_7638,N_7533,N_7537);
xor U7639 (N_7639,N_7597,N_7557);
and U7640 (N_7640,N_7506,N_7553);
nor U7641 (N_7641,N_7528,N_7573);
nor U7642 (N_7642,N_7514,N_7551);
xnor U7643 (N_7643,N_7584,N_7582);
nand U7644 (N_7644,N_7540,N_7563);
nand U7645 (N_7645,N_7547,N_7571);
or U7646 (N_7646,N_7538,N_7583);
nand U7647 (N_7647,N_7515,N_7526);
or U7648 (N_7648,N_7546,N_7534);
nand U7649 (N_7649,N_7591,N_7559);
nor U7650 (N_7650,N_7572,N_7587);
and U7651 (N_7651,N_7507,N_7508);
and U7652 (N_7652,N_7573,N_7586);
nand U7653 (N_7653,N_7596,N_7592);
nor U7654 (N_7654,N_7591,N_7593);
and U7655 (N_7655,N_7532,N_7593);
and U7656 (N_7656,N_7516,N_7555);
nand U7657 (N_7657,N_7533,N_7563);
nand U7658 (N_7658,N_7598,N_7544);
or U7659 (N_7659,N_7543,N_7530);
and U7660 (N_7660,N_7565,N_7508);
nor U7661 (N_7661,N_7533,N_7523);
and U7662 (N_7662,N_7571,N_7521);
or U7663 (N_7663,N_7564,N_7527);
xor U7664 (N_7664,N_7565,N_7539);
and U7665 (N_7665,N_7550,N_7500);
or U7666 (N_7666,N_7515,N_7568);
nand U7667 (N_7667,N_7552,N_7533);
nor U7668 (N_7668,N_7555,N_7563);
or U7669 (N_7669,N_7541,N_7542);
xor U7670 (N_7670,N_7524,N_7528);
nand U7671 (N_7671,N_7515,N_7525);
nand U7672 (N_7672,N_7528,N_7538);
xnor U7673 (N_7673,N_7505,N_7573);
nor U7674 (N_7674,N_7592,N_7575);
nor U7675 (N_7675,N_7532,N_7555);
nor U7676 (N_7676,N_7535,N_7569);
xnor U7677 (N_7677,N_7528,N_7580);
or U7678 (N_7678,N_7584,N_7538);
xor U7679 (N_7679,N_7537,N_7595);
nand U7680 (N_7680,N_7519,N_7529);
xnor U7681 (N_7681,N_7582,N_7515);
nor U7682 (N_7682,N_7583,N_7534);
nor U7683 (N_7683,N_7569,N_7511);
nand U7684 (N_7684,N_7589,N_7514);
nand U7685 (N_7685,N_7576,N_7514);
xnor U7686 (N_7686,N_7586,N_7587);
xnor U7687 (N_7687,N_7546,N_7561);
or U7688 (N_7688,N_7533,N_7595);
and U7689 (N_7689,N_7558,N_7525);
and U7690 (N_7690,N_7597,N_7579);
or U7691 (N_7691,N_7522,N_7585);
and U7692 (N_7692,N_7549,N_7541);
or U7693 (N_7693,N_7591,N_7543);
nand U7694 (N_7694,N_7578,N_7539);
and U7695 (N_7695,N_7510,N_7504);
and U7696 (N_7696,N_7590,N_7505);
and U7697 (N_7697,N_7509,N_7542);
nor U7698 (N_7698,N_7525,N_7566);
and U7699 (N_7699,N_7527,N_7517);
and U7700 (N_7700,N_7655,N_7635);
and U7701 (N_7701,N_7662,N_7648);
and U7702 (N_7702,N_7619,N_7626);
nand U7703 (N_7703,N_7636,N_7631);
or U7704 (N_7704,N_7666,N_7659);
xor U7705 (N_7705,N_7643,N_7678);
nand U7706 (N_7706,N_7601,N_7670);
nand U7707 (N_7707,N_7652,N_7609);
xor U7708 (N_7708,N_7681,N_7660);
and U7709 (N_7709,N_7672,N_7605);
and U7710 (N_7710,N_7606,N_7677);
and U7711 (N_7711,N_7625,N_7639);
and U7712 (N_7712,N_7650,N_7667);
nand U7713 (N_7713,N_7632,N_7696);
or U7714 (N_7714,N_7600,N_7657);
nand U7715 (N_7715,N_7674,N_7620);
nand U7716 (N_7716,N_7630,N_7602);
nand U7717 (N_7717,N_7679,N_7688);
xnor U7718 (N_7718,N_7638,N_7611);
or U7719 (N_7719,N_7604,N_7695);
or U7720 (N_7720,N_7633,N_7675);
and U7721 (N_7721,N_7612,N_7694);
or U7722 (N_7722,N_7687,N_7663);
nand U7723 (N_7723,N_7676,N_7697);
or U7724 (N_7724,N_7653,N_7607);
nor U7725 (N_7725,N_7640,N_7699);
nor U7726 (N_7726,N_7647,N_7685);
or U7727 (N_7727,N_7654,N_7644);
nand U7728 (N_7728,N_7686,N_7698);
nand U7729 (N_7729,N_7668,N_7627);
and U7730 (N_7730,N_7629,N_7603);
and U7731 (N_7731,N_7680,N_7616);
nand U7732 (N_7732,N_7622,N_7658);
nor U7733 (N_7733,N_7683,N_7691);
nand U7734 (N_7734,N_7692,N_7613);
and U7735 (N_7735,N_7634,N_7645);
and U7736 (N_7736,N_7623,N_7651);
or U7737 (N_7737,N_7614,N_7671);
xor U7738 (N_7738,N_7664,N_7656);
nand U7739 (N_7739,N_7624,N_7610);
and U7740 (N_7740,N_7617,N_7641);
nor U7741 (N_7741,N_7673,N_7608);
and U7742 (N_7742,N_7615,N_7689);
and U7743 (N_7743,N_7618,N_7684);
or U7744 (N_7744,N_7690,N_7693);
or U7745 (N_7745,N_7665,N_7649);
and U7746 (N_7746,N_7642,N_7682);
nor U7747 (N_7747,N_7637,N_7646);
or U7748 (N_7748,N_7628,N_7669);
and U7749 (N_7749,N_7621,N_7661);
nor U7750 (N_7750,N_7663,N_7673);
and U7751 (N_7751,N_7684,N_7687);
nand U7752 (N_7752,N_7614,N_7611);
and U7753 (N_7753,N_7607,N_7691);
nor U7754 (N_7754,N_7627,N_7624);
nor U7755 (N_7755,N_7602,N_7687);
or U7756 (N_7756,N_7697,N_7652);
nand U7757 (N_7757,N_7630,N_7665);
xor U7758 (N_7758,N_7637,N_7643);
or U7759 (N_7759,N_7639,N_7653);
and U7760 (N_7760,N_7681,N_7678);
xor U7761 (N_7761,N_7675,N_7682);
or U7762 (N_7762,N_7664,N_7651);
nand U7763 (N_7763,N_7659,N_7638);
nor U7764 (N_7764,N_7679,N_7695);
nand U7765 (N_7765,N_7628,N_7685);
and U7766 (N_7766,N_7623,N_7632);
nand U7767 (N_7767,N_7617,N_7679);
nor U7768 (N_7768,N_7677,N_7626);
or U7769 (N_7769,N_7648,N_7629);
nand U7770 (N_7770,N_7656,N_7668);
and U7771 (N_7771,N_7679,N_7683);
and U7772 (N_7772,N_7679,N_7690);
or U7773 (N_7773,N_7692,N_7645);
nor U7774 (N_7774,N_7626,N_7682);
or U7775 (N_7775,N_7661,N_7622);
xnor U7776 (N_7776,N_7683,N_7601);
nand U7777 (N_7777,N_7688,N_7676);
nand U7778 (N_7778,N_7699,N_7634);
nand U7779 (N_7779,N_7637,N_7648);
and U7780 (N_7780,N_7603,N_7694);
nor U7781 (N_7781,N_7662,N_7630);
and U7782 (N_7782,N_7630,N_7624);
or U7783 (N_7783,N_7614,N_7601);
or U7784 (N_7784,N_7654,N_7634);
or U7785 (N_7785,N_7645,N_7603);
nor U7786 (N_7786,N_7684,N_7635);
nor U7787 (N_7787,N_7640,N_7689);
nor U7788 (N_7788,N_7655,N_7624);
nand U7789 (N_7789,N_7641,N_7695);
and U7790 (N_7790,N_7611,N_7633);
nor U7791 (N_7791,N_7608,N_7641);
nor U7792 (N_7792,N_7632,N_7697);
and U7793 (N_7793,N_7693,N_7645);
nand U7794 (N_7794,N_7693,N_7619);
xnor U7795 (N_7795,N_7653,N_7651);
and U7796 (N_7796,N_7644,N_7607);
nand U7797 (N_7797,N_7682,N_7633);
and U7798 (N_7798,N_7643,N_7697);
or U7799 (N_7799,N_7649,N_7679);
nor U7800 (N_7800,N_7795,N_7743);
nor U7801 (N_7801,N_7761,N_7771);
or U7802 (N_7802,N_7757,N_7701);
and U7803 (N_7803,N_7748,N_7764);
and U7804 (N_7804,N_7782,N_7716);
nand U7805 (N_7805,N_7793,N_7702);
or U7806 (N_7806,N_7739,N_7721);
and U7807 (N_7807,N_7746,N_7778);
and U7808 (N_7808,N_7727,N_7776);
nand U7809 (N_7809,N_7768,N_7753);
nor U7810 (N_7810,N_7762,N_7738);
or U7811 (N_7811,N_7708,N_7728);
nor U7812 (N_7812,N_7774,N_7720);
and U7813 (N_7813,N_7703,N_7737);
or U7814 (N_7814,N_7723,N_7785);
xnor U7815 (N_7815,N_7736,N_7773);
xor U7816 (N_7816,N_7710,N_7713);
nor U7817 (N_7817,N_7724,N_7715);
nor U7818 (N_7818,N_7731,N_7784);
xor U7819 (N_7819,N_7758,N_7726);
xor U7820 (N_7820,N_7797,N_7766);
and U7821 (N_7821,N_7729,N_7730);
and U7822 (N_7822,N_7717,N_7704);
or U7823 (N_7823,N_7790,N_7742);
nor U7824 (N_7824,N_7732,N_7792);
and U7825 (N_7825,N_7765,N_7754);
or U7826 (N_7826,N_7781,N_7794);
nor U7827 (N_7827,N_7751,N_7711);
nand U7828 (N_7828,N_7750,N_7725);
or U7829 (N_7829,N_7712,N_7735);
nand U7830 (N_7830,N_7709,N_7700);
and U7831 (N_7831,N_7770,N_7791);
or U7832 (N_7832,N_7733,N_7719);
nor U7833 (N_7833,N_7789,N_7796);
nor U7834 (N_7834,N_7734,N_7788);
nand U7835 (N_7835,N_7772,N_7755);
nand U7836 (N_7836,N_7786,N_7705);
nor U7837 (N_7837,N_7799,N_7775);
or U7838 (N_7838,N_7756,N_7749);
and U7839 (N_7839,N_7780,N_7718);
or U7840 (N_7840,N_7787,N_7783);
nor U7841 (N_7841,N_7714,N_7769);
xor U7842 (N_7842,N_7747,N_7707);
nor U7843 (N_7843,N_7744,N_7752);
xor U7844 (N_7844,N_7760,N_7745);
or U7845 (N_7845,N_7777,N_7779);
and U7846 (N_7846,N_7706,N_7741);
nand U7847 (N_7847,N_7798,N_7740);
nand U7848 (N_7848,N_7763,N_7759);
xor U7849 (N_7849,N_7722,N_7767);
xor U7850 (N_7850,N_7755,N_7766);
or U7851 (N_7851,N_7730,N_7787);
nand U7852 (N_7852,N_7730,N_7796);
xor U7853 (N_7853,N_7739,N_7795);
xnor U7854 (N_7854,N_7746,N_7745);
nand U7855 (N_7855,N_7720,N_7768);
nand U7856 (N_7856,N_7730,N_7770);
nand U7857 (N_7857,N_7750,N_7774);
nand U7858 (N_7858,N_7781,N_7785);
nor U7859 (N_7859,N_7708,N_7727);
and U7860 (N_7860,N_7797,N_7785);
or U7861 (N_7861,N_7770,N_7704);
and U7862 (N_7862,N_7740,N_7732);
nor U7863 (N_7863,N_7709,N_7797);
and U7864 (N_7864,N_7754,N_7771);
and U7865 (N_7865,N_7798,N_7759);
xor U7866 (N_7866,N_7741,N_7782);
or U7867 (N_7867,N_7712,N_7746);
and U7868 (N_7868,N_7774,N_7752);
and U7869 (N_7869,N_7706,N_7704);
xor U7870 (N_7870,N_7733,N_7763);
or U7871 (N_7871,N_7770,N_7739);
nand U7872 (N_7872,N_7748,N_7743);
and U7873 (N_7873,N_7761,N_7712);
or U7874 (N_7874,N_7711,N_7706);
nand U7875 (N_7875,N_7795,N_7735);
nand U7876 (N_7876,N_7714,N_7744);
xor U7877 (N_7877,N_7717,N_7782);
or U7878 (N_7878,N_7737,N_7771);
nor U7879 (N_7879,N_7785,N_7704);
nor U7880 (N_7880,N_7748,N_7774);
nor U7881 (N_7881,N_7743,N_7764);
nor U7882 (N_7882,N_7798,N_7737);
nand U7883 (N_7883,N_7719,N_7753);
or U7884 (N_7884,N_7720,N_7726);
nor U7885 (N_7885,N_7790,N_7794);
or U7886 (N_7886,N_7784,N_7755);
and U7887 (N_7887,N_7708,N_7715);
and U7888 (N_7888,N_7703,N_7701);
nor U7889 (N_7889,N_7733,N_7724);
nand U7890 (N_7890,N_7740,N_7751);
nor U7891 (N_7891,N_7798,N_7706);
nor U7892 (N_7892,N_7729,N_7775);
nand U7893 (N_7893,N_7747,N_7783);
nand U7894 (N_7894,N_7789,N_7739);
or U7895 (N_7895,N_7792,N_7749);
and U7896 (N_7896,N_7790,N_7741);
and U7897 (N_7897,N_7775,N_7752);
xnor U7898 (N_7898,N_7733,N_7790);
or U7899 (N_7899,N_7712,N_7755);
nor U7900 (N_7900,N_7834,N_7818);
or U7901 (N_7901,N_7888,N_7803);
nand U7902 (N_7902,N_7847,N_7848);
nand U7903 (N_7903,N_7829,N_7853);
xor U7904 (N_7904,N_7895,N_7807);
or U7905 (N_7905,N_7878,N_7822);
or U7906 (N_7906,N_7815,N_7845);
nor U7907 (N_7907,N_7826,N_7855);
nor U7908 (N_7908,N_7814,N_7824);
nand U7909 (N_7909,N_7894,N_7843);
and U7910 (N_7910,N_7879,N_7801);
and U7911 (N_7911,N_7863,N_7832);
and U7912 (N_7912,N_7893,N_7867);
or U7913 (N_7913,N_7817,N_7846);
nor U7914 (N_7914,N_7802,N_7885);
xor U7915 (N_7915,N_7841,N_7865);
nand U7916 (N_7916,N_7821,N_7808);
or U7917 (N_7917,N_7827,N_7820);
nor U7918 (N_7918,N_7881,N_7825);
xnor U7919 (N_7919,N_7839,N_7889);
xor U7920 (N_7920,N_7819,N_7892);
nand U7921 (N_7921,N_7854,N_7874);
and U7922 (N_7922,N_7870,N_7833);
or U7923 (N_7923,N_7868,N_7871);
and U7924 (N_7924,N_7898,N_7837);
nor U7925 (N_7925,N_7828,N_7896);
nand U7926 (N_7926,N_7872,N_7851);
or U7927 (N_7927,N_7852,N_7813);
or U7928 (N_7928,N_7861,N_7890);
or U7929 (N_7929,N_7857,N_7856);
nor U7930 (N_7930,N_7899,N_7876);
and U7931 (N_7931,N_7840,N_7882);
nand U7932 (N_7932,N_7836,N_7884);
or U7933 (N_7933,N_7869,N_7831);
nor U7934 (N_7934,N_7873,N_7858);
nor U7935 (N_7935,N_7897,N_7804);
nand U7936 (N_7936,N_7887,N_7800);
nor U7937 (N_7937,N_7875,N_7880);
and U7938 (N_7938,N_7860,N_7842);
or U7939 (N_7939,N_7849,N_7864);
nand U7940 (N_7940,N_7883,N_7823);
nand U7941 (N_7941,N_7877,N_7830);
or U7942 (N_7942,N_7838,N_7859);
nand U7943 (N_7943,N_7810,N_7866);
and U7944 (N_7944,N_7805,N_7850);
and U7945 (N_7945,N_7812,N_7816);
or U7946 (N_7946,N_7886,N_7811);
nor U7947 (N_7947,N_7835,N_7862);
or U7948 (N_7948,N_7891,N_7809);
nand U7949 (N_7949,N_7844,N_7806);
nand U7950 (N_7950,N_7811,N_7896);
and U7951 (N_7951,N_7878,N_7844);
and U7952 (N_7952,N_7891,N_7856);
nor U7953 (N_7953,N_7803,N_7843);
and U7954 (N_7954,N_7843,N_7845);
and U7955 (N_7955,N_7817,N_7809);
and U7956 (N_7956,N_7818,N_7860);
nand U7957 (N_7957,N_7888,N_7853);
nor U7958 (N_7958,N_7856,N_7863);
and U7959 (N_7959,N_7802,N_7862);
nand U7960 (N_7960,N_7898,N_7880);
and U7961 (N_7961,N_7896,N_7800);
nor U7962 (N_7962,N_7848,N_7865);
nor U7963 (N_7963,N_7872,N_7825);
nand U7964 (N_7964,N_7825,N_7882);
nor U7965 (N_7965,N_7869,N_7876);
nand U7966 (N_7966,N_7894,N_7801);
nor U7967 (N_7967,N_7848,N_7896);
xor U7968 (N_7968,N_7861,N_7835);
nand U7969 (N_7969,N_7802,N_7813);
nand U7970 (N_7970,N_7892,N_7826);
and U7971 (N_7971,N_7855,N_7869);
nand U7972 (N_7972,N_7853,N_7893);
and U7973 (N_7973,N_7857,N_7804);
nand U7974 (N_7974,N_7807,N_7873);
nand U7975 (N_7975,N_7808,N_7835);
or U7976 (N_7976,N_7817,N_7856);
nor U7977 (N_7977,N_7887,N_7883);
or U7978 (N_7978,N_7898,N_7854);
and U7979 (N_7979,N_7800,N_7814);
xor U7980 (N_7980,N_7823,N_7867);
or U7981 (N_7981,N_7873,N_7887);
and U7982 (N_7982,N_7872,N_7888);
or U7983 (N_7983,N_7863,N_7897);
nand U7984 (N_7984,N_7850,N_7823);
and U7985 (N_7985,N_7897,N_7851);
nand U7986 (N_7986,N_7886,N_7832);
and U7987 (N_7987,N_7891,N_7849);
nand U7988 (N_7988,N_7884,N_7888);
and U7989 (N_7989,N_7857,N_7838);
nor U7990 (N_7990,N_7888,N_7838);
and U7991 (N_7991,N_7895,N_7841);
or U7992 (N_7992,N_7821,N_7829);
nor U7993 (N_7993,N_7816,N_7830);
or U7994 (N_7994,N_7877,N_7898);
and U7995 (N_7995,N_7877,N_7854);
and U7996 (N_7996,N_7869,N_7842);
or U7997 (N_7997,N_7845,N_7857);
nand U7998 (N_7998,N_7867,N_7811);
and U7999 (N_7999,N_7811,N_7888);
and U8000 (N_8000,N_7928,N_7990);
or U8001 (N_8001,N_7950,N_7924);
and U8002 (N_8002,N_7920,N_7971);
nor U8003 (N_8003,N_7965,N_7951);
xor U8004 (N_8004,N_7915,N_7952);
nand U8005 (N_8005,N_7985,N_7979);
and U8006 (N_8006,N_7937,N_7983);
nor U8007 (N_8007,N_7930,N_7954);
and U8008 (N_8008,N_7992,N_7977);
nor U8009 (N_8009,N_7963,N_7932);
nand U8010 (N_8010,N_7997,N_7912);
nor U8011 (N_8011,N_7989,N_7940);
nand U8012 (N_8012,N_7976,N_7961);
nor U8013 (N_8013,N_7964,N_7918);
nor U8014 (N_8014,N_7970,N_7933);
and U8015 (N_8015,N_7974,N_7939);
or U8016 (N_8016,N_7973,N_7927);
and U8017 (N_8017,N_7931,N_7929);
and U8018 (N_8018,N_7957,N_7911);
or U8019 (N_8019,N_7978,N_7942);
or U8020 (N_8020,N_7909,N_7945);
or U8021 (N_8021,N_7943,N_7999);
and U8022 (N_8022,N_7935,N_7903);
nor U8023 (N_8023,N_7998,N_7981);
nand U8024 (N_8024,N_7987,N_7902);
and U8025 (N_8025,N_7960,N_7955);
and U8026 (N_8026,N_7938,N_7921);
xnor U8027 (N_8027,N_7980,N_7925);
nor U8028 (N_8028,N_7958,N_7996);
or U8029 (N_8029,N_7994,N_7922);
or U8030 (N_8030,N_7926,N_7914);
nor U8031 (N_8031,N_7962,N_7968);
or U8032 (N_8032,N_7993,N_7966);
nand U8033 (N_8033,N_7906,N_7934);
and U8034 (N_8034,N_7991,N_7947);
nor U8035 (N_8035,N_7984,N_7969);
and U8036 (N_8036,N_7908,N_7967);
or U8037 (N_8037,N_7972,N_7988);
and U8038 (N_8038,N_7995,N_7956);
nand U8039 (N_8039,N_7917,N_7986);
nand U8040 (N_8040,N_7901,N_7948);
nor U8041 (N_8041,N_7904,N_7975);
and U8042 (N_8042,N_7907,N_7949);
nor U8043 (N_8043,N_7953,N_7944);
nand U8044 (N_8044,N_7982,N_7936);
and U8045 (N_8045,N_7905,N_7941);
nor U8046 (N_8046,N_7919,N_7959);
and U8047 (N_8047,N_7923,N_7913);
and U8048 (N_8048,N_7946,N_7910);
nand U8049 (N_8049,N_7900,N_7916);
nor U8050 (N_8050,N_7980,N_7934);
or U8051 (N_8051,N_7955,N_7941);
nor U8052 (N_8052,N_7984,N_7999);
xor U8053 (N_8053,N_7929,N_7921);
nand U8054 (N_8054,N_7930,N_7960);
nand U8055 (N_8055,N_7997,N_7927);
nand U8056 (N_8056,N_7909,N_7954);
and U8057 (N_8057,N_7917,N_7992);
nor U8058 (N_8058,N_7961,N_7995);
nand U8059 (N_8059,N_7998,N_7916);
nand U8060 (N_8060,N_7958,N_7906);
and U8061 (N_8061,N_7956,N_7974);
or U8062 (N_8062,N_7915,N_7985);
or U8063 (N_8063,N_7990,N_7911);
nand U8064 (N_8064,N_7974,N_7995);
nand U8065 (N_8065,N_7905,N_7932);
nand U8066 (N_8066,N_7928,N_7995);
nor U8067 (N_8067,N_7990,N_7998);
and U8068 (N_8068,N_7968,N_7943);
nor U8069 (N_8069,N_7905,N_7901);
and U8070 (N_8070,N_7908,N_7905);
nor U8071 (N_8071,N_7991,N_7989);
and U8072 (N_8072,N_7938,N_7997);
or U8073 (N_8073,N_7990,N_7993);
and U8074 (N_8074,N_7969,N_7933);
nor U8075 (N_8075,N_7923,N_7932);
nor U8076 (N_8076,N_7909,N_7979);
or U8077 (N_8077,N_7956,N_7965);
nand U8078 (N_8078,N_7988,N_7911);
and U8079 (N_8079,N_7920,N_7983);
or U8080 (N_8080,N_7928,N_7974);
nor U8081 (N_8081,N_7955,N_7949);
and U8082 (N_8082,N_7906,N_7917);
nand U8083 (N_8083,N_7947,N_7963);
nand U8084 (N_8084,N_7908,N_7922);
nand U8085 (N_8085,N_7912,N_7915);
and U8086 (N_8086,N_7916,N_7990);
nand U8087 (N_8087,N_7994,N_7978);
and U8088 (N_8088,N_7951,N_7956);
or U8089 (N_8089,N_7979,N_7960);
nand U8090 (N_8090,N_7958,N_7911);
or U8091 (N_8091,N_7920,N_7933);
nand U8092 (N_8092,N_7952,N_7920);
nand U8093 (N_8093,N_7951,N_7986);
nand U8094 (N_8094,N_7940,N_7930);
and U8095 (N_8095,N_7963,N_7902);
nand U8096 (N_8096,N_7993,N_7989);
or U8097 (N_8097,N_7944,N_7972);
nand U8098 (N_8098,N_7904,N_7977);
or U8099 (N_8099,N_7965,N_7913);
or U8100 (N_8100,N_8000,N_8062);
xor U8101 (N_8101,N_8025,N_8058);
and U8102 (N_8102,N_8047,N_8092);
or U8103 (N_8103,N_8035,N_8007);
or U8104 (N_8104,N_8087,N_8078);
nand U8105 (N_8105,N_8086,N_8002);
nor U8106 (N_8106,N_8046,N_8045);
and U8107 (N_8107,N_8032,N_8097);
or U8108 (N_8108,N_8056,N_8026);
or U8109 (N_8109,N_8041,N_8006);
or U8110 (N_8110,N_8014,N_8031);
nor U8111 (N_8111,N_8059,N_8089);
nor U8112 (N_8112,N_8091,N_8090);
nor U8113 (N_8113,N_8080,N_8009);
nand U8114 (N_8114,N_8039,N_8008);
and U8115 (N_8115,N_8005,N_8082);
nor U8116 (N_8116,N_8052,N_8063);
or U8117 (N_8117,N_8060,N_8021);
xor U8118 (N_8118,N_8034,N_8013);
or U8119 (N_8119,N_8094,N_8048);
nor U8120 (N_8120,N_8003,N_8072);
or U8121 (N_8121,N_8027,N_8095);
nor U8122 (N_8122,N_8038,N_8044);
nand U8123 (N_8123,N_8068,N_8053);
xnor U8124 (N_8124,N_8070,N_8024);
or U8125 (N_8125,N_8017,N_8042);
nand U8126 (N_8126,N_8093,N_8030);
xnor U8127 (N_8127,N_8057,N_8033);
nor U8128 (N_8128,N_8077,N_8054);
xor U8129 (N_8129,N_8018,N_8079);
or U8130 (N_8130,N_8022,N_8083);
xnor U8131 (N_8131,N_8040,N_8075);
nand U8132 (N_8132,N_8099,N_8011);
nand U8133 (N_8133,N_8029,N_8073);
xnor U8134 (N_8134,N_8043,N_8019);
xor U8135 (N_8135,N_8065,N_8051);
nand U8136 (N_8136,N_8012,N_8037);
nor U8137 (N_8137,N_8074,N_8049);
nand U8138 (N_8138,N_8088,N_8023);
and U8139 (N_8139,N_8055,N_8001);
nand U8140 (N_8140,N_8036,N_8081);
or U8141 (N_8141,N_8010,N_8098);
nand U8142 (N_8142,N_8076,N_8084);
or U8143 (N_8143,N_8066,N_8085);
or U8144 (N_8144,N_8071,N_8004);
or U8145 (N_8145,N_8028,N_8069);
nand U8146 (N_8146,N_8015,N_8050);
nand U8147 (N_8147,N_8064,N_8061);
xnor U8148 (N_8148,N_8096,N_8067);
nor U8149 (N_8149,N_8016,N_8020);
xor U8150 (N_8150,N_8007,N_8020);
and U8151 (N_8151,N_8077,N_8080);
and U8152 (N_8152,N_8062,N_8022);
nor U8153 (N_8153,N_8059,N_8011);
xor U8154 (N_8154,N_8098,N_8082);
nor U8155 (N_8155,N_8031,N_8023);
xor U8156 (N_8156,N_8008,N_8006);
or U8157 (N_8157,N_8043,N_8036);
nand U8158 (N_8158,N_8074,N_8075);
nor U8159 (N_8159,N_8011,N_8052);
and U8160 (N_8160,N_8047,N_8090);
nand U8161 (N_8161,N_8005,N_8061);
or U8162 (N_8162,N_8031,N_8099);
and U8163 (N_8163,N_8002,N_8083);
nor U8164 (N_8164,N_8005,N_8062);
nor U8165 (N_8165,N_8096,N_8082);
nand U8166 (N_8166,N_8052,N_8022);
nor U8167 (N_8167,N_8065,N_8089);
nor U8168 (N_8168,N_8097,N_8029);
and U8169 (N_8169,N_8021,N_8016);
or U8170 (N_8170,N_8002,N_8029);
nand U8171 (N_8171,N_8060,N_8055);
and U8172 (N_8172,N_8005,N_8078);
or U8173 (N_8173,N_8078,N_8066);
and U8174 (N_8174,N_8016,N_8008);
nor U8175 (N_8175,N_8023,N_8075);
nand U8176 (N_8176,N_8095,N_8025);
nand U8177 (N_8177,N_8074,N_8016);
nand U8178 (N_8178,N_8008,N_8098);
and U8179 (N_8179,N_8023,N_8044);
nand U8180 (N_8180,N_8084,N_8099);
or U8181 (N_8181,N_8049,N_8012);
or U8182 (N_8182,N_8008,N_8095);
nand U8183 (N_8183,N_8058,N_8046);
nand U8184 (N_8184,N_8018,N_8074);
nand U8185 (N_8185,N_8026,N_8001);
or U8186 (N_8186,N_8004,N_8051);
and U8187 (N_8187,N_8027,N_8013);
or U8188 (N_8188,N_8070,N_8099);
nor U8189 (N_8189,N_8047,N_8088);
nor U8190 (N_8190,N_8000,N_8052);
xnor U8191 (N_8191,N_8086,N_8053);
xnor U8192 (N_8192,N_8033,N_8098);
nand U8193 (N_8193,N_8062,N_8036);
nor U8194 (N_8194,N_8035,N_8091);
or U8195 (N_8195,N_8083,N_8042);
and U8196 (N_8196,N_8036,N_8059);
or U8197 (N_8197,N_8006,N_8028);
nand U8198 (N_8198,N_8067,N_8023);
and U8199 (N_8199,N_8083,N_8044);
and U8200 (N_8200,N_8157,N_8125);
nor U8201 (N_8201,N_8131,N_8182);
nand U8202 (N_8202,N_8192,N_8143);
or U8203 (N_8203,N_8109,N_8171);
nand U8204 (N_8204,N_8188,N_8129);
xnor U8205 (N_8205,N_8145,N_8166);
or U8206 (N_8206,N_8116,N_8136);
and U8207 (N_8207,N_8120,N_8132);
nor U8208 (N_8208,N_8100,N_8119);
nor U8209 (N_8209,N_8189,N_8137);
and U8210 (N_8210,N_8193,N_8177);
nand U8211 (N_8211,N_8150,N_8113);
or U8212 (N_8212,N_8183,N_8165);
nand U8213 (N_8213,N_8176,N_8101);
xnor U8214 (N_8214,N_8197,N_8138);
nand U8215 (N_8215,N_8122,N_8186);
or U8216 (N_8216,N_8195,N_8126);
nand U8217 (N_8217,N_8187,N_8154);
and U8218 (N_8218,N_8160,N_8156);
and U8219 (N_8219,N_8163,N_8139);
nor U8220 (N_8220,N_8124,N_8161);
and U8221 (N_8221,N_8191,N_8155);
nor U8222 (N_8222,N_8162,N_8111);
nor U8223 (N_8223,N_8181,N_8148);
xor U8224 (N_8224,N_8151,N_8123);
nand U8225 (N_8225,N_8121,N_8198);
nand U8226 (N_8226,N_8179,N_8142);
or U8227 (N_8227,N_8102,N_8167);
nand U8228 (N_8228,N_8134,N_8133);
xor U8229 (N_8229,N_8178,N_8184);
and U8230 (N_8230,N_8110,N_8115);
and U8231 (N_8231,N_8117,N_8196);
and U8232 (N_8232,N_8112,N_8190);
nor U8233 (N_8233,N_8175,N_8194);
nand U8234 (N_8234,N_8149,N_8114);
nor U8235 (N_8235,N_8103,N_8130);
nand U8236 (N_8236,N_8147,N_8105);
nor U8237 (N_8237,N_8106,N_8158);
or U8238 (N_8238,N_8128,N_8135);
nor U8239 (N_8239,N_8144,N_8140);
or U8240 (N_8240,N_8174,N_8180);
and U8241 (N_8241,N_8107,N_8169);
nor U8242 (N_8242,N_8104,N_8185);
nor U8243 (N_8243,N_8170,N_8159);
nor U8244 (N_8244,N_8199,N_8118);
or U8245 (N_8245,N_8164,N_8141);
nand U8246 (N_8246,N_8152,N_8146);
nand U8247 (N_8247,N_8108,N_8168);
nor U8248 (N_8248,N_8153,N_8172);
or U8249 (N_8249,N_8173,N_8127);
or U8250 (N_8250,N_8174,N_8110);
nor U8251 (N_8251,N_8174,N_8118);
or U8252 (N_8252,N_8135,N_8162);
nand U8253 (N_8253,N_8113,N_8163);
and U8254 (N_8254,N_8177,N_8126);
xnor U8255 (N_8255,N_8182,N_8106);
nand U8256 (N_8256,N_8130,N_8123);
nand U8257 (N_8257,N_8172,N_8178);
nor U8258 (N_8258,N_8133,N_8192);
nand U8259 (N_8259,N_8126,N_8185);
or U8260 (N_8260,N_8182,N_8166);
nor U8261 (N_8261,N_8134,N_8158);
nor U8262 (N_8262,N_8108,N_8135);
and U8263 (N_8263,N_8110,N_8166);
or U8264 (N_8264,N_8156,N_8157);
nor U8265 (N_8265,N_8186,N_8170);
or U8266 (N_8266,N_8165,N_8168);
nor U8267 (N_8267,N_8127,N_8153);
nor U8268 (N_8268,N_8195,N_8198);
and U8269 (N_8269,N_8136,N_8180);
nor U8270 (N_8270,N_8132,N_8139);
nor U8271 (N_8271,N_8189,N_8199);
and U8272 (N_8272,N_8173,N_8151);
nand U8273 (N_8273,N_8154,N_8115);
nand U8274 (N_8274,N_8100,N_8196);
nor U8275 (N_8275,N_8173,N_8145);
nand U8276 (N_8276,N_8108,N_8115);
xnor U8277 (N_8277,N_8195,N_8143);
and U8278 (N_8278,N_8175,N_8153);
or U8279 (N_8279,N_8130,N_8107);
nor U8280 (N_8280,N_8132,N_8118);
nor U8281 (N_8281,N_8152,N_8197);
nand U8282 (N_8282,N_8136,N_8121);
nor U8283 (N_8283,N_8158,N_8141);
or U8284 (N_8284,N_8100,N_8162);
nand U8285 (N_8285,N_8185,N_8167);
and U8286 (N_8286,N_8145,N_8189);
xor U8287 (N_8287,N_8141,N_8103);
nor U8288 (N_8288,N_8104,N_8109);
nor U8289 (N_8289,N_8126,N_8130);
or U8290 (N_8290,N_8171,N_8177);
and U8291 (N_8291,N_8178,N_8185);
or U8292 (N_8292,N_8173,N_8148);
or U8293 (N_8293,N_8103,N_8153);
nand U8294 (N_8294,N_8128,N_8161);
and U8295 (N_8295,N_8171,N_8197);
and U8296 (N_8296,N_8178,N_8100);
nand U8297 (N_8297,N_8198,N_8167);
nand U8298 (N_8298,N_8162,N_8163);
and U8299 (N_8299,N_8185,N_8173);
or U8300 (N_8300,N_8277,N_8204);
nand U8301 (N_8301,N_8263,N_8285);
or U8302 (N_8302,N_8239,N_8258);
and U8303 (N_8303,N_8216,N_8262);
nor U8304 (N_8304,N_8225,N_8281);
and U8305 (N_8305,N_8212,N_8271);
nand U8306 (N_8306,N_8266,N_8254);
xor U8307 (N_8307,N_8252,N_8221);
nor U8308 (N_8308,N_8294,N_8273);
nor U8309 (N_8309,N_8200,N_8268);
xnor U8310 (N_8310,N_8224,N_8282);
nor U8311 (N_8311,N_8207,N_8260);
or U8312 (N_8312,N_8296,N_8238);
nand U8313 (N_8313,N_8249,N_8261);
and U8314 (N_8314,N_8235,N_8203);
nand U8315 (N_8315,N_8209,N_8226);
or U8316 (N_8316,N_8217,N_8259);
and U8317 (N_8317,N_8287,N_8292);
nor U8318 (N_8318,N_8288,N_8233);
nor U8319 (N_8319,N_8295,N_8289);
nand U8320 (N_8320,N_8208,N_8243);
nand U8321 (N_8321,N_8274,N_8297);
nor U8322 (N_8322,N_8213,N_8236);
nor U8323 (N_8323,N_8284,N_8257);
or U8324 (N_8324,N_8230,N_8211);
and U8325 (N_8325,N_8286,N_8220);
or U8326 (N_8326,N_8206,N_8278);
and U8327 (N_8327,N_8223,N_8229);
and U8328 (N_8328,N_8283,N_8241);
nor U8329 (N_8329,N_8231,N_8293);
and U8330 (N_8330,N_8269,N_8215);
or U8331 (N_8331,N_8232,N_8291);
and U8332 (N_8332,N_8255,N_8227);
nor U8333 (N_8333,N_8248,N_8214);
and U8334 (N_8334,N_8251,N_8201);
nor U8335 (N_8335,N_8290,N_8299);
and U8336 (N_8336,N_8246,N_8247);
xor U8337 (N_8337,N_8219,N_8228);
xor U8338 (N_8338,N_8234,N_8202);
nor U8339 (N_8339,N_8280,N_8242);
or U8340 (N_8340,N_8256,N_8240);
nor U8341 (N_8341,N_8250,N_8205);
or U8342 (N_8342,N_8237,N_8270);
xor U8343 (N_8343,N_8264,N_8210);
nor U8344 (N_8344,N_8276,N_8298);
nand U8345 (N_8345,N_8279,N_8267);
nor U8346 (N_8346,N_8244,N_8275);
nand U8347 (N_8347,N_8265,N_8245);
and U8348 (N_8348,N_8218,N_8253);
nor U8349 (N_8349,N_8272,N_8222);
xor U8350 (N_8350,N_8262,N_8254);
nor U8351 (N_8351,N_8229,N_8204);
xor U8352 (N_8352,N_8286,N_8281);
nor U8353 (N_8353,N_8259,N_8267);
or U8354 (N_8354,N_8294,N_8229);
and U8355 (N_8355,N_8289,N_8275);
or U8356 (N_8356,N_8233,N_8249);
nand U8357 (N_8357,N_8206,N_8213);
and U8358 (N_8358,N_8295,N_8200);
or U8359 (N_8359,N_8225,N_8241);
nand U8360 (N_8360,N_8285,N_8225);
and U8361 (N_8361,N_8239,N_8268);
and U8362 (N_8362,N_8217,N_8236);
or U8363 (N_8363,N_8271,N_8286);
nor U8364 (N_8364,N_8200,N_8241);
or U8365 (N_8365,N_8278,N_8210);
nand U8366 (N_8366,N_8254,N_8241);
nor U8367 (N_8367,N_8203,N_8270);
nand U8368 (N_8368,N_8217,N_8252);
xor U8369 (N_8369,N_8274,N_8294);
nor U8370 (N_8370,N_8201,N_8219);
and U8371 (N_8371,N_8205,N_8224);
nand U8372 (N_8372,N_8238,N_8273);
nor U8373 (N_8373,N_8287,N_8260);
and U8374 (N_8374,N_8203,N_8227);
nand U8375 (N_8375,N_8218,N_8255);
xor U8376 (N_8376,N_8280,N_8260);
and U8377 (N_8377,N_8239,N_8273);
nand U8378 (N_8378,N_8237,N_8223);
nor U8379 (N_8379,N_8238,N_8247);
nor U8380 (N_8380,N_8215,N_8218);
nor U8381 (N_8381,N_8222,N_8239);
nand U8382 (N_8382,N_8211,N_8226);
nand U8383 (N_8383,N_8285,N_8222);
and U8384 (N_8384,N_8254,N_8226);
or U8385 (N_8385,N_8251,N_8218);
xor U8386 (N_8386,N_8233,N_8270);
nor U8387 (N_8387,N_8250,N_8230);
and U8388 (N_8388,N_8230,N_8238);
or U8389 (N_8389,N_8293,N_8239);
and U8390 (N_8390,N_8289,N_8262);
nand U8391 (N_8391,N_8274,N_8286);
nand U8392 (N_8392,N_8209,N_8299);
xor U8393 (N_8393,N_8297,N_8246);
or U8394 (N_8394,N_8281,N_8223);
and U8395 (N_8395,N_8213,N_8209);
or U8396 (N_8396,N_8255,N_8205);
or U8397 (N_8397,N_8220,N_8252);
nand U8398 (N_8398,N_8219,N_8260);
xnor U8399 (N_8399,N_8233,N_8225);
nand U8400 (N_8400,N_8317,N_8353);
nand U8401 (N_8401,N_8385,N_8333);
or U8402 (N_8402,N_8312,N_8373);
and U8403 (N_8403,N_8328,N_8378);
or U8404 (N_8404,N_8371,N_8319);
or U8405 (N_8405,N_8310,N_8301);
nand U8406 (N_8406,N_8341,N_8398);
nand U8407 (N_8407,N_8335,N_8379);
or U8408 (N_8408,N_8334,N_8376);
nand U8409 (N_8409,N_8387,N_8368);
xnor U8410 (N_8410,N_8304,N_8347);
nand U8411 (N_8411,N_8309,N_8336);
nand U8412 (N_8412,N_8346,N_8367);
nor U8413 (N_8413,N_8386,N_8354);
and U8414 (N_8414,N_8399,N_8369);
nand U8415 (N_8415,N_8363,N_8308);
nor U8416 (N_8416,N_8372,N_8362);
or U8417 (N_8417,N_8392,N_8396);
and U8418 (N_8418,N_8306,N_8342);
or U8419 (N_8419,N_8359,N_8381);
nand U8420 (N_8420,N_8315,N_8366);
nand U8421 (N_8421,N_8374,N_8394);
or U8422 (N_8422,N_8343,N_8357);
or U8423 (N_8423,N_8303,N_8390);
or U8424 (N_8424,N_8391,N_8300);
nor U8425 (N_8425,N_8397,N_8338);
and U8426 (N_8426,N_8344,N_8380);
and U8427 (N_8427,N_8327,N_8349);
nand U8428 (N_8428,N_8352,N_8318);
xor U8429 (N_8429,N_8360,N_8339);
nand U8430 (N_8430,N_8326,N_8377);
and U8431 (N_8431,N_8355,N_8321);
nor U8432 (N_8432,N_8337,N_8332);
and U8433 (N_8433,N_8330,N_8322);
nor U8434 (N_8434,N_8382,N_8375);
nor U8435 (N_8435,N_8351,N_8395);
nand U8436 (N_8436,N_8350,N_8370);
nand U8437 (N_8437,N_8348,N_8305);
xor U8438 (N_8438,N_8314,N_8389);
nand U8439 (N_8439,N_8302,N_8331);
or U8440 (N_8440,N_8364,N_8323);
nor U8441 (N_8441,N_8388,N_8313);
nand U8442 (N_8442,N_8384,N_8383);
or U8443 (N_8443,N_8316,N_8345);
nor U8444 (N_8444,N_8358,N_8325);
nor U8445 (N_8445,N_8365,N_8307);
nor U8446 (N_8446,N_8356,N_8393);
nor U8447 (N_8447,N_8324,N_8361);
or U8448 (N_8448,N_8320,N_8340);
or U8449 (N_8449,N_8329,N_8311);
and U8450 (N_8450,N_8388,N_8350);
nand U8451 (N_8451,N_8398,N_8374);
nor U8452 (N_8452,N_8304,N_8389);
or U8453 (N_8453,N_8346,N_8310);
nand U8454 (N_8454,N_8386,N_8341);
and U8455 (N_8455,N_8352,N_8363);
and U8456 (N_8456,N_8377,N_8336);
and U8457 (N_8457,N_8393,N_8362);
nand U8458 (N_8458,N_8318,N_8394);
nor U8459 (N_8459,N_8392,N_8327);
and U8460 (N_8460,N_8358,N_8328);
xor U8461 (N_8461,N_8308,N_8367);
nor U8462 (N_8462,N_8377,N_8379);
nand U8463 (N_8463,N_8399,N_8351);
nand U8464 (N_8464,N_8355,N_8343);
and U8465 (N_8465,N_8342,N_8353);
nor U8466 (N_8466,N_8301,N_8359);
nor U8467 (N_8467,N_8340,N_8367);
nor U8468 (N_8468,N_8335,N_8319);
nand U8469 (N_8469,N_8310,N_8378);
nand U8470 (N_8470,N_8349,N_8375);
and U8471 (N_8471,N_8377,N_8328);
and U8472 (N_8472,N_8346,N_8380);
nand U8473 (N_8473,N_8338,N_8352);
or U8474 (N_8474,N_8373,N_8322);
nor U8475 (N_8475,N_8326,N_8305);
nand U8476 (N_8476,N_8365,N_8390);
and U8477 (N_8477,N_8312,N_8332);
nor U8478 (N_8478,N_8323,N_8320);
or U8479 (N_8479,N_8300,N_8379);
and U8480 (N_8480,N_8341,N_8357);
nor U8481 (N_8481,N_8325,N_8359);
nor U8482 (N_8482,N_8333,N_8346);
nor U8483 (N_8483,N_8320,N_8378);
nor U8484 (N_8484,N_8385,N_8377);
nand U8485 (N_8485,N_8322,N_8315);
or U8486 (N_8486,N_8305,N_8317);
or U8487 (N_8487,N_8354,N_8309);
and U8488 (N_8488,N_8310,N_8389);
and U8489 (N_8489,N_8360,N_8355);
nand U8490 (N_8490,N_8361,N_8388);
xor U8491 (N_8491,N_8325,N_8354);
nor U8492 (N_8492,N_8328,N_8351);
nand U8493 (N_8493,N_8320,N_8341);
or U8494 (N_8494,N_8309,N_8303);
nand U8495 (N_8495,N_8344,N_8368);
and U8496 (N_8496,N_8332,N_8345);
and U8497 (N_8497,N_8310,N_8377);
or U8498 (N_8498,N_8372,N_8351);
nand U8499 (N_8499,N_8358,N_8345);
or U8500 (N_8500,N_8408,N_8479);
nand U8501 (N_8501,N_8476,N_8406);
nor U8502 (N_8502,N_8439,N_8488);
xor U8503 (N_8503,N_8413,N_8460);
nand U8504 (N_8504,N_8431,N_8446);
or U8505 (N_8505,N_8466,N_8418);
xnor U8506 (N_8506,N_8483,N_8477);
or U8507 (N_8507,N_8433,N_8401);
or U8508 (N_8508,N_8498,N_8443);
nor U8509 (N_8509,N_8403,N_8407);
and U8510 (N_8510,N_8404,N_8473);
or U8511 (N_8511,N_8487,N_8414);
nand U8512 (N_8512,N_8416,N_8471);
nor U8513 (N_8513,N_8475,N_8428);
nor U8514 (N_8514,N_8456,N_8490);
nand U8515 (N_8515,N_8447,N_8429);
and U8516 (N_8516,N_8400,N_8419);
nand U8517 (N_8517,N_8415,N_8409);
or U8518 (N_8518,N_8421,N_8411);
nor U8519 (N_8519,N_8458,N_8463);
or U8520 (N_8520,N_8492,N_8486);
nand U8521 (N_8521,N_8489,N_8452);
or U8522 (N_8522,N_8449,N_8465);
nor U8523 (N_8523,N_8469,N_8438);
nand U8524 (N_8524,N_8453,N_8457);
or U8525 (N_8525,N_8478,N_8410);
xnor U8526 (N_8526,N_8482,N_8420);
or U8527 (N_8527,N_8424,N_8474);
nand U8528 (N_8528,N_8450,N_8442);
nor U8529 (N_8529,N_8402,N_8491);
and U8530 (N_8530,N_8484,N_8444);
or U8531 (N_8531,N_8441,N_8472);
nor U8532 (N_8532,N_8412,N_8445);
nor U8533 (N_8533,N_8455,N_8494);
xor U8534 (N_8534,N_8481,N_8459);
nor U8535 (N_8535,N_8427,N_8499);
nand U8536 (N_8536,N_8497,N_8461);
xor U8537 (N_8537,N_8436,N_8417);
nand U8538 (N_8538,N_8454,N_8425);
and U8539 (N_8539,N_8422,N_8468);
or U8540 (N_8540,N_8496,N_8485);
nor U8541 (N_8541,N_8434,N_8448);
nor U8542 (N_8542,N_8493,N_8462);
or U8543 (N_8543,N_8426,N_8464);
or U8544 (N_8544,N_8435,N_8467);
nor U8545 (N_8545,N_8432,N_8437);
and U8546 (N_8546,N_8495,N_8423);
xnor U8547 (N_8547,N_8430,N_8405);
nor U8548 (N_8548,N_8440,N_8480);
or U8549 (N_8549,N_8451,N_8470);
nor U8550 (N_8550,N_8498,N_8432);
nand U8551 (N_8551,N_8445,N_8450);
nor U8552 (N_8552,N_8439,N_8495);
nor U8553 (N_8553,N_8470,N_8405);
nand U8554 (N_8554,N_8479,N_8420);
nor U8555 (N_8555,N_8458,N_8464);
nor U8556 (N_8556,N_8402,N_8433);
and U8557 (N_8557,N_8456,N_8463);
or U8558 (N_8558,N_8478,N_8466);
xnor U8559 (N_8559,N_8447,N_8422);
nor U8560 (N_8560,N_8494,N_8408);
and U8561 (N_8561,N_8455,N_8441);
nand U8562 (N_8562,N_8455,N_8422);
or U8563 (N_8563,N_8457,N_8456);
nor U8564 (N_8564,N_8422,N_8473);
and U8565 (N_8565,N_8477,N_8452);
nand U8566 (N_8566,N_8444,N_8423);
xor U8567 (N_8567,N_8425,N_8482);
or U8568 (N_8568,N_8474,N_8469);
or U8569 (N_8569,N_8463,N_8435);
or U8570 (N_8570,N_8448,N_8403);
or U8571 (N_8571,N_8409,N_8417);
nor U8572 (N_8572,N_8472,N_8435);
and U8573 (N_8573,N_8441,N_8480);
xor U8574 (N_8574,N_8465,N_8466);
and U8575 (N_8575,N_8438,N_8477);
xor U8576 (N_8576,N_8408,N_8495);
nor U8577 (N_8577,N_8472,N_8405);
nand U8578 (N_8578,N_8430,N_8418);
nor U8579 (N_8579,N_8466,N_8470);
nor U8580 (N_8580,N_8439,N_8497);
xnor U8581 (N_8581,N_8436,N_8463);
nand U8582 (N_8582,N_8464,N_8406);
nand U8583 (N_8583,N_8490,N_8487);
or U8584 (N_8584,N_8492,N_8467);
nor U8585 (N_8585,N_8444,N_8435);
xnor U8586 (N_8586,N_8480,N_8443);
nand U8587 (N_8587,N_8471,N_8404);
nand U8588 (N_8588,N_8422,N_8450);
or U8589 (N_8589,N_8475,N_8402);
nand U8590 (N_8590,N_8481,N_8430);
xor U8591 (N_8591,N_8469,N_8414);
xnor U8592 (N_8592,N_8467,N_8423);
and U8593 (N_8593,N_8495,N_8470);
nand U8594 (N_8594,N_8457,N_8462);
and U8595 (N_8595,N_8493,N_8427);
nor U8596 (N_8596,N_8496,N_8438);
or U8597 (N_8597,N_8430,N_8462);
nand U8598 (N_8598,N_8460,N_8443);
nand U8599 (N_8599,N_8476,N_8456);
nor U8600 (N_8600,N_8507,N_8505);
or U8601 (N_8601,N_8523,N_8516);
and U8602 (N_8602,N_8589,N_8562);
or U8603 (N_8603,N_8559,N_8577);
or U8604 (N_8604,N_8525,N_8513);
and U8605 (N_8605,N_8584,N_8595);
and U8606 (N_8606,N_8542,N_8528);
nor U8607 (N_8607,N_8566,N_8504);
nor U8608 (N_8608,N_8588,N_8544);
or U8609 (N_8609,N_8586,N_8567);
or U8610 (N_8610,N_8554,N_8565);
nor U8611 (N_8611,N_8521,N_8546);
nand U8612 (N_8612,N_8552,N_8570);
or U8613 (N_8613,N_8550,N_8534);
nor U8614 (N_8614,N_8517,N_8574);
nor U8615 (N_8615,N_8593,N_8548);
and U8616 (N_8616,N_8585,N_8560);
or U8617 (N_8617,N_8512,N_8526);
nand U8618 (N_8618,N_8580,N_8530);
or U8619 (N_8619,N_8578,N_8538);
nand U8620 (N_8620,N_8503,N_8571);
xor U8621 (N_8621,N_8532,N_8535);
xnor U8622 (N_8622,N_8572,N_8555);
nor U8623 (N_8623,N_8583,N_8519);
xnor U8624 (N_8624,N_8592,N_8539);
and U8625 (N_8625,N_8597,N_8502);
nand U8626 (N_8626,N_8582,N_8557);
nor U8627 (N_8627,N_8520,N_8596);
and U8628 (N_8628,N_8533,N_8558);
and U8629 (N_8629,N_8541,N_8551);
and U8630 (N_8630,N_8587,N_8514);
or U8631 (N_8631,N_8594,N_8515);
and U8632 (N_8632,N_8527,N_8561);
or U8633 (N_8633,N_8553,N_8511);
nor U8634 (N_8634,N_8575,N_8518);
and U8635 (N_8635,N_8537,N_8508);
and U8636 (N_8636,N_8599,N_8573);
or U8637 (N_8637,N_8506,N_8524);
or U8638 (N_8638,N_8543,N_8531);
xor U8639 (N_8639,N_8509,N_8556);
nand U8640 (N_8640,N_8563,N_8576);
or U8641 (N_8641,N_8501,N_8568);
nand U8642 (N_8642,N_8549,N_8598);
nor U8643 (N_8643,N_8536,N_8545);
nor U8644 (N_8644,N_8581,N_8529);
nor U8645 (N_8645,N_8540,N_8590);
or U8646 (N_8646,N_8522,N_8547);
and U8647 (N_8647,N_8579,N_8510);
nand U8648 (N_8648,N_8564,N_8591);
nand U8649 (N_8649,N_8569,N_8500);
nand U8650 (N_8650,N_8514,N_8576);
and U8651 (N_8651,N_8518,N_8550);
nand U8652 (N_8652,N_8598,N_8501);
or U8653 (N_8653,N_8586,N_8549);
and U8654 (N_8654,N_8535,N_8548);
or U8655 (N_8655,N_8550,N_8508);
nand U8656 (N_8656,N_8577,N_8528);
nor U8657 (N_8657,N_8596,N_8524);
and U8658 (N_8658,N_8593,N_8523);
nand U8659 (N_8659,N_8516,N_8599);
nand U8660 (N_8660,N_8559,N_8573);
nor U8661 (N_8661,N_8539,N_8545);
nor U8662 (N_8662,N_8542,N_8508);
xor U8663 (N_8663,N_8504,N_8597);
or U8664 (N_8664,N_8577,N_8590);
and U8665 (N_8665,N_8582,N_8501);
nor U8666 (N_8666,N_8505,N_8516);
or U8667 (N_8667,N_8522,N_8554);
nand U8668 (N_8668,N_8546,N_8579);
xnor U8669 (N_8669,N_8533,N_8537);
and U8670 (N_8670,N_8500,N_8570);
nor U8671 (N_8671,N_8533,N_8539);
nor U8672 (N_8672,N_8511,N_8544);
nor U8673 (N_8673,N_8542,N_8592);
or U8674 (N_8674,N_8522,N_8519);
and U8675 (N_8675,N_8551,N_8547);
or U8676 (N_8676,N_8562,N_8550);
and U8677 (N_8677,N_8599,N_8500);
xnor U8678 (N_8678,N_8511,N_8516);
nand U8679 (N_8679,N_8587,N_8504);
or U8680 (N_8680,N_8571,N_8520);
nor U8681 (N_8681,N_8586,N_8533);
or U8682 (N_8682,N_8583,N_8542);
nor U8683 (N_8683,N_8549,N_8581);
and U8684 (N_8684,N_8594,N_8556);
nor U8685 (N_8685,N_8536,N_8520);
nand U8686 (N_8686,N_8584,N_8509);
nand U8687 (N_8687,N_8507,N_8588);
nand U8688 (N_8688,N_8579,N_8561);
or U8689 (N_8689,N_8559,N_8520);
or U8690 (N_8690,N_8560,N_8565);
and U8691 (N_8691,N_8541,N_8540);
nand U8692 (N_8692,N_8546,N_8537);
and U8693 (N_8693,N_8562,N_8503);
and U8694 (N_8694,N_8554,N_8572);
nor U8695 (N_8695,N_8572,N_8576);
and U8696 (N_8696,N_8597,N_8582);
and U8697 (N_8697,N_8580,N_8557);
xor U8698 (N_8698,N_8507,N_8574);
or U8699 (N_8699,N_8573,N_8547);
nand U8700 (N_8700,N_8609,N_8619);
nand U8701 (N_8701,N_8673,N_8694);
or U8702 (N_8702,N_8693,N_8652);
xnor U8703 (N_8703,N_8607,N_8674);
or U8704 (N_8704,N_8698,N_8684);
and U8705 (N_8705,N_8632,N_8608);
or U8706 (N_8706,N_8627,N_8653);
nor U8707 (N_8707,N_8624,N_8649);
and U8708 (N_8708,N_8683,N_8645);
or U8709 (N_8709,N_8614,N_8602);
nor U8710 (N_8710,N_8618,N_8644);
and U8711 (N_8711,N_8696,N_8676);
nand U8712 (N_8712,N_8695,N_8677);
nor U8713 (N_8713,N_8662,N_8605);
nor U8714 (N_8714,N_8625,N_8699);
or U8715 (N_8715,N_8640,N_8621);
or U8716 (N_8716,N_8642,N_8689);
or U8717 (N_8717,N_8616,N_8692);
nor U8718 (N_8718,N_8650,N_8641);
nor U8719 (N_8719,N_8613,N_8623);
and U8720 (N_8720,N_8668,N_8667);
and U8721 (N_8721,N_8680,N_8620);
or U8722 (N_8722,N_8659,N_8665);
and U8723 (N_8723,N_8671,N_8626);
and U8724 (N_8724,N_8681,N_8691);
nor U8725 (N_8725,N_8688,N_8697);
and U8726 (N_8726,N_8651,N_8685);
and U8727 (N_8727,N_8628,N_8647);
or U8728 (N_8728,N_8646,N_8638);
or U8729 (N_8729,N_8656,N_8630);
xor U8730 (N_8730,N_8636,N_8666);
nor U8731 (N_8731,N_8615,N_8655);
nand U8732 (N_8732,N_8690,N_8678);
nand U8733 (N_8733,N_8629,N_8675);
or U8734 (N_8734,N_8648,N_8631);
or U8735 (N_8735,N_8617,N_8679);
xnor U8736 (N_8736,N_8612,N_8634);
or U8737 (N_8737,N_8686,N_8663);
nor U8738 (N_8738,N_8606,N_8643);
and U8739 (N_8739,N_8657,N_8622);
xnor U8740 (N_8740,N_8672,N_8682);
and U8741 (N_8741,N_8603,N_8600);
or U8742 (N_8742,N_8601,N_8604);
nand U8743 (N_8743,N_8661,N_8637);
nor U8744 (N_8744,N_8639,N_8635);
nand U8745 (N_8745,N_8669,N_8660);
nand U8746 (N_8746,N_8658,N_8670);
and U8747 (N_8747,N_8654,N_8664);
or U8748 (N_8748,N_8687,N_8633);
nor U8749 (N_8749,N_8610,N_8611);
nor U8750 (N_8750,N_8693,N_8656);
or U8751 (N_8751,N_8637,N_8616);
nor U8752 (N_8752,N_8656,N_8632);
and U8753 (N_8753,N_8604,N_8690);
nand U8754 (N_8754,N_8642,N_8658);
nand U8755 (N_8755,N_8656,N_8622);
and U8756 (N_8756,N_8651,N_8666);
and U8757 (N_8757,N_8650,N_8676);
and U8758 (N_8758,N_8684,N_8651);
or U8759 (N_8759,N_8682,N_8608);
and U8760 (N_8760,N_8648,N_8697);
nand U8761 (N_8761,N_8664,N_8689);
nor U8762 (N_8762,N_8652,N_8683);
and U8763 (N_8763,N_8624,N_8614);
or U8764 (N_8764,N_8638,N_8685);
xnor U8765 (N_8765,N_8691,N_8693);
xor U8766 (N_8766,N_8615,N_8613);
nand U8767 (N_8767,N_8655,N_8601);
and U8768 (N_8768,N_8671,N_8606);
nor U8769 (N_8769,N_8697,N_8665);
nand U8770 (N_8770,N_8657,N_8669);
nand U8771 (N_8771,N_8656,N_8664);
nand U8772 (N_8772,N_8656,N_8667);
nand U8773 (N_8773,N_8657,N_8650);
or U8774 (N_8774,N_8692,N_8613);
or U8775 (N_8775,N_8693,N_8667);
nand U8776 (N_8776,N_8659,N_8678);
nor U8777 (N_8777,N_8668,N_8627);
nor U8778 (N_8778,N_8680,N_8612);
nand U8779 (N_8779,N_8634,N_8681);
nor U8780 (N_8780,N_8643,N_8650);
nor U8781 (N_8781,N_8680,N_8625);
or U8782 (N_8782,N_8699,N_8655);
or U8783 (N_8783,N_8666,N_8687);
nor U8784 (N_8784,N_8627,N_8649);
nor U8785 (N_8785,N_8693,N_8681);
and U8786 (N_8786,N_8676,N_8659);
xnor U8787 (N_8787,N_8619,N_8661);
xor U8788 (N_8788,N_8698,N_8638);
nand U8789 (N_8789,N_8644,N_8691);
or U8790 (N_8790,N_8606,N_8636);
xor U8791 (N_8791,N_8691,N_8636);
and U8792 (N_8792,N_8676,N_8663);
nor U8793 (N_8793,N_8692,N_8673);
or U8794 (N_8794,N_8692,N_8624);
and U8795 (N_8795,N_8693,N_8607);
nand U8796 (N_8796,N_8647,N_8633);
nor U8797 (N_8797,N_8654,N_8676);
nor U8798 (N_8798,N_8609,N_8627);
nand U8799 (N_8799,N_8658,N_8606);
nor U8800 (N_8800,N_8712,N_8754);
nand U8801 (N_8801,N_8781,N_8723);
or U8802 (N_8802,N_8762,N_8725);
and U8803 (N_8803,N_8748,N_8789);
or U8804 (N_8804,N_8740,N_8744);
and U8805 (N_8805,N_8757,N_8791);
nand U8806 (N_8806,N_8749,N_8769);
nand U8807 (N_8807,N_8731,N_8750);
or U8808 (N_8808,N_8732,N_8768);
xnor U8809 (N_8809,N_8772,N_8738);
or U8810 (N_8810,N_8759,N_8739);
or U8811 (N_8811,N_8798,N_8776);
nand U8812 (N_8812,N_8786,N_8733);
nor U8813 (N_8813,N_8752,N_8718);
xnor U8814 (N_8814,N_8792,N_8705);
or U8815 (N_8815,N_8796,N_8726);
xor U8816 (N_8816,N_8760,N_8734);
and U8817 (N_8817,N_8766,N_8799);
and U8818 (N_8818,N_8746,N_8719);
and U8819 (N_8819,N_8797,N_8735);
nand U8820 (N_8820,N_8706,N_8721);
or U8821 (N_8821,N_8702,N_8761);
nor U8822 (N_8822,N_8770,N_8724);
or U8823 (N_8823,N_8704,N_8755);
or U8824 (N_8824,N_8714,N_8728);
or U8825 (N_8825,N_8707,N_8747);
and U8826 (N_8826,N_8773,N_8742);
nand U8827 (N_8827,N_8758,N_8785);
and U8828 (N_8828,N_8756,N_8763);
nand U8829 (N_8829,N_8775,N_8765);
xor U8830 (N_8830,N_8701,N_8743);
or U8831 (N_8831,N_8793,N_8795);
nand U8832 (N_8832,N_8787,N_8778);
or U8833 (N_8833,N_8794,N_8703);
or U8834 (N_8834,N_8751,N_8709);
nor U8835 (N_8835,N_8716,N_8717);
and U8836 (N_8836,N_8777,N_8782);
nand U8837 (N_8837,N_8730,N_8783);
xnor U8838 (N_8838,N_8764,N_8710);
or U8839 (N_8839,N_8720,N_8779);
or U8840 (N_8840,N_8780,N_8745);
and U8841 (N_8841,N_8713,N_8790);
nand U8842 (N_8842,N_8729,N_8727);
nand U8843 (N_8843,N_8736,N_8711);
xor U8844 (N_8844,N_8737,N_8708);
and U8845 (N_8845,N_8753,N_8788);
and U8846 (N_8846,N_8700,N_8767);
and U8847 (N_8847,N_8715,N_8722);
nand U8848 (N_8848,N_8774,N_8784);
nand U8849 (N_8849,N_8741,N_8771);
or U8850 (N_8850,N_8722,N_8736);
nand U8851 (N_8851,N_8721,N_8700);
nand U8852 (N_8852,N_8771,N_8778);
nand U8853 (N_8853,N_8718,N_8781);
nand U8854 (N_8854,N_8729,N_8717);
nor U8855 (N_8855,N_8796,N_8792);
and U8856 (N_8856,N_8791,N_8744);
and U8857 (N_8857,N_8711,N_8763);
or U8858 (N_8858,N_8784,N_8708);
xor U8859 (N_8859,N_8745,N_8759);
or U8860 (N_8860,N_8703,N_8753);
or U8861 (N_8861,N_8716,N_8762);
nor U8862 (N_8862,N_8700,N_8793);
nand U8863 (N_8863,N_8788,N_8776);
nor U8864 (N_8864,N_8744,N_8765);
or U8865 (N_8865,N_8752,N_8730);
and U8866 (N_8866,N_8755,N_8718);
nor U8867 (N_8867,N_8746,N_8713);
or U8868 (N_8868,N_8727,N_8739);
xnor U8869 (N_8869,N_8791,N_8741);
and U8870 (N_8870,N_8724,N_8799);
nand U8871 (N_8871,N_8706,N_8797);
xnor U8872 (N_8872,N_8774,N_8741);
nand U8873 (N_8873,N_8796,N_8798);
nand U8874 (N_8874,N_8700,N_8710);
nor U8875 (N_8875,N_8769,N_8714);
and U8876 (N_8876,N_8710,N_8776);
and U8877 (N_8877,N_8716,N_8725);
and U8878 (N_8878,N_8740,N_8747);
or U8879 (N_8879,N_8718,N_8746);
nand U8880 (N_8880,N_8745,N_8719);
and U8881 (N_8881,N_8771,N_8722);
nand U8882 (N_8882,N_8736,N_8752);
nor U8883 (N_8883,N_8746,N_8734);
or U8884 (N_8884,N_8719,N_8794);
nor U8885 (N_8885,N_8716,N_8777);
or U8886 (N_8886,N_8705,N_8702);
nand U8887 (N_8887,N_8715,N_8702);
and U8888 (N_8888,N_8701,N_8775);
nand U8889 (N_8889,N_8778,N_8790);
or U8890 (N_8890,N_8742,N_8730);
nor U8891 (N_8891,N_8785,N_8767);
nor U8892 (N_8892,N_8744,N_8795);
and U8893 (N_8893,N_8716,N_8769);
or U8894 (N_8894,N_8739,N_8737);
nor U8895 (N_8895,N_8756,N_8760);
or U8896 (N_8896,N_8700,N_8709);
nor U8897 (N_8897,N_8750,N_8752);
nor U8898 (N_8898,N_8739,N_8712);
and U8899 (N_8899,N_8752,N_8755);
xnor U8900 (N_8900,N_8850,N_8854);
xor U8901 (N_8901,N_8883,N_8869);
or U8902 (N_8902,N_8868,N_8820);
and U8903 (N_8903,N_8802,N_8871);
or U8904 (N_8904,N_8882,N_8898);
and U8905 (N_8905,N_8848,N_8817);
and U8906 (N_8906,N_8856,N_8897);
and U8907 (N_8907,N_8877,N_8865);
xnor U8908 (N_8908,N_8857,N_8805);
or U8909 (N_8909,N_8821,N_8888);
or U8910 (N_8910,N_8803,N_8880);
nor U8911 (N_8911,N_8872,N_8870);
and U8912 (N_8912,N_8825,N_8841);
xor U8913 (N_8913,N_8845,N_8875);
or U8914 (N_8914,N_8840,N_8851);
or U8915 (N_8915,N_8829,N_8858);
nor U8916 (N_8916,N_8835,N_8801);
nor U8917 (N_8917,N_8836,N_8812);
nor U8918 (N_8918,N_8859,N_8837);
nor U8919 (N_8919,N_8804,N_8814);
nand U8920 (N_8920,N_8893,N_8862);
nand U8921 (N_8921,N_8896,N_8800);
or U8922 (N_8922,N_8892,N_8842);
or U8923 (N_8923,N_8806,N_8826);
nor U8924 (N_8924,N_8866,N_8843);
nor U8925 (N_8925,N_8890,N_8822);
nand U8926 (N_8926,N_8807,N_8824);
and U8927 (N_8927,N_8846,N_8816);
nand U8928 (N_8928,N_8878,N_8852);
nor U8929 (N_8929,N_8809,N_8874);
nand U8930 (N_8930,N_8876,N_8864);
or U8931 (N_8931,N_8833,N_8844);
nor U8932 (N_8932,N_8831,N_8873);
and U8933 (N_8933,N_8863,N_8834);
nor U8934 (N_8934,N_8855,N_8815);
nand U8935 (N_8935,N_8887,N_8811);
nand U8936 (N_8936,N_8853,N_8860);
nor U8937 (N_8937,N_8891,N_8832);
nor U8938 (N_8938,N_8894,N_8889);
nand U8939 (N_8939,N_8810,N_8867);
or U8940 (N_8940,N_8895,N_8827);
or U8941 (N_8941,N_8884,N_8879);
and U8942 (N_8942,N_8828,N_8861);
xnor U8943 (N_8943,N_8830,N_8847);
nand U8944 (N_8944,N_8808,N_8839);
nand U8945 (N_8945,N_8813,N_8838);
nand U8946 (N_8946,N_8823,N_8819);
or U8947 (N_8947,N_8881,N_8885);
nor U8948 (N_8948,N_8886,N_8899);
or U8949 (N_8949,N_8849,N_8818);
or U8950 (N_8950,N_8856,N_8808);
and U8951 (N_8951,N_8899,N_8859);
xnor U8952 (N_8952,N_8821,N_8830);
nand U8953 (N_8953,N_8886,N_8803);
or U8954 (N_8954,N_8846,N_8890);
xnor U8955 (N_8955,N_8805,N_8860);
and U8956 (N_8956,N_8832,N_8898);
nor U8957 (N_8957,N_8842,N_8872);
nor U8958 (N_8958,N_8817,N_8838);
nor U8959 (N_8959,N_8813,N_8817);
xnor U8960 (N_8960,N_8845,N_8892);
nor U8961 (N_8961,N_8894,N_8882);
nand U8962 (N_8962,N_8818,N_8805);
nand U8963 (N_8963,N_8842,N_8802);
nor U8964 (N_8964,N_8837,N_8861);
or U8965 (N_8965,N_8829,N_8814);
nor U8966 (N_8966,N_8860,N_8892);
nor U8967 (N_8967,N_8818,N_8828);
or U8968 (N_8968,N_8806,N_8888);
nor U8969 (N_8969,N_8809,N_8871);
nor U8970 (N_8970,N_8829,N_8864);
nand U8971 (N_8971,N_8897,N_8817);
nand U8972 (N_8972,N_8853,N_8844);
nand U8973 (N_8973,N_8806,N_8865);
xor U8974 (N_8974,N_8866,N_8803);
and U8975 (N_8975,N_8889,N_8875);
nor U8976 (N_8976,N_8895,N_8882);
and U8977 (N_8977,N_8893,N_8877);
and U8978 (N_8978,N_8804,N_8829);
nor U8979 (N_8979,N_8897,N_8866);
or U8980 (N_8980,N_8875,N_8804);
or U8981 (N_8981,N_8887,N_8856);
nor U8982 (N_8982,N_8853,N_8863);
nand U8983 (N_8983,N_8894,N_8855);
nand U8984 (N_8984,N_8816,N_8879);
nand U8985 (N_8985,N_8865,N_8856);
xor U8986 (N_8986,N_8864,N_8842);
or U8987 (N_8987,N_8838,N_8844);
nor U8988 (N_8988,N_8808,N_8879);
and U8989 (N_8989,N_8849,N_8874);
and U8990 (N_8990,N_8841,N_8879);
xnor U8991 (N_8991,N_8818,N_8809);
nor U8992 (N_8992,N_8863,N_8884);
nor U8993 (N_8993,N_8825,N_8808);
and U8994 (N_8994,N_8895,N_8800);
nor U8995 (N_8995,N_8813,N_8883);
or U8996 (N_8996,N_8865,N_8848);
or U8997 (N_8997,N_8866,N_8830);
and U8998 (N_8998,N_8834,N_8864);
and U8999 (N_8999,N_8802,N_8832);
nor U9000 (N_9000,N_8966,N_8977);
or U9001 (N_9001,N_8997,N_8924);
nand U9002 (N_9002,N_8945,N_8993);
xnor U9003 (N_9003,N_8959,N_8961);
xor U9004 (N_9004,N_8971,N_8917);
or U9005 (N_9005,N_8952,N_8919);
and U9006 (N_9006,N_8975,N_8903);
or U9007 (N_9007,N_8943,N_8928);
or U9008 (N_9008,N_8989,N_8969);
or U9009 (N_9009,N_8956,N_8921);
and U9010 (N_9010,N_8932,N_8916);
and U9011 (N_9011,N_8996,N_8988);
nor U9012 (N_9012,N_8976,N_8990);
nor U9013 (N_9013,N_8974,N_8980);
nor U9014 (N_9014,N_8962,N_8950);
or U9015 (N_9015,N_8930,N_8955);
nand U9016 (N_9016,N_8948,N_8922);
and U9017 (N_9017,N_8991,N_8939);
or U9018 (N_9018,N_8934,N_8926);
nand U9019 (N_9019,N_8909,N_8904);
or U9020 (N_9020,N_8958,N_8901);
nand U9021 (N_9021,N_8981,N_8914);
nand U9022 (N_9022,N_8972,N_8960);
nor U9023 (N_9023,N_8946,N_8963);
or U9024 (N_9024,N_8949,N_8998);
nand U9025 (N_9025,N_8927,N_8982);
or U9026 (N_9026,N_8992,N_8923);
nor U9027 (N_9027,N_8994,N_8929);
or U9028 (N_9028,N_8940,N_8957);
or U9029 (N_9029,N_8985,N_8906);
and U9030 (N_9030,N_8905,N_8900);
xor U9031 (N_9031,N_8995,N_8984);
nor U9032 (N_9032,N_8913,N_8983);
xnor U9033 (N_9033,N_8936,N_8908);
and U9034 (N_9034,N_8967,N_8915);
and U9035 (N_9035,N_8964,N_8951);
nand U9036 (N_9036,N_8907,N_8954);
nand U9037 (N_9037,N_8942,N_8947);
or U9038 (N_9038,N_8935,N_8973);
nand U9039 (N_9039,N_8999,N_8938);
or U9040 (N_9040,N_8902,N_8968);
or U9041 (N_9041,N_8925,N_8953);
and U9042 (N_9042,N_8970,N_8912);
or U9043 (N_9043,N_8911,N_8920);
and U9044 (N_9044,N_8978,N_8979);
or U9045 (N_9045,N_8965,N_8986);
or U9046 (N_9046,N_8910,N_8987);
nor U9047 (N_9047,N_8933,N_8931);
xnor U9048 (N_9048,N_8944,N_8941);
nor U9049 (N_9049,N_8937,N_8918);
or U9050 (N_9050,N_8964,N_8950);
and U9051 (N_9051,N_8906,N_8912);
nand U9052 (N_9052,N_8968,N_8990);
nor U9053 (N_9053,N_8938,N_8926);
nor U9054 (N_9054,N_8985,N_8980);
and U9055 (N_9055,N_8902,N_8901);
xnor U9056 (N_9056,N_8919,N_8911);
nor U9057 (N_9057,N_8927,N_8957);
or U9058 (N_9058,N_8913,N_8968);
and U9059 (N_9059,N_8914,N_8903);
nand U9060 (N_9060,N_8995,N_8976);
and U9061 (N_9061,N_8956,N_8910);
or U9062 (N_9062,N_8976,N_8900);
nand U9063 (N_9063,N_8989,N_8971);
nor U9064 (N_9064,N_8918,N_8926);
xor U9065 (N_9065,N_8960,N_8940);
nand U9066 (N_9066,N_8939,N_8994);
or U9067 (N_9067,N_8901,N_8988);
or U9068 (N_9068,N_8928,N_8900);
nor U9069 (N_9069,N_8995,N_8917);
or U9070 (N_9070,N_8933,N_8934);
nor U9071 (N_9071,N_8974,N_8909);
xor U9072 (N_9072,N_8966,N_8983);
nand U9073 (N_9073,N_8901,N_8973);
nand U9074 (N_9074,N_8971,N_8969);
nor U9075 (N_9075,N_8902,N_8947);
and U9076 (N_9076,N_8954,N_8959);
nand U9077 (N_9077,N_8930,N_8959);
and U9078 (N_9078,N_8999,N_8977);
nor U9079 (N_9079,N_8947,N_8989);
nor U9080 (N_9080,N_8983,N_8954);
nand U9081 (N_9081,N_8910,N_8948);
and U9082 (N_9082,N_8936,N_8911);
xnor U9083 (N_9083,N_8952,N_8913);
nor U9084 (N_9084,N_8940,N_8988);
and U9085 (N_9085,N_8920,N_8960);
xnor U9086 (N_9086,N_8900,N_8964);
xnor U9087 (N_9087,N_8982,N_8910);
nand U9088 (N_9088,N_8909,N_8963);
nor U9089 (N_9089,N_8978,N_8921);
and U9090 (N_9090,N_8942,N_8939);
nand U9091 (N_9091,N_8976,N_8973);
nor U9092 (N_9092,N_8925,N_8999);
and U9093 (N_9093,N_8915,N_8951);
or U9094 (N_9094,N_8934,N_8968);
nand U9095 (N_9095,N_8927,N_8977);
nor U9096 (N_9096,N_8929,N_8998);
and U9097 (N_9097,N_8995,N_8921);
and U9098 (N_9098,N_8999,N_8933);
and U9099 (N_9099,N_8906,N_8999);
nand U9100 (N_9100,N_9005,N_9055);
nor U9101 (N_9101,N_9058,N_9049);
nand U9102 (N_9102,N_9003,N_9008);
nor U9103 (N_9103,N_9044,N_9098);
or U9104 (N_9104,N_9024,N_9015);
or U9105 (N_9105,N_9086,N_9038);
and U9106 (N_9106,N_9083,N_9050);
nand U9107 (N_9107,N_9062,N_9029);
nand U9108 (N_9108,N_9060,N_9052);
nor U9109 (N_9109,N_9017,N_9028);
nor U9110 (N_9110,N_9064,N_9018);
nor U9111 (N_9111,N_9075,N_9041);
nor U9112 (N_9112,N_9074,N_9000);
and U9113 (N_9113,N_9016,N_9011);
nor U9114 (N_9114,N_9070,N_9037);
nor U9115 (N_9115,N_9097,N_9022);
nor U9116 (N_9116,N_9095,N_9099);
or U9117 (N_9117,N_9032,N_9033);
nor U9118 (N_9118,N_9012,N_9019);
nor U9119 (N_9119,N_9063,N_9035);
and U9120 (N_9120,N_9056,N_9010);
xnor U9121 (N_9121,N_9089,N_9026);
xnor U9122 (N_9122,N_9096,N_9094);
xnor U9123 (N_9123,N_9001,N_9068);
xnor U9124 (N_9124,N_9043,N_9087);
nor U9125 (N_9125,N_9045,N_9013);
nand U9126 (N_9126,N_9080,N_9078);
and U9127 (N_9127,N_9067,N_9002);
nand U9128 (N_9128,N_9091,N_9027);
xor U9129 (N_9129,N_9007,N_9066);
nor U9130 (N_9130,N_9042,N_9065);
nand U9131 (N_9131,N_9093,N_9034);
nand U9132 (N_9132,N_9054,N_9006);
nand U9133 (N_9133,N_9076,N_9077);
and U9134 (N_9134,N_9009,N_9031);
and U9135 (N_9135,N_9021,N_9048);
and U9136 (N_9136,N_9040,N_9073);
nor U9137 (N_9137,N_9039,N_9082);
or U9138 (N_9138,N_9069,N_9081);
nand U9139 (N_9139,N_9036,N_9071);
nand U9140 (N_9140,N_9023,N_9079);
or U9141 (N_9141,N_9084,N_9061);
or U9142 (N_9142,N_9046,N_9030);
and U9143 (N_9143,N_9057,N_9014);
xnor U9144 (N_9144,N_9051,N_9004);
or U9145 (N_9145,N_9020,N_9053);
xor U9146 (N_9146,N_9088,N_9047);
and U9147 (N_9147,N_9072,N_9090);
and U9148 (N_9148,N_9025,N_9085);
or U9149 (N_9149,N_9092,N_9059);
nor U9150 (N_9150,N_9038,N_9045);
and U9151 (N_9151,N_9090,N_9084);
or U9152 (N_9152,N_9087,N_9003);
or U9153 (N_9153,N_9087,N_9066);
or U9154 (N_9154,N_9067,N_9055);
or U9155 (N_9155,N_9056,N_9097);
nand U9156 (N_9156,N_9050,N_9051);
nand U9157 (N_9157,N_9061,N_9016);
or U9158 (N_9158,N_9007,N_9009);
or U9159 (N_9159,N_9041,N_9022);
or U9160 (N_9160,N_9076,N_9072);
and U9161 (N_9161,N_9007,N_9008);
and U9162 (N_9162,N_9027,N_9044);
and U9163 (N_9163,N_9061,N_9017);
nand U9164 (N_9164,N_9074,N_9011);
or U9165 (N_9165,N_9072,N_9018);
or U9166 (N_9166,N_9021,N_9054);
nor U9167 (N_9167,N_9053,N_9012);
nand U9168 (N_9168,N_9024,N_9060);
xnor U9169 (N_9169,N_9034,N_9032);
nor U9170 (N_9170,N_9084,N_9060);
or U9171 (N_9171,N_9016,N_9075);
xnor U9172 (N_9172,N_9078,N_9053);
or U9173 (N_9173,N_9056,N_9025);
and U9174 (N_9174,N_9040,N_9089);
and U9175 (N_9175,N_9039,N_9036);
nand U9176 (N_9176,N_9014,N_9046);
nor U9177 (N_9177,N_9080,N_9075);
or U9178 (N_9178,N_9087,N_9025);
nor U9179 (N_9179,N_9060,N_9078);
nor U9180 (N_9180,N_9076,N_9000);
xnor U9181 (N_9181,N_9013,N_9049);
nor U9182 (N_9182,N_9084,N_9062);
or U9183 (N_9183,N_9094,N_9047);
xor U9184 (N_9184,N_9012,N_9075);
xnor U9185 (N_9185,N_9010,N_9045);
and U9186 (N_9186,N_9037,N_9027);
nor U9187 (N_9187,N_9053,N_9035);
nand U9188 (N_9188,N_9054,N_9041);
nor U9189 (N_9189,N_9048,N_9076);
or U9190 (N_9190,N_9014,N_9018);
nor U9191 (N_9191,N_9086,N_9029);
xnor U9192 (N_9192,N_9079,N_9065);
xnor U9193 (N_9193,N_9035,N_9066);
nand U9194 (N_9194,N_9014,N_9035);
xnor U9195 (N_9195,N_9046,N_9090);
and U9196 (N_9196,N_9063,N_9033);
and U9197 (N_9197,N_9099,N_9018);
nand U9198 (N_9198,N_9004,N_9045);
or U9199 (N_9199,N_9090,N_9088);
nor U9200 (N_9200,N_9165,N_9168);
and U9201 (N_9201,N_9146,N_9145);
and U9202 (N_9202,N_9171,N_9106);
and U9203 (N_9203,N_9152,N_9100);
nand U9204 (N_9204,N_9191,N_9195);
nor U9205 (N_9205,N_9179,N_9154);
and U9206 (N_9206,N_9124,N_9161);
nand U9207 (N_9207,N_9164,N_9134);
nand U9208 (N_9208,N_9169,N_9196);
nor U9209 (N_9209,N_9199,N_9144);
nor U9210 (N_9210,N_9116,N_9198);
and U9211 (N_9211,N_9132,N_9177);
or U9212 (N_9212,N_9193,N_9121);
nor U9213 (N_9213,N_9194,N_9107);
and U9214 (N_9214,N_9162,N_9141);
nor U9215 (N_9215,N_9182,N_9136);
and U9216 (N_9216,N_9142,N_9147);
nor U9217 (N_9217,N_9175,N_9111);
xnor U9218 (N_9218,N_9176,N_9186);
xor U9219 (N_9219,N_9188,N_9155);
nand U9220 (N_9220,N_9131,N_9158);
xor U9221 (N_9221,N_9189,N_9197);
nand U9222 (N_9222,N_9117,N_9187);
and U9223 (N_9223,N_9173,N_9150);
nor U9224 (N_9224,N_9122,N_9153);
and U9225 (N_9225,N_9119,N_9115);
xor U9226 (N_9226,N_9178,N_9105);
nand U9227 (N_9227,N_9112,N_9167);
nand U9228 (N_9228,N_9140,N_9125);
nand U9229 (N_9229,N_9137,N_9166);
or U9230 (N_9230,N_9183,N_9118);
and U9231 (N_9231,N_9128,N_9163);
or U9232 (N_9232,N_9110,N_9103);
and U9233 (N_9233,N_9181,N_9129);
nor U9234 (N_9234,N_9192,N_9139);
nor U9235 (N_9235,N_9104,N_9185);
nand U9236 (N_9236,N_9114,N_9109);
nor U9237 (N_9237,N_9123,N_9148);
or U9238 (N_9238,N_9160,N_9108);
nand U9239 (N_9239,N_9151,N_9159);
xnor U9240 (N_9240,N_9127,N_9157);
nor U9241 (N_9241,N_9156,N_9170);
or U9242 (N_9242,N_9180,N_9138);
and U9243 (N_9243,N_9149,N_9190);
and U9244 (N_9244,N_9102,N_9120);
nand U9245 (N_9245,N_9143,N_9113);
and U9246 (N_9246,N_9101,N_9184);
xor U9247 (N_9247,N_9135,N_9133);
and U9248 (N_9248,N_9172,N_9174);
xor U9249 (N_9249,N_9126,N_9130);
or U9250 (N_9250,N_9187,N_9155);
or U9251 (N_9251,N_9116,N_9112);
nor U9252 (N_9252,N_9155,N_9100);
xor U9253 (N_9253,N_9186,N_9154);
nand U9254 (N_9254,N_9186,N_9158);
or U9255 (N_9255,N_9183,N_9190);
and U9256 (N_9256,N_9184,N_9104);
or U9257 (N_9257,N_9177,N_9198);
nor U9258 (N_9258,N_9136,N_9166);
nor U9259 (N_9259,N_9109,N_9125);
nor U9260 (N_9260,N_9145,N_9179);
nand U9261 (N_9261,N_9185,N_9189);
nand U9262 (N_9262,N_9142,N_9160);
nor U9263 (N_9263,N_9123,N_9139);
nor U9264 (N_9264,N_9157,N_9191);
or U9265 (N_9265,N_9149,N_9133);
or U9266 (N_9266,N_9119,N_9104);
or U9267 (N_9267,N_9170,N_9148);
xor U9268 (N_9268,N_9109,N_9124);
nand U9269 (N_9269,N_9157,N_9118);
xnor U9270 (N_9270,N_9113,N_9172);
nor U9271 (N_9271,N_9179,N_9133);
nand U9272 (N_9272,N_9104,N_9128);
nor U9273 (N_9273,N_9166,N_9199);
and U9274 (N_9274,N_9157,N_9132);
nor U9275 (N_9275,N_9104,N_9161);
nor U9276 (N_9276,N_9131,N_9168);
nand U9277 (N_9277,N_9198,N_9118);
and U9278 (N_9278,N_9185,N_9138);
nor U9279 (N_9279,N_9120,N_9165);
nor U9280 (N_9280,N_9162,N_9122);
nand U9281 (N_9281,N_9123,N_9182);
and U9282 (N_9282,N_9151,N_9170);
xnor U9283 (N_9283,N_9113,N_9149);
or U9284 (N_9284,N_9185,N_9182);
nand U9285 (N_9285,N_9189,N_9199);
or U9286 (N_9286,N_9112,N_9191);
nand U9287 (N_9287,N_9122,N_9172);
nor U9288 (N_9288,N_9113,N_9131);
nand U9289 (N_9289,N_9166,N_9177);
and U9290 (N_9290,N_9119,N_9138);
nor U9291 (N_9291,N_9134,N_9153);
xnor U9292 (N_9292,N_9166,N_9169);
nor U9293 (N_9293,N_9120,N_9121);
and U9294 (N_9294,N_9153,N_9151);
nor U9295 (N_9295,N_9154,N_9122);
nand U9296 (N_9296,N_9151,N_9155);
and U9297 (N_9297,N_9110,N_9145);
and U9298 (N_9298,N_9132,N_9143);
nor U9299 (N_9299,N_9157,N_9159);
nor U9300 (N_9300,N_9285,N_9255);
nor U9301 (N_9301,N_9249,N_9286);
nand U9302 (N_9302,N_9297,N_9295);
and U9303 (N_9303,N_9204,N_9281);
nand U9304 (N_9304,N_9214,N_9226);
and U9305 (N_9305,N_9202,N_9237);
nor U9306 (N_9306,N_9240,N_9293);
nand U9307 (N_9307,N_9222,N_9201);
and U9308 (N_9308,N_9218,N_9270);
xor U9309 (N_9309,N_9275,N_9200);
or U9310 (N_9310,N_9283,N_9277);
nand U9311 (N_9311,N_9241,N_9264);
xor U9312 (N_9312,N_9236,N_9284);
nor U9313 (N_9313,N_9261,N_9260);
nand U9314 (N_9314,N_9271,N_9290);
nand U9315 (N_9315,N_9230,N_9254);
and U9316 (N_9316,N_9258,N_9251);
nor U9317 (N_9317,N_9250,N_9210);
or U9318 (N_9318,N_9265,N_9257);
nand U9319 (N_9319,N_9280,N_9212);
nand U9320 (N_9320,N_9206,N_9263);
and U9321 (N_9321,N_9239,N_9238);
xor U9322 (N_9322,N_9292,N_9245);
xor U9323 (N_9323,N_9228,N_9274);
and U9324 (N_9324,N_9248,N_9243);
nand U9325 (N_9325,N_9227,N_9247);
nand U9326 (N_9326,N_9288,N_9207);
nand U9327 (N_9327,N_9244,N_9296);
or U9328 (N_9328,N_9217,N_9287);
and U9329 (N_9329,N_9233,N_9231);
nand U9330 (N_9330,N_9219,N_9294);
and U9331 (N_9331,N_9267,N_9220);
xnor U9332 (N_9332,N_9234,N_9246);
xor U9333 (N_9333,N_9252,N_9223);
nand U9334 (N_9334,N_9215,N_9259);
nand U9335 (N_9335,N_9266,N_9208);
and U9336 (N_9336,N_9209,N_9256);
or U9337 (N_9337,N_9229,N_9213);
or U9338 (N_9338,N_9235,N_9216);
or U9339 (N_9339,N_9242,N_9272);
nor U9340 (N_9340,N_9279,N_9299);
xnor U9341 (N_9341,N_9221,N_9289);
nor U9342 (N_9342,N_9291,N_9205);
and U9343 (N_9343,N_9225,N_9224);
nor U9344 (N_9344,N_9278,N_9298);
nor U9345 (N_9345,N_9269,N_9268);
nor U9346 (N_9346,N_9253,N_9276);
nor U9347 (N_9347,N_9282,N_9232);
and U9348 (N_9348,N_9203,N_9273);
xnor U9349 (N_9349,N_9211,N_9262);
and U9350 (N_9350,N_9212,N_9205);
or U9351 (N_9351,N_9207,N_9236);
nand U9352 (N_9352,N_9248,N_9255);
and U9353 (N_9353,N_9276,N_9269);
or U9354 (N_9354,N_9235,N_9225);
xnor U9355 (N_9355,N_9208,N_9202);
nand U9356 (N_9356,N_9272,N_9290);
nor U9357 (N_9357,N_9257,N_9234);
nor U9358 (N_9358,N_9252,N_9241);
nand U9359 (N_9359,N_9221,N_9268);
and U9360 (N_9360,N_9258,N_9221);
nand U9361 (N_9361,N_9279,N_9282);
or U9362 (N_9362,N_9246,N_9209);
and U9363 (N_9363,N_9233,N_9296);
nor U9364 (N_9364,N_9295,N_9253);
nor U9365 (N_9365,N_9206,N_9211);
nand U9366 (N_9366,N_9215,N_9231);
nand U9367 (N_9367,N_9253,N_9254);
and U9368 (N_9368,N_9227,N_9279);
and U9369 (N_9369,N_9268,N_9208);
nand U9370 (N_9370,N_9257,N_9278);
or U9371 (N_9371,N_9239,N_9201);
xor U9372 (N_9372,N_9210,N_9283);
nor U9373 (N_9373,N_9299,N_9272);
nor U9374 (N_9374,N_9208,N_9236);
nor U9375 (N_9375,N_9274,N_9205);
and U9376 (N_9376,N_9262,N_9249);
or U9377 (N_9377,N_9279,N_9253);
and U9378 (N_9378,N_9203,N_9242);
xor U9379 (N_9379,N_9227,N_9212);
nor U9380 (N_9380,N_9238,N_9251);
nor U9381 (N_9381,N_9281,N_9222);
and U9382 (N_9382,N_9284,N_9214);
and U9383 (N_9383,N_9242,N_9246);
xor U9384 (N_9384,N_9213,N_9269);
and U9385 (N_9385,N_9281,N_9211);
and U9386 (N_9386,N_9218,N_9277);
and U9387 (N_9387,N_9209,N_9261);
and U9388 (N_9388,N_9229,N_9272);
and U9389 (N_9389,N_9224,N_9256);
and U9390 (N_9390,N_9276,N_9223);
nor U9391 (N_9391,N_9292,N_9251);
and U9392 (N_9392,N_9229,N_9221);
and U9393 (N_9393,N_9291,N_9239);
and U9394 (N_9394,N_9218,N_9205);
nor U9395 (N_9395,N_9234,N_9289);
and U9396 (N_9396,N_9217,N_9268);
nand U9397 (N_9397,N_9278,N_9234);
nor U9398 (N_9398,N_9233,N_9253);
nor U9399 (N_9399,N_9261,N_9219);
nor U9400 (N_9400,N_9372,N_9394);
nand U9401 (N_9401,N_9382,N_9323);
nor U9402 (N_9402,N_9376,N_9331);
or U9403 (N_9403,N_9353,N_9334);
or U9404 (N_9404,N_9301,N_9315);
nor U9405 (N_9405,N_9309,N_9352);
nand U9406 (N_9406,N_9379,N_9362);
nand U9407 (N_9407,N_9359,N_9368);
nor U9408 (N_9408,N_9395,N_9305);
or U9409 (N_9409,N_9348,N_9308);
and U9410 (N_9410,N_9328,N_9312);
xnor U9411 (N_9411,N_9320,N_9314);
nor U9412 (N_9412,N_9391,N_9361);
xnor U9413 (N_9413,N_9399,N_9304);
nand U9414 (N_9414,N_9318,N_9388);
xnor U9415 (N_9415,N_9313,N_9332);
nand U9416 (N_9416,N_9384,N_9370);
or U9417 (N_9417,N_9371,N_9398);
xor U9418 (N_9418,N_9322,N_9397);
nand U9419 (N_9419,N_9326,N_9338);
nor U9420 (N_9420,N_9385,N_9386);
or U9421 (N_9421,N_9364,N_9317);
nor U9422 (N_9422,N_9307,N_9340);
and U9423 (N_9423,N_9381,N_9380);
xnor U9424 (N_9424,N_9390,N_9346);
nand U9425 (N_9425,N_9339,N_9327);
or U9426 (N_9426,N_9393,N_9396);
and U9427 (N_9427,N_9342,N_9343);
nor U9428 (N_9428,N_9347,N_9365);
nand U9429 (N_9429,N_9321,N_9351);
xnor U9430 (N_9430,N_9303,N_9349);
and U9431 (N_9431,N_9392,N_9358);
and U9432 (N_9432,N_9373,N_9374);
and U9433 (N_9433,N_9363,N_9316);
and U9434 (N_9434,N_9378,N_9335);
nand U9435 (N_9435,N_9387,N_9377);
nor U9436 (N_9436,N_9354,N_9375);
or U9437 (N_9437,N_9369,N_9302);
or U9438 (N_9438,N_9360,N_9383);
and U9439 (N_9439,N_9324,N_9356);
and U9440 (N_9440,N_9337,N_9311);
nand U9441 (N_9441,N_9357,N_9341);
and U9442 (N_9442,N_9319,N_9333);
xor U9443 (N_9443,N_9330,N_9336);
nand U9444 (N_9444,N_9310,N_9366);
nor U9445 (N_9445,N_9325,N_9389);
nor U9446 (N_9446,N_9300,N_9367);
and U9447 (N_9447,N_9355,N_9350);
nor U9448 (N_9448,N_9329,N_9344);
nand U9449 (N_9449,N_9306,N_9345);
nor U9450 (N_9450,N_9329,N_9323);
nand U9451 (N_9451,N_9338,N_9387);
nand U9452 (N_9452,N_9392,N_9304);
xor U9453 (N_9453,N_9364,N_9300);
or U9454 (N_9454,N_9354,N_9361);
nand U9455 (N_9455,N_9310,N_9381);
or U9456 (N_9456,N_9373,N_9329);
or U9457 (N_9457,N_9343,N_9360);
nand U9458 (N_9458,N_9308,N_9312);
and U9459 (N_9459,N_9359,N_9396);
and U9460 (N_9460,N_9369,N_9328);
and U9461 (N_9461,N_9344,N_9366);
nor U9462 (N_9462,N_9313,N_9341);
and U9463 (N_9463,N_9330,N_9307);
nor U9464 (N_9464,N_9373,N_9308);
or U9465 (N_9465,N_9343,N_9397);
nand U9466 (N_9466,N_9342,N_9354);
nand U9467 (N_9467,N_9375,N_9344);
nand U9468 (N_9468,N_9379,N_9307);
or U9469 (N_9469,N_9382,N_9393);
and U9470 (N_9470,N_9377,N_9382);
or U9471 (N_9471,N_9332,N_9356);
and U9472 (N_9472,N_9372,N_9304);
nor U9473 (N_9473,N_9347,N_9387);
and U9474 (N_9474,N_9303,N_9362);
nand U9475 (N_9475,N_9349,N_9385);
and U9476 (N_9476,N_9368,N_9304);
or U9477 (N_9477,N_9305,N_9335);
and U9478 (N_9478,N_9335,N_9317);
or U9479 (N_9479,N_9307,N_9344);
nor U9480 (N_9480,N_9354,N_9388);
or U9481 (N_9481,N_9389,N_9384);
xor U9482 (N_9482,N_9323,N_9371);
nor U9483 (N_9483,N_9365,N_9305);
or U9484 (N_9484,N_9358,N_9329);
and U9485 (N_9485,N_9358,N_9349);
nor U9486 (N_9486,N_9387,N_9307);
and U9487 (N_9487,N_9361,N_9325);
and U9488 (N_9488,N_9306,N_9338);
xor U9489 (N_9489,N_9366,N_9307);
and U9490 (N_9490,N_9366,N_9311);
or U9491 (N_9491,N_9317,N_9351);
nor U9492 (N_9492,N_9318,N_9385);
nand U9493 (N_9493,N_9388,N_9384);
nand U9494 (N_9494,N_9360,N_9365);
or U9495 (N_9495,N_9317,N_9300);
nor U9496 (N_9496,N_9334,N_9384);
nand U9497 (N_9497,N_9373,N_9396);
and U9498 (N_9498,N_9343,N_9347);
nor U9499 (N_9499,N_9310,N_9312);
or U9500 (N_9500,N_9459,N_9453);
nand U9501 (N_9501,N_9436,N_9402);
nand U9502 (N_9502,N_9469,N_9466);
and U9503 (N_9503,N_9499,N_9426);
and U9504 (N_9504,N_9488,N_9407);
and U9505 (N_9505,N_9429,N_9465);
or U9506 (N_9506,N_9447,N_9477);
nand U9507 (N_9507,N_9492,N_9431);
nand U9508 (N_9508,N_9484,N_9487);
and U9509 (N_9509,N_9457,N_9490);
or U9510 (N_9510,N_9496,N_9430);
nor U9511 (N_9511,N_9485,N_9461);
xor U9512 (N_9512,N_9467,N_9489);
nand U9513 (N_9513,N_9449,N_9411);
or U9514 (N_9514,N_9495,N_9440);
or U9515 (N_9515,N_9416,N_9423);
and U9516 (N_9516,N_9442,N_9445);
or U9517 (N_9517,N_9486,N_9454);
nor U9518 (N_9518,N_9478,N_9417);
xnor U9519 (N_9519,N_9479,N_9462);
nor U9520 (N_9520,N_9432,N_9433);
and U9521 (N_9521,N_9470,N_9413);
or U9522 (N_9522,N_9448,N_9406);
or U9523 (N_9523,N_9451,N_9420);
xor U9524 (N_9524,N_9481,N_9463);
xnor U9525 (N_9525,N_9419,N_9422);
xnor U9526 (N_9526,N_9491,N_9410);
nor U9527 (N_9527,N_9424,N_9444);
nand U9528 (N_9528,N_9497,N_9455);
nor U9529 (N_9529,N_9498,N_9403);
and U9530 (N_9530,N_9414,N_9474);
nor U9531 (N_9531,N_9472,N_9409);
nor U9532 (N_9532,N_9421,N_9475);
nand U9533 (N_9533,N_9446,N_9401);
and U9534 (N_9534,N_9425,N_9418);
nand U9535 (N_9535,N_9473,N_9464);
and U9536 (N_9536,N_9437,N_9471);
or U9537 (N_9537,N_9458,N_9450);
nand U9538 (N_9538,N_9400,N_9476);
or U9539 (N_9539,N_9434,N_9441);
xnor U9540 (N_9540,N_9482,N_9460);
or U9541 (N_9541,N_9415,N_9493);
nand U9542 (N_9542,N_9408,N_9439);
xor U9543 (N_9543,N_9427,N_9480);
nor U9544 (N_9544,N_9435,N_9404);
and U9545 (N_9545,N_9468,N_9438);
or U9546 (N_9546,N_9483,N_9494);
xnor U9547 (N_9547,N_9452,N_9443);
and U9548 (N_9548,N_9405,N_9428);
nand U9549 (N_9549,N_9412,N_9456);
or U9550 (N_9550,N_9404,N_9441);
and U9551 (N_9551,N_9487,N_9415);
or U9552 (N_9552,N_9455,N_9467);
xnor U9553 (N_9553,N_9403,N_9485);
or U9554 (N_9554,N_9474,N_9482);
nor U9555 (N_9555,N_9448,N_9455);
nand U9556 (N_9556,N_9416,N_9443);
nor U9557 (N_9557,N_9409,N_9494);
or U9558 (N_9558,N_9497,N_9471);
nand U9559 (N_9559,N_9410,N_9421);
nor U9560 (N_9560,N_9409,N_9480);
xnor U9561 (N_9561,N_9454,N_9427);
nor U9562 (N_9562,N_9457,N_9451);
nand U9563 (N_9563,N_9424,N_9415);
nand U9564 (N_9564,N_9407,N_9417);
and U9565 (N_9565,N_9424,N_9422);
and U9566 (N_9566,N_9419,N_9476);
nor U9567 (N_9567,N_9438,N_9439);
or U9568 (N_9568,N_9472,N_9429);
nor U9569 (N_9569,N_9420,N_9465);
or U9570 (N_9570,N_9477,N_9466);
and U9571 (N_9571,N_9428,N_9408);
or U9572 (N_9572,N_9485,N_9438);
and U9573 (N_9573,N_9419,N_9446);
xor U9574 (N_9574,N_9419,N_9436);
nand U9575 (N_9575,N_9485,N_9406);
xor U9576 (N_9576,N_9416,N_9489);
and U9577 (N_9577,N_9419,N_9468);
or U9578 (N_9578,N_9493,N_9403);
nor U9579 (N_9579,N_9408,N_9415);
xor U9580 (N_9580,N_9469,N_9454);
nor U9581 (N_9581,N_9411,N_9468);
nor U9582 (N_9582,N_9478,N_9431);
or U9583 (N_9583,N_9425,N_9466);
nor U9584 (N_9584,N_9487,N_9417);
or U9585 (N_9585,N_9412,N_9470);
and U9586 (N_9586,N_9486,N_9464);
nor U9587 (N_9587,N_9499,N_9406);
and U9588 (N_9588,N_9414,N_9494);
and U9589 (N_9589,N_9487,N_9493);
nand U9590 (N_9590,N_9419,N_9415);
xor U9591 (N_9591,N_9453,N_9409);
and U9592 (N_9592,N_9459,N_9408);
xnor U9593 (N_9593,N_9456,N_9461);
nor U9594 (N_9594,N_9474,N_9434);
nor U9595 (N_9595,N_9462,N_9423);
or U9596 (N_9596,N_9465,N_9413);
and U9597 (N_9597,N_9497,N_9457);
nand U9598 (N_9598,N_9443,N_9425);
or U9599 (N_9599,N_9419,N_9401);
or U9600 (N_9600,N_9562,N_9552);
nand U9601 (N_9601,N_9582,N_9531);
nor U9602 (N_9602,N_9578,N_9527);
nand U9603 (N_9603,N_9536,N_9546);
or U9604 (N_9604,N_9517,N_9590);
nor U9605 (N_9605,N_9542,N_9539);
nand U9606 (N_9606,N_9568,N_9574);
or U9607 (N_9607,N_9535,N_9504);
and U9608 (N_9608,N_9550,N_9588);
or U9609 (N_9609,N_9514,N_9508);
or U9610 (N_9610,N_9577,N_9591);
and U9611 (N_9611,N_9567,N_9511);
nor U9612 (N_9612,N_9579,N_9544);
nor U9613 (N_9613,N_9543,N_9592);
nor U9614 (N_9614,N_9570,N_9503);
xor U9615 (N_9615,N_9500,N_9551);
nor U9616 (N_9616,N_9541,N_9584);
xor U9617 (N_9617,N_9597,N_9532);
and U9618 (N_9618,N_9581,N_9549);
and U9619 (N_9619,N_9554,N_9564);
nand U9620 (N_9620,N_9576,N_9565);
and U9621 (N_9621,N_9507,N_9598);
xnor U9622 (N_9622,N_9594,N_9556);
xor U9623 (N_9623,N_9510,N_9528);
and U9624 (N_9624,N_9583,N_9555);
nand U9625 (N_9625,N_9561,N_9558);
and U9626 (N_9626,N_9566,N_9596);
or U9627 (N_9627,N_9599,N_9553);
and U9628 (N_9628,N_9513,N_9589);
and U9629 (N_9629,N_9560,N_9522);
nor U9630 (N_9630,N_9502,N_9585);
or U9631 (N_9631,N_9580,N_9569);
or U9632 (N_9632,N_9519,N_9559);
or U9633 (N_9633,N_9515,N_9557);
nor U9634 (N_9634,N_9586,N_9525);
nand U9635 (N_9635,N_9524,N_9571);
xor U9636 (N_9636,N_9534,N_9537);
or U9637 (N_9637,N_9538,N_9533);
or U9638 (N_9638,N_9505,N_9506);
nand U9639 (N_9639,N_9512,N_9587);
nand U9640 (N_9640,N_9518,N_9521);
nand U9641 (N_9641,N_9575,N_9509);
nor U9642 (N_9642,N_9545,N_9516);
and U9643 (N_9643,N_9526,N_9540);
nand U9644 (N_9644,N_9573,N_9593);
and U9645 (N_9645,N_9547,N_9523);
and U9646 (N_9646,N_9548,N_9530);
nor U9647 (N_9647,N_9529,N_9572);
nor U9648 (N_9648,N_9563,N_9520);
nor U9649 (N_9649,N_9501,N_9595);
xnor U9650 (N_9650,N_9546,N_9534);
nand U9651 (N_9651,N_9527,N_9546);
and U9652 (N_9652,N_9555,N_9593);
and U9653 (N_9653,N_9500,N_9585);
and U9654 (N_9654,N_9572,N_9516);
and U9655 (N_9655,N_9503,N_9537);
and U9656 (N_9656,N_9580,N_9548);
or U9657 (N_9657,N_9570,N_9580);
nor U9658 (N_9658,N_9598,N_9535);
and U9659 (N_9659,N_9562,N_9558);
nor U9660 (N_9660,N_9515,N_9555);
and U9661 (N_9661,N_9503,N_9550);
or U9662 (N_9662,N_9512,N_9515);
or U9663 (N_9663,N_9543,N_9514);
nand U9664 (N_9664,N_9561,N_9576);
and U9665 (N_9665,N_9587,N_9586);
or U9666 (N_9666,N_9551,N_9570);
or U9667 (N_9667,N_9508,N_9539);
or U9668 (N_9668,N_9532,N_9596);
or U9669 (N_9669,N_9507,N_9544);
or U9670 (N_9670,N_9536,N_9513);
and U9671 (N_9671,N_9528,N_9538);
or U9672 (N_9672,N_9522,N_9515);
and U9673 (N_9673,N_9512,N_9509);
nor U9674 (N_9674,N_9556,N_9549);
and U9675 (N_9675,N_9559,N_9537);
and U9676 (N_9676,N_9595,N_9592);
or U9677 (N_9677,N_9553,N_9536);
nor U9678 (N_9678,N_9529,N_9504);
nand U9679 (N_9679,N_9560,N_9537);
and U9680 (N_9680,N_9587,N_9594);
nor U9681 (N_9681,N_9548,N_9593);
or U9682 (N_9682,N_9502,N_9518);
or U9683 (N_9683,N_9581,N_9570);
xor U9684 (N_9684,N_9536,N_9580);
or U9685 (N_9685,N_9524,N_9591);
and U9686 (N_9686,N_9511,N_9508);
nand U9687 (N_9687,N_9519,N_9569);
nor U9688 (N_9688,N_9514,N_9571);
nand U9689 (N_9689,N_9599,N_9536);
or U9690 (N_9690,N_9579,N_9571);
and U9691 (N_9691,N_9520,N_9575);
nand U9692 (N_9692,N_9581,N_9539);
and U9693 (N_9693,N_9527,N_9589);
nor U9694 (N_9694,N_9542,N_9599);
nor U9695 (N_9695,N_9533,N_9588);
nor U9696 (N_9696,N_9541,N_9531);
nand U9697 (N_9697,N_9540,N_9597);
or U9698 (N_9698,N_9564,N_9527);
or U9699 (N_9699,N_9503,N_9575);
xnor U9700 (N_9700,N_9697,N_9673);
xnor U9701 (N_9701,N_9699,N_9644);
nor U9702 (N_9702,N_9696,N_9646);
nor U9703 (N_9703,N_9652,N_9626);
nor U9704 (N_9704,N_9670,N_9688);
or U9705 (N_9705,N_9665,N_9641);
nor U9706 (N_9706,N_9600,N_9645);
xor U9707 (N_9707,N_9660,N_9686);
or U9708 (N_9708,N_9610,N_9669);
nor U9709 (N_9709,N_9618,N_9601);
and U9710 (N_9710,N_9617,N_9651);
and U9711 (N_9711,N_9614,N_9654);
nand U9712 (N_9712,N_9659,N_9640);
nor U9713 (N_9713,N_9689,N_9625);
and U9714 (N_9714,N_9632,N_9668);
and U9715 (N_9715,N_9642,N_9613);
or U9716 (N_9716,N_9671,N_9623);
xor U9717 (N_9717,N_9607,N_9666);
nand U9718 (N_9718,N_9695,N_9638);
xnor U9719 (N_9719,N_9677,N_9609);
or U9720 (N_9720,N_9657,N_9680);
or U9721 (N_9721,N_9672,N_9616);
nor U9722 (N_9722,N_9636,N_9681);
nor U9723 (N_9723,N_9675,N_9619);
and U9724 (N_9724,N_9629,N_9639);
and U9725 (N_9725,N_9627,N_9608);
xor U9726 (N_9726,N_9631,N_9655);
and U9727 (N_9727,N_9683,N_9647);
and U9728 (N_9728,N_9676,N_9628);
nand U9729 (N_9729,N_9664,N_9662);
nor U9730 (N_9730,N_9687,N_9663);
nand U9731 (N_9731,N_9693,N_9643);
and U9732 (N_9732,N_9694,N_9637);
and U9733 (N_9733,N_9648,N_9621);
and U9734 (N_9734,N_9684,N_9633);
and U9735 (N_9735,N_9604,N_9685);
or U9736 (N_9736,N_9612,N_9656);
nor U9737 (N_9737,N_9692,N_9682);
nor U9738 (N_9738,N_9667,N_9658);
nand U9739 (N_9739,N_9635,N_9653);
or U9740 (N_9740,N_9650,N_9634);
xor U9741 (N_9741,N_9674,N_9615);
or U9742 (N_9742,N_9603,N_9606);
and U9743 (N_9743,N_9602,N_9620);
and U9744 (N_9744,N_9679,N_9630);
nand U9745 (N_9745,N_9691,N_9624);
nor U9746 (N_9746,N_9605,N_9611);
nand U9747 (N_9747,N_9622,N_9678);
or U9748 (N_9748,N_9690,N_9698);
nand U9749 (N_9749,N_9661,N_9649);
nor U9750 (N_9750,N_9637,N_9639);
nor U9751 (N_9751,N_9626,N_9638);
nor U9752 (N_9752,N_9669,N_9627);
nand U9753 (N_9753,N_9680,N_9695);
or U9754 (N_9754,N_9669,N_9603);
xnor U9755 (N_9755,N_9696,N_9692);
xnor U9756 (N_9756,N_9668,N_9665);
xor U9757 (N_9757,N_9601,N_9690);
nor U9758 (N_9758,N_9652,N_9616);
nor U9759 (N_9759,N_9642,N_9636);
nand U9760 (N_9760,N_9626,N_9615);
nor U9761 (N_9761,N_9664,N_9666);
xor U9762 (N_9762,N_9672,N_9608);
nand U9763 (N_9763,N_9613,N_9654);
xnor U9764 (N_9764,N_9623,N_9673);
nor U9765 (N_9765,N_9661,N_9698);
nor U9766 (N_9766,N_9615,N_9645);
or U9767 (N_9767,N_9694,N_9602);
nor U9768 (N_9768,N_9674,N_9665);
and U9769 (N_9769,N_9640,N_9616);
or U9770 (N_9770,N_9675,N_9639);
or U9771 (N_9771,N_9657,N_9608);
nor U9772 (N_9772,N_9656,N_9689);
nor U9773 (N_9773,N_9645,N_9614);
xnor U9774 (N_9774,N_9655,N_9675);
xnor U9775 (N_9775,N_9671,N_9605);
xor U9776 (N_9776,N_9667,N_9684);
nor U9777 (N_9777,N_9662,N_9673);
or U9778 (N_9778,N_9658,N_9665);
nor U9779 (N_9779,N_9678,N_9677);
nand U9780 (N_9780,N_9611,N_9633);
nor U9781 (N_9781,N_9679,N_9606);
nor U9782 (N_9782,N_9685,N_9680);
nor U9783 (N_9783,N_9697,N_9686);
xor U9784 (N_9784,N_9652,N_9686);
and U9785 (N_9785,N_9630,N_9671);
nand U9786 (N_9786,N_9626,N_9677);
nand U9787 (N_9787,N_9627,N_9622);
nand U9788 (N_9788,N_9690,N_9692);
or U9789 (N_9789,N_9643,N_9696);
nor U9790 (N_9790,N_9680,N_9674);
or U9791 (N_9791,N_9668,N_9634);
nand U9792 (N_9792,N_9618,N_9699);
nand U9793 (N_9793,N_9649,N_9642);
and U9794 (N_9794,N_9632,N_9667);
and U9795 (N_9795,N_9654,N_9676);
or U9796 (N_9796,N_9656,N_9645);
xnor U9797 (N_9797,N_9664,N_9620);
or U9798 (N_9798,N_9641,N_9672);
nand U9799 (N_9799,N_9675,N_9616);
nor U9800 (N_9800,N_9748,N_9796);
nor U9801 (N_9801,N_9784,N_9754);
nand U9802 (N_9802,N_9763,N_9771);
nor U9803 (N_9803,N_9715,N_9781);
or U9804 (N_9804,N_9712,N_9780);
or U9805 (N_9805,N_9795,N_9765);
nand U9806 (N_9806,N_9705,N_9737);
xnor U9807 (N_9807,N_9792,N_9730);
and U9808 (N_9808,N_9764,N_9794);
xnor U9809 (N_9809,N_9752,N_9759);
and U9810 (N_9810,N_9710,N_9777);
and U9811 (N_9811,N_9721,N_9704);
or U9812 (N_9812,N_9741,N_9702);
and U9813 (N_9813,N_9776,N_9797);
nand U9814 (N_9814,N_9798,N_9756);
and U9815 (N_9815,N_9724,N_9708);
nand U9816 (N_9816,N_9774,N_9700);
nor U9817 (N_9817,N_9713,N_9709);
xor U9818 (N_9818,N_9782,N_9738);
xnor U9819 (N_9819,N_9740,N_9739);
and U9820 (N_9820,N_9714,N_9703);
nor U9821 (N_9821,N_9734,N_9720);
and U9822 (N_9822,N_9783,N_9729);
nand U9823 (N_9823,N_9768,N_9717);
nand U9824 (N_9824,N_9799,N_9727);
xnor U9825 (N_9825,N_9723,N_9791);
or U9826 (N_9826,N_9707,N_9790);
xor U9827 (N_9827,N_9789,N_9767);
nor U9828 (N_9828,N_9718,N_9722);
or U9829 (N_9829,N_9762,N_9753);
nor U9830 (N_9830,N_9716,N_9725);
nor U9831 (N_9831,N_9755,N_9743);
nand U9832 (N_9832,N_9793,N_9706);
nor U9833 (N_9833,N_9746,N_9751);
or U9834 (N_9834,N_9772,N_9731);
nand U9835 (N_9835,N_9788,N_9775);
and U9836 (N_9836,N_9747,N_9757);
or U9837 (N_9837,N_9787,N_9711);
or U9838 (N_9838,N_9728,N_9766);
nor U9839 (N_9839,N_9719,N_9786);
or U9840 (N_9840,N_9785,N_9744);
or U9841 (N_9841,N_9773,N_9779);
nand U9842 (N_9842,N_9726,N_9733);
xnor U9843 (N_9843,N_9761,N_9732);
or U9844 (N_9844,N_9701,N_9742);
or U9845 (N_9845,N_9735,N_9736);
and U9846 (N_9846,N_9769,N_9749);
or U9847 (N_9847,N_9760,N_9770);
or U9848 (N_9848,N_9758,N_9778);
nand U9849 (N_9849,N_9745,N_9750);
or U9850 (N_9850,N_9705,N_9753);
nand U9851 (N_9851,N_9781,N_9771);
or U9852 (N_9852,N_9757,N_9778);
and U9853 (N_9853,N_9759,N_9708);
nor U9854 (N_9854,N_9751,N_9779);
or U9855 (N_9855,N_9752,N_9734);
nor U9856 (N_9856,N_9723,N_9752);
and U9857 (N_9857,N_9743,N_9776);
or U9858 (N_9858,N_9798,N_9744);
or U9859 (N_9859,N_9767,N_9796);
nand U9860 (N_9860,N_9730,N_9716);
and U9861 (N_9861,N_9729,N_9707);
nor U9862 (N_9862,N_9741,N_9781);
or U9863 (N_9863,N_9796,N_9768);
or U9864 (N_9864,N_9724,N_9705);
nand U9865 (N_9865,N_9791,N_9742);
and U9866 (N_9866,N_9751,N_9702);
nand U9867 (N_9867,N_9784,N_9728);
nor U9868 (N_9868,N_9772,N_9739);
and U9869 (N_9869,N_9764,N_9791);
xnor U9870 (N_9870,N_9737,N_9744);
or U9871 (N_9871,N_9775,N_9784);
nand U9872 (N_9872,N_9731,N_9740);
nor U9873 (N_9873,N_9752,N_9771);
nor U9874 (N_9874,N_9736,N_9762);
nand U9875 (N_9875,N_9702,N_9786);
nand U9876 (N_9876,N_9779,N_9748);
nor U9877 (N_9877,N_9791,N_9795);
nand U9878 (N_9878,N_9733,N_9745);
or U9879 (N_9879,N_9769,N_9713);
nand U9880 (N_9880,N_9788,N_9798);
xor U9881 (N_9881,N_9721,N_9723);
nand U9882 (N_9882,N_9775,N_9787);
nor U9883 (N_9883,N_9705,N_9775);
or U9884 (N_9884,N_9739,N_9765);
nor U9885 (N_9885,N_9769,N_9796);
nor U9886 (N_9886,N_9717,N_9708);
xnor U9887 (N_9887,N_9763,N_9797);
nand U9888 (N_9888,N_9769,N_9740);
nand U9889 (N_9889,N_9794,N_9762);
nor U9890 (N_9890,N_9740,N_9798);
and U9891 (N_9891,N_9706,N_9711);
nand U9892 (N_9892,N_9717,N_9776);
or U9893 (N_9893,N_9715,N_9729);
xnor U9894 (N_9894,N_9712,N_9732);
nand U9895 (N_9895,N_9728,N_9729);
nand U9896 (N_9896,N_9739,N_9779);
nor U9897 (N_9897,N_9757,N_9762);
or U9898 (N_9898,N_9773,N_9742);
nand U9899 (N_9899,N_9703,N_9734);
nand U9900 (N_9900,N_9821,N_9835);
and U9901 (N_9901,N_9800,N_9884);
nor U9902 (N_9902,N_9882,N_9881);
and U9903 (N_9903,N_9829,N_9807);
or U9904 (N_9904,N_9866,N_9859);
and U9905 (N_9905,N_9879,N_9886);
nor U9906 (N_9906,N_9818,N_9885);
nand U9907 (N_9907,N_9880,N_9873);
nand U9908 (N_9908,N_9874,N_9806);
and U9909 (N_9909,N_9809,N_9814);
and U9910 (N_9910,N_9837,N_9867);
nand U9911 (N_9911,N_9825,N_9853);
and U9912 (N_9912,N_9839,N_9832);
or U9913 (N_9913,N_9864,N_9812);
nor U9914 (N_9914,N_9841,N_9815);
and U9915 (N_9915,N_9870,N_9895);
xor U9916 (N_9916,N_9892,N_9869);
or U9917 (N_9917,N_9803,N_9872);
nand U9918 (N_9918,N_9876,N_9877);
nor U9919 (N_9919,N_9858,N_9830);
and U9920 (N_9920,N_9893,N_9819);
and U9921 (N_9921,N_9810,N_9890);
and U9922 (N_9922,N_9848,N_9801);
nand U9923 (N_9923,N_9843,N_9833);
nor U9924 (N_9924,N_9861,N_9888);
nor U9925 (N_9925,N_9871,N_9822);
xor U9926 (N_9926,N_9898,N_9811);
nand U9927 (N_9927,N_9863,N_9852);
nand U9928 (N_9928,N_9891,N_9878);
nand U9929 (N_9929,N_9855,N_9849);
nor U9930 (N_9930,N_9816,N_9862);
or U9931 (N_9931,N_9827,N_9828);
nand U9932 (N_9932,N_9868,N_9817);
and U9933 (N_9933,N_9836,N_9865);
or U9934 (N_9934,N_9857,N_9804);
nor U9935 (N_9935,N_9820,N_9856);
xor U9936 (N_9936,N_9899,N_9813);
and U9937 (N_9937,N_9842,N_9845);
and U9938 (N_9938,N_9851,N_9847);
and U9939 (N_9939,N_9883,N_9805);
nor U9940 (N_9940,N_9834,N_9838);
xor U9941 (N_9941,N_9887,N_9897);
nor U9942 (N_9942,N_9846,N_9896);
or U9943 (N_9943,N_9802,N_9860);
nor U9944 (N_9944,N_9826,N_9889);
nand U9945 (N_9945,N_9854,N_9840);
nor U9946 (N_9946,N_9875,N_9824);
nand U9947 (N_9947,N_9831,N_9894);
or U9948 (N_9948,N_9850,N_9823);
nor U9949 (N_9949,N_9808,N_9844);
and U9950 (N_9950,N_9855,N_9848);
and U9951 (N_9951,N_9877,N_9838);
xnor U9952 (N_9952,N_9866,N_9841);
nor U9953 (N_9953,N_9892,N_9818);
and U9954 (N_9954,N_9813,N_9847);
and U9955 (N_9955,N_9822,N_9882);
and U9956 (N_9956,N_9863,N_9866);
and U9957 (N_9957,N_9828,N_9892);
and U9958 (N_9958,N_9893,N_9843);
and U9959 (N_9959,N_9887,N_9884);
nor U9960 (N_9960,N_9839,N_9805);
and U9961 (N_9961,N_9816,N_9821);
and U9962 (N_9962,N_9849,N_9856);
or U9963 (N_9963,N_9819,N_9826);
nand U9964 (N_9964,N_9841,N_9852);
or U9965 (N_9965,N_9828,N_9856);
nor U9966 (N_9966,N_9852,N_9809);
nand U9967 (N_9967,N_9811,N_9863);
or U9968 (N_9968,N_9860,N_9881);
nor U9969 (N_9969,N_9848,N_9806);
xor U9970 (N_9970,N_9823,N_9879);
or U9971 (N_9971,N_9815,N_9879);
nor U9972 (N_9972,N_9827,N_9885);
and U9973 (N_9973,N_9855,N_9859);
nor U9974 (N_9974,N_9835,N_9817);
xor U9975 (N_9975,N_9862,N_9876);
and U9976 (N_9976,N_9850,N_9886);
nor U9977 (N_9977,N_9894,N_9817);
and U9978 (N_9978,N_9828,N_9872);
or U9979 (N_9979,N_9846,N_9892);
nand U9980 (N_9980,N_9813,N_9868);
xor U9981 (N_9981,N_9852,N_9833);
nor U9982 (N_9982,N_9831,N_9820);
and U9983 (N_9983,N_9873,N_9876);
nor U9984 (N_9984,N_9802,N_9859);
nor U9985 (N_9985,N_9852,N_9828);
or U9986 (N_9986,N_9870,N_9832);
and U9987 (N_9987,N_9808,N_9846);
and U9988 (N_9988,N_9808,N_9891);
or U9989 (N_9989,N_9863,N_9835);
or U9990 (N_9990,N_9803,N_9858);
nand U9991 (N_9991,N_9807,N_9830);
nand U9992 (N_9992,N_9847,N_9890);
nor U9993 (N_9993,N_9804,N_9843);
and U9994 (N_9994,N_9880,N_9881);
nor U9995 (N_9995,N_9850,N_9851);
nand U9996 (N_9996,N_9842,N_9890);
and U9997 (N_9997,N_9806,N_9889);
and U9998 (N_9998,N_9877,N_9837);
or U9999 (N_9999,N_9840,N_9831);
nor UO_0 (O_0,N_9985,N_9962);
nand UO_1 (O_1,N_9945,N_9911);
and UO_2 (O_2,N_9944,N_9908);
nor UO_3 (O_3,N_9990,N_9946);
xor UO_4 (O_4,N_9915,N_9903);
nor UO_5 (O_5,N_9978,N_9984);
nor UO_6 (O_6,N_9969,N_9939);
nand UO_7 (O_7,N_9997,N_9981);
nand UO_8 (O_8,N_9904,N_9953);
or UO_9 (O_9,N_9986,N_9922);
nor UO_10 (O_10,N_9954,N_9974);
nor UO_11 (O_11,N_9947,N_9909);
or UO_12 (O_12,N_9941,N_9987);
or UO_13 (O_13,N_9937,N_9991);
and UO_14 (O_14,N_9914,N_9917);
or UO_15 (O_15,N_9994,N_9973);
xnor UO_16 (O_16,N_9952,N_9967);
xor UO_17 (O_17,N_9966,N_9918);
or UO_18 (O_18,N_9906,N_9907);
nand UO_19 (O_19,N_9976,N_9971);
nor UO_20 (O_20,N_9921,N_9940);
xnor UO_21 (O_21,N_9988,N_9910);
nor UO_22 (O_22,N_9963,N_9905);
or UO_23 (O_23,N_9965,N_9934);
nand UO_24 (O_24,N_9989,N_9960);
and UO_25 (O_25,N_9970,N_9928);
nor UO_26 (O_26,N_9927,N_9929);
nand UO_27 (O_27,N_9935,N_9995);
xnor UO_28 (O_28,N_9900,N_9933);
and UO_29 (O_29,N_9938,N_9996);
and UO_30 (O_30,N_9950,N_9968);
nand UO_31 (O_31,N_9943,N_9916);
and UO_32 (O_32,N_9936,N_9980);
nand UO_33 (O_33,N_9902,N_9979);
or UO_34 (O_34,N_9961,N_9942);
and UO_35 (O_35,N_9993,N_9923);
or UO_36 (O_36,N_9951,N_9925);
or UO_37 (O_37,N_9975,N_9920);
and UO_38 (O_38,N_9999,N_9913);
and UO_39 (O_39,N_9956,N_9926);
nand UO_40 (O_40,N_9977,N_9992);
and UO_41 (O_41,N_9982,N_9983);
xnor UO_42 (O_42,N_9948,N_9957);
and UO_43 (O_43,N_9919,N_9998);
nand UO_44 (O_44,N_9959,N_9930);
nand UO_45 (O_45,N_9912,N_9931);
nor UO_46 (O_46,N_9958,N_9964);
nor UO_47 (O_47,N_9924,N_9949);
or UO_48 (O_48,N_9955,N_9901);
and UO_49 (O_49,N_9932,N_9972);
nand UO_50 (O_50,N_9994,N_9902);
nor UO_51 (O_51,N_9978,N_9925);
or UO_52 (O_52,N_9905,N_9934);
nor UO_53 (O_53,N_9933,N_9912);
and UO_54 (O_54,N_9920,N_9911);
xnor UO_55 (O_55,N_9960,N_9923);
nor UO_56 (O_56,N_9953,N_9985);
xnor UO_57 (O_57,N_9998,N_9996);
or UO_58 (O_58,N_9986,N_9943);
nor UO_59 (O_59,N_9974,N_9991);
nand UO_60 (O_60,N_9903,N_9981);
or UO_61 (O_61,N_9927,N_9947);
nor UO_62 (O_62,N_9934,N_9903);
and UO_63 (O_63,N_9978,N_9918);
xor UO_64 (O_64,N_9948,N_9997);
nor UO_65 (O_65,N_9918,N_9927);
or UO_66 (O_66,N_9950,N_9930);
and UO_67 (O_67,N_9964,N_9940);
or UO_68 (O_68,N_9945,N_9927);
nor UO_69 (O_69,N_9975,N_9969);
nand UO_70 (O_70,N_9940,N_9936);
nand UO_71 (O_71,N_9999,N_9919);
nand UO_72 (O_72,N_9961,N_9937);
or UO_73 (O_73,N_9985,N_9977);
nor UO_74 (O_74,N_9925,N_9975);
nand UO_75 (O_75,N_9945,N_9994);
nand UO_76 (O_76,N_9951,N_9982);
or UO_77 (O_77,N_9903,N_9939);
nand UO_78 (O_78,N_9983,N_9907);
and UO_79 (O_79,N_9996,N_9911);
nor UO_80 (O_80,N_9935,N_9956);
or UO_81 (O_81,N_9928,N_9962);
xor UO_82 (O_82,N_9942,N_9900);
or UO_83 (O_83,N_9909,N_9977);
nor UO_84 (O_84,N_9986,N_9990);
or UO_85 (O_85,N_9968,N_9943);
nor UO_86 (O_86,N_9940,N_9934);
and UO_87 (O_87,N_9937,N_9920);
nor UO_88 (O_88,N_9938,N_9934);
nor UO_89 (O_89,N_9909,N_9940);
xor UO_90 (O_90,N_9927,N_9958);
or UO_91 (O_91,N_9941,N_9901);
nor UO_92 (O_92,N_9915,N_9989);
and UO_93 (O_93,N_9936,N_9979);
nor UO_94 (O_94,N_9959,N_9986);
nand UO_95 (O_95,N_9945,N_9937);
or UO_96 (O_96,N_9986,N_9995);
nor UO_97 (O_97,N_9986,N_9945);
or UO_98 (O_98,N_9964,N_9966);
or UO_99 (O_99,N_9980,N_9955);
nor UO_100 (O_100,N_9954,N_9926);
and UO_101 (O_101,N_9908,N_9961);
nor UO_102 (O_102,N_9942,N_9932);
and UO_103 (O_103,N_9909,N_9957);
or UO_104 (O_104,N_9973,N_9997);
nand UO_105 (O_105,N_9921,N_9906);
nand UO_106 (O_106,N_9903,N_9941);
and UO_107 (O_107,N_9959,N_9995);
nor UO_108 (O_108,N_9911,N_9946);
or UO_109 (O_109,N_9955,N_9969);
and UO_110 (O_110,N_9903,N_9925);
or UO_111 (O_111,N_9972,N_9973);
and UO_112 (O_112,N_9910,N_9921);
or UO_113 (O_113,N_9909,N_9959);
and UO_114 (O_114,N_9937,N_9979);
nor UO_115 (O_115,N_9972,N_9920);
and UO_116 (O_116,N_9995,N_9976);
nand UO_117 (O_117,N_9960,N_9963);
nor UO_118 (O_118,N_9976,N_9957);
nand UO_119 (O_119,N_9981,N_9938);
nand UO_120 (O_120,N_9922,N_9991);
or UO_121 (O_121,N_9916,N_9988);
nand UO_122 (O_122,N_9948,N_9935);
nor UO_123 (O_123,N_9905,N_9909);
or UO_124 (O_124,N_9920,N_9928);
nand UO_125 (O_125,N_9955,N_9945);
nor UO_126 (O_126,N_9982,N_9915);
or UO_127 (O_127,N_9982,N_9924);
and UO_128 (O_128,N_9963,N_9926);
and UO_129 (O_129,N_9959,N_9907);
or UO_130 (O_130,N_9961,N_9936);
and UO_131 (O_131,N_9904,N_9963);
or UO_132 (O_132,N_9944,N_9995);
nor UO_133 (O_133,N_9905,N_9987);
xnor UO_134 (O_134,N_9991,N_9984);
and UO_135 (O_135,N_9968,N_9931);
nand UO_136 (O_136,N_9903,N_9964);
nor UO_137 (O_137,N_9903,N_9989);
nand UO_138 (O_138,N_9985,N_9904);
xnor UO_139 (O_139,N_9935,N_9915);
or UO_140 (O_140,N_9955,N_9989);
nand UO_141 (O_141,N_9930,N_9936);
or UO_142 (O_142,N_9982,N_9901);
and UO_143 (O_143,N_9988,N_9948);
or UO_144 (O_144,N_9967,N_9937);
or UO_145 (O_145,N_9914,N_9972);
nor UO_146 (O_146,N_9906,N_9973);
nor UO_147 (O_147,N_9957,N_9992);
nor UO_148 (O_148,N_9946,N_9989);
nand UO_149 (O_149,N_9998,N_9910);
or UO_150 (O_150,N_9957,N_9932);
or UO_151 (O_151,N_9945,N_9932);
and UO_152 (O_152,N_9967,N_9944);
and UO_153 (O_153,N_9972,N_9979);
nor UO_154 (O_154,N_9916,N_9949);
and UO_155 (O_155,N_9923,N_9989);
nor UO_156 (O_156,N_9969,N_9977);
and UO_157 (O_157,N_9977,N_9974);
nand UO_158 (O_158,N_9974,N_9998);
xor UO_159 (O_159,N_9997,N_9906);
or UO_160 (O_160,N_9979,N_9922);
nor UO_161 (O_161,N_9909,N_9915);
or UO_162 (O_162,N_9945,N_9998);
and UO_163 (O_163,N_9928,N_9957);
xor UO_164 (O_164,N_9930,N_9965);
nor UO_165 (O_165,N_9961,N_9934);
xnor UO_166 (O_166,N_9948,N_9917);
nor UO_167 (O_167,N_9959,N_9926);
xnor UO_168 (O_168,N_9985,N_9905);
or UO_169 (O_169,N_9944,N_9950);
or UO_170 (O_170,N_9902,N_9920);
nor UO_171 (O_171,N_9916,N_9992);
or UO_172 (O_172,N_9917,N_9988);
nand UO_173 (O_173,N_9979,N_9920);
xnor UO_174 (O_174,N_9931,N_9976);
nand UO_175 (O_175,N_9957,N_9963);
nand UO_176 (O_176,N_9979,N_9983);
nor UO_177 (O_177,N_9994,N_9913);
or UO_178 (O_178,N_9902,N_9967);
nand UO_179 (O_179,N_9977,N_9907);
nor UO_180 (O_180,N_9924,N_9976);
nand UO_181 (O_181,N_9923,N_9982);
or UO_182 (O_182,N_9968,N_9992);
and UO_183 (O_183,N_9969,N_9930);
xor UO_184 (O_184,N_9908,N_9997);
nand UO_185 (O_185,N_9912,N_9979);
or UO_186 (O_186,N_9936,N_9906);
and UO_187 (O_187,N_9906,N_9971);
and UO_188 (O_188,N_9946,N_9903);
nor UO_189 (O_189,N_9909,N_9943);
xor UO_190 (O_190,N_9919,N_9948);
xor UO_191 (O_191,N_9970,N_9993);
nand UO_192 (O_192,N_9973,N_9969);
or UO_193 (O_193,N_9981,N_9998);
or UO_194 (O_194,N_9962,N_9967);
nor UO_195 (O_195,N_9988,N_9926);
or UO_196 (O_196,N_9924,N_9937);
or UO_197 (O_197,N_9987,N_9985);
xor UO_198 (O_198,N_9968,N_9944);
and UO_199 (O_199,N_9917,N_9989);
nand UO_200 (O_200,N_9985,N_9954);
nand UO_201 (O_201,N_9914,N_9950);
nand UO_202 (O_202,N_9943,N_9939);
or UO_203 (O_203,N_9919,N_9982);
and UO_204 (O_204,N_9942,N_9960);
and UO_205 (O_205,N_9900,N_9995);
and UO_206 (O_206,N_9900,N_9971);
nand UO_207 (O_207,N_9927,N_9901);
xnor UO_208 (O_208,N_9916,N_9941);
nand UO_209 (O_209,N_9983,N_9915);
nor UO_210 (O_210,N_9940,N_9960);
xnor UO_211 (O_211,N_9997,N_9952);
and UO_212 (O_212,N_9959,N_9943);
or UO_213 (O_213,N_9920,N_9908);
nand UO_214 (O_214,N_9990,N_9917);
xnor UO_215 (O_215,N_9985,N_9944);
nand UO_216 (O_216,N_9934,N_9955);
or UO_217 (O_217,N_9946,N_9910);
and UO_218 (O_218,N_9918,N_9910);
nor UO_219 (O_219,N_9911,N_9919);
and UO_220 (O_220,N_9912,N_9900);
nor UO_221 (O_221,N_9906,N_9964);
nor UO_222 (O_222,N_9997,N_9936);
and UO_223 (O_223,N_9915,N_9947);
or UO_224 (O_224,N_9910,N_9995);
xor UO_225 (O_225,N_9954,N_9930);
xnor UO_226 (O_226,N_9982,N_9929);
and UO_227 (O_227,N_9942,N_9996);
or UO_228 (O_228,N_9917,N_9980);
nand UO_229 (O_229,N_9986,N_9955);
or UO_230 (O_230,N_9920,N_9906);
and UO_231 (O_231,N_9982,N_9909);
or UO_232 (O_232,N_9922,N_9988);
nand UO_233 (O_233,N_9935,N_9901);
xnor UO_234 (O_234,N_9948,N_9920);
and UO_235 (O_235,N_9999,N_9990);
or UO_236 (O_236,N_9980,N_9934);
xnor UO_237 (O_237,N_9934,N_9942);
and UO_238 (O_238,N_9946,N_9994);
and UO_239 (O_239,N_9908,N_9971);
and UO_240 (O_240,N_9968,N_9971);
xnor UO_241 (O_241,N_9972,N_9912);
or UO_242 (O_242,N_9931,N_9922);
nand UO_243 (O_243,N_9972,N_9950);
and UO_244 (O_244,N_9925,N_9917);
nand UO_245 (O_245,N_9900,N_9903);
xor UO_246 (O_246,N_9938,N_9940);
and UO_247 (O_247,N_9904,N_9951);
or UO_248 (O_248,N_9908,N_9914);
nand UO_249 (O_249,N_9953,N_9974);
and UO_250 (O_250,N_9917,N_9924);
nand UO_251 (O_251,N_9987,N_9918);
or UO_252 (O_252,N_9999,N_9997);
and UO_253 (O_253,N_9977,N_9991);
and UO_254 (O_254,N_9959,N_9997);
and UO_255 (O_255,N_9904,N_9917);
nor UO_256 (O_256,N_9919,N_9910);
nand UO_257 (O_257,N_9901,N_9995);
nand UO_258 (O_258,N_9992,N_9920);
and UO_259 (O_259,N_9902,N_9915);
nor UO_260 (O_260,N_9975,N_9931);
nor UO_261 (O_261,N_9969,N_9927);
nor UO_262 (O_262,N_9975,N_9990);
and UO_263 (O_263,N_9996,N_9952);
nand UO_264 (O_264,N_9993,N_9949);
nor UO_265 (O_265,N_9918,N_9938);
xor UO_266 (O_266,N_9931,N_9989);
and UO_267 (O_267,N_9907,N_9925);
and UO_268 (O_268,N_9986,N_9984);
nor UO_269 (O_269,N_9950,N_9973);
nor UO_270 (O_270,N_9971,N_9987);
nand UO_271 (O_271,N_9968,N_9929);
and UO_272 (O_272,N_9932,N_9975);
xor UO_273 (O_273,N_9968,N_9961);
nor UO_274 (O_274,N_9941,N_9913);
nand UO_275 (O_275,N_9932,N_9968);
nor UO_276 (O_276,N_9936,N_9946);
or UO_277 (O_277,N_9953,N_9943);
nand UO_278 (O_278,N_9909,N_9965);
nor UO_279 (O_279,N_9947,N_9901);
nor UO_280 (O_280,N_9997,N_9946);
nor UO_281 (O_281,N_9925,N_9912);
nand UO_282 (O_282,N_9921,N_9914);
xnor UO_283 (O_283,N_9944,N_9981);
and UO_284 (O_284,N_9978,N_9948);
nor UO_285 (O_285,N_9944,N_9970);
and UO_286 (O_286,N_9997,N_9985);
nor UO_287 (O_287,N_9941,N_9994);
nor UO_288 (O_288,N_9922,N_9992);
and UO_289 (O_289,N_9984,N_9947);
or UO_290 (O_290,N_9992,N_9900);
nor UO_291 (O_291,N_9942,N_9923);
nand UO_292 (O_292,N_9985,N_9975);
nor UO_293 (O_293,N_9912,N_9992);
nor UO_294 (O_294,N_9923,N_9932);
nand UO_295 (O_295,N_9950,N_9929);
and UO_296 (O_296,N_9934,N_9974);
nor UO_297 (O_297,N_9911,N_9949);
or UO_298 (O_298,N_9965,N_9990);
or UO_299 (O_299,N_9916,N_9908);
or UO_300 (O_300,N_9901,N_9926);
or UO_301 (O_301,N_9965,N_9977);
or UO_302 (O_302,N_9930,N_9942);
xnor UO_303 (O_303,N_9905,N_9941);
nand UO_304 (O_304,N_9983,N_9959);
and UO_305 (O_305,N_9918,N_9965);
or UO_306 (O_306,N_9972,N_9977);
nor UO_307 (O_307,N_9970,N_9945);
nand UO_308 (O_308,N_9931,N_9927);
nand UO_309 (O_309,N_9901,N_9962);
and UO_310 (O_310,N_9990,N_9914);
nand UO_311 (O_311,N_9900,N_9905);
nand UO_312 (O_312,N_9960,N_9993);
nor UO_313 (O_313,N_9902,N_9980);
or UO_314 (O_314,N_9907,N_9919);
and UO_315 (O_315,N_9994,N_9966);
or UO_316 (O_316,N_9936,N_9996);
xor UO_317 (O_317,N_9929,N_9989);
and UO_318 (O_318,N_9916,N_9917);
or UO_319 (O_319,N_9947,N_9965);
nor UO_320 (O_320,N_9968,N_9970);
nor UO_321 (O_321,N_9995,N_9938);
xnor UO_322 (O_322,N_9981,N_9941);
and UO_323 (O_323,N_9969,N_9984);
and UO_324 (O_324,N_9913,N_9912);
and UO_325 (O_325,N_9957,N_9977);
and UO_326 (O_326,N_9952,N_9980);
nand UO_327 (O_327,N_9928,N_9999);
and UO_328 (O_328,N_9916,N_9940);
nand UO_329 (O_329,N_9987,N_9975);
xor UO_330 (O_330,N_9983,N_9998);
nor UO_331 (O_331,N_9980,N_9916);
and UO_332 (O_332,N_9909,N_9983);
or UO_333 (O_333,N_9981,N_9969);
or UO_334 (O_334,N_9949,N_9900);
or UO_335 (O_335,N_9907,N_9944);
or UO_336 (O_336,N_9979,N_9957);
or UO_337 (O_337,N_9994,N_9972);
and UO_338 (O_338,N_9970,N_9908);
or UO_339 (O_339,N_9983,N_9928);
and UO_340 (O_340,N_9972,N_9974);
nor UO_341 (O_341,N_9917,N_9906);
nor UO_342 (O_342,N_9921,N_9978);
or UO_343 (O_343,N_9912,N_9915);
and UO_344 (O_344,N_9921,N_9961);
nor UO_345 (O_345,N_9931,N_9994);
nor UO_346 (O_346,N_9951,N_9973);
and UO_347 (O_347,N_9933,N_9906);
nand UO_348 (O_348,N_9956,N_9979);
nand UO_349 (O_349,N_9939,N_9934);
nor UO_350 (O_350,N_9948,N_9921);
and UO_351 (O_351,N_9953,N_9983);
nor UO_352 (O_352,N_9984,N_9905);
nor UO_353 (O_353,N_9996,N_9915);
nor UO_354 (O_354,N_9977,N_9936);
or UO_355 (O_355,N_9938,N_9931);
nand UO_356 (O_356,N_9987,N_9969);
nand UO_357 (O_357,N_9956,N_9984);
nor UO_358 (O_358,N_9907,N_9999);
and UO_359 (O_359,N_9986,N_9999);
nor UO_360 (O_360,N_9963,N_9977);
or UO_361 (O_361,N_9975,N_9902);
xnor UO_362 (O_362,N_9953,N_9986);
nand UO_363 (O_363,N_9924,N_9960);
xnor UO_364 (O_364,N_9967,N_9983);
nor UO_365 (O_365,N_9976,N_9992);
nor UO_366 (O_366,N_9992,N_9959);
nand UO_367 (O_367,N_9930,N_9924);
nand UO_368 (O_368,N_9915,N_9970);
xnor UO_369 (O_369,N_9980,N_9931);
or UO_370 (O_370,N_9974,N_9961);
or UO_371 (O_371,N_9986,N_9985);
and UO_372 (O_372,N_9942,N_9910);
nor UO_373 (O_373,N_9972,N_9999);
or UO_374 (O_374,N_9948,N_9901);
nand UO_375 (O_375,N_9957,N_9959);
nor UO_376 (O_376,N_9981,N_9970);
nand UO_377 (O_377,N_9932,N_9907);
or UO_378 (O_378,N_9913,N_9940);
and UO_379 (O_379,N_9994,N_9992);
nor UO_380 (O_380,N_9937,N_9974);
and UO_381 (O_381,N_9948,N_9964);
xnor UO_382 (O_382,N_9916,N_9956);
nand UO_383 (O_383,N_9996,N_9976);
and UO_384 (O_384,N_9997,N_9902);
nand UO_385 (O_385,N_9902,N_9908);
nand UO_386 (O_386,N_9935,N_9963);
and UO_387 (O_387,N_9948,N_9973);
or UO_388 (O_388,N_9971,N_9958);
or UO_389 (O_389,N_9997,N_9965);
or UO_390 (O_390,N_9992,N_9974);
nand UO_391 (O_391,N_9944,N_9923);
and UO_392 (O_392,N_9930,N_9994);
nand UO_393 (O_393,N_9989,N_9954);
nand UO_394 (O_394,N_9935,N_9902);
nor UO_395 (O_395,N_9955,N_9960);
or UO_396 (O_396,N_9907,N_9903);
or UO_397 (O_397,N_9997,N_9945);
nor UO_398 (O_398,N_9910,N_9974);
nand UO_399 (O_399,N_9929,N_9992);
nand UO_400 (O_400,N_9942,N_9914);
nand UO_401 (O_401,N_9938,N_9939);
and UO_402 (O_402,N_9971,N_9917);
or UO_403 (O_403,N_9963,N_9934);
nor UO_404 (O_404,N_9905,N_9975);
nor UO_405 (O_405,N_9931,N_9920);
and UO_406 (O_406,N_9965,N_9938);
or UO_407 (O_407,N_9962,N_9919);
and UO_408 (O_408,N_9926,N_9971);
nor UO_409 (O_409,N_9932,N_9936);
or UO_410 (O_410,N_9940,N_9930);
or UO_411 (O_411,N_9941,N_9960);
and UO_412 (O_412,N_9908,N_9956);
or UO_413 (O_413,N_9905,N_9954);
or UO_414 (O_414,N_9940,N_9985);
and UO_415 (O_415,N_9941,N_9958);
or UO_416 (O_416,N_9968,N_9997);
nand UO_417 (O_417,N_9908,N_9934);
or UO_418 (O_418,N_9947,N_9938);
and UO_419 (O_419,N_9997,N_9914);
or UO_420 (O_420,N_9974,N_9999);
xnor UO_421 (O_421,N_9967,N_9928);
and UO_422 (O_422,N_9978,N_9907);
or UO_423 (O_423,N_9973,N_9960);
or UO_424 (O_424,N_9963,N_9981);
or UO_425 (O_425,N_9984,N_9937);
nand UO_426 (O_426,N_9958,N_9924);
or UO_427 (O_427,N_9904,N_9905);
and UO_428 (O_428,N_9979,N_9903);
xor UO_429 (O_429,N_9991,N_9944);
or UO_430 (O_430,N_9966,N_9985);
and UO_431 (O_431,N_9987,N_9997);
nor UO_432 (O_432,N_9913,N_9988);
nand UO_433 (O_433,N_9988,N_9923);
or UO_434 (O_434,N_9942,N_9925);
or UO_435 (O_435,N_9942,N_9990);
nand UO_436 (O_436,N_9932,N_9935);
or UO_437 (O_437,N_9946,N_9907);
nor UO_438 (O_438,N_9963,N_9997);
or UO_439 (O_439,N_9964,N_9918);
xnor UO_440 (O_440,N_9905,N_9976);
nand UO_441 (O_441,N_9926,N_9906);
xor UO_442 (O_442,N_9941,N_9952);
or UO_443 (O_443,N_9993,N_9988);
or UO_444 (O_444,N_9903,N_9927);
or UO_445 (O_445,N_9993,N_9953);
nor UO_446 (O_446,N_9933,N_9975);
and UO_447 (O_447,N_9910,N_9977);
or UO_448 (O_448,N_9911,N_9999);
and UO_449 (O_449,N_9977,N_9979);
or UO_450 (O_450,N_9916,N_9929);
nor UO_451 (O_451,N_9990,N_9928);
and UO_452 (O_452,N_9977,N_9954);
or UO_453 (O_453,N_9914,N_9998);
nor UO_454 (O_454,N_9902,N_9931);
nor UO_455 (O_455,N_9907,N_9936);
nor UO_456 (O_456,N_9906,N_9953);
and UO_457 (O_457,N_9961,N_9964);
nor UO_458 (O_458,N_9925,N_9998);
and UO_459 (O_459,N_9967,N_9931);
xor UO_460 (O_460,N_9955,N_9928);
and UO_461 (O_461,N_9907,N_9904);
nand UO_462 (O_462,N_9940,N_9990);
or UO_463 (O_463,N_9994,N_9952);
and UO_464 (O_464,N_9945,N_9919);
nor UO_465 (O_465,N_9917,N_9956);
nor UO_466 (O_466,N_9910,N_9923);
nand UO_467 (O_467,N_9952,N_9939);
xnor UO_468 (O_468,N_9937,N_9905);
and UO_469 (O_469,N_9999,N_9985);
or UO_470 (O_470,N_9987,N_9991);
nor UO_471 (O_471,N_9913,N_9909);
xor UO_472 (O_472,N_9927,N_9909);
and UO_473 (O_473,N_9925,N_9914);
nand UO_474 (O_474,N_9990,N_9960);
or UO_475 (O_475,N_9919,N_9952);
or UO_476 (O_476,N_9920,N_9985);
or UO_477 (O_477,N_9953,N_9905);
nor UO_478 (O_478,N_9983,N_9924);
or UO_479 (O_479,N_9910,N_9978);
xnor UO_480 (O_480,N_9994,N_9978);
and UO_481 (O_481,N_9942,N_9989);
nand UO_482 (O_482,N_9925,N_9908);
and UO_483 (O_483,N_9917,N_9981);
and UO_484 (O_484,N_9952,N_9977);
nand UO_485 (O_485,N_9987,N_9955);
nor UO_486 (O_486,N_9932,N_9965);
nor UO_487 (O_487,N_9944,N_9990);
or UO_488 (O_488,N_9925,N_9986);
nor UO_489 (O_489,N_9924,N_9999);
and UO_490 (O_490,N_9970,N_9936);
and UO_491 (O_491,N_9975,N_9957);
nor UO_492 (O_492,N_9982,N_9989);
nor UO_493 (O_493,N_9968,N_9980);
nor UO_494 (O_494,N_9961,N_9913);
and UO_495 (O_495,N_9951,N_9943);
nand UO_496 (O_496,N_9960,N_9981);
nand UO_497 (O_497,N_9945,N_9980);
xnor UO_498 (O_498,N_9934,N_9956);
nand UO_499 (O_499,N_9970,N_9960);
nand UO_500 (O_500,N_9900,N_9932);
and UO_501 (O_501,N_9905,N_9959);
nand UO_502 (O_502,N_9926,N_9915);
and UO_503 (O_503,N_9974,N_9908);
or UO_504 (O_504,N_9922,N_9999);
or UO_505 (O_505,N_9928,N_9914);
and UO_506 (O_506,N_9916,N_9902);
or UO_507 (O_507,N_9939,N_9967);
and UO_508 (O_508,N_9926,N_9982);
and UO_509 (O_509,N_9951,N_9990);
and UO_510 (O_510,N_9968,N_9938);
xor UO_511 (O_511,N_9928,N_9988);
nor UO_512 (O_512,N_9909,N_9945);
or UO_513 (O_513,N_9993,N_9945);
or UO_514 (O_514,N_9982,N_9936);
xor UO_515 (O_515,N_9938,N_9915);
nor UO_516 (O_516,N_9991,N_9989);
or UO_517 (O_517,N_9937,N_9910);
or UO_518 (O_518,N_9908,N_9988);
and UO_519 (O_519,N_9978,N_9967);
nor UO_520 (O_520,N_9987,N_9995);
nor UO_521 (O_521,N_9965,N_9928);
nor UO_522 (O_522,N_9930,N_9948);
nand UO_523 (O_523,N_9934,N_9957);
nor UO_524 (O_524,N_9977,N_9929);
nand UO_525 (O_525,N_9957,N_9939);
xnor UO_526 (O_526,N_9980,N_9900);
and UO_527 (O_527,N_9945,N_9963);
and UO_528 (O_528,N_9924,N_9970);
nor UO_529 (O_529,N_9961,N_9967);
nor UO_530 (O_530,N_9997,N_9994);
and UO_531 (O_531,N_9917,N_9983);
xor UO_532 (O_532,N_9941,N_9949);
or UO_533 (O_533,N_9948,N_9958);
or UO_534 (O_534,N_9972,N_9928);
xor UO_535 (O_535,N_9965,N_9962);
nand UO_536 (O_536,N_9993,N_9925);
nand UO_537 (O_537,N_9936,N_9999);
and UO_538 (O_538,N_9988,N_9934);
nand UO_539 (O_539,N_9975,N_9916);
nor UO_540 (O_540,N_9964,N_9939);
or UO_541 (O_541,N_9995,N_9956);
nor UO_542 (O_542,N_9931,N_9957);
nand UO_543 (O_543,N_9904,N_9927);
nand UO_544 (O_544,N_9935,N_9925);
nand UO_545 (O_545,N_9970,N_9976);
and UO_546 (O_546,N_9996,N_9925);
or UO_547 (O_547,N_9940,N_9914);
nor UO_548 (O_548,N_9971,N_9930);
or UO_549 (O_549,N_9928,N_9971);
and UO_550 (O_550,N_9922,N_9980);
and UO_551 (O_551,N_9981,N_9945);
and UO_552 (O_552,N_9927,N_9957);
or UO_553 (O_553,N_9910,N_9997);
xor UO_554 (O_554,N_9941,N_9957);
nand UO_555 (O_555,N_9972,N_9991);
and UO_556 (O_556,N_9912,N_9930);
or UO_557 (O_557,N_9975,N_9953);
and UO_558 (O_558,N_9982,N_9942);
nand UO_559 (O_559,N_9926,N_9984);
nor UO_560 (O_560,N_9941,N_9997);
or UO_561 (O_561,N_9958,N_9930);
and UO_562 (O_562,N_9979,N_9974);
nand UO_563 (O_563,N_9910,N_9980);
nor UO_564 (O_564,N_9938,N_9984);
or UO_565 (O_565,N_9919,N_9968);
nor UO_566 (O_566,N_9964,N_9992);
nor UO_567 (O_567,N_9986,N_9907);
nand UO_568 (O_568,N_9902,N_9998);
nand UO_569 (O_569,N_9942,N_9939);
nand UO_570 (O_570,N_9948,N_9961);
or UO_571 (O_571,N_9954,N_9950);
nor UO_572 (O_572,N_9969,N_9936);
and UO_573 (O_573,N_9951,N_9968);
nor UO_574 (O_574,N_9920,N_9934);
nand UO_575 (O_575,N_9994,N_9901);
nor UO_576 (O_576,N_9957,N_9970);
nand UO_577 (O_577,N_9909,N_9971);
or UO_578 (O_578,N_9962,N_9989);
nand UO_579 (O_579,N_9939,N_9956);
or UO_580 (O_580,N_9983,N_9919);
nand UO_581 (O_581,N_9934,N_9948);
nor UO_582 (O_582,N_9900,N_9963);
nand UO_583 (O_583,N_9956,N_9972);
and UO_584 (O_584,N_9994,N_9940);
and UO_585 (O_585,N_9908,N_9964);
nor UO_586 (O_586,N_9982,N_9968);
or UO_587 (O_587,N_9900,N_9924);
nor UO_588 (O_588,N_9930,N_9970);
or UO_589 (O_589,N_9945,N_9914);
or UO_590 (O_590,N_9952,N_9943);
xnor UO_591 (O_591,N_9939,N_9947);
or UO_592 (O_592,N_9900,N_9941);
xnor UO_593 (O_593,N_9986,N_9908);
nand UO_594 (O_594,N_9962,N_9956);
nand UO_595 (O_595,N_9926,N_9916);
xnor UO_596 (O_596,N_9928,N_9935);
nor UO_597 (O_597,N_9936,N_9955);
and UO_598 (O_598,N_9950,N_9974);
and UO_599 (O_599,N_9916,N_9935);
nor UO_600 (O_600,N_9944,N_9941);
or UO_601 (O_601,N_9921,N_9970);
or UO_602 (O_602,N_9943,N_9995);
nand UO_603 (O_603,N_9922,N_9929);
nor UO_604 (O_604,N_9928,N_9997);
nand UO_605 (O_605,N_9912,N_9961);
and UO_606 (O_606,N_9980,N_9915);
xor UO_607 (O_607,N_9910,N_9962);
nor UO_608 (O_608,N_9976,N_9987);
or UO_609 (O_609,N_9953,N_9942);
nand UO_610 (O_610,N_9994,N_9936);
nor UO_611 (O_611,N_9994,N_9965);
nor UO_612 (O_612,N_9956,N_9987);
and UO_613 (O_613,N_9911,N_9943);
xor UO_614 (O_614,N_9943,N_9919);
and UO_615 (O_615,N_9961,N_9986);
nor UO_616 (O_616,N_9900,N_9977);
and UO_617 (O_617,N_9991,N_9992);
nor UO_618 (O_618,N_9905,N_9929);
or UO_619 (O_619,N_9986,N_9914);
nor UO_620 (O_620,N_9972,N_9967);
or UO_621 (O_621,N_9901,N_9996);
nand UO_622 (O_622,N_9911,N_9990);
nand UO_623 (O_623,N_9902,N_9951);
nand UO_624 (O_624,N_9938,N_9921);
nor UO_625 (O_625,N_9978,N_9927);
and UO_626 (O_626,N_9942,N_9924);
nor UO_627 (O_627,N_9960,N_9976);
nor UO_628 (O_628,N_9988,N_9977);
or UO_629 (O_629,N_9975,N_9965);
nor UO_630 (O_630,N_9948,N_9942);
nor UO_631 (O_631,N_9983,N_9901);
nand UO_632 (O_632,N_9941,N_9991);
or UO_633 (O_633,N_9983,N_9977);
or UO_634 (O_634,N_9954,N_9982);
nor UO_635 (O_635,N_9989,N_9975);
nand UO_636 (O_636,N_9952,N_9968);
nor UO_637 (O_637,N_9999,N_9975);
nor UO_638 (O_638,N_9971,N_9956);
or UO_639 (O_639,N_9941,N_9998);
or UO_640 (O_640,N_9953,N_9963);
and UO_641 (O_641,N_9950,N_9981);
nand UO_642 (O_642,N_9912,N_9993);
or UO_643 (O_643,N_9916,N_9951);
nor UO_644 (O_644,N_9988,N_9932);
and UO_645 (O_645,N_9918,N_9906);
nand UO_646 (O_646,N_9933,N_9934);
xor UO_647 (O_647,N_9981,N_9991);
nor UO_648 (O_648,N_9919,N_9958);
nand UO_649 (O_649,N_9971,N_9953);
nand UO_650 (O_650,N_9974,N_9900);
or UO_651 (O_651,N_9918,N_9903);
nand UO_652 (O_652,N_9991,N_9913);
and UO_653 (O_653,N_9903,N_9924);
xor UO_654 (O_654,N_9998,N_9984);
or UO_655 (O_655,N_9943,N_9999);
or UO_656 (O_656,N_9993,N_9922);
nor UO_657 (O_657,N_9954,N_9994);
and UO_658 (O_658,N_9940,N_9924);
or UO_659 (O_659,N_9983,N_9997);
nand UO_660 (O_660,N_9902,N_9904);
nor UO_661 (O_661,N_9971,N_9984);
and UO_662 (O_662,N_9925,N_9959);
xor UO_663 (O_663,N_9969,N_9956);
nand UO_664 (O_664,N_9940,N_9954);
xor UO_665 (O_665,N_9935,N_9967);
xnor UO_666 (O_666,N_9975,N_9955);
nand UO_667 (O_667,N_9922,N_9951);
nand UO_668 (O_668,N_9921,N_9947);
and UO_669 (O_669,N_9982,N_9905);
xor UO_670 (O_670,N_9984,N_9949);
or UO_671 (O_671,N_9956,N_9906);
nor UO_672 (O_672,N_9963,N_9980);
nor UO_673 (O_673,N_9951,N_9920);
or UO_674 (O_674,N_9945,N_9942);
xnor UO_675 (O_675,N_9946,N_9905);
nand UO_676 (O_676,N_9971,N_9923);
xnor UO_677 (O_677,N_9914,N_9973);
or UO_678 (O_678,N_9969,N_9931);
or UO_679 (O_679,N_9996,N_9957);
nand UO_680 (O_680,N_9994,N_9921);
or UO_681 (O_681,N_9990,N_9980);
and UO_682 (O_682,N_9987,N_9932);
or UO_683 (O_683,N_9994,N_9975);
or UO_684 (O_684,N_9988,N_9980);
nor UO_685 (O_685,N_9939,N_9980);
and UO_686 (O_686,N_9932,N_9933);
nor UO_687 (O_687,N_9933,N_9905);
or UO_688 (O_688,N_9999,N_9959);
xnor UO_689 (O_689,N_9915,N_9984);
or UO_690 (O_690,N_9929,N_9913);
or UO_691 (O_691,N_9988,N_9940);
nor UO_692 (O_692,N_9964,N_9953);
or UO_693 (O_693,N_9982,N_9944);
nor UO_694 (O_694,N_9911,N_9925);
nand UO_695 (O_695,N_9902,N_9974);
nor UO_696 (O_696,N_9964,N_9944);
nand UO_697 (O_697,N_9983,N_9985);
or UO_698 (O_698,N_9942,N_9913);
or UO_699 (O_699,N_9995,N_9979);
nor UO_700 (O_700,N_9974,N_9990);
nand UO_701 (O_701,N_9985,N_9980);
nor UO_702 (O_702,N_9954,N_9964);
nor UO_703 (O_703,N_9923,N_9901);
or UO_704 (O_704,N_9945,N_9991);
nor UO_705 (O_705,N_9935,N_9993);
and UO_706 (O_706,N_9971,N_9964);
or UO_707 (O_707,N_9972,N_9910);
nor UO_708 (O_708,N_9979,N_9948);
and UO_709 (O_709,N_9996,N_9969);
and UO_710 (O_710,N_9923,N_9951);
or UO_711 (O_711,N_9921,N_9977);
nor UO_712 (O_712,N_9991,N_9935);
or UO_713 (O_713,N_9951,N_9970);
nor UO_714 (O_714,N_9914,N_9964);
and UO_715 (O_715,N_9933,N_9954);
or UO_716 (O_716,N_9933,N_9910);
xor UO_717 (O_717,N_9940,N_9951);
and UO_718 (O_718,N_9982,N_9979);
xnor UO_719 (O_719,N_9957,N_9906);
nand UO_720 (O_720,N_9995,N_9942);
nor UO_721 (O_721,N_9985,N_9931);
or UO_722 (O_722,N_9901,N_9919);
nor UO_723 (O_723,N_9978,N_9913);
nor UO_724 (O_724,N_9969,N_9986);
or UO_725 (O_725,N_9991,N_9918);
or UO_726 (O_726,N_9931,N_9935);
or UO_727 (O_727,N_9936,N_9941);
nor UO_728 (O_728,N_9959,N_9968);
and UO_729 (O_729,N_9933,N_9971);
nand UO_730 (O_730,N_9937,N_9973);
xnor UO_731 (O_731,N_9976,N_9952);
nor UO_732 (O_732,N_9935,N_9981);
and UO_733 (O_733,N_9971,N_9913);
nand UO_734 (O_734,N_9958,N_9961);
or UO_735 (O_735,N_9948,N_9936);
or UO_736 (O_736,N_9999,N_9942);
xnor UO_737 (O_737,N_9957,N_9995);
nand UO_738 (O_738,N_9947,N_9953);
nand UO_739 (O_739,N_9992,N_9983);
and UO_740 (O_740,N_9912,N_9997);
and UO_741 (O_741,N_9960,N_9907);
nand UO_742 (O_742,N_9922,N_9985);
nand UO_743 (O_743,N_9959,N_9965);
and UO_744 (O_744,N_9902,N_9964);
nand UO_745 (O_745,N_9993,N_9946);
nor UO_746 (O_746,N_9997,N_9998);
nand UO_747 (O_747,N_9920,N_9945);
and UO_748 (O_748,N_9922,N_9983);
or UO_749 (O_749,N_9916,N_9942);
nor UO_750 (O_750,N_9900,N_9957);
or UO_751 (O_751,N_9926,N_9957);
nand UO_752 (O_752,N_9957,N_9925);
xor UO_753 (O_753,N_9956,N_9965);
or UO_754 (O_754,N_9978,N_9939);
and UO_755 (O_755,N_9907,N_9905);
or UO_756 (O_756,N_9954,N_9904);
and UO_757 (O_757,N_9931,N_9998);
and UO_758 (O_758,N_9987,N_9999);
xor UO_759 (O_759,N_9936,N_9974);
or UO_760 (O_760,N_9937,N_9929);
nor UO_761 (O_761,N_9957,N_9986);
nor UO_762 (O_762,N_9915,N_9934);
and UO_763 (O_763,N_9935,N_9945);
and UO_764 (O_764,N_9915,N_9914);
and UO_765 (O_765,N_9997,N_9917);
or UO_766 (O_766,N_9964,N_9975);
or UO_767 (O_767,N_9930,N_9904);
or UO_768 (O_768,N_9910,N_9913);
nor UO_769 (O_769,N_9949,N_9931);
or UO_770 (O_770,N_9954,N_9967);
and UO_771 (O_771,N_9988,N_9924);
nand UO_772 (O_772,N_9921,N_9993);
nand UO_773 (O_773,N_9931,N_9906);
nand UO_774 (O_774,N_9947,N_9943);
nor UO_775 (O_775,N_9962,N_9916);
or UO_776 (O_776,N_9957,N_9999);
xor UO_777 (O_777,N_9969,N_9992);
nor UO_778 (O_778,N_9996,N_9917);
and UO_779 (O_779,N_9987,N_9913);
nand UO_780 (O_780,N_9978,N_9904);
and UO_781 (O_781,N_9906,N_9988);
and UO_782 (O_782,N_9990,N_9932);
xnor UO_783 (O_783,N_9904,N_9970);
nand UO_784 (O_784,N_9949,N_9962);
and UO_785 (O_785,N_9920,N_9961);
and UO_786 (O_786,N_9912,N_9954);
nor UO_787 (O_787,N_9900,N_9930);
or UO_788 (O_788,N_9914,N_9957);
or UO_789 (O_789,N_9944,N_9932);
and UO_790 (O_790,N_9923,N_9921);
nand UO_791 (O_791,N_9922,N_9965);
or UO_792 (O_792,N_9919,N_9928);
and UO_793 (O_793,N_9992,N_9933);
and UO_794 (O_794,N_9930,N_9995);
or UO_795 (O_795,N_9971,N_9994);
xnor UO_796 (O_796,N_9958,N_9906);
nand UO_797 (O_797,N_9945,N_9965);
xnor UO_798 (O_798,N_9969,N_9938);
or UO_799 (O_799,N_9903,N_9935);
nor UO_800 (O_800,N_9924,N_9936);
and UO_801 (O_801,N_9964,N_9980);
xor UO_802 (O_802,N_9933,N_9938);
xor UO_803 (O_803,N_9912,N_9924);
and UO_804 (O_804,N_9967,N_9992);
nor UO_805 (O_805,N_9994,N_9903);
and UO_806 (O_806,N_9918,N_9940);
nand UO_807 (O_807,N_9953,N_9945);
nor UO_808 (O_808,N_9992,N_9932);
xnor UO_809 (O_809,N_9956,N_9923);
or UO_810 (O_810,N_9939,N_9910);
nor UO_811 (O_811,N_9945,N_9900);
xor UO_812 (O_812,N_9954,N_9946);
nor UO_813 (O_813,N_9930,N_9907);
and UO_814 (O_814,N_9998,N_9926);
or UO_815 (O_815,N_9900,N_9968);
and UO_816 (O_816,N_9993,N_9991);
xnor UO_817 (O_817,N_9966,N_9921);
xnor UO_818 (O_818,N_9933,N_9917);
nor UO_819 (O_819,N_9922,N_9966);
nor UO_820 (O_820,N_9962,N_9972);
nor UO_821 (O_821,N_9918,N_9958);
nor UO_822 (O_822,N_9950,N_9963);
nand UO_823 (O_823,N_9957,N_9984);
and UO_824 (O_824,N_9927,N_9946);
nand UO_825 (O_825,N_9983,N_9932);
nand UO_826 (O_826,N_9971,N_9952);
or UO_827 (O_827,N_9939,N_9902);
or UO_828 (O_828,N_9958,N_9973);
nor UO_829 (O_829,N_9967,N_9958);
and UO_830 (O_830,N_9902,N_9976);
nor UO_831 (O_831,N_9916,N_9901);
nand UO_832 (O_832,N_9914,N_9954);
and UO_833 (O_833,N_9964,N_9910);
and UO_834 (O_834,N_9911,N_9908);
and UO_835 (O_835,N_9954,N_9916);
xor UO_836 (O_836,N_9943,N_9996);
xor UO_837 (O_837,N_9975,N_9971);
nand UO_838 (O_838,N_9982,N_9916);
and UO_839 (O_839,N_9945,N_9936);
nor UO_840 (O_840,N_9921,N_9949);
xnor UO_841 (O_841,N_9965,N_9978);
and UO_842 (O_842,N_9903,N_9913);
and UO_843 (O_843,N_9983,N_9911);
nor UO_844 (O_844,N_9964,N_9911);
and UO_845 (O_845,N_9950,N_9916);
xnor UO_846 (O_846,N_9982,N_9946);
nor UO_847 (O_847,N_9996,N_9950);
nand UO_848 (O_848,N_9997,N_9909);
and UO_849 (O_849,N_9935,N_9917);
and UO_850 (O_850,N_9950,N_9969);
nand UO_851 (O_851,N_9924,N_9922);
xnor UO_852 (O_852,N_9910,N_9971);
or UO_853 (O_853,N_9973,N_9978);
and UO_854 (O_854,N_9944,N_9911);
nor UO_855 (O_855,N_9923,N_9947);
or UO_856 (O_856,N_9970,N_9961);
xor UO_857 (O_857,N_9995,N_9918);
nor UO_858 (O_858,N_9926,N_9907);
nand UO_859 (O_859,N_9961,N_9950);
nand UO_860 (O_860,N_9930,N_9996);
nor UO_861 (O_861,N_9973,N_9953);
and UO_862 (O_862,N_9975,N_9942);
nand UO_863 (O_863,N_9980,N_9951);
nor UO_864 (O_864,N_9948,N_9994);
and UO_865 (O_865,N_9931,N_9937);
nor UO_866 (O_866,N_9971,N_9929);
nand UO_867 (O_867,N_9987,N_9963);
nand UO_868 (O_868,N_9983,N_9920);
nand UO_869 (O_869,N_9968,N_9956);
nor UO_870 (O_870,N_9937,N_9960);
nand UO_871 (O_871,N_9931,N_9963);
or UO_872 (O_872,N_9948,N_9944);
xor UO_873 (O_873,N_9940,N_9970);
xnor UO_874 (O_874,N_9979,N_9989);
nand UO_875 (O_875,N_9926,N_9985);
and UO_876 (O_876,N_9955,N_9925);
xnor UO_877 (O_877,N_9957,N_9973);
and UO_878 (O_878,N_9955,N_9957);
xor UO_879 (O_879,N_9934,N_9992);
nor UO_880 (O_880,N_9961,N_9976);
nand UO_881 (O_881,N_9972,N_9949);
or UO_882 (O_882,N_9903,N_9933);
or UO_883 (O_883,N_9931,N_9908);
xor UO_884 (O_884,N_9995,N_9920);
or UO_885 (O_885,N_9962,N_9969);
nand UO_886 (O_886,N_9900,N_9927);
nor UO_887 (O_887,N_9961,N_9947);
xor UO_888 (O_888,N_9925,N_9983);
nor UO_889 (O_889,N_9908,N_9994);
nand UO_890 (O_890,N_9959,N_9921);
and UO_891 (O_891,N_9954,N_9958);
and UO_892 (O_892,N_9902,N_9929);
or UO_893 (O_893,N_9958,N_9975);
and UO_894 (O_894,N_9983,N_9913);
and UO_895 (O_895,N_9915,N_9940);
nand UO_896 (O_896,N_9913,N_9927);
xor UO_897 (O_897,N_9951,N_9924);
nor UO_898 (O_898,N_9943,N_9956);
and UO_899 (O_899,N_9908,N_9947);
nand UO_900 (O_900,N_9969,N_9911);
or UO_901 (O_901,N_9946,N_9975);
nand UO_902 (O_902,N_9923,N_9934);
xnor UO_903 (O_903,N_9995,N_9908);
nand UO_904 (O_904,N_9972,N_9942);
nand UO_905 (O_905,N_9901,N_9959);
nor UO_906 (O_906,N_9900,N_9943);
and UO_907 (O_907,N_9919,N_9956);
or UO_908 (O_908,N_9923,N_9957);
nand UO_909 (O_909,N_9954,N_9951);
and UO_910 (O_910,N_9910,N_9945);
nor UO_911 (O_911,N_9940,N_9942);
and UO_912 (O_912,N_9981,N_9926);
and UO_913 (O_913,N_9997,N_9903);
or UO_914 (O_914,N_9972,N_9995);
and UO_915 (O_915,N_9959,N_9993);
and UO_916 (O_916,N_9905,N_9903);
and UO_917 (O_917,N_9993,N_9994);
and UO_918 (O_918,N_9909,N_9967);
nand UO_919 (O_919,N_9987,N_9901);
or UO_920 (O_920,N_9932,N_9949);
nor UO_921 (O_921,N_9928,N_9977);
or UO_922 (O_922,N_9923,N_9985);
nand UO_923 (O_923,N_9918,N_9926);
and UO_924 (O_924,N_9950,N_9994);
nand UO_925 (O_925,N_9968,N_9995);
or UO_926 (O_926,N_9909,N_9904);
xnor UO_927 (O_927,N_9935,N_9955);
nand UO_928 (O_928,N_9966,N_9939);
nand UO_929 (O_929,N_9965,N_9948);
nand UO_930 (O_930,N_9937,N_9928);
nand UO_931 (O_931,N_9926,N_9905);
or UO_932 (O_932,N_9926,N_9980);
nand UO_933 (O_933,N_9933,N_9965);
nor UO_934 (O_934,N_9927,N_9974);
nor UO_935 (O_935,N_9949,N_9933);
nand UO_936 (O_936,N_9963,N_9914);
nor UO_937 (O_937,N_9968,N_9930);
or UO_938 (O_938,N_9916,N_9915);
and UO_939 (O_939,N_9923,N_9918);
and UO_940 (O_940,N_9995,N_9985);
nor UO_941 (O_941,N_9946,N_9969);
and UO_942 (O_942,N_9968,N_9949);
and UO_943 (O_943,N_9917,N_9961);
or UO_944 (O_944,N_9919,N_9921);
nand UO_945 (O_945,N_9959,N_9954);
or UO_946 (O_946,N_9904,N_9991);
nand UO_947 (O_947,N_9949,N_9975);
or UO_948 (O_948,N_9962,N_9921);
and UO_949 (O_949,N_9958,N_9962);
xnor UO_950 (O_950,N_9994,N_9985);
or UO_951 (O_951,N_9921,N_9901);
or UO_952 (O_952,N_9974,N_9918);
nor UO_953 (O_953,N_9925,N_9995);
nor UO_954 (O_954,N_9947,N_9917);
nor UO_955 (O_955,N_9942,N_9976);
or UO_956 (O_956,N_9978,N_9966);
and UO_957 (O_957,N_9992,N_9948);
or UO_958 (O_958,N_9984,N_9954);
or UO_959 (O_959,N_9909,N_9975);
and UO_960 (O_960,N_9947,N_9905);
or UO_961 (O_961,N_9945,N_9959);
nor UO_962 (O_962,N_9991,N_9949);
or UO_963 (O_963,N_9973,N_9920);
or UO_964 (O_964,N_9955,N_9911);
and UO_965 (O_965,N_9937,N_9999);
or UO_966 (O_966,N_9932,N_9969);
and UO_967 (O_967,N_9918,N_9954);
nand UO_968 (O_968,N_9987,N_9972);
xnor UO_969 (O_969,N_9962,N_9931);
or UO_970 (O_970,N_9949,N_9939);
nand UO_971 (O_971,N_9919,N_9961);
nor UO_972 (O_972,N_9970,N_9925);
nor UO_973 (O_973,N_9977,N_9984);
or UO_974 (O_974,N_9942,N_9915);
nand UO_975 (O_975,N_9917,N_9902);
nand UO_976 (O_976,N_9904,N_9969);
nor UO_977 (O_977,N_9965,N_9999);
xor UO_978 (O_978,N_9932,N_9912);
and UO_979 (O_979,N_9930,N_9989);
nor UO_980 (O_980,N_9983,N_9981);
and UO_981 (O_981,N_9988,N_9901);
nor UO_982 (O_982,N_9941,N_9922);
nand UO_983 (O_983,N_9929,N_9936);
nand UO_984 (O_984,N_9961,N_9924);
nand UO_985 (O_985,N_9951,N_9919);
or UO_986 (O_986,N_9917,N_9907);
or UO_987 (O_987,N_9968,N_9969);
nand UO_988 (O_988,N_9907,N_9968);
nand UO_989 (O_989,N_9908,N_9953);
and UO_990 (O_990,N_9939,N_9955);
nor UO_991 (O_991,N_9991,N_9930);
and UO_992 (O_992,N_9935,N_9979);
or UO_993 (O_993,N_9929,N_9966);
xnor UO_994 (O_994,N_9912,N_9955);
or UO_995 (O_995,N_9921,N_9912);
nor UO_996 (O_996,N_9937,N_9922);
and UO_997 (O_997,N_9921,N_9934);
nor UO_998 (O_998,N_9981,N_9995);
nor UO_999 (O_999,N_9996,N_9944);
nand UO_1000 (O_1000,N_9952,N_9965);
nand UO_1001 (O_1001,N_9939,N_9909);
and UO_1002 (O_1002,N_9953,N_9949);
and UO_1003 (O_1003,N_9919,N_9967);
or UO_1004 (O_1004,N_9934,N_9902);
nand UO_1005 (O_1005,N_9937,N_9944);
and UO_1006 (O_1006,N_9958,N_9969);
nor UO_1007 (O_1007,N_9955,N_9996);
and UO_1008 (O_1008,N_9931,N_9971);
and UO_1009 (O_1009,N_9967,N_9925);
nand UO_1010 (O_1010,N_9921,N_9933);
nor UO_1011 (O_1011,N_9954,N_9915);
nor UO_1012 (O_1012,N_9959,N_9933);
and UO_1013 (O_1013,N_9999,N_9984);
and UO_1014 (O_1014,N_9917,N_9966);
nor UO_1015 (O_1015,N_9933,N_9969);
and UO_1016 (O_1016,N_9981,N_9921);
nor UO_1017 (O_1017,N_9983,N_9951);
nand UO_1018 (O_1018,N_9971,N_9947);
and UO_1019 (O_1019,N_9908,N_9924);
xor UO_1020 (O_1020,N_9994,N_9935);
and UO_1021 (O_1021,N_9968,N_9928);
xor UO_1022 (O_1022,N_9999,N_9983);
nand UO_1023 (O_1023,N_9909,N_9926);
nand UO_1024 (O_1024,N_9933,N_9904);
and UO_1025 (O_1025,N_9936,N_9989);
nand UO_1026 (O_1026,N_9994,N_9933);
nand UO_1027 (O_1027,N_9927,N_9992);
and UO_1028 (O_1028,N_9927,N_9902);
nor UO_1029 (O_1029,N_9980,N_9942);
and UO_1030 (O_1030,N_9920,N_9914);
nand UO_1031 (O_1031,N_9968,N_9941);
or UO_1032 (O_1032,N_9912,N_9944);
nand UO_1033 (O_1033,N_9954,N_9902);
nor UO_1034 (O_1034,N_9973,N_9924);
xnor UO_1035 (O_1035,N_9924,N_9931);
and UO_1036 (O_1036,N_9913,N_9990);
or UO_1037 (O_1037,N_9949,N_9990);
xor UO_1038 (O_1038,N_9968,N_9993);
or UO_1039 (O_1039,N_9961,N_9960);
nor UO_1040 (O_1040,N_9900,N_9921);
nand UO_1041 (O_1041,N_9961,N_9935);
or UO_1042 (O_1042,N_9915,N_9955);
nand UO_1043 (O_1043,N_9965,N_9986);
and UO_1044 (O_1044,N_9930,N_9967);
or UO_1045 (O_1045,N_9959,N_9981);
and UO_1046 (O_1046,N_9913,N_9945);
xnor UO_1047 (O_1047,N_9946,N_9914);
or UO_1048 (O_1048,N_9964,N_9924);
and UO_1049 (O_1049,N_9976,N_9937);
nor UO_1050 (O_1050,N_9929,N_9943);
nor UO_1051 (O_1051,N_9963,N_9928);
or UO_1052 (O_1052,N_9955,N_9981);
and UO_1053 (O_1053,N_9982,N_9980);
and UO_1054 (O_1054,N_9954,N_9957);
or UO_1055 (O_1055,N_9922,N_9948);
nand UO_1056 (O_1056,N_9999,N_9991);
and UO_1057 (O_1057,N_9910,N_9983);
xnor UO_1058 (O_1058,N_9906,N_9923);
or UO_1059 (O_1059,N_9970,N_9989);
and UO_1060 (O_1060,N_9970,N_9965);
nor UO_1061 (O_1061,N_9941,N_9924);
and UO_1062 (O_1062,N_9984,N_9916);
nand UO_1063 (O_1063,N_9966,N_9949);
nor UO_1064 (O_1064,N_9908,N_9913);
or UO_1065 (O_1065,N_9913,N_9992);
or UO_1066 (O_1066,N_9964,N_9974);
nand UO_1067 (O_1067,N_9912,N_9975);
nor UO_1068 (O_1068,N_9937,N_9916);
and UO_1069 (O_1069,N_9969,N_9966);
nand UO_1070 (O_1070,N_9934,N_9970);
xnor UO_1071 (O_1071,N_9945,N_9992);
nor UO_1072 (O_1072,N_9983,N_9973);
and UO_1073 (O_1073,N_9922,N_9947);
nand UO_1074 (O_1074,N_9965,N_9998);
or UO_1075 (O_1075,N_9910,N_9905);
nand UO_1076 (O_1076,N_9938,N_9935);
xnor UO_1077 (O_1077,N_9933,N_9940);
nor UO_1078 (O_1078,N_9995,N_9912);
nand UO_1079 (O_1079,N_9916,N_9989);
nand UO_1080 (O_1080,N_9981,N_9927);
and UO_1081 (O_1081,N_9974,N_9917);
or UO_1082 (O_1082,N_9958,N_9946);
nor UO_1083 (O_1083,N_9967,N_9941);
nor UO_1084 (O_1084,N_9923,N_9940);
nor UO_1085 (O_1085,N_9916,N_9986);
or UO_1086 (O_1086,N_9943,N_9989);
nand UO_1087 (O_1087,N_9998,N_9976);
and UO_1088 (O_1088,N_9941,N_9966);
nor UO_1089 (O_1089,N_9965,N_9921);
nand UO_1090 (O_1090,N_9987,N_9921);
or UO_1091 (O_1091,N_9993,N_9914);
and UO_1092 (O_1092,N_9977,N_9949);
nand UO_1093 (O_1093,N_9955,N_9961);
nand UO_1094 (O_1094,N_9931,N_9996);
or UO_1095 (O_1095,N_9980,N_9947);
and UO_1096 (O_1096,N_9994,N_9924);
nand UO_1097 (O_1097,N_9991,N_9916);
nand UO_1098 (O_1098,N_9974,N_9905);
or UO_1099 (O_1099,N_9937,N_9997);
and UO_1100 (O_1100,N_9947,N_9935);
and UO_1101 (O_1101,N_9989,N_9995);
xor UO_1102 (O_1102,N_9940,N_9986);
nand UO_1103 (O_1103,N_9985,N_9989);
xnor UO_1104 (O_1104,N_9910,N_9908);
nor UO_1105 (O_1105,N_9996,N_9961);
or UO_1106 (O_1106,N_9982,N_9995);
nor UO_1107 (O_1107,N_9935,N_9970);
nand UO_1108 (O_1108,N_9984,N_9952);
nor UO_1109 (O_1109,N_9966,N_9911);
nand UO_1110 (O_1110,N_9963,N_9998);
and UO_1111 (O_1111,N_9909,N_9903);
nand UO_1112 (O_1112,N_9982,N_9932);
xor UO_1113 (O_1113,N_9940,N_9937);
nor UO_1114 (O_1114,N_9920,N_9996);
nor UO_1115 (O_1115,N_9974,N_9938);
nand UO_1116 (O_1116,N_9964,N_9982);
xor UO_1117 (O_1117,N_9920,N_9994);
nor UO_1118 (O_1118,N_9965,N_9991);
xor UO_1119 (O_1119,N_9916,N_9966);
nor UO_1120 (O_1120,N_9948,N_9925);
nor UO_1121 (O_1121,N_9903,N_9965);
and UO_1122 (O_1122,N_9926,N_9965);
or UO_1123 (O_1123,N_9940,N_9943);
or UO_1124 (O_1124,N_9997,N_9964);
and UO_1125 (O_1125,N_9957,N_9903);
or UO_1126 (O_1126,N_9908,N_9937);
nor UO_1127 (O_1127,N_9916,N_9987);
and UO_1128 (O_1128,N_9921,N_9972);
nor UO_1129 (O_1129,N_9967,N_9966);
or UO_1130 (O_1130,N_9952,N_9929);
or UO_1131 (O_1131,N_9982,N_9939);
or UO_1132 (O_1132,N_9940,N_9908);
nand UO_1133 (O_1133,N_9972,N_9952);
nand UO_1134 (O_1134,N_9921,N_9935);
and UO_1135 (O_1135,N_9907,N_9942);
and UO_1136 (O_1136,N_9949,N_9943);
xnor UO_1137 (O_1137,N_9985,N_9906);
and UO_1138 (O_1138,N_9932,N_9948);
and UO_1139 (O_1139,N_9941,N_9906);
nand UO_1140 (O_1140,N_9927,N_9936);
and UO_1141 (O_1141,N_9920,N_9993);
nor UO_1142 (O_1142,N_9957,N_9907);
nor UO_1143 (O_1143,N_9921,N_9992);
nand UO_1144 (O_1144,N_9996,N_9985);
and UO_1145 (O_1145,N_9991,N_9921);
or UO_1146 (O_1146,N_9937,N_9925);
xnor UO_1147 (O_1147,N_9968,N_9957);
nor UO_1148 (O_1148,N_9933,N_9963);
and UO_1149 (O_1149,N_9969,N_9970);
nand UO_1150 (O_1150,N_9981,N_9993);
nor UO_1151 (O_1151,N_9909,N_9936);
nand UO_1152 (O_1152,N_9951,N_9961);
nor UO_1153 (O_1153,N_9957,N_9951);
or UO_1154 (O_1154,N_9943,N_9925);
xnor UO_1155 (O_1155,N_9955,N_9910);
and UO_1156 (O_1156,N_9914,N_9952);
nor UO_1157 (O_1157,N_9955,N_9913);
xnor UO_1158 (O_1158,N_9986,N_9918);
nor UO_1159 (O_1159,N_9944,N_9938);
nand UO_1160 (O_1160,N_9914,N_9936);
and UO_1161 (O_1161,N_9954,N_9921);
nor UO_1162 (O_1162,N_9928,N_9982);
nor UO_1163 (O_1163,N_9968,N_9926);
and UO_1164 (O_1164,N_9943,N_9979);
nand UO_1165 (O_1165,N_9900,N_9998);
nor UO_1166 (O_1166,N_9935,N_9904);
nand UO_1167 (O_1167,N_9927,N_9983);
nor UO_1168 (O_1168,N_9936,N_9981);
and UO_1169 (O_1169,N_9946,N_9956);
nor UO_1170 (O_1170,N_9986,N_9932);
xor UO_1171 (O_1171,N_9998,N_9912);
or UO_1172 (O_1172,N_9990,N_9921);
or UO_1173 (O_1173,N_9997,N_9992);
xor UO_1174 (O_1174,N_9992,N_9982);
or UO_1175 (O_1175,N_9936,N_9938);
nor UO_1176 (O_1176,N_9950,N_9948);
and UO_1177 (O_1177,N_9944,N_9900);
or UO_1178 (O_1178,N_9905,N_9948);
or UO_1179 (O_1179,N_9925,N_9931);
nand UO_1180 (O_1180,N_9959,N_9969);
or UO_1181 (O_1181,N_9946,N_9906);
or UO_1182 (O_1182,N_9908,N_9991);
xor UO_1183 (O_1183,N_9970,N_9954);
and UO_1184 (O_1184,N_9996,N_9914);
and UO_1185 (O_1185,N_9991,N_9997);
nand UO_1186 (O_1186,N_9989,N_9906);
nand UO_1187 (O_1187,N_9927,N_9930);
and UO_1188 (O_1188,N_9919,N_9970);
nand UO_1189 (O_1189,N_9927,N_9963);
and UO_1190 (O_1190,N_9913,N_9986);
and UO_1191 (O_1191,N_9958,N_9994);
nor UO_1192 (O_1192,N_9989,N_9959);
xnor UO_1193 (O_1193,N_9954,N_9952);
nand UO_1194 (O_1194,N_9929,N_9963);
nand UO_1195 (O_1195,N_9944,N_9979);
or UO_1196 (O_1196,N_9986,N_9971);
nor UO_1197 (O_1197,N_9915,N_9975);
nand UO_1198 (O_1198,N_9982,N_9957);
or UO_1199 (O_1199,N_9945,N_9948);
nand UO_1200 (O_1200,N_9933,N_9977);
nor UO_1201 (O_1201,N_9947,N_9906);
xor UO_1202 (O_1202,N_9967,N_9904);
nor UO_1203 (O_1203,N_9990,N_9936);
nor UO_1204 (O_1204,N_9922,N_9940);
nor UO_1205 (O_1205,N_9988,N_9976);
nor UO_1206 (O_1206,N_9977,N_9947);
nand UO_1207 (O_1207,N_9925,N_9990);
nand UO_1208 (O_1208,N_9913,N_9953);
and UO_1209 (O_1209,N_9997,N_9958);
nand UO_1210 (O_1210,N_9912,N_9996);
nor UO_1211 (O_1211,N_9950,N_9932);
nor UO_1212 (O_1212,N_9910,N_9996);
or UO_1213 (O_1213,N_9927,N_9914);
xnor UO_1214 (O_1214,N_9927,N_9948);
nand UO_1215 (O_1215,N_9914,N_9922);
xor UO_1216 (O_1216,N_9959,N_9922);
or UO_1217 (O_1217,N_9943,N_9981);
nand UO_1218 (O_1218,N_9934,N_9985);
and UO_1219 (O_1219,N_9945,N_9929);
or UO_1220 (O_1220,N_9963,N_9954);
or UO_1221 (O_1221,N_9945,N_9975);
xnor UO_1222 (O_1222,N_9902,N_9955);
nand UO_1223 (O_1223,N_9990,N_9947);
nand UO_1224 (O_1224,N_9927,N_9997);
nor UO_1225 (O_1225,N_9941,N_9942);
and UO_1226 (O_1226,N_9911,N_9940);
and UO_1227 (O_1227,N_9932,N_9993);
nor UO_1228 (O_1228,N_9929,N_9991);
nor UO_1229 (O_1229,N_9967,N_9995);
or UO_1230 (O_1230,N_9992,N_9995);
and UO_1231 (O_1231,N_9954,N_9943);
nand UO_1232 (O_1232,N_9948,N_9998);
and UO_1233 (O_1233,N_9952,N_9949);
nor UO_1234 (O_1234,N_9908,N_9906);
xnor UO_1235 (O_1235,N_9992,N_9962);
or UO_1236 (O_1236,N_9932,N_9976);
or UO_1237 (O_1237,N_9976,N_9969);
xnor UO_1238 (O_1238,N_9991,N_9902);
or UO_1239 (O_1239,N_9903,N_9974);
nand UO_1240 (O_1240,N_9955,N_9991);
nand UO_1241 (O_1241,N_9963,N_9992);
nand UO_1242 (O_1242,N_9971,N_9940);
xor UO_1243 (O_1243,N_9985,N_9957);
nand UO_1244 (O_1244,N_9948,N_9969);
and UO_1245 (O_1245,N_9987,N_9980);
and UO_1246 (O_1246,N_9904,N_9921);
and UO_1247 (O_1247,N_9949,N_9964);
or UO_1248 (O_1248,N_9943,N_9923);
or UO_1249 (O_1249,N_9908,N_9909);
and UO_1250 (O_1250,N_9990,N_9919);
nand UO_1251 (O_1251,N_9971,N_9920);
or UO_1252 (O_1252,N_9972,N_9931);
or UO_1253 (O_1253,N_9984,N_9944);
nor UO_1254 (O_1254,N_9943,N_9998);
nor UO_1255 (O_1255,N_9901,N_9956);
or UO_1256 (O_1256,N_9934,N_9962);
nor UO_1257 (O_1257,N_9997,N_9978);
nand UO_1258 (O_1258,N_9987,N_9900);
or UO_1259 (O_1259,N_9900,N_9976);
and UO_1260 (O_1260,N_9912,N_9987);
nand UO_1261 (O_1261,N_9959,N_9988);
nor UO_1262 (O_1262,N_9965,N_9939);
or UO_1263 (O_1263,N_9996,N_9977);
or UO_1264 (O_1264,N_9901,N_9934);
nand UO_1265 (O_1265,N_9921,N_9995);
and UO_1266 (O_1266,N_9941,N_9992);
nand UO_1267 (O_1267,N_9909,N_9972);
nand UO_1268 (O_1268,N_9941,N_9910);
and UO_1269 (O_1269,N_9989,N_9926);
nand UO_1270 (O_1270,N_9951,N_9987);
nand UO_1271 (O_1271,N_9979,N_9968);
and UO_1272 (O_1272,N_9956,N_9970);
nor UO_1273 (O_1273,N_9904,N_9920);
and UO_1274 (O_1274,N_9934,N_9936);
nand UO_1275 (O_1275,N_9902,N_9922);
nand UO_1276 (O_1276,N_9945,N_9915);
nor UO_1277 (O_1277,N_9910,N_9934);
or UO_1278 (O_1278,N_9999,N_9967);
nor UO_1279 (O_1279,N_9981,N_9974);
and UO_1280 (O_1280,N_9938,N_9901);
xor UO_1281 (O_1281,N_9978,N_9975);
or UO_1282 (O_1282,N_9962,N_9943);
nand UO_1283 (O_1283,N_9960,N_9967);
nand UO_1284 (O_1284,N_9975,N_9970);
or UO_1285 (O_1285,N_9918,N_9944);
or UO_1286 (O_1286,N_9928,N_9961);
nor UO_1287 (O_1287,N_9901,N_9912);
nand UO_1288 (O_1288,N_9917,N_9991);
and UO_1289 (O_1289,N_9911,N_9939);
or UO_1290 (O_1290,N_9926,N_9948);
nor UO_1291 (O_1291,N_9944,N_9906);
nand UO_1292 (O_1292,N_9972,N_9905);
and UO_1293 (O_1293,N_9906,N_9961);
nand UO_1294 (O_1294,N_9907,N_9974);
or UO_1295 (O_1295,N_9969,N_9954);
and UO_1296 (O_1296,N_9945,N_9925);
nor UO_1297 (O_1297,N_9959,N_9914);
xnor UO_1298 (O_1298,N_9979,N_9980);
nand UO_1299 (O_1299,N_9926,N_9966);
nor UO_1300 (O_1300,N_9921,N_9964);
and UO_1301 (O_1301,N_9973,N_9911);
nand UO_1302 (O_1302,N_9982,N_9970);
and UO_1303 (O_1303,N_9971,N_9943);
nor UO_1304 (O_1304,N_9947,N_9982);
or UO_1305 (O_1305,N_9990,N_9920);
nand UO_1306 (O_1306,N_9919,N_9994);
or UO_1307 (O_1307,N_9987,N_9909);
xnor UO_1308 (O_1308,N_9943,N_9965);
nand UO_1309 (O_1309,N_9996,N_9989);
or UO_1310 (O_1310,N_9979,N_9916);
or UO_1311 (O_1311,N_9937,N_9950);
or UO_1312 (O_1312,N_9944,N_9913);
nand UO_1313 (O_1313,N_9903,N_9920);
nand UO_1314 (O_1314,N_9941,N_9912);
nor UO_1315 (O_1315,N_9939,N_9990);
nand UO_1316 (O_1316,N_9999,N_9904);
nand UO_1317 (O_1317,N_9913,N_9966);
and UO_1318 (O_1318,N_9950,N_9915);
and UO_1319 (O_1319,N_9993,N_9924);
nand UO_1320 (O_1320,N_9948,N_9977);
nor UO_1321 (O_1321,N_9937,N_9903);
and UO_1322 (O_1322,N_9927,N_9917);
xnor UO_1323 (O_1323,N_9931,N_9929);
xor UO_1324 (O_1324,N_9931,N_9991);
or UO_1325 (O_1325,N_9953,N_9977);
and UO_1326 (O_1326,N_9941,N_9954);
nor UO_1327 (O_1327,N_9957,N_9942);
nand UO_1328 (O_1328,N_9932,N_9903);
xor UO_1329 (O_1329,N_9919,N_9903);
and UO_1330 (O_1330,N_9924,N_9955);
nor UO_1331 (O_1331,N_9909,N_9938);
nor UO_1332 (O_1332,N_9958,N_9980);
or UO_1333 (O_1333,N_9979,N_9966);
nor UO_1334 (O_1334,N_9956,N_9974);
xnor UO_1335 (O_1335,N_9918,N_9911);
nand UO_1336 (O_1336,N_9982,N_9959);
nor UO_1337 (O_1337,N_9980,N_9959);
nor UO_1338 (O_1338,N_9930,N_9922);
and UO_1339 (O_1339,N_9904,N_9961);
nand UO_1340 (O_1340,N_9946,N_9901);
or UO_1341 (O_1341,N_9906,N_9993);
and UO_1342 (O_1342,N_9945,N_9922);
or UO_1343 (O_1343,N_9954,N_9962);
and UO_1344 (O_1344,N_9963,N_9955);
or UO_1345 (O_1345,N_9979,N_9945);
and UO_1346 (O_1346,N_9964,N_9986);
nand UO_1347 (O_1347,N_9938,N_9927);
nor UO_1348 (O_1348,N_9952,N_9902);
xor UO_1349 (O_1349,N_9944,N_9972);
nor UO_1350 (O_1350,N_9951,N_9913);
and UO_1351 (O_1351,N_9947,N_9918);
and UO_1352 (O_1352,N_9991,N_9943);
or UO_1353 (O_1353,N_9940,N_9944);
nand UO_1354 (O_1354,N_9934,N_9935);
nor UO_1355 (O_1355,N_9908,N_9949);
or UO_1356 (O_1356,N_9948,N_9904);
nand UO_1357 (O_1357,N_9935,N_9918);
or UO_1358 (O_1358,N_9949,N_9961);
xnor UO_1359 (O_1359,N_9979,N_9925);
or UO_1360 (O_1360,N_9946,N_9900);
and UO_1361 (O_1361,N_9947,N_9979);
and UO_1362 (O_1362,N_9933,N_9979);
and UO_1363 (O_1363,N_9976,N_9994);
nand UO_1364 (O_1364,N_9946,N_9995);
and UO_1365 (O_1365,N_9973,N_9956);
and UO_1366 (O_1366,N_9992,N_9923);
or UO_1367 (O_1367,N_9920,N_9960);
xnor UO_1368 (O_1368,N_9941,N_9920);
or UO_1369 (O_1369,N_9960,N_9984);
and UO_1370 (O_1370,N_9948,N_9924);
and UO_1371 (O_1371,N_9937,N_9926);
nor UO_1372 (O_1372,N_9925,N_9950);
or UO_1373 (O_1373,N_9967,N_9979);
xnor UO_1374 (O_1374,N_9947,N_9988);
nand UO_1375 (O_1375,N_9952,N_9953);
and UO_1376 (O_1376,N_9924,N_9928);
and UO_1377 (O_1377,N_9904,N_9983);
nand UO_1378 (O_1378,N_9984,N_9993);
or UO_1379 (O_1379,N_9928,N_9995);
or UO_1380 (O_1380,N_9911,N_9962);
nor UO_1381 (O_1381,N_9928,N_9979);
nor UO_1382 (O_1382,N_9912,N_9994);
or UO_1383 (O_1383,N_9942,N_9929);
or UO_1384 (O_1384,N_9913,N_9926);
nor UO_1385 (O_1385,N_9950,N_9962);
or UO_1386 (O_1386,N_9916,N_9968);
or UO_1387 (O_1387,N_9974,N_9988);
nor UO_1388 (O_1388,N_9950,N_9913);
nor UO_1389 (O_1389,N_9932,N_9920);
xor UO_1390 (O_1390,N_9960,N_9985);
or UO_1391 (O_1391,N_9999,N_9994);
nand UO_1392 (O_1392,N_9953,N_9967);
and UO_1393 (O_1393,N_9957,N_9905);
and UO_1394 (O_1394,N_9926,N_9902);
or UO_1395 (O_1395,N_9922,N_9943);
or UO_1396 (O_1396,N_9996,N_9995);
nand UO_1397 (O_1397,N_9908,N_9900);
xor UO_1398 (O_1398,N_9932,N_9928);
nor UO_1399 (O_1399,N_9922,N_9933);
and UO_1400 (O_1400,N_9947,N_9963);
or UO_1401 (O_1401,N_9929,N_9932);
or UO_1402 (O_1402,N_9925,N_9922);
xor UO_1403 (O_1403,N_9925,N_9909);
nor UO_1404 (O_1404,N_9919,N_9995);
or UO_1405 (O_1405,N_9971,N_9942);
nor UO_1406 (O_1406,N_9911,N_9981);
xor UO_1407 (O_1407,N_9973,N_9931);
nand UO_1408 (O_1408,N_9997,N_9904);
nor UO_1409 (O_1409,N_9960,N_9966);
nand UO_1410 (O_1410,N_9911,N_9980);
nor UO_1411 (O_1411,N_9978,N_9989);
nand UO_1412 (O_1412,N_9922,N_9984);
xnor UO_1413 (O_1413,N_9907,N_9971);
xor UO_1414 (O_1414,N_9923,N_9911);
nor UO_1415 (O_1415,N_9954,N_9987);
and UO_1416 (O_1416,N_9987,N_9922);
nor UO_1417 (O_1417,N_9989,N_9947);
xnor UO_1418 (O_1418,N_9973,N_9915);
nand UO_1419 (O_1419,N_9900,N_9923);
and UO_1420 (O_1420,N_9989,N_9998);
nand UO_1421 (O_1421,N_9938,N_9975);
and UO_1422 (O_1422,N_9976,N_9947);
and UO_1423 (O_1423,N_9920,N_9989);
nor UO_1424 (O_1424,N_9900,N_9981);
or UO_1425 (O_1425,N_9962,N_9959);
xnor UO_1426 (O_1426,N_9977,N_9930);
nor UO_1427 (O_1427,N_9938,N_9943);
and UO_1428 (O_1428,N_9902,N_9983);
or UO_1429 (O_1429,N_9944,N_9909);
nand UO_1430 (O_1430,N_9949,N_9926);
nor UO_1431 (O_1431,N_9971,N_9918);
and UO_1432 (O_1432,N_9976,N_9967);
and UO_1433 (O_1433,N_9944,N_9916);
and UO_1434 (O_1434,N_9994,N_9929);
and UO_1435 (O_1435,N_9964,N_9926);
nor UO_1436 (O_1436,N_9930,N_9919);
or UO_1437 (O_1437,N_9965,N_9953);
nand UO_1438 (O_1438,N_9974,N_9922);
nor UO_1439 (O_1439,N_9976,N_9943);
nand UO_1440 (O_1440,N_9982,N_9934);
nand UO_1441 (O_1441,N_9935,N_9978);
nand UO_1442 (O_1442,N_9923,N_9922);
nand UO_1443 (O_1443,N_9974,N_9996);
nand UO_1444 (O_1444,N_9978,N_9957);
nor UO_1445 (O_1445,N_9962,N_9960);
or UO_1446 (O_1446,N_9968,N_9977);
nand UO_1447 (O_1447,N_9938,N_9982);
or UO_1448 (O_1448,N_9913,N_9963);
nor UO_1449 (O_1449,N_9941,N_9978);
and UO_1450 (O_1450,N_9981,N_9953);
and UO_1451 (O_1451,N_9998,N_9980);
and UO_1452 (O_1452,N_9949,N_9956);
and UO_1453 (O_1453,N_9948,N_9960);
nor UO_1454 (O_1454,N_9996,N_9972);
nand UO_1455 (O_1455,N_9990,N_9962);
or UO_1456 (O_1456,N_9966,N_9931);
and UO_1457 (O_1457,N_9940,N_9976);
or UO_1458 (O_1458,N_9980,N_9997);
or UO_1459 (O_1459,N_9905,N_9945);
and UO_1460 (O_1460,N_9957,N_9933);
or UO_1461 (O_1461,N_9905,N_9942);
and UO_1462 (O_1462,N_9989,N_9972);
xor UO_1463 (O_1463,N_9900,N_9909);
nand UO_1464 (O_1464,N_9986,N_9901);
xor UO_1465 (O_1465,N_9951,N_9950);
or UO_1466 (O_1466,N_9908,N_9918);
and UO_1467 (O_1467,N_9919,N_9917);
or UO_1468 (O_1468,N_9966,N_9980);
nand UO_1469 (O_1469,N_9975,N_9982);
nor UO_1470 (O_1470,N_9910,N_9909);
xor UO_1471 (O_1471,N_9990,N_9910);
xor UO_1472 (O_1472,N_9905,N_9994);
xor UO_1473 (O_1473,N_9921,N_9989);
and UO_1474 (O_1474,N_9995,N_9909);
or UO_1475 (O_1475,N_9956,N_9942);
nor UO_1476 (O_1476,N_9929,N_9940);
and UO_1477 (O_1477,N_9914,N_9966);
and UO_1478 (O_1478,N_9934,N_9919);
xor UO_1479 (O_1479,N_9962,N_9999);
nor UO_1480 (O_1480,N_9934,N_9904);
nor UO_1481 (O_1481,N_9927,N_9972);
and UO_1482 (O_1482,N_9936,N_9976);
xnor UO_1483 (O_1483,N_9964,N_9972);
or UO_1484 (O_1484,N_9998,N_9966);
or UO_1485 (O_1485,N_9929,N_9980);
xnor UO_1486 (O_1486,N_9972,N_9901);
xor UO_1487 (O_1487,N_9968,N_9912);
and UO_1488 (O_1488,N_9976,N_9986);
nand UO_1489 (O_1489,N_9917,N_9999);
or UO_1490 (O_1490,N_9907,N_9973);
nor UO_1491 (O_1491,N_9950,N_9908);
nor UO_1492 (O_1492,N_9979,N_9997);
nor UO_1493 (O_1493,N_9902,N_9907);
nor UO_1494 (O_1494,N_9915,N_9910);
nand UO_1495 (O_1495,N_9917,N_9942);
or UO_1496 (O_1496,N_9989,N_9937);
nand UO_1497 (O_1497,N_9979,N_9926);
or UO_1498 (O_1498,N_9925,N_9972);
or UO_1499 (O_1499,N_9933,N_9908);
endmodule