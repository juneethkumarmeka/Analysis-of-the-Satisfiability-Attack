module basic_500_3000_500_6_levels_5xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_431,In_97);
or U1 (N_1,In_166,In_290);
nand U2 (N_2,In_164,In_465);
nor U3 (N_3,In_47,In_128);
and U4 (N_4,In_466,In_67);
nor U5 (N_5,In_124,In_358);
or U6 (N_6,In_69,In_120);
or U7 (N_7,In_132,In_178);
nand U8 (N_8,In_84,In_262);
nor U9 (N_9,In_20,In_103);
nand U10 (N_10,In_375,In_188);
nand U11 (N_11,In_207,In_353);
nor U12 (N_12,In_180,In_0);
xor U13 (N_13,In_364,In_244);
or U14 (N_14,In_352,In_169);
nand U15 (N_15,In_165,In_469);
nor U16 (N_16,In_393,In_109);
nand U17 (N_17,In_298,In_36);
nor U18 (N_18,In_77,In_446);
nor U19 (N_19,In_57,In_331);
nor U20 (N_20,In_237,In_195);
or U21 (N_21,In_492,In_223);
and U22 (N_22,In_425,In_496);
and U23 (N_23,In_283,In_250);
and U24 (N_24,In_40,In_367);
and U25 (N_25,In_398,In_285);
nand U26 (N_26,In_216,In_155);
xnor U27 (N_27,In_487,In_481);
or U28 (N_28,In_76,In_72);
and U29 (N_29,In_86,In_498);
nand U30 (N_30,In_122,In_133);
or U31 (N_31,In_260,In_483);
xor U32 (N_32,In_211,In_127);
nor U33 (N_33,In_177,In_362);
nor U34 (N_34,In_63,In_130);
nand U35 (N_35,In_389,In_87);
nand U36 (N_36,In_28,In_117);
and U37 (N_37,In_332,In_248);
nand U38 (N_38,In_312,In_288);
xor U39 (N_39,In_82,In_279);
nand U40 (N_40,In_58,In_25);
or U41 (N_41,In_236,In_340);
or U42 (N_42,In_246,In_476);
nor U43 (N_43,In_255,In_175);
nand U44 (N_44,In_239,In_380);
nand U45 (N_45,In_454,In_105);
and U46 (N_46,In_320,In_489);
and U47 (N_47,In_327,In_281);
nand U48 (N_48,In_245,In_61);
or U49 (N_49,In_444,In_43);
nand U50 (N_50,In_346,In_2);
or U51 (N_51,In_123,In_74);
or U52 (N_52,In_297,In_261);
xor U53 (N_53,In_418,In_194);
and U54 (N_54,In_107,In_140);
xnor U55 (N_55,In_95,In_83);
nand U56 (N_56,In_277,In_486);
nor U57 (N_57,In_1,In_464);
nor U58 (N_58,In_394,In_263);
or U59 (N_59,In_354,In_210);
or U60 (N_60,In_447,In_435);
and U61 (N_61,In_342,In_171);
and U62 (N_62,In_403,In_462);
nand U63 (N_63,In_493,In_280);
nand U64 (N_64,In_173,In_313);
xor U65 (N_65,In_348,In_150);
nor U66 (N_66,In_247,In_70);
or U67 (N_67,In_160,In_268);
and U68 (N_68,In_186,In_409);
or U69 (N_69,In_34,In_92);
nand U70 (N_70,In_46,In_322);
xnor U71 (N_71,In_142,In_345);
nor U72 (N_72,In_491,In_391);
and U73 (N_73,In_151,In_271);
or U74 (N_74,In_60,In_439);
and U75 (N_75,In_51,In_220);
or U76 (N_76,In_448,In_114);
and U77 (N_77,In_264,In_181);
nand U78 (N_78,In_480,In_372);
xor U79 (N_79,In_126,In_197);
or U80 (N_80,In_33,In_406);
and U81 (N_81,In_416,In_470);
nor U82 (N_82,In_295,In_162);
nor U83 (N_83,In_8,In_225);
or U84 (N_84,In_484,In_282);
and U85 (N_85,In_401,In_4);
and U86 (N_86,In_26,In_89);
nor U87 (N_87,In_205,In_6);
or U88 (N_88,In_318,In_330);
nor U89 (N_89,In_427,In_347);
and U90 (N_90,In_185,In_52);
nor U91 (N_91,In_184,In_218);
nor U92 (N_92,In_350,In_110);
nor U93 (N_93,In_78,In_256);
or U94 (N_94,In_414,In_229);
or U95 (N_95,In_198,In_112);
or U96 (N_96,In_19,In_306);
or U97 (N_97,In_287,In_208);
nand U98 (N_98,In_485,In_232);
and U99 (N_99,In_10,In_324);
nor U100 (N_100,In_302,In_49);
and U101 (N_101,In_59,In_235);
or U102 (N_102,In_265,In_479);
nor U103 (N_103,In_121,In_168);
and U104 (N_104,In_240,In_407);
and U105 (N_105,In_118,In_81);
nand U106 (N_106,In_284,In_148);
nand U107 (N_107,In_432,In_7);
or U108 (N_108,In_16,In_317);
or U109 (N_109,In_228,In_495);
and U110 (N_110,In_349,In_385);
xnor U111 (N_111,In_199,In_286);
or U112 (N_112,In_471,In_278);
nor U113 (N_113,In_412,In_292);
or U114 (N_114,In_193,In_338);
and U115 (N_115,In_440,In_450);
and U116 (N_116,In_434,In_377);
or U117 (N_117,In_88,In_259);
nor U118 (N_118,In_215,In_68);
or U119 (N_119,In_80,In_91);
nand U120 (N_120,In_390,In_366);
nand U121 (N_121,In_399,In_191);
or U122 (N_122,In_341,In_326);
or U123 (N_123,In_23,In_293);
and U124 (N_124,In_299,In_159);
and U125 (N_125,In_337,In_189);
nand U126 (N_126,In_3,In_101);
or U127 (N_127,In_386,In_314);
nor U128 (N_128,In_417,In_316);
nand U129 (N_129,In_339,In_45);
or U130 (N_130,In_217,In_9);
or U131 (N_131,In_149,In_368);
and U132 (N_132,In_145,In_424);
xor U133 (N_133,In_397,In_272);
and U134 (N_134,In_359,In_41);
or U135 (N_135,In_116,In_29);
xor U136 (N_136,In_309,In_163);
nand U137 (N_137,In_307,In_463);
and U138 (N_138,In_176,In_275);
or U139 (N_139,In_413,In_323);
nor U140 (N_140,In_94,In_451);
or U141 (N_141,In_442,In_50);
nor U142 (N_142,In_54,In_460);
nand U143 (N_143,In_161,In_154);
and U144 (N_144,In_66,In_443);
xor U145 (N_145,In_104,In_141);
xor U146 (N_146,In_333,In_482);
nand U147 (N_147,In_294,In_325);
nor U148 (N_148,In_497,In_422);
nand U149 (N_149,In_289,In_137);
and U150 (N_150,In_300,In_405);
and U151 (N_151,In_230,In_429);
nor U152 (N_152,In_182,In_379);
nand U153 (N_153,In_301,In_304);
and U154 (N_154,In_35,In_310);
nand U155 (N_155,In_98,In_455);
or U156 (N_156,In_421,In_461);
nor U157 (N_157,In_321,In_231);
nand U158 (N_158,In_381,In_305);
nand U159 (N_159,In_363,In_212);
nor U160 (N_160,In_38,In_308);
xnor U161 (N_161,In_125,In_62);
xnor U162 (N_162,In_488,In_274);
or U163 (N_163,In_222,In_370);
or U164 (N_164,In_241,In_219);
or U165 (N_165,In_378,In_31);
and U166 (N_166,In_373,In_113);
xor U167 (N_167,In_419,In_5);
or U168 (N_168,In_64,In_190);
nand U169 (N_169,In_388,In_226);
nand U170 (N_170,In_200,In_172);
and U171 (N_171,In_315,In_430);
nand U172 (N_172,In_257,In_201);
or U173 (N_173,In_192,In_473);
or U174 (N_174,In_170,In_392);
and U175 (N_175,In_179,In_39);
or U176 (N_176,In_65,In_146);
and U177 (N_177,In_355,In_18);
and U178 (N_178,In_213,In_108);
or U179 (N_179,In_85,In_356);
or U180 (N_180,In_227,In_79);
and U181 (N_181,In_343,In_458);
nand U182 (N_182,In_144,In_404);
and U183 (N_183,In_267,In_73);
xor U184 (N_184,In_344,In_15);
nor U185 (N_185,In_396,In_291);
or U186 (N_186,In_402,In_11);
or U187 (N_187,In_100,In_93);
nor U188 (N_188,In_99,In_303);
nand U189 (N_189,In_209,In_328);
and U190 (N_190,In_369,In_472);
nor U191 (N_191,In_351,In_249);
xor U192 (N_192,In_428,In_90);
nor U193 (N_193,In_233,In_410);
or U194 (N_194,In_253,In_203);
or U195 (N_195,In_468,In_361);
xnor U196 (N_196,In_30,In_420);
xnor U197 (N_197,In_129,In_478);
nor U198 (N_198,In_258,In_311);
nor U199 (N_199,In_329,In_234);
or U200 (N_200,In_21,In_187);
and U201 (N_201,In_37,In_365);
and U202 (N_202,In_436,In_376);
nand U203 (N_203,In_445,In_13);
nand U204 (N_204,In_336,In_136);
or U205 (N_205,In_152,In_174);
nand U206 (N_206,In_96,In_252);
nand U207 (N_207,In_449,In_467);
nand U208 (N_208,In_499,In_243);
or U209 (N_209,In_17,In_131);
or U210 (N_210,In_56,In_474);
nand U211 (N_211,In_156,In_374);
or U212 (N_212,In_204,In_296);
and U213 (N_213,In_55,In_395);
nor U214 (N_214,In_106,In_433);
and U215 (N_215,In_102,In_242);
or U216 (N_216,In_360,In_251);
nor U217 (N_217,In_266,In_224);
nor U218 (N_218,In_270,In_371);
nor U219 (N_219,In_139,In_276);
or U220 (N_220,In_456,In_457);
and U221 (N_221,In_415,In_384);
or U222 (N_222,In_453,In_441);
and U223 (N_223,In_238,In_138);
or U224 (N_224,In_143,In_75);
nor U225 (N_225,In_158,In_452);
and U226 (N_226,In_147,In_71);
or U227 (N_227,In_115,In_153);
nor U228 (N_228,In_423,In_167);
or U229 (N_229,In_32,In_157);
nand U230 (N_230,In_44,In_494);
and U231 (N_231,In_382,In_438);
and U232 (N_232,In_42,In_22);
nand U233 (N_233,In_411,In_319);
nand U234 (N_234,In_214,In_119);
or U235 (N_235,In_134,In_357);
nand U236 (N_236,In_111,In_269);
or U237 (N_237,In_335,In_196);
nor U238 (N_238,In_408,In_53);
nand U239 (N_239,In_221,In_383);
nor U240 (N_240,In_426,In_48);
nor U241 (N_241,In_183,In_202);
nor U242 (N_242,In_334,In_387);
and U243 (N_243,In_437,In_206);
nor U244 (N_244,In_490,In_27);
xnor U245 (N_245,In_135,In_477);
nor U246 (N_246,In_273,In_24);
nor U247 (N_247,In_14,In_459);
nor U248 (N_248,In_475,In_400);
xnor U249 (N_249,In_12,In_254);
and U250 (N_250,In_212,In_95);
nor U251 (N_251,In_186,In_453);
nand U252 (N_252,In_404,In_65);
nand U253 (N_253,In_45,In_157);
and U254 (N_254,In_116,In_419);
or U255 (N_255,In_315,In_14);
nor U256 (N_256,In_390,In_320);
nand U257 (N_257,In_456,In_319);
or U258 (N_258,In_479,In_267);
nor U259 (N_259,In_149,In_137);
nand U260 (N_260,In_475,In_487);
nor U261 (N_261,In_389,In_304);
nor U262 (N_262,In_72,In_46);
nor U263 (N_263,In_302,In_427);
nand U264 (N_264,In_378,In_128);
nor U265 (N_265,In_60,In_201);
and U266 (N_266,In_97,In_452);
or U267 (N_267,In_410,In_205);
nor U268 (N_268,In_330,In_158);
or U269 (N_269,In_445,In_245);
or U270 (N_270,In_216,In_323);
and U271 (N_271,In_212,In_477);
or U272 (N_272,In_361,In_23);
nor U273 (N_273,In_145,In_189);
nand U274 (N_274,In_211,In_160);
and U275 (N_275,In_261,In_31);
and U276 (N_276,In_2,In_413);
and U277 (N_277,In_282,In_214);
nand U278 (N_278,In_444,In_343);
or U279 (N_279,In_411,In_290);
or U280 (N_280,In_472,In_197);
nand U281 (N_281,In_116,In_365);
nor U282 (N_282,In_161,In_31);
xor U283 (N_283,In_236,In_20);
or U284 (N_284,In_316,In_77);
or U285 (N_285,In_380,In_171);
and U286 (N_286,In_133,In_495);
nor U287 (N_287,In_243,In_35);
nand U288 (N_288,In_445,In_364);
or U289 (N_289,In_250,In_465);
or U290 (N_290,In_241,In_85);
nand U291 (N_291,In_74,In_356);
and U292 (N_292,In_276,In_409);
nor U293 (N_293,In_52,In_422);
xor U294 (N_294,In_4,In_112);
and U295 (N_295,In_313,In_477);
nor U296 (N_296,In_21,In_40);
nor U297 (N_297,In_339,In_104);
xnor U298 (N_298,In_83,In_284);
nand U299 (N_299,In_301,In_371);
nor U300 (N_300,In_126,In_57);
or U301 (N_301,In_290,In_450);
nor U302 (N_302,In_248,In_387);
or U303 (N_303,In_205,In_33);
nand U304 (N_304,In_398,In_392);
or U305 (N_305,In_192,In_370);
or U306 (N_306,In_188,In_12);
nor U307 (N_307,In_351,In_292);
nor U308 (N_308,In_352,In_197);
nor U309 (N_309,In_311,In_23);
or U310 (N_310,In_344,In_229);
and U311 (N_311,In_78,In_484);
and U312 (N_312,In_491,In_454);
xnor U313 (N_313,In_224,In_127);
and U314 (N_314,In_139,In_386);
or U315 (N_315,In_87,In_362);
xnor U316 (N_316,In_280,In_475);
nand U317 (N_317,In_37,In_143);
and U318 (N_318,In_136,In_372);
or U319 (N_319,In_438,In_461);
nor U320 (N_320,In_170,In_52);
and U321 (N_321,In_416,In_119);
nor U322 (N_322,In_335,In_237);
or U323 (N_323,In_409,In_166);
nand U324 (N_324,In_418,In_499);
xor U325 (N_325,In_360,In_113);
and U326 (N_326,In_456,In_68);
nor U327 (N_327,In_416,In_259);
or U328 (N_328,In_290,In_461);
nand U329 (N_329,In_393,In_118);
or U330 (N_330,In_272,In_485);
and U331 (N_331,In_332,In_101);
or U332 (N_332,In_480,In_255);
xor U333 (N_333,In_5,In_425);
xor U334 (N_334,In_226,In_349);
or U335 (N_335,In_411,In_185);
and U336 (N_336,In_83,In_295);
nand U337 (N_337,In_118,In_120);
or U338 (N_338,In_468,In_466);
or U339 (N_339,In_269,In_127);
and U340 (N_340,In_25,In_235);
nand U341 (N_341,In_461,In_392);
nor U342 (N_342,In_104,In_113);
nor U343 (N_343,In_147,In_98);
nor U344 (N_344,In_245,In_457);
and U345 (N_345,In_43,In_22);
nor U346 (N_346,In_347,In_121);
or U347 (N_347,In_435,In_55);
nand U348 (N_348,In_366,In_198);
and U349 (N_349,In_191,In_45);
nand U350 (N_350,In_295,In_186);
nor U351 (N_351,In_398,In_407);
nor U352 (N_352,In_288,In_404);
or U353 (N_353,In_255,In_257);
nand U354 (N_354,In_98,In_483);
nand U355 (N_355,In_96,In_291);
nor U356 (N_356,In_457,In_47);
and U357 (N_357,In_30,In_82);
nor U358 (N_358,In_371,In_433);
xnor U359 (N_359,In_311,In_457);
or U360 (N_360,In_180,In_477);
nand U361 (N_361,In_346,In_90);
nand U362 (N_362,In_394,In_358);
nor U363 (N_363,In_355,In_281);
nand U364 (N_364,In_280,In_269);
nand U365 (N_365,In_338,In_222);
xnor U366 (N_366,In_344,In_35);
and U367 (N_367,In_214,In_339);
nand U368 (N_368,In_175,In_189);
or U369 (N_369,In_450,In_421);
and U370 (N_370,In_313,In_262);
nor U371 (N_371,In_231,In_100);
or U372 (N_372,In_406,In_325);
nor U373 (N_373,In_159,In_258);
and U374 (N_374,In_59,In_206);
nor U375 (N_375,In_171,In_151);
nor U376 (N_376,In_167,In_190);
or U377 (N_377,In_421,In_280);
xor U378 (N_378,In_295,In_159);
xor U379 (N_379,In_395,In_339);
or U380 (N_380,In_229,In_325);
or U381 (N_381,In_347,In_384);
nand U382 (N_382,In_270,In_214);
and U383 (N_383,In_207,In_391);
nand U384 (N_384,In_131,In_247);
xor U385 (N_385,In_154,In_446);
nor U386 (N_386,In_484,In_185);
nor U387 (N_387,In_133,In_199);
xor U388 (N_388,In_316,In_94);
nor U389 (N_389,In_445,In_190);
or U390 (N_390,In_91,In_206);
or U391 (N_391,In_462,In_159);
nor U392 (N_392,In_291,In_334);
nand U393 (N_393,In_462,In_270);
or U394 (N_394,In_334,In_270);
nor U395 (N_395,In_238,In_79);
nor U396 (N_396,In_26,In_245);
nor U397 (N_397,In_177,In_449);
nor U398 (N_398,In_296,In_219);
nand U399 (N_399,In_405,In_162);
or U400 (N_400,In_455,In_82);
nand U401 (N_401,In_80,In_60);
and U402 (N_402,In_245,In_294);
or U403 (N_403,In_40,In_157);
nor U404 (N_404,In_100,In_65);
or U405 (N_405,In_54,In_440);
and U406 (N_406,In_63,In_482);
xnor U407 (N_407,In_21,In_134);
and U408 (N_408,In_217,In_359);
or U409 (N_409,In_316,In_442);
and U410 (N_410,In_20,In_26);
nor U411 (N_411,In_404,In_176);
nor U412 (N_412,In_241,In_305);
and U413 (N_413,In_156,In_346);
or U414 (N_414,In_321,In_412);
and U415 (N_415,In_225,In_66);
and U416 (N_416,In_148,In_406);
nand U417 (N_417,In_2,In_165);
and U418 (N_418,In_90,In_405);
nand U419 (N_419,In_288,In_260);
or U420 (N_420,In_398,In_433);
or U421 (N_421,In_176,In_108);
and U422 (N_422,In_484,In_358);
and U423 (N_423,In_472,In_331);
nand U424 (N_424,In_99,In_476);
nor U425 (N_425,In_464,In_357);
and U426 (N_426,In_305,In_124);
nor U427 (N_427,In_99,In_39);
or U428 (N_428,In_9,In_487);
or U429 (N_429,In_57,In_311);
or U430 (N_430,In_434,In_345);
and U431 (N_431,In_363,In_292);
or U432 (N_432,In_146,In_144);
or U433 (N_433,In_142,In_48);
nand U434 (N_434,In_186,In_259);
nand U435 (N_435,In_301,In_442);
and U436 (N_436,In_180,In_343);
or U437 (N_437,In_345,In_292);
nand U438 (N_438,In_52,In_6);
nor U439 (N_439,In_101,In_70);
and U440 (N_440,In_279,In_347);
nor U441 (N_441,In_140,In_214);
xor U442 (N_442,In_84,In_88);
xnor U443 (N_443,In_178,In_303);
nor U444 (N_444,In_228,In_323);
and U445 (N_445,In_332,In_410);
or U446 (N_446,In_121,In_332);
and U447 (N_447,In_407,In_474);
and U448 (N_448,In_268,In_312);
and U449 (N_449,In_209,In_287);
and U450 (N_450,In_388,In_444);
or U451 (N_451,In_146,In_5);
nor U452 (N_452,In_144,In_264);
nor U453 (N_453,In_330,In_371);
and U454 (N_454,In_69,In_396);
and U455 (N_455,In_58,In_94);
or U456 (N_456,In_48,In_94);
and U457 (N_457,In_464,In_137);
and U458 (N_458,In_406,In_27);
nor U459 (N_459,In_289,In_197);
or U460 (N_460,In_267,In_265);
nand U461 (N_461,In_333,In_248);
nor U462 (N_462,In_300,In_4);
or U463 (N_463,In_46,In_35);
nand U464 (N_464,In_101,In_476);
nor U465 (N_465,In_427,In_384);
nor U466 (N_466,In_345,In_155);
or U467 (N_467,In_491,In_98);
nor U468 (N_468,In_478,In_180);
nor U469 (N_469,In_457,In_277);
or U470 (N_470,In_328,In_310);
nor U471 (N_471,In_254,In_446);
or U472 (N_472,In_51,In_202);
xor U473 (N_473,In_228,In_462);
nor U474 (N_474,In_90,In_3);
or U475 (N_475,In_144,In_366);
xor U476 (N_476,In_141,In_174);
nand U477 (N_477,In_400,In_349);
and U478 (N_478,In_23,In_358);
nor U479 (N_479,In_73,In_227);
or U480 (N_480,In_1,In_94);
and U481 (N_481,In_185,In_424);
nand U482 (N_482,In_116,In_158);
nor U483 (N_483,In_485,In_391);
or U484 (N_484,In_311,In_485);
nand U485 (N_485,In_63,In_246);
nand U486 (N_486,In_347,In_263);
nor U487 (N_487,In_186,In_135);
nand U488 (N_488,In_354,In_496);
or U489 (N_489,In_142,In_356);
nand U490 (N_490,In_89,In_230);
nand U491 (N_491,In_326,In_15);
or U492 (N_492,In_359,In_368);
nor U493 (N_493,In_330,In_203);
nor U494 (N_494,In_263,In_248);
or U495 (N_495,In_190,In_309);
xnor U496 (N_496,In_448,In_290);
xnor U497 (N_497,In_454,In_385);
or U498 (N_498,In_264,In_236);
nor U499 (N_499,In_391,In_380);
xnor U500 (N_500,N_370,N_262);
and U501 (N_501,N_30,N_192);
and U502 (N_502,N_329,N_267);
nand U503 (N_503,N_495,N_249);
and U504 (N_504,N_282,N_280);
nor U505 (N_505,N_472,N_85);
and U506 (N_506,N_106,N_420);
or U507 (N_507,N_298,N_250);
nor U508 (N_508,N_166,N_448);
nor U509 (N_509,N_492,N_176);
or U510 (N_510,N_22,N_43);
nand U511 (N_511,N_428,N_94);
and U512 (N_512,N_376,N_345);
xnor U513 (N_513,N_175,N_456);
xor U514 (N_514,N_463,N_398);
nor U515 (N_515,N_159,N_139);
nor U516 (N_516,N_226,N_169);
nor U517 (N_517,N_443,N_1);
nand U518 (N_518,N_58,N_287);
nor U519 (N_519,N_78,N_349);
nor U520 (N_520,N_227,N_450);
nand U521 (N_521,N_427,N_328);
nand U522 (N_522,N_423,N_89);
xor U523 (N_523,N_95,N_231);
nor U524 (N_524,N_454,N_440);
or U525 (N_525,N_236,N_147);
nor U526 (N_526,N_90,N_86);
or U527 (N_527,N_323,N_102);
and U528 (N_528,N_105,N_103);
or U529 (N_529,N_441,N_21);
nand U530 (N_530,N_145,N_317);
xor U531 (N_531,N_120,N_331);
or U532 (N_532,N_339,N_109);
or U533 (N_533,N_395,N_392);
and U534 (N_534,N_372,N_322);
or U535 (N_535,N_452,N_144);
or U536 (N_536,N_464,N_410);
xor U537 (N_537,N_430,N_297);
or U538 (N_538,N_218,N_238);
and U539 (N_539,N_32,N_68);
or U540 (N_540,N_351,N_332);
or U541 (N_541,N_379,N_397);
and U542 (N_542,N_325,N_158);
nand U543 (N_543,N_67,N_88);
and U544 (N_544,N_467,N_63);
nor U545 (N_545,N_4,N_148);
and U546 (N_546,N_152,N_256);
or U547 (N_547,N_26,N_112);
nor U548 (N_548,N_37,N_98);
and U549 (N_549,N_125,N_275);
xor U550 (N_550,N_178,N_404);
and U551 (N_551,N_38,N_377);
nand U552 (N_552,N_140,N_12);
nand U553 (N_553,N_9,N_433);
and U554 (N_554,N_243,N_39);
and U555 (N_555,N_260,N_278);
nand U556 (N_556,N_354,N_342);
nand U557 (N_557,N_59,N_274);
nand U558 (N_558,N_299,N_465);
xor U559 (N_559,N_264,N_284);
and U560 (N_560,N_437,N_10);
nand U561 (N_561,N_183,N_493);
or U562 (N_562,N_419,N_19);
or U563 (N_563,N_358,N_453);
nor U564 (N_564,N_247,N_401);
xnor U565 (N_565,N_435,N_458);
and U566 (N_566,N_16,N_424);
or U567 (N_567,N_45,N_131);
nand U568 (N_568,N_115,N_242);
and U569 (N_569,N_205,N_479);
nand U570 (N_570,N_241,N_20);
or U571 (N_571,N_214,N_407);
and U572 (N_572,N_172,N_173);
nand U573 (N_573,N_52,N_422);
and U574 (N_574,N_389,N_484);
xnor U575 (N_575,N_28,N_330);
nand U576 (N_576,N_113,N_359);
and U577 (N_577,N_170,N_228);
and U578 (N_578,N_283,N_213);
or U579 (N_579,N_27,N_321);
nand U580 (N_580,N_151,N_117);
nand U581 (N_581,N_223,N_224);
and U582 (N_582,N_219,N_7);
xor U583 (N_583,N_327,N_72);
nand U584 (N_584,N_201,N_432);
or U585 (N_585,N_266,N_305);
nand U586 (N_586,N_107,N_303);
nor U587 (N_587,N_82,N_498);
or U588 (N_588,N_204,N_100);
nand U589 (N_589,N_348,N_200);
and U590 (N_590,N_391,N_385);
and U591 (N_591,N_439,N_455);
nor U592 (N_592,N_14,N_483);
and U593 (N_593,N_235,N_56);
and U594 (N_594,N_77,N_251);
nor U595 (N_595,N_333,N_253);
nor U596 (N_596,N_234,N_451);
nor U597 (N_597,N_476,N_80);
nor U598 (N_598,N_347,N_50);
xnor U599 (N_599,N_135,N_184);
or U600 (N_600,N_296,N_17);
and U601 (N_601,N_289,N_124);
and U602 (N_602,N_373,N_336);
or U603 (N_603,N_0,N_3);
or U604 (N_604,N_365,N_315);
nor U605 (N_605,N_108,N_460);
and U606 (N_606,N_360,N_216);
nor U607 (N_607,N_269,N_215);
nand U608 (N_608,N_44,N_486);
nand U609 (N_609,N_134,N_74);
or U610 (N_610,N_6,N_421);
xor U611 (N_611,N_302,N_362);
nand U612 (N_612,N_64,N_411);
nor U613 (N_613,N_132,N_314);
xnor U614 (N_614,N_62,N_301);
and U615 (N_615,N_5,N_119);
nor U616 (N_616,N_23,N_11);
and U617 (N_617,N_255,N_61);
or U618 (N_618,N_149,N_319);
or U619 (N_619,N_118,N_79);
or U620 (N_620,N_101,N_384);
and U621 (N_621,N_245,N_368);
xor U622 (N_622,N_473,N_71);
and U623 (N_623,N_248,N_313);
nor U624 (N_624,N_304,N_265);
and U625 (N_625,N_48,N_364);
or U626 (N_626,N_188,N_163);
and U627 (N_627,N_55,N_335);
or U628 (N_628,N_8,N_346);
and U629 (N_629,N_344,N_292);
or U630 (N_630,N_165,N_261);
nor U631 (N_631,N_499,N_168);
or U632 (N_632,N_185,N_426);
and U633 (N_633,N_459,N_308);
or U634 (N_634,N_312,N_133);
xor U635 (N_635,N_233,N_116);
and U636 (N_636,N_374,N_121);
nor U637 (N_637,N_340,N_246);
nand U638 (N_638,N_399,N_127);
and U639 (N_639,N_155,N_154);
xnor U640 (N_640,N_445,N_66);
and U641 (N_641,N_300,N_320);
or U642 (N_642,N_309,N_29);
xor U643 (N_643,N_488,N_18);
nor U644 (N_644,N_177,N_53);
nor U645 (N_645,N_180,N_99);
or U646 (N_646,N_198,N_271);
nand U647 (N_647,N_475,N_478);
and U648 (N_648,N_489,N_257);
or U649 (N_649,N_356,N_326);
and U650 (N_650,N_137,N_84);
nor U651 (N_651,N_123,N_191);
xnor U652 (N_652,N_156,N_202);
or U653 (N_653,N_457,N_306);
nand U654 (N_654,N_468,N_469);
and U655 (N_655,N_111,N_294);
and U656 (N_656,N_466,N_291);
nand U657 (N_657,N_381,N_217);
or U658 (N_658,N_485,N_161);
nand U659 (N_659,N_114,N_334);
xor U660 (N_660,N_491,N_254);
xor U661 (N_661,N_279,N_222);
or U662 (N_662,N_409,N_211);
nor U663 (N_663,N_481,N_136);
and U664 (N_664,N_371,N_295);
nand U665 (N_665,N_199,N_174);
and U666 (N_666,N_57,N_229);
or U667 (N_667,N_24,N_497);
nand U668 (N_668,N_193,N_225);
and U669 (N_669,N_438,N_157);
nand U670 (N_670,N_341,N_436);
nor U671 (N_671,N_138,N_15);
and U672 (N_672,N_153,N_142);
nor U673 (N_673,N_51,N_353);
nor U674 (N_674,N_337,N_104);
xnor U675 (N_675,N_390,N_13);
and U676 (N_676,N_276,N_418);
and U677 (N_677,N_442,N_128);
or U678 (N_678,N_244,N_25);
or U679 (N_679,N_146,N_355);
nor U680 (N_680,N_240,N_367);
nand U681 (N_681,N_190,N_496);
nand U682 (N_682,N_447,N_417);
and U683 (N_683,N_110,N_209);
or U684 (N_684,N_273,N_141);
nand U685 (N_685,N_167,N_393);
or U686 (N_686,N_474,N_75);
and U687 (N_687,N_210,N_87);
and U688 (N_688,N_277,N_350);
or U689 (N_689,N_316,N_46);
nand U690 (N_690,N_434,N_413);
nor U691 (N_691,N_307,N_416);
nand U692 (N_692,N_408,N_31);
and U693 (N_693,N_293,N_162);
xor U694 (N_694,N_93,N_187);
and U695 (N_695,N_318,N_487);
nand U696 (N_696,N_324,N_494);
and U697 (N_697,N_396,N_194);
nand U698 (N_698,N_286,N_268);
and U699 (N_699,N_285,N_164);
and U700 (N_700,N_406,N_160);
or U701 (N_701,N_73,N_252);
nor U702 (N_702,N_338,N_361);
or U703 (N_703,N_363,N_263);
or U704 (N_704,N_387,N_40);
nand U705 (N_705,N_383,N_207);
nor U706 (N_706,N_446,N_212);
and U707 (N_707,N_36,N_414);
or U708 (N_708,N_378,N_415);
xnor U709 (N_709,N_237,N_189);
nor U710 (N_710,N_34,N_83);
nand U711 (N_711,N_311,N_81);
and U712 (N_712,N_366,N_288);
or U713 (N_713,N_461,N_412);
nor U714 (N_714,N_179,N_259);
nor U715 (N_715,N_480,N_203);
nor U716 (N_716,N_65,N_91);
or U717 (N_717,N_54,N_402);
nand U718 (N_718,N_92,N_122);
nand U719 (N_719,N_290,N_208);
nor U720 (N_720,N_33,N_182);
nand U721 (N_721,N_310,N_272);
nand U722 (N_722,N_171,N_42);
nand U723 (N_723,N_126,N_76);
nor U724 (N_724,N_357,N_425);
and U725 (N_725,N_181,N_130);
or U726 (N_726,N_380,N_369);
or U727 (N_727,N_47,N_477);
or U728 (N_728,N_431,N_70);
xor U729 (N_729,N_206,N_232);
and U730 (N_730,N_69,N_186);
or U731 (N_731,N_462,N_490);
or U732 (N_732,N_375,N_429);
nor U733 (N_733,N_394,N_2);
or U734 (N_734,N_197,N_96);
xnor U735 (N_735,N_221,N_388);
and U736 (N_736,N_482,N_150);
and U737 (N_737,N_281,N_352);
or U738 (N_738,N_405,N_41);
xnor U739 (N_739,N_60,N_270);
nand U740 (N_740,N_195,N_343);
and U741 (N_741,N_49,N_444);
nand U742 (N_742,N_449,N_400);
or U743 (N_743,N_382,N_35);
nor U744 (N_744,N_97,N_471);
nand U745 (N_745,N_258,N_129);
nand U746 (N_746,N_470,N_386);
xnor U747 (N_747,N_403,N_196);
nor U748 (N_748,N_220,N_239);
or U749 (N_749,N_230,N_143);
and U750 (N_750,N_275,N_238);
or U751 (N_751,N_3,N_402);
or U752 (N_752,N_489,N_418);
nor U753 (N_753,N_219,N_330);
and U754 (N_754,N_40,N_48);
or U755 (N_755,N_79,N_219);
nand U756 (N_756,N_78,N_409);
and U757 (N_757,N_453,N_469);
xor U758 (N_758,N_22,N_454);
nand U759 (N_759,N_164,N_308);
nor U760 (N_760,N_257,N_462);
xor U761 (N_761,N_427,N_16);
nand U762 (N_762,N_423,N_90);
nand U763 (N_763,N_490,N_104);
or U764 (N_764,N_124,N_496);
or U765 (N_765,N_44,N_282);
and U766 (N_766,N_138,N_182);
or U767 (N_767,N_413,N_52);
nor U768 (N_768,N_498,N_246);
nor U769 (N_769,N_159,N_215);
and U770 (N_770,N_400,N_28);
and U771 (N_771,N_71,N_191);
xnor U772 (N_772,N_454,N_225);
nand U773 (N_773,N_311,N_12);
nor U774 (N_774,N_72,N_1);
nand U775 (N_775,N_182,N_143);
nor U776 (N_776,N_86,N_152);
nor U777 (N_777,N_57,N_148);
nor U778 (N_778,N_374,N_477);
nand U779 (N_779,N_429,N_171);
and U780 (N_780,N_347,N_334);
and U781 (N_781,N_240,N_56);
nor U782 (N_782,N_62,N_314);
nand U783 (N_783,N_95,N_227);
and U784 (N_784,N_467,N_290);
or U785 (N_785,N_389,N_279);
nor U786 (N_786,N_1,N_26);
nand U787 (N_787,N_470,N_170);
nor U788 (N_788,N_469,N_441);
nand U789 (N_789,N_232,N_407);
or U790 (N_790,N_77,N_440);
or U791 (N_791,N_326,N_245);
xor U792 (N_792,N_418,N_221);
nor U793 (N_793,N_1,N_319);
and U794 (N_794,N_434,N_334);
and U795 (N_795,N_272,N_369);
or U796 (N_796,N_27,N_8);
and U797 (N_797,N_91,N_154);
nand U798 (N_798,N_423,N_307);
nand U799 (N_799,N_69,N_230);
or U800 (N_800,N_240,N_434);
xor U801 (N_801,N_229,N_388);
nor U802 (N_802,N_251,N_70);
nor U803 (N_803,N_91,N_166);
nand U804 (N_804,N_309,N_479);
and U805 (N_805,N_64,N_306);
or U806 (N_806,N_358,N_499);
xnor U807 (N_807,N_441,N_340);
nor U808 (N_808,N_430,N_257);
or U809 (N_809,N_115,N_13);
and U810 (N_810,N_140,N_83);
nor U811 (N_811,N_78,N_306);
or U812 (N_812,N_60,N_315);
nor U813 (N_813,N_472,N_442);
nand U814 (N_814,N_495,N_496);
xor U815 (N_815,N_257,N_175);
or U816 (N_816,N_493,N_306);
nor U817 (N_817,N_382,N_29);
nand U818 (N_818,N_229,N_96);
or U819 (N_819,N_49,N_425);
nor U820 (N_820,N_97,N_61);
nand U821 (N_821,N_187,N_104);
nor U822 (N_822,N_403,N_356);
and U823 (N_823,N_141,N_96);
or U824 (N_824,N_346,N_304);
nand U825 (N_825,N_40,N_449);
or U826 (N_826,N_159,N_347);
nand U827 (N_827,N_286,N_79);
or U828 (N_828,N_21,N_471);
or U829 (N_829,N_167,N_293);
nor U830 (N_830,N_227,N_48);
nand U831 (N_831,N_48,N_403);
nand U832 (N_832,N_28,N_196);
nor U833 (N_833,N_140,N_132);
nor U834 (N_834,N_347,N_469);
nor U835 (N_835,N_282,N_128);
or U836 (N_836,N_446,N_43);
nand U837 (N_837,N_243,N_148);
or U838 (N_838,N_16,N_219);
and U839 (N_839,N_204,N_263);
or U840 (N_840,N_272,N_239);
or U841 (N_841,N_57,N_311);
nor U842 (N_842,N_454,N_91);
or U843 (N_843,N_447,N_67);
and U844 (N_844,N_437,N_88);
nor U845 (N_845,N_96,N_179);
or U846 (N_846,N_302,N_471);
or U847 (N_847,N_453,N_343);
or U848 (N_848,N_272,N_37);
nor U849 (N_849,N_457,N_255);
or U850 (N_850,N_73,N_30);
and U851 (N_851,N_84,N_214);
and U852 (N_852,N_498,N_14);
nor U853 (N_853,N_212,N_254);
nor U854 (N_854,N_416,N_140);
or U855 (N_855,N_236,N_275);
or U856 (N_856,N_375,N_27);
nor U857 (N_857,N_78,N_243);
or U858 (N_858,N_126,N_465);
nor U859 (N_859,N_12,N_209);
and U860 (N_860,N_470,N_419);
or U861 (N_861,N_84,N_408);
and U862 (N_862,N_435,N_489);
and U863 (N_863,N_300,N_185);
and U864 (N_864,N_433,N_133);
or U865 (N_865,N_283,N_316);
nand U866 (N_866,N_135,N_252);
or U867 (N_867,N_314,N_204);
and U868 (N_868,N_348,N_133);
and U869 (N_869,N_133,N_292);
or U870 (N_870,N_188,N_88);
nor U871 (N_871,N_327,N_102);
nor U872 (N_872,N_431,N_424);
or U873 (N_873,N_46,N_450);
nor U874 (N_874,N_384,N_376);
and U875 (N_875,N_278,N_267);
or U876 (N_876,N_339,N_81);
nor U877 (N_877,N_26,N_357);
and U878 (N_878,N_197,N_251);
nand U879 (N_879,N_283,N_358);
nand U880 (N_880,N_215,N_496);
nor U881 (N_881,N_299,N_477);
and U882 (N_882,N_16,N_81);
or U883 (N_883,N_222,N_186);
nor U884 (N_884,N_102,N_475);
or U885 (N_885,N_86,N_308);
nand U886 (N_886,N_285,N_10);
nor U887 (N_887,N_200,N_314);
xnor U888 (N_888,N_403,N_24);
nand U889 (N_889,N_59,N_138);
or U890 (N_890,N_138,N_349);
or U891 (N_891,N_313,N_295);
or U892 (N_892,N_397,N_125);
nor U893 (N_893,N_493,N_256);
xor U894 (N_894,N_208,N_411);
or U895 (N_895,N_92,N_88);
xnor U896 (N_896,N_113,N_340);
nand U897 (N_897,N_468,N_387);
or U898 (N_898,N_271,N_388);
xor U899 (N_899,N_271,N_371);
nor U900 (N_900,N_299,N_366);
nand U901 (N_901,N_223,N_295);
and U902 (N_902,N_416,N_306);
and U903 (N_903,N_315,N_163);
or U904 (N_904,N_228,N_87);
and U905 (N_905,N_344,N_305);
nor U906 (N_906,N_3,N_369);
and U907 (N_907,N_37,N_11);
or U908 (N_908,N_450,N_120);
or U909 (N_909,N_404,N_310);
xor U910 (N_910,N_178,N_450);
or U911 (N_911,N_401,N_117);
nor U912 (N_912,N_264,N_431);
nand U913 (N_913,N_428,N_183);
or U914 (N_914,N_312,N_39);
and U915 (N_915,N_417,N_441);
xor U916 (N_916,N_183,N_66);
and U917 (N_917,N_297,N_96);
or U918 (N_918,N_63,N_340);
or U919 (N_919,N_205,N_173);
nand U920 (N_920,N_329,N_459);
nand U921 (N_921,N_24,N_133);
nand U922 (N_922,N_275,N_112);
xor U923 (N_923,N_255,N_397);
and U924 (N_924,N_270,N_59);
nor U925 (N_925,N_142,N_418);
and U926 (N_926,N_280,N_486);
and U927 (N_927,N_480,N_345);
nand U928 (N_928,N_85,N_357);
or U929 (N_929,N_245,N_361);
nand U930 (N_930,N_348,N_244);
or U931 (N_931,N_418,N_487);
nand U932 (N_932,N_142,N_319);
and U933 (N_933,N_206,N_133);
or U934 (N_934,N_108,N_271);
xor U935 (N_935,N_427,N_391);
nand U936 (N_936,N_85,N_311);
and U937 (N_937,N_156,N_29);
nor U938 (N_938,N_469,N_210);
nor U939 (N_939,N_480,N_416);
nor U940 (N_940,N_371,N_290);
nor U941 (N_941,N_394,N_320);
nor U942 (N_942,N_373,N_293);
nor U943 (N_943,N_1,N_96);
or U944 (N_944,N_165,N_461);
nor U945 (N_945,N_157,N_495);
nor U946 (N_946,N_279,N_408);
and U947 (N_947,N_327,N_461);
or U948 (N_948,N_225,N_449);
and U949 (N_949,N_421,N_292);
or U950 (N_950,N_427,N_207);
nor U951 (N_951,N_201,N_204);
nor U952 (N_952,N_404,N_41);
and U953 (N_953,N_60,N_494);
and U954 (N_954,N_159,N_298);
nand U955 (N_955,N_266,N_242);
nor U956 (N_956,N_114,N_361);
nor U957 (N_957,N_319,N_304);
nor U958 (N_958,N_84,N_380);
or U959 (N_959,N_457,N_11);
and U960 (N_960,N_339,N_17);
xor U961 (N_961,N_254,N_140);
nand U962 (N_962,N_10,N_414);
or U963 (N_963,N_435,N_44);
nand U964 (N_964,N_483,N_170);
or U965 (N_965,N_127,N_294);
nor U966 (N_966,N_21,N_224);
nand U967 (N_967,N_385,N_486);
or U968 (N_968,N_307,N_467);
xor U969 (N_969,N_384,N_11);
and U970 (N_970,N_168,N_160);
or U971 (N_971,N_263,N_118);
or U972 (N_972,N_248,N_309);
xnor U973 (N_973,N_217,N_45);
or U974 (N_974,N_445,N_368);
or U975 (N_975,N_74,N_21);
and U976 (N_976,N_411,N_42);
or U977 (N_977,N_308,N_44);
xor U978 (N_978,N_223,N_154);
or U979 (N_979,N_296,N_459);
or U980 (N_980,N_483,N_464);
and U981 (N_981,N_262,N_215);
nand U982 (N_982,N_407,N_81);
nor U983 (N_983,N_422,N_291);
xor U984 (N_984,N_110,N_291);
xnor U985 (N_985,N_169,N_419);
xor U986 (N_986,N_491,N_86);
xor U987 (N_987,N_214,N_158);
nor U988 (N_988,N_491,N_147);
xor U989 (N_989,N_92,N_175);
or U990 (N_990,N_365,N_200);
nor U991 (N_991,N_463,N_155);
or U992 (N_992,N_53,N_65);
nand U993 (N_993,N_93,N_225);
nand U994 (N_994,N_105,N_292);
nand U995 (N_995,N_179,N_171);
and U996 (N_996,N_79,N_437);
or U997 (N_997,N_354,N_492);
or U998 (N_998,N_20,N_259);
or U999 (N_999,N_30,N_14);
nand U1000 (N_1000,N_778,N_957);
or U1001 (N_1001,N_539,N_536);
and U1002 (N_1002,N_954,N_515);
and U1003 (N_1003,N_906,N_933);
and U1004 (N_1004,N_971,N_698);
and U1005 (N_1005,N_689,N_828);
nand U1006 (N_1006,N_719,N_656);
or U1007 (N_1007,N_584,N_932);
or U1008 (N_1008,N_592,N_648);
or U1009 (N_1009,N_973,N_585);
nand U1010 (N_1010,N_830,N_702);
and U1011 (N_1011,N_647,N_559);
or U1012 (N_1012,N_683,N_696);
nand U1013 (N_1013,N_996,N_629);
nor U1014 (N_1014,N_734,N_995);
and U1015 (N_1015,N_975,N_739);
and U1016 (N_1016,N_746,N_628);
and U1017 (N_1017,N_606,N_994);
and U1018 (N_1018,N_791,N_888);
nor U1019 (N_1019,N_573,N_985);
and U1020 (N_1020,N_969,N_833);
or U1021 (N_1021,N_652,N_547);
or U1022 (N_1022,N_821,N_999);
or U1023 (N_1023,N_605,N_674);
or U1024 (N_1024,N_760,N_820);
and U1025 (N_1025,N_521,N_890);
or U1026 (N_1026,N_646,N_838);
nor U1027 (N_1027,N_776,N_849);
or U1028 (N_1028,N_787,N_618);
nand U1029 (N_1029,N_621,N_765);
nand U1030 (N_1030,N_854,N_958);
nand U1031 (N_1031,N_750,N_844);
and U1032 (N_1032,N_793,N_917);
nor U1033 (N_1033,N_856,N_633);
nand U1034 (N_1034,N_612,N_721);
nand U1035 (N_1035,N_553,N_679);
nand U1036 (N_1036,N_916,N_617);
nor U1037 (N_1037,N_927,N_964);
nand U1038 (N_1038,N_540,N_896);
and U1039 (N_1039,N_625,N_865);
nand U1040 (N_1040,N_915,N_759);
or U1041 (N_1041,N_563,N_730);
and U1042 (N_1042,N_587,N_538);
or U1043 (N_1043,N_703,N_792);
or U1044 (N_1044,N_593,N_567);
nand U1045 (N_1045,N_959,N_818);
nor U1046 (N_1046,N_529,N_526);
nand U1047 (N_1047,N_517,N_744);
nor U1048 (N_1048,N_962,N_518);
nand U1049 (N_1049,N_986,N_914);
and U1050 (N_1050,N_913,N_904);
nor U1051 (N_1051,N_556,N_837);
or U1052 (N_1052,N_983,N_903);
nor U1053 (N_1053,N_641,N_666);
nor U1054 (N_1054,N_723,N_998);
nor U1055 (N_1055,N_832,N_626);
and U1056 (N_1056,N_525,N_823);
xor U1057 (N_1057,N_619,N_937);
and U1058 (N_1058,N_875,N_551);
or U1059 (N_1059,N_852,N_535);
nor U1060 (N_1060,N_966,N_813);
nand U1061 (N_1061,N_943,N_910);
or U1062 (N_1062,N_727,N_543);
nand U1063 (N_1063,N_976,N_511);
and U1064 (N_1064,N_694,N_700);
nand U1065 (N_1065,N_705,N_710);
and U1066 (N_1066,N_632,N_790);
or U1067 (N_1067,N_729,N_816);
and U1068 (N_1068,N_970,N_968);
nor U1069 (N_1069,N_627,N_835);
or U1070 (N_1070,N_767,N_575);
nor U1071 (N_1071,N_921,N_939);
nand U1072 (N_1072,N_747,N_523);
and U1073 (N_1073,N_610,N_850);
or U1074 (N_1074,N_794,N_686);
or U1075 (N_1075,N_918,N_659);
nand U1076 (N_1076,N_631,N_501);
or U1077 (N_1077,N_929,N_909);
nor U1078 (N_1078,N_931,N_675);
nor U1079 (N_1079,N_984,N_819);
nor U1080 (N_1080,N_634,N_616);
or U1081 (N_1081,N_578,N_831);
nor U1082 (N_1082,N_953,N_722);
and U1083 (N_1083,N_800,N_944);
nand U1084 (N_1084,N_745,N_712);
nor U1085 (N_1085,N_718,N_545);
or U1086 (N_1086,N_691,N_684);
or U1087 (N_1087,N_766,N_615);
xor U1088 (N_1088,N_881,N_528);
and U1089 (N_1089,N_770,N_560);
and U1090 (N_1090,N_795,N_542);
nor U1091 (N_1091,N_952,N_704);
nor U1092 (N_1092,N_609,N_841);
nor U1093 (N_1093,N_640,N_847);
and U1094 (N_1094,N_965,N_869);
nor U1095 (N_1095,N_548,N_506);
nand U1096 (N_1096,N_512,N_514);
nor U1097 (N_1097,N_822,N_855);
nor U1098 (N_1098,N_980,N_599);
or U1099 (N_1099,N_639,N_733);
xnor U1100 (N_1100,N_873,N_576);
or U1101 (N_1101,N_902,N_851);
xnor U1102 (N_1102,N_789,N_907);
nand U1103 (N_1103,N_591,N_503);
nor U1104 (N_1104,N_509,N_596);
nand U1105 (N_1105,N_643,N_868);
nand U1106 (N_1106,N_737,N_784);
xor U1107 (N_1107,N_665,N_711);
nand U1108 (N_1108,N_565,N_883);
and U1109 (N_1109,N_668,N_751);
nor U1110 (N_1110,N_663,N_961);
or U1111 (N_1111,N_658,N_842);
nand U1112 (N_1112,N_775,N_810);
nor U1113 (N_1113,N_546,N_798);
and U1114 (N_1114,N_895,N_552);
and U1115 (N_1115,N_699,N_589);
nand U1116 (N_1116,N_924,N_945);
or U1117 (N_1117,N_877,N_992);
or U1118 (N_1118,N_814,N_566);
and U1119 (N_1119,N_504,N_845);
or U1120 (N_1120,N_912,N_779);
xor U1121 (N_1121,N_678,N_987);
xor U1122 (N_1122,N_951,N_701);
and U1123 (N_1123,N_595,N_935);
xnor U1124 (N_1124,N_754,N_941);
nand U1125 (N_1125,N_908,N_872);
and U1126 (N_1126,N_717,N_843);
nor U1127 (N_1127,N_581,N_669);
and U1128 (N_1128,N_682,N_500);
and U1129 (N_1129,N_502,N_714);
and U1130 (N_1130,N_786,N_748);
nand U1131 (N_1131,N_812,N_728);
nor U1132 (N_1132,N_863,N_649);
nand U1133 (N_1133,N_796,N_861);
nand U1134 (N_1134,N_622,N_756);
and U1135 (N_1135,N_771,N_857);
and U1136 (N_1136,N_724,N_860);
or U1137 (N_1137,N_706,N_799);
nand U1138 (N_1138,N_879,N_803);
or U1139 (N_1139,N_804,N_802);
nand U1140 (N_1140,N_695,N_527);
or U1141 (N_1141,N_541,N_967);
and U1142 (N_1142,N_726,N_707);
nand U1143 (N_1143,N_732,N_809);
nor U1144 (N_1144,N_664,N_922);
xor U1145 (N_1145,N_555,N_769);
nor U1146 (N_1146,N_533,N_570);
xnor U1147 (N_1147,N_989,N_824);
nor U1148 (N_1148,N_571,N_955);
nor U1149 (N_1149,N_624,N_940);
xnor U1150 (N_1150,N_513,N_781);
xnor U1151 (N_1151,N_900,N_887);
or U1152 (N_1152,N_607,N_763);
and U1153 (N_1153,N_884,N_600);
xor U1154 (N_1154,N_716,N_697);
or U1155 (N_1155,N_797,N_720);
xnor U1156 (N_1156,N_758,N_742);
nand U1157 (N_1157,N_774,N_738);
nor U1158 (N_1158,N_508,N_956);
xnor U1159 (N_1159,N_550,N_885);
nand U1160 (N_1160,N_840,N_544);
and U1161 (N_1161,N_685,N_898);
nand U1162 (N_1162,N_590,N_979);
nand U1163 (N_1163,N_761,N_806);
and U1164 (N_1164,N_532,N_637);
or U1165 (N_1165,N_653,N_926);
xor U1166 (N_1166,N_558,N_715);
nand U1167 (N_1167,N_782,N_892);
and U1168 (N_1168,N_897,N_755);
or U1169 (N_1169,N_708,N_925);
nand U1170 (N_1170,N_725,N_709);
and U1171 (N_1171,N_601,N_692);
nor U1172 (N_1172,N_825,N_598);
or U1173 (N_1173,N_524,N_537);
nand U1174 (N_1174,N_583,N_805);
or U1175 (N_1175,N_645,N_894);
nand U1176 (N_1176,N_911,N_671);
nand U1177 (N_1177,N_650,N_562);
nor U1178 (N_1178,N_839,N_569);
nor U1179 (N_1179,N_807,N_834);
or U1180 (N_1180,N_977,N_549);
nand U1181 (N_1181,N_743,N_949);
nor U1182 (N_1182,N_923,N_990);
nor U1183 (N_1183,N_870,N_773);
nand U1184 (N_1184,N_928,N_871);
or U1185 (N_1185,N_602,N_811);
xor U1186 (N_1186,N_777,N_862);
and U1187 (N_1187,N_530,N_950);
or U1188 (N_1188,N_880,N_801);
or U1189 (N_1189,N_772,N_946);
xor U1190 (N_1190,N_846,N_505);
nor U1191 (N_1191,N_693,N_853);
and U1192 (N_1192,N_905,N_597);
and U1193 (N_1193,N_938,N_919);
or U1194 (N_1194,N_808,N_687);
nand U1195 (N_1195,N_981,N_673);
xor U1196 (N_1196,N_901,N_564);
or U1197 (N_1197,N_878,N_613);
nand U1198 (N_1198,N_608,N_690);
nor U1199 (N_1199,N_997,N_749);
nand U1200 (N_1200,N_866,N_623);
nor U1201 (N_1201,N_603,N_561);
or U1202 (N_1202,N_815,N_635);
and U1203 (N_1203,N_594,N_736);
or U1204 (N_1204,N_672,N_768);
or U1205 (N_1205,N_620,N_757);
and U1206 (N_1206,N_630,N_788);
nand U1207 (N_1207,N_582,N_507);
and U1208 (N_1208,N_522,N_660);
or U1209 (N_1209,N_762,N_670);
and U1210 (N_1210,N_579,N_920);
or U1211 (N_1211,N_572,N_882);
or U1212 (N_1212,N_604,N_519);
xnor U1213 (N_1213,N_817,N_848);
or U1214 (N_1214,N_642,N_886);
or U1215 (N_1215,N_586,N_826);
or U1216 (N_1216,N_752,N_942);
and U1217 (N_1217,N_991,N_574);
nor U1218 (N_1218,N_948,N_753);
nand U1219 (N_1219,N_899,N_876);
and U1220 (N_1220,N_614,N_936);
nor U1221 (N_1221,N_829,N_534);
nor U1222 (N_1222,N_974,N_988);
and U1223 (N_1223,N_993,N_520);
nor U1224 (N_1224,N_662,N_972);
xnor U1225 (N_1225,N_651,N_735);
or U1226 (N_1226,N_681,N_531);
nor U1227 (N_1227,N_731,N_982);
nor U1228 (N_1228,N_516,N_661);
and U1229 (N_1229,N_891,N_780);
nor U1230 (N_1230,N_588,N_611);
or U1231 (N_1231,N_568,N_654);
nand U1232 (N_1232,N_836,N_783);
and U1233 (N_1233,N_688,N_580);
nor U1234 (N_1234,N_554,N_859);
nand U1235 (N_1235,N_963,N_644);
xnor U1236 (N_1236,N_867,N_930);
and U1237 (N_1237,N_858,N_785);
and U1238 (N_1238,N_657,N_636);
and U1239 (N_1239,N_889,N_960);
nor U1240 (N_1240,N_655,N_557);
or U1241 (N_1241,N_740,N_676);
nand U1242 (N_1242,N_947,N_978);
or U1243 (N_1243,N_741,N_827);
and U1244 (N_1244,N_893,N_680);
nand U1245 (N_1245,N_764,N_874);
nand U1246 (N_1246,N_667,N_677);
nand U1247 (N_1247,N_510,N_638);
nor U1248 (N_1248,N_864,N_713);
nand U1249 (N_1249,N_577,N_934);
nand U1250 (N_1250,N_666,N_606);
or U1251 (N_1251,N_531,N_860);
nand U1252 (N_1252,N_968,N_602);
nor U1253 (N_1253,N_519,N_830);
and U1254 (N_1254,N_865,N_964);
nor U1255 (N_1255,N_783,N_883);
and U1256 (N_1256,N_925,N_585);
xor U1257 (N_1257,N_530,N_534);
nor U1258 (N_1258,N_721,N_869);
and U1259 (N_1259,N_911,N_702);
xnor U1260 (N_1260,N_946,N_794);
nor U1261 (N_1261,N_870,N_724);
nand U1262 (N_1262,N_862,N_744);
or U1263 (N_1263,N_930,N_773);
and U1264 (N_1264,N_627,N_883);
nand U1265 (N_1265,N_565,N_561);
and U1266 (N_1266,N_609,N_566);
and U1267 (N_1267,N_880,N_883);
nand U1268 (N_1268,N_556,N_955);
nand U1269 (N_1269,N_568,N_687);
and U1270 (N_1270,N_538,N_660);
nor U1271 (N_1271,N_737,N_730);
nand U1272 (N_1272,N_737,N_752);
xor U1273 (N_1273,N_567,N_902);
and U1274 (N_1274,N_511,N_711);
nor U1275 (N_1275,N_681,N_931);
nand U1276 (N_1276,N_787,N_659);
nor U1277 (N_1277,N_908,N_835);
and U1278 (N_1278,N_930,N_863);
and U1279 (N_1279,N_585,N_629);
xnor U1280 (N_1280,N_531,N_932);
xor U1281 (N_1281,N_737,N_528);
nor U1282 (N_1282,N_580,N_563);
and U1283 (N_1283,N_923,N_905);
and U1284 (N_1284,N_811,N_899);
nor U1285 (N_1285,N_784,N_616);
or U1286 (N_1286,N_790,N_967);
nand U1287 (N_1287,N_627,N_766);
and U1288 (N_1288,N_803,N_936);
nor U1289 (N_1289,N_723,N_700);
nor U1290 (N_1290,N_619,N_584);
and U1291 (N_1291,N_625,N_964);
nand U1292 (N_1292,N_675,N_636);
xor U1293 (N_1293,N_617,N_823);
or U1294 (N_1294,N_824,N_914);
and U1295 (N_1295,N_649,N_620);
nand U1296 (N_1296,N_640,N_645);
nand U1297 (N_1297,N_839,N_998);
nand U1298 (N_1298,N_667,N_596);
nor U1299 (N_1299,N_524,N_841);
nor U1300 (N_1300,N_804,N_526);
and U1301 (N_1301,N_707,N_513);
nand U1302 (N_1302,N_724,N_884);
nand U1303 (N_1303,N_950,N_932);
and U1304 (N_1304,N_820,N_620);
xnor U1305 (N_1305,N_520,N_565);
nor U1306 (N_1306,N_881,N_642);
and U1307 (N_1307,N_502,N_654);
nand U1308 (N_1308,N_714,N_882);
nand U1309 (N_1309,N_939,N_603);
xnor U1310 (N_1310,N_527,N_614);
or U1311 (N_1311,N_525,N_575);
and U1312 (N_1312,N_992,N_934);
and U1313 (N_1313,N_896,N_998);
nor U1314 (N_1314,N_959,N_995);
nor U1315 (N_1315,N_961,N_918);
and U1316 (N_1316,N_544,N_805);
and U1317 (N_1317,N_506,N_848);
nor U1318 (N_1318,N_769,N_785);
nand U1319 (N_1319,N_811,N_506);
and U1320 (N_1320,N_998,N_784);
and U1321 (N_1321,N_881,N_856);
nand U1322 (N_1322,N_954,N_585);
or U1323 (N_1323,N_850,N_915);
nand U1324 (N_1324,N_813,N_972);
xnor U1325 (N_1325,N_709,N_620);
and U1326 (N_1326,N_721,N_784);
nor U1327 (N_1327,N_855,N_788);
nand U1328 (N_1328,N_823,N_652);
and U1329 (N_1329,N_513,N_833);
or U1330 (N_1330,N_836,N_802);
or U1331 (N_1331,N_829,N_650);
xnor U1332 (N_1332,N_881,N_781);
nor U1333 (N_1333,N_663,N_633);
or U1334 (N_1334,N_889,N_618);
nor U1335 (N_1335,N_728,N_718);
xnor U1336 (N_1336,N_797,N_601);
nor U1337 (N_1337,N_555,N_882);
and U1338 (N_1338,N_903,N_558);
or U1339 (N_1339,N_822,N_760);
xor U1340 (N_1340,N_727,N_705);
or U1341 (N_1341,N_995,N_540);
nand U1342 (N_1342,N_897,N_823);
nor U1343 (N_1343,N_950,N_851);
and U1344 (N_1344,N_529,N_648);
xnor U1345 (N_1345,N_934,N_675);
nand U1346 (N_1346,N_530,N_539);
and U1347 (N_1347,N_787,N_670);
nor U1348 (N_1348,N_673,N_537);
xor U1349 (N_1349,N_662,N_526);
or U1350 (N_1350,N_915,N_920);
xnor U1351 (N_1351,N_958,N_960);
nand U1352 (N_1352,N_905,N_688);
and U1353 (N_1353,N_512,N_566);
and U1354 (N_1354,N_728,N_813);
nand U1355 (N_1355,N_884,N_898);
or U1356 (N_1356,N_681,N_508);
nand U1357 (N_1357,N_983,N_751);
nor U1358 (N_1358,N_671,N_615);
or U1359 (N_1359,N_700,N_982);
xor U1360 (N_1360,N_742,N_831);
and U1361 (N_1361,N_725,N_754);
and U1362 (N_1362,N_787,N_509);
or U1363 (N_1363,N_594,N_767);
or U1364 (N_1364,N_611,N_599);
or U1365 (N_1365,N_631,N_948);
nand U1366 (N_1366,N_708,N_897);
nor U1367 (N_1367,N_866,N_535);
or U1368 (N_1368,N_753,N_623);
nand U1369 (N_1369,N_566,N_922);
or U1370 (N_1370,N_831,N_878);
or U1371 (N_1371,N_672,N_800);
nand U1372 (N_1372,N_539,N_931);
nor U1373 (N_1373,N_589,N_760);
and U1374 (N_1374,N_927,N_692);
xor U1375 (N_1375,N_652,N_609);
or U1376 (N_1376,N_591,N_860);
nand U1377 (N_1377,N_758,N_964);
or U1378 (N_1378,N_521,N_769);
and U1379 (N_1379,N_892,N_737);
or U1380 (N_1380,N_905,N_574);
nand U1381 (N_1381,N_868,N_536);
nand U1382 (N_1382,N_647,N_540);
or U1383 (N_1383,N_981,N_789);
and U1384 (N_1384,N_879,N_817);
nor U1385 (N_1385,N_753,N_761);
or U1386 (N_1386,N_978,N_990);
or U1387 (N_1387,N_609,N_688);
or U1388 (N_1388,N_839,N_647);
and U1389 (N_1389,N_824,N_822);
or U1390 (N_1390,N_535,N_631);
nand U1391 (N_1391,N_647,N_552);
nand U1392 (N_1392,N_558,N_634);
and U1393 (N_1393,N_623,N_908);
nor U1394 (N_1394,N_784,N_913);
xor U1395 (N_1395,N_528,N_754);
nand U1396 (N_1396,N_813,N_603);
nand U1397 (N_1397,N_753,N_594);
nor U1398 (N_1398,N_588,N_790);
nand U1399 (N_1399,N_930,N_685);
nand U1400 (N_1400,N_736,N_660);
nand U1401 (N_1401,N_993,N_839);
nand U1402 (N_1402,N_784,N_752);
and U1403 (N_1403,N_803,N_640);
xor U1404 (N_1404,N_882,N_540);
and U1405 (N_1405,N_709,N_795);
nand U1406 (N_1406,N_871,N_952);
nor U1407 (N_1407,N_893,N_974);
nor U1408 (N_1408,N_661,N_619);
or U1409 (N_1409,N_731,N_898);
nor U1410 (N_1410,N_509,N_965);
nor U1411 (N_1411,N_643,N_636);
nand U1412 (N_1412,N_570,N_526);
or U1413 (N_1413,N_565,N_998);
xnor U1414 (N_1414,N_777,N_583);
nor U1415 (N_1415,N_778,N_898);
and U1416 (N_1416,N_937,N_692);
or U1417 (N_1417,N_923,N_881);
nand U1418 (N_1418,N_591,N_529);
nor U1419 (N_1419,N_812,N_971);
or U1420 (N_1420,N_931,N_829);
or U1421 (N_1421,N_658,N_970);
nand U1422 (N_1422,N_704,N_567);
and U1423 (N_1423,N_837,N_573);
nand U1424 (N_1424,N_532,N_547);
nor U1425 (N_1425,N_650,N_550);
or U1426 (N_1426,N_729,N_904);
nand U1427 (N_1427,N_716,N_740);
and U1428 (N_1428,N_823,N_925);
nand U1429 (N_1429,N_823,N_779);
nand U1430 (N_1430,N_639,N_833);
nor U1431 (N_1431,N_698,N_513);
or U1432 (N_1432,N_632,N_651);
nor U1433 (N_1433,N_948,N_975);
nor U1434 (N_1434,N_930,N_660);
or U1435 (N_1435,N_817,N_703);
nand U1436 (N_1436,N_649,N_693);
nor U1437 (N_1437,N_995,N_547);
xnor U1438 (N_1438,N_984,N_930);
and U1439 (N_1439,N_755,N_678);
nand U1440 (N_1440,N_896,N_723);
or U1441 (N_1441,N_532,N_628);
and U1442 (N_1442,N_532,N_905);
and U1443 (N_1443,N_722,N_741);
nor U1444 (N_1444,N_781,N_784);
xnor U1445 (N_1445,N_781,N_643);
nand U1446 (N_1446,N_857,N_518);
and U1447 (N_1447,N_750,N_885);
and U1448 (N_1448,N_811,N_532);
nor U1449 (N_1449,N_871,N_809);
and U1450 (N_1450,N_555,N_919);
nor U1451 (N_1451,N_663,N_722);
xnor U1452 (N_1452,N_701,N_914);
and U1453 (N_1453,N_843,N_840);
and U1454 (N_1454,N_968,N_788);
and U1455 (N_1455,N_898,N_604);
nor U1456 (N_1456,N_641,N_774);
nand U1457 (N_1457,N_587,N_950);
or U1458 (N_1458,N_966,N_848);
nor U1459 (N_1459,N_897,N_693);
and U1460 (N_1460,N_911,N_592);
or U1461 (N_1461,N_894,N_581);
nand U1462 (N_1462,N_593,N_912);
nor U1463 (N_1463,N_887,N_631);
or U1464 (N_1464,N_709,N_819);
nand U1465 (N_1465,N_654,N_624);
xnor U1466 (N_1466,N_651,N_664);
and U1467 (N_1467,N_764,N_880);
nor U1468 (N_1468,N_594,N_835);
and U1469 (N_1469,N_810,N_740);
nor U1470 (N_1470,N_752,N_890);
xnor U1471 (N_1471,N_947,N_765);
and U1472 (N_1472,N_799,N_889);
and U1473 (N_1473,N_802,N_555);
or U1474 (N_1474,N_591,N_546);
nor U1475 (N_1475,N_991,N_662);
and U1476 (N_1476,N_824,N_564);
nand U1477 (N_1477,N_690,N_839);
and U1478 (N_1478,N_879,N_585);
and U1479 (N_1479,N_517,N_729);
or U1480 (N_1480,N_558,N_717);
nand U1481 (N_1481,N_949,N_919);
or U1482 (N_1482,N_644,N_823);
or U1483 (N_1483,N_905,N_782);
nor U1484 (N_1484,N_944,N_537);
or U1485 (N_1485,N_828,N_840);
nor U1486 (N_1486,N_916,N_735);
nand U1487 (N_1487,N_653,N_959);
nand U1488 (N_1488,N_694,N_987);
nand U1489 (N_1489,N_998,N_877);
nand U1490 (N_1490,N_708,N_618);
or U1491 (N_1491,N_815,N_978);
nand U1492 (N_1492,N_831,N_859);
and U1493 (N_1493,N_530,N_628);
nor U1494 (N_1494,N_819,N_584);
nand U1495 (N_1495,N_515,N_545);
xor U1496 (N_1496,N_620,N_890);
nor U1497 (N_1497,N_573,N_938);
xnor U1498 (N_1498,N_516,N_645);
nand U1499 (N_1499,N_895,N_664);
nor U1500 (N_1500,N_1125,N_1254);
nand U1501 (N_1501,N_1466,N_1001);
and U1502 (N_1502,N_1338,N_1468);
nand U1503 (N_1503,N_1285,N_1036);
or U1504 (N_1504,N_1240,N_1180);
nand U1505 (N_1505,N_1273,N_1141);
and U1506 (N_1506,N_1089,N_1078);
xor U1507 (N_1507,N_1485,N_1426);
nand U1508 (N_1508,N_1386,N_1226);
nand U1509 (N_1509,N_1146,N_1460);
nor U1510 (N_1510,N_1073,N_1081);
nor U1511 (N_1511,N_1454,N_1390);
nand U1512 (N_1512,N_1418,N_1373);
xnor U1513 (N_1513,N_1147,N_1067);
nor U1514 (N_1514,N_1217,N_1307);
and U1515 (N_1515,N_1463,N_1409);
nor U1516 (N_1516,N_1308,N_1289);
or U1517 (N_1517,N_1145,N_1387);
and U1518 (N_1518,N_1206,N_1372);
nand U1519 (N_1519,N_1114,N_1247);
nand U1520 (N_1520,N_1100,N_1408);
and U1521 (N_1521,N_1119,N_1484);
xnor U1522 (N_1522,N_1221,N_1498);
or U1523 (N_1523,N_1276,N_1019);
nor U1524 (N_1524,N_1395,N_1382);
and U1525 (N_1525,N_1002,N_1261);
xor U1526 (N_1526,N_1295,N_1123);
and U1527 (N_1527,N_1300,N_1381);
and U1528 (N_1528,N_1269,N_1122);
and U1529 (N_1529,N_1199,N_1405);
and U1530 (N_1530,N_1057,N_1438);
nand U1531 (N_1531,N_1317,N_1369);
nand U1532 (N_1532,N_1437,N_1355);
nand U1533 (N_1533,N_1054,N_1026);
nand U1534 (N_1534,N_1050,N_1354);
nor U1535 (N_1535,N_1425,N_1106);
nor U1536 (N_1536,N_1434,N_1228);
nand U1537 (N_1537,N_1477,N_1190);
nor U1538 (N_1538,N_1275,N_1008);
and U1539 (N_1539,N_1197,N_1441);
nor U1540 (N_1540,N_1415,N_1065);
or U1541 (N_1541,N_1155,N_1037);
nand U1542 (N_1542,N_1350,N_1031);
nand U1543 (N_1543,N_1212,N_1222);
nor U1544 (N_1544,N_1284,N_1375);
and U1545 (N_1545,N_1492,N_1207);
nor U1546 (N_1546,N_1432,N_1393);
nand U1547 (N_1547,N_1262,N_1299);
nor U1548 (N_1548,N_1175,N_1274);
nand U1549 (N_1549,N_1430,N_1062);
and U1550 (N_1550,N_1227,N_1132);
and U1551 (N_1551,N_1322,N_1150);
nor U1552 (N_1552,N_1118,N_1185);
or U1553 (N_1553,N_1267,N_1076);
or U1554 (N_1554,N_1204,N_1191);
or U1555 (N_1555,N_1278,N_1263);
or U1556 (N_1556,N_1166,N_1052);
xnor U1557 (N_1557,N_1461,N_1332);
or U1558 (N_1558,N_1084,N_1211);
nor U1559 (N_1559,N_1178,N_1033);
nand U1560 (N_1560,N_1032,N_1245);
xnor U1561 (N_1561,N_1394,N_1069);
nand U1562 (N_1562,N_1347,N_1099);
nor U1563 (N_1563,N_1164,N_1007);
and U1564 (N_1564,N_1163,N_1096);
nand U1565 (N_1565,N_1324,N_1015);
and U1566 (N_1566,N_1223,N_1005);
and U1567 (N_1567,N_1287,N_1021);
and U1568 (N_1568,N_1348,N_1140);
xnor U1569 (N_1569,N_1170,N_1366);
or U1570 (N_1570,N_1205,N_1329);
or U1571 (N_1571,N_1494,N_1358);
and U1572 (N_1572,N_1041,N_1256);
and U1573 (N_1573,N_1156,N_1174);
xnor U1574 (N_1574,N_1169,N_1027);
nand U1575 (N_1575,N_1326,N_1202);
nand U1576 (N_1576,N_1234,N_1298);
and U1577 (N_1577,N_1391,N_1328);
or U1578 (N_1578,N_1231,N_1384);
nand U1579 (N_1579,N_1310,N_1412);
xor U1580 (N_1580,N_1377,N_1116);
or U1581 (N_1581,N_1229,N_1182);
xnor U1582 (N_1582,N_1286,N_1124);
and U1583 (N_1583,N_1060,N_1055);
and U1584 (N_1584,N_1104,N_1203);
nand U1585 (N_1585,N_1351,N_1220);
nand U1586 (N_1586,N_1362,N_1070);
and U1587 (N_1587,N_1135,N_1165);
nor U1588 (N_1588,N_1105,N_1490);
nand U1589 (N_1589,N_1445,N_1480);
nand U1590 (N_1590,N_1396,N_1277);
or U1591 (N_1591,N_1109,N_1340);
nor U1592 (N_1592,N_1149,N_1216);
or U1593 (N_1593,N_1473,N_1266);
nand U1594 (N_1594,N_1115,N_1148);
nand U1595 (N_1595,N_1143,N_1176);
nand U1596 (N_1596,N_1380,N_1092);
and U1597 (N_1597,N_1242,N_1399);
xnor U1598 (N_1598,N_1077,N_1435);
xnor U1599 (N_1599,N_1456,N_1080);
or U1600 (N_1600,N_1248,N_1499);
and U1601 (N_1601,N_1496,N_1359);
nor U1602 (N_1602,N_1258,N_1268);
nand U1603 (N_1603,N_1038,N_1431);
nor U1604 (N_1604,N_1043,N_1474);
nor U1605 (N_1605,N_1087,N_1194);
xnor U1606 (N_1606,N_1264,N_1016);
or U1607 (N_1607,N_1012,N_1424);
and U1608 (N_1608,N_1225,N_1341);
or U1609 (N_1609,N_1091,N_1304);
nor U1610 (N_1610,N_1028,N_1446);
nand U1611 (N_1611,N_1337,N_1257);
xor U1612 (N_1612,N_1422,N_1279);
nor U1613 (N_1613,N_1113,N_1379);
nand U1614 (N_1614,N_1058,N_1400);
and U1615 (N_1615,N_1365,N_1401);
and U1616 (N_1616,N_1112,N_1051);
nor U1617 (N_1617,N_1406,N_1253);
and U1618 (N_1618,N_1068,N_1283);
or U1619 (N_1619,N_1158,N_1160);
and U1620 (N_1620,N_1196,N_1029);
and U1621 (N_1621,N_1093,N_1181);
or U1622 (N_1622,N_1357,N_1108);
nor U1623 (N_1623,N_1018,N_1364);
nand U1624 (N_1624,N_1459,N_1318);
and U1625 (N_1625,N_1342,N_1288);
nor U1626 (N_1626,N_1173,N_1239);
or U1627 (N_1627,N_1294,N_1404);
or U1628 (N_1628,N_1361,N_1339);
or U1629 (N_1629,N_1030,N_1352);
nor U1630 (N_1630,N_1013,N_1309);
or U1631 (N_1631,N_1088,N_1133);
nor U1632 (N_1632,N_1320,N_1259);
and U1633 (N_1633,N_1255,N_1376);
and U1634 (N_1634,N_1414,N_1045);
xnor U1635 (N_1635,N_1230,N_1444);
xor U1636 (N_1636,N_1171,N_1440);
nor U1637 (N_1637,N_1144,N_1172);
and U1638 (N_1638,N_1004,N_1235);
nor U1639 (N_1639,N_1271,N_1388);
nor U1640 (N_1640,N_1331,N_1048);
nor U1641 (N_1641,N_1243,N_1383);
nand U1642 (N_1642,N_1327,N_1233);
and U1643 (N_1643,N_1035,N_1022);
nor U1644 (N_1644,N_1017,N_1210);
and U1645 (N_1645,N_1086,N_1291);
nor U1646 (N_1646,N_1407,N_1471);
nand U1647 (N_1647,N_1345,N_1218);
nor U1648 (N_1648,N_1046,N_1305);
nor U1649 (N_1649,N_1039,N_1385);
xor U1650 (N_1650,N_1064,N_1389);
or U1651 (N_1651,N_1419,N_1107);
and U1652 (N_1652,N_1198,N_1421);
and U1653 (N_1653,N_1465,N_1134);
and U1654 (N_1654,N_1486,N_1201);
nand U1655 (N_1655,N_1219,N_1209);
and U1656 (N_1656,N_1398,N_1493);
nand U1657 (N_1657,N_1478,N_1292);
or U1658 (N_1658,N_1270,N_1168);
nand U1659 (N_1659,N_1489,N_1138);
or U1660 (N_1660,N_1189,N_1157);
nand U1661 (N_1661,N_1436,N_1397);
nand U1662 (N_1662,N_1470,N_1102);
nor U1663 (N_1663,N_1006,N_1334);
or U1664 (N_1664,N_1469,N_1371);
nor U1665 (N_1665,N_1392,N_1303);
nor U1666 (N_1666,N_1402,N_1323);
and U1667 (N_1667,N_1413,N_1117);
or U1668 (N_1668,N_1244,N_1000);
xnor U1669 (N_1669,N_1250,N_1416);
or U1670 (N_1670,N_1479,N_1301);
nand U1671 (N_1671,N_1442,N_1333);
or U1672 (N_1672,N_1097,N_1003);
or U1673 (N_1673,N_1159,N_1183);
nand U1674 (N_1674,N_1136,N_1154);
and U1675 (N_1675,N_1049,N_1251);
nor U1676 (N_1676,N_1495,N_1103);
nor U1677 (N_1677,N_1417,N_1040);
nor U1678 (N_1678,N_1177,N_1448);
nor U1679 (N_1679,N_1346,N_1137);
nand U1680 (N_1680,N_1410,N_1316);
and U1681 (N_1681,N_1467,N_1314);
or U1682 (N_1682,N_1186,N_1367);
or U1683 (N_1683,N_1451,N_1429);
nand U1684 (N_1684,N_1014,N_1293);
nor U1685 (N_1685,N_1455,N_1472);
and U1686 (N_1686,N_1192,N_1476);
or U1687 (N_1687,N_1142,N_1208);
nor U1688 (N_1688,N_1297,N_1025);
nor U1689 (N_1689,N_1457,N_1462);
or U1690 (N_1690,N_1311,N_1187);
and U1691 (N_1691,N_1120,N_1330);
or U1692 (N_1692,N_1296,N_1433);
nand U1693 (N_1693,N_1010,N_1075);
or U1694 (N_1694,N_1281,N_1428);
nand U1695 (N_1695,N_1056,N_1335);
xor U1696 (N_1696,N_1167,N_1024);
xor U1697 (N_1697,N_1047,N_1153);
nand U1698 (N_1698,N_1129,N_1059);
and U1699 (N_1699,N_1249,N_1127);
and U1700 (N_1700,N_1082,N_1312);
xnor U1701 (N_1701,N_1272,N_1403);
or U1702 (N_1702,N_1237,N_1265);
and U1703 (N_1703,N_1363,N_1184);
nor U1704 (N_1704,N_1370,N_1213);
nand U1705 (N_1705,N_1095,N_1193);
nand U1706 (N_1706,N_1356,N_1321);
or U1707 (N_1707,N_1121,N_1344);
nor U1708 (N_1708,N_1319,N_1343);
and U1709 (N_1709,N_1487,N_1475);
or U1710 (N_1710,N_1483,N_1491);
nand U1711 (N_1711,N_1071,N_1450);
or U1712 (N_1712,N_1290,N_1034);
or U1713 (N_1713,N_1053,N_1368);
and U1714 (N_1714,N_1110,N_1325);
nor U1715 (N_1715,N_1161,N_1306);
xnor U1716 (N_1716,N_1481,N_1411);
and U1717 (N_1717,N_1151,N_1083);
or U1718 (N_1718,N_1280,N_1066);
and U1719 (N_1719,N_1179,N_1315);
or U1720 (N_1720,N_1200,N_1488);
and U1721 (N_1721,N_1313,N_1360);
and U1722 (N_1722,N_1111,N_1302);
xor U1723 (N_1723,N_1098,N_1464);
or U1724 (N_1724,N_1238,N_1232);
and U1725 (N_1725,N_1374,N_1353);
nor U1726 (N_1726,N_1152,N_1139);
xnor U1727 (N_1727,N_1128,N_1447);
nor U1728 (N_1728,N_1215,N_1252);
nand U1729 (N_1729,N_1009,N_1427);
nand U1730 (N_1730,N_1042,N_1453);
and U1731 (N_1731,N_1282,N_1236);
nor U1732 (N_1732,N_1101,N_1336);
or U1733 (N_1733,N_1423,N_1126);
nor U1734 (N_1734,N_1072,N_1214);
or U1735 (N_1735,N_1131,N_1094);
and U1736 (N_1736,N_1130,N_1378);
nand U1737 (N_1737,N_1452,N_1241);
nor U1738 (N_1738,N_1090,N_1420);
and U1739 (N_1739,N_1224,N_1085);
nand U1740 (N_1740,N_1074,N_1439);
or U1741 (N_1741,N_1497,N_1195);
nor U1742 (N_1742,N_1246,N_1449);
nor U1743 (N_1743,N_1023,N_1044);
nand U1744 (N_1744,N_1349,N_1061);
and U1745 (N_1745,N_1162,N_1063);
nand U1746 (N_1746,N_1443,N_1458);
or U1747 (N_1747,N_1482,N_1079);
and U1748 (N_1748,N_1020,N_1011);
and U1749 (N_1749,N_1188,N_1260);
and U1750 (N_1750,N_1433,N_1263);
or U1751 (N_1751,N_1468,N_1414);
nand U1752 (N_1752,N_1012,N_1035);
xnor U1753 (N_1753,N_1487,N_1189);
nand U1754 (N_1754,N_1348,N_1209);
nor U1755 (N_1755,N_1282,N_1437);
xor U1756 (N_1756,N_1075,N_1338);
nor U1757 (N_1757,N_1367,N_1047);
nor U1758 (N_1758,N_1165,N_1003);
nor U1759 (N_1759,N_1460,N_1000);
or U1760 (N_1760,N_1219,N_1281);
or U1761 (N_1761,N_1121,N_1271);
nor U1762 (N_1762,N_1110,N_1455);
nor U1763 (N_1763,N_1355,N_1230);
nand U1764 (N_1764,N_1277,N_1264);
or U1765 (N_1765,N_1470,N_1176);
nor U1766 (N_1766,N_1082,N_1202);
nor U1767 (N_1767,N_1276,N_1230);
xnor U1768 (N_1768,N_1009,N_1432);
or U1769 (N_1769,N_1140,N_1471);
nand U1770 (N_1770,N_1101,N_1058);
or U1771 (N_1771,N_1425,N_1342);
and U1772 (N_1772,N_1374,N_1132);
nor U1773 (N_1773,N_1257,N_1329);
and U1774 (N_1774,N_1332,N_1274);
nand U1775 (N_1775,N_1480,N_1034);
nor U1776 (N_1776,N_1342,N_1107);
nor U1777 (N_1777,N_1130,N_1123);
or U1778 (N_1778,N_1219,N_1449);
nor U1779 (N_1779,N_1098,N_1447);
and U1780 (N_1780,N_1413,N_1324);
or U1781 (N_1781,N_1258,N_1434);
or U1782 (N_1782,N_1387,N_1165);
nand U1783 (N_1783,N_1049,N_1025);
nand U1784 (N_1784,N_1041,N_1430);
nor U1785 (N_1785,N_1096,N_1098);
nand U1786 (N_1786,N_1429,N_1473);
or U1787 (N_1787,N_1082,N_1034);
and U1788 (N_1788,N_1461,N_1044);
nor U1789 (N_1789,N_1298,N_1205);
or U1790 (N_1790,N_1207,N_1124);
and U1791 (N_1791,N_1245,N_1311);
nor U1792 (N_1792,N_1293,N_1323);
nor U1793 (N_1793,N_1296,N_1088);
and U1794 (N_1794,N_1263,N_1194);
and U1795 (N_1795,N_1479,N_1096);
nand U1796 (N_1796,N_1132,N_1326);
nor U1797 (N_1797,N_1081,N_1399);
or U1798 (N_1798,N_1228,N_1295);
or U1799 (N_1799,N_1146,N_1016);
nand U1800 (N_1800,N_1380,N_1160);
nor U1801 (N_1801,N_1289,N_1414);
nand U1802 (N_1802,N_1091,N_1348);
xor U1803 (N_1803,N_1333,N_1001);
nand U1804 (N_1804,N_1167,N_1235);
nand U1805 (N_1805,N_1384,N_1274);
nand U1806 (N_1806,N_1014,N_1320);
and U1807 (N_1807,N_1281,N_1111);
or U1808 (N_1808,N_1308,N_1160);
and U1809 (N_1809,N_1445,N_1341);
and U1810 (N_1810,N_1189,N_1004);
nor U1811 (N_1811,N_1409,N_1156);
nor U1812 (N_1812,N_1194,N_1473);
nand U1813 (N_1813,N_1286,N_1062);
xnor U1814 (N_1814,N_1037,N_1371);
nand U1815 (N_1815,N_1444,N_1104);
nand U1816 (N_1816,N_1253,N_1256);
or U1817 (N_1817,N_1223,N_1055);
nor U1818 (N_1818,N_1492,N_1483);
nor U1819 (N_1819,N_1343,N_1494);
nand U1820 (N_1820,N_1388,N_1457);
or U1821 (N_1821,N_1464,N_1306);
or U1822 (N_1822,N_1242,N_1112);
nand U1823 (N_1823,N_1362,N_1433);
nand U1824 (N_1824,N_1114,N_1027);
or U1825 (N_1825,N_1101,N_1132);
nand U1826 (N_1826,N_1289,N_1494);
and U1827 (N_1827,N_1220,N_1273);
nor U1828 (N_1828,N_1332,N_1474);
and U1829 (N_1829,N_1495,N_1283);
nor U1830 (N_1830,N_1260,N_1147);
or U1831 (N_1831,N_1249,N_1365);
nand U1832 (N_1832,N_1315,N_1168);
nor U1833 (N_1833,N_1161,N_1223);
nor U1834 (N_1834,N_1402,N_1320);
or U1835 (N_1835,N_1493,N_1235);
and U1836 (N_1836,N_1234,N_1288);
nand U1837 (N_1837,N_1242,N_1150);
nand U1838 (N_1838,N_1117,N_1012);
or U1839 (N_1839,N_1164,N_1011);
xnor U1840 (N_1840,N_1325,N_1045);
and U1841 (N_1841,N_1072,N_1067);
and U1842 (N_1842,N_1382,N_1007);
nand U1843 (N_1843,N_1227,N_1405);
or U1844 (N_1844,N_1155,N_1172);
and U1845 (N_1845,N_1381,N_1295);
xor U1846 (N_1846,N_1297,N_1435);
nand U1847 (N_1847,N_1428,N_1461);
nand U1848 (N_1848,N_1426,N_1279);
or U1849 (N_1849,N_1103,N_1297);
nand U1850 (N_1850,N_1191,N_1475);
nor U1851 (N_1851,N_1104,N_1188);
or U1852 (N_1852,N_1451,N_1265);
nand U1853 (N_1853,N_1413,N_1394);
nor U1854 (N_1854,N_1372,N_1183);
and U1855 (N_1855,N_1331,N_1024);
or U1856 (N_1856,N_1420,N_1294);
or U1857 (N_1857,N_1498,N_1408);
or U1858 (N_1858,N_1078,N_1307);
and U1859 (N_1859,N_1279,N_1148);
nor U1860 (N_1860,N_1007,N_1290);
nand U1861 (N_1861,N_1015,N_1040);
and U1862 (N_1862,N_1264,N_1146);
and U1863 (N_1863,N_1320,N_1152);
nor U1864 (N_1864,N_1190,N_1218);
and U1865 (N_1865,N_1121,N_1455);
nor U1866 (N_1866,N_1157,N_1402);
nor U1867 (N_1867,N_1203,N_1136);
nor U1868 (N_1868,N_1362,N_1438);
nor U1869 (N_1869,N_1297,N_1284);
nor U1870 (N_1870,N_1250,N_1045);
nand U1871 (N_1871,N_1069,N_1492);
or U1872 (N_1872,N_1443,N_1493);
and U1873 (N_1873,N_1440,N_1262);
nand U1874 (N_1874,N_1394,N_1496);
and U1875 (N_1875,N_1414,N_1128);
or U1876 (N_1876,N_1206,N_1351);
or U1877 (N_1877,N_1147,N_1499);
nand U1878 (N_1878,N_1194,N_1327);
nand U1879 (N_1879,N_1253,N_1287);
and U1880 (N_1880,N_1162,N_1174);
and U1881 (N_1881,N_1313,N_1413);
and U1882 (N_1882,N_1156,N_1129);
nand U1883 (N_1883,N_1231,N_1207);
and U1884 (N_1884,N_1205,N_1069);
and U1885 (N_1885,N_1264,N_1324);
nor U1886 (N_1886,N_1077,N_1069);
nand U1887 (N_1887,N_1022,N_1312);
and U1888 (N_1888,N_1195,N_1391);
and U1889 (N_1889,N_1303,N_1388);
nor U1890 (N_1890,N_1209,N_1154);
nor U1891 (N_1891,N_1277,N_1028);
and U1892 (N_1892,N_1439,N_1213);
nand U1893 (N_1893,N_1431,N_1165);
or U1894 (N_1894,N_1439,N_1391);
and U1895 (N_1895,N_1281,N_1464);
nand U1896 (N_1896,N_1311,N_1294);
or U1897 (N_1897,N_1161,N_1139);
and U1898 (N_1898,N_1417,N_1232);
and U1899 (N_1899,N_1355,N_1038);
and U1900 (N_1900,N_1173,N_1316);
xnor U1901 (N_1901,N_1290,N_1141);
xnor U1902 (N_1902,N_1259,N_1403);
or U1903 (N_1903,N_1410,N_1336);
nor U1904 (N_1904,N_1228,N_1315);
or U1905 (N_1905,N_1489,N_1362);
and U1906 (N_1906,N_1390,N_1245);
nor U1907 (N_1907,N_1136,N_1491);
nand U1908 (N_1908,N_1484,N_1141);
nand U1909 (N_1909,N_1288,N_1082);
nand U1910 (N_1910,N_1253,N_1429);
nand U1911 (N_1911,N_1424,N_1040);
or U1912 (N_1912,N_1245,N_1055);
nor U1913 (N_1913,N_1161,N_1112);
or U1914 (N_1914,N_1341,N_1339);
nand U1915 (N_1915,N_1004,N_1280);
and U1916 (N_1916,N_1233,N_1250);
and U1917 (N_1917,N_1050,N_1331);
nand U1918 (N_1918,N_1353,N_1133);
nand U1919 (N_1919,N_1404,N_1491);
nand U1920 (N_1920,N_1151,N_1091);
and U1921 (N_1921,N_1212,N_1469);
or U1922 (N_1922,N_1025,N_1219);
nand U1923 (N_1923,N_1475,N_1291);
nor U1924 (N_1924,N_1158,N_1370);
nand U1925 (N_1925,N_1272,N_1459);
xnor U1926 (N_1926,N_1101,N_1051);
or U1927 (N_1927,N_1326,N_1176);
or U1928 (N_1928,N_1372,N_1141);
nor U1929 (N_1929,N_1248,N_1489);
nand U1930 (N_1930,N_1246,N_1083);
or U1931 (N_1931,N_1494,N_1254);
nor U1932 (N_1932,N_1473,N_1038);
or U1933 (N_1933,N_1393,N_1024);
nand U1934 (N_1934,N_1365,N_1460);
and U1935 (N_1935,N_1293,N_1104);
nand U1936 (N_1936,N_1499,N_1392);
and U1937 (N_1937,N_1304,N_1181);
nand U1938 (N_1938,N_1071,N_1348);
xor U1939 (N_1939,N_1131,N_1177);
nand U1940 (N_1940,N_1328,N_1344);
or U1941 (N_1941,N_1430,N_1266);
or U1942 (N_1942,N_1453,N_1237);
or U1943 (N_1943,N_1020,N_1084);
nor U1944 (N_1944,N_1065,N_1402);
or U1945 (N_1945,N_1238,N_1202);
or U1946 (N_1946,N_1428,N_1221);
xnor U1947 (N_1947,N_1096,N_1273);
and U1948 (N_1948,N_1143,N_1471);
nor U1949 (N_1949,N_1297,N_1274);
or U1950 (N_1950,N_1126,N_1449);
nand U1951 (N_1951,N_1463,N_1370);
nor U1952 (N_1952,N_1366,N_1294);
xor U1953 (N_1953,N_1096,N_1305);
and U1954 (N_1954,N_1018,N_1166);
nor U1955 (N_1955,N_1335,N_1389);
or U1956 (N_1956,N_1382,N_1376);
and U1957 (N_1957,N_1462,N_1467);
nand U1958 (N_1958,N_1499,N_1247);
nand U1959 (N_1959,N_1420,N_1038);
or U1960 (N_1960,N_1351,N_1300);
nand U1961 (N_1961,N_1002,N_1182);
or U1962 (N_1962,N_1060,N_1402);
or U1963 (N_1963,N_1225,N_1296);
or U1964 (N_1964,N_1383,N_1321);
xnor U1965 (N_1965,N_1112,N_1279);
and U1966 (N_1966,N_1103,N_1104);
nand U1967 (N_1967,N_1408,N_1441);
and U1968 (N_1968,N_1410,N_1248);
xor U1969 (N_1969,N_1284,N_1113);
or U1970 (N_1970,N_1387,N_1427);
and U1971 (N_1971,N_1466,N_1495);
or U1972 (N_1972,N_1483,N_1165);
and U1973 (N_1973,N_1299,N_1219);
or U1974 (N_1974,N_1089,N_1086);
and U1975 (N_1975,N_1370,N_1157);
and U1976 (N_1976,N_1414,N_1190);
or U1977 (N_1977,N_1240,N_1167);
nor U1978 (N_1978,N_1389,N_1357);
or U1979 (N_1979,N_1441,N_1335);
nor U1980 (N_1980,N_1169,N_1297);
or U1981 (N_1981,N_1411,N_1026);
and U1982 (N_1982,N_1360,N_1372);
and U1983 (N_1983,N_1202,N_1015);
and U1984 (N_1984,N_1171,N_1076);
nor U1985 (N_1985,N_1249,N_1308);
and U1986 (N_1986,N_1439,N_1264);
nor U1987 (N_1987,N_1477,N_1094);
nand U1988 (N_1988,N_1071,N_1230);
nor U1989 (N_1989,N_1284,N_1280);
and U1990 (N_1990,N_1428,N_1184);
nor U1991 (N_1991,N_1432,N_1181);
and U1992 (N_1992,N_1349,N_1394);
nand U1993 (N_1993,N_1481,N_1320);
nor U1994 (N_1994,N_1164,N_1075);
xnor U1995 (N_1995,N_1412,N_1122);
and U1996 (N_1996,N_1204,N_1491);
or U1997 (N_1997,N_1119,N_1235);
nor U1998 (N_1998,N_1074,N_1131);
or U1999 (N_1999,N_1035,N_1414);
nand U2000 (N_2000,N_1517,N_1601);
or U2001 (N_2001,N_1902,N_1520);
nand U2002 (N_2002,N_1782,N_1528);
nor U2003 (N_2003,N_1732,N_1534);
or U2004 (N_2004,N_1752,N_1717);
nor U2005 (N_2005,N_1816,N_1635);
nor U2006 (N_2006,N_1718,N_1956);
and U2007 (N_2007,N_1770,N_1771);
or U2008 (N_2008,N_1990,N_1598);
or U2009 (N_2009,N_1772,N_1536);
or U2010 (N_2010,N_1998,N_1865);
nor U2011 (N_2011,N_1632,N_1693);
nor U2012 (N_2012,N_1648,N_1863);
or U2013 (N_2013,N_1791,N_1574);
and U2014 (N_2014,N_1906,N_1814);
nand U2015 (N_2015,N_1750,N_1530);
nand U2016 (N_2016,N_1868,N_1954);
nand U2017 (N_2017,N_1897,N_1636);
nor U2018 (N_2018,N_1774,N_1503);
xor U2019 (N_2019,N_1886,N_1871);
nand U2020 (N_2020,N_1920,N_1657);
or U2021 (N_2021,N_1812,N_1555);
nand U2022 (N_2022,N_1795,N_1662);
nand U2023 (N_2023,N_1987,N_1725);
xnor U2024 (N_2024,N_1653,N_1899);
nor U2025 (N_2025,N_1842,N_1753);
or U2026 (N_2026,N_1896,N_1714);
nand U2027 (N_2027,N_1834,N_1595);
nor U2028 (N_2028,N_1828,N_1959);
nor U2029 (N_2029,N_1720,N_1594);
nor U2030 (N_2030,N_1824,N_1641);
nor U2031 (N_2031,N_1997,N_1850);
nor U2032 (N_2032,N_1889,N_1739);
and U2033 (N_2033,N_1529,N_1869);
nand U2034 (N_2034,N_1887,N_1908);
or U2035 (N_2035,N_1845,N_1599);
and U2036 (N_2036,N_1973,N_1966);
nand U2037 (N_2037,N_1822,N_1736);
or U2038 (N_2038,N_1805,N_1874);
and U2039 (N_2039,N_1619,N_1836);
nor U2040 (N_2040,N_1958,N_1832);
xor U2041 (N_2041,N_1769,N_1557);
nand U2042 (N_2042,N_1623,N_1751);
nand U2043 (N_2043,N_1553,N_1875);
or U2044 (N_2044,N_1661,N_1705);
and U2045 (N_2045,N_1934,N_1674);
or U2046 (N_2046,N_1811,N_1540);
and U2047 (N_2047,N_1737,N_1668);
nand U2048 (N_2048,N_1986,N_1999);
nand U2049 (N_2049,N_1846,N_1700);
and U2050 (N_2050,N_1904,N_1565);
nor U2051 (N_2051,N_1698,N_1515);
or U2052 (N_2052,N_1537,N_1918);
nor U2053 (N_2053,N_1708,N_1792);
nor U2054 (N_2054,N_1793,N_1633);
or U2055 (N_2055,N_1531,N_1905);
nand U2056 (N_2056,N_1643,N_1608);
nor U2057 (N_2057,N_1687,N_1963);
nor U2058 (N_2058,N_1734,N_1815);
and U2059 (N_2059,N_1640,N_1860);
or U2060 (N_2060,N_1600,N_1722);
or U2061 (N_2061,N_1511,N_1941);
nand U2062 (N_2062,N_1932,N_1937);
xor U2063 (N_2063,N_1981,N_1843);
or U2064 (N_2064,N_1803,N_1768);
nor U2065 (N_2065,N_1879,N_1820);
or U2066 (N_2066,N_1676,N_1888);
and U2067 (N_2067,N_1776,N_1525);
nor U2068 (N_2068,N_1796,N_1710);
and U2069 (N_2069,N_1799,N_1882);
and U2070 (N_2070,N_1677,N_1802);
or U2071 (N_2071,N_1910,N_1707);
or U2072 (N_2072,N_1898,N_1609);
nand U2073 (N_2073,N_1507,N_1764);
and U2074 (N_2074,N_1506,N_1585);
xor U2075 (N_2075,N_1561,N_1575);
or U2076 (N_2076,N_1929,N_1712);
nand U2077 (N_2077,N_1994,N_1983);
and U2078 (N_2078,N_1518,N_1709);
and U2079 (N_2079,N_1502,N_1829);
and U2080 (N_2080,N_1978,N_1762);
or U2081 (N_2081,N_1780,N_1819);
nand U2082 (N_2082,N_1616,N_1790);
nor U2083 (N_2083,N_1942,N_1613);
nand U2084 (N_2084,N_1610,N_1781);
or U2085 (N_2085,N_1852,N_1629);
or U2086 (N_2086,N_1991,N_1532);
and U2087 (N_2087,N_1590,N_1581);
xnor U2088 (N_2088,N_1833,N_1509);
nor U2089 (N_2089,N_1678,N_1578);
and U2090 (N_2090,N_1808,N_1579);
and U2091 (N_2091,N_1965,N_1731);
or U2092 (N_2092,N_1697,N_1719);
xor U2093 (N_2093,N_1630,N_1961);
nor U2094 (N_2094,N_1622,N_1873);
nand U2095 (N_2095,N_1658,N_1851);
nor U2096 (N_2096,N_1522,N_1542);
or U2097 (N_2097,N_1703,N_1759);
or U2098 (N_2098,N_1947,N_1858);
and U2099 (N_2099,N_1746,N_1827);
and U2100 (N_2100,N_1938,N_1901);
or U2101 (N_2101,N_1713,N_1556);
and U2102 (N_2102,N_1749,N_1952);
nor U2103 (N_2103,N_1686,N_1597);
and U2104 (N_2104,N_1931,N_1784);
and U2105 (N_2105,N_1683,N_1501);
and U2106 (N_2106,N_1951,N_1779);
nand U2107 (N_2107,N_1651,N_1625);
and U2108 (N_2108,N_1924,N_1979);
nor U2109 (N_2109,N_1883,N_1925);
nor U2110 (N_2110,N_1554,N_1831);
or U2111 (N_2111,N_1618,N_1847);
and U2112 (N_2112,N_1809,N_1785);
and U2113 (N_2113,N_1583,N_1928);
and U2114 (N_2114,N_1996,N_1968);
or U2115 (N_2115,N_1923,N_1969);
nor U2116 (N_2116,N_1577,N_1587);
nor U2117 (N_2117,N_1558,N_1611);
and U2118 (N_2118,N_1573,N_1562);
and U2119 (N_2119,N_1706,N_1867);
xnor U2120 (N_2120,N_1605,N_1907);
nor U2121 (N_2121,N_1945,N_1870);
or U2122 (N_2122,N_1591,N_1624);
nand U2123 (N_2123,N_1724,N_1620);
and U2124 (N_2124,N_1637,N_1631);
and U2125 (N_2125,N_1786,N_1716);
or U2126 (N_2126,N_1754,N_1854);
or U2127 (N_2127,N_1733,N_1543);
or U2128 (N_2128,N_1593,N_1545);
and U2129 (N_2129,N_1549,N_1756);
nor U2130 (N_2130,N_1895,N_1841);
or U2131 (N_2131,N_1681,N_1992);
nand U2132 (N_2132,N_1919,N_1612);
nand U2133 (N_2133,N_1989,N_1659);
nand U2134 (N_2134,N_1500,N_1665);
and U2135 (N_2135,N_1894,N_1626);
xnor U2136 (N_2136,N_1670,N_1943);
nand U2137 (N_2137,N_1566,N_1933);
and U2138 (N_2138,N_1711,N_1589);
nor U2139 (N_2139,N_1950,N_1614);
or U2140 (N_2140,N_1917,N_1721);
or U2141 (N_2141,N_1984,N_1855);
or U2142 (N_2142,N_1849,N_1830);
nor U2143 (N_2143,N_1767,N_1813);
nand U2144 (N_2144,N_1976,N_1758);
nor U2145 (N_2145,N_1970,N_1604);
or U2146 (N_2146,N_1563,N_1881);
or U2147 (N_2147,N_1508,N_1837);
and U2148 (N_2148,N_1726,N_1539);
and U2149 (N_2149,N_1744,N_1663);
nor U2150 (N_2150,N_1794,N_1909);
nor U2151 (N_2151,N_1957,N_1864);
or U2152 (N_2152,N_1944,N_1922);
and U2153 (N_2153,N_1695,N_1946);
nor U2154 (N_2154,N_1660,N_1694);
or U2155 (N_2155,N_1513,N_1877);
nand U2156 (N_2156,N_1835,N_1747);
and U2157 (N_2157,N_1646,N_1582);
nand U2158 (N_2158,N_1916,N_1972);
nand U2159 (N_2159,N_1914,N_1738);
nand U2160 (N_2160,N_1757,N_1584);
nand U2161 (N_2161,N_1818,N_1891);
or U2162 (N_2162,N_1890,N_1804);
nor U2163 (N_2163,N_1866,N_1642);
and U2164 (N_2164,N_1729,N_1592);
xnor U2165 (N_2165,N_1655,N_1702);
nand U2166 (N_2166,N_1995,N_1826);
nand U2167 (N_2167,N_1519,N_1844);
nand U2168 (N_2168,N_1892,N_1621);
or U2169 (N_2169,N_1823,N_1948);
or U2170 (N_2170,N_1634,N_1701);
or U2171 (N_2171,N_1921,N_1541);
xor U2172 (N_2172,N_1735,N_1748);
nor U2173 (N_2173,N_1505,N_1940);
nor U2174 (N_2174,N_1760,N_1912);
nand U2175 (N_2175,N_1699,N_1967);
or U2176 (N_2176,N_1672,N_1872);
and U2177 (N_2177,N_1862,N_1740);
nand U2178 (N_2178,N_1654,N_1690);
nand U2179 (N_2179,N_1988,N_1730);
nand U2180 (N_2180,N_1962,N_1533);
nor U2181 (N_2181,N_1666,N_1569);
nand U2182 (N_2182,N_1885,N_1688);
nor U2183 (N_2183,N_1806,N_1807);
nand U2184 (N_2184,N_1568,N_1971);
nand U2185 (N_2185,N_1656,N_1913);
nand U2186 (N_2186,N_1572,N_1810);
or U2187 (N_2187,N_1783,N_1673);
and U2188 (N_2188,N_1607,N_1664);
nand U2189 (N_2189,N_1787,N_1848);
xnor U2190 (N_2190,N_1627,N_1975);
and U2191 (N_2191,N_1544,N_1715);
nand U2192 (N_2192,N_1982,N_1761);
nand U2193 (N_2193,N_1953,N_1580);
and U2194 (N_2194,N_1884,N_1588);
and U2195 (N_2195,N_1977,N_1876);
nand U2196 (N_2196,N_1689,N_1777);
and U2197 (N_2197,N_1801,N_1974);
nor U2198 (N_2198,N_1667,N_1857);
or U2199 (N_2199,N_1685,N_1900);
nand U2200 (N_2200,N_1853,N_1949);
nor U2201 (N_2201,N_1838,N_1617);
nor U2202 (N_2202,N_1684,N_1504);
xnor U2203 (N_2203,N_1644,N_1559);
nand U2204 (N_2204,N_1880,N_1742);
nor U2205 (N_2205,N_1727,N_1915);
or U2206 (N_2206,N_1980,N_1548);
nand U2207 (N_2207,N_1510,N_1669);
or U2208 (N_2208,N_1798,N_1741);
nor U2209 (N_2209,N_1650,N_1955);
or U2210 (N_2210,N_1516,N_1535);
xnor U2211 (N_2211,N_1586,N_1527);
and U2212 (N_2212,N_1765,N_1692);
and U2213 (N_2213,N_1723,N_1512);
nor U2214 (N_2214,N_1745,N_1691);
nand U2215 (N_2215,N_1679,N_1839);
or U2216 (N_2216,N_1766,N_1960);
xor U2217 (N_2217,N_1817,N_1645);
nor U2218 (N_2218,N_1936,N_1671);
nand U2219 (N_2219,N_1821,N_1606);
nand U2220 (N_2220,N_1524,N_1800);
nor U2221 (N_2221,N_1675,N_1680);
or U2222 (N_2222,N_1570,N_1514);
or U2223 (N_2223,N_1704,N_1840);
or U2224 (N_2224,N_1538,N_1521);
and U2225 (N_2225,N_1523,N_1985);
xor U2226 (N_2226,N_1893,N_1927);
or U2227 (N_2227,N_1571,N_1775);
and U2228 (N_2228,N_1926,N_1550);
nand U2229 (N_2229,N_1547,N_1564);
nand U2230 (N_2230,N_1773,N_1576);
or U2231 (N_2231,N_1560,N_1859);
nand U2232 (N_2232,N_1789,N_1649);
and U2233 (N_2233,N_1825,N_1743);
and U2234 (N_2234,N_1552,N_1911);
and U2235 (N_2235,N_1652,N_1567);
and U2236 (N_2236,N_1551,N_1696);
xnor U2237 (N_2237,N_1763,N_1546);
nand U2238 (N_2238,N_1856,N_1647);
nor U2239 (N_2239,N_1728,N_1993);
nor U2240 (N_2240,N_1964,N_1861);
xnor U2241 (N_2241,N_1682,N_1639);
nand U2242 (N_2242,N_1797,N_1526);
nand U2243 (N_2243,N_1603,N_1615);
and U2244 (N_2244,N_1778,N_1939);
or U2245 (N_2245,N_1930,N_1596);
and U2246 (N_2246,N_1788,N_1935);
nor U2247 (N_2247,N_1602,N_1628);
nor U2248 (N_2248,N_1755,N_1638);
nor U2249 (N_2249,N_1878,N_1903);
or U2250 (N_2250,N_1966,N_1597);
nor U2251 (N_2251,N_1764,N_1980);
nor U2252 (N_2252,N_1848,N_1528);
and U2253 (N_2253,N_1674,N_1548);
or U2254 (N_2254,N_1788,N_1776);
or U2255 (N_2255,N_1688,N_1744);
nor U2256 (N_2256,N_1829,N_1596);
nand U2257 (N_2257,N_1617,N_1761);
nor U2258 (N_2258,N_1714,N_1764);
or U2259 (N_2259,N_1952,N_1875);
nand U2260 (N_2260,N_1583,N_1863);
nor U2261 (N_2261,N_1637,N_1602);
nand U2262 (N_2262,N_1894,N_1827);
nor U2263 (N_2263,N_1985,N_1533);
nand U2264 (N_2264,N_1894,N_1608);
or U2265 (N_2265,N_1896,N_1803);
or U2266 (N_2266,N_1566,N_1980);
nand U2267 (N_2267,N_1527,N_1658);
xor U2268 (N_2268,N_1930,N_1791);
and U2269 (N_2269,N_1554,N_1514);
nor U2270 (N_2270,N_1684,N_1549);
nor U2271 (N_2271,N_1706,N_1905);
or U2272 (N_2272,N_1548,N_1560);
or U2273 (N_2273,N_1978,N_1967);
nor U2274 (N_2274,N_1808,N_1632);
xnor U2275 (N_2275,N_1979,N_1961);
xnor U2276 (N_2276,N_1615,N_1851);
or U2277 (N_2277,N_1907,N_1893);
or U2278 (N_2278,N_1899,N_1505);
nor U2279 (N_2279,N_1987,N_1824);
nor U2280 (N_2280,N_1895,N_1668);
xor U2281 (N_2281,N_1568,N_1682);
nor U2282 (N_2282,N_1835,N_1584);
or U2283 (N_2283,N_1873,N_1942);
or U2284 (N_2284,N_1579,N_1948);
nand U2285 (N_2285,N_1671,N_1568);
and U2286 (N_2286,N_1736,N_1664);
xor U2287 (N_2287,N_1866,N_1973);
and U2288 (N_2288,N_1597,N_1923);
or U2289 (N_2289,N_1830,N_1837);
nand U2290 (N_2290,N_1585,N_1842);
nand U2291 (N_2291,N_1737,N_1736);
and U2292 (N_2292,N_1723,N_1728);
or U2293 (N_2293,N_1712,N_1593);
and U2294 (N_2294,N_1906,N_1846);
nand U2295 (N_2295,N_1708,N_1802);
and U2296 (N_2296,N_1990,N_1861);
and U2297 (N_2297,N_1577,N_1836);
or U2298 (N_2298,N_1996,N_1771);
nand U2299 (N_2299,N_1591,N_1948);
nand U2300 (N_2300,N_1904,N_1751);
xor U2301 (N_2301,N_1923,N_1993);
or U2302 (N_2302,N_1805,N_1959);
or U2303 (N_2303,N_1505,N_1710);
and U2304 (N_2304,N_1947,N_1974);
nand U2305 (N_2305,N_1626,N_1517);
nor U2306 (N_2306,N_1606,N_1793);
and U2307 (N_2307,N_1883,N_1908);
nor U2308 (N_2308,N_1949,N_1667);
and U2309 (N_2309,N_1828,N_1791);
nand U2310 (N_2310,N_1904,N_1731);
or U2311 (N_2311,N_1692,N_1539);
nor U2312 (N_2312,N_1782,N_1883);
nand U2313 (N_2313,N_1636,N_1535);
nor U2314 (N_2314,N_1513,N_1790);
and U2315 (N_2315,N_1948,N_1842);
and U2316 (N_2316,N_1970,N_1534);
nand U2317 (N_2317,N_1778,N_1528);
xnor U2318 (N_2318,N_1543,N_1652);
or U2319 (N_2319,N_1603,N_1745);
nor U2320 (N_2320,N_1828,N_1686);
and U2321 (N_2321,N_1524,N_1638);
xor U2322 (N_2322,N_1556,N_1509);
and U2323 (N_2323,N_1570,N_1766);
nor U2324 (N_2324,N_1532,N_1797);
nor U2325 (N_2325,N_1539,N_1652);
nand U2326 (N_2326,N_1901,N_1524);
nor U2327 (N_2327,N_1837,N_1587);
nand U2328 (N_2328,N_1769,N_1957);
nand U2329 (N_2329,N_1551,N_1820);
nor U2330 (N_2330,N_1676,N_1867);
or U2331 (N_2331,N_1768,N_1523);
and U2332 (N_2332,N_1789,N_1500);
and U2333 (N_2333,N_1507,N_1877);
nand U2334 (N_2334,N_1812,N_1510);
nor U2335 (N_2335,N_1765,N_1885);
nor U2336 (N_2336,N_1733,N_1648);
nor U2337 (N_2337,N_1870,N_1725);
nand U2338 (N_2338,N_1826,N_1505);
or U2339 (N_2339,N_1561,N_1513);
and U2340 (N_2340,N_1964,N_1745);
or U2341 (N_2341,N_1540,N_1757);
nor U2342 (N_2342,N_1695,N_1670);
and U2343 (N_2343,N_1616,N_1820);
xnor U2344 (N_2344,N_1776,N_1860);
and U2345 (N_2345,N_1923,N_1717);
nand U2346 (N_2346,N_1596,N_1635);
or U2347 (N_2347,N_1889,N_1599);
or U2348 (N_2348,N_1918,N_1523);
and U2349 (N_2349,N_1619,N_1665);
nor U2350 (N_2350,N_1678,N_1922);
nand U2351 (N_2351,N_1584,N_1843);
or U2352 (N_2352,N_1652,N_1844);
xnor U2353 (N_2353,N_1631,N_1804);
nor U2354 (N_2354,N_1501,N_1860);
or U2355 (N_2355,N_1740,N_1767);
and U2356 (N_2356,N_1842,N_1713);
nor U2357 (N_2357,N_1652,N_1723);
or U2358 (N_2358,N_1685,N_1932);
xnor U2359 (N_2359,N_1593,N_1625);
xnor U2360 (N_2360,N_1639,N_1603);
and U2361 (N_2361,N_1935,N_1659);
and U2362 (N_2362,N_1580,N_1685);
nand U2363 (N_2363,N_1567,N_1617);
nand U2364 (N_2364,N_1763,N_1858);
or U2365 (N_2365,N_1755,N_1634);
or U2366 (N_2366,N_1946,N_1809);
nand U2367 (N_2367,N_1717,N_1676);
nor U2368 (N_2368,N_1618,N_1898);
xor U2369 (N_2369,N_1998,N_1548);
and U2370 (N_2370,N_1700,N_1602);
and U2371 (N_2371,N_1594,N_1797);
nand U2372 (N_2372,N_1648,N_1663);
and U2373 (N_2373,N_1795,N_1523);
nor U2374 (N_2374,N_1827,N_1842);
or U2375 (N_2375,N_1805,N_1592);
nor U2376 (N_2376,N_1924,N_1558);
nand U2377 (N_2377,N_1759,N_1728);
and U2378 (N_2378,N_1550,N_1501);
xor U2379 (N_2379,N_1949,N_1562);
xnor U2380 (N_2380,N_1605,N_1891);
nor U2381 (N_2381,N_1509,N_1506);
and U2382 (N_2382,N_1736,N_1827);
and U2383 (N_2383,N_1520,N_1911);
or U2384 (N_2384,N_1587,N_1943);
nor U2385 (N_2385,N_1619,N_1528);
nor U2386 (N_2386,N_1705,N_1766);
or U2387 (N_2387,N_1536,N_1631);
nor U2388 (N_2388,N_1747,N_1746);
nor U2389 (N_2389,N_1512,N_1916);
nand U2390 (N_2390,N_1829,N_1656);
nand U2391 (N_2391,N_1674,N_1894);
and U2392 (N_2392,N_1982,N_1639);
and U2393 (N_2393,N_1729,N_1948);
and U2394 (N_2394,N_1946,N_1959);
xor U2395 (N_2395,N_1680,N_1972);
xor U2396 (N_2396,N_1749,N_1921);
and U2397 (N_2397,N_1541,N_1984);
or U2398 (N_2398,N_1903,N_1851);
or U2399 (N_2399,N_1884,N_1821);
and U2400 (N_2400,N_1779,N_1814);
nor U2401 (N_2401,N_1721,N_1641);
nor U2402 (N_2402,N_1908,N_1865);
nand U2403 (N_2403,N_1526,N_1624);
nand U2404 (N_2404,N_1763,N_1660);
nor U2405 (N_2405,N_1989,N_1965);
nor U2406 (N_2406,N_1738,N_1962);
and U2407 (N_2407,N_1895,N_1520);
and U2408 (N_2408,N_1901,N_1971);
nor U2409 (N_2409,N_1844,N_1766);
xnor U2410 (N_2410,N_1507,N_1967);
or U2411 (N_2411,N_1658,N_1554);
nand U2412 (N_2412,N_1731,N_1532);
nand U2413 (N_2413,N_1526,N_1713);
or U2414 (N_2414,N_1951,N_1673);
and U2415 (N_2415,N_1941,N_1784);
and U2416 (N_2416,N_1988,N_1856);
or U2417 (N_2417,N_1637,N_1817);
nand U2418 (N_2418,N_1939,N_1921);
nand U2419 (N_2419,N_1999,N_1716);
nand U2420 (N_2420,N_1627,N_1614);
or U2421 (N_2421,N_1725,N_1896);
nand U2422 (N_2422,N_1931,N_1655);
and U2423 (N_2423,N_1579,N_1673);
nor U2424 (N_2424,N_1854,N_1619);
nor U2425 (N_2425,N_1507,N_1851);
nand U2426 (N_2426,N_1607,N_1676);
and U2427 (N_2427,N_1909,N_1835);
nor U2428 (N_2428,N_1707,N_1695);
nor U2429 (N_2429,N_1795,N_1574);
or U2430 (N_2430,N_1820,N_1593);
or U2431 (N_2431,N_1747,N_1939);
and U2432 (N_2432,N_1831,N_1763);
nand U2433 (N_2433,N_1639,N_1946);
nor U2434 (N_2434,N_1810,N_1882);
nand U2435 (N_2435,N_1645,N_1580);
xnor U2436 (N_2436,N_1652,N_1685);
xnor U2437 (N_2437,N_1786,N_1742);
nand U2438 (N_2438,N_1860,N_1972);
nor U2439 (N_2439,N_1697,N_1814);
xor U2440 (N_2440,N_1823,N_1909);
nor U2441 (N_2441,N_1953,N_1746);
nand U2442 (N_2442,N_1874,N_1809);
nand U2443 (N_2443,N_1736,N_1527);
nor U2444 (N_2444,N_1737,N_1567);
or U2445 (N_2445,N_1538,N_1678);
and U2446 (N_2446,N_1996,N_1824);
or U2447 (N_2447,N_1773,N_1690);
or U2448 (N_2448,N_1891,N_1663);
and U2449 (N_2449,N_1796,N_1531);
xor U2450 (N_2450,N_1700,N_1956);
nor U2451 (N_2451,N_1948,N_1568);
and U2452 (N_2452,N_1670,N_1919);
nor U2453 (N_2453,N_1572,N_1829);
or U2454 (N_2454,N_1740,N_1689);
and U2455 (N_2455,N_1756,N_1843);
or U2456 (N_2456,N_1968,N_1970);
xnor U2457 (N_2457,N_1634,N_1838);
nand U2458 (N_2458,N_1702,N_1882);
nor U2459 (N_2459,N_1943,N_1754);
and U2460 (N_2460,N_1835,N_1665);
nor U2461 (N_2461,N_1752,N_1979);
xnor U2462 (N_2462,N_1726,N_1980);
nand U2463 (N_2463,N_1637,N_1808);
xor U2464 (N_2464,N_1781,N_1989);
and U2465 (N_2465,N_1964,N_1566);
nor U2466 (N_2466,N_1655,N_1530);
or U2467 (N_2467,N_1861,N_1598);
or U2468 (N_2468,N_1855,N_1870);
nor U2469 (N_2469,N_1748,N_1917);
nor U2470 (N_2470,N_1769,N_1624);
and U2471 (N_2471,N_1738,N_1830);
nand U2472 (N_2472,N_1866,N_1806);
nand U2473 (N_2473,N_1965,N_1888);
and U2474 (N_2474,N_1902,N_1749);
and U2475 (N_2475,N_1869,N_1573);
and U2476 (N_2476,N_1741,N_1524);
and U2477 (N_2477,N_1674,N_1541);
and U2478 (N_2478,N_1941,N_1580);
and U2479 (N_2479,N_1990,N_1915);
nand U2480 (N_2480,N_1726,N_1586);
and U2481 (N_2481,N_1605,N_1827);
or U2482 (N_2482,N_1937,N_1734);
or U2483 (N_2483,N_1854,N_1772);
and U2484 (N_2484,N_1822,N_1967);
nor U2485 (N_2485,N_1629,N_1597);
nor U2486 (N_2486,N_1531,N_1743);
xnor U2487 (N_2487,N_1649,N_1556);
nand U2488 (N_2488,N_1537,N_1873);
or U2489 (N_2489,N_1522,N_1643);
or U2490 (N_2490,N_1693,N_1590);
and U2491 (N_2491,N_1692,N_1782);
and U2492 (N_2492,N_1515,N_1660);
or U2493 (N_2493,N_1708,N_1761);
or U2494 (N_2494,N_1885,N_1833);
or U2495 (N_2495,N_1986,N_1732);
nor U2496 (N_2496,N_1744,N_1759);
and U2497 (N_2497,N_1860,N_1740);
or U2498 (N_2498,N_1512,N_1807);
and U2499 (N_2499,N_1566,N_1901);
nor U2500 (N_2500,N_2392,N_2015);
and U2501 (N_2501,N_2470,N_2151);
or U2502 (N_2502,N_2379,N_2361);
or U2503 (N_2503,N_2398,N_2100);
and U2504 (N_2504,N_2125,N_2449);
or U2505 (N_2505,N_2251,N_2194);
nand U2506 (N_2506,N_2074,N_2047);
nand U2507 (N_2507,N_2069,N_2090);
and U2508 (N_2508,N_2186,N_2054);
nand U2509 (N_2509,N_2331,N_2312);
or U2510 (N_2510,N_2055,N_2488);
nand U2511 (N_2511,N_2080,N_2436);
nor U2512 (N_2512,N_2463,N_2082);
xnor U2513 (N_2513,N_2044,N_2363);
or U2514 (N_2514,N_2152,N_2423);
nor U2515 (N_2515,N_2387,N_2328);
nand U2516 (N_2516,N_2264,N_2322);
and U2517 (N_2517,N_2109,N_2282);
and U2518 (N_2518,N_2123,N_2099);
and U2519 (N_2519,N_2349,N_2342);
and U2520 (N_2520,N_2014,N_2477);
nor U2521 (N_2521,N_2433,N_2106);
or U2522 (N_2522,N_2017,N_2405);
nand U2523 (N_2523,N_2475,N_2011);
nor U2524 (N_2524,N_2023,N_2027);
and U2525 (N_2525,N_2499,N_2163);
nor U2526 (N_2526,N_2112,N_2207);
and U2527 (N_2527,N_2494,N_2372);
nor U2528 (N_2528,N_2330,N_2235);
or U2529 (N_2529,N_2496,N_2242);
and U2530 (N_2530,N_2244,N_2323);
nor U2531 (N_2531,N_2297,N_2350);
and U2532 (N_2532,N_2348,N_2183);
nand U2533 (N_2533,N_2401,N_2130);
or U2534 (N_2534,N_2215,N_2386);
nand U2535 (N_2535,N_2158,N_2190);
or U2536 (N_2536,N_2059,N_2126);
and U2537 (N_2537,N_2335,N_2284);
or U2538 (N_2538,N_2421,N_2239);
nor U2539 (N_2539,N_2198,N_2346);
xor U2540 (N_2540,N_2155,N_2028);
and U2541 (N_2541,N_2443,N_2310);
xnor U2542 (N_2542,N_2424,N_2138);
and U2543 (N_2543,N_2365,N_2142);
nor U2544 (N_2544,N_2381,N_2431);
xnor U2545 (N_2545,N_2233,N_2077);
xor U2546 (N_2546,N_2049,N_2199);
nand U2547 (N_2547,N_2225,N_2202);
nor U2548 (N_2548,N_2139,N_2079);
or U2549 (N_2549,N_2291,N_2184);
nand U2550 (N_2550,N_2094,N_2232);
xnor U2551 (N_2551,N_2147,N_2238);
xnor U2552 (N_2552,N_2294,N_2218);
xnor U2553 (N_2553,N_2060,N_2088);
and U2554 (N_2554,N_2033,N_2408);
and U2555 (N_2555,N_2275,N_2181);
or U2556 (N_2556,N_2143,N_2241);
nor U2557 (N_2557,N_2168,N_2355);
xor U2558 (N_2558,N_2344,N_2473);
xor U2559 (N_2559,N_2256,N_2287);
nand U2560 (N_2560,N_2292,N_2117);
nand U2561 (N_2561,N_2351,N_2110);
nor U2562 (N_2562,N_2428,N_2131);
nand U2563 (N_2563,N_2179,N_2465);
nor U2564 (N_2564,N_2360,N_2356);
nor U2565 (N_2565,N_2396,N_2093);
and U2566 (N_2566,N_2434,N_2065);
nor U2567 (N_2567,N_2252,N_2309);
xnor U2568 (N_2568,N_2382,N_2249);
nand U2569 (N_2569,N_2277,N_2270);
nand U2570 (N_2570,N_2279,N_2299);
and U2571 (N_2571,N_2039,N_2013);
nand U2572 (N_2572,N_2283,N_2347);
and U2573 (N_2573,N_2036,N_2020);
nand U2574 (N_2574,N_2461,N_2324);
nand U2575 (N_2575,N_2224,N_2352);
and U2576 (N_2576,N_2373,N_2162);
nand U2577 (N_2577,N_2001,N_2257);
nand U2578 (N_2578,N_2076,N_2050);
or U2579 (N_2579,N_2305,N_2371);
or U2580 (N_2580,N_2263,N_2133);
and U2581 (N_2581,N_2266,N_2402);
nand U2582 (N_2582,N_2144,N_2478);
nand U2583 (N_2583,N_2010,N_2319);
xnor U2584 (N_2584,N_2317,N_2229);
and U2585 (N_2585,N_2145,N_2164);
and U2586 (N_2586,N_2046,N_2389);
nor U2587 (N_2587,N_2150,N_2493);
xor U2588 (N_2588,N_2458,N_2084);
nor U2589 (N_2589,N_2097,N_2000);
nor U2590 (N_2590,N_2228,N_2154);
nor U2591 (N_2591,N_2022,N_2078);
and U2592 (N_2592,N_2311,N_2453);
nor U2593 (N_2593,N_2073,N_2192);
xor U2594 (N_2594,N_2467,N_2129);
and U2595 (N_2595,N_2114,N_2037);
nor U2596 (N_2596,N_2188,N_2417);
and U2597 (N_2597,N_2214,N_2438);
or U2598 (N_2598,N_2153,N_2306);
xnor U2599 (N_2599,N_2092,N_2378);
nand U2600 (N_2600,N_2315,N_2081);
or U2601 (N_2601,N_2116,N_2107);
or U2602 (N_2602,N_2087,N_2182);
and U2603 (N_2603,N_2211,N_2432);
nor U2604 (N_2604,N_2327,N_2440);
nor U2605 (N_2605,N_2300,N_2083);
nand U2606 (N_2606,N_2469,N_2180);
nor U2607 (N_2607,N_2197,N_2255);
or U2608 (N_2608,N_2318,N_2062);
nand U2609 (N_2609,N_2149,N_2262);
or U2610 (N_2610,N_2212,N_2172);
and U2611 (N_2611,N_2018,N_2273);
nand U2612 (N_2612,N_2068,N_2380);
nor U2613 (N_2613,N_2095,N_2165);
nor U2614 (N_2614,N_2410,N_2167);
or U2615 (N_2615,N_2429,N_2240);
or U2616 (N_2616,N_2272,N_2450);
or U2617 (N_2617,N_2486,N_2177);
or U2618 (N_2618,N_2205,N_2267);
and U2619 (N_2619,N_2040,N_2425);
nor U2620 (N_2620,N_2329,N_2326);
nor U2621 (N_2621,N_2113,N_2254);
nor U2622 (N_2622,N_2189,N_2103);
nor U2623 (N_2623,N_2213,N_2217);
xnor U2624 (N_2624,N_2446,N_2383);
xnor U2625 (N_2625,N_2206,N_2456);
xnor U2626 (N_2626,N_2422,N_2419);
or U2627 (N_2627,N_2340,N_2220);
nor U2628 (N_2628,N_2271,N_2427);
nor U2629 (N_2629,N_2176,N_2245);
and U2630 (N_2630,N_2464,N_2159);
or U2631 (N_2631,N_2261,N_2048);
nand U2632 (N_2632,N_2089,N_2032);
and U2633 (N_2633,N_2343,N_2295);
and U2634 (N_2634,N_2231,N_2406);
or U2635 (N_2635,N_2485,N_2358);
nor U2636 (N_2636,N_2170,N_2368);
and U2637 (N_2637,N_2169,N_2135);
or U2638 (N_2638,N_2430,N_2070);
xnor U2639 (N_2639,N_2171,N_2320);
and U2640 (N_2640,N_2276,N_2411);
nand U2641 (N_2641,N_2246,N_2064);
or U2642 (N_2642,N_2426,N_2136);
nor U2643 (N_2643,N_2259,N_2490);
xor U2644 (N_2644,N_2399,N_2481);
or U2645 (N_2645,N_2203,N_2435);
and U2646 (N_2646,N_2376,N_2196);
xnor U2647 (N_2647,N_2004,N_2281);
or U2648 (N_2648,N_2035,N_2302);
and U2649 (N_2649,N_2075,N_2045);
nand U2650 (N_2650,N_2191,N_2071);
or U2651 (N_2651,N_2293,N_2003);
and U2652 (N_2652,N_2395,N_2210);
and U2653 (N_2653,N_2053,N_2104);
nor U2654 (N_2654,N_2471,N_2445);
nor U2655 (N_2655,N_2390,N_2012);
and U2656 (N_2656,N_2057,N_2115);
or U2657 (N_2657,N_2029,N_2394);
nor U2658 (N_2658,N_2332,N_2222);
nor U2659 (N_2659,N_2487,N_2400);
nor U2660 (N_2660,N_2479,N_2321);
nand U2661 (N_2661,N_2298,N_2121);
and U2662 (N_2662,N_2333,N_2007);
or U2663 (N_2663,N_2021,N_2460);
xnor U2664 (N_2664,N_2226,N_2454);
and U2665 (N_2665,N_2407,N_2026);
nand U2666 (N_2666,N_2141,N_2280);
nor U2667 (N_2667,N_2124,N_2412);
nor U2668 (N_2668,N_2457,N_2034);
and U2669 (N_2669,N_2223,N_2384);
or U2670 (N_2670,N_2375,N_2274);
nor U2671 (N_2671,N_2413,N_2146);
xnor U2672 (N_2672,N_2474,N_2128);
and U2673 (N_2673,N_2120,N_2303);
or U2674 (N_2674,N_2391,N_2268);
xor U2675 (N_2675,N_2316,N_2019);
and U2676 (N_2676,N_2489,N_2286);
nor U2677 (N_2677,N_2414,N_2385);
nand U2678 (N_2678,N_2448,N_2056);
and U2679 (N_2679,N_2404,N_2237);
nor U2680 (N_2680,N_2166,N_2006);
nand U2681 (N_2681,N_2250,N_2096);
or U2682 (N_2682,N_2403,N_2009);
nand U2683 (N_2683,N_2442,N_2416);
nor U2684 (N_2684,N_2236,N_2370);
nor U2685 (N_2685,N_2296,N_2483);
xnor U2686 (N_2686,N_2038,N_2174);
nand U2687 (N_2687,N_2441,N_2148);
nand U2688 (N_2688,N_2393,N_2193);
and U2689 (N_2689,N_2025,N_2132);
nor U2690 (N_2690,N_2043,N_2051);
nand U2691 (N_2691,N_2418,N_2337);
nor U2692 (N_2692,N_2314,N_2452);
nand U2693 (N_2693,N_2357,N_2498);
and U2694 (N_2694,N_2462,N_2313);
or U2695 (N_2695,N_2497,N_2216);
and U2696 (N_2696,N_2127,N_2157);
nand U2697 (N_2697,N_2415,N_2278);
and U2698 (N_2698,N_2098,N_2016);
nand U2699 (N_2699,N_2227,N_2451);
or U2700 (N_2700,N_2230,N_2052);
and U2701 (N_2701,N_2364,N_2173);
and U2702 (N_2702,N_2439,N_2409);
nand U2703 (N_2703,N_2369,N_2397);
nor U2704 (N_2704,N_2063,N_2156);
or U2705 (N_2705,N_2334,N_2253);
nor U2706 (N_2706,N_2243,N_2492);
nor U2707 (N_2707,N_2341,N_2288);
nor U2708 (N_2708,N_2388,N_2290);
and U2709 (N_2709,N_2265,N_2325);
nand U2710 (N_2710,N_2248,N_2377);
nand U2711 (N_2711,N_2195,N_2061);
nor U2712 (N_2712,N_2105,N_2108);
nor U2713 (N_2713,N_2459,N_2354);
nand U2714 (N_2714,N_2200,N_2476);
or U2715 (N_2715,N_2301,N_2111);
nand U2716 (N_2716,N_2058,N_2118);
or U2717 (N_2717,N_2482,N_2005);
nand U2718 (N_2718,N_2119,N_2366);
or U2719 (N_2719,N_2208,N_2221);
nand U2720 (N_2720,N_2234,N_2444);
xor U2721 (N_2721,N_2134,N_2187);
nand U2722 (N_2722,N_2359,N_2204);
nand U2723 (N_2723,N_2030,N_2367);
or U2724 (N_2724,N_2289,N_2160);
nor U2725 (N_2725,N_2178,N_2362);
nand U2726 (N_2726,N_2219,N_2002);
xor U2727 (N_2727,N_2338,N_2420);
nand U2728 (N_2728,N_2086,N_2067);
or U2729 (N_2729,N_2031,N_2345);
nand U2730 (N_2730,N_2480,N_2466);
or U2731 (N_2731,N_2455,N_2140);
nor U2732 (N_2732,N_2085,N_2353);
and U2733 (N_2733,N_2185,N_2258);
and U2734 (N_2734,N_2468,N_2209);
nor U2735 (N_2735,N_2102,N_2304);
nand U2736 (N_2736,N_2161,N_2122);
nand U2737 (N_2737,N_2201,N_2260);
nor U2738 (N_2738,N_2091,N_2472);
nor U2739 (N_2739,N_2336,N_2437);
or U2740 (N_2740,N_2491,N_2175);
and U2741 (N_2741,N_2247,N_2137);
and U2742 (N_2742,N_2042,N_2447);
and U2743 (N_2743,N_2041,N_2307);
xnor U2744 (N_2744,N_2101,N_2024);
or U2745 (N_2745,N_2374,N_2269);
nand U2746 (N_2746,N_2008,N_2484);
nor U2747 (N_2747,N_2072,N_2495);
nand U2748 (N_2748,N_2066,N_2339);
nor U2749 (N_2749,N_2308,N_2285);
nor U2750 (N_2750,N_2452,N_2027);
or U2751 (N_2751,N_2245,N_2483);
or U2752 (N_2752,N_2051,N_2282);
nand U2753 (N_2753,N_2345,N_2239);
and U2754 (N_2754,N_2047,N_2357);
xnor U2755 (N_2755,N_2298,N_2255);
nor U2756 (N_2756,N_2281,N_2270);
nand U2757 (N_2757,N_2444,N_2250);
and U2758 (N_2758,N_2241,N_2499);
or U2759 (N_2759,N_2366,N_2401);
nand U2760 (N_2760,N_2095,N_2421);
nor U2761 (N_2761,N_2145,N_2241);
nor U2762 (N_2762,N_2158,N_2221);
and U2763 (N_2763,N_2166,N_2100);
or U2764 (N_2764,N_2326,N_2211);
and U2765 (N_2765,N_2013,N_2426);
nor U2766 (N_2766,N_2166,N_2221);
nand U2767 (N_2767,N_2217,N_2189);
nand U2768 (N_2768,N_2094,N_2385);
or U2769 (N_2769,N_2212,N_2025);
nand U2770 (N_2770,N_2021,N_2400);
nor U2771 (N_2771,N_2034,N_2415);
nand U2772 (N_2772,N_2118,N_2205);
xor U2773 (N_2773,N_2459,N_2349);
and U2774 (N_2774,N_2167,N_2488);
nor U2775 (N_2775,N_2050,N_2166);
nand U2776 (N_2776,N_2411,N_2051);
nor U2777 (N_2777,N_2474,N_2388);
nor U2778 (N_2778,N_2417,N_2238);
or U2779 (N_2779,N_2079,N_2419);
nand U2780 (N_2780,N_2088,N_2176);
nand U2781 (N_2781,N_2049,N_2010);
nand U2782 (N_2782,N_2324,N_2276);
nand U2783 (N_2783,N_2416,N_2261);
or U2784 (N_2784,N_2158,N_2458);
nor U2785 (N_2785,N_2039,N_2299);
and U2786 (N_2786,N_2223,N_2121);
and U2787 (N_2787,N_2104,N_2095);
nor U2788 (N_2788,N_2297,N_2138);
nand U2789 (N_2789,N_2484,N_2363);
or U2790 (N_2790,N_2223,N_2338);
or U2791 (N_2791,N_2369,N_2074);
nand U2792 (N_2792,N_2133,N_2498);
nor U2793 (N_2793,N_2330,N_2025);
nor U2794 (N_2794,N_2103,N_2332);
xnor U2795 (N_2795,N_2169,N_2448);
nor U2796 (N_2796,N_2227,N_2045);
xnor U2797 (N_2797,N_2221,N_2440);
nor U2798 (N_2798,N_2446,N_2376);
and U2799 (N_2799,N_2016,N_2008);
xor U2800 (N_2800,N_2437,N_2451);
or U2801 (N_2801,N_2374,N_2011);
xnor U2802 (N_2802,N_2333,N_2364);
xor U2803 (N_2803,N_2482,N_2159);
nor U2804 (N_2804,N_2071,N_2422);
nand U2805 (N_2805,N_2033,N_2386);
nor U2806 (N_2806,N_2155,N_2241);
nand U2807 (N_2807,N_2248,N_2244);
nor U2808 (N_2808,N_2259,N_2014);
nor U2809 (N_2809,N_2358,N_2413);
nor U2810 (N_2810,N_2064,N_2313);
nor U2811 (N_2811,N_2182,N_2493);
nand U2812 (N_2812,N_2189,N_2183);
nor U2813 (N_2813,N_2419,N_2219);
nand U2814 (N_2814,N_2439,N_2444);
xor U2815 (N_2815,N_2456,N_2296);
nor U2816 (N_2816,N_2068,N_2155);
nand U2817 (N_2817,N_2142,N_2103);
nand U2818 (N_2818,N_2334,N_2285);
and U2819 (N_2819,N_2136,N_2498);
nand U2820 (N_2820,N_2444,N_2176);
or U2821 (N_2821,N_2430,N_2103);
nand U2822 (N_2822,N_2207,N_2470);
nor U2823 (N_2823,N_2433,N_2347);
nand U2824 (N_2824,N_2014,N_2288);
and U2825 (N_2825,N_2411,N_2421);
and U2826 (N_2826,N_2034,N_2237);
nand U2827 (N_2827,N_2022,N_2249);
nand U2828 (N_2828,N_2037,N_2439);
and U2829 (N_2829,N_2121,N_2449);
nor U2830 (N_2830,N_2211,N_2023);
and U2831 (N_2831,N_2478,N_2263);
and U2832 (N_2832,N_2096,N_2091);
or U2833 (N_2833,N_2111,N_2430);
nor U2834 (N_2834,N_2099,N_2027);
nor U2835 (N_2835,N_2102,N_2062);
nand U2836 (N_2836,N_2072,N_2158);
and U2837 (N_2837,N_2393,N_2058);
and U2838 (N_2838,N_2219,N_2377);
nor U2839 (N_2839,N_2146,N_2071);
and U2840 (N_2840,N_2016,N_2472);
nor U2841 (N_2841,N_2060,N_2048);
nor U2842 (N_2842,N_2413,N_2348);
nand U2843 (N_2843,N_2090,N_2370);
or U2844 (N_2844,N_2428,N_2254);
or U2845 (N_2845,N_2014,N_2388);
or U2846 (N_2846,N_2426,N_2134);
nand U2847 (N_2847,N_2241,N_2469);
and U2848 (N_2848,N_2287,N_2432);
and U2849 (N_2849,N_2040,N_2491);
or U2850 (N_2850,N_2071,N_2121);
xnor U2851 (N_2851,N_2361,N_2485);
nand U2852 (N_2852,N_2065,N_2017);
nor U2853 (N_2853,N_2023,N_2480);
nand U2854 (N_2854,N_2469,N_2053);
or U2855 (N_2855,N_2035,N_2018);
xnor U2856 (N_2856,N_2360,N_2011);
or U2857 (N_2857,N_2178,N_2034);
nand U2858 (N_2858,N_2429,N_2089);
xnor U2859 (N_2859,N_2184,N_2256);
nand U2860 (N_2860,N_2296,N_2195);
and U2861 (N_2861,N_2200,N_2048);
and U2862 (N_2862,N_2127,N_2017);
nor U2863 (N_2863,N_2030,N_2349);
and U2864 (N_2864,N_2451,N_2310);
or U2865 (N_2865,N_2249,N_2024);
or U2866 (N_2866,N_2194,N_2066);
and U2867 (N_2867,N_2012,N_2247);
nand U2868 (N_2868,N_2128,N_2149);
and U2869 (N_2869,N_2165,N_2197);
xnor U2870 (N_2870,N_2386,N_2126);
or U2871 (N_2871,N_2071,N_2091);
or U2872 (N_2872,N_2469,N_2439);
xor U2873 (N_2873,N_2289,N_2169);
nand U2874 (N_2874,N_2290,N_2410);
nand U2875 (N_2875,N_2497,N_2119);
and U2876 (N_2876,N_2025,N_2472);
xor U2877 (N_2877,N_2381,N_2498);
and U2878 (N_2878,N_2442,N_2198);
and U2879 (N_2879,N_2475,N_2122);
nand U2880 (N_2880,N_2479,N_2104);
or U2881 (N_2881,N_2171,N_2089);
or U2882 (N_2882,N_2023,N_2273);
nor U2883 (N_2883,N_2389,N_2255);
nor U2884 (N_2884,N_2190,N_2028);
nand U2885 (N_2885,N_2397,N_2043);
nand U2886 (N_2886,N_2375,N_2292);
nand U2887 (N_2887,N_2257,N_2313);
nor U2888 (N_2888,N_2214,N_2419);
nor U2889 (N_2889,N_2013,N_2300);
and U2890 (N_2890,N_2491,N_2207);
nand U2891 (N_2891,N_2331,N_2153);
or U2892 (N_2892,N_2265,N_2112);
and U2893 (N_2893,N_2329,N_2428);
nor U2894 (N_2894,N_2110,N_2410);
nor U2895 (N_2895,N_2053,N_2321);
nand U2896 (N_2896,N_2080,N_2176);
and U2897 (N_2897,N_2036,N_2174);
or U2898 (N_2898,N_2037,N_2002);
or U2899 (N_2899,N_2478,N_2058);
and U2900 (N_2900,N_2417,N_2233);
or U2901 (N_2901,N_2261,N_2203);
or U2902 (N_2902,N_2150,N_2138);
nor U2903 (N_2903,N_2179,N_2409);
and U2904 (N_2904,N_2496,N_2019);
nor U2905 (N_2905,N_2214,N_2300);
and U2906 (N_2906,N_2465,N_2051);
and U2907 (N_2907,N_2146,N_2354);
nand U2908 (N_2908,N_2006,N_2252);
and U2909 (N_2909,N_2440,N_2097);
nor U2910 (N_2910,N_2397,N_2252);
and U2911 (N_2911,N_2178,N_2148);
and U2912 (N_2912,N_2359,N_2450);
nor U2913 (N_2913,N_2173,N_2384);
nor U2914 (N_2914,N_2142,N_2322);
and U2915 (N_2915,N_2258,N_2365);
and U2916 (N_2916,N_2459,N_2192);
or U2917 (N_2917,N_2418,N_2037);
or U2918 (N_2918,N_2126,N_2160);
nor U2919 (N_2919,N_2126,N_2112);
and U2920 (N_2920,N_2283,N_2003);
or U2921 (N_2921,N_2048,N_2336);
xor U2922 (N_2922,N_2335,N_2008);
nand U2923 (N_2923,N_2157,N_2339);
and U2924 (N_2924,N_2160,N_2272);
or U2925 (N_2925,N_2204,N_2040);
nand U2926 (N_2926,N_2376,N_2344);
nand U2927 (N_2927,N_2038,N_2251);
and U2928 (N_2928,N_2068,N_2286);
or U2929 (N_2929,N_2080,N_2243);
and U2930 (N_2930,N_2441,N_2149);
and U2931 (N_2931,N_2271,N_2104);
and U2932 (N_2932,N_2052,N_2093);
or U2933 (N_2933,N_2498,N_2305);
xnor U2934 (N_2934,N_2290,N_2089);
nand U2935 (N_2935,N_2489,N_2325);
xnor U2936 (N_2936,N_2372,N_2227);
or U2937 (N_2937,N_2122,N_2137);
or U2938 (N_2938,N_2168,N_2003);
nor U2939 (N_2939,N_2435,N_2377);
nor U2940 (N_2940,N_2367,N_2331);
nor U2941 (N_2941,N_2170,N_2259);
or U2942 (N_2942,N_2414,N_2416);
or U2943 (N_2943,N_2379,N_2007);
and U2944 (N_2944,N_2127,N_2200);
nand U2945 (N_2945,N_2433,N_2361);
or U2946 (N_2946,N_2113,N_2013);
and U2947 (N_2947,N_2357,N_2260);
or U2948 (N_2948,N_2323,N_2426);
or U2949 (N_2949,N_2484,N_2097);
nand U2950 (N_2950,N_2427,N_2460);
and U2951 (N_2951,N_2484,N_2237);
and U2952 (N_2952,N_2075,N_2291);
nor U2953 (N_2953,N_2143,N_2077);
nand U2954 (N_2954,N_2480,N_2403);
or U2955 (N_2955,N_2040,N_2372);
and U2956 (N_2956,N_2303,N_2004);
nand U2957 (N_2957,N_2140,N_2009);
or U2958 (N_2958,N_2246,N_2009);
and U2959 (N_2959,N_2082,N_2088);
nand U2960 (N_2960,N_2083,N_2185);
or U2961 (N_2961,N_2081,N_2092);
nand U2962 (N_2962,N_2384,N_2098);
and U2963 (N_2963,N_2301,N_2377);
and U2964 (N_2964,N_2389,N_2069);
nor U2965 (N_2965,N_2122,N_2411);
or U2966 (N_2966,N_2142,N_2069);
and U2967 (N_2967,N_2423,N_2408);
and U2968 (N_2968,N_2404,N_2139);
nand U2969 (N_2969,N_2435,N_2354);
and U2970 (N_2970,N_2324,N_2293);
nand U2971 (N_2971,N_2408,N_2202);
and U2972 (N_2972,N_2346,N_2395);
nand U2973 (N_2973,N_2308,N_2003);
or U2974 (N_2974,N_2044,N_2181);
and U2975 (N_2975,N_2316,N_2484);
nor U2976 (N_2976,N_2097,N_2006);
nand U2977 (N_2977,N_2337,N_2194);
xor U2978 (N_2978,N_2055,N_2417);
nor U2979 (N_2979,N_2396,N_2331);
and U2980 (N_2980,N_2138,N_2203);
or U2981 (N_2981,N_2071,N_2055);
xor U2982 (N_2982,N_2247,N_2297);
nand U2983 (N_2983,N_2444,N_2287);
or U2984 (N_2984,N_2317,N_2493);
nor U2985 (N_2985,N_2423,N_2279);
xor U2986 (N_2986,N_2476,N_2160);
and U2987 (N_2987,N_2489,N_2288);
nand U2988 (N_2988,N_2302,N_2284);
and U2989 (N_2989,N_2034,N_2158);
xnor U2990 (N_2990,N_2099,N_2343);
xnor U2991 (N_2991,N_2467,N_2400);
and U2992 (N_2992,N_2333,N_2286);
and U2993 (N_2993,N_2216,N_2183);
xor U2994 (N_2994,N_2380,N_2125);
and U2995 (N_2995,N_2496,N_2060);
xnor U2996 (N_2996,N_2488,N_2475);
nor U2997 (N_2997,N_2201,N_2096);
nand U2998 (N_2998,N_2171,N_2333);
or U2999 (N_2999,N_2474,N_2215);
or UO_0 (O_0,N_2663,N_2584);
nor UO_1 (O_1,N_2648,N_2601);
nor UO_2 (O_2,N_2613,N_2804);
and UO_3 (O_3,N_2963,N_2808);
nor UO_4 (O_4,N_2664,N_2824);
or UO_5 (O_5,N_2796,N_2600);
nor UO_6 (O_6,N_2978,N_2854);
and UO_7 (O_7,N_2774,N_2834);
nor UO_8 (O_8,N_2517,N_2645);
or UO_9 (O_9,N_2863,N_2518);
xnor UO_10 (O_10,N_2729,N_2593);
nand UO_11 (O_11,N_2853,N_2913);
or UO_12 (O_12,N_2515,N_2948);
nor UO_13 (O_13,N_2975,N_2710);
nand UO_14 (O_14,N_2894,N_2655);
nand UO_15 (O_15,N_2903,N_2790);
or UO_16 (O_16,N_2884,N_2882);
nor UO_17 (O_17,N_2507,N_2723);
or UO_18 (O_18,N_2835,N_2526);
nor UO_19 (O_19,N_2772,N_2839);
nor UO_20 (O_20,N_2706,N_2512);
nand UO_21 (O_21,N_2879,N_2956);
nand UO_22 (O_22,N_2800,N_2656);
or UO_23 (O_23,N_2803,N_2533);
xnor UO_24 (O_24,N_2862,N_2757);
nand UO_25 (O_25,N_2717,N_2509);
and UO_26 (O_26,N_2747,N_2881);
xor UO_27 (O_27,N_2618,N_2597);
and UO_28 (O_28,N_2551,N_2749);
xnor UO_29 (O_29,N_2599,N_2638);
xnor UO_30 (O_30,N_2641,N_2845);
or UO_31 (O_31,N_2791,N_2691);
nor UO_32 (O_32,N_2654,N_2928);
and UO_33 (O_33,N_2525,N_2646);
nor UO_34 (O_34,N_2633,N_2625);
and UO_35 (O_35,N_2912,N_2728);
nor UO_36 (O_36,N_2787,N_2642);
nor UO_37 (O_37,N_2871,N_2883);
nor UO_38 (O_38,N_2754,N_2589);
or UO_39 (O_39,N_2877,N_2671);
or UO_40 (O_40,N_2698,N_2616);
xor UO_41 (O_41,N_2976,N_2983);
nand UO_42 (O_42,N_2636,N_2500);
nor UO_43 (O_43,N_2732,N_2842);
and UO_44 (O_44,N_2586,N_2895);
and UO_45 (O_45,N_2659,N_2611);
and UO_46 (O_46,N_2935,N_2994);
nor UO_47 (O_47,N_2847,N_2812);
nor UO_48 (O_48,N_2741,N_2738);
or UO_49 (O_49,N_2650,N_2521);
nand UO_50 (O_50,N_2987,N_2534);
nand UO_51 (O_51,N_2991,N_2936);
xnor UO_52 (O_52,N_2579,N_2857);
or UO_53 (O_53,N_2590,N_2891);
nor UO_54 (O_54,N_2662,N_2795);
xor UO_55 (O_55,N_2657,N_2964);
nand UO_56 (O_56,N_2554,N_2966);
or UO_57 (O_57,N_2680,N_2627);
or UO_58 (O_58,N_2773,N_2933);
nand UO_59 (O_59,N_2561,N_2524);
or UO_60 (O_60,N_2621,N_2694);
xnor UO_61 (O_61,N_2907,N_2575);
xor UO_62 (O_62,N_2667,N_2643);
xor UO_63 (O_63,N_2825,N_2875);
or UO_64 (O_64,N_2727,N_2878);
xnor UO_65 (O_65,N_2510,N_2814);
nand UO_66 (O_66,N_2789,N_2559);
nor UO_67 (O_67,N_2690,N_2753);
xnor UO_68 (O_68,N_2637,N_2563);
nor UO_69 (O_69,N_2969,N_2631);
and UO_70 (O_70,N_2892,N_2595);
nor UO_71 (O_71,N_2904,N_2763);
or UO_72 (O_72,N_2955,N_2736);
xor UO_73 (O_73,N_2911,N_2817);
and UO_74 (O_74,N_2940,N_2954);
and UO_75 (O_75,N_2609,N_2622);
and UO_76 (O_76,N_2992,N_2916);
or UO_77 (O_77,N_2914,N_2651);
and UO_78 (O_78,N_2675,N_2982);
xnor UO_79 (O_79,N_2957,N_2813);
nand UO_80 (O_80,N_2666,N_2527);
and UO_81 (O_81,N_2755,N_2899);
or UO_82 (O_82,N_2861,N_2921);
nor UO_83 (O_83,N_2931,N_2677);
and UO_84 (O_84,N_2565,N_2557);
or UO_85 (O_85,N_2793,N_2668);
nor UO_86 (O_86,N_2750,N_2560);
nor UO_87 (O_87,N_2759,N_2831);
or UO_88 (O_88,N_2827,N_2821);
and UO_89 (O_89,N_2567,N_2615);
nor UO_90 (O_90,N_2828,N_2799);
and UO_91 (O_91,N_2665,N_2902);
xor UO_92 (O_92,N_2923,N_2829);
nor UO_93 (O_93,N_2591,N_2910);
and UO_94 (O_94,N_2640,N_2783);
xnor UO_95 (O_95,N_2602,N_2697);
nand UO_96 (O_96,N_2746,N_2767);
and UO_97 (O_97,N_2573,N_2644);
nand UO_98 (O_98,N_2927,N_2777);
and UO_99 (O_99,N_2805,N_2617);
and UO_100 (O_100,N_2535,N_2999);
or UO_101 (O_101,N_2695,N_2528);
nor UO_102 (O_102,N_2979,N_2612);
and UO_103 (O_103,N_2959,N_2961);
and UO_104 (O_104,N_2583,N_2720);
nor UO_105 (O_105,N_2700,N_2544);
or UO_106 (O_106,N_2603,N_2626);
or UO_107 (O_107,N_2674,N_2730);
nor UO_108 (O_108,N_2532,N_2908);
nand UO_109 (O_109,N_2809,N_2873);
xor UO_110 (O_110,N_2553,N_2820);
nand UO_111 (O_111,N_2718,N_2807);
nor UO_112 (O_112,N_2592,N_2909);
or UO_113 (O_113,N_2762,N_2930);
and UO_114 (O_114,N_2962,N_2505);
or UO_115 (O_115,N_2685,N_2826);
or UO_116 (O_116,N_2836,N_2761);
and UO_117 (O_117,N_2968,N_2596);
nand UO_118 (O_118,N_2708,N_2922);
xnor UO_119 (O_119,N_2776,N_2890);
nand UO_120 (O_120,N_2770,N_2974);
xnor UO_121 (O_121,N_2538,N_2926);
nor UO_122 (O_122,N_2905,N_2840);
nand UO_123 (O_123,N_2558,N_2632);
or UO_124 (O_124,N_2806,N_2769);
or UO_125 (O_125,N_2744,N_2610);
or UO_126 (O_126,N_2540,N_2819);
or UO_127 (O_127,N_2766,N_2541);
and UO_128 (O_128,N_2856,N_2833);
or UO_129 (O_129,N_2511,N_2623);
and UO_130 (O_130,N_2798,N_2506);
and UO_131 (O_131,N_2570,N_2855);
xnor UO_132 (O_132,N_2702,N_2900);
or UO_133 (O_133,N_2849,N_2726);
or UO_134 (O_134,N_2764,N_2996);
xor UO_135 (O_135,N_2859,N_2858);
xor UO_136 (O_136,N_2660,N_2945);
and UO_137 (O_137,N_2925,N_2830);
nand UO_138 (O_138,N_2737,N_2519);
nor UO_139 (O_139,N_2571,N_2548);
and UO_140 (O_140,N_2993,N_2681);
nor UO_141 (O_141,N_2782,N_2693);
and UO_142 (O_142,N_2546,N_2688);
and UO_143 (O_143,N_2887,N_2876);
nor UO_144 (O_144,N_2545,N_2932);
or UO_145 (O_145,N_2823,N_2568);
nor UO_146 (O_146,N_2973,N_2536);
and UO_147 (O_147,N_2739,N_2815);
nand UO_148 (O_148,N_2598,N_2712);
nand UO_149 (O_149,N_2658,N_2550);
or UO_150 (O_150,N_2607,N_2582);
or UO_151 (O_151,N_2542,N_2822);
xnor UO_152 (O_152,N_2984,N_2786);
nand UO_153 (O_153,N_2722,N_2647);
or UO_154 (O_154,N_2713,N_2715);
nor UO_155 (O_155,N_2639,N_2846);
xor UO_156 (O_156,N_2941,N_2619);
and UO_157 (O_157,N_2503,N_2947);
nor UO_158 (O_158,N_2543,N_2952);
or UO_159 (O_159,N_2520,N_2797);
or UO_160 (O_160,N_2699,N_2965);
nand UO_161 (O_161,N_2868,N_2620);
nand UO_162 (O_162,N_2985,N_2679);
nand UO_163 (O_163,N_2889,N_2946);
nand UO_164 (O_164,N_2686,N_2724);
and UO_165 (O_165,N_2530,N_2844);
nand UO_166 (O_166,N_2634,N_2745);
or UO_167 (O_167,N_2917,N_2802);
or UO_168 (O_168,N_2816,N_2587);
or UO_169 (O_169,N_2841,N_2949);
nand UO_170 (O_170,N_2661,N_2604);
or UO_171 (O_171,N_2683,N_2578);
nand UO_172 (O_172,N_2980,N_2880);
nor UO_173 (O_173,N_2537,N_2733);
nor UO_174 (O_174,N_2672,N_2972);
and UO_175 (O_175,N_2635,N_2709);
xnor UO_176 (O_176,N_2758,N_2630);
or UO_177 (O_177,N_2838,N_2860);
or UO_178 (O_178,N_2864,N_2705);
nand UO_179 (O_179,N_2539,N_2760);
xnor UO_180 (O_180,N_2942,N_2811);
nand UO_181 (O_181,N_2522,N_2735);
nor UO_182 (O_182,N_2742,N_2549);
and UO_183 (O_183,N_2516,N_2788);
nor UO_184 (O_184,N_2896,N_2939);
or UO_185 (O_185,N_2832,N_2779);
or UO_186 (O_186,N_2934,N_2673);
nand UO_187 (O_187,N_2501,N_2986);
and UO_188 (O_188,N_2555,N_2508);
or UO_189 (O_189,N_2707,N_2676);
or UO_190 (O_190,N_2867,N_2970);
nor UO_191 (O_191,N_2608,N_2703);
nand UO_192 (O_192,N_2513,N_2566);
nand UO_193 (O_193,N_2901,N_2514);
nor UO_194 (O_194,N_2775,N_2924);
nor UO_195 (O_195,N_2851,N_2780);
nor UO_196 (O_196,N_2848,N_2624);
or UO_197 (O_197,N_2564,N_2725);
and UO_198 (O_198,N_2950,N_2938);
or UO_199 (O_199,N_2778,N_2898);
nor UO_200 (O_200,N_2751,N_2605);
and UO_201 (O_201,N_2971,N_2906);
xor UO_202 (O_202,N_2740,N_2678);
nand UO_203 (O_203,N_2687,N_2581);
nand UO_204 (O_204,N_2670,N_2574);
or UO_205 (O_205,N_2628,N_2653);
and UO_206 (O_206,N_2756,N_2711);
nand UO_207 (O_207,N_2997,N_2765);
nor UO_208 (O_208,N_2850,N_2734);
nor UO_209 (O_209,N_2748,N_2810);
nor UO_210 (O_210,N_2652,N_2870);
or UO_211 (O_211,N_2801,N_2523);
nand UO_212 (O_212,N_2569,N_2872);
or UO_213 (O_213,N_2953,N_2704);
nor UO_214 (O_214,N_2929,N_2629);
nand UO_215 (O_215,N_2869,N_2606);
and UO_216 (O_216,N_2714,N_2874);
nand UO_217 (O_217,N_2944,N_2684);
nor UO_218 (O_218,N_2731,N_2784);
nand UO_219 (O_219,N_2531,N_2843);
or UO_220 (O_220,N_2852,N_2614);
nand UO_221 (O_221,N_2866,N_2918);
and UO_222 (O_222,N_2943,N_2577);
nor UO_223 (O_223,N_2701,N_2818);
nand UO_224 (O_224,N_2794,N_2981);
nand UO_225 (O_225,N_2837,N_2716);
or UO_226 (O_226,N_2669,N_2502);
xnor UO_227 (O_227,N_2885,N_2990);
nor UO_228 (O_228,N_2781,N_2919);
and UO_229 (O_229,N_2504,N_2989);
nand UO_230 (O_230,N_2692,N_2958);
xnor UO_231 (O_231,N_2576,N_2547);
nor UO_232 (O_232,N_2556,N_2689);
xor UO_233 (O_233,N_2785,N_2580);
or UO_234 (O_234,N_2588,N_2995);
and UO_235 (O_235,N_2649,N_2886);
nand UO_236 (O_236,N_2937,N_2719);
nor UO_237 (O_237,N_2977,N_2960);
or UO_238 (O_238,N_2915,N_2743);
xnor UO_239 (O_239,N_2888,N_2529);
or UO_240 (O_240,N_2988,N_2682);
and UO_241 (O_241,N_2792,N_2897);
nand UO_242 (O_242,N_2893,N_2572);
or UO_243 (O_243,N_2771,N_2768);
nor UO_244 (O_244,N_2967,N_2865);
nor UO_245 (O_245,N_2920,N_2594);
nor UO_246 (O_246,N_2721,N_2998);
nand UO_247 (O_247,N_2562,N_2696);
nor UO_248 (O_248,N_2752,N_2552);
nand UO_249 (O_249,N_2951,N_2585);
xnor UO_250 (O_250,N_2634,N_2774);
or UO_251 (O_251,N_2841,N_2621);
and UO_252 (O_252,N_2731,N_2894);
or UO_253 (O_253,N_2523,N_2908);
and UO_254 (O_254,N_2900,N_2547);
or UO_255 (O_255,N_2967,N_2776);
nand UO_256 (O_256,N_2511,N_2899);
nor UO_257 (O_257,N_2551,N_2878);
and UO_258 (O_258,N_2907,N_2596);
nor UO_259 (O_259,N_2609,N_2598);
and UO_260 (O_260,N_2778,N_2673);
nor UO_261 (O_261,N_2674,N_2594);
and UO_262 (O_262,N_2668,N_2735);
or UO_263 (O_263,N_2632,N_2650);
nand UO_264 (O_264,N_2733,N_2631);
nand UO_265 (O_265,N_2691,N_2823);
nand UO_266 (O_266,N_2884,N_2649);
nor UO_267 (O_267,N_2571,N_2740);
nand UO_268 (O_268,N_2689,N_2937);
nor UO_269 (O_269,N_2588,N_2823);
nand UO_270 (O_270,N_2768,N_2737);
xnor UO_271 (O_271,N_2970,N_2866);
or UO_272 (O_272,N_2994,N_2650);
nand UO_273 (O_273,N_2788,N_2997);
nor UO_274 (O_274,N_2966,N_2553);
nand UO_275 (O_275,N_2583,N_2861);
nand UO_276 (O_276,N_2949,N_2953);
xnor UO_277 (O_277,N_2566,N_2595);
or UO_278 (O_278,N_2989,N_2651);
xnor UO_279 (O_279,N_2789,N_2758);
or UO_280 (O_280,N_2993,N_2958);
or UO_281 (O_281,N_2772,N_2505);
and UO_282 (O_282,N_2707,N_2928);
and UO_283 (O_283,N_2616,N_2677);
or UO_284 (O_284,N_2553,N_2755);
or UO_285 (O_285,N_2510,N_2980);
or UO_286 (O_286,N_2850,N_2780);
xnor UO_287 (O_287,N_2831,N_2811);
nor UO_288 (O_288,N_2816,N_2826);
xor UO_289 (O_289,N_2754,N_2966);
or UO_290 (O_290,N_2527,N_2655);
nand UO_291 (O_291,N_2960,N_2886);
and UO_292 (O_292,N_2979,N_2768);
and UO_293 (O_293,N_2733,N_2652);
nor UO_294 (O_294,N_2703,N_2682);
xnor UO_295 (O_295,N_2605,N_2805);
or UO_296 (O_296,N_2779,N_2534);
or UO_297 (O_297,N_2637,N_2968);
and UO_298 (O_298,N_2896,N_2763);
nor UO_299 (O_299,N_2884,N_2691);
and UO_300 (O_300,N_2962,N_2640);
or UO_301 (O_301,N_2583,N_2508);
or UO_302 (O_302,N_2597,N_2603);
nor UO_303 (O_303,N_2626,N_2996);
and UO_304 (O_304,N_2820,N_2613);
or UO_305 (O_305,N_2928,N_2805);
and UO_306 (O_306,N_2732,N_2795);
or UO_307 (O_307,N_2613,N_2867);
or UO_308 (O_308,N_2957,N_2699);
xor UO_309 (O_309,N_2583,N_2980);
and UO_310 (O_310,N_2674,N_2956);
and UO_311 (O_311,N_2816,N_2539);
or UO_312 (O_312,N_2921,N_2559);
and UO_313 (O_313,N_2731,N_2644);
or UO_314 (O_314,N_2528,N_2789);
and UO_315 (O_315,N_2801,N_2787);
xnor UO_316 (O_316,N_2750,N_2566);
and UO_317 (O_317,N_2740,N_2894);
or UO_318 (O_318,N_2954,N_2741);
nor UO_319 (O_319,N_2565,N_2527);
nor UO_320 (O_320,N_2944,N_2697);
nand UO_321 (O_321,N_2606,N_2694);
or UO_322 (O_322,N_2962,N_2932);
or UO_323 (O_323,N_2657,N_2768);
or UO_324 (O_324,N_2778,N_2787);
and UO_325 (O_325,N_2947,N_2684);
or UO_326 (O_326,N_2850,N_2810);
or UO_327 (O_327,N_2988,N_2719);
or UO_328 (O_328,N_2633,N_2505);
or UO_329 (O_329,N_2957,N_2763);
or UO_330 (O_330,N_2785,N_2962);
and UO_331 (O_331,N_2500,N_2789);
or UO_332 (O_332,N_2618,N_2742);
or UO_333 (O_333,N_2658,N_2614);
nor UO_334 (O_334,N_2893,N_2651);
nor UO_335 (O_335,N_2624,N_2662);
or UO_336 (O_336,N_2765,N_2926);
nand UO_337 (O_337,N_2772,N_2754);
xnor UO_338 (O_338,N_2862,N_2837);
nor UO_339 (O_339,N_2849,N_2644);
xnor UO_340 (O_340,N_2559,N_2643);
nor UO_341 (O_341,N_2509,N_2626);
and UO_342 (O_342,N_2512,N_2828);
or UO_343 (O_343,N_2676,N_2917);
xnor UO_344 (O_344,N_2862,N_2923);
nor UO_345 (O_345,N_2958,N_2833);
nor UO_346 (O_346,N_2824,N_2967);
nand UO_347 (O_347,N_2987,N_2925);
nand UO_348 (O_348,N_2756,N_2921);
and UO_349 (O_349,N_2574,N_2774);
and UO_350 (O_350,N_2884,N_2903);
nor UO_351 (O_351,N_2567,N_2882);
nand UO_352 (O_352,N_2995,N_2857);
nor UO_353 (O_353,N_2599,N_2869);
nor UO_354 (O_354,N_2744,N_2908);
nand UO_355 (O_355,N_2783,N_2560);
nor UO_356 (O_356,N_2887,N_2601);
nand UO_357 (O_357,N_2604,N_2707);
or UO_358 (O_358,N_2809,N_2985);
and UO_359 (O_359,N_2643,N_2700);
xnor UO_360 (O_360,N_2802,N_2894);
or UO_361 (O_361,N_2755,N_2819);
and UO_362 (O_362,N_2551,N_2632);
nor UO_363 (O_363,N_2797,N_2630);
xnor UO_364 (O_364,N_2727,N_2871);
nor UO_365 (O_365,N_2718,N_2965);
or UO_366 (O_366,N_2916,N_2761);
or UO_367 (O_367,N_2976,N_2767);
nor UO_368 (O_368,N_2798,N_2896);
xor UO_369 (O_369,N_2572,N_2800);
nor UO_370 (O_370,N_2534,N_2795);
or UO_371 (O_371,N_2947,N_2744);
or UO_372 (O_372,N_2851,N_2659);
xnor UO_373 (O_373,N_2506,N_2578);
and UO_374 (O_374,N_2580,N_2849);
nand UO_375 (O_375,N_2709,N_2834);
nand UO_376 (O_376,N_2983,N_2981);
nor UO_377 (O_377,N_2503,N_2596);
xnor UO_378 (O_378,N_2502,N_2980);
or UO_379 (O_379,N_2947,N_2896);
nand UO_380 (O_380,N_2768,N_2908);
nor UO_381 (O_381,N_2906,N_2635);
nor UO_382 (O_382,N_2953,N_2875);
nor UO_383 (O_383,N_2573,N_2589);
or UO_384 (O_384,N_2978,N_2998);
or UO_385 (O_385,N_2631,N_2598);
nor UO_386 (O_386,N_2803,N_2765);
and UO_387 (O_387,N_2890,N_2967);
nor UO_388 (O_388,N_2889,N_2973);
or UO_389 (O_389,N_2649,N_2552);
nor UO_390 (O_390,N_2936,N_2790);
nor UO_391 (O_391,N_2717,N_2753);
or UO_392 (O_392,N_2598,N_2851);
nand UO_393 (O_393,N_2602,N_2582);
xor UO_394 (O_394,N_2996,N_2619);
nor UO_395 (O_395,N_2634,N_2809);
xor UO_396 (O_396,N_2527,N_2680);
and UO_397 (O_397,N_2502,N_2857);
and UO_398 (O_398,N_2623,N_2515);
nor UO_399 (O_399,N_2580,N_2591);
nand UO_400 (O_400,N_2865,N_2521);
or UO_401 (O_401,N_2848,N_2797);
and UO_402 (O_402,N_2717,N_2570);
and UO_403 (O_403,N_2728,N_2840);
or UO_404 (O_404,N_2769,N_2878);
nand UO_405 (O_405,N_2928,N_2956);
or UO_406 (O_406,N_2747,N_2861);
and UO_407 (O_407,N_2505,N_2861);
and UO_408 (O_408,N_2518,N_2688);
nand UO_409 (O_409,N_2541,N_2746);
or UO_410 (O_410,N_2686,N_2963);
nor UO_411 (O_411,N_2810,N_2819);
nor UO_412 (O_412,N_2753,N_2824);
and UO_413 (O_413,N_2684,N_2830);
xnor UO_414 (O_414,N_2809,N_2820);
xnor UO_415 (O_415,N_2534,N_2639);
or UO_416 (O_416,N_2809,N_2548);
and UO_417 (O_417,N_2530,N_2809);
nor UO_418 (O_418,N_2502,N_2737);
or UO_419 (O_419,N_2892,N_2928);
or UO_420 (O_420,N_2887,N_2627);
nor UO_421 (O_421,N_2651,N_2755);
or UO_422 (O_422,N_2838,N_2544);
or UO_423 (O_423,N_2793,N_2840);
nor UO_424 (O_424,N_2537,N_2718);
or UO_425 (O_425,N_2793,N_2981);
nand UO_426 (O_426,N_2694,N_2699);
or UO_427 (O_427,N_2841,N_2825);
nand UO_428 (O_428,N_2738,N_2903);
nand UO_429 (O_429,N_2904,N_2602);
xnor UO_430 (O_430,N_2893,N_2584);
or UO_431 (O_431,N_2890,N_2802);
xnor UO_432 (O_432,N_2596,N_2836);
xor UO_433 (O_433,N_2816,N_2631);
nand UO_434 (O_434,N_2785,N_2700);
nor UO_435 (O_435,N_2966,N_2851);
and UO_436 (O_436,N_2744,N_2910);
xnor UO_437 (O_437,N_2637,N_2864);
nor UO_438 (O_438,N_2902,N_2519);
xnor UO_439 (O_439,N_2820,N_2865);
nand UO_440 (O_440,N_2552,N_2588);
nor UO_441 (O_441,N_2937,N_2955);
or UO_442 (O_442,N_2836,N_2732);
nor UO_443 (O_443,N_2955,N_2669);
or UO_444 (O_444,N_2779,N_2971);
nor UO_445 (O_445,N_2824,N_2843);
and UO_446 (O_446,N_2675,N_2741);
and UO_447 (O_447,N_2794,N_2977);
nand UO_448 (O_448,N_2592,N_2979);
nor UO_449 (O_449,N_2816,N_2524);
nor UO_450 (O_450,N_2640,N_2637);
nor UO_451 (O_451,N_2796,N_2602);
nand UO_452 (O_452,N_2703,N_2974);
or UO_453 (O_453,N_2595,N_2629);
and UO_454 (O_454,N_2735,N_2911);
nand UO_455 (O_455,N_2855,N_2586);
nand UO_456 (O_456,N_2697,N_2584);
and UO_457 (O_457,N_2649,N_2877);
or UO_458 (O_458,N_2785,N_2670);
nand UO_459 (O_459,N_2636,N_2716);
and UO_460 (O_460,N_2895,N_2797);
nor UO_461 (O_461,N_2955,N_2523);
nor UO_462 (O_462,N_2978,N_2674);
or UO_463 (O_463,N_2682,N_2810);
and UO_464 (O_464,N_2975,N_2717);
nor UO_465 (O_465,N_2979,N_2839);
nand UO_466 (O_466,N_2588,N_2907);
or UO_467 (O_467,N_2590,N_2950);
nand UO_468 (O_468,N_2756,N_2750);
nand UO_469 (O_469,N_2835,N_2855);
nor UO_470 (O_470,N_2831,N_2936);
or UO_471 (O_471,N_2733,N_2579);
or UO_472 (O_472,N_2502,N_2731);
nand UO_473 (O_473,N_2764,N_2648);
and UO_474 (O_474,N_2500,N_2681);
nor UO_475 (O_475,N_2580,N_2741);
nand UO_476 (O_476,N_2910,N_2543);
nand UO_477 (O_477,N_2834,N_2657);
nor UO_478 (O_478,N_2899,N_2986);
nor UO_479 (O_479,N_2903,N_2894);
and UO_480 (O_480,N_2851,N_2751);
nor UO_481 (O_481,N_2862,N_2626);
and UO_482 (O_482,N_2932,N_2956);
xor UO_483 (O_483,N_2637,N_2739);
nor UO_484 (O_484,N_2566,N_2653);
nand UO_485 (O_485,N_2750,N_2715);
nand UO_486 (O_486,N_2591,N_2872);
and UO_487 (O_487,N_2936,N_2992);
nand UO_488 (O_488,N_2929,N_2649);
and UO_489 (O_489,N_2631,N_2533);
nand UO_490 (O_490,N_2539,N_2619);
nor UO_491 (O_491,N_2675,N_2758);
nand UO_492 (O_492,N_2782,N_2981);
or UO_493 (O_493,N_2586,N_2700);
and UO_494 (O_494,N_2526,N_2753);
nor UO_495 (O_495,N_2882,N_2841);
nor UO_496 (O_496,N_2523,N_2696);
and UO_497 (O_497,N_2780,N_2713);
nand UO_498 (O_498,N_2674,N_2632);
nand UO_499 (O_499,N_2840,N_2651);
endmodule