module basic_1000_10000_1500_100_levels_5xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nor U0 (N_0,In_40,In_653);
or U1 (N_1,In_31,In_476);
nor U2 (N_2,In_844,In_981);
and U3 (N_3,In_353,In_718);
nor U4 (N_4,In_479,In_542);
and U5 (N_5,In_944,In_57);
xnor U6 (N_6,In_722,In_909);
and U7 (N_7,In_261,In_229);
or U8 (N_8,In_879,In_558);
nand U9 (N_9,In_764,In_552);
or U10 (N_10,In_478,In_395);
or U11 (N_11,In_267,In_543);
or U12 (N_12,In_915,In_382);
and U13 (N_13,In_784,In_239);
and U14 (N_14,In_309,In_54);
and U15 (N_15,In_562,In_390);
or U16 (N_16,In_929,In_398);
nand U17 (N_17,In_787,In_882);
xnor U18 (N_18,In_607,In_958);
nand U19 (N_19,In_186,In_775);
and U20 (N_20,In_172,In_689);
and U21 (N_21,In_702,In_743);
or U22 (N_22,In_978,In_564);
nor U23 (N_23,In_497,In_582);
or U24 (N_24,In_532,In_703);
nand U25 (N_25,In_394,In_484);
or U26 (N_26,In_374,In_594);
and U27 (N_27,In_603,In_131);
or U28 (N_28,In_328,In_366);
nor U29 (N_29,In_585,In_126);
nor U30 (N_30,In_156,In_461);
nor U31 (N_31,In_52,In_575);
nand U32 (N_32,In_723,In_280);
nor U33 (N_33,In_822,In_505);
nor U34 (N_34,In_886,In_572);
or U35 (N_35,In_616,In_530);
nand U36 (N_36,In_533,In_826);
nand U37 (N_37,In_165,In_742);
xnor U38 (N_38,In_363,In_690);
nor U39 (N_39,In_7,In_643);
nand U40 (N_40,In_860,In_574);
or U41 (N_41,In_486,In_214);
nor U42 (N_42,In_525,In_684);
and U43 (N_43,In_902,In_633);
nor U44 (N_44,In_244,In_134);
and U45 (N_45,In_122,In_794);
or U46 (N_46,In_231,In_135);
nor U47 (N_47,In_514,In_622);
or U48 (N_48,In_521,In_628);
or U49 (N_49,In_713,In_977);
nand U50 (N_50,In_597,In_284);
or U51 (N_51,In_389,In_454);
nand U52 (N_52,In_881,In_350);
nand U53 (N_53,In_602,In_460);
or U54 (N_54,In_618,In_788);
nand U55 (N_55,In_320,In_121);
and U56 (N_56,In_220,In_841);
xor U57 (N_57,In_265,In_474);
and U58 (N_58,In_636,In_254);
or U59 (N_59,In_931,In_963);
nor U60 (N_60,In_817,In_998);
nor U61 (N_61,In_277,In_235);
and U62 (N_62,In_59,In_71);
nand U63 (N_63,In_502,In_746);
or U64 (N_64,In_921,In_178);
and U65 (N_65,In_279,In_839);
and U66 (N_66,In_438,In_696);
nor U67 (N_67,In_419,In_922);
nor U68 (N_68,In_606,In_835);
nand U69 (N_69,In_615,In_767);
and U70 (N_70,In_880,In_369);
nor U71 (N_71,In_90,In_272);
or U72 (N_72,In_21,In_85);
nand U73 (N_73,In_544,In_301);
xnor U74 (N_74,In_691,In_845);
xor U75 (N_75,In_330,In_660);
nand U76 (N_76,In_424,In_276);
nor U77 (N_77,In_992,In_979);
xnor U78 (N_78,In_207,In_295);
xnor U79 (N_79,In_458,In_162);
or U80 (N_80,In_924,In_311);
and U81 (N_81,In_549,In_409);
nand U82 (N_82,In_682,In_766);
nor U83 (N_83,In_733,In_114);
nor U84 (N_84,In_506,In_967);
or U85 (N_85,In_571,In_34);
and U86 (N_86,In_440,In_570);
nor U87 (N_87,In_517,In_82);
xnor U88 (N_88,In_348,In_30);
xor U89 (N_89,In_119,In_983);
nand U90 (N_90,In_180,In_687);
and U91 (N_91,In_827,In_700);
or U92 (N_92,In_905,In_446);
and U93 (N_93,In_730,In_432);
nand U94 (N_94,In_972,In_230);
nand U95 (N_95,In_536,In_26);
nand U96 (N_96,In_298,In_355);
nor U97 (N_97,In_125,In_495);
or U98 (N_98,In_185,In_74);
xnor U99 (N_99,In_117,In_107);
and U100 (N_100,In_953,In_406);
or U101 (N_101,In_588,In_737);
nand U102 (N_102,N_12,N_75);
and U103 (N_103,N_96,In_305);
and U104 (N_104,In_782,In_601);
nor U105 (N_105,In_332,In_926);
nor U106 (N_106,In_200,In_205);
or U107 (N_107,In_216,In_412);
and U108 (N_108,N_88,In_55);
and U109 (N_109,In_0,In_193);
nor U110 (N_110,In_555,In_673);
and U111 (N_111,N_80,In_566);
nand U112 (N_112,N_25,In_580);
nand U113 (N_113,In_793,In_890);
xor U114 (N_114,In_403,In_397);
nor U115 (N_115,In_526,In_83);
nor U116 (N_116,In_170,In_413);
nor U117 (N_117,N_92,In_147);
nand U118 (N_118,In_138,In_211);
nand U119 (N_119,In_504,In_725);
nand U120 (N_120,In_511,In_393);
nor U121 (N_121,In_509,In_97);
nand U122 (N_122,In_176,In_747);
or U123 (N_123,In_686,In_133);
nor U124 (N_124,In_187,In_183);
nand U125 (N_125,In_213,In_2);
nor U126 (N_126,In_891,In_589);
nor U127 (N_127,In_892,In_73);
nand U128 (N_128,N_43,N_78);
and U129 (N_129,In_518,N_49);
and U130 (N_130,In_955,In_294);
or U131 (N_131,In_949,In_577);
nor U132 (N_132,In_810,In_415);
or U133 (N_133,In_593,In_539);
and U134 (N_134,In_334,In_318);
or U135 (N_135,In_857,N_73);
nor U136 (N_136,In_975,In_867);
nand U137 (N_137,In_245,N_62);
and U138 (N_138,In_217,In_657);
and U139 (N_139,In_993,In_798);
and U140 (N_140,In_4,In_257);
or U141 (N_141,In_136,In_275);
xnor U142 (N_142,In_300,In_443);
or U143 (N_143,In_58,In_223);
nand U144 (N_144,N_22,In_98);
and U145 (N_145,N_69,In_876);
or U146 (N_146,N_50,In_251);
or U147 (N_147,N_19,In_990);
xor U148 (N_148,In_286,In_473);
or U149 (N_149,In_523,In_654);
and U150 (N_150,N_38,In_510);
or U151 (N_151,In_584,In_417);
nand U152 (N_152,In_838,In_351);
nor U153 (N_153,N_23,N_59);
nor U154 (N_154,N_97,In_222);
and U155 (N_155,In_635,In_896);
and U156 (N_156,In_828,In_19);
nand U157 (N_157,In_120,In_604);
or U158 (N_158,In_695,In_319);
nand U159 (N_159,In_989,In_154);
nor U160 (N_160,N_93,In_883);
nand U161 (N_161,In_937,In_596);
nor U162 (N_162,In_538,N_45);
nor U163 (N_163,In_499,In_51);
and U164 (N_164,In_435,In_789);
or U165 (N_165,In_760,In_24);
and U166 (N_166,In_400,In_729);
or U167 (N_167,In_559,In_43);
or U168 (N_168,In_388,N_74);
or U169 (N_169,In_528,In_168);
and U170 (N_170,In_488,N_81);
nand U171 (N_171,In_966,In_242);
nand U172 (N_172,In_489,In_802);
nand U173 (N_173,In_316,In_236);
or U174 (N_174,In_155,In_60);
nor U175 (N_175,In_141,In_237);
nor U176 (N_176,In_195,In_666);
and U177 (N_177,In_675,In_67);
nand U178 (N_178,In_785,N_57);
or U179 (N_179,In_551,In_545);
or U180 (N_180,In_333,In_496);
nand U181 (N_181,In_386,In_144);
and U182 (N_182,In_865,In_641);
and U183 (N_183,In_541,In_270);
xor U184 (N_184,In_697,In_592);
or U185 (N_185,In_938,In_677);
nor U186 (N_186,In_91,In_201);
nand U187 (N_187,In_898,In_112);
nor U188 (N_188,In_964,In_611);
nor U189 (N_189,In_976,In_665);
or U190 (N_190,In_66,N_53);
and U191 (N_191,In_825,N_55);
or U192 (N_192,In_226,In_77);
or U193 (N_193,In_901,In_175);
xnor U194 (N_194,In_469,In_823);
nand U195 (N_195,In_44,In_961);
nand U196 (N_196,In_973,In_491);
or U197 (N_197,In_848,In_87);
nand U198 (N_198,In_342,In_765);
and U199 (N_199,In_221,In_158);
or U200 (N_200,In_317,N_135);
or U201 (N_201,In_965,In_262);
or U202 (N_202,In_281,N_70);
and U203 (N_203,In_368,In_816);
nor U204 (N_204,N_124,In_357);
and U205 (N_205,In_581,In_161);
and U206 (N_206,In_888,In_932);
nand U207 (N_207,In_53,In_293);
xnor U208 (N_208,N_60,In_380);
nor U209 (N_209,In_913,In_86);
or U210 (N_210,N_64,In_347);
nand U211 (N_211,In_290,In_630);
and U212 (N_212,N_155,In_727);
nor U213 (N_213,N_182,In_797);
xnor U214 (N_214,N_98,In_110);
xnor U215 (N_215,In_916,In_359);
or U216 (N_216,N_156,In_656);
and U217 (N_217,In_296,N_95);
nand U218 (N_218,In_847,N_101);
xor U219 (N_219,In_724,N_148);
or U220 (N_220,In_819,In_379);
nand U221 (N_221,In_741,In_774);
and U222 (N_222,In_269,In_352);
nor U223 (N_223,In_315,N_6);
and U224 (N_224,In_407,In_331);
nor U225 (N_225,In_149,In_649);
xor U226 (N_226,In_501,In_439);
nand U227 (N_227,In_971,In_402);
nor U228 (N_228,In_401,In_445);
and U229 (N_229,In_314,In_619);
xnor U230 (N_230,In_863,In_35);
nor U231 (N_231,In_621,N_159);
and U232 (N_232,In_232,In_451);
nor U233 (N_233,N_146,In_706);
nand U234 (N_234,N_67,In_763);
nor U235 (N_235,In_171,In_598);
nand U236 (N_236,In_970,In_820);
or U237 (N_237,In_959,N_189);
nor U238 (N_238,In_781,In_805);
or U239 (N_239,In_32,N_47);
nand U240 (N_240,In_659,In_988);
nand U241 (N_241,In_292,In_70);
and U242 (N_242,In_47,In_285);
and U243 (N_243,In_834,In_197);
nand U244 (N_244,In_508,In_934);
nor U245 (N_245,In_247,In_994);
nor U246 (N_246,In_493,In_768);
and U247 (N_247,In_645,In_814);
nand U248 (N_248,In_462,In_6);
or U249 (N_249,N_130,In_132);
nor U250 (N_250,In_431,In_153);
nand U251 (N_251,N_176,N_180);
and U252 (N_252,In_65,N_36);
nor U253 (N_253,In_408,In_92);
or U254 (N_254,N_161,N_10);
nand U255 (N_255,In_336,In_465);
nor U256 (N_256,In_591,In_312);
xor U257 (N_257,In_206,In_321);
and U258 (N_258,In_10,In_106);
xnor U259 (N_259,In_910,N_151);
or U260 (N_260,In_1,N_195);
and U261 (N_261,In_524,In_731);
nor U262 (N_262,In_701,N_100);
and U263 (N_263,In_914,In_456);
nand U264 (N_264,In_864,In_288);
xor U265 (N_265,In_227,In_668);
xor U266 (N_266,In_821,N_114);
nand U267 (N_267,In_780,In_837);
nand U268 (N_268,N_132,In_167);
nor U269 (N_269,In_776,In_253);
nand U270 (N_270,In_739,In_25);
or U271 (N_271,In_980,In_349);
nor U272 (N_272,N_193,In_629);
or U273 (N_273,N_108,In_411);
and U274 (N_274,In_507,N_13);
and U275 (N_275,In_343,In_557);
nor U276 (N_276,In_225,N_51);
or U277 (N_277,N_178,N_83);
nand U278 (N_278,In_118,N_16);
xor U279 (N_279,In_906,In_999);
or U280 (N_280,In_260,N_192);
nand U281 (N_281,N_18,In_189);
or U282 (N_282,In_907,In_772);
nor U283 (N_283,In_383,In_875);
nand U284 (N_284,N_9,In_670);
and U285 (N_285,In_579,N_82);
nand U286 (N_286,In_278,In_770);
and U287 (N_287,In_322,In_95);
and U288 (N_288,N_28,N_77);
xor U289 (N_289,N_42,N_186);
nor U290 (N_290,In_639,In_418);
and U291 (N_291,In_792,In_116);
nor U292 (N_292,In_655,N_72);
or U293 (N_293,N_136,In_410);
xnor U294 (N_294,In_783,N_165);
nor U295 (N_295,In_648,In_9);
nand U296 (N_296,N_133,In_215);
nor U297 (N_297,In_843,In_68);
xor U298 (N_298,N_160,N_103);
nand U299 (N_299,In_283,N_166);
nor U300 (N_300,In_799,N_140);
or U301 (N_301,N_169,N_39);
nand U302 (N_302,In_777,In_851);
or U303 (N_303,In_303,In_856);
xor U304 (N_304,In_11,N_234);
nand U305 (N_305,In_266,N_190);
nand U306 (N_306,In_519,In_853);
nor U307 (N_307,In_33,In_920);
and U308 (N_308,N_79,N_137);
nand U309 (N_309,N_52,N_84);
xor U310 (N_310,N_107,In_425);
nor U311 (N_311,In_234,N_58);
and U312 (N_312,In_69,In_813);
xor U313 (N_313,In_671,N_215);
nand U314 (N_314,N_54,In_5);
nand U315 (N_315,In_323,In_627);
or U316 (N_316,N_202,In_849);
or U317 (N_317,N_94,In_928);
xnor U318 (N_318,In_769,N_219);
or U319 (N_319,N_260,N_56);
nor U320 (N_320,N_90,In_459);
nor U321 (N_321,In_480,In_84);
or U322 (N_322,N_232,N_210);
nor U323 (N_323,In_846,In_75);
xor U324 (N_324,N_71,In_855);
nor U325 (N_325,In_81,In_996);
or U326 (N_326,In_634,In_302);
and U327 (N_327,In_483,N_194);
and U328 (N_328,In_145,In_680);
xor U329 (N_329,In_72,In_751);
or U330 (N_330,In_487,In_282);
and U331 (N_331,In_362,N_282);
or U332 (N_332,N_243,In_885);
nand U333 (N_333,N_157,N_24);
xor U334 (N_334,In_762,In_482);
nor U335 (N_335,N_200,N_209);
nor U336 (N_336,N_286,In_664);
and U337 (N_337,N_281,In_744);
or U338 (N_338,In_626,N_191);
nand U339 (N_339,In_800,In_356);
or U340 (N_340,In_109,N_113);
nand U341 (N_341,N_150,In_943);
or U342 (N_342,In_586,N_276);
and U343 (N_343,In_694,In_946);
and U344 (N_344,In_128,N_239);
or U345 (N_345,In_948,N_168);
nand U346 (N_346,In_99,In_877);
nor U347 (N_347,N_222,In_918);
nand U348 (N_348,N_206,In_831);
and U349 (N_349,In_537,In_866);
or U350 (N_350,N_162,In_516);
nor U351 (N_351,In_704,In_248);
and U352 (N_352,In_199,In_164);
and U353 (N_353,In_143,In_854);
nor U354 (N_354,In_307,In_39);
and U355 (N_355,In_354,In_950);
and U356 (N_356,In_177,In_893);
nor U357 (N_357,In_732,In_632);
nand U358 (N_358,In_255,In_416);
or U359 (N_359,In_693,In_27);
and U360 (N_360,In_803,In_712);
nor U361 (N_361,In_801,In_553);
nor U362 (N_362,In_194,In_674);
and U363 (N_363,In_908,In_139);
or U364 (N_364,N_227,N_241);
or U365 (N_365,In_137,In_360);
nand U366 (N_366,In_726,N_121);
xnor U367 (N_367,N_66,In_373);
nor U368 (N_368,In_754,In_858);
or U369 (N_369,In_995,In_748);
nor U370 (N_370,In_917,N_86);
nand U371 (N_371,In_399,N_289);
nand U372 (N_372,In_709,N_258);
and U373 (N_373,In_587,In_859);
or U374 (N_374,N_257,N_235);
nor U375 (N_375,N_35,In_683);
and U376 (N_376,In_576,In_16);
nor U377 (N_377,N_120,In_246);
nand U378 (N_378,In_287,N_207);
nor U379 (N_379,In_590,In_108);
nand U380 (N_380,In_273,In_749);
nand U381 (N_381,In_46,In_925);
nand U382 (N_382,In_830,In_494);
nor U383 (N_383,In_361,In_750);
xnor U384 (N_384,In_159,In_637);
and U385 (N_385,N_299,In_662);
and U386 (N_386,N_40,N_283);
nand U387 (N_387,In_61,N_170);
nand U388 (N_388,N_17,In_364);
nor U389 (N_389,N_218,In_644);
nand U390 (N_390,In_753,In_740);
or U391 (N_391,In_939,In_378);
nor U392 (N_392,In_985,In_196);
and U393 (N_393,N_290,In_919);
nor U394 (N_394,In_338,In_535);
and U395 (N_395,In_101,In_450);
nand U396 (N_396,In_927,In_738);
xnor U397 (N_397,N_30,N_261);
nand U398 (N_398,In_578,N_119);
or U399 (N_399,In_599,In_150);
or U400 (N_400,In_204,N_310);
nand U401 (N_401,In_113,In_640);
or U402 (N_402,N_138,In_678);
nor U403 (N_403,N_185,In_426);
and U404 (N_404,In_452,N_320);
nor U405 (N_405,In_911,N_347);
nand U406 (N_406,In_531,In_982);
and U407 (N_407,N_158,In_142);
nor U408 (N_408,In_808,In_468);
and U409 (N_409,N_181,In_475);
and U410 (N_410,N_167,N_153);
or U411 (N_411,N_389,In_62);
or U412 (N_412,In_872,N_212);
or U413 (N_413,In_889,In_850);
nor U414 (N_414,N_305,N_233);
xor U415 (N_415,In_48,N_267);
xnor U416 (N_416,N_164,In_466);
and U417 (N_417,N_127,In_852);
nand U418 (N_418,In_17,N_109);
and U419 (N_419,In_667,In_699);
nand U420 (N_420,N_251,N_3);
nand U421 (N_421,N_145,N_271);
nand U422 (N_422,N_339,In_540);
nor U423 (N_423,N_244,N_313);
and U424 (N_424,In_313,N_152);
or U425 (N_425,N_99,N_223);
and U426 (N_426,In_870,In_608);
xor U427 (N_427,In_812,In_447);
or U428 (N_428,In_271,In_49);
nor U429 (N_429,In_954,In_492);
nor U430 (N_430,In_151,N_317);
and U431 (N_431,N_360,In_651);
xnor U432 (N_432,N_297,In_923);
and U433 (N_433,N_341,In_795);
nor U434 (N_434,In_289,N_1);
nand U435 (N_435,In_376,N_106);
and U436 (N_436,In_182,N_291);
nand U437 (N_437,In_481,N_380);
nand U438 (N_438,N_346,N_225);
nand U439 (N_439,N_323,In_111);
or U440 (N_440,In_652,In_427);
and U441 (N_441,In_663,In_500);
nand U442 (N_442,In_734,In_42);
or U443 (N_443,In_771,N_328);
nand U444 (N_444,In_428,In_962);
and U445 (N_445,N_358,In_610);
or U446 (N_446,In_710,In_735);
nand U447 (N_447,In_94,N_8);
nand U448 (N_448,In_941,In_614);
nor U449 (N_449,N_300,In_984);
nor U450 (N_450,In_884,N_179);
or U451 (N_451,N_231,N_333);
xor U452 (N_452,In_811,N_221);
or U453 (N_453,In_952,In_513);
nor U454 (N_454,N_245,In_88);
and U455 (N_455,In_372,In_455);
nor U456 (N_456,N_87,N_230);
nand U457 (N_457,N_369,In_173);
xor U458 (N_458,In_676,N_349);
nand U459 (N_459,N_366,In_15);
and U460 (N_460,In_688,N_368);
and U461 (N_461,In_707,In_3);
or U462 (N_462,N_361,In_20);
and U463 (N_463,In_471,N_265);
nand U464 (N_464,N_263,In_202);
nand U465 (N_465,In_933,In_631);
nor U466 (N_466,In_498,N_353);
nor U467 (N_467,In_335,N_27);
nor U468 (N_468,In_711,N_104);
or U469 (N_469,In_124,N_177);
nor U470 (N_470,In_105,N_247);
nor U471 (N_471,N_115,In_22);
nor U472 (N_472,N_375,N_329);
or U473 (N_473,In_672,N_144);
xor U474 (N_474,In_396,In_661);
nand U475 (N_475,In_472,In_218);
nor U476 (N_476,In_371,In_986);
and U477 (N_477,N_278,In_609);
xnor U478 (N_478,In_512,In_642);
nand U479 (N_479,In_96,In_840);
and U480 (N_480,In_160,In_554);
nor U481 (N_481,In_829,In_241);
and U482 (N_482,In_951,In_940);
nor U483 (N_483,N_279,N_122);
nand U484 (N_484,In_370,N_270);
and U485 (N_485,N_4,In_930);
nor U486 (N_486,N_392,In_717);
nor U487 (N_487,In_679,In_377);
xnor U488 (N_488,In_947,N_105);
nand U489 (N_489,In_250,N_370);
nand U490 (N_490,In_887,N_201);
nor U491 (N_491,N_336,In_436);
nor U492 (N_492,N_48,In_759);
nand U493 (N_493,In_894,In_470);
nor U494 (N_494,N_292,In_624);
nor U495 (N_495,N_268,N_102);
xor U496 (N_496,In_8,In_969);
nor U497 (N_497,N_354,N_362);
or U498 (N_498,In_605,In_779);
and U499 (N_499,In_548,N_33);
or U500 (N_500,In_752,N_29);
nand U501 (N_501,N_401,In_174);
xor U502 (N_502,N_312,In_560);
xor U503 (N_503,N_430,N_183);
nor U504 (N_504,N_21,N_229);
or U505 (N_505,In_367,N_469);
xor U506 (N_506,N_126,In_715);
or U507 (N_507,N_345,N_112);
or U508 (N_508,N_302,In_720);
or U509 (N_509,In_297,In_324);
and U510 (N_510,N_129,N_388);
nor U511 (N_511,N_211,In_692);
nand U512 (N_512,N_26,In_14);
nand U513 (N_513,In_546,N_175);
and U514 (N_514,N_493,In_935);
nand U515 (N_515,In_429,In_756);
and U516 (N_516,In_600,N_421);
nor U517 (N_517,N_259,N_236);
nor U518 (N_518,N_378,In_184);
or U519 (N_519,In_129,In_453);
or U520 (N_520,In_568,N_449);
nor U521 (N_521,N_385,In_212);
nand U522 (N_522,In_904,In_874);
nand U523 (N_523,In_329,In_895);
and U524 (N_524,In_358,In_344);
nand U525 (N_525,N_32,In_130);
nand U526 (N_526,N_416,N_444);
nand U527 (N_527,In_146,N_249);
nand U528 (N_528,In_243,N_497);
or U529 (N_529,N_437,In_669);
nand U530 (N_530,N_141,In_249);
nand U531 (N_531,In_422,N_85);
nor U532 (N_532,N_63,N_208);
or U533 (N_533,N_205,In_224);
nor U534 (N_534,N_473,N_487);
nor U535 (N_535,N_197,In_623);
and U536 (N_536,N_496,N_316);
nor U537 (N_537,In_203,N_335);
and U538 (N_538,N_142,N_338);
and U539 (N_539,In_897,N_15);
or U540 (N_540,N_242,N_373);
nor U541 (N_541,N_255,N_428);
and U542 (N_542,N_226,In_547);
nand U543 (N_543,In_179,In_719);
nor U544 (N_544,In_268,In_942);
and U545 (N_545,In_522,N_455);
and U546 (N_546,N_116,In_341);
nor U547 (N_547,In_405,N_284);
or U548 (N_548,N_171,N_44);
nor U549 (N_549,N_31,N_438);
and U550 (N_550,N_163,N_348);
nand U551 (N_551,In_681,In_89);
nor U552 (N_552,N_149,N_376);
or U553 (N_553,N_415,N_383);
nor U554 (N_554,In_658,In_912);
nand U555 (N_555,N_371,In_12);
xor U556 (N_556,N_384,N_408);
and U557 (N_557,N_427,N_187);
nand U558 (N_558,N_327,In_104);
and U559 (N_559,N_466,N_293);
nand U560 (N_560,N_365,N_452);
or U561 (N_561,N_68,N_390);
and U562 (N_562,N_479,N_447);
nor U563 (N_563,N_425,In_38);
nand U564 (N_564,N_475,In_100);
or U565 (N_565,In_327,In_299);
nor U566 (N_566,In_263,N_311);
or U567 (N_567,N_342,In_716);
nor U568 (N_568,N_314,In_228);
nand U569 (N_569,In_325,N_448);
or U570 (N_570,In_467,N_198);
nor U571 (N_571,In_375,In_448);
nor U572 (N_572,N_275,In_638);
nand U573 (N_573,N_399,N_322);
nor U574 (N_574,In_583,N_91);
nor U575 (N_575,In_127,N_318);
xnor U576 (N_576,In_326,N_445);
or U577 (N_577,N_463,In_45);
or U578 (N_578,N_393,In_93);
nand U579 (N_579,N_435,N_266);
nand U580 (N_580,N_307,N_407);
nor U581 (N_581,N_443,N_472);
nor U582 (N_582,N_432,In_103);
nor U583 (N_583,In_903,N_214);
nor U584 (N_584,In_157,In_728);
or U585 (N_585,N_468,N_340);
or U586 (N_586,N_213,N_134);
or U587 (N_587,In_758,In_78);
nand U588 (N_588,In_337,N_471);
or U589 (N_589,In_842,N_14);
and U590 (N_590,N_173,N_417);
or U591 (N_591,N_488,N_220);
or U592 (N_592,N_306,N_499);
nor U593 (N_593,In_404,In_650);
or U594 (N_594,In_233,N_332);
or U595 (N_595,In_869,In_209);
and U596 (N_596,In_63,N_324);
nor U597 (N_597,N_89,N_461);
nand U598 (N_598,In_809,N_381);
nor U599 (N_599,N_216,In_818);
xor U600 (N_600,N_503,N_409);
or U601 (N_601,N_555,N_41);
nor U602 (N_602,N_295,N_539);
nor U603 (N_603,N_248,N_523);
nor U604 (N_604,N_379,In_13);
nor U605 (N_605,In_256,In_392);
and U606 (N_606,N_454,N_334);
and U607 (N_607,N_436,N_351);
or U608 (N_608,N_557,N_571);
nand U609 (N_609,N_174,N_565);
nor U610 (N_610,In_414,N_564);
xnor U611 (N_611,N_422,N_501);
nand U612 (N_612,In_804,In_833);
nand U613 (N_613,In_520,N_462);
xnor U614 (N_614,N_489,N_595);
or U615 (N_615,N_442,In_464);
and U616 (N_616,In_191,N_535);
nor U617 (N_617,N_543,N_131);
nor U618 (N_618,In_188,N_294);
xor U619 (N_619,In_346,N_397);
nand U620 (N_620,N_596,N_598);
and U621 (N_621,N_586,N_544);
or U622 (N_622,In_791,In_550);
or U623 (N_623,In_573,N_429);
and U624 (N_624,N_572,N_363);
nor U625 (N_625,N_538,In_595);
and U626 (N_626,N_567,N_413);
nor U627 (N_627,N_431,In_274);
nor U628 (N_628,N_382,N_128);
and U629 (N_629,N_285,N_514);
nand U630 (N_630,N_424,In_166);
nor U631 (N_631,N_391,N_46);
nand U632 (N_632,N_534,N_238);
nor U633 (N_633,N_518,N_524);
nand U634 (N_634,N_277,In_755);
nand U635 (N_635,In_23,N_542);
nand U636 (N_636,N_480,N_331);
nor U637 (N_637,N_528,N_326);
nor U638 (N_638,N_350,N_355);
or U639 (N_639,In_878,N_330);
and U640 (N_640,In_259,In_708);
and U641 (N_641,In_18,In_365);
nor U642 (N_642,N_592,N_520);
nor U643 (N_643,N_575,N_554);
xor U644 (N_644,In_806,In_968);
nand U645 (N_645,N_404,N_356);
and U646 (N_646,In_102,N_504);
or U647 (N_647,In_430,In_463);
nor U648 (N_648,N_117,N_395);
and U649 (N_649,N_545,In_36);
xnor U650 (N_650,N_439,In_871);
nor U651 (N_651,N_453,N_511);
nand U652 (N_652,In_721,N_485);
nor U653 (N_653,In_987,N_203);
or U654 (N_654,N_477,In_862);
or U655 (N_655,N_254,N_498);
xor U656 (N_656,In_625,N_588);
nand U657 (N_657,In_527,N_325);
or U658 (N_658,N_147,N_143);
or U659 (N_659,N_7,N_593);
and U660 (N_660,N_537,N_224);
nor U661 (N_661,In_423,In_900);
xnor U662 (N_662,N_541,In_477);
nand U663 (N_663,N_204,N_367);
nand U664 (N_664,N_552,N_502);
nand U665 (N_665,N_506,N_298);
nor U666 (N_666,In_80,In_442);
and U667 (N_667,N_184,N_563);
and U668 (N_668,In_64,In_181);
nor U669 (N_669,N_364,N_400);
and U670 (N_670,N_188,In_37);
and U671 (N_671,N_446,In_647);
or U672 (N_672,In_123,In_796);
and U673 (N_673,In_28,In_345);
or U674 (N_674,N_406,N_199);
nor U675 (N_675,N_478,In_381);
and U676 (N_676,In_387,In_252);
nor U677 (N_677,N_457,N_599);
or U678 (N_678,N_578,In_391);
nor U679 (N_679,In_773,N_526);
nor U680 (N_680,In_308,N_246);
or U681 (N_681,N_516,N_154);
and U682 (N_682,N_2,In_79);
nor U683 (N_683,In_873,N_490);
nand U684 (N_684,N_581,N_519);
nand U685 (N_685,In_441,N_540);
and U686 (N_686,In_503,N_296);
or U687 (N_687,N_303,In_957);
nand U688 (N_688,N_492,N_486);
nor U689 (N_689,N_460,N_508);
or U690 (N_690,N_589,N_11);
nor U691 (N_691,N_301,N_252);
or U692 (N_692,In_264,In_163);
nor U693 (N_693,In_304,In_807);
nand U694 (N_694,N_434,N_217);
and U695 (N_695,In_210,In_832);
and U696 (N_696,In_190,In_339);
and U697 (N_697,N_110,In_534);
and U698 (N_698,N_403,In_790);
or U699 (N_699,N_548,N_560);
or U700 (N_700,In_41,N_631);
nor U701 (N_701,N_604,N_450);
and U702 (N_702,N_309,In_529);
nand U703 (N_703,N_343,N_549);
and U704 (N_704,N_686,N_250);
nand U705 (N_705,N_522,N_580);
nor U706 (N_706,In_778,N_617);
and U707 (N_707,N_546,N_482);
or U708 (N_708,In_490,In_714);
or U709 (N_709,N_605,N_653);
xor U710 (N_710,N_695,N_663);
or U711 (N_711,N_517,In_421);
nor U712 (N_712,N_670,N_619);
nor U713 (N_713,N_440,N_111);
nand U714 (N_714,N_319,N_411);
or U715 (N_715,In_310,N_402);
and U716 (N_716,N_612,N_256);
nand U717 (N_717,N_691,N_673);
and U718 (N_718,N_590,N_602);
nor U719 (N_719,N_240,N_562);
or U720 (N_720,N_262,In_515);
and U721 (N_721,N_682,N_584);
nand U722 (N_722,In_449,N_669);
nand U723 (N_723,N_414,In_786);
nor U724 (N_724,N_608,N_253);
xor U725 (N_725,N_606,N_272);
xor U726 (N_726,In_698,N_579);
nor U727 (N_727,N_610,In_219);
nand U728 (N_728,N_597,N_139);
nor U729 (N_729,N_577,N_681);
nand U730 (N_730,N_576,N_643);
and U731 (N_731,N_683,N_566);
and U732 (N_732,In_736,N_685);
nor U733 (N_733,N_237,N_618);
and U734 (N_734,N_172,N_65);
or U735 (N_735,N_573,N_529);
nand U736 (N_736,N_591,N_650);
and U737 (N_737,N_649,N_396);
or U738 (N_738,N_627,N_521);
xor U739 (N_739,N_646,N_558);
nand U740 (N_740,In_685,N_377);
or U741 (N_741,N_196,N_568);
and U742 (N_742,N_507,N_405);
xor U743 (N_743,N_359,In_620);
nor U744 (N_744,N_500,N_659);
or U745 (N_745,In_258,N_637);
and U746 (N_746,In_563,N_505);
nand U747 (N_747,N_441,N_654);
or U748 (N_748,N_601,In_238);
and U749 (N_749,N_690,N_536);
and U750 (N_750,N_76,In_974);
or U751 (N_751,N_456,N_613);
nand U752 (N_752,N_5,N_315);
xnor U753 (N_753,In_434,In_433);
or U754 (N_754,N_684,N_594);
and U755 (N_755,N_614,In_291);
nor U756 (N_756,N_672,N_509);
nor U757 (N_757,N_352,N_668);
and U758 (N_758,N_625,In_485);
nand U759 (N_759,In_861,In_936);
nor U760 (N_760,N_616,N_675);
nand U761 (N_761,N_556,N_386);
or U762 (N_762,N_624,N_274);
nand U763 (N_763,N_433,N_623);
or U764 (N_764,In_815,N_470);
nand U765 (N_765,In_569,N_658);
or U766 (N_766,N_666,N_525);
or U767 (N_767,N_530,In_757);
or U768 (N_768,N_694,In_306);
xor U769 (N_769,N_228,N_337);
and U770 (N_770,N_287,In_617);
or U771 (N_771,N_633,N_288);
and U772 (N_772,In_991,N_280);
nor U773 (N_773,N_664,In_457);
xnor U774 (N_774,In_824,N_394);
or U775 (N_775,N_665,In_956);
nand U776 (N_776,N_645,N_420);
or U777 (N_777,N_344,N_264);
nand U778 (N_778,In_437,N_321);
and U779 (N_779,In_945,N_603);
or U780 (N_780,N_551,N_34);
or U781 (N_781,N_512,N_620);
nor U782 (N_782,N_611,N_638);
or U783 (N_783,In_612,N_626);
and U784 (N_784,N_398,N_372);
nor U785 (N_785,N_467,N_465);
nor U786 (N_786,N_678,N_634);
or U787 (N_787,N_585,N_533);
and U788 (N_788,N_412,N_688);
or U789 (N_789,In_148,N_547);
nor U790 (N_790,N_458,N_644);
xor U791 (N_791,N_642,N_125);
nand U792 (N_792,N_510,N_513);
and U793 (N_793,N_600,In_420);
nor U794 (N_794,In_556,N_615);
and U795 (N_795,N_474,In_152);
or U796 (N_796,N_459,N_582);
or U797 (N_797,N_689,In_646);
or U798 (N_798,N_495,N_677);
xor U799 (N_799,N_476,N_531);
and U800 (N_800,N_676,N_744);
or U801 (N_801,N_778,N_712);
or U802 (N_802,N_721,N_628);
and U803 (N_803,N_709,N_652);
or U804 (N_804,In_761,N_789);
xnor U805 (N_805,N_410,N_733);
or U806 (N_806,N_769,N_491);
nor U807 (N_807,In_192,N_630);
nor U808 (N_808,N_703,N_797);
nand U809 (N_809,N_737,N_374);
and U810 (N_810,N_799,N_749);
nand U811 (N_811,N_622,N_738);
or U812 (N_812,N_308,N_648);
nand U813 (N_813,N_569,In_29);
or U814 (N_814,N_640,N_426);
nand U815 (N_815,N_718,N_61);
and U816 (N_816,N_731,N_776);
or U817 (N_817,N_719,N_704);
nor U818 (N_818,N_722,N_742);
or U819 (N_819,N_760,N_387);
xnor U820 (N_820,N_609,N_680);
or U821 (N_821,N_780,N_657);
nor U822 (N_822,N_790,N_553);
and U823 (N_823,N_788,N_118);
or U824 (N_824,N_736,N_783);
xnor U825 (N_825,N_481,N_768);
and U826 (N_826,N_754,In_115);
or U827 (N_827,N_418,N_660);
and U828 (N_828,N_782,N_745);
or U829 (N_829,In_899,N_759);
nor U830 (N_830,N_357,N_671);
nor U831 (N_831,N_792,N_269);
nor U832 (N_832,N_734,N_750);
or U833 (N_833,N_661,N_707);
nor U834 (N_834,N_798,N_693);
and U835 (N_835,N_647,N_674);
and U836 (N_836,N_777,N_717);
and U837 (N_837,N_729,In_567);
and U838 (N_838,In_745,N_451);
nand U839 (N_839,N_767,In_240);
or U840 (N_840,N_755,N_710);
nor U841 (N_841,N_727,N_550);
and U842 (N_842,N_762,N_743);
and U843 (N_843,N_705,N_785);
and U844 (N_844,N_656,N_20);
or U845 (N_845,N_720,N_696);
xnor U846 (N_846,N_781,N_651);
nor U847 (N_847,N_796,N_667);
or U848 (N_848,N_583,N_735);
nor U849 (N_849,N_728,In_385);
or U850 (N_850,In_76,N_715);
nor U851 (N_851,N_779,N_723);
nand U852 (N_852,N_773,N_570);
xnor U853 (N_853,N_787,N_770);
nor U854 (N_854,N_716,In_565);
nor U855 (N_855,N_700,N_639);
nand U856 (N_856,N_698,N_795);
nor U857 (N_857,In_705,N_532);
nand U858 (N_858,In_50,N_632);
or U859 (N_859,N_304,In_960);
nand U860 (N_860,N_679,N_123);
and U861 (N_861,N_711,N_756);
nor U862 (N_862,N_771,N_774);
nor U863 (N_863,N_741,N_494);
nand U864 (N_864,N_687,N_746);
and U865 (N_865,N_764,In_198);
or U866 (N_866,In_997,In_613);
nor U867 (N_867,In_561,N_641);
nand U868 (N_868,N_635,In_169);
nor U869 (N_869,In_444,N_702);
and U870 (N_870,N_713,N_464);
nand U871 (N_871,In_140,N_793);
or U872 (N_872,N_636,N_739);
nor U873 (N_873,N_706,In_56);
and U874 (N_874,N_662,N_607);
nand U875 (N_875,N_730,N_587);
and U876 (N_876,N_629,N_527);
or U877 (N_877,N_725,In_384);
or U878 (N_878,N_559,N_794);
nor U879 (N_879,N_515,N_740);
xnor U880 (N_880,N_0,N_726);
nor U881 (N_881,N_763,N_753);
nor U882 (N_882,In_208,N_701);
or U883 (N_883,N_273,N_775);
or U884 (N_884,N_766,N_574);
or U885 (N_885,N_758,N_655);
nor U886 (N_886,N_752,N_786);
nor U887 (N_887,N_37,N_484);
nand U888 (N_888,N_561,In_868);
and U889 (N_889,N_732,N_761);
nor U890 (N_890,N_747,In_836);
or U891 (N_891,In_340,N_708);
or U892 (N_892,N_483,N_751);
nand U893 (N_893,N_419,N_699);
and U894 (N_894,N_765,N_772);
and U895 (N_895,N_757,N_714);
xnor U896 (N_896,N_692,N_724);
nor U897 (N_897,N_697,N_423);
nand U898 (N_898,N_791,N_621);
and U899 (N_899,N_748,N_784);
nor U900 (N_900,N_888,N_883);
or U901 (N_901,N_848,N_830);
and U902 (N_902,N_871,N_864);
xor U903 (N_903,N_890,N_811);
and U904 (N_904,N_858,N_826);
xnor U905 (N_905,N_840,N_851);
or U906 (N_906,N_849,N_842);
or U907 (N_907,N_859,N_839);
and U908 (N_908,N_855,N_879);
nand U909 (N_909,N_832,N_887);
and U910 (N_910,N_816,N_850);
and U911 (N_911,N_813,N_868);
nor U912 (N_912,N_854,N_852);
and U913 (N_913,N_800,N_857);
nor U914 (N_914,N_812,N_892);
or U915 (N_915,N_877,N_893);
and U916 (N_916,N_807,N_894);
nor U917 (N_917,N_806,N_819);
and U918 (N_918,N_815,N_817);
xnor U919 (N_919,N_873,N_876);
nand U920 (N_920,N_820,N_886);
nand U921 (N_921,N_818,N_809);
or U922 (N_922,N_829,N_860);
nor U923 (N_923,N_880,N_865);
or U924 (N_924,N_824,N_833);
nand U925 (N_925,N_889,N_835);
xor U926 (N_926,N_821,N_856);
and U927 (N_927,N_828,N_884);
or U928 (N_928,N_899,N_836);
nor U929 (N_929,N_897,N_823);
or U930 (N_930,N_898,N_891);
or U931 (N_931,N_875,N_838);
nor U932 (N_932,N_814,N_853);
and U933 (N_933,N_827,N_885);
and U934 (N_934,N_805,N_810);
and U935 (N_935,N_882,N_870);
and U936 (N_936,N_841,N_834);
or U937 (N_937,N_895,N_869);
or U938 (N_938,N_874,N_822);
nor U939 (N_939,N_872,N_845);
nor U940 (N_940,N_802,N_825);
and U941 (N_941,N_837,N_831);
nor U942 (N_942,N_843,N_847);
or U943 (N_943,N_878,N_866);
and U944 (N_944,N_803,N_804);
xnor U945 (N_945,N_801,N_896);
and U946 (N_946,N_867,N_844);
and U947 (N_947,N_863,N_846);
nor U948 (N_948,N_862,N_861);
xnor U949 (N_949,N_881,N_808);
nor U950 (N_950,N_897,N_873);
nand U951 (N_951,N_817,N_847);
xnor U952 (N_952,N_852,N_822);
nand U953 (N_953,N_884,N_833);
and U954 (N_954,N_800,N_847);
or U955 (N_955,N_859,N_853);
nor U956 (N_956,N_811,N_894);
or U957 (N_957,N_872,N_884);
nor U958 (N_958,N_864,N_893);
and U959 (N_959,N_875,N_893);
or U960 (N_960,N_852,N_889);
nor U961 (N_961,N_803,N_881);
and U962 (N_962,N_809,N_832);
nand U963 (N_963,N_868,N_858);
nor U964 (N_964,N_807,N_821);
or U965 (N_965,N_806,N_800);
nand U966 (N_966,N_898,N_885);
or U967 (N_967,N_876,N_831);
and U968 (N_968,N_835,N_896);
xor U969 (N_969,N_867,N_814);
xor U970 (N_970,N_874,N_816);
nor U971 (N_971,N_815,N_847);
nor U972 (N_972,N_822,N_838);
nor U973 (N_973,N_852,N_801);
nor U974 (N_974,N_818,N_852);
nor U975 (N_975,N_802,N_835);
xor U976 (N_976,N_835,N_898);
or U977 (N_977,N_880,N_858);
or U978 (N_978,N_896,N_832);
and U979 (N_979,N_862,N_813);
nor U980 (N_980,N_884,N_895);
or U981 (N_981,N_875,N_880);
and U982 (N_982,N_823,N_864);
or U983 (N_983,N_850,N_844);
nor U984 (N_984,N_844,N_834);
or U985 (N_985,N_803,N_859);
and U986 (N_986,N_836,N_867);
nor U987 (N_987,N_834,N_837);
xor U988 (N_988,N_829,N_876);
and U989 (N_989,N_821,N_826);
or U990 (N_990,N_810,N_875);
and U991 (N_991,N_879,N_892);
nand U992 (N_992,N_829,N_804);
nand U993 (N_993,N_832,N_867);
nor U994 (N_994,N_844,N_863);
and U995 (N_995,N_892,N_804);
and U996 (N_996,N_869,N_802);
nand U997 (N_997,N_875,N_873);
nor U998 (N_998,N_824,N_860);
nor U999 (N_999,N_817,N_895);
or U1000 (N_1000,N_950,N_977);
nand U1001 (N_1001,N_997,N_987);
nor U1002 (N_1002,N_923,N_973);
xnor U1003 (N_1003,N_995,N_904);
xnor U1004 (N_1004,N_934,N_932);
xnor U1005 (N_1005,N_986,N_985);
and U1006 (N_1006,N_928,N_979);
nor U1007 (N_1007,N_922,N_951);
xor U1008 (N_1008,N_967,N_981);
and U1009 (N_1009,N_918,N_917);
nor U1010 (N_1010,N_912,N_925);
or U1011 (N_1011,N_901,N_954);
nor U1012 (N_1012,N_938,N_921);
nor U1013 (N_1013,N_943,N_966);
nor U1014 (N_1014,N_957,N_914);
nand U1015 (N_1015,N_935,N_947);
nor U1016 (N_1016,N_910,N_926);
nand U1017 (N_1017,N_992,N_970);
or U1018 (N_1018,N_974,N_964);
and U1019 (N_1019,N_909,N_903);
nor U1020 (N_1020,N_937,N_993);
nor U1021 (N_1021,N_933,N_968);
nand U1022 (N_1022,N_902,N_905);
nor U1023 (N_1023,N_948,N_939);
nor U1024 (N_1024,N_972,N_924);
and U1025 (N_1025,N_942,N_998);
or U1026 (N_1026,N_991,N_959);
or U1027 (N_1027,N_965,N_988);
nand U1028 (N_1028,N_920,N_982);
and U1029 (N_1029,N_963,N_953);
nand U1030 (N_1030,N_944,N_927);
nand U1031 (N_1031,N_911,N_990);
or U1032 (N_1032,N_949,N_931);
or U1033 (N_1033,N_916,N_956);
and U1034 (N_1034,N_996,N_929);
nor U1035 (N_1035,N_978,N_936);
nor U1036 (N_1036,N_983,N_930);
and U1037 (N_1037,N_961,N_994);
nor U1038 (N_1038,N_946,N_969);
nand U1039 (N_1039,N_952,N_984);
or U1040 (N_1040,N_975,N_908);
or U1041 (N_1041,N_958,N_945);
and U1042 (N_1042,N_940,N_955);
and U1043 (N_1043,N_906,N_971);
or U1044 (N_1044,N_913,N_941);
and U1045 (N_1045,N_915,N_962);
and U1046 (N_1046,N_960,N_989);
and U1047 (N_1047,N_976,N_919);
nand U1048 (N_1048,N_900,N_907);
nor U1049 (N_1049,N_999,N_980);
or U1050 (N_1050,N_987,N_999);
or U1051 (N_1051,N_931,N_999);
xor U1052 (N_1052,N_984,N_963);
nand U1053 (N_1053,N_926,N_950);
nand U1054 (N_1054,N_968,N_915);
or U1055 (N_1055,N_921,N_945);
nand U1056 (N_1056,N_936,N_941);
or U1057 (N_1057,N_900,N_976);
nor U1058 (N_1058,N_984,N_992);
nor U1059 (N_1059,N_971,N_950);
nor U1060 (N_1060,N_940,N_972);
nor U1061 (N_1061,N_965,N_913);
or U1062 (N_1062,N_957,N_982);
and U1063 (N_1063,N_905,N_937);
or U1064 (N_1064,N_902,N_991);
and U1065 (N_1065,N_980,N_949);
nor U1066 (N_1066,N_969,N_912);
and U1067 (N_1067,N_981,N_957);
or U1068 (N_1068,N_970,N_943);
nand U1069 (N_1069,N_963,N_944);
xor U1070 (N_1070,N_958,N_998);
nor U1071 (N_1071,N_920,N_987);
and U1072 (N_1072,N_969,N_931);
nor U1073 (N_1073,N_929,N_960);
nor U1074 (N_1074,N_986,N_941);
nor U1075 (N_1075,N_907,N_937);
or U1076 (N_1076,N_941,N_990);
and U1077 (N_1077,N_900,N_918);
and U1078 (N_1078,N_967,N_954);
or U1079 (N_1079,N_926,N_979);
nand U1080 (N_1080,N_924,N_966);
nor U1081 (N_1081,N_925,N_981);
xnor U1082 (N_1082,N_967,N_958);
and U1083 (N_1083,N_968,N_999);
or U1084 (N_1084,N_924,N_977);
and U1085 (N_1085,N_987,N_953);
nand U1086 (N_1086,N_994,N_917);
nor U1087 (N_1087,N_953,N_941);
xor U1088 (N_1088,N_972,N_929);
or U1089 (N_1089,N_907,N_964);
nor U1090 (N_1090,N_955,N_989);
nand U1091 (N_1091,N_911,N_932);
and U1092 (N_1092,N_929,N_917);
or U1093 (N_1093,N_933,N_929);
and U1094 (N_1094,N_944,N_909);
or U1095 (N_1095,N_982,N_945);
nand U1096 (N_1096,N_907,N_920);
nand U1097 (N_1097,N_932,N_908);
and U1098 (N_1098,N_919,N_943);
or U1099 (N_1099,N_953,N_973);
or U1100 (N_1100,N_1093,N_1076);
nor U1101 (N_1101,N_1084,N_1077);
nand U1102 (N_1102,N_1079,N_1046);
or U1103 (N_1103,N_1021,N_1019);
nor U1104 (N_1104,N_1095,N_1036);
or U1105 (N_1105,N_1074,N_1059);
nor U1106 (N_1106,N_1049,N_1043);
nor U1107 (N_1107,N_1000,N_1035);
or U1108 (N_1108,N_1067,N_1055);
or U1109 (N_1109,N_1038,N_1053);
xor U1110 (N_1110,N_1014,N_1003);
nor U1111 (N_1111,N_1022,N_1032);
xnor U1112 (N_1112,N_1086,N_1018);
or U1113 (N_1113,N_1031,N_1065);
nand U1114 (N_1114,N_1033,N_1020);
nor U1115 (N_1115,N_1081,N_1091);
nand U1116 (N_1116,N_1060,N_1094);
nand U1117 (N_1117,N_1042,N_1088);
xnor U1118 (N_1118,N_1073,N_1083);
nand U1119 (N_1119,N_1099,N_1092);
xnor U1120 (N_1120,N_1039,N_1051);
and U1121 (N_1121,N_1029,N_1027);
or U1122 (N_1122,N_1013,N_1087);
xnor U1123 (N_1123,N_1098,N_1045);
nor U1124 (N_1124,N_1052,N_1089);
or U1125 (N_1125,N_1037,N_1006);
and U1126 (N_1126,N_1056,N_1072);
nor U1127 (N_1127,N_1030,N_1071);
or U1128 (N_1128,N_1061,N_1004);
nand U1129 (N_1129,N_1062,N_1008);
and U1130 (N_1130,N_1068,N_1025);
nor U1131 (N_1131,N_1001,N_1090);
nor U1132 (N_1132,N_1026,N_1002);
or U1133 (N_1133,N_1097,N_1075);
or U1134 (N_1134,N_1005,N_1078);
and U1135 (N_1135,N_1044,N_1017);
xnor U1136 (N_1136,N_1010,N_1028);
or U1137 (N_1137,N_1070,N_1040);
nand U1138 (N_1138,N_1058,N_1082);
or U1139 (N_1139,N_1063,N_1012);
nor U1140 (N_1140,N_1085,N_1057);
nand U1141 (N_1141,N_1048,N_1054);
and U1142 (N_1142,N_1023,N_1016);
nor U1143 (N_1143,N_1011,N_1096);
nand U1144 (N_1144,N_1047,N_1034);
nand U1145 (N_1145,N_1041,N_1007);
and U1146 (N_1146,N_1069,N_1024);
and U1147 (N_1147,N_1080,N_1064);
nor U1148 (N_1148,N_1066,N_1015);
nand U1149 (N_1149,N_1050,N_1009);
nand U1150 (N_1150,N_1016,N_1043);
nand U1151 (N_1151,N_1068,N_1062);
or U1152 (N_1152,N_1012,N_1073);
nand U1153 (N_1153,N_1079,N_1016);
and U1154 (N_1154,N_1086,N_1035);
nand U1155 (N_1155,N_1071,N_1061);
and U1156 (N_1156,N_1083,N_1028);
or U1157 (N_1157,N_1095,N_1087);
or U1158 (N_1158,N_1007,N_1072);
or U1159 (N_1159,N_1093,N_1054);
xor U1160 (N_1160,N_1060,N_1050);
nand U1161 (N_1161,N_1088,N_1081);
nand U1162 (N_1162,N_1066,N_1029);
nand U1163 (N_1163,N_1018,N_1095);
nor U1164 (N_1164,N_1092,N_1036);
and U1165 (N_1165,N_1080,N_1007);
or U1166 (N_1166,N_1047,N_1039);
and U1167 (N_1167,N_1010,N_1046);
nor U1168 (N_1168,N_1022,N_1064);
nand U1169 (N_1169,N_1095,N_1039);
and U1170 (N_1170,N_1053,N_1092);
nand U1171 (N_1171,N_1073,N_1060);
or U1172 (N_1172,N_1057,N_1090);
and U1173 (N_1173,N_1077,N_1015);
nor U1174 (N_1174,N_1090,N_1012);
nor U1175 (N_1175,N_1062,N_1040);
and U1176 (N_1176,N_1085,N_1063);
or U1177 (N_1177,N_1087,N_1003);
or U1178 (N_1178,N_1073,N_1067);
nand U1179 (N_1179,N_1087,N_1019);
or U1180 (N_1180,N_1079,N_1058);
nand U1181 (N_1181,N_1002,N_1004);
nor U1182 (N_1182,N_1094,N_1008);
xnor U1183 (N_1183,N_1034,N_1076);
nand U1184 (N_1184,N_1039,N_1006);
or U1185 (N_1185,N_1035,N_1040);
or U1186 (N_1186,N_1064,N_1094);
nand U1187 (N_1187,N_1076,N_1069);
or U1188 (N_1188,N_1095,N_1060);
or U1189 (N_1189,N_1063,N_1028);
nand U1190 (N_1190,N_1077,N_1082);
or U1191 (N_1191,N_1025,N_1003);
nor U1192 (N_1192,N_1077,N_1036);
xor U1193 (N_1193,N_1049,N_1072);
or U1194 (N_1194,N_1021,N_1008);
and U1195 (N_1195,N_1063,N_1026);
and U1196 (N_1196,N_1053,N_1073);
nand U1197 (N_1197,N_1083,N_1002);
or U1198 (N_1198,N_1037,N_1070);
nand U1199 (N_1199,N_1057,N_1036);
nand U1200 (N_1200,N_1192,N_1180);
or U1201 (N_1201,N_1118,N_1143);
or U1202 (N_1202,N_1105,N_1132);
or U1203 (N_1203,N_1179,N_1123);
nor U1204 (N_1204,N_1121,N_1160);
nor U1205 (N_1205,N_1133,N_1102);
nor U1206 (N_1206,N_1163,N_1187);
nand U1207 (N_1207,N_1131,N_1145);
or U1208 (N_1208,N_1106,N_1150);
nor U1209 (N_1209,N_1147,N_1198);
or U1210 (N_1210,N_1127,N_1188);
xor U1211 (N_1211,N_1164,N_1162);
nor U1212 (N_1212,N_1182,N_1167);
or U1213 (N_1213,N_1138,N_1175);
nor U1214 (N_1214,N_1185,N_1136);
and U1215 (N_1215,N_1169,N_1171);
xnor U1216 (N_1216,N_1156,N_1193);
or U1217 (N_1217,N_1154,N_1149);
nor U1218 (N_1218,N_1122,N_1197);
nor U1219 (N_1219,N_1166,N_1174);
and U1220 (N_1220,N_1117,N_1191);
nand U1221 (N_1221,N_1135,N_1129);
and U1222 (N_1222,N_1114,N_1140);
and U1223 (N_1223,N_1184,N_1157);
nor U1224 (N_1224,N_1161,N_1168);
or U1225 (N_1225,N_1176,N_1142);
and U1226 (N_1226,N_1177,N_1116);
nand U1227 (N_1227,N_1141,N_1120);
nor U1228 (N_1228,N_1119,N_1165);
and U1229 (N_1229,N_1152,N_1158);
or U1230 (N_1230,N_1109,N_1108);
nor U1231 (N_1231,N_1144,N_1112);
and U1232 (N_1232,N_1111,N_1130);
or U1233 (N_1233,N_1148,N_1125);
nor U1234 (N_1234,N_1137,N_1153);
nand U1235 (N_1235,N_1172,N_1101);
nor U1236 (N_1236,N_1194,N_1124);
nor U1237 (N_1237,N_1113,N_1170);
or U1238 (N_1238,N_1134,N_1183);
or U1239 (N_1239,N_1155,N_1199);
nor U1240 (N_1240,N_1100,N_1173);
or U1241 (N_1241,N_1103,N_1115);
or U1242 (N_1242,N_1196,N_1139);
nor U1243 (N_1243,N_1107,N_1190);
nand U1244 (N_1244,N_1146,N_1110);
and U1245 (N_1245,N_1178,N_1151);
nand U1246 (N_1246,N_1189,N_1159);
or U1247 (N_1247,N_1104,N_1195);
nand U1248 (N_1248,N_1126,N_1128);
or U1249 (N_1249,N_1181,N_1186);
nor U1250 (N_1250,N_1110,N_1190);
nor U1251 (N_1251,N_1150,N_1122);
nor U1252 (N_1252,N_1186,N_1157);
nand U1253 (N_1253,N_1196,N_1191);
nand U1254 (N_1254,N_1159,N_1117);
nand U1255 (N_1255,N_1105,N_1159);
and U1256 (N_1256,N_1112,N_1198);
or U1257 (N_1257,N_1184,N_1196);
nor U1258 (N_1258,N_1102,N_1191);
and U1259 (N_1259,N_1155,N_1186);
and U1260 (N_1260,N_1191,N_1115);
nand U1261 (N_1261,N_1174,N_1185);
or U1262 (N_1262,N_1141,N_1154);
nor U1263 (N_1263,N_1170,N_1150);
or U1264 (N_1264,N_1181,N_1185);
nor U1265 (N_1265,N_1154,N_1159);
nor U1266 (N_1266,N_1159,N_1110);
nor U1267 (N_1267,N_1120,N_1185);
and U1268 (N_1268,N_1188,N_1113);
and U1269 (N_1269,N_1115,N_1146);
and U1270 (N_1270,N_1136,N_1143);
xnor U1271 (N_1271,N_1117,N_1114);
or U1272 (N_1272,N_1174,N_1171);
or U1273 (N_1273,N_1172,N_1134);
xnor U1274 (N_1274,N_1176,N_1112);
and U1275 (N_1275,N_1163,N_1102);
nor U1276 (N_1276,N_1153,N_1197);
nand U1277 (N_1277,N_1115,N_1184);
nand U1278 (N_1278,N_1198,N_1145);
nand U1279 (N_1279,N_1193,N_1185);
nor U1280 (N_1280,N_1185,N_1145);
nor U1281 (N_1281,N_1199,N_1180);
and U1282 (N_1282,N_1144,N_1140);
or U1283 (N_1283,N_1178,N_1156);
xor U1284 (N_1284,N_1100,N_1107);
xor U1285 (N_1285,N_1153,N_1191);
xor U1286 (N_1286,N_1145,N_1173);
or U1287 (N_1287,N_1162,N_1146);
nand U1288 (N_1288,N_1144,N_1194);
nand U1289 (N_1289,N_1146,N_1188);
or U1290 (N_1290,N_1105,N_1123);
and U1291 (N_1291,N_1189,N_1164);
or U1292 (N_1292,N_1183,N_1171);
nor U1293 (N_1293,N_1107,N_1172);
nor U1294 (N_1294,N_1194,N_1117);
and U1295 (N_1295,N_1104,N_1150);
xor U1296 (N_1296,N_1186,N_1129);
xnor U1297 (N_1297,N_1141,N_1158);
nor U1298 (N_1298,N_1181,N_1121);
and U1299 (N_1299,N_1129,N_1173);
and U1300 (N_1300,N_1207,N_1202);
and U1301 (N_1301,N_1250,N_1211);
nor U1302 (N_1302,N_1255,N_1238);
or U1303 (N_1303,N_1280,N_1213);
nor U1304 (N_1304,N_1226,N_1251);
and U1305 (N_1305,N_1212,N_1221);
and U1306 (N_1306,N_1246,N_1263);
xnor U1307 (N_1307,N_1292,N_1243);
nor U1308 (N_1308,N_1293,N_1296);
nand U1309 (N_1309,N_1286,N_1262);
nand U1310 (N_1310,N_1259,N_1297);
or U1311 (N_1311,N_1256,N_1275);
nor U1312 (N_1312,N_1294,N_1281);
xnor U1313 (N_1313,N_1288,N_1236);
nor U1314 (N_1314,N_1261,N_1248);
nand U1315 (N_1315,N_1219,N_1247);
or U1316 (N_1316,N_1244,N_1241);
nand U1317 (N_1317,N_1274,N_1205);
nor U1318 (N_1318,N_1204,N_1242);
xor U1319 (N_1319,N_1214,N_1231);
nor U1320 (N_1320,N_1253,N_1279);
and U1321 (N_1321,N_1267,N_1229);
nor U1322 (N_1322,N_1257,N_1249);
or U1323 (N_1323,N_1284,N_1218);
nand U1324 (N_1324,N_1287,N_1271);
nor U1325 (N_1325,N_1278,N_1210);
and U1326 (N_1326,N_1215,N_1264);
xor U1327 (N_1327,N_1299,N_1295);
xor U1328 (N_1328,N_1220,N_1254);
nand U1329 (N_1329,N_1222,N_1225);
nand U1330 (N_1330,N_1240,N_1270);
and U1331 (N_1331,N_1228,N_1230);
nand U1332 (N_1332,N_1239,N_1216);
or U1333 (N_1333,N_1260,N_1282);
and U1334 (N_1334,N_1203,N_1208);
or U1335 (N_1335,N_1283,N_1232);
nor U1336 (N_1336,N_1273,N_1298);
nand U1337 (N_1337,N_1258,N_1201);
nand U1338 (N_1338,N_1223,N_1224);
nand U1339 (N_1339,N_1235,N_1206);
nor U1340 (N_1340,N_1291,N_1289);
nor U1341 (N_1341,N_1265,N_1277);
nand U1342 (N_1342,N_1237,N_1276);
or U1343 (N_1343,N_1217,N_1227);
or U1344 (N_1344,N_1268,N_1285);
nand U1345 (N_1345,N_1272,N_1290);
nor U1346 (N_1346,N_1209,N_1269);
nor U1347 (N_1347,N_1200,N_1233);
and U1348 (N_1348,N_1266,N_1245);
xnor U1349 (N_1349,N_1252,N_1234);
or U1350 (N_1350,N_1213,N_1265);
xor U1351 (N_1351,N_1203,N_1284);
or U1352 (N_1352,N_1280,N_1285);
and U1353 (N_1353,N_1243,N_1272);
and U1354 (N_1354,N_1248,N_1290);
nand U1355 (N_1355,N_1278,N_1242);
and U1356 (N_1356,N_1232,N_1203);
nor U1357 (N_1357,N_1223,N_1231);
and U1358 (N_1358,N_1228,N_1280);
or U1359 (N_1359,N_1236,N_1216);
nand U1360 (N_1360,N_1262,N_1200);
xnor U1361 (N_1361,N_1237,N_1283);
xor U1362 (N_1362,N_1254,N_1262);
and U1363 (N_1363,N_1282,N_1204);
nand U1364 (N_1364,N_1274,N_1217);
xnor U1365 (N_1365,N_1206,N_1239);
nor U1366 (N_1366,N_1239,N_1297);
nand U1367 (N_1367,N_1298,N_1285);
or U1368 (N_1368,N_1255,N_1280);
or U1369 (N_1369,N_1230,N_1203);
nor U1370 (N_1370,N_1298,N_1245);
nor U1371 (N_1371,N_1242,N_1216);
and U1372 (N_1372,N_1234,N_1264);
or U1373 (N_1373,N_1264,N_1254);
nand U1374 (N_1374,N_1216,N_1264);
or U1375 (N_1375,N_1205,N_1238);
nand U1376 (N_1376,N_1212,N_1249);
or U1377 (N_1377,N_1247,N_1242);
or U1378 (N_1378,N_1246,N_1295);
or U1379 (N_1379,N_1263,N_1230);
and U1380 (N_1380,N_1273,N_1288);
nor U1381 (N_1381,N_1237,N_1282);
nor U1382 (N_1382,N_1258,N_1271);
nor U1383 (N_1383,N_1263,N_1209);
nor U1384 (N_1384,N_1282,N_1267);
or U1385 (N_1385,N_1206,N_1273);
nor U1386 (N_1386,N_1225,N_1290);
and U1387 (N_1387,N_1205,N_1272);
nand U1388 (N_1388,N_1230,N_1257);
and U1389 (N_1389,N_1253,N_1268);
nand U1390 (N_1390,N_1222,N_1241);
or U1391 (N_1391,N_1268,N_1292);
and U1392 (N_1392,N_1220,N_1222);
nor U1393 (N_1393,N_1267,N_1263);
or U1394 (N_1394,N_1265,N_1205);
or U1395 (N_1395,N_1254,N_1238);
and U1396 (N_1396,N_1277,N_1243);
and U1397 (N_1397,N_1288,N_1207);
or U1398 (N_1398,N_1245,N_1223);
nand U1399 (N_1399,N_1279,N_1223);
and U1400 (N_1400,N_1373,N_1367);
nor U1401 (N_1401,N_1375,N_1346);
nor U1402 (N_1402,N_1314,N_1302);
nor U1403 (N_1403,N_1307,N_1325);
and U1404 (N_1404,N_1322,N_1301);
or U1405 (N_1405,N_1377,N_1386);
nor U1406 (N_1406,N_1315,N_1394);
or U1407 (N_1407,N_1390,N_1328);
or U1408 (N_1408,N_1323,N_1310);
xor U1409 (N_1409,N_1398,N_1319);
or U1410 (N_1410,N_1330,N_1355);
or U1411 (N_1411,N_1313,N_1333);
nor U1412 (N_1412,N_1337,N_1353);
or U1413 (N_1413,N_1343,N_1397);
and U1414 (N_1414,N_1363,N_1356);
nand U1415 (N_1415,N_1344,N_1352);
and U1416 (N_1416,N_1336,N_1350);
nor U1417 (N_1417,N_1360,N_1385);
nor U1418 (N_1418,N_1393,N_1321);
nor U1419 (N_1419,N_1389,N_1304);
nor U1420 (N_1420,N_1349,N_1364);
or U1421 (N_1421,N_1388,N_1306);
xnor U1422 (N_1422,N_1361,N_1391);
nand U1423 (N_1423,N_1354,N_1387);
and U1424 (N_1424,N_1308,N_1311);
xnor U1425 (N_1425,N_1327,N_1326);
nor U1426 (N_1426,N_1317,N_1396);
xor U1427 (N_1427,N_1334,N_1358);
nand U1428 (N_1428,N_1342,N_1320);
or U1429 (N_1429,N_1303,N_1345);
or U1430 (N_1430,N_1347,N_1376);
nand U1431 (N_1431,N_1300,N_1369);
or U1432 (N_1432,N_1324,N_1331);
xor U1433 (N_1433,N_1332,N_1399);
and U1434 (N_1434,N_1374,N_1329);
nand U1435 (N_1435,N_1368,N_1340);
or U1436 (N_1436,N_1359,N_1362);
nor U1437 (N_1437,N_1372,N_1339);
xnor U1438 (N_1438,N_1309,N_1382);
nand U1439 (N_1439,N_1395,N_1341);
or U1440 (N_1440,N_1366,N_1348);
nor U1441 (N_1441,N_1380,N_1383);
nor U1442 (N_1442,N_1365,N_1378);
nor U1443 (N_1443,N_1312,N_1381);
xnor U1444 (N_1444,N_1338,N_1392);
nand U1445 (N_1445,N_1371,N_1384);
nand U1446 (N_1446,N_1357,N_1335);
nor U1447 (N_1447,N_1316,N_1318);
and U1448 (N_1448,N_1379,N_1305);
and U1449 (N_1449,N_1370,N_1351);
and U1450 (N_1450,N_1313,N_1307);
nor U1451 (N_1451,N_1378,N_1373);
nor U1452 (N_1452,N_1310,N_1369);
or U1453 (N_1453,N_1309,N_1307);
nand U1454 (N_1454,N_1318,N_1306);
and U1455 (N_1455,N_1354,N_1300);
nor U1456 (N_1456,N_1301,N_1365);
xnor U1457 (N_1457,N_1367,N_1335);
nand U1458 (N_1458,N_1334,N_1364);
nand U1459 (N_1459,N_1373,N_1395);
nand U1460 (N_1460,N_1344,N_1308);
and U1461 (N_1461,N_1321,N_1305);
nand U1462 (N_1462,N_1391,N_1314);
and U1463 (N_1463,N_1352,N_1394);
xor U1464 (N_1464,N_1326,N_1387);
nor U1465 (N_1465,N_1388,N_1383);
nor U1466 (N_1466,N_1335,N_1342);
nand U1467 (N_1467,N_1303,N_1318);
nand U1468 (N_1468,N_1376,N_1395);
nand U1469 (N_1469,N_1376,N_1325);
nor U1470 (N_1470,N_1341,N_1330);
nand U1471 (N_1471,N_1396,N_1355);
or U1472 (N_1472,N_1372,N_1303);
and U1473 (N_1473,N_1343,N_1379);
nand U1474 (N_1474,N_1323,N_1300);
nand U1475 (N_1475,N_1332,N_1373);
and U1476 (N_1476,N_1383,N_1386);
nor U1477 (N_1477,N_1376,N_1333);
or U1478 (N_1478,N_1303,N_1391);
nand U1479 (N_1479,N_1338,N_1357);
nand U1480 (N_1480,N_1363,N_1340);
or U1481 (N_1481,N_1324,N_1337);
xor U1482 (N_1482,N_1378,N_1330);
and U1483 (N_1483,N_1343,N_1380);
and U1484 (N_1484,N_1319,N_1321);
nor U1485 (N_1485,N_1396,N_1390);
nor U1486 (N_1486,N_1392,N_1334);
nor U1487 (N_1487,N_1309,N_1357);
xnor U1488 (N_1488,N_1373,N_1312);
and U1489 (N_1489,N_1339,N_1343);
nor U1490 (N_1490,N_1388,N_1395);
nand U1491 (N_1491,N_1352,N_1343);
nor U1492 (N_1492,N_1302,N_1385);
and U1493 (N_1493,N_1328,N_1335);
and U1494 (N_1494,N_1324,N_1341);
or U1495 (N_1495,N_1373,N_1340);
or U1496 (N_1496,N_1349,N_1392);
and U1497 (N_1497,N_1372,N_1300);
or U1498 (N_1498,N_1302,N_1350);
and U1499 (N_1499,N_1373,N_1322);
and U1500 (N_1500,N_1482,N_1453);
nor U1501 (N_1501,N_1449,N_1416);
nor U1502 (N_1502,N_1494,N_1441);
nor U1503 (N_1503,N_1408,N_1488);
or U1504 (N_1504,N_1429,N_1431);
nand U1505 (N_1505,N_1409,N_1450);
or U1506 (N_1506,N_1452,N_1443);
nor U1507 (N_1507,N_1402,N_1499);
or U1508 (N_1508,N_1444,N_1470);
nor U1509 (N_1509,N_1442,N_1497);
nor U1510 (N_1510,N_1465,N_1405);
nor U1511 (N_1511,N_1472,N_1483);
nand U1512 (N_1512,N_1463,N_1466);
nand U1513 (N_1513,N_1457,N_1477);
nor U1514 (N_1514,N_1435,N_1404);
nor U1515 (N_1515,N_1401,N_1460);
nor U1516 (N_1516,N_1490,N_1438);
or U1517 (N_1517,N_1403,N_1471);
and U1518 (N_1518,N_1493,N_1485);
nor U1519 (N_1519,N_1489,N_1418);
nand U1520 (N_1520,N_1479,N_1458);
nand U1521 (N_1521,N_1478,N_1400);
nand U1522 (N_1522,N_1439,N_1422);
xor U1523 (N_1523,N_1469,N_1445);
or U1524 (N_1524,N_1446,N_1423);
and U1525 (N_1525,N_1414,N_1424);
nor U1526 (N_1526,N_1498,N_1476);
or U1527 (N_1527,N_1406,N_1407);
or U1528 (N_1528,N_1459,N_1415);
xor U1529 (N_1529,N_1474,N_1433);
or U1530 (N_1530,N_1495,N_1484);
or U1531 (N_1531,N_1492,N_1454);
or U1532 (N_1532,N_1426,N_1491);
nand U1533 (N_1533,N_1487,N_1421);
or U1534 (N_1534,N_1486,N_1481);
xnor U1535 (N_1535,N_1437,N_1468);
or U1536 (N_1536,N_1447,N_1448);
xor U1537 (N_1537,N_1462,N_1425);
or U1538 (N_1538,N_1464,N_1413);
nand U1539 (N_1539,N_1411,N_1467);
nor U1540 (N_1540,N_1420,N_1456);
or U1541 (N_1541,N_1455,N_1461);
or U1542 (N_1542,N_1430,N_1440);
and U1543 (N_1543,N_1432,N_1417);
nand U1544 (N_1544,N_1436,N_1410);
nor U1545 (N_1545,N_1434,N_1412);
nand U1546 (N_1546,N_1427,N_1419);
and U1547 (N_1547,N_1480,N_1473);
and U1548 (N_1548,N_1496,N_1428);
nor U1549 (N_1549,N_1451,N_1475);
xnor U1550 (N_1550,N_1491,N_1481);
nor U1551 (N_1551,N_1448,N_1459);
and U1552 (N_1552,N_1442,N_1474);
or U1553 (N_1553,N_1498,N_1496);
or U1554 (N_1554,N_1496,N_1475);
and U1555 (N_1555,N_1438,N_1448);
and U1556 (N_1556,N_1417,N_1422);
xnor U1557 (N_1557,N_1431,N_1476);
and U1558 (N_1558,N_1416,N_1481);
nor U1559 (N_1559,N_1481,N_1412);
nand U1560 (N_1560,N_1433,N_1442);
nand U1561 (N_1561,N_1434,N_1455);
xor U1562 (N_1562,N_1468,N_1422);
and U1563 (N_1563,N_1494,N_1442);
xnor U1564 (N_1564,N_1478,N_1466);
or U1565 (N_1565,N_1493,N_1436);
xor U1566 (N_1566,N_1461,N_1481);
nor U1567 (N_1567,N_1451,N_1462);
nor U1568 (N_1568,N_1492,N_1420);
nor U1569 (N_1569,N_1425,N_1448);
xnor U1570 (N_1570,N_1414,N_1417);
nor U1571 (N_1571,N_1458,N_1443);
and U1572 (N_1572,N_1465,N_1425);
xnor U1573 (N_1573,N_1409,N_1459);
xnor U1574 (N_1574,N_1433,N_1439);
nor U1575 (N_1575,N_1480,N_1477);
and U1576 (N_1576,N_1431,N_1489);
nor U1577 (N_1577,N_1459,N_1410);
or U1578 (N_1578,N_1423,N_1456);
nand U1579 (N_1579,N_1490,N_1475);
nand U1580 (N_1580,N_1432,N_1405);
and U1581 (N_1581,N_1495,N_1431);
nor U1582 (N_1582,N_1445,N_1441);
nor U1583 (N_1583,N_1484,N_1407);
nor U1584 (N_1584,N_1401,N_1473);
and U1585 (N_1585,N_1427,N_1495);
or U1586 (N_1586,N_1422,N_1432);
and U1587 (N_1587,N_1444,N_1489);
and U1588 (N_1588,N_1450,N_1405);
nand U1589 (N_1589,N_1407,N_1495);
and U1590 (N_1590,N_1412,N_1443);
nor U1591 (N_1591,N_1467,N_1429);
nor U1592 (N_1592,N_1447,N_1495);
or U1593 (N_1593,N_1421,N_1445);
or U1594 (N_1594,N_1429,N_1448);
or U1595 (N_1595,N_1498,N_1430);
or U1596 (N_1596,N_1492,N_1486);
nor U1597 (N_1597,N_1463,N_1485);
or U1598 (N_1598,N_1457,N_1439);
nor U1599 (N_1599,N_1405,N_1440);
or U1600 (N_1600,N_1586,N_1543);
nor U1601 (N_1601,N_1596,N_1595);
and U1602 (N_1602,N_1560,N_1588);
nand U1603 (N_1603,N_1549,N_1551);
nand U1604 (N_1604,N_1507,N_1515);
xor U1605 (N_1605,N_1555,N_1517);
nand U1606 (N_1606,N_1525,N_1538);
or U1607 (N_1607,N_1541,N_1535);
nand U1608 (N_1608,N_1561,N_1574);
nor U1609 (N_1609,N_1562,N_1573);
nor U1610 (N_1610,N_1524,N_1556);
nand U1611 (N_1611,N_1542,N_1548);
nand U1612 (N_1612,N_1532,N_1563);
nand U1613 (N_1613,N_1554,N_1572);
nand U1614 (N_1614,N_1502,N_1504);
xor U1615 (N_1615,N_1570,N_1585);
nand U1616 (N_1616,N_1501,N_1534);
and U1617 (N_1617,N_1559,N_1568);
or U1618 (N_1618,N_1576,N_1581);
and U1619 (N_1619,N_1516,N_1506);
nand U1620 (N_1620,N_1567,N_1587);
nand U1621 (N_1621,N_1545,N_1510);
or U1622 (N_1622,N_1583,N_1584);
nand U1623 (N_1623,N_1527,N_1566);
or U1624 (N_1624,N_1552,N_1571);
and U1625 (N_1625,N_1591,N_1521);
or U1626 (N_1626,N_1536,N_1597);
nor U1627 (N_1627,N_1500,N_1557);
and U1628 (N_1628,N_1590,N_1528);
nand U1629 (N_1629,N_1533,N_1553);
nand U1630 (N_1630,N_1592,N_1544);
or U1631 (N_1631,N_1531,N_1580);
nand U1632 (N_1632,N_1582,N_1508);
xnor U1633 (N_1633,N_1514,N_1577);
xnor U1634 (N_1634,N_1579,N_1518);
or U1635 (N_1635,N_1513,N_1511);
nor U1636 (N_1636,N_1503,N_1594);
or U1637 (N_1637,N_1599,N_1537);
xnor U1638 (N_1638,N_1558,N_1509);
or U1639 (N_1639,N_1539,N_1520);
and U1640 (N_1640,N_1564,N_1598);
or U1641 (N_1641,N_1512,N_1530);
and U1642 (N_1642,N_1540,N_1505);
nand U1643 (N_1643,N_1523,N_1575);
and U1644 (N_1644,N_1546,N_1529);
xor U1645 (N_1645,N_1547,N_1550);
and U1646 (N_1646,N_1565,N_1593);
nor U1647 (N_1647,N_1522,N_1526);
nor U1648 (N_1648,N_1578,N_1519);
or U1649 (N_1649,N_1569,N_1589);
xnor U1650 (N_1650,N_1517,N_1519);
nor U1651 (N_1651,N_1593,N_1580);
nor U1652 (N_1652,N_1598,N_1501);
and U1653 (N_1653,N_1507,N_1591);
or U1654 (N_1654,N_1537,N_1584);
nor U1655 (N_1655,N_1559,N_1510);
or U1656 (N_1656,N_1525,N_1566);
xor U1657 (N_1657,N_1589,N_1532);
or U1658 (N_1658,N_1506,N_1501);
or U1659 (N_1659,N_1565,N_1503);
nor U1660 (N_1660,N_1501,N_1551);
nand U1661 (N_1661,N_1592,N_1509);
and U1662 (N_1662,N_1597,N_1573);
nand U1663 (N_1663,N_1516,N_1575);
nor U1664 (N_1664,N_1556,N_1586);
and U1665 (N_1665,N_1521,N_1566);
or U1666 (N_1666,N_1555,N_1515);
or U1667 (N_1667,N_1581,N_1519);
or U1668 (N_1668,N_1568,N_1560);
or U1669 (N_1669,N_1566,N_1569);
nand U1670 (N_1670,N_1540,N_1533);
and U1671 (N_1671,N_1508,N_1593);
xor U1672 (N_1672,N_1513,N_1562);
nand U1673 (N_1673,N_1514,N_1580);
nand U1674 (N_1674,N_1547,N_1505);
nor U1675 (N_1675,N_1587,N_1510);
or U1676 (N_1676,N_1521,N_1596);
and U1677 (N_1677,N_1570,N_1575);
or U1678 (N_1678,N_1526,N_1517);
and U1679 (N_1679,N_1587,N_1502);
nor U1680 (N_1680,N_1503,N_1551);
and U1681 (N_1681,N_1510,N_1561);
nor U1682 (N_1682,N_1540,N_1517);
or U1683 (N_1683,N_1573,N_1552);
nand U1684 (N_1684,N_1574,N_1505);
and U1685 (N_1685,N_1538,N_1518);
or U1686 (N_1686,N_1599,N_1538);
and U1687 (N_1687,N_1566,N_1570);
nor U1688 (N_1688,N_1547,N_1501);
nor U1689 (N_1689,N_1581,N_1540);
nor U1690 (N_1690,N_1525,N_1500);
or U1691 (N_1691,N_1514,N_1566);
nor U1692 (N_1692,N_1521,N_1547);
nand U1693 (N_1693,N_1500,N_1518);
or U1694 (N_1694,N_1580,N_1511);
and U1695 (N_1695,N_1549,N_1596);
or U1696 (N_1696,N_1580,N_1578);
nand U1697 (N_1697,N_1540,N_1539);
or U1698 (N_1698,N_1548,N_1560);
nor U1699 (N_1699,N_1586,N_1580);
and U1700 (N_1700,N_1615,N_1644);
nor U1701 (N_1701,N_1690,N_1653);
nor U1702 (N_1702,N_1607,N_1673);
nand U1703 (N_1703,N_1637,N_1624);
nor U1704 (N_1704,N_1601,N_1697);
nand U1705 (N_1705,N_1654,N_1619);
or U1706 (N_1706,N_1694,N_1617);
and U1707 (N_1707,N_1630,N_1614);
nand U1708 (N_1708,N_1600,N_1659);
xor U1709 (N_1709,N_1698,N_1610);
and U1710 (N_1710,N_1667,N_1687);
xnor U1711 (N_1711,N_1678,N_1662);
xnor U1712 (N_1712,N_1603,N_1666);
and U1713 (N_1713,N_1646,N_1629);
nand U1714 (N_1714,N_1650,N_1685);
or U1715 (N_1715,N_1648,N_1665);
and U1716 (N_1716,N_1649,N_1693);
xnor U1717 (N_1717,N_1608,N_1691);
or U1718 (N_1718,N_1627,N_1657);
xnor U1719 (N_1719,N_1626,N_1641);
xor U1720 (N_1720,N_1620,N_1605);
nand U1721 (N_1721,N_1651,N_1609);
or U1722 (N_1722,N_1677,N_1639);
xor U1723 (N_1723,N_1602,N_1622);
nor U1724 (N_1724,N_1632,N_1664);
xnor U1725 (N_1725,N_1671,N_1660);
or U1726 (N_1726,N_1613,N_1640);
and U1727 (N_1727,N_1672,N_1606);
nand U1728 (N_1728,N_1633,N_1686);
nor U1729 (N_1729,N_1699,N_1623);
or U1730 (N_1730,N_1611,N_1628);
xor U1731 (N_1731,N_1669,N_1621);
xnor U1732 (N_1732,N_1642,N_1638);
nor U1733 (N_1733,N_1604,N_1674);
nor U1734 (N_1734,N_1696,N_1635);
nand U1735 (N_1735,N_1680,N_1661);
and U1736 (N_1736,N_1652,N_1663);
xnor U1737 (N_1737,N_1647,N_1618);
nor U1738 (N_1738,N_1679,N_1634);
xor U1739 (N_1739,N_1675,N_1683);
or U1740 (N_1740,N_1656,N_1612);
and U1741 (N_1741,N_1668,N_1631);
nor U1742 (N_1742,N_1682,N_1645);
or U1743 (N_1743,N_1636,N_1625);
and U1744 (N_1744,N_1676,N_1643);
or U1745 (N_1745,N_1655,N_1616);
nor U1746 (N_1746,N_1688,N_1670);
and U1747 (N_1747,N_1695,N_1689);
or U1748 (N_1748,N_1684,N_1658);
nor U1749 (N_1749,N_1681,N_1692);
nor U1750 (N_1750,N_1666,N_1647);
and U1751 (N_1751,N_1609,N_1660);
nor U1752 (N_1752,N_1603,N_1674);
xor U1753 (N_1753,N_1612,N_1660);
or U1754 (N_1754,N_1635,N_1655);
xor U1755 (N_1755,N_1606,N_1651);
xor U1756 (N_1756,N_1631,N_1659);
nand U1757 (N_1757,N_1644,N_1661);
and U1758 (N_1758,N_1601,N_1625);
nor U1759 (N_1759,N_1623,N_1657);
nor U1760 (N_1760,N_1626,N_1638);
nand U1761 (N_1761,N_1606,N_1691);
nor U1762 (N_1762,N_1689,N_1616);
and U1763 (N_1763,N_1631,N_1644);
or U1764 (N_1764,N_1661,N_1635);
and U1765 (N_1765,N_1673,N_1663);
or U1766 (N_1766,N_1631,N_1653);
nand U1767 (N_1767,N_1686,N_1643);
nor U1768 (N_1768,N_1608,N_1634);
nand U1769 (N_1769,N_1624,N_1682);
and U1770 (N_1770,N_1626,N_1624);
and U1771 (N_1771,N_1686,N_1683);
nor U1772 (N_1772,N_1638,N_1687);
and U1773 (N_1773,N_1630,N_1678);
nand U1774 (N_1774,N_1624,N_1694);
and U1775 (N_1775,N_1620,N_1660);
nand U1776 (N_1776,N_1675,N_1695);
xnor U1777 (N_1777,N_1646,N_1685);
and U1778 (N_1778,N_1685,N_1671);
nor U1779 (N_1779,N_1639,N_1624);
xnor U1780 (N_1780,N_1604,N_1663);
and U1781 (N_1781,N_1654,N_1685);
nand U1782 (N_1782,N_1642,N_1633);
and U1783 (N_1783,N_1651,N_1655);
or U1784 (N_1784,N_1635,N_1622);
and U1785 (N_1785,N_1681,N_1654);
nand U1786 (N_1786,N_1608,N_1683);
xor U1787 (N_1787,N_1653,N_1695);
and U1788 (N_1788,N_1652,N_1619);
and U1789 (N_1789,N_1668,N_1609);
and U1790 (N_1790,N_1665,N_1623);
xor U1791 (N_1791,N_1674,N_1666);
nor U1792 (N_1792,N_1676,N_1608);
and U1793 (N_1793,N_1640,N_1628);
xnor U1794 (N_1794,N_1605,N_1631);
and U1795 (N_1795,N_1626,N_1614);
nand U1796 (N_1796,N_1641,N_1663);
nand U1797 (N_1797,N_1614,N_1603);
nand U1798 (N_1798,N_1696,N_1650);
nand U1799 (N_1799,N_1604,N_1645);
and U1800 (N_1800,N_1763,N_1766);
or U1801 (N_1801,N_1714,N_1750);
nand U1802 (N_1802,N_1724,N_1742);
and U1803 (N_1803,N_1701,N_1787);
and U1804 (N_1804,N_1770,N_1708);
xnor U1805 (N_1805,N_1751,N_1722);
xor U1806 (N_1806,N_1798,N_1749);
xnor U1807 (N_1807,N_1719,N_1728);
or U1808 (N_1808,N_1717,N_1703);
nor U1809 (N_1809,N_1760,N_1761);
xor U1810 (N_1810,N_1793,N_1744);
or U1811 (N_1811,N_1773,N_1738);
nand U1812 (N_1812,N_1780,N_1727);
nand U1813 (N_1813,N_1791,N_1764);
and U1814 (N_1814,N_1765,N_1733);
and U1815 (N_1815,N_1720,N_1759);
xor U1816 (N_1816,N_1711,N_1753);
nand U1817 (N_1817,N_1746,N_1707);
or U1818 (N_1818,N_1799,N_1739);
nor U1819 (N_1819,N_1758,N_1704);
nor U1820 (N_1820,N_1789,N_1771);
nand U1821 (N_1821,N_1754,N_1737);
nand U1822 (N_1822,N_1729,N_1716);
nor U1823 (N_1823,N_1777,N_1774);
or U1824 (N_1824,N_1775,N_1776);
and U1825 (N_1825,N_1752,N_1755);
or U1826 (N_1826,N_1783,N_1796);
nand U1827 (N_1827,N_1730,N_1778);
nand U1828 (N_1828,N_1762,N_1781);
or U1829 (N_1829,N_1710,N_1706);
nand U1830 (N_1830,N_1732,N_1757);
nand U1831 (N_1831,N_1745,N_1715);
and U1832 (N_1832,N_1794,N_1702);
nor U1833 (N_1833,N_1792,N_1782);
nor U1834 (N_1834,N_1731,N_1743);
xor U1835 (N_1835,N_1784,N_1734);
nand U1836 (N_1836,N_1705,N_1726);
and U1837 (N_1837,N_1788,N_1740);
or U1838 (N_1838,N_1718,N_1786);
and U1839 (N_1839,N_1769,N_1785);
or U1840 (N_1840,N_1713,N_1712);
nand U1841 (N_1841,N_1779,N_1795);
and U1842 (N_1842,N_1725,N_1736);
nor U1843 (N_1843,N_1709,N_1723);
nand U1844 (N_1844,N_1797,N_1756);
and U1845 (N_1845,N_1790,N_1768);
nand U1846 (N_1846,N_1767,N_1735);
or U1847 (N_1847,N_1700,N_1772);
and U1848 (N_1848,N_1741,N_1747);
xnor U1849 (N_1849,N_1748,N_1721);
or U1850 (N_1850,N_1756,N_1763);
or U1851 (N_1851,N_1727,N_1758);
and U1852 (N_1852,N_1703,N_1708);
nand U1853 (N_1853,N_1722,N_1765);
or U1854 (N_1854,N_1784,N_1712);
and U1855 (N_1855,N_1782,N_1781);
and U1856 (N_1856,N_1798,N_1745);
or U1857 (N_1857,N_1713,N_1759);
or U1858 (N_1858,N_1739,N_1742);
nand U1859 (N_1859,N_1731,N_1786);
and U1860 (N_1860,N_1798,N_1750);
nor U1861 (N_1861,N_1775,N_1717);
and U1862 (N_1862,N_1737,N_1722);
nand U1863 (N_1863,N_1717,N_1758);
nor U1864 (N_1864,N_1775,N_1706);
and U1865 (N_1865,N_1708,N_1761);
nand U1866 (N_1866,N_1722,N_1795);
nand U1867 (N_1867,N_1795,N_1717);
nand U1868 (N_1868,N_1790,N_1776);
or U1869 (N_1869,N_1799,N_1754);
xnor U1870 (N_1870,N_1759,N_1765);
and U1871 (N_1871,N_1722,N_1756);
and U1872 (N_1872,N_1784,N_1749);
and U1873 (N_1873,N_1745,N_1794);
nand U1874 (N_1874,N_1779,N_1784);
and U1875 (N_1875,N_1740,N_1726);
or U1876 (N_1876,N_1797,N_1779);
nand U1877 (N_1877,N_1738,N_1751);
nand U1878 (N_1878,N_1760,N_1786);
nor U1879 (N_1879,N_1773,N_1720);
nand U1880 (N_1880,N_1766,N_1770);
nor U1881 (N_1881,N_1777,N_1799);
nor U1882 (N_1882,N_1758,N_1733);
nand U1883 (N_1883,N_1715,N_1763);
nand U1884 (N_1884,N_1712,N_1754);
nor U1885 (N_1885,N_1748,N_1779);
nor U1886 (N_1886,N_1713,N_1782);
or U1887 (N_1887,N_1763,N_1798);
nor U1888 (N_1888,N_1749,N_1770);
and U1889 (N_1889,N_1762,N_1771);
or U1890 (N_1890,N_1749,N_1763);
nand U1891 (N_1891,N_1748,N_1731);
nand U1892 (N_1892,N_1796,N_1707);
nor U1893 (N_1893,N_1799,N_1716);
nand U1894 (N_1894,N_1762,N_1750);
nand U1895 (N_1895,N_1798,N_1788);
nor U1896 (N_1896,N_1700,N_1723);
nand U1897 (N_1897,N_1771,N_1748);
nand U1898 (N_1898,N_1781,N_1710);
or U1899 (N_1899,N_1764,N_1721);
or U1900 (N_1900,N_1837,N_1882);
nor U1901 (N_1901,N_1851,N_1834);
nand U1902 (N_1902,N_1850,N_1823);
or U1903 (N_1903,N_1864,N_1832);
or U1904 (N_1904,N_1858,N_1841);
nor U1905 (N_1905,N_1867,N_1830);
nor U1906 (N_1906,N_1838,N_1822);
nand U1907 (N_1907,N_1894,N_1859);
nor U1908 (N_1908,N_1805,N_1886);
or U1909 (N_1909,N_1809,N_1854);
nand U1910 (N_1910,N_1895,N_1857);
and U1911 (N_1911,N_1814,N_1802);
nand U1912 (N_1912,N_1807,N_1896);
nand U1913 (N_1913,N_1806,N_1884);
and U1914 (N_1914,N_1874,N_1892);
nand U1915 (N_1915,N_1828,N_1852);
or U1916 (N_1916,N_1803,N_1835);
nand U1917 (N_1917,N_1849,N_1875);
and U1918 (N_1918,N_1831,N_1813);
or U1919 (N_1919,N_1825,N_1848);
nor U1920 (N_1920,N_1898,N_1808);
xnor U1921 (N_1921,N_1820,N_1817);
nor U1922 (N_1922,N_1833,N_1826);
nand U1923 (N_1923,N_1870,N_1843);
or U1924 (N_1924,N_1887,N_1891);
and U1925 (N_1925,N_1866,N_1880);
and U1926 (N_1926,N_1893,N_1844);
or U1927 (N_1927,N_1873,N_1876);
nand U1928 (N_1928,N_1804,N_1871);
nand U1929 (N_1929,N_1872,N_1862);
nor U1930 (N_1930,N_1861,N_1865);
nor U1931 (N_1931,N_1869,N_1812);
nor U1932 (N_1932,N_1889,N_1897);
nand U1933 (N_1933,N_1836,N_1824);
and U1934 (N_1934,N_1800,N_1810);
and U1935 (N_1935,N_1890,N_1815);
nor U1936 (N_1936,N_1856,N_1879);
or U1937 (N_1937,N_1863,N_1811);
or U1938 (N_1938,N_1801,N_1816);
and U1939 (N_1939,N_1855,N_1881);
nand U1940 (N_1940,N_1868,N_1846);
and U1941 (N_1941,N_1842,N_1829);
or U1942 (N_1942,N_1860,N_1827);
or U1943 (N_1943,N_1840,N_1877);
nand U1944 (N_1944,N_1818,N_1853);
nor U1945 (N_1945,N_1883,N_1845);
or U1946 (N_1946,N_1839,N_1878);
xor U1947 (N_1947,N_1819,N_1885);
or U1948 (N_1948,N_1888,N_1847);
and U1949 (N_1949,N_1899,N_1821);
and U1950 (N_1950,N_1872,N_1812);
and U1951 (N_1951,N_1898,N_1899);
or U1952 (N_1952,N_1889,N_1824);
and U1953 (N_1953,N_1869,N_1862);
and U1954 (N_1954,N_1896,N_1802);
nand U1955 (N_1955,N_1821,N_1886);
and U1956 (N_1956,N_1829,N_1817);
nand U1957 (N_1957,N_1810,N_1849);
and U1958 (N_1958,N_1841,N_1884);
and U1959 (N_1959,N_1855,N_1830);
and U1960 (N_1960,N_1826,N_1809);
or U1961 (N_1961,N_1886,N_1808);
nand U1962 (N_1962,N_1812,N_1892);
and U1963 (N_1963,N_1855,N_1821);
and U1964 (N_1964,N_1832,N_1870);
and U1965 (N_1965,N_1889,N_1821);
nand U1966 (N_1966,N_1855,N_1835);
xnor U1967 (N_1967,N_1800,N_1826);
xnor U1968 (N_1968,N_1849,N_1887);
and U1969 (N_1969,N_1830,N_1837);
nor U1970 (N_1970,N_1838,N_1876);
nor U1971 (N_1971,N_1895,N_1809);
nor U1972 (N_1972,N_1862,N_1894);
and U1973 (N_1973,N_1817,N_1832);
and U1974 (N_1974,N_1867,N_1806);
and U1975 (N_1975,N_1842,N_1889);
nand U1976 (N_1976,N_1806,N_1837);
nor U1977 (N_1977,N_1853,N_1852);
xnor U1978 (N_1978,N_1884,N_1816);
nand U1979 (N_1979,N_1850,N_1895);
or U1980 (N_1980,N_1896,N_1894);
xnor U1981 (N_1981,N_1850,N_1893);
and U1982 (N_1982,N_1801,N_1802);
nand U1983 (N_1983,N_1815,N_1854);
or U1984 (N_1984,N_1890,N_1843);
nand U1985 (N_1985,N_1833,N_1892);
and U1986 (N_1986,N_1896,N_1855);
or U1987 (N_1987,N_1860,N_1840);
nor U1988 (N_1988,N_1835,N_1845);
nand U1989 (N_1989,N_1812,N_1888);
or U1990 (N_1990,N_1855,N_1847);
or U1991 (N_1991,N_1812,N_1876);
nor U1992 (N_1992,N_1808,N_1802);
nand U1993 (N_1993,N_1869,N_1899);
or U1994 (N_1994,N_1856,N_1838);
and U1995 (N_1995,N_1863,N_1896);
nor U1996 (N_1996,N_1824,N_1879);
and U1997 (N_1997,N_1825,N_1883);
and U1998 (N_1998,N_1899,N_1884);
nand U1999 (N_1999,N_1882,N_1871);
or U2000 (N_2000,N_1912,N_1923);
or U2001 (N_2001,N_1909,N_1953);
nor U2002 (N_2002,N_1969,N_1908);
nand U2003 (N_2003,N_1967,N_1996);
nand U2004 (N_2004,N_1907,N_1966);
or U2005 (N_2005,N_1951,N_1934);
and U2006 (N_2006,N_1994,N_1919);
and U2007 (N_2007,N_1927,N_1900);
nand U2008 (N_2008,N_1988,N_1992);
nor U2009 (N_2009,N_1942,N_1957);
and U2010 (N_2010,N_1903,N_1930);
and U2011 (N_2011,N_1965,N_1901);
nand U2012 (N_2012,N_1933,N_1925);
or U2013 (N_2013,N_1920,N_1911);
and U2014 (N_2014,N_1939,N_1941);
nor U2015 (N_2015,N_1928,N_1982);
nor U2016 (N_2016,N_1998,N_1981);
nand U2017 (N_2017,N_1945,N_1987);
nand U2018 (N_2018,N_1980,N_1932);
or U2019 (N_2019,N_1955,N_1976);
nand U2020 (N_2020,N_1958,N_1962);
nor U2021 (N_2021,N_1915,N_1947);
nor U2022 (N_2022,N_1940,N_1959);
and U2023 (N_2023,N_1999,N_1902);
and U2024 (N_2024,N_1956,N_1917);
or U2025 (N_2025,N_1970,N_1950);
nand U2026 (N_2026,N_1937,N_1910);
or U2027 (N_2027,N_1936,N_1926);
nand U2028 (N_2028,N_1963,N_1979);
nor U2029 (N_2029,N_1914,N_1991);
and U2030 (N_2030,N_1972,N_1968);
nand U2031 (N_2031,N_1931,N_1993);
nand U2032 (N_2032,N_1971,N_1983);
nand U2033 (N_2033,N_1948,N_1904);
or U2034 (N_2034,N_1978,N_1995);
xnor U2035 (N_2035,N_1949,N_1944);
xnor U2036 (N_2036,N_1924,N_1961);
or U2037 (N_2037,N_1938,N_1964);
or U2038 (N_2038,N_1905,N_1984);
and U2039 (N_2039,N_1989,N_1943);
xnor U2040 (N_2040,N_1977,N_1954);
nor U2041 (N_2041,N_1975,N_1974);
nand U2042 (N_2042,N_1986,N_1985);
nor U2043 (N_2043,N_1952,N_1973);
nand U2044 (N_2044,N_1916,N_1918);
and U2045 (N_2045,N_1921,N_1997);
nand U2046 (N_2046,N_1946,N_1990);
nand U2047 (N_2047,N_1906,N_1929);
or U2048 (N_2048,N_1960,N_1935);
or U2049 (N_2049,N_1922,N_1913);
or U2050 (N_2050,N_1974,N_1967);
xnor U2051 (N_2051,N_1929,N_1947);
and U2052 (N_2052,N_1968,N_1928);
nand U2053 (N_2053,N_1905,N_1958);
and U2054 (N_2054,N_1972,N_1998);
nand U2055 (N_2055,N_1991,N_1988);
and U2056 (N_2056,N_1973,N_1951);
or U2057 (N_2057,N_1965,N_1962);
nor U2058 (N_2058,N_1960,N_1996);
nand U2059 (N_2059,N_1997,N_1952);
and U2060 (N_2060,N_1967,N_1978);
nand U2061 (N_2061,N_1905,N_1903);
nor U2062 (N_2062,N_1965,N_1945);
nand U2063 (N_2063,N_1943,N_1991);
nand U2064 (N_2064,N_1960,N_1947);
nand U2065 (N_2065,N_1965,N_1932);
xnor U2066 (N_2066,N_1914,N_1933);
nor U2067 (N_2067,N_1940,N_1991);
and U2068 (N_2068,N_1946,N_1944);
nor U2069 (N_2069,N_1988,N_1953);
and U2070 (N_2070,N_1970,N_1925);
nor U2071 (N_2071,N_1984,N_1931);
and U2072 (N_2072,N_1981,N_1966);
nor U2073 (N_2073,N_1922,N_1937);
nand U2074 (N_2074,N_1951,N_1980);
and U2075 (N_2075,N_1965,N_1969);
nor U2076 (N_2076,N_1924,N_1996);
and U2077 (N_2077,N_1962,N_1977);
or U2078 (N_2078,N_1961,N_1939);
and U2079 (N_2079,N_1997,N_1979);
nand U2080 (N_2080,N_1910,N_1925);
or U2081 (N_2081,N_1929,N_1915);
and U2082 (N_2082,N_1960,N_1930);
nand U2083 (N_2083,N_1940,N_1923);
nand U2084 (N_2084,N_1910,N_1994);
nand U2085 (N_2085,N_1925,N_1981);
nor U2086 (N_2086,N_1929,N_1980);
nor U2087 (N_2087,N_1913,N_1955);
or U2088 (N_2088,N_1952,N_1972);
nand U2089 (N_2089,N_1995,N_1983);
and U2090 (N_2090,N_1974,N_1979);
or U2091 (N_2091,N_1900,N_1918);
and U2092 (N_2092,N_1988,N_1979);
or U2093 (N_2093,N_1918,N_1987);
or U2094 (N_2094,N_1917,N_1984);
xnor U2095 (N_2095,N_1965,N_1913);
nand U2096 (N_2096,N_1921,N_1952);
nand U2097 (N_2097,N_1902,N_1950);
nand U2098 (N_2098,N_1974,N_1938);
nor U2099 (N_2099,N_1975,N_1936);
nor U2100 (N_2100,N_2040,N_2043);
xnor U2101 (N_2101,N_2071,N_2097);
and U2102 (N_2102,N_2030,N_2062);
xnor U2103 (N_2103,N_2073,N_2024);
and U2104 (N_2104,N_2055,N_2023);
or U2105 (N_2105,N_2044,N_2057);
or U2106 (N_2106,N_2098,N_2060);
nand U2107 (N_2107,N_2018,N_2006);
nand U2108 (N_2108,N_2016,N_2058);
nor U2109 (N_2109,N_2011,N_2028);
nor U2110 (N_2110,N_2088,N_2029);
nand U2111 (N_2111,N_2004,N_2064);
or U2112 (N_2112,N_2091,N_2069);
or U2113 (N_2113,N_2054,N_2079);
or U2114 (N_2114,N_2019,N_2038);
or U2115 (N_2115,N_2086,N_2005);
or U2116 (N_2116,N_2012,N_2090);
nand U2117 (N_2117,N_2007,N_2052);
nor U2118 (N_2118,N_2095,N_2008);
and U2119 (N_2119,N_2065,N_2059);
and U2120 (N_2120,N_2042,N_2068);
nand U2121 (N_2121,N_2096,N_2049);
or U2122 (N_2122,N_2045,N_2020);
or U2123 (N_2123,N_2072,N_2081);
and U2124 (N_2124,N_2035,N_2092);
xnor U2125 (N_2125,N_2047,N_2032);
nand U2126 (N_2126,N_2075,N_2056);
and U2127 (N_2127,N_2046,N_2034);
nand U2128 (N_2128,N_2000,N_2041);
or U2129 (N_2129,N_2083,N_2022);
xor U2130 (N_2130,N_2027,N_2070);
nand U2131 (N_2131,N_2015,N_2010);
nor U2132 (N_2132,N_2001,N_2099);
xor U2133 (N_2133,N_2067,N_2066);
nand U2134 (N_2134,N_2026,N_2077);
nand U2135 (N_2135,N_2033,N_2050);
nor U2136 (N_2136,N_2036,N_2003);
nand U2137 (N_2137,N_2078,N_2021);
nand U2138 (N_2138,N_2009,N_2080);
nor U2139 (N_2139,N_2014,N_2017);
nor U2140 (N_2140,N_2025,N_2085);
nand U2141 (N_2141,N_2094,N_2039);
xor U2142 (N_2142,N_2087,N_2013);
nand U2143 (N_2143,N_2002,N_2061);
and U2144 (N_2144,N_2089,N_2084);
nor U2145 (N_2145,N_2053,N_2031);
xor U2146 (N_2146,N_2048,N_2082);
nand U2147 (N_2147,N_2076,N_2074);
and U2148 (N_2148,N_2051,N_2093);
or U2149 (N_2149,N_2037,N_2063);
nor U2150 (N_2150,N_2033,N_2053);
nor U2151 (N_2151,N_2048,N_2090);
nor U2152 (N_2152,N_2074,N_2008);
nand U2153 (N_2153,N_2015,N_2083);
and U2154 (N_2154,N_2019,N_2062);
and U2155 (N_2155,N_2064,N_2048);
nand U2156 (N_2156,N_2024,N_2053);
nand U2157 (N_2157,N_2040,N_2069);
and U2158 (N_2158,N_2016,N_2089);
xor U2159 (N_2159,N_2008,N_2027);
or U2160 (N_2160,N_2009,N_2072);
or U2161 (N_2161,N_2064,N_2025);
nor U2162 (N_2162,N_2017,N_2058);
nor U2163 (N_2163,N_2043,N_2067);
nand U2164 (N_2164,N_2084,N_2087);
and U2165 (N_2165,N_2051,N_2080);
nand U2166 (N_2166,N_2044,N_2017);
or U2167 (N_2167,N_2062,N_2001);
nand U2168 (N_2168,N_2050,N_2028);
xor U2169 (N_2169,N_2037,N_2025);
nand U2170 (N_2170,N_2050,N_2084);
or U2171 (N_2171,N_2011,N_2069);
nor U2172 (N_2172,N_2023,N_2039);
nor U2173 (N_2173,N_2002,N_2099);
xnor U2174 (N_2174,N_2010,N_2048);
or U2175 (N_2175,N_2071,N_2006);
nor U2176 (N_2176,N_2086,N_2053);
nor U2177 (N_2177,N_2004,N_2086);
and U2178 (N_2178,N_2086,N_2094);
and U2179 (N_2179,N_2065,N_2028);
or U2180 (N_2180,N_2084,N_2024);
or U2181 (N_2181,N_2024,N_2093);
nor U2182 (N_2182,N_2036,N_2017);
nand U2183 (N_2183,N_2035,N_2019);
or U2184 (N_2184,N_2022,N_2013);
nand U2185 (N_2185,N_2010,N_2056);
nor U2186 (N_2186,N_2033,N_2045);
nand U2187 (N_2187,N_2070,N_2010);
nand U2188 (N_2188,N_2024,N_2017);
nand U2189 (N_2189,N_2042,N_2002);
or U2190 (N_2190,N_2072,N_2007);
and U2191 (N_2191,N_2003,N_2043);
or U2192 (N_2192,N_2004,N_2045);
nand U2193 (N_2193,N_2006,N_2028);
and U2194 (N_2194,N_2005,N_2076);
nor U2195 (N_2195,N_2082,N_2039);
nor U2196 (N_2196,N_2031,N_2085);
and U2197 (N_2197,N_2034,N_2033);
nand U2198 (N_2198,N_2024,N_2043);
xor U2199 (N_2199,N_2094,N_2008);
or U2200 (N_2200,N_2116,N_2173);
nor U2201 (N_2201,N_2104,N_2169);
nor U2202 (N_2202,N_2127,N_2162);
and U2203 (N_2203,N_2160,N_2120);
nor U2204 (N_2204,N_2154,N_2176);
and U2205 (N_2205,N_2103,N_2178);
nor U2206 (N_2206,N_2135,N_2150);
nand U2207 (N_2207,N_2138,N_2111);
or U2208 (N_2208,N_2145,N_2128);
or U2209 (N_2209,N_2119,N_2121);
or U2210 (N_2210,N_2110,N_2112);
or U2211 (N_2211,N_2107,N_2199);
nor U2212 (N_2212,N_2186,N_2157);
nor U2213 (N_2213,N_2122,N_2123);
nand U2214 (N_2214,N_2167,N_2161);
nand U2215 (N_2215,N_2194,N_2106);
and U2216 (N_2216,N_2153,N_2180);
nor U2217 (N_2217,N_2144,N_2170);
or U2218 (N_2218,N_2155,N_2134);
nand U2219 (N_2219,N_2195,N_2183);
nand U2220 (N_2220,N_2172,N_2114);
nor U2221 (N_2221,N_2189,N_2164);
and U2222 (N_2222,N_2102,N_2175);
nand U2223 (N_2223,N_2137,N_2129);
nor U2224 (N_2224,N_2156,N_2197);
nand U2225 (N_2225,N_2117,N_2124);
nand U2226 (N_2226,N_2130,N_2152);
and U2227 (N_2227,N_2190,N_2198);
and U2228 (N_2228,N_2146,N_2131);
nand U2229 (N_2229,N_2147,N_2177);
nor U2230 (N_2230,N_2181,N_2118);
nor U2231 (N_2231,N_2196,N_2168);
nand U2232 (N_2232,N_2105,N_2132);
xnor U2233 (N_2233,N_2140,N_2100);
nand U2234 (N_2234,N_2184,N_2142);
nor U2235 (N_2235,N_2141,N_2187);
nand U2236 (N_2236,N_2192,N_2174);
nor U2237 (N_2237,N_2185,N_2166);
xor U2238 (N_2238,N_2182,N_2151);
nor U2239 (N_2239,N_2159,N_2139);
and U2240 (N_2240,N_2126,N_2136);
nor U2241 (N_2241,N_2149,N_2125);
xor U2242 (N_2242,N_2115,N_2191);
xor U2243 (N_2243,N_2148,N_2193);
xnor U2244 (N_2244,N_2133,N_2188);
nor U2245 (N_2245,N_2101,N_2158);
nor U2246 (N_2246,N_2113,N_2143);
or U2247 (N_2247,N_2108,N_2163);
nor U2248 (N_2248,N_2179,N_2109);
nand U2249 (N_2249,N_2165,N_2171);
nor U2250 (N_2250,N_2180,N_2186);
nor U2251 (N_2251,N_2106,N_2156);
or U2252 (N_2252,N_2101,N_2178);
nand U2253 (N_2253,N_2146,N_2182);
nand U2254 (N_2254,N_2131,N_2164);
xnor U2255 (N_2255,N_2111,N_2118);
nor U2256 (N_2256,N_2144,N_2118);
or U2257 (N_2257,N_2192,N_2124);
and U2258 (N_2258,N_2106,N_2108);
xor U2259 (N_2259,N_2185,N_2102);
or U2260 (N_2260,N_2113,N_2188);
nor U2261 (N_2261,N_2187,N_2138);
nor U2262 (N_2262,N_2171,N_2147);
or U2263 (N_2263,N_2159,N_2170);
xor U2264 (N_2264,N_2118,N_2191);
or U2265 (N_2265,N_2138,N_2196);
nor U2266 (N_2266,N_2159,N_2199);
or U2267 (N_2267,N_2174,N_2146);
xor U2268 (N_2268,N_2164,N_2107);
and U2269 (N_2269,N_2160,N_2107);
nor U2270 (N_2270,N_2180,N_2175);
nor U2271 (N_2271,N_2136,N_2145);
nand U2272 (N_2272,N_2163,N_2164);
and U2273 (N_2273,N_2113,N_2179);
nor U2274 (N_2274,N_2162,N_2161);
xor U2275 (N_2275,N_2173,N_2159);
nor U2276 (N_2276,N_2194,N_2100);
nor U2277 (N_2277,N_2185,N_2189);
nand U2278 (N_2278,N_2168,N_2178);
nor U2279 (N_2279,N_2159,N_2174);
or U2280 (N_2280,N_2166,N_2195);
xnor U2281 (N_2281,N_2190,N_2129);
xor U2282 (N_2282,N_2101,N_2116);
and U2283 (N_2283,N_2187,N_2191);
nor U2284 (N_2284,N_2149,N_2152);
or U2285 (N_2285,N_2133,N_2154);
xor U2286 (N_2286,N_2164,N_2171);
nand U2287 (N_2287,N_2126,N_2150);
or U2288 (N_2288,N_2188,N_2152);
and U2289 (N_2289,N_2107,N_2115);
xor U2290 (N_2290,N_2120,N_2140);
or U2291 (N_2291,N_2161,N_2144);
or U2292 (N_2292,N_2107,N_2180);
nor U2293 (N_2293,N_2101,N_2196);
and U2294 (N_2294,N_2193,N_2191);
nand U2295 (N_2295,N_2107,N_2156);
nor U2296 (N_2296,N_2189,N_2193);
nand U2297 (N_2297,N_2164,N_2113);
and U2298 (N_2298,N_2124,N_2178);
or U2299 (N_2299,N_2149,N_2148);
or U2300 (N_2300,N_2296,N_2264);
nand U2301 (N_2301,N_2249,N_2236);
nand U2302 (N_2302,N_2275,N_2200);
and U2303 (N_2303,N_2260,N_2235);
and U2304 (N_2304,N_2291,N_2294);
nand U2305 (N_2305,N_2225,N_2232);
nand U2306 (N_2306,N_2240,N_2212);
or U2307 (N_2307,N_2277,N_2227);
or U2308 (N_2308,N_2228,N_2286);
nand U2309 (N_2309,N_2205,N_2209);
and U2310 (N_2310,N_2245,N_2254);
xnor U2311 (N_2311,N_2268,N_2261);
xor U2312 (N_2312,N_2217,N_2231);
and U2313 (N_2313,N_2242,N_2239);
nor U2314 (N_2314,N_2215,N_2266);
or U2315 (N_2315,N_2219,N_2267);
or U2316 (N_2316,N_2211,N_2262);
and U2317 (N_2317,N_2226,N_2259);
nand U2318 (N_2318,N_2233,N_2270);
and U2319 (N_2319,N_2253,N_2281);
nor U2320 (N_2320,N_2288,N_2282);
or U2321 (N_2321,N_2251,N_2250);
nor U2322 (N_2322,N_2237,N_2284);
or U2323 (N_2323,N_2299,N_2252);
and U2324 (N_2324,N_2223,N_2273);
nand U2325 (N_2325,N_2213,N_2248);
or U2326 (N_2326,N_2269,N_2230);
nand U2327 (N_2327,N_2216,N_2214);
or U2328 (N_2328,N_2234,N_2210);
and U2329 (N_2329,N_2295,N_2255);
nor U2330 (N_2330,N_2283,N_2202);
or U2331 (N_2331,N_2297,N_2285);
xor U2332 (N_2332,N_2274,N_2224);
and U2333 (N_2333,N_2208,N_2289);
and U2334 (N_2334,N_2265,N_2203);
xor U2335 (N_2335,N_2280,N_2222);
xnor U2336 (N_2336,N_2258,N_2244);
nand U2337 (N_2337,N_2276,N_2204);
or U2338 (N_2338,N_2292,N_2271);
xnor U2339 (N_2339,N_2241,N_2218);
nand U2340 (N_2340,N_2206,N_2220);
xor U2341 (N_2341,N_2293,N_2272);
xor U2342 (N_2342,N_2246,N_2247);
or U2343 (N_2343,N_2229,N_2256);
and U2344 (N_2344,N_2243,N_2290);
nor U2345 (N_2345,N_2257,N_2201);
nor U2346 (N_2346,N_2287,N_2238);
nor U2347 (N_2347,N_2263,N_2221);
and U2348 (N_2348,N_2278,N_2207);
nor U2349 (N_2349,N_2279,N_2298);
nand U2350 (N_2350,N_2222,N_2245);
nor U2351 (N_2351,N_2235,N_2299);
nor U2352 (N_2352,N_2218,N_2272);
or U2353 (N_2353,N_2216,N_2297);
nand U2354 (N_2354,N_2233,N_2285);
xor U2355 (N_2355,N_2256,N_2278);
nand U2356 (N_2356,N_2296,N_2280);
or U2357 (N_2357,N_2268,N_2226);
nand U2358 (N_2358,N_2277,N_2274);
xnor U2359 (N_2359,N_2267,N_2251);
and U2360 (N_2360,N_2250,N_2289);
nor U2361 (N_2361,N_2268,N_2201);
or U2362 (N_2362,N_2250,N_2227);
nor U2363 (N_2363,N_2232,N_2254);
nand U2364 (N_2364,N_2298,N_2227);
and U2365 (N_2365,N_2239,N_2292);
and U2366 (N_2366,N_2231,N_2245);
and U2367 (N_2367,N_2294,N_2253);
nor U2368 (N_2368,N_2255,N_2283);
xnor U2369 (N_2369,N_2250,N_2212);
nor U2370 (N_2370,N_2259,N_2267);
or U2371 (N_2371,N_2221,N_2254);
and U2372 (N_2372,N_2213,N_2289);
nand U2373 (N_2373,N_2222,N_2242);
or U2374 (N_2374,N_2291,N_2257);
and U2375 (N_2375,N_2226,N_2275);
nor U2376 (N_2376,N_2223,N_2260);
nor U2377 (N_2377,N_2272,N_2289);
nor U2378 (N_2378,N_2220,N_2224);
nor U2379 (N_2379,N_2237,N_2267);
or U2380 (N_2380,N_2224,N_2253);
xor U2381 (N_2381,N_2265,N_2252);
or U2382 (N_2382,N_2259,N_2263);
or U2383 (N_2383,N_2221,N_2249);
nand U2384 (N_2384,N_2212,N_2273);
and U2385 (N_2385,N_2285,N_2299);
nor U2386 (N_2386,N_2294,N_2212);
nor U2387 (N_2387,N_2248,N_2201);
xnor U2388 (N_2388,N_2292,N_2277);
and U2389 (N_2389,N_2292,N_2275);
or U2390 (N_2390,N_2271,N_2237);
or U2391 (N_2391,N_2266,N_2202);
or U2392 (N_2392,N_2250,N_2224);
or U2393 (N_2393,N_2252,N_2230);
or U2394 (N_2394,N_2259,N_2200);
and U2395 (N_2395,N_2214,N_2261);
nor U2396 (N_2396,N_2247,N_2217);
nand U2397 (N_2397,N_2277,N_2261);
or U2398 (N_2398,N_2227,N_2209);
nand U2399 (N_2399,N_2201,N_2263);
nand U2400 (N_2400,N_2322,N_2373);
nor U2401 (N_2401,N_2398,N_2356);
nand U2402 (N_2402,N_2335,N_2321);
nor U2403 (N_2403,N_2358,N_2357);
and U2404 (N_2404,N_2395,N_2369);
or U2405 (N_2405,N_2380,N_2340);
nand U2406 (N_2406,N_2364,N_2330);
or U2407 (N_2407,N_2314,N_2325);
or U2408 (N_2408,N_2312,N_2302);
nor U2409 (N_2409,N_2390,N_2391);
nor U2410 (N_2410,N_2361,N_2393);
nand U2411 (N_2411,N_2304,N_2366);
or U2412 (N_2412,N_2328,N_2307);
or U2413 (N_2413,N_2367,N_2353);
or U2414 (N_2414,N_2336,N_2315);
or U2415 (N_2415,N_2348,N_2338);
nor U2416 (N_2416,N_2331,N_2308);
nor U2417 (N_2417,N_2389,N_2392);
nand U2418 (N_2418,N_2365,N_2327);
nand U2419 (N_2419,N_2386,N_2344);
nand U2420 (N_2420,N_2363,N_2313);
and U2421 (N_2421,N_2316,N_2379);
or U2422 (N_2422,N_2326,N_2396);
or U2423 (N_2423,N_2354,N_2329);
nor U2424 (N_2424,N_2384,N_2347);
nand U2425 (N_2425,N_2318,N_2349);
and U2426 (N_2426,N_2301,N_2323);
and U2427 (N_2427,N_2372,N_2311);
nor U2428 (N_2428,N_2360,N_2374);
nand U2429 (N_2429,N_2397,N_2300);
and U2430 (N_2430,N_2341,N_2383);
and U2431 (N_2431,N_2376,N_2320);
xnor U2432 (N_2432,N_2355,N_2350);
or U2433 (N_2433,N_2381,N_2375);
nand U2434 (N_2434,N_2362,N_2399);
or U2435 (N_2435,N_2343,N_2334);
nand U2436 (N_2436,N_2352,N_2310);
nor U2437 (N_2437,N_2317,N_2345);
and U2438 (N_2438,N_2319,N_2339);
xor U2439 (N_2439,N_2359,N_2378);
or U2440 (N_2440,N_2394,N_2377);
and U2441 (N_2441,N_2332,N_2324);
nand U2442 (N_2442,N_2303,N_2371);
nand U2443 (N_2443,N_2337,N_2351);
nand U2444 (N_2444,N_2346,N_2306);
nand U2445 (N_2445,N_2387,N_2305);
and U2446 (N_2446,N_2342,N_2370);
nor U2447 (N_2447,N_2368,N_2333);
or U2448 (N_2448,N_2309,N_2385);
nand U2449 (N_2449,N_2388,N_2382);
nor U2450 (N_2450,N_2371,N_2398);
xor U2451 (N_2451,N_2327,N_2311);
nor U2452 (N_2452,N_2387,N_2365);
nand U2453 (N_2453,N_2328,N_2304);
nand U2454 (N_2454,N_2367,N_2382);
and U2455 (N_2455,N_2386,N_2398);
or U2456 (N_2456,N_2396,N_2386);
nor U2457 (N_2457,N_2375,N_2372);
xnor U2458 (N_2458,N_2397,N_2312);
or U2459 (N_2459,N_2379,N_2398);
nand U2460 (N_2460,N_2305,N_2393);
nand U2461 (N_2461,N_2307,N_2314);
nor U2462 (N_2462,N_2333,N_2339);
nand U2463 (N_2463,N_2360,N_2319);
xor U2464 (N_2464,N_2340,N_2362);
xnor U2465 (N_2465,N_2335,N_2370);
nor U2466 (N_2466,N_2320,N_2361);
nand U2467 (N_2467,N_2305,N_2312);
nor U2468 (N_2468,N_2310,N_2336);
nand U2469 (N_2469,N_2360,N_2333);
or U2470 (N_2470,N_2307,N_2374);
nor U2471 (N_2471,N_2301,N_2315);
nor U2472 (N_2472,N_2390,N_2386);
nand U2473 (N_2473,N_2380,N_2399);
xnor U2474 (N_2474,N_2375,N_2358);
and U2475 (N_2475,N_2338,N_2368);
and U2476 (N_2476,N_2360,N_2358);
xnor U2477 (N_2477,N_2363,N_2392);
nand U2478 (N_2478,N_2328,N_2308);
xor U2479 (N_2479,N_2359,N_2379);
nor U2480 (N_2480,N_2324,N_2377);
or U2481 (N_2481,N_2323,N_2313);
and U2482 (N_2482,N_2300,N_2307);
nor U2483 (N_2483,N_2300,N_2348);
or U2484 (N_2484,N_2313,N_2393);
nand U2485 (N_2485,N_2386,N_2324);
or U2486 (N_2486,N_2362,N_2330);
nand U2487 (N_2487,N_2314,N_2381);
and U2488 (N_2488,N_2393,N_2390);
and U2489 (N_2489,N_2338,N_2385);
and U2490 (N_2490,N_2366,N_2330);
nor U2491 (N_2491,N_2394,N_2386);
and U2492 (N_2492,N_2303,N_2374);
or U2493 (N_2493,N_2310,N_2383);
nor U2494 (N_2494,N_2332,N_2346);
xor U2495 (N_2495,N_2384,N_2326);
or U2496 (N_2496,N_2386,N_2338);
or U2497 (N_2497,N_2322,N_2369);
and U2498 (N_2498,N_2392,N_2374);
nand U2499 (N_2499,N_2388,N_2341);
or U2500 (N_2500,N_2480,N_2477);
and U2501 (N_2501,N_2461,N_2426);
nor U2502 (N_2502,N_2428,N_2422);
nor U2503 (N_2503,N_2433,N_2406);
and U2504 (N_2504,N_2474,N_2441);
and U2505 (N_2505,N_2453,N_2458);
or U2506 (N_2506,N_2405,N_2479);
and U2507 (N_2507,N_2448,N_2416);
and U2508 (N_2508,N_2485,N_2491);
or U2509 (N_2509,N_2430,N_2459);
nand U2510 (N_2510,N_2411,N_2496);
and U2511 (N_2511,N_2463,N_2417);
xor U2512 (N_2512,N_2420,N_2499);
or U2513 (N_2513,N_2407,N_2478);
or U2514 (N_2514,N_2408,N_2414);
nor U2515 (N_2515,N_2452,N_2432);
nor U2516 (N_2516,N_2443,N_2442);
nor U2517 (N_2517,N_2415,N_2436);
nand U2518 (N_2518,N_2454,N_2427);
or U2519 (N_2519,N_2409,N_2412);
or U2520 (N_2520,N_2494,N_2423);
xnor U2521 (N_2521,N_2421,N_2465);
and U2522 (N_2522,N_2487,N_2482);
nor U2523 (N_2523,N_2456,N_2418);
xor U2524 (N_2524,N_2460,N_2488);
and U2525 (N_2525,N_2492,N_2447);
and U2526 (N_2526,N_2473,N_2413);
and U2527 (N_2527,N_2472,N_2400);
nor U2528 (N_2528,N_2437,N_2438);
nand U2529 (N_2529,N_2489,N_2449);
or U2530 (N_2530,N_2490,N_2434);
or U2531 (N_2531,N_2467,N_2431);
xnor U2532 (N_2532,N_2446,N_2468);
and U2533 (N_2533,N_2475,N_2451);
nor U2534 (N_2534,N_2495,N_2471);
or U2535 (N_2535,N_2498,N_2457);
xor U2536 (N_2536,N_2470,N_2404);
xor U2537 (N_2537,N_2450,N_2435);
and U2538 (N_2538,N_2419,N_2403);
nand U2539 (N_2539,N_2455,N_2476);
nor U2540 (N_2540,N_2469,N_2429);
or U2541 (N_2541,N_2486,N_2497);
and U2542 (N_2542,N_2402,N_2440);
and U2543 (N_2543,N_2445,N_2444);
or U2544 (N_2544,N_2462,N_2481);
and U2545 (N_2545,N_2483,N_2464);
nand U2546 (N_2546,N_2484,N_2424);
or U2547 (N_2547,N_2401,N_2466);
or U2548 (N_2548,N_2439,N_2425);
nor U2549 (N_2549,N_2410,N_2493);
nor U2550 (N_2550,N_2494,N_2427);
nand U2551 (N_2551,N_2486,N_2473);
nand U2552 (N_2552,N_2492,N_2465);
or U2553 (N_2553,N_2427,N_2459);
nor U2554 (N_2554,N_2466,N_2434);
nor U2555 (N_2555,N_2470,N_2459);
and U2556 (N_2556,N_2449,N_2443);
nor U2557 (N_2557,N_2440,N_2423);
and U2558 (N_2558,N_2427,N_2410);
or U2559 (N_2559,N_2497,N_2441);
or U2560 (N_2560,N_2496,N_2424);
and U2561 (N_2561,N_2435,N_2457);
or U2562 (N_2562,N_2465,N_2450);
and U2563 (N_2563,N_2418,N_2432);
nor U2564 (N_2564,N_2472,N_2491);
or U2565 (N_2565,N_2404,N_2447);
xnor U2566 (N_2566,N_2451,N_2467);
or U2567 (N_2567,N_2485,N_2409);
nor U2568 (N_2568,N_2448,N_2433);
and U2569 (N_2569,N_2497,N_2402);
nand U2570 (N_2570,N_2440,N_2441);
or U2571 (N_2571,N_2437,N_2465);
nor U2572 (N_2572,N_2451,N_2435);
nor U2573 (N_2573,N_2458,N_2412);
or U2574 (N_2574,N_2421,N_2410);
nor U2575 (N_2575,N_2493,N_2403);
and U2576 (N_2576,N_2411,N_2493);
and U2577 (N_2577,N_2401,N_2462);
xnor U2578 (N_2578,N_2410,N_2488);
and U2579 (N_2579,N_2441,N_2495);
and U2580 (N_2580,N_2420,N_2406);
nand U2581 (N_2581,N_2421,N_2489);
nor U2582 (N_2582,N_2424,N_2408);
nand U2583 (N_2583,N_2404,N_2420);
or U2584 (N_2584,N_2439,N_2432);
or U2585 (N_2585,N_2474,N_2430);
nand U2586 (N_2586,N_2468,N_2474);
and U2587 (N_2587,N_2452,N_2464);
nor U2588 (N_2588,N_2458,N_2443);
or U2589 (N_2589,N_2443,N_2437);
and U2590 (N_2590,N_2498,N_2464);
xnor U2591 (N_2591,N_2407,N_2498);
nor U2592 (N_2592,N_2455,N_2417);
nand U2593 (N_2593,N_2495,N_2475);
and U2594 (N_2594,N_2432,N_2460);
nand U2595 (N_2595,N_2437,N_2416);
nor U2596 (N_2596,N_2479,N_2420);
xnor U2597 (N_2597,N_2448,N_2438);
and U2598 (N_2598,N_2420,N_2413);
nor U2599 (N_2599,N_2465,N_2466);
and U2600 (N_2600,N_2571,N_2508);
nand U2601 (N_2601,N_2528,N_2512);
nand U2602 (N_2602,N_2559,N_2548);
or U2603 (N_2603,N_2521,N_2533);
nand U2604 (N_2604,N_2558,N_2522);
nand U2605 (N_2605,N_2573,N_2543);
or U2606 (N_2606,N_2503,N_2535);
nor U2607 (N_2607,N_2532,N_2516);
and U2608 (N_2608,N_2506,N_2501);
xnor U2609 (N_2609,N_2569,N_2529);
and U2610 (N_2610,N_2549,N_2593);
and U2611 (N_2611,N_2564,N_2557);
nor U2612 (N_2612,N_2589,N_2547);
nor U2613 (N_2613,N_2582,N_2597);
nand U2614 (N_2614,N_2513,N_2585);
nor U2615 (N_2615,N_2552,N_2575);
nand U2616 (N_2616,N_2541,N_2598);
and U2617 (N_2617,N_2504,N_2568);
xnor U2618 (N_2618,N_2500,N_2587);
or U2619 (N_2619,N_2550,N_2561);
or U2620 (N_2620,N_2525,N_2594);
nor U2621 (N_2621,N_2524,N_2572);
and U2622 (N_2622,N_2539,N_2537);
nor U2623 (N_2623,N_2517,N_2507);
and U2624 (N_2624,N_2565,N_2526);
or U2625 (N_2625,N_2514,N_2584);
or U2626 (N_2626,N_2530,N_2540);
nor U2627 (N_2627,N_2505,N_2544);
nand U2628 (N_2628,N_2579,N_2560);
or U2629 (N_2629,N_2546,N_2527);
nand U2630 (N_2630,N_2545,N_2583);
or U2631 (N_2631,N_2534,N_2580);
nand U2632 (N_2632,N_2566,N_2502);
nand U2633 (N_2633,N_2578,N_2536);
and U2634 (N_2634,N_2562,N_2590);
or U2635 (N_2635,N_2519,N_2518);
and U2636 (N_2636,N_2542,N_2555);
nand U2637 (N_2637,N_2599,N_2509);
xnor U2638 (N_2638,N_2551,N_2576);
and U2639 (N_2639,N_2563,N_2592);
nand U2640 (N_2640,N_2531,N_2570);
or U2641 (N_2641,N_2538,N_2591);
nor U2642 (N_2642,N_2515,N_2595);
xnor U2643 (N_2643,N_2586,N_2577);
and U2644 (N_2644,N_2523,N_2596);
xor U2645 (N_2645,N_2556,N_2574);
or U2646 (N_2646,N_2581,N_2567);
nor U2647 (N_2647,N_2553,N_2511);
and U2648 (N_2648,N_2520,N_2554);
and U2649 (N_2649,N_2588,N_2510);
and U2650 (N_2650,N_2593,N_2594);
nor U2651 (N_2651,N_2502,N_2576);
nor U2652 (N_2652,N_2562,N_2571);
and U2653 (N_2653,N_2522,N_2570);
and U2654 (N_2654,N_2570,N_2556);
nor U2655 (N_2655,N_2584,N_2503);
nand U2656 (N_2656,N_2518,N_2583);
or U2657 (N_2657,N_2508,N_2564);
or U2658 (N_2658,N_2569,N_2591);
nand U2659 (N_2659,N_2509,N_2594);
and U2660 (N_2660,N_2581,N_2576);
nand U2661 (N_2661,N_2512,N_2572);
and U2662 (N_2662,N_2534,N_2553);
and U2663 (N_2663,N_2541,N_2561);
and U2664 (N_2664,N_2514,N_2586);
xnor U2665 (N_2665,N_2574,N_2530);
xor U2666 (N_2666,N_2597,N_2563);
or U2667 (N_2667,N_2530,N_2578);
nand U2668 (N_2668,N_2527,N_2554);
nor U2669 (N_2669,N_2519,N_2565);
nand U2670 (N_2670,N_2548,N_2570);
nand U2671 (N_2671,N_2516,N_2506);
xor U2672 (N_2672,N_2564,N_2582);
or U2673 (N_2673,N_2500,N_2514);
nor U2674 (N_2674,N_2522,N_2539);
nor U2675 (N_2675,N_2579,N_2534);
nor U2676 (N_2676,N_2536,N_2511);
xor U2677 (N_2677,N_2559,N_2504);
nand U2678 (N_2678,N_2512,N_2536);
nor U2679 (N_2679,N_2514,N_2569);
nor U2680 (N_2680,N_2561,N_2559);
and U2681 (N_2681,N_2503,N_2528);
nor U2682 (N_2682,N_2583,N_2549);
and U2683 (N_2683,N_2575,N_2528);
or U2684 (N_2684,N_2577,N_2560);
nor U2685 (N_2685,N_2518,N_2529);
nand U2686 (N_2686,N_2517,N_2530);
nand U2687 (N_2687,N_2560,N_2535);
xor U2688 (N_2688,N_2561,N_2506);
nand U2689 (N_2689,N_2566,N_2517);
or U2690 (N_2690,N_2509,N_2539);
nor U2691 (N_2691,N_2555,N_2544);
nand U2692 (N_2692,N_2572,N_2563);
or U2693 (N_2693,N_2519,N_2541);
or U2694 (N_2694,N_2521,N_2592);
nand U2695 (N_2695,N_2598,N_2568);
and U2696 (N_2696,N_2537,N_2581);
and U2697 (N_2697,N_2552,N_2594);
or U2698 (N_2698,N_2531,N_2591);
or U2699 (N_2699,N_2582,N_2579);
or U2700 (N_2700,N_2677,N_2642);
xnor U2701 (N_2701,N_2655,N_2654);
or U2702 (N_2702,N_2694,N_2616);
and U2703 (N_2703,N_2653,N_2683);
nand U2704 (N_2704,N_2632,N_2673);
xor U2705 (N_2705,N_2675,N_2668);
xor U2706 (N_2706,N_2657,N_2663);
nand U2707 (N_2707,N_2609,N_2631);
xnor U2708 (N_2708,N_2699,N_2666);
or U2709 (N_2709,N_2624,N_2669);
or U2710 (N_2710,N_2630,N_2656);
or U2711 (N_2711,N_2672,N_2614);
or U2712 (N_2712,N_2648,N_2687);
and U2713 (N_2713,N_2639,N_2644);
nor U2714 (N_2714,N_2612,N_2617);
nand U2715 (N_2715,N_2660,N_2601);
nand U2716 (N_2716,N_2693,N_2633);
nand U2717 (N_2717,N_2627,N_2661);
nor U2718 (N_2718,N_2610,N_2618);
nand U2719 (N_2719,N_2606,N_2604);
and U2720 (N_2720,N_2638,N_2621);
or U2721 (N_2721,N_2646,N_2625);
or U2722 (N_2722,N_2615,N_2658);
or U2723 (N_2723,N_2695,N_2674);
nor U2724 (N_2724,N_2628,N_2652);
or U2725 (N_2725,N_2698,N_2662);
and U2726 (N_2726,N_2619,N_2620);
nand U2727 (N_2727,N_2600,N_2607);
or U2728 (N_2728,N_2636,N_2670);
nand U2729 (N_2729,N_2641,N_2651);
xnor U2730 (N_2730,N_2647,N_2686);
and U2731 (N_2731,N_2685,N_2691);
or U2732 (N_2732,N_2664,N_2667);
nor U2733 (N_2733,N_2679,N_2626);
nand U2734 (N_2734,N_2645,N_2684);
nor U2735 (N_2735,N_2602,N_2622);
nand U2736 (N_2736,N_2688,N_2605);
nand U2737 (N_2737,N_2637,N_2629);
or U2738 (N_2738,N_2613,N_2623);
and U2739 (N_2739,N_2692,N_2697);
nand U2740 (N_2740,N_2696,N_2689);
nor U2741 (N_2741,N_2649,N_2640);
nor U2742 (N_2742,N_2676,N_2659);
and U2743 (N_2743,N_2678,N_2608);
or U2744 (N_2744,N_2682,N_2634);
and U2745 (N_2745,N_2671,N_2643);
nor U2746 (N_2746,N_2650,N_2635);
nand U2747 (N_2747,N_2690,N_2665);
xor U2748 (N_2748,N_2681,N_2680);
nand U2749 (N_2749,N_2603,N_2611);
or U2750 (N_2750,N_2614,N_2667);
nand U2751 (N_2751,N_2658,N_2662);
and U2752 (N_2752,N_2639,N_2622);
nor U2753 (N_2753,N_2686,N_2642);
and U2754 (N_2754,N_2614,N_2617);
nand U2755 (N_2755,N_2618,N_2605);
or U2756 (N_2756,N_2644,N_2693);
or U2757 (N_2757,N_2657,N_2653);
nor U2758 (N_2758,N_2684,N_2694);
and U2759 (N_2759,N_2634,N_2619);
and U2760 (N_2760,N_2653,N_2698);
or U2761 (N_2761,N_2621,N_2676);
nand U2762 (N_2762,N_2674,N_2682);
or U2763 (N_2763,N_2681,N_2691);
and U2764 (N_2764,N_2606,N_2635);
nor U2765 (N_2765,N_2647,N_2680);
nor U2766 (N_2766,N_2656,N_2686);
xor U2767 (N_2767,N_2687,N_2647);
and U2768 (N_2768,N_2627,N_2682);
and U2769 (N_2769,N_2614,N_2648);
or U2770 (N_2770,N_2652,N_2646);
nand U2771 (N_2771,N_2637,N_2614);
and U2772 (N_2772,N_2617,N_2694);
and U2773 (N_2773,N_2660,N_2604);
xnor U2774 (N_2774,N_2651,N_2602);
and U2775 (N_2775,N_2656,N_2623);
nor U2776 (N_2776,N_2608,N_2610);
and U2777 (N_2777,N_2671,N_2633);
and U2778 (N_2778,N_2676,N_2680);
xor U2779 (N_2779,N_2605,N_2662);
nor U2780 (N_2780,N_2606,N_2664);
or U2781 (N_2781,N_2605,N_2694);
nand U2782 (N_2782,N_2652,N_2645);
xnor U2783 (N_2783,N_2658,N_2622);
nor U2784 (N_2784,N_2674,N_2650);
nor U2785 (N_2785,N_2657,N_2605);
or U2786 (N_2786,N_2675,N_2680);
nor U2787 (N_2787,N_2647,N_2659);
xor U2788 (N_2788,N_2658,N_2644);
nand U2789 (N_2789,N_2679,N_2610);
xnor U2790 (N_2790,N_2617,N_2669);
nor U2791 (N_2791,N_2653,N_2613);
xor U2792 (N_2792,N_2693,N_2682);
nand U2793 (N_2793,N_2661,N_2642);
nand U2794 (N_2794,N_2631,N_2646);
nand U2795 (N_2795,N_2659,N_2617);
nor U2796 (N_2796,N_2632,N_2694);
xor U2797 (N_2797,N_2678,N_2617);
xnor U2798 (N_2798,N_2648,N_2696);
nor U2799 (N_2799,N_2676,N_2685);
or U2800 (N_2800,N_2778,N_2708);
and U2801 (N_2801,N_2782,N_2785);
or U2802 (N_2802,N_2787,N_2719);
or U2803 (N_2803,N_2770,N_2756);
nand U2804 (N_2804,N_2753,N_2747);
nand U2805 (N_2805,N_2763,N_2722);
nor U2806 (N_2806,N_2779,N_2727);
and U2807 (N_2807,N_2709,N_2731);
and U2808 (N_2808,N_2766,N_2786);
or U2809 (N_2809,N_2714,N_2742);
xor U2810 (N_2810,N_2774,N_2755);
or U2811 (N_2811,N_2754,N_2768);
and U2812 (N_2812,N_2701,N_2797);
and U2813 (N_2813,N_2744,N_2791);
and U2814 (N_2814,N_2749,N_2759);
xnor U2815 (N_2815,N_2741,N_2724);
or U2816 (N_2816,N_2767,N_2734);
xnor U2817 (N_2817,N_2703,N_2798);
or U2818 (N_2818,N_2745,N_2783);
and U2819 (N_2819,N_2737,N_2750);
and U2820 (N_2820,N_2775,N_2769);
or U2821 (N_2821,N_2764,N_2748);
nand U2822 (N_2822,N_2712,N_2772);
or U2823 (N_2823,N_2796,N_2725);
and U2824 (N_2824,N_2777,N_2721);
or U2825 (N_2825,N_2700,N_2702);
nor U2826 (N_2826,N_2717,N_2784);
xnor U2827 (N_2827,N_2743,N_2762);
and U2828 (N_2828,N_2765,N_2790);
nand U2829 (N_2829,N_2780,N_2716);
or U2830 (N_2830,N_2726,N_2760);
or U2831 (N_2831,N_2752,N_2728);
or U2832 (N_2832,N_2799,N_2792);
or U2833 (N_2833,N_2781,N_2771);
nor U2834 (N_2834,N_2706,N_2705);
nand U2835 (N_2835,N_2713,N_2735);
nor U2836 (N_2836,N_2751,N_2788);
and U2837 (N_2837,N_2732,N_2746);
or U2838 (N_2838,N_2793,N_2733);
nor U2839 (N_2839,N_2757,N_2758);
nand U2840 (N_2840,N_2707,N_2730);
nand U2841 (N_2841,N_2776,N_2720);
and U2842 (N_2842,N_2729,N_2773);
xnor U2843 (N_2843,N_2794,N_2715);
nor U2844 (N_2844,N_2723,N_2795);
and U2845 (N_2845,N_2740,N_2718);
and U2846 (N_2846,N_2736,N_2711);
nand U2847 (N_2847,N_2738,N_2704);
nand U2848 (N_2848,N_2789,N_2761);
xnor U2849 (N_2849,N_2739,N_2710);
or U2850 (N_2850,N_2726,N_2794);
and U2851 (N_2851,N_2712,N_2778);
nand U2852 (N_2852,N_2729,N_2703);
or U2853 (N_2853,N_2724,N_2785);
nand U2854 (N_2854,N_2780,N_2726);
nor U2855 (N_2855,N_2758,N_2726);
or U2856 (N_2856,N_2765,N_2772);
nor U2857 (N_2857,N_2771,N_2766);
nor U2858 (N_2858,N_2720,N_2725);
xnor U2859 (N_2859,N_2733,N_2719);
and U2860 (N_2860,N_2743,N_2771);
and U2861 (N_2861,N_2772,N_2770);
or U2862 (N_2862,N_2760,N_2781);
nand U2863 (N_2863,N_2751,N_2715);
and U2864 (N_2864,N_2788,N_2735);
nor U2865 (N_2865,N_2749,N_2703);
nor U2866 (N_2866,N_2741,N_2714);
xor U2867 (N_2867,N_2739,N_2717);
nand U2868 (N_2868,N_2753,N_2782);
nand U2869 (N_2869,N_2751,N_2759);
and U2870 (N_2870,N_2725,N_2736);
nor U2871 (N_2871,N_2714,N_2783);
and U2872 (N_2872,N_2746,N_2759);
and U2873 (N_2873,N_2705,N_2757);
nand U2874 (N_2874,N_2709,N_2749);
nand U2875 (N_2875,N_2716,N_2765);
or U2876 (N_2876,N_2759,N_2756);
xor U2877 (N_2877,N_2763,N_2729);
and U2878 (N_2878,N_2725,N_2734);
and U2879 (N_2879,N_2748,N_2784);
nand U2880 (N_2880,N_2717,N_2751);
and U2881 (N_2881,N_2767,N_2713);
and U2882 (N_2882,N_2722,N_2717);
or U2883 (N_2883,N_2720,N_2797);
and U2884 (N_2884,N_2762,N_2729);
nor U2885 (N_2885,N_2735,N_2777);
nand U2886 (N_2886,N_2762,N_2700);
nor U2887 (N_2887,N_2702,N_2778);
nand U2888 (N_2888,N_2785,N_2773);
nand U2889 (N_2889,N_2777,N_2784);
and U2890 (N_2890,N_2761,N_2707);
xor U2891 (N_2891,N_2720,N_2740);
nor U2892 (N_2892,N_2742,N_2709);
nor U2893 (N_2893,N_2799,N_2784);
or U2894 (N_2894,N_2709,N_2717);
nand U2895 (N_2895,N_2751,N_2770);
and U2896 (N_2896,N_2797,N_2775);
nand U2897 (N_2897,N_2744,N_2723);
or U2898 (N_2898,N_2724,N_2777);
nor U2899 (N_2899,N_2767,N_2729);
nand U2900 (N_2900,N_2842,N_2821);
and U2901 (N_2901,N_2868,N_2833);
or U2902 (N_2902,N_2875,N_2890);
nand U2903 (N_2903,N_2835,N_2800);
nor U2904 (N_2904,N_2831,N_2845);
nand U2905 (N_2905,N_2824,N_2822);
nor U2906 (N_2906,N_2850,N_2826);
nand U2907 (N_2907,N_2847,N_2840);
or U2908 (N_2908,N_2805,N_2887);
xor U2909 (N_2909,N_2860,N_2878);
and U2910 (N_2910,N_2818,N_2883);
or U2911 (N_2911,N_2819,N_2872);
and U2912 (N_2912,N_2863,N_2852);
or U2913 (N_2913,N_2857,N_2886);
and U2914 (N_2914,N_2859,N_2884);
nand U2915 (N_2915,N_2877,N_2893);
nor U2916 (N_2916,N_2856,N_2885);
or U2917 (N_2917,N_2892,N_2849);
or U2918 (N_2918,N_2820,N_2825);
nor U2919 (N_2919,N_2843,N_2844);
nand U2920 (N_2920,N_2827,N_2891);
and U2921 (N_2921,N_2839,N_2836);
or U2922 (N_2922,N_2817,N_2816);
nand U2923 (N_2923,N_2804,N_2898);
nor U2924 (N_2924,N_2828,N_2874);
and U2925 (N_2925,N_2889,N_2851);
nand U2926 (N_2926,N_2834,N_2808);
or U2927 (N_2927,N_2866,N_2801);
nor U2928 (N_2928,N_2865,N_2858);
nand U2929 (N_2929,N_2854,N_2806);
nor U2930 (N_2930,N_2812,N_2837);
or U2931 (N_2931,N_2807,N_2811);
or U2932 (N_2932,N_2838,N_2888);
nand U2933 (N_2933,N_2830,N_2809);
xnor U2934 (N_2934,N_2873,N_2862);
and U2935 (N_2935,N_2895,N_2867);
nor U2936 (N_2936,N_2803,N_2861);
nand U2937 (N_2937,N_2853,N_2813);
and U2938 (N_2938,N_2832,N_2869);
and U2939 (N_2939,N_2870,N_2899);
nand U2940 (N_2940,N_2810,N_2896);
or U2941 (N_2941,N_2814,N_2881);
or U2942 (N_2942,N_2848,N_2871);
nor U2943 (N_2943,N_2876,N_2882);
and U2944 (N_2944,N_2841,N_2879);
and U2945 (N_2945,N_2829,N_2897);
xnor U2946 (N_2946,N_2802,N_2880);
nor U2947 (N_2947,N_2823,N_2894);
nor U2948 (N_2948,N_2815,N_2855);
and U2949 (N_2949,N_2846,N_2864);
or U2950 (N_2950,N_2862,N_2810);
and U2951 (N_2951,N_2848,N_2834);
nor U2952 (N_2952,N_2899,N_2873);
or U2953 (N_2953,N_2818,N_2832);
nor U2954 (N_2954,N_2818,N_2836);
or U2955 (N_2955,N_2899,N_2853);
or U2956 (N_2956,N_2852,N_2859);
or U2957 (N_2957,N_2819,N_2892);
or U2958 (N_2958,N_2831,N_2894);
and U2959 (N_2959,N_2833,N_2825);
nand U2960 (N_2960,N_2840,N_2873);
or U2961 (N_2961,N_2829,N_2854);
or U2962 (N_2962,N_2820,N_2898);
nand U2963 (N_2963,N_2849,N_2850);
and U2964 (N_2964,N_2803,N_2889);
nor U2965 (N_2965,N_2806,N_2872);
and U2966 (N_2966,N_2870,N_2821);
nor U2967 (N_2967,N_2848,N_2885);
nand U2968 (N_2968,N_2839,N_2866);
or U2969 (N_2969,N_2878,N_2865);
nor U2970 (N_2970,N_2894,N_2857);
nor U2971 (N_2971,N_2837,N_2880);
nor U2972 (N_2972,N_2832,N_2850);
nand U2973 (N_2973,N_2840,N_2869);
nor U2974 (N_2974,N_2835,N_2855);
nor U2975 (N_2975,N_2874,N_2827);
nor U2976 (N_2976,N_2881,N_2847);
xnor U2977 (N_2977,N_2896,N_2873);
and U2978 (N_2978,N_2830,N_2821);
and U2979 (N_2979,N_2871,N_2849);
nor U2980 (N_2980,N_2877,N_2895);
or U2981 (N_2981,N_2891,N_2863);
or U2982 (N_2982,N_2822,N_2895);
xor U2983 (N_2983,N_2838,N_2865);
nand U2984 (N_2984,N_2871,N_2813);
nand U2985 (N_2985,N_2831,N_2874);
and U2986 (N_2986,N_2878,N_2892);
nor U2987 (N_2987,N_2899,N_2801);
nand U2988 (N_2988,N_2852,N_2837);
nor U2989 (N_2989,N_2892,N_2873);
and U2990 (N_2990,N_2810,N_2811);
nand U2991 (N_2991,N_2861,N_2872);
or U2992 (N_2992,N_2818,N_2892);
and U2993 (N_2993,N_2803,N_2821);
or U2994 (N_2994,N_2825,N_2883);
and U2995 (N_2995,N_2891,N_2832);
and U2996 (N_2996,N_2861,N_2834);
or U2997 (N_2997,N_2832,N_2830);
or U2998 (N_2998,N_2892,N_2864);
and U2999 (N_2999,N_2830,N_2820);
xor U3000 (N_3000,N_2916,N_2909);
nand U3001 (N_3001,N_2945,N_2969);
nor U3002 (N_3002,N_2938,N_2998);
and U3003 (N_3003,N_2994,N_2977);
nand U3004 (N_3004,N_2927,N_2947);
nor U3005 (N_3005,N_2958,N_2979);
nand U3006 (N_3006,N_2954,N_2937);
nand U3007 (N_3007,N_2991,N_2974);
nor U3008 (N_3008,N_2972,N_2962);
nor U3009 (N_3009,N_2960,N_2997);
xnor U3010 (N_3010,N_2939,N_2934);
nand U3011 (N_3011,N_2956,N_2907);
or U3012 (N_3012,N_2982,N_2935);
xor U3013 (N_3013,N_2913,N_2924);
xor U3014 (N_3014,N_2946,N_2957);
or U3015 (N_3015,N_2908,N_2953);
or U3016 (N_3016,N_2901,N_2985);
nor U3017 (N_3017,N_2920,N_2900);
nor U3018 (N_3018,N_2989,N_2967);
and U3019 (N_3019,N_2968,N_2910);
and U3020 (N_3020,N_2949,N_2914);
nand U3021 (N_3021,N_2988,N_2943);
or U3022 (N_3022,N_2975,N_2993);
nor U3023 (N_3023,N_2990,N_2983);
nor U3024 (N_3024,N_2922,N_2941);
nand U3025 (N_3025,N_2948,N_2932);
nand U3026 (N_3026,N_2940,N_2930);
nand U3027 (N_3027,N_2919,N_2952);
nor U3028 (N_3028,N_2976,N_2951);
nand U3029 (N_3029,N_2961,N_2931);
nand U3030 (N_3030,N_2923,N_2942);
nand U3031 (N_3031,N_2987,N_2921);
and U3032 (N_3032,N_2965,N_2973);
nor U3033 (N_3033,N_2995,N_2964);
or U3034 (N_3034,N_2959,N_2929);
nand U3035 (N_3035,N_2905,N_2950);
nor U3036 (N_3036,N_2980,N_2902);
nor U3037 (N_3037,N_2903,N_2963);
or U3038 (N_3038,N_2999,N_2966);
nor U3039 (N_3039,N_2971,N_2992);
nor U3040 (N_3040,N_2911,N_2912);
or U3041 (N_3041,N_2978,N_2936);
nor U3042 (N_3042,N_2984,N_2904);
and U3043 (N_3043,N_2926,N_2915);
xor U3044 (N_3044,N_2928,N_2986);
nor U3045 (N_3045,N_2955,N_2944);
nand U3046 (N_3046,N_2933,N_2925);
nand U3047 (N_3047,N_2970,N_2981);
and U3048 (N_3048,N_2917,N_2996);
or U3049 (N_3049,N_2918,N_2906);
nor U3050 (N_3050,N_2906,N_2998);
xor U3051 (N_3051,N_2948,N_2958);
nor U3052 (N_3052,N_2946,N_2967);
and U3053 (N_3053,N_2948,N_2913);
nor U3054 (N_3054,N_2946,N_2945);
nor U3055 (N_3055,N_2925,N_2961);
or U3056 (N_3056,N_2979,N_2924);
nor U3057 (N_3057,N_2931,N_2913);
and U3058 (N_3058,N_2979,N_2934);
nor U3059 (N_3059,N_2909,N_2905);
nand U3060 (N_3060,N_2945,N_2919);
or U3061 (N_3061,N_2987,N_2977);
or U3062 (N_3062,N_2994,N_2967);
nor U3063 (N_3063,N_2953,N_2983);
and U3064 (N_3064,N_2938,N_2950);
nand U3065 (N_3065,N_2939,N_2902);
or U3066 (N_3066,N_2940,N_2963);
nand U3067 (N_3067,N_2916,N_2955);
and U3068 (N_3068,N_2902,N_2970);
xnor U3069 (N_3069,N_2977,N_2933);
and U3070 (N_3070,N_2996,N_2924);
nand U3071 (N_3071,N_2908,N_2927);
nor U3072 (N_3072,N_2902,N_2995);
nand U3073 (N_3073,N_2903,N_2912);
nand U3074 (N_3074,N_2917,N_2913);
xnor U3075 (N_3075,N_2952,N_2953);
or U3076 (N_3076,N_2908,N_2988);
xnor U3077 (N_3077,N_2991,N_2962);
nor U3078 (N_3078,N_2995,N_2923);
nor U3079 (N_3079,N_2914,N_2927);
xnor U3080 (N_3080,N_2972,N_2983);
or U3081 (N_3081,N_2932,N_2939);
or U3082 (N_3082,N_2901,N_2905);
xnor U3083 (N_3083,N_2929,N_2932);
nand U3084 (N_3084,N_2927,N_2952);
or U3085 (N_3085,N_2983,N_2947);
nand U3086 (N_3086,N_2921,N_2993);
and U3087 (N_3087,N_2909,N_2939);
or U3088 (N_3088,N_2926,N_2973);
xnor U3089 (N_3089,N_2993,N_2925);
nand U3090 (N_3090,N_2986,N_2905);
or U3091 (N_3091,N_2926,N_2969);
or U3092 (N_3092,N_2904,N_2910);
nor U3093 (N_3093,N_2948,N_2943);
and U3094 (N_3094,N_2963,N_2952);
nor U3095 (N_3095,N_2959,N_2923);
or U3096 (N_3096,N_2948,N_2954);
xnor U3097 (N_3097,N_2964,N_2974);
nor U3098 (N_3098,N_2907,N_2996);
nor U3099 (N_3099,N_2951,N_2974);
and U3100 (N_3100,N_3064,N_3082);
and U3101 (N_3101,N_3059,N_3029);
or U3102 (N_3102,N_3073,N_3021);
and U3103 (N_3103,N_3058,N_3062);
and U3104 (N_3104,N_3028,N_3051);
and U3105 (N_3105,N_3001,N_3002);
nand U3106 (N_3106,N_3008,N_3072);
or U3107 (N_3107,N_3093,N_3017);
or U3108 (N_3108,N_3066,N_3039);
xor U3109 (N_3109,N_3096,N_3025);
xor U3110 (N_3110,N_3015,N_3003);
and U3111 (N_3111,N_3010,N_3035);
and U3112 (N_3112,N_3049,N_3014);
xnor U3113 (N_3113,N_3032,N_3009);
and U3114 (N_3114,N_3084,N_3056);
or U3115 (N_3115,N_3006,N_3071);
nor U3116 (N_3116,N_3036,N_3026);
nand U3117 (N_3117,N_3092,N_3076);
nor U3118 (N_3118,N_3050,N_3098);
and U3119 (N_3119,N_3011,N_3068);
nor U3120 (N_3120,N_3048,N_3075);
xnor U3121 (N_3121,N_3054,N_3020);
nor U3122 (N_3122,N_3090,N_3085);
nor U3123 (N_3123,N_3018,N_3043);
and U3124 (N_3124,N_3079,N_3030);
or U3125 (N_3125,N_3069,N_3024);
and U3126 (N_3126,N_3094,N_3061);
and U3127 (N_3127,N_3040,N_3078);
nor U3128 (N_3128,N_3099,N_3000);
and U3129 (N_3129,N_3097,N_3004);
nor U3130 (N_3130,N_3022,N_3044);
and U3131 (N_3131,N_3019,N_3037);
and U3132 (N_3132,N_3038,N_3070);
nor U3133 (N_3133,N_3042,N_3041);
and U3134 (N_3134,N_3033,N_3034);
nand U3135 (N_3135,N_3005,N_3053);
or U3136 (N_3136,N_3023,N_3060);
nor U3137 (N_3137,N_3057,N_3065);
and U3138 (N_3138,N_3012,N_3083);
or U3139 (N_3139,N_3086,N_3007);
nand U3140 (N_3140,N_3013,N_3046);
xnor U3141 (N_3141,N_3091,N_3016);
and U3142 (N_3142,N_3031,N_3074);
xnor U3143 (N_3143,N_3027,N_3067);
and U3144 (N_3144,N_3095,N_3045);
or U3145 (N_3145,N_3088,N_3047);
or U3146 (N_3146,N_3055,N_3052);
and U3147 (N_3147,N_3063,N_3087);
nor U3148 (N_3148,N_3077,N_3080);
nor U3149 (N_3149,N_3081,N_3089);
xor U3150 (N_3150,N_3062,N_3065);
nor U3151 (N_3151,N_3034,N_3017);
nand U3152 (N_3152,N_3036,N_3006);
nor U3153 (N_3153,N_3047,N_3025);
nor U3154 (N_3154,N_3018,N_3086);
nor U3155 (N_3155,N_3046,N_3048);
or U3156 (N_3156,N_3058,N_3011);
nor U3157 (N_3157,N_3050,N_3070);
nor U3158 (N_3158,N_3067,N_3058);
nand U3159 (N_3159,N_3005,N_3070);
nor U3160 (N_3160,N_3099,N_3058);
nand U3161 (N_3161,N_3086,N_3040);
nor U3162 (N_3162,N_3036,N_3040);
nand U3163 (N_3163,N_3044,N_3001);
or U3164 (N_3164,N_3057,N_3085);
xnor U3165 (N_3165,N_3053,N_3072);
nand U3166 (N_3166,N_3026,N_3020);
xnor U3167 (N_3167,N_3075,N_3052);
xor U3168 (N_3168,N_3034,N_3036);
and U3169 (N_3169,N_3008,N_3090);
or U3170 (N_3170,N_3038,N_3074);
and U3171 (N_3171,N_3037,N_3007);
or U3172 (N_3172,N_3016,N_3030);
nor U3173 (N_3173,N_3086,N_3062);
or U3174 (N_3174,N_3041,N_3059);
or U3175 (N_3175,N_3095,N_3032);
xor U3176 (N_3176,N_3063,N_3064);
or U3177 (N_3177,N_3083,N_3080);
xor U3178 (N_3178,N_3057,N_3074);
nand U3179 (N_3179,N_3011,N_3064);
and U3180 (N_3180,N_3049,N_3043);
xor U3181 (N_3181,N_3064,N_3031);
nand U3182 (N_3182,N_3042,N_3070);
or U3183 (N_3183,N_3079,N_3094);
and U3184 (N_3184,N_3042,N_3061);
nor U3185 (N_3185,N_3088,N_3016);
nand U3186 (N_3186,N_3097,N_3001);
and U3187 (N_3187,N_3096,N_3012);
or U3188 (N_3188,N_3050,N_3080);
nand U3189 (N_3189,N_3034,N_3079);
or U3190 (N_3190,N_3081,N_3085);
nand U3191 (N_3191,N_3084,N_3001);
and U3192 (N_3192,N_3030,N_3003);
and U3193 (N_3193,N_3015,N_3080);
and U3194 (N_3194,N_3046,N_3034);
or U3195 (N_3195,N_3012,N_3098);
nand U3196 (N_3196,N_3093,N_3068);
nor U3197 (N_3197,N_3083,N_3093);
and U3198 (N_3198,N_3007,N_3071);
nand U3199 (N_3199,N_3057,N_3041);
nor U3200 (N_3200,N_3182,N_3142);
nor U3201 (N_3201,N_3169,N_3132);
nor U3202 (N_3202,N_3187,N_3114);
nor U3203 (N_3203,N_3147,N_3136);
and U3204 (N_3204,N_3190,N_3155);
and U3205 (N_3205,N_3143,N_3118);
and U3206 (N_3206,N_3111,N_3141);
or U3207 (N_3207,N_3102,N_3161);
and U3208 (N_3208,N_3140,N_3146);
xor U3209 (N_3209,N_3157,N_3144);
and U3210 (N_3210,N_3123,N_3103);
and U3211 (N_3211,N_3180,N_3110);
nor U3212 (N_3212,N_3167,N_3129);
and U3213 (N_3213,N_3189,N_3191);
nor U3214 (N_3214,N_3122,N_3130);
nor U3215 (N_3215,N_3174,N_3100);
nor U3216 (N_3216,N_3153,N_3178);
nor U3217 (N_3217,N_3115,N_3168);
nand U3218 (N_3218,N_3109,N_3158);
nand U3219 (N_3219,N_3116,N_3193);
nor U3220 (N_3220,N_3131,N_3192);
nor U3221 (N_3221,N_3112,N_3134);
nand U3222 (N_3222,N_3170,N_3176);
and U3223 (N_3223,N_3166,N_3175);
and U3224 (N_3224,N_3198,N_3183);
or U3225 (N_3225,N_3117,N_3188);
nor U3226 (N_3226,N_3186,N_3108);
or U3227 (N_3227,N_3120,N_3151);
nand U3228 (N_3228,N_3159,N_3162);
nand U3229 (N_3229,N_3152,N_3139);
or U3230 (N_3230,N_3199,N_3126);
xnor U3231 (N_3231,N_3154,N_3119);
or U3232 (N_3232,N_3156,N_3160);
and U3233 (N_3233,N_3172,N_3163);
and U3234 (N_3234,N_3164,N_3177);
nor U3235 (N_3235,N_3150,N_3104);
and U3236 (N_3236,N_3181,N_3194);
and U3237 (N_3237,N_3106,N_3128);
nand U3238 (N_3238,N_3135,N_3145);
nor U3239 (N_3239,N_3121,N_3105);
or U3240 (N_3240,N_3185,N_3138);
or U3241 (N_3241,N_3173,N_3133);
or U3242 (N_3242,N_3184,N_3179);
xnor U3243 (N_3243,N_3197,N_3171);
and U3244 (N_3244,N_3149,N_3107);
nand U3245 (N_3245,N_3148,N_3124);
or U3246 (N_3246,N_3137,N_3125);
nor U3247 (N_3247,N_3127,N_3101);
nand U3248 (N_3248,N_3165,N_3196);
or U3249 (N_3249,N_3195,N_3113);
and U3250 (N_3250,N_3114,N_3197);
and U3251 (N_3251,N_3177,N_3104);
and U3252 (N_3252,N_3112,N_3120);
or U3253 (N_3253,N_3191,N_3126);
or U3254 (N_3254,N_3102,N_3153);
nand U3255 (N_3255,N_3144,N_3153);
or U3256 (N_3256,N_3164,N_3154);
nand U3257 (N_3257,N_3153,N_3114);
xor U3258 (N_3258,N_3117,N_3198);
or U3259 (N_3259,N_3125,N_3193);
nor U3260 (N_3260,N_3198,N_3152);
nand U3261 (N_3261,N_3149,N_3156);
nor U3262 (N_3262,N_3191,N_3167);
nor U3263 (N_3263,N_3120,N_3116);
nor U3264 (N_3264,N_3151,N_3117);
nor U3265 (N_3265,N_3116,N_3151);
nand U3266 (N_3266,N_3114,N_3148);
xnor U3267 (N_3267,N_3148,N_3167);
or U3268 (N_3268,N_3135,N_3143);
or U3269 (N_3269,N_3154,N_3113);
xnor U3270 (N_3270,N_3119,N_3168);
or U3271 (N_3271,N_3124,N_3128);
nand U3272 (N_3272,N_3184,N_3138);
nand U3273 (N_3273,N_3102,N_3156);
and U3274 (N_3274,N_3133,N_3117);
or U3275 (N_3275,N_3180,N_3148);
or U3276 (N_3276,N_3121,N_3165);
nand U3277 (N_3277,N_3120,N_3165);
nor U3278 (N_3278,N_3174,N_3164);
nor U3279 (N_3279,N_3144,N_3106);
nor U3280 (N_3280,N_3103,N_3104);
nand U3281 (N_3281,N_3164,N_3172);
nor U3282 (N_3282,N_3105,N_3112);
nand U3283 (N_3283,N_3132,N_3141);
and U3284 (N_3284,N_3185,N_3168);
or U3285 (N_3285,N_3181,N_3163);
nand U3286 (N_3286,N_3199,N_3128);
nor U3287 (N_3287,N_3194,N_3157);
or U3288 (N_3288,N_3116,N_3192);
nand U3289 (N_3289,N_3180,N_3149);
or U3290 (N_3290,N_3161,N_3125);
nor U3291 (N_3291,N_3182,N_3135);
nand U3292 (N_3292,N_3130,N_3105);
nand U3293 (N_3293,N_3110,N_3181);
and U3294 (N_3294,N_3111,N_3158);
nand U3295 (N_3295,N_3199,N_3185);
nor U3296 (N_3296,N_3133,N_3140);
and U3297 (N_3297,N_3158,N_3184);
and U3298 (N_3298,N_3110,N_3172);
nor U3299 (N_3299,N_3192,N_3198);
nor U3300 (N_3300,N_3271,N_3289);
or U3301 (N_3301,N_3220,N_3205);
and U3302 (N_3302,N_3252,N_3245);
nor U3303 (N_3303,N_3284,N_3224);
xor U3304 (N_3304,N_3275,N_3261);
nor U3305 (N_3305,N_3251,N_3296);
and U3306 (N_3306,N_3223,N_3201);
or U3307 (N_3307,N_3255,N_3290);
and U3308 (N_3308,N_3202,N_3231);
and U3309 (N_3309,N_3269,N_3226);
nand U3310 (N_3310,N_3288,N_3221);
xor U3311 (N_3311,N_3265,N_3240);
or U3312 (N_3312,N_3227,N_3277);
nor U3313 (N_3313,N_3238,N_3276);
or U3314 (N_3314,N_3232,N_3279);
nand U3315 (N_3315,N_3236,N_3292);
nand U3316 (N_3316,N_3200,N_3213);
or U3317 (N_3317,N_3273,N_3299);
xnor U3318 (N_3318,N_3249,N_3264);
nor U3319 (N_3319,N_3263,N_3295);
or U3320 (N_3320,N_3243,N_3237);
nor U3321 (N_3321,N_3222,N_3297);
or U3322 (N_3322,N_3247,N_3229);
and U3323 (N_3323,N_3212,N_3286);
nand U3324 (N_3324,N_3241,N_3203);
nor U3325 (N_3325,N_3262,N_3266);
xor U3326 (N_3326,N_3294,N_3230);
or U3327 (N_3327,N_3235,N_3283);
nand U3328 (N_3328,N_3270,N_3211);
and U3329 (N_3329,N_3259,N_3228);
and U3330 (N_3330,N_3272,N_3210);
or U3331 (N_3331,N_3248,N_3257);
or U3332 (N_3332,N_3287,N_3285);
and U3333 (N_3333,N_3268,N_3282);
or U3334 (N_3334,N_3274,N_3239);
xnor U3335 (N_3335,N_3250,N_3217);
or U3336 (N_3336,N_3216,N_3209);
xor U3337 (N_3337,N_3206,N_3234);
or U3338 (N_3338,N_3258,N_3215);
or U3339 (N_3339,N_3218,N_3278);
nand U3340 (N_3340,N_3253,N_3246);
nor U3341 (N_3341,N_3256,N_3208);
or U3342 (N_3342,N_3207,N_3242);
or U3343 (N_3343,N_3293,N_3298);
nand U3344 (N_3344,N_3214,N_3280);
nand U3345 (N_3345,N_3225,N_3281);
nor U3346 (N_3346,N_3254,N_3291);
and U3347 (N_3347,N_3260,N_3204);
nand U3348 (N_3348,N_3267,N_3233);
and U3349 (N_3349,N_3219,N_3244);
nand U3350 (N_3350,N_3290,N_3280);
nand U3351 (N_3351,N_3214,N_3204);
or U3352 (N_3352,N_3223,N_3215);
and U3353 (N_3353,N_3205,N_3275);
and U3354 (N_3354,N_3206,N_3253);
nand U3355 (N_3355,N_3268,N_3249);
or U3356 (N_3356,N_3297,N_3208);
and U3357 (N_3357,N_3290,N_3218);
and U3358 (N_3358,N_3273,N_3264);
and U3359 (N_3359,N_3295,N_3212);
and U3360 (N_3360,N_3281,N_3299);
nand U3361 (N_3361,N_3214,N_3266);
and U3362 (N_3362,N_3286,N_3217);
or U3363 (N_3363,N_3213,N_3222);
or U3364 (N_3364,N_3274,N_3232);
xor U3365 (N_3365,N_3211,N_3230);
nor U3366 (N_3366,N_3292,N_3228);
and U3367 (N_3367,N_3223,N_3242);
xor U3368 (N_3368,N_3266,N_3279);
or U3369 (N_3369,N_3207,N_3226);
nand U3370 (N_3370,N_3250,N_3266);
nand U3371 (N_3371,N_3229,N_3239);
and U3372 (N_3372,N_3213,N_3294);
and U3373 (N_3373,N_3295,N_3220);
nand U3374 (N_3374,N_3205,N_3269);
and U3375 (N_3375,N_3291,N_3236);
or U3376 (N_3376,N_3287,N_3249);
nor U3377 (N_3377,N_3277,N_3256);
nor U3378 (N_3378,N_3223,N_3299);
nand U3379 (N_3379,N_3255,N_3247);
nor U3380 (N_3380,N_3298,N_3232);
and U3381 (N_3381,N_3248,N_3235);
nor U3382 (N_3382,N_3205,N_3291);
or U3383 (N_3383,N_3277,N_3239);
or U3384 (N_3384,N_3203,N_3264);
nand U3385 (N_3385,N_3285,N_3205);
and U3386 (N_3386,N_3226,N_3261);
and U3387 (N_3387,N_3290,N_3247);
or U3388 (N_3388,N_3223,N_3288);
xnor U3389 (N_3389,N_3298,N_3281);
or U3390 (N_3390,N_3286,N_3267);
or U3391 (N_3391,N_3230,N_3292);
and U3392 (N_3392,N_3200,N_3250);
nand U3393 (N_3393,N_3250,N_3242);
and U3394 (N_3394,N_3213,N_3254);
nor U3395 (N_3395,N_3261,N_3241);
or U3396 (N_3396,N_3265,N_3225);
nand U3397 (N_3397,N_3297,N_3282);
nand U3398 (N_3398,N_3217,N_3230);
xor U3399 (N_3399,N_3267,N_3287);
nand U3400 (N_3400,N_3341,N_3387);
and U3401 (N_3401,N_3395,N_3312);
or U3402 (N_3402,N_3365,N_3347);
or U3403 (N_3403,N_3376,N_3360);
or U3404 (N_3404,N_3328,N_3335);
and U3405 (N_3405,N_3397,N_3325);
xnor U3406 (N_3406,N_3350,N_3316);
or U3407 (N_3407,N_3385,N_3396);
and U3408 (N_3408,N_3363,N_3375);
nor U3409 (N_3409,N_3367,N_3300);
and U3410 (N_3410,N_3393,N_3379);
nor U3411 (N_3411,N_3369,N_3313);
nand U3412 (N_3412,N_3355,N_3326);
and U3413 (N_3413,N_3380,N_3336);
nand U3414 (N_3414,N_3329,N_3314);
and U3415 (N_3415,N_3361,N_3392);
nand U3416 (N_3416,N_3366,N_3370);
and U3417 (N_3417,N_3337,N_3389);
nand U3418 (N_3418,N_3340,N_3384);
and U3419 (N_3419,N_3318,N_3374);
nor U3420 (N_3420,N_3372,N_3399);
or U3421 (N_3421,N_3327,N_3373);
and U3422 (N_3422,N_3382,N_3331);
or U3423 (N_3423,N_3343,N_3345);
and U3424 (N_3424,N_3332,N_3352);
or U3425 (N_3425,N_3304,N_3351);
nand U3426 (N_3426,N_3319,N_3348);
and U3427 (N_3427,N_3330,N_3324);
or U3428 (N_3428,N_3323,N_3354);
and U3429 (N_3429,N_3388,N_3307);
nor U3430 (N_3430,N_3383,N_3377);
nor U3431 (N_3431,N_3386,N_3356);
xnor U3432 (N_3432,N_3305,N_3309);
nand U3433 (N_3433,N_3346,N_3315);
xnor U3434 (N_3434,N_3362,N_3378);
nor U3435 (N_3435,N_3353,N_3381);
nand U3436 (N_3436,N_3364,N_3357);
and U3437 (N_3437,N_3371,N_3339);
or U3438 (N_3438,N_3391,N_3349);
and U3439 (N_3439,N_3302,N_3306);
xnor U3440 (N_3440,N_3359,N_3333);
and U3441 (N_3441,N_3368,N_3358);
and U3442 (N_3442,N_3390,N_3301);
nor U3443 (N_3443,N_3322,N_3303);
nand U3444 (N_3444,N_3398,N_3317);
or U3445 (N_3445,N_3344,N_3311);
nor U3446 (N_3446,N_3310,N_3394);
xnor U3447 (N_3447,N_3338,N_3321);
or U3448 (N_3448,N_3342,N_3308);
nor U3449 (N_3449,N_3320,N_3334);
nor U3450 (N_3450,N_3304,N_3341);
xnor U3451 (N_3451,N_3373,N_3311);
or U3452 (N_3452,N_3393,N_3377);
and U3453 (N_3453,N_3346,N_3386);
nand U3454 (N_3454,N_3364,N_3362);
nand U3455 (N_3455,N_3308,N_3335);
nand U3456 (N_3456,N_3327,N_3344);
nand U3457 (N_3457,N_3378,N_3352);
and U3458 (N_3458,N_3360,N_3353);
nor U3459 (N_3459,N_3334,N_3390);
and U3460 (N_3460,N_3313,N_3316);
and U3461 (N_3461,N_3328,N_3375);
nand U3462 (N_3462,N_3368,N_3332);
nand U3463 (N_3463,N_3328,N_3393);
nand U3464 (N_3464,N_3300,N_3371);
or U3465 (N_3465,N_3399,N_3379);
or U3466 (N_3466,N_3383,N_3399);
nor U3467 (N_3467,N_3385,N_3317);
nor U3468 (N_3468,N_3328,N_3313);
or U3469 (N_3469,N_3380,N_3375);
and U3470 (N_3470,N_3390,N_3367);
and U3471 (N_3471,N_3377,N_3318);
and U3472 (N_3472,N_3331,N_3348);
or U3473 (N_3473,N_3387,N_3303);
nand U3474 (N_3474,N_3372,N_3322);
and U3475 (N_3475,N_3353,N_3312);
or U3476 (N_3476,N_3382,N_3396);
and U3477 (N_3477,N_3323,N_3394);
nand U3478 (N_3478,N_3334,N_3337);
or U3479 (N_3479,N_3326,N_3387);
and U3480 (N_3480,N_3311,N_3304);
nand U3481 (N_3481,N_3327,N_3332);
or U3482 (N_3482,N_3383,N_3396);
or U3483 (N_3483,N_3372,N_3358);
nand U3484 (N_3484,N_3345,N_3389);
and U3485 (N_3485,N_3341,N_3394);
or U3486 (N_3486,N_3316,N_3302);
or U3487 (N_3487,N_3319,N_3328);
or U3488 (N_3488,N_3391,N_3388);
xnor U3489 (N_3489,N_3305,N_3313);
and U3490 (N_3490,N_3397,N_3380);
nand U3491 (N_3491,N_3348,N_3386);
nand U3492 (N_3492,N_3378,N_3310);
and U3493 (N_3493,N_3340,N_3389);
and U3494 (N_3494,N_3315,N_3352);
or U3495 (N_3495,N_3302,N_3349);
nor U3496 (N_3496,N_3333,N_3344);
or U3497 (N_3497,N_3393,N_3363);
or U3498 (N_3498,N_3330,N_3398);
nor U3499 (N_3499,N_3365,N_3326);
nand U3500 (N_3500,N_3476,N_3442);
or U3501 (N_3501,N_3474,N_3447);
nand U3502 (N_3502,N_3415,N_3446);
nor U3503 (N_3503,N_3427,N_3429);
or U3504 (N_3504,N_3469,N_3481);
or U3505 (N_3505,N_3484,N_3457);
and U3506 (N_3506,N_3406,N_3443);
nor U3507 (N_3507,N_3438,N_3471);
nor U3508 (N_3508,N_3467,N_3436);
nand U3509 (N_3509,N_3489,N_3488);
and U3510 (N_3510,N_3405,N_3465);
nand U3511 (N_3511,N_3459,N_3485);
and U3512 (N_3512,N_3463,N_3437);
nor U3513 (N_3513,N_3497,N_3490);
nand U3514 (N_3514,N_3466,N_3448);
or U3515 (N_3515,N_3409,N_3453);
nor U3516 (N_3516,N_3482,N_3462);
or U3517 (N_3517,N_3424,N_3495);
nand U3518 (N_3518,N_3426,N_3483);
nand U3519 (N_3519,N_3445,N_3428);
and U3520 (N_3520,N_3475,N_3449);
nor U3521 (N_3521,N_3477,N_3499);
nand U3522 (N_3522,N_3458,N_3423);
nand U3523 (N_3523,N_3425,N_3473);
nor U3524 (N_3524,N_3404,N_3400);
and U3525 (N_3525,N_3472,N_3444);
nor U3526 (N_3526,N_3410,N_3419);
and U3527 (N_3527,N_3416,N_3480);
and U3528 (N_3528,N_3408,N_3487);
nor U3529 (N_3529,N_3479,N_3454);
nand U3530 (N_3530,N_3493,N_3403);
and U3531 (N_3531,N_3464,N_3422);
nor U3532 (N_3532,N_3434,N_3468);
nor U3533 (N_3533,N_3432,N_3413);
nand U3534 (N_3534,N_3402,N_3492);
or U3535 (N_3535,N_3418,N_3421);
and U3536 (N_3536,N_3430,N_3452);
or U3537 (N_3537,N_3417,N_3433);
and U3538 (N_3538,N_3439,N_3401);
nor U3539 (N_3539,N_3412,N_3407);
and U3540 (N_3540,N_3451,N_3440);
and U3541 (N_3541,N_3491,N_3494);
xnor U3542 (N_3542,N_3486,N_3456);
nand U3543 (N_3543,N_3498,N_3431);
or U3544 (N_3544,N_3460,N_3441);
xor U3545 (N_3545,N_3478,N_3435);
or U3546 (N_3546,N_3455,N_3461);
and U3547 (N_3547,N_3411,N_3420);
nand U3548 (N_3548,N_3450,N_3470);
nand U3549 (N_3549,N_3414,N_3496);
nand U3550 (N_3550,N_3448,N_3419);
or U3551 (N_3551,N_3443,N_3427);
and U3552 (N_3552,N_3469,N_3445);
and U3553 (N_3553,N_3445,N_3435);
nor U3554 (N_3554,N_3497,N_3469);
nand U3555 (N_3555,N_3469,N_3496);
xnor U3556 (N_3556,N_3464,N_3480);
nand U3557 (N_3557,N_3404,N_3494);
nand U3558 (N_3558,N_3439,N_3418);
nand U3559 (N_3559,N_3462,N_3475);
nand U3560 (N_3560,N_3415,N_3454);
or U3561 (N_3561,N_3432,N_3410);
xor U3562 (N_3562,N_3466,N_3493);
nand U3563 (N_3563,N_3485,N_3481);
nor U3564 (N_3564,N_3497,N_3495);
nor U3565 (N_3565,N_3402,N_3474);
nor U3566 (N_3566,N_3453,N_3458);
nand U3567 (N_3567,N_3461,N_3495);
nand U3568 (N_3568,N_3479,N_3417);
nor U3569 (N_3569,N_3420,N_3402);
nor U3570 (N_3570,N_3470,N_3459);
or U3571 (N_3571,N_3432,N_3457);
nand U3572 (N_3572,N_3481,N_3470);
nor U3573 (N_3573,N_3411,N_3477);
or U3574 (N_3574,N_3471,N_3441);
and U3575 (N_3575,N_3450,N_3433);
or U3576 (N_3576,N_3408,N_3497);
nand U3577 (N_3577,N_3411,N_3422);
nor U3578 (N_3578,N_3413,N_3438);
xnor U3579 (N_3579,N_3466,N_3415);
and U3580 (N_3580,N_3457,N_3460);
nand U3581 (N_3581,N_3474,N_3488);
xor U3582 (N_3582,N_3490,N_3402);
nand U3583 (N_3583,N_3461,N_3403);
or U3584 (N_3584,N_3451,N_3405);
nand U3585 (N_3585,N_3455,N_3437);
and U3586 (N_3586,N_3405,N_3422);
nor U3587 (N_3587,N_3412,N_3468);
and U3588 (N_3588,N_3447,N_3486);
nand U3589 (N_3589,N_3473,N_3433);
nand U3590 (N_3590,N_3473,N_3456);
nor U3591 (N_3591,N_3463,N_3474);
or U3592 (N_3592,N_3408,N_3453);
and U3593 (N_3593,N_3477,N_3487);
nand U3594 (N_3594,N_3438,N_3420);
nand U3595 (N_3595,N_3417,N_3421);
nor U3596 (N_3596,N_3457,N_3420);
nor U3597 (N_3597,N_3429,N_3470);
nor U3598 (N_3598,N_3449,N_3484);
nor U3599 (N_3599,N_3406,N_3473);
nand U3600 (N_3600,N_3589,N_3538);
xor U3601 (N_3601,N_3556,N_3505);
xnor U3602 (N_3602,N_3516,N_3528);
nand U3603 (N_3603,N_3583,N_3558);
nor U3604 (N_3604,N_3551,N_3517);
nor U3605 (N_3605,N_3501,N_3552);
xor U3606 (N_3606,N_3567,N_3550);
and U3607 (N_3607,N_3593,N_3579);
xnor U3608 (N_3608,N_3563,N_3568);
and U3609 (N_3609,N_3539,N_3561);
xnor U3610 (N_3610,N_3519,N_3584);
nand U3611 (N_3611,N_3590,N_3592);
or U3612 (N_3612,N_3520,N_3504);
nand U3613 (N_3613,N_3506,N_3597);
and U3614 (N_3614,N_3525,N_3581);
nand U3615 (N_3615,N_3596,N_3565);
or U3616 (N_3616,N_3523,N_3549);
and U3617 (N_3617,N_3503,N_3573);
or U3618 (N_3618,N_3514,N_3532);
nand U3619 (N_3619,N_3502,N_3559);
nor U3620 (N_3620,N_3513,N_3598);
or U3621 (N_3621,N_3570,N_3574);
nand U3622 (N_3622,N_3533,N_3543);
or U3623 (N_3623,N_3591,N_3531);
nor U3624 (N_3624,N_3569,N_3509);
or U3625 (N_3625,N_3511,N_3535);
and U3626 (N_3626,N_3580,N_3546);
nor U3627 (N_3627,N_3544,N_3545);
and U3628 (N_3628,N_3577,N_3541);
nand U3629 (N_3629,N_3529,N_3526);
nor U3630 (N_3630,N_3547,N_3508);
and U3631 (N_3631,N_3571,N_3534);
nand U3632 (N_3632,N_3527,N_3522);
nor U3633 (N_3633,N_3518,N_3557);
nor U3634 (N_3634,N_3566,N_3515);
nor U3635 (N_3635,N_3536,N_3530);
and U3636 (N_3636,N_3512,N_3572);
or U3637 (N_3637,N_3540,N_3585);
nand U3638 (N_3638,N_3587,N_3500);
and U3639 (N_3639,N_3548,N_3553);
xnor U3640 (N_3640,N_3554,N_3576);
and U3641 (N_3641,N_3595,N_3562);
or U3642 (N_3642,N_3582,N_3524);
or U3643 (N_3643,N_3560,N_3510);
xor U3644 (N_3644,N_3507,N_3594);
nor U3645 (N_3645,N_3555,N_3599);
or U3646 (N_3646,N_3586,N_3537);
xnor U3647 (N_3647,N_3564,N_3588);
and U3648 (N_3648,N_3521,N_3542);
or U3649 (N_3649,N_3578,N_3575);
nand U3650 (N_3650,N_3588,N_3599);
nand U3651 (N_3651,N_3502,N_3588);
nand U3652 (N_3652,N_3599,N_3574);
and U3653 (N_3653,N_3572,N_3502);
xor U3654 (N_3654,N_3507,N_3540);
xnor U3655 (N_3655,N_3566,N_3557);
and U3656 (N_3656,N_3561,N_3502);
nand U3657 (N_3657,N_3518,N_3532);
nand U3658 (N_3658,N_3568,N_3536);
nand U3659 (N_3659,N_3593,N_3551);
nor U3660 (N_3660,N_3519,N_3555);
and U3661 (N_3661,N_3525,N_3593);
nor U3662 (N_3662,N_3567,N_3575);
or U3663 (N_3663,N_3539,N_3574);
nand U3664 (N_3664,N_3517,N_3560);
or U3665 (N_3665,N_3519,N_3530);
nand U3666 (N_3666,N_3532,N_3580);
and U3667 (N_3667,N_3509,N_3528);
nand U3668 (N_3668,N_3596,N_3585);
nand U3669 (N_3669,N_3576,N_3555);
or U3670 (N_3670,N_3507,N_3549);
or U3671 (N_3671,N_3579,N_3573);
xor U3672 (N_3672,N_3550,N_3579);
nand U3673 (N_3673,N_3505,N_3580);
nand U3674 (N_3674,N_3528,N_3594);
nor U3675 (N_3675,N_3539,N_3541);
nand U3676 (N_3676,N_3526,N_3508);
or U3677 (N_3677,N_3542,N_3548);
and U3678 (N_3678,N_3575,N_3512);
or U3679 (N_3679,N_3593,N_3519);
nor U3680 (N_3680,N_3520,N_3573);
nand U3681 (N_3681,N_3517,N_3574);
nand U3682 (N_3682,N_3544,N_3580);
or U3683 (N_3683,N_3540,N_3554);
or U3684 (N_3684,N_3584,N_3596);
and U3685 (N_3685,N_3544,N_3589);
and U3686 (N_3686,N_3597,N_3569);
xnor U3687 (N_3687,N_3525,N_3567);
or U3688 (N_3688,N_3543,N_3522);
and U3689 (N_3689,N_3583,N_3541);
nand U3690 (N_3690,N_3546,N_3530);
or U3691 (N_3691,N_3581,N_3560);
nand U3692 (N_3692,N_3546,N_3517);
and U3693 (N_3693,N_3537,N_3514);
and U3694 (N_3694,N_3568,N_3552);
nor U3695 (N_3695,N_3575,N_3598);
or U3696 (N_3696,N_3502,N_3509);
nor U3697 (N_3697,N_3538,N_3508);
xnor U3698 (N_3698,N_3501,N_3571);
xor U3699 (N_3699,N_3511,N_3562);
and U3700 (N_3700,N_3693,N_3623);
and U3701 (N_3701,N_3682,N_3639);
or U3702 (N_3702,N_3626,N_3619);
xnor U3703 (N_3703,N_3646,N_3667);
nand U3704 (N_3704,N_3630,N_3676);
or U3705 (N_3705,N_3681,N_3645);
nor U3706 (N_3706,N_3652,N_3612);
nor U3707 (N_3707,N_3662,N_3611);
nor U3708 (N_3708,N_3698,N_3608);
and U3709 (N_3709,N_3643,N_3697);
nand U3710 (N_3710,N_3624,N_3672);
nand U3711 (N_3711,N_3655,N_3658);
nand U3712 (N_3712,N_3636,N_3678);
nand U3713 (N_3713,N_3673,N_3691);
nor U3714 (N_3714,N_3677,N_3651);
or U3715 (N_3715,N_3654,N_3625);
or U3716 (N_3716,N_3695,N_3670);
nand U3717 (N_3717,N_3656,N_3661);
nand U3718 (N_3718,N_3650,N_3627);
or U3719 (N_3719,N_3694,N_3688);
or U3720 (N_3720,N_3660,N_3601);
and U3721 (N_3721,N_3692,N_3629);
or U3722 (N_3722,N_3615,N_3634);
and U3723 (N_3723,N_3685,N_3640);
and U3724 (N_3724,N_3603,N_3657);
or U3725 (N_3725,N_3613,N_3617);
or U3726 (N_3726,N_3664,N_3642);
nor U3727 (N_3727,N_3637,N_3609);
nor U3728 (N_3728,N_3659,N_3631);
nand U3729 (N_3729,N_3605,N_3638);
nor U3730 (N_3730,N_3665,N_3618);
and U3731 (N_3731,N_3690,N_3616);
xor U3732 (N_3732,N_3696,N_3680);
and U3733 (N_3733,N_3632,N_3628);
or U3734 (N_3734,N_3666,N_3699);
or U3735 (N_3735,N_3621,N_3648);
or U3736 (N_3736,N_3641,N_3683);
nor U3737 (N_3737,N_3644,N_3610);
nor U3738 (N_3738,N_3620,N_3679);
nand U3739 (N_3739,N_3669,N_3602);
xor U3740 (N_3740,N_3686,N_3668);
or U3741 (N_3741,N_3675,N_3604);
xor U3742 (N_3742,N_3647,N_3614);
nor U3743 (N_3743,N_3622,N_3663);
xor U3744 (N_3744,N_3689,N_3606);
nand U3745 (N_3745,N_3633,N_3674);
xnor U3746 (N_3746,N_3653,N_3684);
or U3747 (N_3747,N_3600,N_3687);
nor U3748 (N_3748,N_3607,N_3649);
or U3749 (N_3749,N_3635,N_3671);
nand U3750 (N_3750,N_3653,N_3647);
and U3751 (N_3751,N_3661,N_3633);
nand U3752 (N_3752,N_3609,N_3602);
and U3753 (N_3753,N_3624,N_3648);
nand U3754 (N_3754,N_3690,N_3645);
nand U3755 (N_3755,N_3669,N_3690);
nor U3756 (N_3756,N_3688,N_3682);
nand U3757 (N_3757,N_3654,N_3634);
or U3758 (N_3758,N_3611,N_3652);
nand U3759 (N_3759,N_3644,N_3678);
and U3760 (N_3760,N_3674,N_3670);
nor U3761 (N_3761,N_3620,N_3631);
and U3762 (N_3762,N_3613,N_3659);
xor U3763 (N_3763,N_3602,N_3664);
and U3764 (N_3764,N_3654,N_3633);
and U3765 (N_3765,N_3654,N_3646);
nand U3766 (N_3766,N_3600,N_3686);
nand U3767 (N_3767,N_3616,N_3661);
nor U3768 (N_3768,N_3675,N_3627);
and U3769 (N_3769,N_3666,N_3603);
nor U3770 (N_3770,N_3624,N_3649);
and U3771 (N_3771,N_3677,N_3682);
nand U3772 (N_3772,N_3643,N_3656);
nor U3773 (N_3773,N_3618,N_3699);
or U3774 (N_3774,N_3676,N_3666);
or U3775 (N_3775,N_3670,N_3696);
nand U3776 (N_3776,N_3682,N_3692);
nand U3777 (N_3777,N_3674,N_3616);
nand U3778 (N_3778,N_3687,N_3692);
and U3779 (N_3779,N_3649,N_3680);
and U3780 (N_3780,N_3669,N_3647);
or U3781 (N_3781,N_3667,N_3680);
or U3782 (N_3782,N_3605,N_3627);
and U3783 (N_3783,N_3676,N_3631);
or U3784 (N_3784,N_3651,N_3618);
xnor U3785 (N_3785,N_3645,N_3696);
and U3786 (N_3786,N_3656,N_3653);
and U3787 (N_3787,N_3622,N_3671);
xor U3788 (N_3788,N_3688,N_3647);
or U3789 (N_3789,N_3696,N_3618);
and U3790 (N_3790,N_3679,N_3678);
nor U3791 (N_3791,N_3685,N_3676);
or U3792 (N_3792,N_3671,N_3658);
xnor U3793 (N_3793,N_3658,N_3694);
or U3794 (N_3794,N_3693,N_3609);
nand U3795 (N_3795,N_3676,N_3680);
xnor U3796 (N_3796,N_3650,N_3655);
and U3797 (N_3797,N_3604,N_3642);
xor U3798 (N_3798,N_3619,N_3635);
or U3799 (N_3799,N_3632,N_3630);
nor U3800 (N_3800,N_3786,N_3751);
nand U3801 (N_3801,N_3706,N_3796);
nand U3802 (N_3802,N_3754,N_3799);
xor U3803 (N_3803,N_3716,N_3730);
nand U3804 (N_3804,N_3776,N_3791);
nor U3805 (N_3805,N_3768,N_3752);
nand U3806 (N_3806,N_3766,N_3753);
and U3807 (N_3807,N_3794,N_3729);
or U3808 (N_3808,N_3763,N_3719);
or U3809 (N_3809,N_3780,N_3724);
xnor U3810 (N_3810,N_3737,N_3772);
or U3811 (N_3811,N_3721,N_3784);
or U3812 (N_3812,N_3762,N_3727);
and U3813 (N_3813,N_3707,N_3733);
nand U3814 (N_3814,N_3702,N_3755);
and U3815 (N_3815,N_3769,N_3718);
nor U3816 (N_3816,N_3735,N_3742);
nor U3817 (N_3817,N_3723,N_3795);
nor U3818 (N_3818,N_3748,N_3728);
or U3819 (N_3819,N_3725,N_3777);
nor U3820 (N_3820,N_3720,N_3767);
and U3821 (N_3821,N_3739,N_3743);
or U3822 (N_3822,N_3787,N_3788);
nor U3823 (N_3823,N_3793,N_3722);
nor U3824 (N_3824,N_3759,N_3798);
and U3825 (N_3825,N_3709,N_3781);
or U3826 (N_3826,N_3783,N_3792);
nand U3827 (N_3827,N_3703,N_3711);
nor U3828 (N_3828,N_3770,N_3764);
or U3829 (N_3829,N_3771,N_3785);
nor U3830 (N_3830,N_3744,N_3705);
nand U3831 (N_3831,N_3741,N_3778);
nor U3832 (N_3832,N_3761,N_3715);
and U3833 (N_3833,N_3782,N_3738);
xor U3834 (N_3834,N_3745,N_3717);
xnor U3835 (N_3835,N_3736,N_3731);
nand U3836 (N_3836,N_3779,N_3700);
nor U3837 (N_3837,N_3701,N_3732);
nand U3838 (N_3838,N_3756,N_3797);
nor U3839 (N_3839,N_3746,N_3708);
nand U3840 (N_3840,N_3749,N_3775);
or U3841 (N_3841,N_3774,N_3773);
nand U3842 (N_3842,N_3710,N_3750);
and U3843 (N_3843,N_3758,N_3765);
and U3844 (N_3844,N_3760,N_3740);
nand U3845 (N_3845,N_3713,N_3790);
nand U3846 (N_3846,N_3734,N_3757);
or U3847 (N_3847,N_3712,N_3714);
nor U3848 (N_3848,N_3726,N_3747);
nand U3849 (N_3849,N_3789,N_3704);
and U3850 (N_3850,N_3776,N_3734);
xnor U3851 (N_3851,N_3740,N_3705);
xor U3852 (N_3852,N_3746,N_3777);
nand U3853 (N_3853,N_3769,N_3724);
nor U3854 (N_3854,N_3705,N_3777);
and U3855 (N_3855,N_3798,N_3774);
nor U3856 (N_3856,N_3708,N_3738);
and U3857 (N_3857,N_3798,N_3796);
xnor U3858 (N_3858,N_3758,N_3706);
nand U3859 (N_3859,N_3793,N_3773);
nor U3860 (N_3860,N_3797,N_3776);
nand U3861 (N_3861,N_3792,N_3751);
and U3862 (N_3862,N_3732,N_3753);
xor U3863 (N_3863,N_3764,N_3700);
or U3864 (N_3864,N_3756,N_3700);
or U3865 (N_3865,N_3783,N_3795);
and U3866 (N_3866,N_3708,N_3782);
and U3867 (N_3867,N_3727,N_3786);
nand U3868 (N_3868,N_3789,N_3726);
nand U3869 (N_3869,N_3733,N_3732);
or U3870 (N_3870,N_3785,N_3705);
or U3871 (N_3871,N_3741,N_3751);
or U3872 (N_3872,N_3779,N_3702);
and U3873 (N_3873,N_3734,N_3723);
and U3874 (N_3874,N_3771,N_3788);
and U3875 (N_3875,N_3738,N_3703);
and U3876 (N_3876,N_3754,N_3760);
nor U3877 (N_3877,N_3734,N_3788);
nor U3878 (N_3878,N_3739,N_3760);
or U3879 (N_3879,N_3747,N_3737);
and U3880 (N_3880,N_3790,N_3734);
nand U3881 (N_3881,N_3729,N_3730);
nand U3882 (N_3882,N_3798,N_3752);
xor U3883 (N_3883,N_3787,N_3738);
and U3884 (N_3884,N_3716,N_3765);
and U3885 (N_3885,N_3759,N_3715);
and U3886 (N_3886,N_3745,N_3775);
or U3887 (N_3887,N_3700,N_3743);
or U3888 (N_3888,N_3747,N_3788);
xor U3889 (N_3889,N_3792,N_3756);
or U3890 (N_3890,N_3752,N_3797);
nor U3891 (N_3891,N_3786,N_3764);
nor U3892 (N_3892,N_3745,N_3781);
nor U3893 (N_3893,N_3783,N_3718);
nand U3894 (N_3894,N_3736,N_3783);
nor U3895 (N_3895,N_3758,N_3792);
nor U3896 (N_3896,N_3712,N_3720);
nand U3897 (N_3897,N_3724,N_3742);
nor U3898 (N_3898,N_3719,N_3723);
and U3899 (N_3899,N_3744,N_3781);
or U3900 (N_3900,N_3872,N_3889);
or U3901 (N_3901,N_3880,N_3881);
or U3902 (N_3902,N_3847,N_3812);
nor U3903 (N_3903,N_3800,N_3840);
nand U3904 (N_3904,N_3876,N_3879);
xnor U3905 (N_3905,N_3838,N_3875);
and U3906 (N_3906,N_3882,N_3888);
nand U3907 (N_3907,N_3824,N_3844);
and U3908 (N_3908,N_3825,N_3828);
or U3909 (N_3909,N_3821,N_3829);
or U3910 (N_3910,N_3865,N_3868);
nand U3911 (N_3911,N_3891,N_3867);
nand U3912 (N_3912,N_3805,N_3848);
nand U3913 (N_3913,N_3851,N_3898);
nand U3914 (N_3914,N_3818,N_3813);
xor U3915 (N_3915,N_3853,N_3859);
nand U3916 (N_3916,N_3832,N_3820);
nor U3917 (N_3917,N_3827,N_3811);
nor U3918 (N_3918,N_3819,N_3895);
and U3919 (N_3919,N_3877,N_3855);
xor U3920 (N_3920,N_3830,N_3816);
xnor U3921 (N_3921,N_3841,N_3804);
nor U3922 (N_3922,N_3849,N_3822);
nor U3923 (N_3923,N_3864,N_3837);
nand U3924 (N_3924,N_3870,N_3897);
xnor U3925 (N_3925,N_3843,N_3863);
and U3926 (N_3926,N_3842,N_3831);
nand U3927 (N_3927,N_3846,N_3886);
xnor U3928 (N_3928,N_3893,N_3806);
and U3929 (N_3929,N_3807,N_3833);
xor U3930 (N_3930,N_3861,N_3808);
xor U3931 (N_3931,N_3852,N_3860);
or U3932 (N_3932,N_3823,N_3878);
and U3933 (N_3933,N_3885,N_3826);
or U3934 (N_3934,N_3845,N_3856);
nor U3935 (N_3935,N_3809,N_3802);
nand U3936 (N_3936,N_3892,N_3896);
nor U3937 (N_3937,N_3858,N_3871);
nand U3938 (N_3938,N_3894,N_3884);
and U3939 (N_3939,N_3873,N_3850);
or U3940 (N_3940,N_3869,N_3883);
xor U3941 (N_3941,N_3814,N_3899);
or U3942 (N_3942,N_3835,N_3887);
nand U3943 (N_3943,N_3834,N_3890);
nor U3944 (N_3944,N_3854,N_3839);
or U3945 (N_3945,N_3810,N_3801);
and U3946 (N_3946,N_3874,N_3803);
or U3947 (N_3947,N_3817,N_3862);
and U3948 (N_3948,N_3857,N_3836);
and U3949 (N_3949,N_3866,N_3815);
nand U3950 (N_3950,N_3858,N_3801);
nand U3951 (N_3951,N_3856,N_3830);
xnor U3952 (N_3952,N_3830,N_3823);
nand U3953 (N_3953,N_3851,N_3873);
nor U3954 (N_3954,N_3860,N_3869);
nand U3955 (N_3955,N_3857,N_3889);
xor U3956 (N_3956,N_3873,N_3848);
or U3957 (N_3957,N_3891,N_3810);
or U3958 (N_3958,N_3820,N_3895);
nor U3959 (N_3959,N_3883,N_3864);
or U3960 (N_3960,N_3824,N_3854);
and U3961 (N_3961,N_3855,N_3867);
nor U3962 (N_3962,N_3854,N_3882);
nor U3963 (N_3963,N_3815,N_3860);
nand U3964 (N_3964,N_3868,N_3898);
or U3965 (N_3965,N_3890,N_3852);
or U3966 (N_3966,N_3809,N_3815);
nor U3967 (N_3967,N_3877,N_3850);
nand U3968 (N_3968,N_3883,N_3822);
and U3969 (N_3969,N_3892,N_3829);
or U3970 (N_3970,N_3853,N_3860);
nand U3971 (N_3971,N_3800,N_3851);
nor U3972 (N_3972,N_3845,N_3802);
and U3973 (N_3973,N_3841,N_3851);
nand U3974 (N_3974,N_3805,N_3835);
or U3975 (N_3975,N_3827,N_3887);
nor U3976 (N_3976,N_3834,N_3809);
nand U3977 (N_3977,N_3826,N_3868);
or U3978 (N_3978,N_3822,N_3874);
and U3979 (N_3979,N_3879,N_3889);
and U3980 (N_3980,N_3836,N_3844);
and U3981 (N_3981,N_3857,N_3831);
or U3982 (N_3982,N_3805,N_3872);
nor U3983 (N_3983,N_3879,N_3859);
nor U3984 (N_3984,N_3812,N_3895);
and U3985 (N_3985,N_3858,N_3890);
nor U3986 (N_3986,N_3879,N_3887);
nand U3987 (N_3987,N_3866,N_3897);
nor U3988 (N_3988,N_3832,N_3843);
nand U3989 (N_3989,N_3896,N_3865);
and U3990 (N_3990,N_3896,N_3897);
xnor U3991 (N_3991,N_3804,N_3802);
and U3992 (N_3992,N_3869,N_3888);
nor U3993 (N_3993,N_3895,N_3896);
nor U3994 (N_3994,N_3886,N_3816);
xor U3995 (N_3995,N_3867,N_3822);
nand U3996 (N_3996,N_3841,N_3852);
nor U3997 (N_3997,N_3850,N_3810);
or U3998 (N_3998,N_3858,N_3808);
and U3999 (N_3999,N_3839,N_3825);
or U4000 (N_4000,N_3913,N_3907);
and U4001 (N_4001,N_3979,N_3936);
xnor U4002 (N_4002,N_3947,N_3966);
nor U4003 (N_4003,N_3943,N_3935);
or U4004 (N_4004,N_3965,N_3909);
or U4005 (N_4005,N_3993,N_3949);
or U4006 (N_4006,N_3985,N_3989);
or U4007 (N_4007,N_3967,N_3924);
and U4008 (N_4008,N_3970,N_3923);
or U4009 (N_4009,N_3946,N_3964);
nand U4010 (N_4010,N_3975,N_3968);
or U4011 (N_4011,N_3982,N_3981);
nand U4012 (N_4012,N_3916,N_3906);
nor U4013 (N_4013,N_3958,N_3944);
nand U4014 (N_4014,N_3976,N_3918);
nor U4015 (N_4015,N_3977,N_3917);
nand U4016 (N_4016,N_3998,N_3956);
or U4017 (N_4017,N_3940,N_3900);
or U4018 (N_4018,N_3983,N_3990);
and U4019 (N_4019,N_3997,N_3905);
nand U4020 (N_4020,N_3933,N_3915);
nor U4021 (N_4021,N_3992,N_3962);
or U4022 (N_4022,N_3929,N_3926);
or U4023 (N_4023,N_3922,N_3930);
nand U4024 (N_4024,N_3996,N_3954);
nand U4025 (N_4025,N_3972,N_3948);
and U4026 (N_4026,N_3974,N_3960);
nand U4027 (N_4027,N_3901,N_3932);
and U4028 (N_4028,N_3927,N_3921);
nand U4029 (N_4029,N_3904,N_3908);
and U4030 (N_4030,N_3910,N_3984);
nor U4031 (N_4031,N_3971,N_3912);
nand U4032 (N_4032,N_3914,N_3978);
nand U4033 (N_4033,N_3991,N_3955);
nor U4034 (N_4034,N_3920,N_3903);
or U4035 (N_4035,N_3973,N_3951);
or U4036 (N_4036,N_3995,N_3953);
and U4037 (N_4037,N_3931,N_3945);
xor U4038 (N_4038,N_3952,N_3986);
and U4039 (N_4039,N_3988,N_3994);
or U4040 (N_4040,N_3937,N_3999);
nand U4041 (N_4041,N_3987,N_3928);
or U4042 (N_4042,N_3980,N_3950);
nand U4043 (N_4043,N_3963,N_3961);
xnor U4044 (N_4044,N_3957,N_3959);
and U4045 (N_4045,N_3919,N_3939);
nand U4046 (N_4046,N_3969,N_3934);
nand U4047 (N_4047,N_3911,N_3941);
xnor U4048 (N_4048,N_3925,N_3938);
xnor U4049 (N_4049,N_3942,N_3902);
nand U4050 (N_4050,N_3927,N_3962);
nor U4051 (N_4051,N_3985,N_3959);
and U4052 (N_4052,N_3946,N_3945);
or U4053 (N_4053,N_3989,N_3945);
nand U4054 (N_4054,N_3956,N_3918);
and U4055 (N_4055,N_3979,N_3956);
and U4056 (N_4056,N_3965,N_3961);
or U4057 (N_4057,N_3908,N_3944);
and U4058 (N_4058,N_3971,N_3905);
or U4059 (N_4059,N_3992,N_3948);
nand U4060 (N_4060,N_3977,N_3959);
and U4061 (N_4061,N_3926,N_3937);
nand U4062 (N_4062,N_3976,N_3929);
or U4063 (N_4063,N_3941,N_3971);
nor U4064 (N_4064,N_3945,N_3910);
or U4065 (N_4065,N_3969,N_3960);
xnor U4066 (N_4066,N_3910,N_3931);
nand U4067 (N_4067,N_3919,N_3950);
and U4068 (N_4068,N_3916,N_3921);
xor U4069 (N_4069,N_3940,N_3996);
nor U4070 (N_4070,N_3962,N_3933);
nor U4071 (N_4071,N_3933,N_3981);
nor U4072 (N_4072,N_3973,N_3955);
nand U4073 (N_4073,N_3919,N_3918);
or U4074 (N_4074,N_3980,N_3970);
xor U4075 (N_4075,N_3910,N_3959);
nor U4076 (N_4076,N_3994,N_3953);
or U4077 (N_4077,N_3975,N_3929);
and U4078 (N_4078,N_3907,N_3922);
or U4079 (N_4079,N_3986,N_3901);
xnor U4080 (N_4080,N_3919,N_3977);
or U4081 (N_4081,N_3967,N_3939);
nor U4082 (N_4082,N_3917,N_3919);
nor U4083 (N_4083,N_3984,N_3952);
and U4084 (N_4084,N_3950,N_3956);
nand U4085 (N_4085,N_3917,N_3992);
nor U4086 (N_4086,N_3915,N_3978);
and U4087 (N_4087,N_3998,N_3983);
nor U4088 (N_4088,N_3924,N_3922);
or U4089 (N_4089,N_3915,N_3922);
nand U4090 (N_4090,N_3966,N_3910);
nand U4091 (N_4091,N_3964,N_3994);
or U4092 (N_4092,N_3954,N_3998);
or U4093 (N_4093,N_3900,N_3976);
or U4094 (N_4094,N_3917,N_3995);
nor U4095 (N_4095,N_3921,N_3908);
nor U4096 (N_4096,N_3931,N_3976);
and U4097 (N_4097,N_3908,N_3911);
and U4098 (N_4098,N_3942,N_3960);
nor U4099 (N_4099,N_3941,N_3910);
or U4100 (N_4100,N_4003,N_4046);
nand U4101 (N_4101,N_4041,N_4033);
or U4102 (N_4102,N_4066,N_4077);
and U4103 (N_4103,N_4055,N_4071);
nand U4104 (N_4104,N_4024,N_4097);
or U4105 (N_4105,N_4064,N_4009);
nor U4106 (N_4106,N_4095,N_4062);
xor U4107 (N_4107,N_4065,N_4023);
and U4108 (N_4108,N_4015,N_4019);
and U4109 (N_4109,N_4021,N_4070);
nor U4110 (N_4110,N_4083,N_4049);
nand U4111 (N_4111,N_4048,N_4027);
and U4112 (N_4112,N_4000,N_4005);
and U4113 (N_4113,N_4044,N_4073);
and U4114 (N_4114,N_4022,N_4004);
nand U4115 (N_4115,N_4031,N_4084);
or U4116 (N_4116,N_4085,N_4008);
or U4117 (N_4117,N_4030,N_4012);
and U4118 (N_4118,N_4075,N_4050);
nor U4119 (N_4119,N_4092,N_4053);
nor U4120 (N_4120,N_4091,N_4052);
and U4121 (N_4121,N_4036,N_4068);
xor U4122 (N_4122,N_4032,N_4054);
nand U4123 (N_4123,N_4020,N_4026);
and U4124 (N_4124,N_4002,N_4017);
or U4125 (N_4125,N_4072,N_4038);
nor U4126 (N_4126,N_4094,N_4011);
and U4127 (N_4127,N_4063,N_4013);
nand U4128 (N_4128,N_4001,N_4018);
or U4129 (N_4129,N_4059,N_4057);
or U4130 (N_4130,N_4007,N_4074);
xnor U4131 (N_4131,N_4016,N_4076);
xor U4132 (N_4132,N_4087,N_4037);
or U4133 (N_4133,N_4058,N_4069);
nand U4134 (N_4134,N_4088,N_4034);
or U4135 (N_4135,N_4060,N_4079);
or U4136 (N_4136,N_4093,N_4067);
and U4137 (N_4137,N_4086,N_4098);
or U4138 (N_4138,N_4090,N_4025);
or U4139 (N_4139,N_4061,N_4056);
nor U4140 (N_4140,N_4089,N_4081);
nand U4141 (N_4141,N_4082,N_4006);
nor U4142 (N_4142,N_4096,N_4078);
or U4143 (N_4143,N_4045,N_4051);
nand U4144 (N_4144,N_4080,N_4010);
and U4145 (N_4145,N_4029,N_4035);
nand U4146 (N_4146,N_4039,N_4042);
or U4147 (N_4147,N_4043,N_4099);
xnor U4148 (N_4148,N_4040,N_4014);
or U4149 (N_4149,N_4047,N_4028);
and U4150 (N_4150,N_4071,N_4063);
nor U4151 (N_4151,N_4060,N_4090);
nor U4152 (N_4152,N_4038,N_4026);
or U4153 (N_4153,N_4022,N_4056);
and U4154 (N_4154,N_4018,N_4077);
and U4155 (N_4155,N_4045,N_4037);
nor U4156 (N_4156,N_4037,N_4036);
or U4157 (N_4157,N_4078,N_4079);
or U4158 (N_4158,N_4033,N_4091);
nand U4159 (N_4159,N_4077,N_4061);
or U4160 (N_4160,N_4038,N_4064);
and U4161 (N_4161,N_4018,N_4032);
or U4162 (N_4162,N_4007,N_4045);
and U4163 (N_4163,N_4032,N_4075);
nand U4164 (N_4164,N_4003,N_4092);
or U4165 (N_4165,N_4097,N_4090);
or U4166 (N_4166,N_4000,N_4087);
and U4167 (N_4167,N_4072,N_4055);
or U4168 (N_4168,N_4098,N_4018);
and U4169 (N_4169,N_4009,N_4085);
and U4170 (N_4170,N_4003,N_4095);
nand U4171 (N_4171,N_4073,N_4037);
and U4172 (N_4172,N_4093,N_4054);
or U4173 (N_4173,N_4028,N_4042);
or U4174 (N_4174,N_4001,N_4050);
nand U4175 (N_4175,N_4074,N_4089);
and U4176 (N_4176,N_4072,N_4050);
or U4177 (N_4177,N_4031,N_4061);
and U4178 (N_4178,N_4040,N_4016);
nand U4179 (N_4179,N_4034,N_4069);
nor U4180 (N_4180,N_4028,N_4052);
or U4181 (N_4181,N_4012,N_4013);
or U4182 (N_4182,N_4050,N_4057);
nand U4183 (N_4183,N_4058,N_4064);
nor U4184 (N_4184,N_4090,N_4070);
nor U4185 (N_4185,N_4023,N_4080);
nand U4186 (N_4186,N_4058,N_4056);
or U4187 (N_4187,N_4088,N_4003);
nand U4188 (N_4188,N_4066,N_4033);
or U4189 (N_4189,N_4033,N_4075);
and U4190 (N_4190,N_4066,N_4092);
or U4191 (N_4191,N_4095,N_4024);
and U4192 (N_4192,N_4042,N_4025);
nand U4193 (N_4193,N_4075,N_4044);
nand U4194 (N_4194,N_4003,N_4044);
or U4195 (N_4195,N_4094,N_4053);
nand U4196 (N_4196,N_4018,N_4064);
and U4197 (N_4197,N_4011,N_4056);
nor U4198 (N_4198,N_4088,N_4000);
and U4199 (N_4199,N_4027,N_4025);
or U4200 (N_4200,N_4150,N_4173);
xnor U4201 (N_4201,N_4197,N_4179);
or U4202 (N_4202,N_4152,N_4133);
xor U4203 (N_4203,N_4129,N_4162);
and U4204 (N_4204,N_4172,N_4175);
and U4205 (N_4205,N_4141,N_4146);
and U4206 (N_4206,N_4130,N_4110);
or U4207 (N_4207,N_4187,N_4196);
nand U4208 (N_4208,N_4134,N_4164);
nor U4209 (N_4209,N_4193,N_4140);
nand U4210 (N_4210,N_4183,N_4144);
nand U4211 (N_4211,N_4192,N_4127);
nand U4212 (N_4212,N_4168,N_4190);
or U4213 (N_4213,N_4131,N_4106);
nor U4214 (N_4214,N_4116,N_4161);
nor U4215 (N_4215,N_4100,N_4142);
xnor U4216 (N_4216,N_4107,N_4123);
or U4217 (N_4217,N_4194,N_4135);
xor U4218 (N_4218,N_4189,N_4149);
nor U4219 (N_4219,N_4125,N_4126);
and U4220 (N_4220,N_4111,N_4124);
and U4221 (N_4221,N_4128,N_4158);
nor U4222 (N_4222,N_4109,N_4169);
nor U4223 (N_4223,N_4122,N_4171);
nand U4224 (N_4224,N_4114,N_4138);
xor U4225 (N_4225,N_4188,N_4163);
and U4226 (N_4226,N_4180,N_4165);
nand U4227 (N_4227,N_4104,N_4139);
nor U4228 (N_4228,N_4121,N_4143);
xnor U4229 (N_4229,N_4115,N_4102);
nand U4230 (N_4230,N_4113,N_4160);
xor U4231 (N_4231,N_4156,N_4176);
nand U4232 (N_4232,N_4119,N_4198);
nand U4233 (N_4233,N_4195,N_4177);
nor U4234 (N_4234,N_4174,N_4136);
and U4235 (N_4235,N_4155,N_4151);
nor U4236 (N_4236,N_4167,N_4120);
and U4237 (N_4237,N_4101,N_4181);
nand U4238 (N_4238,N_4153,N_4103);
or U4239 (N_4239,N_4191,N_4159);
xor U4240 (N_4240,N_4184,N_4185);
xnor U4241 (N_4241,N_4157,N_4137);
and U4242 (N_4242,N_4145,N_4105);
xor U4243 (N_4243,N_4148,N_4186);
nand U4244 (N_4244,N_4182,N_4118);
or U4245 (N_4245,N_4112,N_4178);
nor U4246 (N_4246,N_4166,N_4117);
nor U4247 (N_4247,N_4108,N_4132);
and U4248 (N_4248,N_4170,N_4154);
and U4249 (N_4249,N_4147,N_4199);
nor U4250 (N_4250,N_4127,N_4133);
and U4251 (N_4251,N_4187,N_4199);
nand U4252 (N_4252,N_4171,N_4148);
or U4253 (N_4253,N_4118,N_4108);
nand U4254 (N_4254,N_4130,N_4155);
and U4255 (N_4255,N_4119,N_4139);
or U4256 (N_4256,N_4164,N_4115);
nor U4257 (N_4257,N_4175,N_4168);
and U4258 (N_4258,N_4162,N_4111);
and U4259 (N_4259,N_4169,N_4127);
nand U4260 (N_4260,N_4168,N_4134);
and U4261 (N_4261,N_4128,N_4118);
or U4262 (N_4262,N_4100,N_4139);
or U4263 (N_4263,N_4129,N_4197);
and U4264 (N_4264,N_4166,N_4180);
nor U4265 (N_4265,N_4138,N_4127);
nor U4266 (N_4266,N_4162,N_4169);
or U4267 (N_4267,N_4195,N_4109);
or U4268 (N_4268,N_4144,N_4122);
nand U4269 (N_4269,N_4190,N_4116);
and U4270 (N_4270,N_4118,N_4174);
nand U4271 (N_4271,N_4164,N_4158);
nor U4272 (N_4272,N_4131,N_4181);
nand U4273 (N_4273,N_4100,N_4158);
or U4274 (N_4274,N_4166,N_4113);
nand U4275 (N_4275,N_4120,N_4146);
and U4276 (N_4276,N_4121,N_4196);
or U4277 (N_4277,N_4179,N_4122);
xnor U4278 (N_4278,N_4119,N_4175);
and U4279 (N_4279,N_4139,N_4101);
and U4280 (N_4280,N_4136,N_4148);
nand U4281 (N_4281,N_4106,N_4199);
xor U4282 (N_4282,N_4108,N_4113);
or U4283 (N_4283,N_4158,N_4138);
xnor U4284 (N_4284,N_4134,N_4119);
and U4285 (N_4285,N_4123,N_4153);
nand U4286 (N_4286,N_4181,N_4169);
nor U4287 (N_4287,N_4117,N_4172);
and U4288 (N_4288,N_4189,N_4118);
and U4289 (N_4289,N_4113,N_4107);
and U4290 (N_4290,N_4153,N_4115);
nand U4291 (N_4291,N_4110,N_4101);
and U4292 (N_4292,N_4157,N_4129);
or U4293 (N_4293,N_4113,N_4159);
or U4294 (N_4294,N_4157,N_4134);
xor U4295 (N_4295,N_4112,N_4167);
nand U4296 (N_4296,N_4175,N_4106);
nor U4297 (N_4297,N_4165,N_4111);
or U4298 (N_4298,N_4157,N_4185);
xnor U4299 (N_4299,N_4168,N_4140);
and U4300 (N_4300,N_4250,N_4246);
nand U4301 (N_4301,N_4230,N_4251);
and U4302 (N_4302,N_4216,N_4284);
and U4303 (N_4303,N_4244,N_4256);
nand U4304 (N_4304,N_4289,N_4260);
nand U4305 (N_4305,N_4226,N_4217);
or U4306 (N_4306,N_4257,N_4255);
nor U4307 (N_4307,N_4228,N_4268);
xor U4308 (N_4308,N_4219,N_4221);
and U4309 (N_4309,N_4227,N_4215);
or U4310 (N_4310,N_4274,N_4299);
or U4311 (N_4311,N_4294,N_4214);
xnor U4312 (N_4312,N_4285,N_4258);
xnor U4313 (N_4313,N_4283,N_4212);
nand U4314 (N_4314,N_4273,N_4281);
and U4315 (N_4315,N_4272,N_4276);
xor U4316 (N_4316,N_4287,N_4269);
nand U4317 (N_4317,N_4267,N_4265);
nand U4318 (N_4318,N_4253,N_4293);
nor U4319 (N_4319,N_4296,N_4233);
nor U4320 (N_4320,N_4213,N_4241);
or U4321 (N_4321,N_4220,N_4205);
or U4322 (N_4322,N_4280,N_4262);
and U4323 (N_4323,N_4263,N_4224);
nand U4324 (N_4324,N_4290,N_4211);
or U4325 (N_4325,N_4245,N_4201);
nor U4326 (N_4326,N_4200,N_4286);
nand U4327 (N_4327,N_4252,N_4292);
and U4328 (N_4328,N_4243,N_4277);
nand U4329 (N_4329,N_4297,N_4259);
nand U4330 (N_4330,N_4225,N_4218);
xor U4331 (N_4331,N_4247,N_4239);
or U4332 (N_4332,N_4248,N_4210);
xor U4333 (N_4333,N_4282,N_4295);
nor U4334 (N_4334,N_4264,N_4232);
and U4335 (N_4335,N_4298,N_4208);
nor U4336 (N_4336,N_4261,N_4222);
and U4337 (N_4337,N_4291,N_4235);
and U4338 (N_4338,N_4223,N_4288);
and U4339 (N_4339,N_4206,N_4203);
and U4340 (N_4340,N_4275,N_4202);
nor U4341 (N_4341,N_4249,N_4242);
and U4342 (N_4342,N_4270,N_4207);
or U4343 (N_4343,N_4237,N_4278);
nand U4344 (N_4344,N_4209,N_4254);
nand U4345 (N_4345,N_4236,N_4204);
and U4346 (N_4346,N_4234,N_4231);
and U4347 (N_4347,N_4229,N_4238);
or U4348 (N_4348,N_4279,N_4266);
nand U4349 (N_4349,N_4271,N_4240);
nor U4350 (N_4350,N_4293,N_4282);
nor U4351 (N_4351,N_4251,N_4205);
or U4352 (N_4352,N_4242,N_4271);
nor U4353 (N_4353,N_4243,N_4220);
nor U4354 (N_4354,N_4268,N_4277);
and U4355 (N_4355,N_4264,N_4213);
and U4356 (N_4356,N_4263,N_4220);
or U4357 (N_4357,N_4245,N_4259);
nor U4358 (N_4358,N_4234,N_4274);
xor U4359 (N_4359,N_4236,N_4249);
or U4360 (N_4360,N_4278,N_4203);
and U4361 (N_4361,N_4252,N_4283);
nand U4362 (N_4362,N_4281,N_4234);
and U4363 (N_4363,N_4284,N_4229);
nand U4364 (N_4364,N_4239,N_4220);
nor U4365 (N_4365,N_4230,N_4238);
nor U4366 (N_4366,N_4266,N_4236);
nor U4367 (N_4367,N_4283,N_4298);
and U4368 (N_4368,N_4200,N_4296);
or U4369 (N_4369,N_4251,N_4269);
and U4370 (N_4370,N_4255,N_4219);
nand U4371 (N_4371,N_4295,N_4208);
nand U4372 (N_4372,N_4239,N_4246);
nand U4373 (N_4373,N_4295,N_4245);
and U4374 (N_4374,N_4278,N_4281);
nand U4375 (N_4375,N_4259,N_4250);
nand U4376 (N_4376,N_4214,N_4273);
nor U4377 (N_4377,N_4273,N_4242);
and U4378 (N_4378,N_4203,N_4282);
nor U4379 (N_4379,N_4208,N_4249);
or U4380 (N_4380,N_4253,N_4213);
nand U4381 (N_4381,N_4267,N_4254);
and U4382 (N_4382,N_4264,N_4242);
nand U4383 (N_4383,N_4214,N_4270);
nor U4384 (N_4384,N_4255,N_4209);
xnor U4385 (N_4385,N_4292,N_4287);
nand U4386 (N_4386,N_4248,N_4255);
nand U4387 (N_4387,N_4248,N_4218);
nor U4388 (N_4388,N_4225,N_4260);
nor U4389 (N_4389,N_4275,N_4296);
xor U4390 (N_4390,N_4227,N_4220);
and U4391 (N_4391,N_4264,N_4220);
or U4392 (N_4392,N_4239,N_4219);
and U4393 (N_4393,N_4266,N_4257);
and U4394 (N_4394,N_4249,N_4284);
or U4395 (N_4395,N_4273,N_4208);
nand U4396 (N_4396,N_4292,N_4291);
nand U4397 (N_4397,N_4291,N_4216);
nand U4398 (N_4398,N_4264,N_4215);
and U4399 (N_4399,N_4203,N_4216);
nor U4400 (N_4400,N_4379,N_4370);
and U4401 (N_4401,N_4315,N_4349);
or U4402 (N_4402,N_4371,N_4372);
or U4403 (N_4403,N_4316,N_4375);
or U4404 (N_4404,N_4328,N_4398);
nor U4405 (N_4405,N_4364,N_4310);
and U4406 (N_4406,N_4333,N_4305);
or U4407 (N_4407,N_4321,N_4347);
and U4408 (N_4408,N_4373,N_4318);
xnor U4409 (N_4409,N_4312,N_4309);
or U4410 (N_4410,N_4319,N_4317);
or U4411 (N_4411,N_4322,N_4323);
xnor U4412 (N_4412,N_4377,N_4302);
xnor U4413 (N_4413,N_4397,N_4329);
nand U4414 (N_4414,N_4388,N_4369);
nor U4415 (N_4415,N_4343,N_4332);
xor U4416 (N_4416,N_4387,N_4300);
nand U4417 (N_4417,N_4352,N_4389);
nor U4418 (N_4418,N_4354,N_4358);
or U4419 (N_4419,N_4361,N_4381);
nand U4420 (N_4420,N_4380,N_4338);
nand U4421 (N_4421,N_4355,N_4301);
or U4422 (N_4422,N_4360,N_4350);
xor U4423 (N_4423,N_4337,N_4344);
nand U4424 (N_4424,N_4346,N_4365);
and U4425 (N_4425,N_4351,N_4335);
xnor U4426 (N_4426,N_4386,N_4367);
nor U4427 (N_4427,N_4391,N_4308);
or U4428 (N_4428,N_4326,N_4399);
and U4429 (N_4429,N_4324,N_4366);
nor U4430 (N_4430,N_4394,N_4382);
and U4431 (N_4431,N_4353,N_4307);
nand U4432 (N_4432,N_4378,N_4339);
xnor U4433 (N_4433,N_4342,N_4363);
nand U4434 (N_4434,N_4303,N_4345);
nor U4435 (N_4435,N_4340,N_4336);
nor U4436 (N_4436,N_4385,N_4395);
xnor U4437 (N_4437,N_4362,N_4348);
nand U4438 (N_4438,N_4311,N_4384);
nand U4439 (N_4439,N_4331,N_4325);
and U4440 (N_4440,N_4327,N_4383);
nor U4441 (N_4441,N_4359,N_4357);
xnor U4442 (N_4442,N_4306,N_4314);
nor U4443 (N_4443,N_4392,N_4368);
nand U4444 (N_4444,N_4304,N_4393);
and U4445 (N_4445,N_4396,N_4356);
and U4446 (N_4446,N_4320,N_4390);
and U4447 (N_4447,N_4341,N_4330);
or U4448 (N_4448,N_4334,N_4313);
and U4449 (N_4449,N_4376,N_4374);
or U4450 (N_4450,N_4391,N_4333);
and U4451 (N_4451,N_4395,N_4329);
xnor U4452 (N_4452,N_4369,N_4363);
and U4453 (N_4453,N_4326,N_4387);
and U4454 (N_4454,N_4388,N_4313);
and U4455 (N_4455,N_4347,N_4315);
and U4456 (N_4456,N_4335,N_4363);
xor U4457 (N_4457,N_4333,N_4373);
nor U4458 (N_4458,N_4321,N_4383);
and U4459 (N_4459,N_4308,N_4338);
nor U4460 (N_4460,N_4340,N_4388);
xor U4461 (N_4461,N_4325,N_4359);
and U4462 (N_4462,N_4369,N_4314);
nor U4463 (N_4463,N_4330,N_4391);
nand U4464 (N_4464,N_4332,N_4317);
nand U4465 (N_4465,N_4351,N_4316);
and U4466 (N_4466,N_4398,N_4343);
nand U4467 (N_4467,N_4356,N_4393);
xnor U4468 (N_4468,N_4370,N_4381);
nand U4469 (N_4469,N_4317,N_4369);
xor U4470 (N_4470,N_4351,N_4346);
nor U4471 (N_4471,N_4313,N_4370);
nand U4472 (N_4472,N_4319,N_4330);
nand U4473 (N_4473,N_4340,N_4300);
and U4474 (N_4474,N_4320,N_4359);
nor U4475 (N_4475,N_4362,N_4302);
nor U4476 (N_4476,N_4329,N_4322);
nand U4477 (N_4477,N_4386,N_4384);
nand U4478 (N_4478,N_4317,N_4337);
or U4479 (N_4479,N_4300,N_4376);
xor U4480 (N_4480,N_4360,N_4395);
and U4481 (N_4481,N_4382,N_4389);
or U4482 (N_4482,N_4349,N_4364);
nand U4483 (N_4483,N_4381,N_4330);
or U4484 (N_4484,N_4389,N_4308);
or U4485 (N_4485,N_4388,N_4367);
nor U4486 (N_4486,N_4382,N_4387);
and U4487 (N_4487,N_4337,N_4374);
xnor U4488 (N_4488,N_4322,N_4319);
nand U4489 (N_4489,N_4399,N_4336);
nor U4490 (N_4490,N_4312,N_4361);
or U4491 (N_4491,N_4342,N_4396);
nand U4492 (N_4492,N_4345,N_4335);
xor U4493 (N_4493,N_4309,N_4372);
and U4494 (N_4494,N_4348,N_4300);
or U4495 (N_4495,N_4342,N_4388);
and U4496 (N_4496,N_4399,N_4311);
nand U4497 (N_4497,N_4319,N_4314);
and U4498 (N_4498,N_4398,N_4332);
or U4499 (N_4499,N_4373,N_4308);
xnor U4500 (N_4500,N_4483,N_4417);
or U4501 (N_4501,N_4456,N_4479);
or U4502 (N_4502,N_4453,N_4486);
xor U4503 (N_4503,N_4433,N_4423);
and U4504 (N_4504,N_4404,N_4430);
nand U4505 (N_4505,N_4450,N_4452);
nand U4506 (N_4506,N_4458,N_4457);
nand U4507 (N_4507,N_4401,N_4403);
or U4508 (N_4508,N_4439,N_4448);
and U4509 (N_4509,N_4478,N_4491);
or U4510 (N_4510,N_4400,N_4424);
nand U4511 (N_4511,N_4487,N_4415);
and U4512 (N_4512,N_4492,N_4446);
xor U4513 (N_4513,N_4489,N_4480);
xnor U4514 (N_4514,N_4465,N_4470);
nor U4515 (N_4515,N_4472,N_4496);
and U4516 (N_4516,N_4451,N_4429);
nor U4517 (N_4517,N_4406,N_4402);
nand U4518 (N_4518,N_4419,N_4405);
and U4519 (N_4519,N_4428,N_4412);
nor U4520 (N_4520,N_4494,N_4481);
xor U4521 (N_4521,N_4482,N_4462);
and U4522 (N_4522,N_4416,N_4436);
nand U4523 (N_4523,N_4455,N_4408);
nor U4524 (N_4524,N_4437,N_4473);
and U4525 (N_4525,N_4432,N_4476);
xor U4526 (N_4526,N_4431,N_4407);
and U4527 (N_4527,N_4477,N_4425);
or U4528 (N_4528,N_4410,N_4447);
nand U4529 (N_4529,N_4443,N_4454);
nand U4530 (N_4530,N_4497,N_4490);
nand U4531 (N_4531,N_4499,N_4421);
nor U4532 (N_4532,N_4466,N_4435);
nand U4533 (N_4533,N_4413,N_4464);
nand U4534 (N_4534,N_4468,N_4495);
and U4535 (N_4535,N_4474,N_4471);
or U4536 (N_4536,N_4475,N_4414);
or U4537 (N_4537,N_4440,N_4460);
nand U4538 (N_4538,N_4438,N_4449);
and U4539 (N_4539,N_4418,N_4461);
nand U4540 (N_4540,N_4488,N_4445);
xor U4541 (N_4541,N_4467,N_4434);
nor U4542 (N_4542,N_4422,N_4463);
and U4543 (N_4543,N_4459,N_4444);
or U4544 (N_4544,N_4442,N_4411);
or U4545 (N_4545,N_4427,N_4420);
nand U4546 (N_4546,N_4485,N_4498);
and U4547 (N_4547,N_4493,N_4469);
and U4548 (N_4548,N_4426,N_4484);
and U4549 (N_4549,N_4409,N_4441);
or U4550 (N_4550,N_4483,N_4428);
nand U4551 (N_4551,N_4452,N_4404);
or U4552 (N_4552,N_4491,N_4446);
or U4553 (N_4553,N_4478,N_4423);
or U4554 (N_4554,N_4439,N_4447);
nor U4555 (N_4555,N_4447,N_4459);
nand U4556 (N_4556,N_4420,N_4401);
or U4557 (N_4557,N_4460,N_4421);
nor U4558 (N_4558,N_4423,N_4455);
nor U4559 (N_4559,N_4441,N_4404);
nand U4560 (N_4560,N_4401,N_4443);
nand U4561 (N_4561,N_4425,N_4437);
nand U4562 (N_4562,N_4404,N_4498);
and U4563 (N_4563,N_4448,N_4400);
xnor U4564 (N_4564,N_4468,N_4481);
nor U4565 (N_4565,N_4473,N_4435);
nor U4566 (N_4566,N_4461,N_4458);
and U4567 (N_4567,N_4415,N_4433);
and U4568 (N_4568,N_4410,N_4425);
nor U4569 (N_4569,N_4480,N_4433);
or U4570 (N_4570,N_4405,N_4455);
or U4571 (N_4571,N_4470,N_4455);
or U4572 (N_4572,N_4422,N_4431);
xnor U4573 (N_4573,N_4435,N_4411);
nor U4574 (N_4574,N_4431,N_4410);
and U4575 (N_4575,N_4414,N_4484);
and U4576 (N_4576,N_4451,N_4497);
or U4577 (N_4577,N_4483,N_4491);
or U4578 (N_4578,N_4414,N_4429);
nor U4579 (N_4579,N_4491,N_4432);
or U4580 (N_4580,N_4439,N_4475);
nor U4581 (N_4581,N_4467,N_4495);
xor U4582 (N_4582,N_4452,N_4422);
or U4583 (N_4583,N_4439,N_4493);
nand U4584 (N_4584,N_4438,N_4494);
and U4585 (N_4585,N_4483,N_4490);
and U4586 (N_4586,N_4489,N_4441);
nand U4587 (N_4587,N_4458,N_4406);
and U4588 (N_4588,N_4400,N_4484);
or U4589 (N_4589,N_4414,N_4412);
nor U4590 (N_4590,N_4481,N_4425);
nor U4591 (N_4591,N_4458,N_4437);
nor U4592 (N_4592,N_4428,N_4478);
and U4593 (N_4593,N_4423,N_4417);
and U4594 (N_4594,N_4404,N_4431);
nor U4595 (N_4595,N_4409,N_4439);
and U4596 (N_4596,N_4491,N_4428);
xor U4597 (N_4597,N_4474,N_4472);
nor U4598 (N_4598,N_4468,N_4456);
nor U4599 (N_4599,N_4415,N_4470);
nand U4600 (N_4600,N_4558,N_4597);
nor U4601 (N_4601,N_4502,N_4566);
nand U4602 (N_4602,N_4527,N_4500);
nor U4603 (N_4603,N_4592,N_4565);
xnor U4604 (N_4604,N_4506,N_4546);
nor U4605 (N_4605,N_4516,N_4518);
nor U4606 (N_4606,N_4578,N_4582);
and U4607 (N_4607,N_4526,N_4567);
and U4608 (N_4608,N_4523,N_4579);
nor U4609 (N_4609,N_4521,N_4573);
nor U4610 (N_4610,N_4510,N_4569);
nor U4611 (N_4611,N_4515,N_4596);
nand U4612 (N_4612,N_4501,N_4551);
and U4613 (N_4613,N_4548,N_4561);
nand U4614 (N_4614,N_4590,N_4520);
nand U4615 (N_4615,N_4503,N_4513);
nor U4616 (N_4616,N_4563,N_4581);
nor U4617 (N_4617,N_4542,N_4544);
and U4618 (N_4618,N_4530,N_4505);
nand U4619 (N_4619,N_4564,N_4538);
nand U4620 (N_4620,N_4512,N_4560);
nor U4621 (N_4621,N_4508,N_4529);
or U4622 (N_4622,N_4519,N_4535);
nor U4623 (N_4623,N_4528,N_4532);
and U4624 (N_4624,N_4550,N_4553);
or U4625 (N_4625,N_4580,N_4545);
and U4626 (N_4626,N_4577,N_4525);
nand U4627 (N_4627,N_4509,N_4514);
nor U4628 (N_4628,N_4593,N_4594);
or U4629 (N_4629,N_4555,N_4595);
nand U4630 (N_4630,N_4504,N_4522);
nor U4631 (N_4631,N_4571,N_4562);
or U4632 (N_4632,N_4589,N_4507);
nor U4633 (N_4633,N_4534,N_4570);
or U4634 (N_4634,N_4588,N_4554);
and U4635 (N_4635,N_4587,N_4552);
nor U4636 (N_4636,N_4539,N_4598);
and U4637 (N_4637,N_4557,N_4547);
and U4638 (N_4638,N_4572,N_4586);
nand U4639 (N_4639,N_4541,N_4533);
or U4640 (N_4640,N_4584,N_4576);
nor U4641 (N_4641,N_4591,N_4549);
or U4642 (N_4642,N_4540,N_4583);
or U4643 (N_4643,N_4517,N_4556);
xor U4644 (N_4644,N_4575,N_4559);
nor U4645 (N_4645,N_4524,N_4568);
and U4646 (N_4646,N_4599,N_4585);
nand U4647 (N_4647,N_4537,N_4531);
xor U4648 (N_4648,N_4511,N_4536);
nor U4649 (N_4649,N_4574,N_4543);
or U4650 (N_4650,N_4531,N_4572);
or U4651 (N_4651,N_4518,N_4540);
nand U4652 (N_4652,N_4598,N_4555);
and U4653 (N_4653,N_4564,N_4507);
nand U4654 (N_4654,N_4508,N_4520);
nand U4655 (N_4655,N_4574,N_4532);
nor U4656 (N_4656,N_4580,N_4582);
nor U4657 (N_4657,N_4558,N_4510);
and U4658 (N_4658,N_4510,N_4572);
nor U4659 (N_4659,N_4575,N_4530);
nand U4660 (N_4660,N_4504,N_4531);
or U4661 (N_4661,N_4553,N_4531);
xnor U4662 (N_4662,N_4501,N_4523);
xor U4663 (N_4663,N_4548,N_4546);
nor U4664 (N_4664,N_4518,N_4566);
nand U4665 (N_4665,N_4594,N_4553);
and U4666 (N_4666,N_4542,N_4515);
nor U4667 (N_4667,N_4549,N_4575);
and U4668 (N_4668,N_4573,N_4547);
nand U4669 (N_4669,N_4568,N_4573);
nand U4670 (N_4670,N_4538,N_4558);
nor U4671 (N_4671,N_4540,N_4501);
and U4672 (N_4672,N_4570,N_4520);
nor U4673 (N_4673,N_4559,N_4573);
or U4674 (N_4674,N_4514,N_4569);
nand U4675 (N_4675,N_4508,N_4552);
nor U4676 (N_4676,N_4590,N_4576);
or U4677 (N_4677,N_4543,N_4565);
or U4678 (N_4678,N_4558,N_4564);
nor U4679 (N_4679,N_4537,N_4517);
or U4680 (N_4680,N_4516,N_4568);
nor U4681 (N_4681,N_4522,N_4593);
nand U4682 (N_4682,N_4505,N_4501);
or U4683 (N_4683,N_4531,N_4586);
nand U4684 (N_4684,N_4596,N_4512);
and U4685 (N_4685,N_4598,N_4557);
and U4686 (N_4686,N_4503,N_4528);
nor U4687 (N_4687,N_4525,N_4598);
and U4688 (N_4688,N_4525,N_4546);
and U4689 (N_4689,N_4542,N_4518);
nor U4690 (N_4690,N_4579,N_4561);
and U4691 (N_4691,N_4548,N_4542);
and U4692 (N_4692,N_4573,N_4524);
nand U4693 (N_4693,N_4507,N_4540);
nand U4694 (N_4694,N_4587,N_4501);
and U4695 (N_4695,N_4523,N_4586);
nand U4696 (N_4696,N_4548,N_4552);
nor U4697 (N_4697,N_4548,N_4584);
and U4698 (N_4698,N_4562,N_4591);
nor U4699 (N_4699,N_4585,N_4509);
nand U4700 (N_4700,N_4663,N_4699);
nor U4701 (N_4701,N_4681,N_4636);
or U4702 (N_4702,N_4618,N_4695);
or U4703 (N_4703,N_4696,N_4633);
or U4704 (N_4704,N_4649,N_4611);
or U4705 (N_4705,N_4668,N_4609);
or U4706 (N_4706,N_4682,N_4625);
or U4707 (N_4707,N_4679,N_4688);
or U4708 (N_4708,N_4675,N_4652);
or U4709 (N_4709,N_4674,N_4641);
nor U4710 (N_4710,N_4639,N_4672);
xor U4711 (N_4711,N_4677,N_4647);
xor U4712 (N_4712,N_4676,N_4685);
nor U4713 (N_4713,N_4607,N_4623);
xnor U4714 (N_4714,N_4622,N_4643);
xnor U4715 (N_4715,N_4610,N_4693);
nor U4716 (N_4716,N_4673,N_4660);
nor U4717 (N_4717,N_4645,N_4698);
nand U4718 (N_4718,N_4644,N_4640);
xor U4719 (N_4719,N_4608,N_4613);
and U4720 (N_4720,N_4616,N_4691);
or U4721 (N_4721,N_4683,N_4628);
nand U4722 (N_4722,N_4666,N_4651);
and U4723 (N_4723,N_4621,N_4642);
nor U4724 (N_4724,N_4626,N_4614);
nand U4725 (N_4725,N_4662,N_4612);
or U4726 (N_4726,N_4637,N_4606);
or U4727 (N_4727,N_4678,N_4635);
and U4728 (N_4728,N_4670,N_4600);
and U4729 (N_4729,N_4619,N_4680);
nand U4730 (N_4730,N_4605,N_4689);
or U4731 (N_4731,N_4667,N_4631);
xor U4732 (N_4732,N_4632,N_4658);
or U4733 (N_4733,N_4657,N_4601);
or U4734 (N_4734,N_4654,N_4694);
or U4735 (N_4735,N_4665,N_4615);
nand U4736 (N_4736,N_4655,N_4617);
and U4737 (N_4737,N_4650,N_4692);
nor U4738 (N_4738,N_4664,N_4697);
and U4739 (N_4739,N_4629,N_4656);
and U4740 (N_4740,N_4603,N_4627);
xor U4741 (N_4741,N_4659,N_4671);
nor U4742 (N_4742,N_4634,N_4684);
nand U4743 (N_4743,N_4602,N_4648);
nand U4744 (N_4744,N_4630,N_4686);
nor U4745 (N_4745,N_4638,N_4687);
and U4746 (N_4746,N_4620,N_4604);
xnor U4747 (N_4747,N_4669,N_4646);
nor U4748 (N_4748,N_4661,N_4624);
nor U4749 (N_4749,N_4653,N_4690);
nor U4750 (N_4750,N_4620,N_4649);
or U4751 (N_4751,N_4637,N_4635);
xor U4752 (N_4752,N_4649,N_4641);
nand U4753 (N_4753,N_4661,N_4610);
xnor U4754 (N_4754,N_4672,N_4612);
nor U4755 (N_4755,N_4609,N_4618);
and U4756 (N_4756,N_4630,N_4695);
nand U4757 (N_4757,N_4673,N_4689);
nand U4758 (N_4758,N_4688,N_4603);
nor U4759 (N_4759,N_4629,N_4657);
or U4760 (N_4760,N_4634,N_4688);
nor U4761 (N_4761,N_4670,N_4615);
nor U4762 (N_4762,N_4623,N_4681);
xnor U4763 (N_4763,N_4627,N_4674);
nand U4764 (N_4764,N_4616,N_4625);
and U4765 (N_4765,N_4602,N_4665);
nor U4766 (N_4766,N_4647,N_4676);
xor U4767 (N_4767,N_4675,N_4640);
or U4768 (N_4768,N_4616,N_4604);
and U4769 (N_4769,N_4646,N_4691);
nor U4770 (N_4770,N_4698,N_4670);
nand U4771 (N_4771,N_4666,N_4673);
xnor U4772 (N_4772,N_4673,N_4657);
and U4773 (N_4773,N_4668,N_4677);
nand U4774 (N_4774,N_4654,N_4653);
or U4775 (N_4775,N_4632,N_4666);
nand U4776 (N_4776,N_4614,N_4634);
nor U4777 (N_4777,N_4680,N_4681);
nor U4778 (N_4778,N_4684,N_4636);
and U4779 (N_4779,N_4695,N_4628);
nand U4780 (N_4780,N_4652,N_4609);
or U4781 (N_4781,N_4602,N_4677);
nor U4782 (N_4782,N_4620,N_4692);
or U4783 (N_4783,N_4626,N_4604);
nor U4784 (N_4784,N_4639,N_4625);
xnor U4785 (N_4785,N_4607,N_4696);
and U4786 (N_4786,N_4647,N_4659);
nand U4787 (N_4787,N_4667,N_4649);
nor U4788 (N_4788,N_4664,N_4603);
nand U4789 (N_4789,N_4609,N_4669);
xnor U4790 (N_4790,N_4678,N_4672);
nand U4791 (N_4791,N_4668,N_4681);
nand U4792 (N_4792,N_4605,N_4687);
nor U4793 (N_4793,N_4650,N_4645);
nor U4794 (N_4794,N_4618,N_4621);
and U4795 (N_4795,N_4648,N_4622);
nor U4796 (N_4796,N_4629,N_4658);
nor U4797 (N_4797,N_4622,N_4696);
or U4798 (N_4798,N_4630,N_4623);
and U4799 (N_4799,N_4620,N_4641);
and U4800 (N_4800,N_4708,N_4749);
and U4801 (N_4801,N_4780,N_4763);
and U4802 (N_4802,N_4740,N_4774);
and U4803 (N_4803,N_4765,N_4782);
and U4804 (N_4804,N_4790,N_4752);
or U4805 (N_4805,N_4796,N_4716);
or U4806 (N_4806,N_4704,N_4721);
or U4807 (N_4807,N_4703,N_4776);
xnor U4808 (N_4808,N_4739,N_4746);
nor U4809 (N_4809,N_4729,N_4702);
nor U4810 (N_4810,N_4715,N_4748);
and U4811 (N_4811,N_4726,N_4755);
nand U4812 (N_4812,N_4725,N_4760);
nor U4813 (N_4813,N_4786,N_4727);
nand U4814 (N_4814,N_4728,N_4733);
nand U4815 (N_4815,N_4743,N_4754);
nand U4816 (N_4816,N_4747,N_4722);
or U4817 (N_4817,N_4718,N_4798);
and U4818 (N_4818,N_4730,N_4738);
or U4819 (N_4819,N_4745,N_4764);
nand U4820 (N_4820,N_4719,N_4756);
or U4821 (N_4821,N_4735,N_4714);
nand U4822 (N_4822,N_4758,N_4709);
xor U4823 (N_4823,N_4705,N_4791);
and U4824 (N_4824,N_4797,N_4766);
nand U4825 (N_4825,N_4794,N_4770);
or U4826 (N_4826,N_4731,N_4707);
and U4827 (N_4827,N_4779,N_4751);
xor U4828 (N_4828,N_4717,N_4710);
xnor U4829 (N_4829,N_4723,N_4783);
and U4830 (N_4830,N_4769,N_4789);
and U4831 (N_4831,N_4767,N_4788);
or U4832 (N_4832,N_4732,N_4762);
or U4833 (N_4833,N_4737,N_4724);
or U4834 (N_4834,N_4701,N_4775);
or U4835 (N_4835,N_4772,N_4712);
nor U4836 (N_4836,N_4771,N_4734);
nor U4837 (N_4837,N_4784,N_4795);
or U4838 (N_4838,N_4706,N_4773);
and U4839 (N_4839,N_4759,N_4741);
nand U4840 (N_4840,N_4781,N_4700);
xor U4841 (N_4841,N_4744,N_4736);
or U4842 (N_4842,N_4711,N_4750);
and U4843 (N_4843,N_4778,N_4777);
xor U4844 (N_4844,N_4720,N_4787);
and U4845 (N_4845,N_4761,N_4799);
nand U4846 (N_4846,N_4753,N_4757);
or U4847 (N_4847,N_4713,N_4768);
nor U4848 (N_4848,N_4785,N_4793);
or U4849 (N_4849,N_4792,N_4742);
nand U4850 (N_4850,N_4742,N_4780);
or U4851 (N_4851,N_4788,N_4747);
nand U4852 (N_4852,N_4763,N_4792);
and U4853 (N_4853,N_4711,N_4715);
nand U4854 (N_4854,N_4734,N_4797);
nand U4855 (N_4855,N_4718,N_4758);
or U4856 (N_4856,N_4787,N_4768);
and U4857 (N_4857,N_4742,N_4711);
and U4858 (N_4858,N_4768,N_4724);
nand U4859 (N_4859,N_4709,N_4732);
and U4860 (N_4860,N_4756,N_4781);
and U4861 (N_4861,N_4785,N_4753);
nand U4862 (N_4862,N_4757,N_4781);
or U4863 (N_4863,N_4714,N_4773);
nor U4864 (N_4864,N_4788,N_4754);
and U4865 (N_4865,N_4794,N_4711);
and U4866 (N_4866,N_4760,N_4742);
nand U4867 (N_4867,N_4785,N_4795);
nor U4868 (N_4868,N_4752,N_4727);
nor U4869 (N_4869,N_4722,N_4706);
xor U4870 (N_4870,N_4774,N_4750);
xor U4871 (N_4871,N_4788,N_4769);
xor U4872 (N_4872,N_4713,N_4775);
and U4873 (N_4873,N_4758,N_4739);
nand U4874 (N_4874,N_4700,N_4786);
nand U4875 (N_4875,N_4729,N_4774);
nand U4876 (N_4876,N_4762,N_4781);
xnor U4877 (N_4877,N_4711,N_4799);
or U4878 (N_4878,N_4797,N_4715);
xnor U4879 (N_4879,N_4769,N_4724);
nand U4880 (N_4880,N_4721,N_4724);
nand U4881 (N_4881,N_4742,N_4778);
nand U4882 (N_4882,N_4719,N_4796);
or U4883 (N_4883,N_4757,N_4784);
nor U4884 (N_4884,N_4780,N_4736);
and U4885 (N_4885,N_4796,N_4755);
nand U4886 (N_4886,N_4776,N_4738);
and U4887 (N_4887,N_4736,N_4798);
nand U4888 (N_4888,N_4773,N_4792);
or U4889 (N_4889,N_4767,N_4734);
nand U4890 (N_4890,N_4751,N_4750);
nor U4891 (N_4891,N_4754,N_4774);
nor U4892 (N_4892,N_4711,N_4762);
and U4893 (N_4893,N_4757,N_4715);
nand U4894 (N_4894,N_4777,N_4743);
nand U4895 (N_4895,N_4726,N_4764);
nor U4896 (N_4896,N_4754,N_4755);
and U4897 (N_4897,N_4748,N_4756);
nand U4898 (N_4898,N_4736,N_4727);
and U4899 (N_4899,N_4734,N_4730);
xor U4900 (N_4900,N_4850,N_4847);
xor U4901 (N_4901,N_4840,N_4880);
nor U4902 (N_4902,N_4829,N_4889);
or U4903 (N_4903,N_4874,N_4837);
and U4904 (N_4904,N_4828,N_4863);
or U4905 (N_4905,N_4876,N_4814);
nand U4906 (N_4906,N_4879,N_4877);
nor U4907 (N_4907,N_4864,N_4807);
nor U4908 (N_4908,N_4812,N_4816);
nand U4909 (N_4909,N_4805,N_4857);
xor U4910 (N_4910,N_4819,N_4804);
nand U4911 (N_4911,N_4859,N_4854);
and U4912 (N_4912,N_4852,N_4867);
or U4913 (N_4913,N_4820,N_4825);
and U4914 (N_4914,N_4878,N_4842);
and U4915 (N_4915,N_4885,N_4873);
or U4916 (N_4916,N_4849,N_4886);
and U4917 (N_4917,N_4895,N_4898);
nand U4918 (N_4918,N_4891,N_4836);
nand U4919 (N_4919,N_4810,N_4835);
nor U4920 (N_4920,N_4802,N_4893);
or U4921 (N_4921,N_4843,N_4848);
nand U4922 (N_4922,N_4826,N_4887);
xor U4923 (N_4923,N_4821,N_4856);
or U4924 (N_4924,N_4888,N_4831);
and U4925 (N_4925,N_4830,N_4803);
nor U4926 (N_4926,N_4806,N_4851);
and U4927 (N_4927,N_4818,N_4823);
or U4928 (N_4928,N_4865,N_4882);
and U4929 (N_4929,N_4890,N_4861);
nand U4930 (N_4930,N_4875,N_4862);
nand U4931 (N_4931,N_4871,N_4884);
nand U4932 (N_4932,N_4853,N_4811);
nor U4933 (N_4933,N_4800,N_4834);
nand U4934 (N_4934,N_4881,N_4866);
nand U4935 (N_4935,N_4896,N_4869);
nand U4936 (N_4936,N_4860,N_4832);
and U4937 (N_4937,N_4817,N_4883);
or U4938 (N_4938,N_4868,N_4841);
or U4939 (N_4939,N_4855,N_4894);
nand U4940 (N_4940,N_4824,N_4838);
and U4941 (N_4941,N_4813,N_4801);
nand U4942 (N_4942,N_4897,N_4822);
nor U4943 (N_4943,N_4839,N_4845);
nor U4944 (N_4944,N_4899,N_4808);
nand U4945 (N_4945,N_4833,N_4858);
nor U4946 (N_4946,N_4892,N_4809);
or U4947 (N_4947,N_4844,N_4846);
nand U4948 (N_4948,N_4827,N_4872);
nor U4949 (N_4949,N_4870,N_4815);
nand U4950 (N_4950,N_4883,N_4875);
nand U4951 (N_4951,N_4858,N_4836);
and U4952 (N_4952,N_4853,N_4883);
nand U4953 (N_4953,N_4895,N_4810);
nand U4954 (N_4954,N_4824,N_4815);
xor U4955 (N_4955,N_4894,N_4856);
and U4956 (N_4956,N_4803,N_4801);
and U4957 (N_4957,N_4845,N_4804);
nand U4958 (N_4958,N_4816,N_4840);
and U4959 (N_4959,N_4812,N_4801);
and U4960 (N_4960,N_4868,N_4852);
nand U4961 (N_4961,N_4897,N_4856);
xor U4962 (N_4962,N_4884,N_4885);
and U4963 (N_4963,N_4853,N_4880);
nor U4964 (N_4964,N_4846,N_4843);
nand U4965 (N_4965,N_4835,N_4842);
nor U4966 (N_4966,N_4846,N_4808);
and U4967 (N_4967,N_4871,N_4835);
nor U4968 (N_4968,N_4863,N_4885);
xor U4969 (N_4969,N_4824,N_4870);
nor U4970 (N_4970,N_4866,N_4814);
xnor U4971 (N_4971,N_4831,N_4801);
and U4972 (N_4972,N_4824,N_4867);
nor U4973 (N_4973,N_4818,N_4824);
nand U4974 (N_4974,N_4853,N_4806);
nor U4975 (N_4975,N_4834,N_4806);
or U4976 (N_4976,N_4810,N_4866);
and U4977 (N_4977,N_4844,N_4895);
or U4978 (N_4978,N_4886,N_4845);
xor U4979 (N_4979,N_4859,N_4827);
nand U4980 (N_4980,N_4848,N_4831);
or U4981 (N_4981,N_4840,N_4813);
xor U4982 (N_4982,N_4836,N_4830);
xnor U4983 (N_4983,N_4849,N_4847);
and U4984 (N_4984,N_4817,N_4808);
nand U4985 (N_4985,N_4870,N_4879);
or U4986 (N_4986,N_4842,N_4802);
nor U4987 (N_4987,N_4877,N_4837);
and U4988 (N_4988,N_4824,N_4803);
nor U4989 (N_4989,N_4858,N_4870);
and U4990 (N_4990,N_4866,N_4889);
and U4991 (N_4991,N_4831,N_4817);
and U4992 (N_4992,N_4889,N_4834);
or U4993 (N_4993,N_4867,N_4865);
and U4994 (N_4994,N_4890,N_4837);
nand U4995 (N_4995,N_4863,N_4847);
or U4996 (N_4996,N_4833,N_4869);
and U4997 (N_4997,N_4898,N_4863);
or U4998 (N_4998,N_4828,N_4880);
nand U4999 (N_4999,N_4859,N_4885);
nor U5000 (N_5000,N_4947,N_4913);
or U5001 (N_5001,N_4986,N_4981);
nor U5002 (N_5002,N_4988,N_4967);
or U5003 (N_5003,N_4973,N_4952);
or U5004 (N_5004,N_4995,N_4983);
nor U5005 (N_5005,N_4919,N_4931);
nand U5006 (N_5006,N_4962,N_4950);
and U5007 (N_5007,N_4917,N_4900);
or U5008 (N_5008,N_4909,N_4978);
nor U5009 (N_5009,N_4956,N_4963);
nand U5010 (N_5010,N_4916,N_4996);
xor U5011 (N_5011,N_4915,N_4907);
nand U5012 (N_5012,N_4966,N_4987);
nand U5013 (N_5013,N_4980,N_4975);
and U5014 (N_5014,N_4935,N_4911);
nor U5015 (N_5015,N_4905,N_4968);
nand U5016 (N_5016,N_4985,N_4903);
and U5017 (N_5017,N_4937,N_4974);
nor U5018 (N_5018,N_4940,N_4920);
or U5019 (N_5019,N_4918,N_4925);
or U5020 (N_5020,N_4939,N_4926);
nand U5021 (N_5021,N_4998,N_4902);
nand U5022 (N_5022,N_4906,N_4958);
nand U5023 (N_5023,N_4994,N_4960);
nor U5024 (N_5024,N_4999,N_4972);
or U5025 (N_5025,N_4961,N_4979);
nand U5026 (N_5026,N_4921,N_4982);
and U5027 (N_5027,N_4989,N_4928);
or U5028 (N_5028,N_4970,N_4951);
or U5029 (N_5029,N_4930,N_4922);
or U5030 (N_5030,N_4993,N_4969);
nand U5031 (N_5031,N_4959,N_4929);
nand U5032 (N_5032,N_4908,N_4945);
and U5033 (N_5033,N_4965,N_4914);
or U5034 (N_5034,N_4932,N_4944);
xor U5035 (N_5035,N_4942,N_4955);
or U5036 (N_5036,N_4954,N_4964);
xnor U5037 (N_5037,N_4946,N_4924);
nor U5038 (N_5038,N_4901,N_4990);
and U5039 (N_5039,N_4991,N_4927);
and U5040 (N_5040,N_4984,N_4923);
or U5041 (N_5041,N_4936,N_4948);
or U5042 (N_5042,N_4943,N_4933);
nand U5043 (N_5043,N_4971,N_4941);
or U5044 (N_5044,N_4977,N_4912);
or U5045 (N_5045,N_4976,N_4904);
xnor U5046 (N_5046,N_4910,N_4953);
or U5047 (N_5047,N_4997,N_4949);
nand U5048 (N_5048,N_4934,N_4992);
or U5049 (N_5049,N_4938,N_4957);
nand U5050 (N_5050,N_4904,N_4911);
or U5051 (N_5051,N_4973,N_4974);
or U5052 (N_5052,N_4918,N_4919);
nand U5053 (N_5053,N_4902,N_4980);
or U5054 (N_5054,N_4907,N_4917);
nor U5055 (N_5055,N_4992,N_4984);
and U5056 (N_5056,N_4965,N_4958);
or U5057 (N_5057,N_4980,N_4987);
nand U5058 (N_5058,N_4919,N_4936);
nor U5059 (N_5059,N_4926,N_4917);
or U5060 (N_5060,N_4991,N_4918);
and U5061 (N_5061,N_4998,N_4939);
and U5062 (N_5062,N_4994,N_4980);
nor U5063 (N_5063,N_4902,N_4977);
or U5064 (N_5064,N_4982,N_4919);
nor U5065 (N_5065,N_4975,N_4947);
xor U5066 (N_5066,N_4982,N_4905);
or U5067 (N_5067,N_4938,N_4966);
or U5068 (N_5068,N_4931,N_4943);
nor U5069 (N_5069,N_4911,N_4995);
or U5070 (N_5070,N_4963,N_4908);
and U5071 (N_5071,N_4934,N_4943);
and U5072 (N_5072,N_4978,N_4927);
nand U5073 (N_5073,N_4923,N_4977);
or U5074 (N_5074,N_4941,N_4997);
nor U5075 (N_5075,N_4926,N_4951);
and U5076 (N_5076,N_4906,N_4962);
and U5077 (N_5077,N_4910,N_4908);
nand U5078 (N_5078,N_4926,N_4979);
nor U5079 (N_5079,N_4901,N_4946);
nor U5080 (N_5080,N_4995,N_4947);
and U5081 (N_5081,N_4931,N_4994);
nor U5082 (N_5082,N_4921,N_4933);
nand U5083 (N_5083,N_4914,N_4916);
nand U5084 (N_5084,N_4987,N_4989);
and U5085 (N_5085,N_4958,N_4948);
xnor U5086 (N_5086,N_4981,N_4992);
or U5087 (N_5087,N_4942,N_4905);
and U5088 (N_5088,N_4964,N_4924);
or U5089 (N_5089,N_4990,N_4972);
nand U5090 (N_5090,N_4998,N_4978);
and U5091 (N_5091,N_4932,N_4931);
nor U5092 (N_5092,N_4997,N_4977);
nand U5093 (N_5093,N_4961,N_4939);
xnor U5094 (N_5094,N_4936,N_4929);
or U5095 (N_5095,N_4951,N_4999);
and U5096 (N_5096,N_4920,N_4944);
or U5097 (N_5097,N_4918,N_4915);
and U5098 (N_5098,N_4944,N_4926);
nand U5099 (N_5099,N_4964,N_4913);
nor U5100 (N_5100,N_5044,N_5083);
and U5101 (N_5101,N_5065,N_5006);
xor U5102 (N_5102,N_5096,N_5075);
or U5103 (N_5103,N_5073,N_5047);
nand U5104 (N_5104,N_5018,N_5068);
or U5105 (N_5105,N_5041,N_5021);
or U5106 (N_5106,N_5040,N_5059);
nor U5107 (N_5107,N_5055,N_5099);
nor U5108 (N_5108,N_5010,N_5048);
or U5109 (N_5109,N_5093,N_5060);
and U5110 (N_5110,N_5008,N_5042);
and U5111 (N_5111,N_5011,N_5032);
nor U5112 (N_5112,N_5023,N_5033);
xnor U5113 (N_5113,N_5038,N_5090);
nor U5114 (N_5114,N_5019,N_5081);
nor U5115 (N_5115,N_5017,N_5085);
or U5116 (N_5116,N_5094,N_5082);
nand U5117 (N_5117,N_5064,N_5031);
nand U5118 (N_5118,N_5098,N_5045);
nand U5119 (N_5119,N_5077,N_5028);
nand U5120 (N_5120,N_5052,N_5016);
nand U5121 (N_5121,N_5034,N_5062);
nor U5122 (N_5122,N_5080,N_5054);
nor U5123 (N_5123,N_5035,N_5097);
or U5124 (N_5124,N_5001,N_5087);
xnor U5125 (N_5125,N_5057,N_5004);
nand U5126 (N_5126,N_5029,N_5027);
nand U5127 (N_5127,N_5070,N_5092);
and U5128 (N_5128,N_5079,N_5022);
nor U5129 (N_5129,N_5037,N_5072);
or U5130 (N_5130,N_5078,N_5088);
or U5131 (N_5131,N_5061,N_5053);
or U5132 (N_5132,N_5046,N_5024);
and U5133 (N_5133,N_5013,N_5091);
nand U5134 (N_5134,N_5076,N_5084);
xor U5135 (N_5135,N_5074,N_5049);
and U5136 (N_5136,N_5030,N_5063);
and U5137 (N_5137,N_5095,N_5039);
and U5138 (N_5138,N_5007,N_5071);
or U5139 (N_5139,N_5003,N_5066);
and U5140 (N_5140,N_5086,N_5051);
or U5141 (N_5141,N_5020,N_5036);
nor U5142 (N_5142,N_5043,N_5005);
or U5143 (N_5143,N_5089,N_5000);
nand U5144 (N_5144,N_5002,N_5056);
nand U5145 (N_5145,N_5058,N_5069);
and U5146 (N_5146,N_5025,N_5050);
nand U5147 (N_5147,N_5026,N_5067);
or U5148 (N_5148,N_5015,N_5012);
nor U5149 (N_5149,N_5009,N_5014);
and U5150 (N_5150,N_5094,N_5021);
and U5151 (N_5151,N_5038,N_5019);
nor U5152 (N_5152,N_5099,N_5010);
nor U5153 (N_5153,N_5054,N_5077);
nor U5154 (N_5154,N_5001,N_5060);
or U5155 (N_5155,N_5051,N_5094);
nand U5156 (N_5156,N_5012,N_5059);
or U5157 (N_5157,N_5075,N_5065);
nor U5158 (N_5158,N_5054,N_5051);
or U5159 (N_5159,N_5030,N_5006);
nor U5160 (N_5160,N_5028,N_5020);
nor U5161 (N_5161,N_5007,N_5063);
and U5162 (N_5162,N_5002,N_5091);
or U5163 (N_5163,N_5041,N_5006);
and U5164 (N_5164,N_5078,N_5057);
and U5165 (N_5165,N_5075,N_5026);
and U5166 (N_5166,N_5013,N_5036);
nand U5167 (N_5167,N_5092,N_5020);
or U5168 (N_5168,N_5090,N_5058);
nand U5169 (N_5169,N_5025,N_5077);
or U5170 (N_5170,N_5031,N_5081);
nand U5171 (N_5171,N_5078,N_5028);
and U5172 (N_5172,N_5075,N_5015);
nor U5173 (N_5173,N_5010,N_5095);
nor U5174 (N_5174,N_5057,N_5009);
nor U5175 (N_5175,N_5088,N_5074);
nand U5176 (N_5176,N_5076,N_5050);
xor U5177 (N_5177,N_5075,N_5019);
and U5178 (N_5178,N_5081,N_5046);
nor U5179 (N_5179,N_5059,N_5096);
nor U5180 (N_5180,N_5043,N_5014);
nor U5181 (N_5181,N_5058,N_5027);
nor U5182 (N_5182,N_5068,N_5042);
nor U5183 (N_5183,N_5097,N_5063);
and U5184 (N_5184,N_5057,N_5014);
or U5185 (N_5185,N_5045,N_5070);
nand U5186 (N_5186,N_5019,N_5079);
xor U5187 (N_5187,N_5001,N_5065);
or U5188 (N_5188,N_5056,N_5018);
nor U5189 (N_5189,N_5061,N_5015);
and U5190 (N_5190,N_5095,N_5054);
nor U5191 (N_5191,N_5021,N_5086);
nand U5192 (N_5192,N_5037,N_5098);
nand U5193 (N_5193,N_5008,N_5076);
xnor U5194 (N_5194,N_5040,N_5058);
or U5195 (N_5195,N_5097,N_5099);
or U5196 (N_5196,N_5029,N_5096);
nor U5197 (N_5197,N_5040,N_5098);
and U5198 (N_5198,N_5073,N_5035);
or U5199 (N_5199,N_5091,N_5024);
nand U5200 (N_5200,N_5138,N_5135);
xnor U5201 (N_5201,N_5112,N_5175);
xor U5202 (N_5202,N_5182,N_5196);
or U5203 (N_5203,N_5194,N_5111);
or U5204 (N_5204,N_5103,N_5152);
and U5205 (N_5205,N_5173,N_5189);
nor U5206 (N_5206,N_5150,N_5113);
nand U5207 (N_5207,N_5123,N_5117);
or U5208 (N_5208,N_5100,N_5174);
or U5209 (N_5209,N_5153,N_5180);
and U5210 (N_5210,N_5129,N_5140);
and U5211 (N_5211,N_5118,N_5102);
and U5212 (N_5212,N_5158,N_5149);
nand U5213 (N_5213,N_5165,N_5162);
nor U5214 (N_5214,N_5166,N_5172);
or U5215 (N_5215,N_5198,N_5116);
xnor U5216 (N_5216,N_5107,N_5195);
or U5217 (N_5217,N_5147,N_5191);
nand U5218 (N_5218,N_5114,N_5197);
and U5219 (N_5219,N_5132,N_5125);
and U5220 (N_5220,N_5156,N_5109);
or U5221 (N_5221,N_5122,N_5168);
nor U5222 (N_5222,N_5130,N_5178);
nor U5223 (N_5223,N_5154,N_5142);
or U5224 (N_5224,N_5137,N_5139);
nand U5225 (N_5225,N_5101,N_5126);
nand U5226 (N_5226,N_5186,N_5144);
nand U5227 (N_5227,N_5185,N_5151);
and U5228 (N_5228,N_5167,N_5176);
or U5229 (N_5229,N_5192,N_5124);
xnor U5230 (N_5230,N_5105,N_5183);
nor U5231 (N_5231,N_5148,N_5187);
or U5232 (N_5232,N_5179,N_5155);
nand U5233 (N_5233,N_5120,N_5161);
nor U5234 (N_5234,N_5127,N_5121);
and U5235 (N_5235,N_5110,N_5108);
xnor U5236 (N_5236,N_5169,N_5119);
or U5237 (N_5237,N_5160,N_5131);
and U5238 (N_5238,N_5141,N_5134);
xor U5239 (N_5239,N_5163,N_5157);
or U5240 (N_5240,N_5104,N_5136);
and U5241 (N_5241,N_5181,N_5171);
or U5242 (N_5242,N_5164,N_5145);
or U5243 (N_5243,N_5133,N_5146);
and U5244 (N_5244,N_5199,N_5193);
nand U5245 (N_5245,N_5177,N_5170);
xnor U5246 (N_5246,N_5143,N_5188);
and U5247 (N_5247,N_5190,N_5159);
nand U5248 (N_5248,N_5184,N_5106);
nor U5249 (N_5249,N_5115,N_5128);
or U5250 (N_5250,N_5198,N_5187);
nand U5251 (N_5251,N_5107,N_5147);
or U5252 (N_5252,N_5192,N_5160);
and U5253 (N_5253,N_5111,N_5130);
or U5254 (N_5254,N_5172,N_5187);
nor U5255 (N_5255,N_5140,N_5174);
or U5256 (N_5256,N_5159,N_5109);
and U5257 (N_5257,N_5183,N_5122);
xor U5258 (N_5258,N_5128,N_5129);
or U5259 (N_5259,N_5192,N_5187);
nand U5260 (N_5260,N_5153,N_5106);
and U5261 (N_5261,N_5198,N_5163);
nand U5262 (N_5262,N_5175,N_5177);
or U5263 (N_5263,N_5161,N_5114);
and U5264 (N_5264,N_5125,N_5145);
nand U5265 (N_5265,N_5193,N_5180);
nand U5266 (N_5266,N_5188,N_5151);
nand U5267 (N_5267,N_5118,N_5180);
nor U5268 (N_5268,N_5110,N_5119);
and U5269 (N_5269,N_5123,N_5120);
and U5270 (N_5270,N_5197,N_5138);
xnor U5271 (N_5271,N_5133,N_5109);
and U5272 (N_5272,N_5153,N_5109);
or U5273 (N_5273,N_5192,N_5113);
and U5274 (N_5274,N_5169,N_5164);
xnor U5275 (N_5275,N_5135,N_5195);
nor U5276 (N_5276,N_5172,N_5131);
nor U5277 (N_5277,N_5171,N_5179);
nand U5278 (N_5278,N_5187,N_5167);
xnor U5279 (N_5279,N_5183,N_5148);
nor U5280 (N_5280,N_5184,N_5115);
and U5281 (N_5281,N_5166,N_5127);
and U5282 (N_5282,N_5111,N_5178);
and U5283 (N_5283,N_5140,N_5156);
or U5284 (N_5284,N_5152,N_5164);
or U5285 (N_5285,N_5101,N_5144);
or U5286 (N_5286,N_5188,N_5139);
nor U5287 (N_5287,N_5106,N_5122);
nor U5288 (N_5288,N_5187,N_5116);
nand U5289 (N_5289,N_5123,N_5102);
xor U5290 (N_5290,N_5108,N_5186);
or U5291 (N_5291,N_5135,N_5169);
or U5292 (N_5292,N_5117,N_5135);
or U5293 (N_5293,N_5191,N_5137);
nand U5294 (N_5294,N_5160,N_5196);
xnor U5295 (N_5295,N_5130,N_5102);
xor U5296 (N_5296,N_5149,N_5130);
and U5297 (N_5297,N_5150,N_5160);
and U5298 (N_5298,N_5113,N_5114);
xnor U5299 (N_5299,N_5112,N_5160);
nor U5300 (N_5300,N_5236,N_5255);
nand U5301 (N_5301,N_5215,N_5246);
xor U5302 (N_5302,N_5249,N_5222);
nor U5303 (N_5303,N_5290,N_5221);
or U5304 (N_5304,N_5228,N_5245);
nand U5305 (N_5305,N_5267,N_5227);
nand U5306 (N_5306,N_5217,N_5284);
nor U5307 (N_5307,N_5223,N_5293);
and U5308 (N_5308,N_5295,N_5209);
nor U5309 (N_5309,N_5212,N_5204);
or U5310 (N_5310,N_5272,N_5234);
nor U5311 (N_5311,N_5297,N_5211);
nor U5312 (N_5312,N_5260,N_5271);
and U5313 (N_5313,N_5216,N_5237);
nor U5314 (N_5314,N_5218,N_5273);
and U5315 (N_5315,N_5231,N_5241);
and U5316 (N_5316,N_5288,N_5263);
or U5317 (N_5317,N_5205,N_5282);
nand U5318 (N_5318,N_5250,N_5247);
xnor U5319 (N_5319,N_5213,N_5281);
nand U5320 (N_5320,N_5232,N_5278);
and U5321 (N_5321,N_5275,N_5240);
and U5322 (N_5322,N_5287,N_5226);
or U5323 (N_5323,N_5268,N_5252);
and U5324 (N_5324,N_5254,N_5279);
or U5325 (N_5325,N_5292,N_5266);
xor U5326 (N_5326,N_5283,N_5270);
nor U5327 (N_5327,N_5207,N_5276);
nand U5328 (N_5328,N_5208,N_5233);
nor U5329 (N_5329,N_5220,N_5265);
nor U5330 (N_5330,N_5235,N_5243);
or U5331 (N_5331,N_5294,N_5225);
nor U5332 (N_5332,N_5201,N_5248);
nor U5333 (N_5333,N_5229,N_5202);
or U5334 (N_5334,N_5230,N_5261);
and U5335 (N_5335,N_5291,N_5251);
nor U5336 (N_5336,N_5214,N_5203);
nor U5337 (N_5337,N_5206,N_5258);
nor U5338 (N_5338,N_5238,N_5224);
nor U5339 (N_5339,N_5253,N_5210);
and U5340 (N_5340,N_5296,N_5259);
or U5341 (N_5341,N_5274,N_5244);
or U5342 (N_5342,N_5242,N_5262);
nor U5343 (N_5343,N_5286,N_5299);
nand U5344 (N_5344,N_5257,N_5277);
and U5345 (N_5345,N_5219,N_5289);
xnor U5346 (N_5346,N_5269,N_5280);
and U5347 (N_5347,N_5285,N_5264);
or U5348 (N_5348,N_5298,N_5200);
or U5349 (N_5349,N_5239,N_5256);
and U5350 (N_5350,N_5261,N_5226);
nand U5351 (N_5351,N_5244,N_5277);
nand U5352 (N_5352,N_5217,N_5267);
nand U5353 (N_5353,N_5253,N_5205);
nand U5354 (N_5354,N_5297,N_5216);
or U5355 (N_5355,N_5287,N_5242);
nor U5356 (N_5356,N_5229,N_5287);
and U5357 (N_5357,N_5218,N_5204);
nand U5358 (N_5358,N_5260,N_5245);
xnor U5359 (N_5359,N_5244,N_5291);
nor U5360 (N_5360,N_5266,N_5240);
nand U5361 (N_5361,N_5204,N_5265);
or U5362 (N_5362,N_5207,N_5278);
nand U5363 (N_5363,N_5224,N_5292);
or U5364 (N_5364,N_5200,N_5280);
nor U5365 (N_5365,N_5203,N_5225);
or U5366 (N_5366,N_5270,N_5217);
or U5367 (N_5367,N_5297,N_5224);
or U5368 (N_5368,N_5231,N_5290);
or U5369 (N_5369,N_5285,N_5201);
or U5370 (N_5370,N_5292,N_5207);
and U5371 (N_5371,N_5298,N_5286);
xor U5372 (N_5372,N_5271,N_5220);
and U5373 (N_5373,N_5214,N_5253);
xor U5374 (N_5374,N_5254,N_5292);
nor U5375 (N_5375,N_5215,N_5256);
or U5376 (N_5376,N_5230,N_5259);
nor U5377 (N_5377,N_5210,N_5291);
nor U5378 (N_5378,N_5211,N_5283);
nor U5379 (N_5379,N_5295,N_5293);
nand U5380 (N_5380,N_5240,N_5282);
or U5381 (N_5381,N_5255,N_5220);
nand U5382 (N_5382,N_5242,N_5219);
and U5383 (N_5383,N_5216,N_5293);
nand U5384 (N_5384,N_5280,N_5294);
xor U5385 (N_5385,N_5287,N_5271);
and U5386 (N_5386,N_5236,N_5260);
or U5387 (N_5387,N_5203,N_5249);
nand U5388 (N_5388,N_5243,N_5251);
nand U5389 (N_5389,N_5262,N_5298);
and U5390 (N_5390,N_5214,N_5204);
xnor U5391 (N_5391,N_5255,N_5295);
or U5392 (N_5392,N_5220,N_5203);
or U5393 (N_5393,N_5210,N_5280);
nor U5394 (N_5394,N_5202,N_5251);
or U5395 (N_5395,N_5205,N_5256);
and U5396 (N_5396,N_5201,N_5292);
and U5397 (N_5397,N_5209,N_5270);
or U5398 (N_5398,N_5243,N_5234);
nand U5399 (N_5399,N_5211,N_5219);
and U5400 (N_5400,N_5337,N_5331);
xnor U5401 (N_5401,N_5381,N_5359);
xor U5402 (N_5402,N_5357,N_5374);
or U5403 (N_5403,N_5308,N_5365);
nor U5404 (N_5404,N_5378,N_5327);
nand U5405 (N_5405,N_5347,N_5305);
nor U5406 (N_5406,N_5349,N_5340);
nor U5407 (N_5407,N_5319,N_5313);
nand U5408 (N_5408,N_5363,N_5391);
nand U5409 (N_5409,N_5325,N_5335);
xnor U5410 (N_5410,N_5332,N_5302);
nor U5411 (N_5411,N_5330,N_5309);
nor U5412 (N_5412,N_5304,N_5338);
nor U5413 (N_5413,N_5360,N_5311);
or U5414 (N_5414,N_5315,N_5396);
or U5415 (N_5415,N_5326,N_5367);
nor U5416 (N_5416,N_5353,N_5352);
and U5417 (N_5417,N_5385,N_5393);
xnor U5418 (N_5418,N_5355,N_5377);
nand U5419 (N_5419,N_5371,N_5364);
nor U5420 (N_5420,N_5301,N_5379);
and U5421 (N_5421,N_5320,N_5376);
and U5422 (N_5422,N_5350,N_5390);
nor U5423 (N_5423,N_5399,N_5369);
or U5424 (N_5424,N_5346,N_5339);
or U5425 (N_5425,N_5310,N_5321);
nor U5426 (N_5426,N_5372,N_5384);
or U5427 (N_5427,N_5388,N_5345);
nor U5428 (N_5428,N_5375,N_5361);
and U5429 (N_5429,N_5317,N_5366);
and U5430 (N_5430,N_5322,N_5392);
or U5431 (N_5431,N_5336,N_5316);
and U5432 (N_5432,N_5387,N_5368);
xnor U5433 (N_5433,N_5358,N_5351);
nand U5434 (N_5434,N_5383,N_5300);
nor U5435 (N_5435,N_5323,N_5333);
nor U5436 (N_5436,N_5362,N_5354);
nor U5437 (N_5437,N_5324,N_5356);
or U5438 (N_5438,N_5307,N_5386);
and U5439 (N_5439,N_5348,N_5398);
or U5440 (N_5440,N_5303,N_5373);
nor U5441 (N_5441,N_5312,N_5314);
or U5442 (N_5442,N_5343,N_5382);
or U5443 (N_5443,N_5380,N_5344);
xor U5444 (N_5444,N_5318,N_5394);
or U5445 (N_5445,N_5329,N_5397);
nor U5446 (N_5446,N_5389,N_5306);
nor U5447 (N_5447,N_5341,N_5342);
and U5448 (N_5448,N_5328,N_5370);
xnor U5449 (N_5449,N_5395,N_5334);
or U5450 (N_5450,N_5351,N_5312);
nand U5451 (N_5451,N_5351,N_5313);
and U5452 (N_5452,N_5372,N_5393);
nand U5453 (N_5453,N_5397,N_5367);
or U5454 (N_5454,N_5320,N_5305);
nand U5455 (N_5455,N_5306,N_5397);
nor U5456 (N_5456,N_5313,N_5393);
nand U5457 (N_5457,N_5330,N_5354);
nor U5458 (N_5458,N_5301,N_5325);
nor U5459 (N_5459,N_5335,N_5381);
and U5460 (N_5460,N_5328,N_5386);
xor U5461 (N_5461,N_5346,N_5356);
nand U5462 (N_5462,N_5355,N_5334);
nand U5463 (N_5463,N_5352,N_5364);
xnor U5464 (N_5464,N_5329,N_5309);
nor U5465 (N_5465,N_5301,N_5375);
or U5466 (N_5466,N_5357,N_5392);
xnor U5467 (N_5467,N_5381,N_5372);
and U5468 (N_5468,N_5391,N_5312);
and U5469 (N_5469,N_5366,N_5362);
nor U5470 (N_5470,N_5360,N_5340);
nor U5471 (N_5471,N_5365,N_5396);
and U5472 (N_5472,N_5356,N_5313);
or U5473 (N_5473,N_5363,N_5336);
nor U5474 (N_5474,N_5308,N_5319);
or U5475 (N_5475,N_5396,N_5355);
and U5476 (N_5476,N_5300,N_5325);
or U5477 (N_5477,N_5394,N_5351);
nand U5478 (N_5478,N_5328,N_5394);
nand U5479 (N_5479,N_5351,N_5306);
nand U5480 (N_5480,N_5336,N_5398);
and U5481 (N_5481,N_5390,N_5398);
or U5482 (N_5482,N_5349,N_5348);
and U5483 (N_5483,N_5313,N_5324);
and U5484 (N_5484,N_5313,N_5348);
nor U5485 (N_5485,N_5361,N_5386);
nand U5486 (N_5486,N_5377,N_5382);
nor U5487 (N_5487,N_5331,N_5338);
or U5488 (N_5488,N_5300,N_5333);
nor U5489 (N_5489,N_5335,N_5307);
or U5490 (N_5490,N_5339,N_5394);
and U5491 (N_5491,N_5370,N_5389);
and U5492 (N_5492,N_5381,N_5338);
or U5493 (N_5493,N_5342,N_5344);
nand U5494 (N_5494,N_5357,N_5315);
nand U5495 (N_5495,N_5313,N_5328);
nand U5496 (N_5496,N_5369,N_5371);
and U5497 (N_5497,N_5353,N_5357);
xor U5498 (N_5498,N_5363,N_5384);
nand U5499 (N_5499,N_5378,N_5394);
and U5500 (N_5500,N_5408,N_5460);
or U5501 (N_5501,N_5406,N_5447);
nor U5502 (N_5502,N_5400,N_5402);
and U5503 (N_5503,N_5457,N_5473);
nand U5504 (N_5504,N_5441,N_5498);
and U5505 (N_5505,N_5428,N_5465);
and U5506 (N_5506,N_5418,N_5421);
xnor U5507 (N_5507,N_5442,N_5467);
and U5508 (N_5508,N_5464,N_5476);
xnor U5509 (N_5509,N_5492,N_5490);
and U5510 (N_5510,N_5471,N_5401);
or U5511 (N_5511,N_5416,N_5444);
or U5512 (N_5512,N_5485,N_5452);
nor U5513 (N_5513,N_5413,N_5474);
nor U5514 (N_5514,N_5431,N_5432);
nor U5515 (N_5515,N_5411,N_5445);
and U5516 (N_5516,N_5463,N_5427);
and U5517 (N_5517,N_5494,N_5412);
nand U5518 (N_5518,N_5440,N_5420);
xnor U5519 (N_5519,N_5486,N_5491);
nand U5520 (N_5520,N_5497,N_5433);
nand U5521 (N_5521,N_5468,N_5438);
or U5522 (N_5522,N_5478,N_5407);
nand U5523 (N_5523,N_5435,N_5493);
nor U5524 (N_5524,N_5458,N_5422);
nand U5525 (N_5525,N_5403,N_5410);
nor U5526 (N_5526,N_5415,N_5488);
and U5527 (N_5527,N_5429,N_5450);
nor U5528 (N_5528,N_5414,N_5462);
nand U5529 (N_5529,N_5472,N_5453);
nor U5530 (N_5530,N_5417,N_5482);
nand U5531 (N_5531,N_5499,N_5459);
and U5532 (N_5532,N_5484,N_5404);
nor U5533 (N_5533,N_5443,N_5430);
nand U5534 (N_5534,N_5446,N_5454);
or U5535 (N_5535,N_5461,N_5469);
nand U5536 (N_5536,N_5423,N_5425);
and U5537 (N_5537,N_5405,N_5449);
or U5538 (N_5538,N_5437,N_5455);
nor U5539 (N_5539,N_5496,N_5489);
nor U5540 (N_5540,N_5487,N_5477);
or U5541 (N_5541,N_5436,N_5466);
nor U5542 (N_5542,N_5481,N_5448);
or U5543 (N_5543,N_5426,N_5424);
nor U5544 (N_5544,N_5480,N_5483);
nand U5545 (N_5545,N_5419,N_5456);
nor U5546 (N_5546,N_5409,N_5495);
and U5547 (N_5547,N_5434,N_5475);
nor U5548 (N_5548,N_5479,N_5451);
nor U5549 (N_5549,N_5470,N_5439);
nand U5550 (N_5550,N_5485,N_5460);
nand U5551 (N_5551,N_5496,N_5477);
and U5552 (N_5552,N_5407,N_5425);
and U5553 (N_5553,N_5412,N_5438);
or U5554 (N_5554,N_5489,N_5411);
and U5555 (N_5555,N_5432,N_5402);
nand U5556 (N_5556,N_5437,N_5432);
nor U5557 (N_5557,N_5459,N_5407);
nand U5558 (N_5558,N_5448,N_5465);
or U5559 (N_5559,N_5460,N_5438);
and U5560 (N_5560,N_5481,N_5449);
nor U5561 (N_5561,N_5462,N_5433);
or U5562 (N_5562,N_5442,N_5423);
and U5563 (N_5563,N_5456,N_5408);
nand U5564 (N_5564,N_5486,N_5482);
and U5565 (N_5565,N_5447,N_5486);
xnor U5566 (N_5566,N_5487,N_5402);
and U5567 (N_5567,N_5452,N_5444);
nor U5568 (N_5568,N_5485,N_5499);
xor U5569 (N_5569,N_5449,N_5416);
nor U5570 (N_5570,N_5433,N_5485);
and U5571 (N_5571,N_5433,N_5404);
nand U5572 (N_5572,N_5480,N_5489);
nor U5573 (N_5573,N_5438,N_5481);
nor U5574 (N_5574,N_5429,N_5495);
nor U5575 (N_5575,N_5458,N_5402);
and U5576 (N_5576,N_5470,N_5459);
xor U5577 (N_5577,N_5423,N_5430);
nor U5578 (N_5578,N_5459,N_5490);
nand U5579 (N_5579,N_5496,N_5465);
and U5580 (N_5580,N_5473,N_5436);
or U5581 (N_5581,N_5403,N_5402);
nand U5582 (N_5582,N_5470,N_5408);
and U5583 (N_5583,N_5474,N_5412);
xnor U5584 (N_5584,N_5404,N_5451);
or U5585 (N_5585,N_5445,N_5418);
and U5586 (N_5586,N_5452,N_5401);
nand U5587 (N_5587,N_5476,N_5470);
and U5588 (N_5588,N_5491,N_5496);
nor U5589 (N_5589,N_5484,N_5453);
and U5590 (N_5590,N_5431,N_5420);
nand U5591 (N_5591,N_5448,N_5450);
xor U5592 (N_5592,N_5480,N_5460);
and U5593 (N_5593,N_5448,N_5447);
nor U5594 (N_5594,N_5491,N_5411);
nor U5595 (N_5595,N_5470,N_5449);
nor U5596 (N_5596,N_5429,N_5465);
and U5597 (N_5597,N_5423,N_5447);
and U5598 (N_5598,N_5415,N_5412);
xor U5599 (N_5599,N_5440,N_5436);
or U5600 (N_5600,N_5565,N_5510);
nand U5601 (N_5601,N_5593,N_5511);
or U5602 (N_5602,N_5556,N_5529);
or U5603 (N_5603,N_5516,N_5591);
nor U5604 (N_5604,N_5544,N_5595);
nor U5605 (N_5605,N_5520,N_5584);
nor U5606 (N_5606,N_5522,N_5555);
and U5607 (N_5607,N_5585,N_5501);
nor U5608 (N_5608,N_5559,N_5535);
and U5609 (N_5609,N_5581,N_5503);
or U5610 (N_5610,N_5509,N_5539);
xnor U5611 (N_5611,N_5517,N_5596);
nor U5612 (N_5612,N_5580,N_5571);
nor U5613 (N_5613,N_5527,N_5572);
nor U5614 (N_5614,N_5548,N_5545);
and U5615 (N_5615,N_5518,N_5582);
nor U5616 (N_5616,N_5576,N_5579);
or U5617 (N_5617,N_5505,N_5549);
or U5618 (N_5618,N_5590,N_5570);
nand U5619 (N_5619,N_5553,N_5563);
nand U5620 (N_5620,N_5546,N_5534);
nor U5621 (N_5621,N_5561,N_5514);
xnor U5622 (N_5622,N_5562,N_5554);
nand U5623 (N_5623,N_5575,N_5526);
xnor U5624 (N_5624,N_5574,N_5543);
or U5625 (N_5625,N_5524,N_5531);
or U5626 (N_5626,N_5500,N_5557);
or U5627 (N_5627,N_5564,N_5541);
and U5628 (N_5628,N_5504,N_5578);
nor U5629 (N_5629,N_5512,N_5550);
nor U5630 (N_5630,N_5599,N_5530);
and U5631 (N_5631,N_5587,N_5519);
and U5632 (N_5632,N_5506,N_5589);
nand U5633 (N_5633,N_5558,N_5597);
nor U5634 (N_5634,N_5568,N_5540);
or U5635 (N_5635,N_5538,N_5586);
nor U5636 (N_5636,N_5573,N_5502);
nand U5637 (N_5637,N_5569,N_5537);
and U5638 (N_5638,N_5532,N_5598);
or U5639 (N_5639,N_5507,N_5525);
nand U5640 (N_5640,N_5588,N_5594);
nor U5641 (N_5641,N_5560,N_5521);
nand U5642 (N_5642,N_5547,N_5528);
or U5643 (N_5643,N_5577,N_5552);
nor U5644 (N_5644,N_5583,N_5592);
xnor U5645 (N_5645,N_5523,N_5551);
or U5646 (N_5646,N_5513,N_5515);
nand U5647 (N_5647,N_5567,N_5508);
or U5648 (N_5648,N_5542,N_5536);
nand U5649 (N_5649,N_5533,N_5566);
nor U5650 (N_5650,N_5552,N_5583);
and U5651 (N_5651,N_5589,N_5562);
or U5652 (N_5652,N_5534,N_5598);
nand U5653 (N_5653,N_5570,N_5502);
nor U5654 (N_5654,N_5583,N_5570);
nor U5655 (N_5655,N_5534,N_5541);
nand U5656 (N_5656,N_5561,N_5556);
and U5657 (N_5657,N_5591,N_5559);
or U5658 (N_5658,N_5519,N_5500);
nand U5659 (N_5659,N_5507,N_5563);
and U5660 (N_5660,N_5508,N_5591);
or U5661 (N_5661,N_5565,N_5561);
nor U5662 (N_5662,N_5505,N_5532);
nand U5663 (N_5663,N_5544,N_5579);
or U5664 (N_5664,N_5543,N_5591);
xnor U5665 (N_5665,N_5598,N_5585);
nand U5666 (N_5666,N_5598,N_5595);
or U5667 (N_5667,N_5512,N_5564);
or U5668 (N_5668,N_5584,N_5531);
and U5669 (N_5669,N_5585,N_5595);
and U5670 (N_5670,N_5535,N_5527);
xnor U5671 (N_5671,N_5577,N_5593);
nand U5672 (N_5672,N_5522,N_5533);
nand U5673 (N_5673,N_5526,N_5586);
and U5674 (N_5674,N_5508,N_5507);
and U5675 (N_5675,N_5523,N_5518);
nand U5676 (N_5676,N_5573,N_5594);
or U5677 (N_5677,N_5544,N_5505);
and U5678 (N_5678,N_5530,N_5525);
nand U5679 (N_5679,N_5538,N_5529);
and U5680 (N_5680,N_5507,N_5565);
nand U5681 (N_5681,N_5579,N_5523);
nor U5682 (N_5682,N_5526,N_5500);
xor U5683 (N_5683,N_5542,N_5558);
nor U5684 (N_5684,N_5546,N_5539);
or U5685 (N_5685,N_5595,N_5516);
xnor U5686 (N_5686,N_5525,N_5543);
nor U5687 (N_5687,N_5551,N_5563);
nor U5688 (N_5688,N_5549,N_5577);
or U5689 (N_5689,N_5566,N_5512);
or U5690 (N_5690,N_5577,N_5568);
nor U5691 (N_5691,N_5570,N_5531);
or U5692 (N_5692,N_5575,N_5501);
xnor U5693 (N_5693,N_5550,N_5507);
or U5694 (N_5694,N_5577,N_5534);
and U5695 (N_5695,N_5500,N_5510);
nor U5696 (N_5696,N_5555,N_5584);
xnor U5697 (N_5697,N_5549,N_5580);
nor U5698 (N_5698,N_5580,N_5598);
and U5699 (N_5699,N_5580,N_5577);
or U5700 (N_5700,N_5655,N_5603);
and U5701 (N_5701,N_5629,N_5647);
nor U5702 (N_5702,N_5638,N_5685);
nand U5703 (N_5703,N_5618,N_5632);
nor U5704 (N_5704,N_5696,N_5621);
nor U5705 (N_5705,N_5658,N_5608);
nand U5706 (N_5706,N_5690,N_5606);
and U5707 (N_5707,N_5630,N_5668);
nand U5708 (N_5708,N_5692,N_5631);
and U5709 (N_5709,N_5648,N_5610);
nand U5710 (N_5710,N_5677,N_5625);
nand U5711 (N_5711,N_5612,N_5669);
nor U5712 (N_5712,N_5626,N_5649);
and U5713 (N_5713,N_5661,N_5650);
nand U5714 (N_5714,N_5682,N_5611);
nand U5715 (N_5715,N_5665,N_5673);
nand U5716 (N_5716,N_5688,N_5693);
nand U5717 (N_5717,N_5604,N_5678);
nand U5718 (N_5718,N_5634,N_5637);
nand U5719 (N_5719,N_5623,N_5664);
nor U5720 (N_5720,N_5691,N_5662);
nor U5721 (N_5721,N_5635,N_5651);
nor U5722 (N_5722,N_5657,N_5666);
xnor U5723 (N_5723,N_5689,N_5699);
nand U5724 (N_5724,N_5694,N_5656);
nand U5725 (N_5725,N_5601,N_5641);
and U5726 (N_5726,N_5679,N_5659);
nand U5727 (N_5727,N_5663,N_5617);
or U5728 (N_5728,N_5633,N_5680);
or U5729 (N_5729,N_5695,N_5640);
nand U5730 (N_5730,N_5642,N_5674);
and U5731 (N_5731,N_5686,N_5698);
nand U5732 (N_5732,N_5675,N_5654);
nor U5733 (N_5733,N_5602,N_5667);
nand U5734 (N_5734,N_5643,N_5660);
or U5735 (N_5735,N_5672,N_5622);
nor U5736 (N_5736,N_5687,N_5607);
or U5737 (N_5737,N_5609,N_5670);
and U5738 (N_5738,N_5628,N_5624);
and U5739 (N_5739,N_5620,N_5613);
and U5740 (N_5740,N_5653,N_5615);
nand U5741 (N_5741,N_5676,N_5646);
and U5742 (N_5742,N_5697,N_5600);
nor U5743 (N_5743,N_5645,N_5652);
xor U5744 (N_5744,N_5616,N_5636);
nand U5745 (N_5745,N_5614,N_5681);
nor U5746 (N_5746,N_5627,N_5639);
or U5747 (N_5747,N_5619,N_5671);
nor U5748 (N_5748,N_5683,N_5684);
nor U5749 (N_5749,N_5644,N_5605);
and U5750 (N_5750,N_5682,N_5681);
or U5751 (N_5751,N_5602,N_5675);
nor U5752 (N_5752,N_5678,N_5613);
nand U5753 (N_5753,N_5618,N_5613);
nand U5754 (N_5754,N_5645,N_5677);
or U5755 (N_5755,N_5691,N_5664);
and U5756 (N_5756,N_5601,N_5669);
nand U5757 (N_5757,N_5673,N_5629);
nand U5758 (N_5758,N_5694,N_5621);
or U5759 (N_5759,N_5698,N_5643);
or U5760 (N_5760,N_5694,N_5652);
and U5761 (N_5761,N_5643,N_5640);
xnor U5762 (N_5762,N_5664,N_5642);
nand U5763 (N_5763,N_5680,N_5649);
nor U5764 (N_5764,N_5626,N_5688);
nor U5765 (N_5765,N_5620,N_5689);
nor U5766 (N_5766,N_5669,N_5693);
nor U5767 (N_5767,N_5600,N_5688);
or U5768 (N_5768,N_5693,N_5664);
xor U5769 (N_5769,N_5613,N_5671);
nor U5770 (N_5770,N_5651,N_5650);
or U5771 (N_5771,N_5653,N_5683);
nand U5772 (N_5772,N_5686,N_5622);
or U5773 (N_5773,N_5634,N_5697);
xor U5774 (N_5774,N_5630,N_5635);
or U5775 (N_5775,N_5630,N_5658);
nor U5776 (N_5776,N_5689,N_5692);
or U5777 (N_5777,N_5666,N_5608);
nand U5778 (N_5778,N_5661,N_5655);
or U5779 (N_5779,N_5665,N_5682);
or U5780 (N_5780,N_5610,N_5631);
nor U5781 (N_5781,N_5644,N_5676);
and U5782 (N_5782,N_5625,N_5624);
xor U5783 (N_5783,N_5674,N_5694);
nor U5784 (N_5784,N_5676,N_5620);
nand U5785 (N_5785,N_5641,N_5626);
nor U5786 (N_5786,N_5659,N_5611);
nor U5787 (N_5787,N_5671,N_5636);
or U5788 (N_5788,N_5675,N_5659);
nand U5789 (N_5789,N_5661,N_5620);
xor U5790 (N_5790,N_5611,N_5689);
and U5791 (N_5791,N_5631,N_5633);
or U5792 (N_5792,N_5663,N_5695);
nand U5793 (N_5793,N_5637,N_5628);
or U5794 (N_5794,N_5627,N_5652);
or U5795 (N_5795,N_5639,N_5601);
nand U5796 (N_5796,N_5648,N_5639);
or U5797 (N_5797,N_5697,N_5667);
or U5798 (N_5798,N_5631,N_5678);
and U5799 (N_5799,N_5689,N_5639);
nor U5800 (N_5800,N_5783,N_5773);
or U5801 (N_5801,N_5709,N_5763);
nor U5802 (N_5802,N_5727,N_5721);
or U5803 (N_5803,N_5719,N_5715);
nand U5804 (N_5804,N_5718,N_5716);
nand U5805 (N_5805,N_5778,N_5729);
or U5806 (N_5806,N_5785,N_5758);
nand U5807 (N_5807,N_5701,N_5752);
or U5808 (N_5808,N_5775,N_5741);
and U5809 (N_5809,N_5734,N_5789);
nor U5810 (N_5810,N_5708,N_5743);
nand U5811 (N_5811,N_5792,N_5740);
nand U5812 (N_5812,N_5714,N_5705);
nand U5813 (N_5813,N_5761,N_5787);
or U5814 (N_5814,N_5760,N_5796);
nor U5815 (N_5815,N_5764,N_5755);
xor U5816 (N_5816,N_5711,N_5745);
nor U5817 (N_5817,N_5756,N_5724);
and U5818 (N_5818,N_5777,N_5725);
xnor U5819 (N_5819,N_5704,N_5742);
or U5820 (N_5820,N_5768,N_5780);
and U5821 (N_5821,N_5784,N_5791);
xnor U5822 (N_5822,N_5772,N_5757);
and U5823 (N_5823,N_5736,N_5748);
nand U5824 (N_5824,N_5767,N_5774);
nand U5825 (N_5825,N_5703,N_5735);
nand U5826 (N_5826,N_5788,N_5790);
xor U5827 (N_5827,N_5733,N_5749);
and U5828 (N_5828,N_5726,N_5720);
and U5829 (N_5829,N_5759,N_5712);
and U5830 (N_5830,N_5751,N_5707);
and U5831 (N_5831,N_5771,N_5770);
nand U5832 (N_5832,N_5779,N_5738);
nor U5833 (N_5833,N_5753,N_5744);
or U5834 (N_5834,N_5739,N_5766);
nand U5835 (N_5835,N_5737,N_5776);
or U5836 (N_5836,N_5794,N_5798);
nor U5837 (N_5837,N_5713,N_5702);
nor U5838 (N_5838,N_5795,N_5730);
nor U5839 (N_5839,N_5710,N_5728);
nor U5840 (N_5840,N_5722,N_5762);
nand U5841 (N_5841,N_5723,N_5706);
nand U5842 (N_5842,N_5781,N_5799);
or U5843 (N_5843,N_5700,N_5717);
nand U5844 (N_5844,N_5786,N_5732);
nand U5845 (N_5845,N_5731,N_5750);
nor U5846 (N_5846,N_5793,N_5769);
or U5847 (N_5847,N_5765,N_5747);
nand U5848 (N_5848,N_5754,N_5746);
nor U5849 (N_5849,N_5797,N_5782);
and U5850 (N_5850,N_5756,N_5723);
or U5851 (N_5851,N_5722,N_5707);
and U5852 (N_5852,N_5740,N_5744);
or U5853 (N_5853,N_5782,N_5769);
xor U5854 (N_5854,N_5700,N_5737);
or U5855 (N_5855,N_5771,N_5765);
nand U5856 (N_5856,N_5709,N_5755);
and U5857 (N_5857,N_5774,N_5726);
nor U5858 (N_5858,N_5720,N_5779);
nor U5859 (N_5859,N_5794,N_5736);
nor U5860 (N_5860,N_5735,N_5720);
or U5861 (N_5861,N_5773,N_5722);
and U5862 (N_5862,N_5786,N_5775);
nor U5863 (N_5863,N_5763,N_5743);
nand U5864 (N_5864,N_5767,N_5795);
nand U5865 (N_5865,N_5749,N_5767);
nand U5866 (N_5866,N_5719,N_5791);
xnor U5867 (N_5867,N_5745,N_5751);
nor U5868 (N_5868,N_5736,N_5732);
nor U5869 (N_5869,N_5782,N_5733);
and U5870 (N_5870,N_5738,N_5739);
nor U5871 (N_5871,N_5739,N_5743);
nand U5872 (N_5872,N_5795,N_5785);
or U5873 (N_5873,N_5730,N_5735);
xnor U5874 (N_5874,N_5797,N_5783);
and U5875 (N_5875,N_5747,N_5795);
and U5876 (N_5876,N_5751,N_5767);
or U5877 (N_5877,N_5727,N_5735);
and U5878 (N_5878,N_5791,N_5757);
xnor U5879 (N_5879,N_5782,N_5766);
or U5880 (N_5880,N_5795,N_5798);
nand U5881 (N_5881,N_5703,N_5736);
or U5882 (N_5882,N_5715,N_5748);
nor U5883 (N_5883,N_5744,N_5737);
nand U5884 (N_5884,N_5775,N_5748);
or U5885 (N_5885,N_5757,N_5748);
nand U5886 (N_5886,N_5780,N_5762);
or U5887 (N_5887,N_5777,N_5724);
and U5888 (N_5888,N_5700,N_5769);
and U5889 (N_5889,N_5720,N_5743);
nand U5890 (N_5890,N_5778,N_5734);
or U5891 (N_5891,N_5713,N_5708);
xnor U5892 (N_5892,N_5732,N_5739);
or U5893 (N_5893,N_5718,N_5709);
and U5894 (N_5894,N_5721,N_5778);
and U5895 (N_5895,N_5783,N_5718);
and U5896 (N_5896,N_5795,N_5759);
and U5897 (N_5897,N_5753,N_5797);
or U5898 (N_5898,N_5754,N_5744);
nand U5899 (N_5899,N_5789,N_5771);
and U5900 (N_5900,N_5889,N_5848);
or U5901 (N_5901,N_5808,N_5845);
nand U5902 (N_5902,N_5873,N_5829);
nor U5903 (N_5903,N_5811,N_5804);
or U5904 (N_5904,N_5896,N_5813);
nand U5905 (N_5905,N_5898,N_5865);
or U5906 (N_5906,N_5840,N_5823);
and U5907 (N_5907,N_5876,N_5849);
nand U5908 (N_5908,N_5884,N_5836);
or U5909 (N_5909,N_5844,N_5872);
nand U5910 (N_5910,N_5824,N_5892);
or U5911 (N_5911,N_5877,N_5886);
nor U5912 (N_5912,N_5837,N_5891);
nand U5913 (N_5913,N_5821,N_5838);
nor U5914 (N_5914,N_5828,N_5825);
nor U5915 (N_5915,N_5893,N_5846);
and U5916 (N_5916,N_5858,N_5875);
and U5917 (N_5917,N_5806,N_5860);
and U5918 (N_5918,N_5810,N_5812);
or U5919 (N_5919,N_5887,N_5835);
and U5920 (N_5920,N_5850,N_5847);
nand U5921 (N_5921,N_5897,N_5874);
nor U5922 (N_5922,N_5853,N_5899);
xnor U5923 (N_5923,N_5816,N_5834);
nor U5924 (N_5924,N_5843,N_5805);
and U5925 (N_5925,N_5832,N_5826);
or U5926 (N_5926,N_5862,N_5841);
or U5927 (N_5927,N_5807,N_5867);
xor U5928 (N_5928,N_5815,N_5868);
or U5929 (N_5929,N_5883,N_5861);
or U5930 (N_5930,N_5851,N_5819);
nor U5931 (N_5931,N_5856,N_5839);
nor U5932 (N_5932,N_5820,N_5830);
nand U5933 (N_5933,N_5833,N_5880);
and U5934 (N_5934,N_5818,N_5817);
nor U5935 (N_5935,N_5800,N_5885);
and U5936 (N_5936,N_5801,N_5803);
nand U5937 (N_5937,N_5831,N_5802);
and U5938 (N_5938,N_5870,N_5888);
nand U5939 (N_5939,N_5882,N_5895);
and U5940 (N_5940,N_5890,N_5852);
and U5941 (N_5941,N_5871,N_5855);
nor U5942 (N_5942,N_5827,N_5866);
or U5943 (N_5943,N_5822,N_5842);
nor U5944 (N_5944,N_5869,N_5881);
or U5945 (N_5945,N_5854,N_5859);
and U5946 (N_5946,N_5863,N_5879);
nand U5947 (N_5947,N_5814,N_5857);
nand U5948 (N_5948,N_5864,N_5894);
nor U5949 (N_5949,N_5809,N_5878);
nor U5950 (N_5950,N_5876,N_5840);
nor U5951 (N_5951,N_5832,N_5858);
or U5952 (N_5952,N_5812,N_5856);
nand U5953 (N_5953,N_5825,N_5884);
or U5954 (N_5954,N_5810,N_5839);
or U5955 (N_5955,N_5812,N_5825);
and U5956 (N_5956,N_5818,N_5833);
and U5957 (N_5957,N_5812,N_5898);
nand U5958 (N_5958,N_5874,N_5840);
nor U5959 (N_5959,N_5873,N_5864);
or U5960 (N_5960,N_5805,N_5862);
nand U5961 (N_5961,N_5869,N_5802);
and U5962 (N_5962,N_5825,N_5800);
and U5963 (N_5963,N_5897,N_5846);
nand U5964 (N_5964,N_5859,N_5895);
and U5965 (N_5965,N_5886,N_5830);
and U5966 (N_5966,N_5865,N_5874);
and U5967 (N_5967,N_5898,N_5855);
xnor U5968 (N_5968,N_5852,N_5872);
and U5969 (N_5969,N_5845,N_5802);
nand U5970 (N_5970,N_5861,N_5847);
nor U5971 (N_5971,N_5871,N_5836);
nand U5972 (N_5972,N_5835,N_5871);
nor U5973 (N_5973,N_5876,N_5804);
or U5974 (N_5974,N_5857,N_5856);
and U5975 (N_5975,N_5871,N_5890);
xnor U5976 (N_5976,N_5825,N_5861);
and U5977 (N_5977,N_5860,N_5819);
or U5978 (N_5978,N_5811,N_5864);
nor U5979 (N_5979,N_5877,N_5818);
nor U5980 (N_5980,N_5834,N_5862);
or U5981 (N_5981,N_5894,N_5800);
or U5982 (N_5982,N_5836,N_5856);
or U5983 (N_5983,N_5839,N_5804);
and U5984 (N_5984,N_5816,N_5870);
nand U5985 (N_5985,N_5888,N_5860);
or U5986 (N_5986,N_5886,N_5810);
xor U5987 (N_5987,N_5871,N_5898);
or U5988 (N_5988,N_5812,N_5822);
nor U5989 (N_5989,N_5863,N_5857);
or U5990 (N_5990,N_5858,N_5855);
nor U5991 (N_5991,N_5873,N_5825);
or U5992 (N_5992,N_5869,N_5837);
or U5993 (N_5993,N_5867,N_5802);
xor U5994 (N_5994,N_5807,N_5808);
nand U5995 (N_5995,N_5875,N_5882);
nand U5996 (N_5996,N_5824,N_5835);
nor U5997 (N_5997,N_5852,N_5813);
xor U5998 (N_5998,N_5807,N_5869);
or U5999 (N_5999,N_5885,N_5817);
xnor U6000 (N_6000,N_5930,N_5918);
nor U6001 (N_6001,N_5905,N_5965);
nor U6002 (N_6002,N_5944,N_5984);
or U6003 (N_6003,N_5921,N_5909);
or U6004 (N_6004,N_5995,N_5939);
or U6005 (N_6005,N_5949,N_5912);
nand U6006 (N_6006,N_5997,N_5989);
and U6007 (N_6007,N_5910,N_5928);
and U6008 (N_6008,N_5968,N_5991);
or U6009 (N_6009,N_5990,N_5996);
nand U6010 (N_6010,N_5943,N_5938);
nor U6011 (N_6011,N_5941,N_5994);
nor U6012 (N_6012,N_5957,N_5926);
nand U6013 (N_6013,N_5919,N_5931);
nor U6014 (N_6014,N_5967,N_5988);
and U6015 (N_6015,N_5987,N_5973);
xor U6016 (N_6016,N_5917,N_5974);
xnor U6017 (N_6017,N_5915,N_5908);
and U6018 (N_6018,N_5986,N_5954);
and U6019 (N_6019,N_5972,N_5964);
nor U6020 (N_6020,N_5950,N_5947);
or U6021 (N_6021,N_5907,N_5992);
nor U6022 (N_6022,N_5927,N_5937);
nor U6023 (N_6023,N_5911,N_5904);
nand U6024 (N_6024,N_5906,N_5951);
nor U6025 (N_6025,N_5955,N_5932);
and U6026 (N_6026,N_5923,N_5913);
nor U6027 (N_6027,N_5922,N_5936);
nand U6028 (N_6028,N_5958,N_5916);
and U6029 (N_6029,N_5981,N_5975);
nand U6030 (N_6030,N_5977,N_5960);
or U6031 (N_6031,N_5948,N_5980);
or U6032 (N_6032,N_5985,N_5946);
nand U6033 (N_6033,N_5982,N_5933);
and U6034 (N_6034,N_5962,N_5993);
and U6035 (N_6035,N_5966,N_5983);
xor U6036 (N_6036,N_5998,N_5935);
or U6037 (N_6037,N_5999,N_5942);
xnor U6038 (N_6038,N_5929,N_5920);
xor U6039 (N_6039,N_5961,N_5976);
and U6040 (N_6040,N_5945,N_5924);
nor U6041 (N_6041,N_5901,N_5969);
and U6042 (N_6042,N_5925,N_5978);
nand U6043 (N_6043,N_5956,N_5959);
nand U6044 (N_6044,N_5914,N_5952);
or U6045 (N_6045,N_5979,N_5900);
or U6046 (N_6046,N_5963,N_5970);
nand U6047 (N_6047,N_5971,N_5902);
nand U6048 (N_6048,N_5903,N_5934);
nand U6049 (N_6049,N_5953,N_5940);
nor U6050 (N_6050,N_5953,N_5948);
or U6051 (N_6051,N_5926,N_5960);
xor U6052 (N_6052,N_5946,N_5940);
nand U6053 (N_6053,N_5997,N_5908);
nand U6054 (N_6054,N_5994,N_5972);
and U6055 (N_6055,N_5959,N_5994);
xnor U6056 (N_6056,N_5952,N_5925);
or U6057 (N_6057,N_5975,N_5967);
or U6058 (N_6058,N_5941,N_5912);
or U6059 (N_6059,N_5937,N_5979);
xor U6060 (N_6060,N_5911,N_5914);
or U6061 (N_6061,N_5957,N_5969);
or U6062 (N_6062,N_5955,N_5913);
and U6063 (N_6063,N_5950,N_5992);
nor U6064 (N_6064,N_5908,N_5942);
nor U6065 (N_6065,N_5904,N_5961);
and U6066 (N_6066,N_5945,N_5973);
xnor U6067 (N_6067,N_5935,N_5945);
nand U6068 (N_6068,N_5946,N_5984);
nand U6069 (N_6069,N_5987,N_5957);
nor U6070 (N_6070,N_5989,N_5923);
nor U6071 (N_6071,N_5986,N_5939);
and U6072 (N_6072,N_5993,N_5924);
nor U6073 (N_6073,N_5953,N_5946);
and U6074 (N_6074,N_5915,N_5907);
and U6075 (N_6075,N_5969,N_5932);
nand U6076 (N_6076,N_5907,N_5988);
nand U6077 (N_6077,N_5931,N_5998);
nand U6078 (N_6078,N_5979,N_5931);
xor U6079 (N_6079,N_5979,N_5943);
and U6080 (N_6080,N_5903,N_5955);
nand U6081 (N_6081,N_5912,N_5921);
or U6082 (N_6082,N_5961,N_5938);
and U6083 (N_6083,N_5992,N_5929);
nand U6084 (N_6084,N_5909,N_5927);
nand U6085 (N_6085,N_5986,N_5924);
or U6086 (N_6086,N_5975,N_5924);
and U6087 (N_6087,N_5975,N_5943);
and U6088 (N_6088,N_5949,N_5911);
nand U6089 (N_6089,N_5996,N_5980);
nor U6090 (N_6090,N_5995,N_5963);
or U6091 (N_6091,N_5996,N_5921);
and U6092 (N_6092,N_5937,N_5926);
or U6093 (N_6093,N_5900,N_5906);
nor U6094 (N_6094,N_5907,N_5917);
nand U6095 (N_6095,N_5915,N_5900);
xnor U6096 (N_6096,N_5922,N_5967);
nand U6097 (N_6097,N_5947,N_5911);
and U6098 (N_6098,N_5984,N_5922);
nor U6099 (N_6099,N_5914,N_5954);
or U6100 (N_6100,N_6028,N_6064);
or U6101 (N_6101,N_6043,N_6025);
nand U6102 (N_6102,N_6088,N_6058);
nor U6103 (N_6103,N_6010,N_6065);
nor U6104 (N_6104,N_6067,N_6008);
nand U6105 (N_6105,N_6002,N_6042);
xor U6106 (N_6106,N_6012,N_6082);
or U6107 (N_6107,N_6059,N_6031);
or U6108 (N_6108,N_6081,N_6039);
or U6109 (N_6109,N_6015,N_6027);
nor U6110 (N_6110,N_6011,N_6083);
nand U6111 (N_6111,N_6084,N_6001);
or U6112 (N_6112,N_6038,N_6078);
nand U6113 (N_6113,N_6089,N_6087);
nor U6114 (N_6114,N_6071,N_6006);
or U6115 (N_6115,N_6099,N_6068);
nor U6116 (N_6116,N_6020,N_6005);
or U6117 (N_6117,N_6062,N_6090);
or U6118 (N_6118,N_6056,N_6014);
xor U6119 (N_6119,N_6053,N_6029);
or U6120 (N_6120,N_6032,N_6009);
or U6121 (N_6121,N_6092,N_6075);
or U6122 (N_6122,N_6045,N_6050);
and U6123 (N_6123,N_6023,N_6085);
nand U6124 (N_6124,N_6049,N_6036);
nand U6125 (N_6125,N_6026,N_6057);
nor U6126 (N_6126,N_6072,N_6003);
or U6127 (N_6127,N_6018,N_6073);
and U6128 (N_6128,N_6048,N_6022);
nand U6129 (N_6129,N_6034,N_6074);
nor U6130 (N_6130,N_6055,N_6052);
or U6131 (N_6131,N_6004,N_6066);
and U6132 (N_6132,N_6047,N_6037);
nor U6133 (N_6133,N_6021,N_6061);
nand U6134 (N_6134,N_6096,N_6063);
nand U6135 (N_6135,N_6093,N_6007);
nand U6136 (N_6136,N_6044,N_6041);
nand U6137 (N_6137,N_6097,N_6080);
xor U6138 (N_6138,N_6095,N_6017);
nor U6139 (N_6139,N_6040,N_6013);
nor U6140 (N_6140,N_6060,N_6046);
and U6141 (N_6141,N_6024,N_6051);
xor U6142 (N_6142,N_6077,N_6070);
and U6143 (N_6143,N_6019,N_6035);
or U6144 (N_6144,N_6030,N_6091);
nand U6145 (N_6145,N_6016,N_6033);
nand U6146 (N_6146,N_6094,N_6098);
nand U6147 (N_6147,N_6076,N_6069);
nor U6148 (N_6148,N_6000,N_6079);
or U6149 (N_6149,N_6054,N_6086);
and U6150 (N_6150,N_6033,N_6037);
nand U6151 (N_6151,N_6005,N_6076);
nor U6152 (N_6152,N_6078,N_6066);
and U6153 (N_6153,N_6048,N_6065);
and U6154 (N_6154,N_6091,N_6050);
xnor U6155 (N_6155,N_6095,N_6097);
nand U6156 (N_6156,N_6020,N_6025);
nand U6157 (N_6157,N_6099,N_6039);
and U6158 (N_6158,N_6021,N_6050);
xnor U6159 (N_6159,N_6027,N_6046);
and U6160 (N_6160,N_6091,N_6081);
nor U6161 (N_6161,N_6065,N_6069);
nand U6162 (N_6162,N_6041,N_6097);
nand U6163 (N_6163,N_6026,N_6022);
nand U6164 (N_6164,N_6033,N_6012);
or U6165 (N_6165,N_6066,N_6014);
or U6166 (N_6166,N_6030,N_6024);
nor U6167 (N_6167,N_6063,N_6043);
and U6168 (N_6168,N_6006,N_6064);
or U6169 (N_6169,N_6006,N_6079);
nand U6170 (N_6170,N_6045,N_6031);
and U6171 (N_6171,N_6030,N_6072);
nand U6172 (N_6172,N_6055,N_6003);
or U6173 (N_6173,N_6072,N_6069);
nand U6174 (N_6174,N_6006,N_6000);
nand U6175 (N_6175,N_6073,N_6001);
nand U6176 (N_6176,N_6053,N_6059);
nor U6177 (N_6177,N_6042,N_6036);
or U6178 (N_6178,N_6071,N_6088);
nand U6179 (N_6179,N_6000,N_6090);
and U6180 (N_6180,N_6003,N_6043);
nand U6181 (N_6181,N_6041,N_6071);
nand U6182 (N_6182,N_6059,N_6027);
or U6183 (N_6183,N_6052,N_6000);
and U6184 (N_6184,N_6076,N_6039);
xnor U6185 (N_6185,N_6041,N_6033);
xor U6186 (N_6186,N_6045,N_6067);
and U6187 (N_6187,N_6091,N_6057);
nand U6188 (N_6188,N_6049,N_6074);
nor U6189 (N_6189,N_6066,N_6044);
nor U6190 (N_6190,N_6042,N_6063);
and U6191 (N_6191,N_6068,N_6065);
nor U6192 (N_6192,N_6086,N_6097);
and U6193 (N_6193,N_6066,N_6013);
or U6194 (N_6194,N_6043,N_6011);
and U6195 (N_6195,N_6002,N_6045);
or U6196 (N_6196,N_6024,N_6066);
and U6197 (N_6197,N_6035,N_6099);
nand U6198 (N_6198,N_6044,N_6093);
and U6199 (N_6199,N_6029,N_6071);
nand U6200 (N_6200,N_6181,N_6183);
xor U6201 (N_6201,N_6115,N_6199);
xnor U6202 (N_6202,N_6188,N_6100);
nand U6203 (N_6203,N_6174,N_6103);
nor U6204 (N_6204,N_6120,N_6109);
nor U6205 (N_6205,N_6104,N_6141);
nand U6206 (N_6206,N_6142,N_6134);
and U6207 (N_6207,N_6127,N_6119);
and U6208 (N_6208,N_6157,N_6117);
or U6209 (N_6209,N_6111,N_6168);
xor U6210 (N_6210,N_6153,N_6133);
nor U6211 (N_6211,N_6189,N_6148);
or U6212 (N_6212,N_6143,N_6110);
xor U6213 (N_6213,N_6114,N_6122);
nor U6214 (N_6214,N_6164,N_6149);
nor U6215 (N_6215,N_6190,N_6193);
xor U6216 (N_6216,N_6178,N_6140);
nand U6217 (N_6217,N_6118,N_6136);
and U6218 (N_6218,N_6124,N_6137);
nand U6219 (N_6219,N_6112,N_6172);
and U6220 (N_6220,N_6177,N_6123);
and U6221 (N_6221,N_6171,N_6196);
nand U6222 (N_6222,N_6107,N_6102);
or U6223 (N_6223,N_6160,N_6158);
nor U6224 (N_6224,N_6176,N_6185);
nand U6225 (N_6225,N_6152,N_6182);
nand U6226 (N_6226,N_6132,N_6167);
xor U6227 (N_6227,N_6162,N_6165);
and U6228 (N_6228,N_6139,N_6159);
nand U6229 (N_6229,N_6186,N_6192);
and U6230 (N_6230,N_6146,N_6126);
nand U6231 (N_6231,N_6147,N_6179);
nand U6232 (N_6232,N_6194,N_6128);
or U6233 (N_6233,N_6161,N_6187);
nand U6234 (N_6234,N_6135,N_6195);
and U6235 (N_6235,N_6163,N_6191);
nand U6236 (N_6236,N_6145,N_6138);
or U6237 (N_6237,N_6129,N_6197);
or U6238 (N_6238,N_6169,N_6125);
or U6239 (N_6239,N_6198,N_6121);
or U6240 (N_6240,N_6180,N_6155);
xnor U6241 (N_6241,N_6170,N_6130);
nor U6242 (N_6242,N_6106,N_6166);
or U6243 (N_6243,N_6184,N_6151);
or U6244 (N_6244,N_6108,N_6101);
nand U6245 (N_6245,N_6156,N_6175);
or U6246 (N_6246,N_6116,N_6144);
nand U6247 (N_6247,N_6154,N_6150);
or U6248 (N_6248,N_6113,N_6105);
and U6249 (N_6249,N_6173,N_6131);
or U6250 (N_6250,N_6106,N_6104);
nand U6251 (N_6251,N_6177,N_6166);
and U6252 (N_6252,N_6124,N_6189);
nor U6253 (N_6253,N_6179,N_6148);
nand U6254 (N_6254,N_6104,N_6188);
nor U6255 (N_6255,N_6137,N_6126);
nand U6256 (N_6256,N_6127,N_6174);
xnor U6257 (N_6257,N_6193,N_6189);
and U6258 (N_6258,N_6164,N_6176);
nand U6259 (N_6259,N_6157,N_6185);
or U6260 (N_6260,N_6180,N_6169);
xor U6261 (N_6261,N_6127,N_6192);
or U6262 (N_6262,N_6113,N_6185);
or U6263 (N_6263,N_6126,N_6125);
and U6264 (N_6264,N_6121,N_6166);
xor U6265 (N_6265,N_6196,N_6181);
nand U6266 (N_6266,N_6174,N_6169);
nand U6267 (N_6267,N_6180,N_6197);
nor U6268 (N_6268,N_6193,N_6111);
nand U6269 (N_6269,N_6168,N_6112);
or U6270 (N_6270,N_6121,N_6119);
nor U6271 (N_6271,N_6186,N_6145);
and U6272 (N_6272,N_6170,N_6178);
or U6273 (N_6273,N_6169,N_6105);
and U6274 (N_6274,N_6186,N_6135);
or U6275 (N_6275,N_6146,N_6131);
nor U6276 (N_6276,N_6192,N_6136);
nand U6277 (N_6277,N_6138,N_6175);
xor U6278 (N_6278,N_6120,N_6102);
and U6279 (N_6279,N_6123,N_6147);
nand U6280 (N_6280,N_6187,N_6115);
xnor U6281 (N_6281,N_6186,N_6154);
or U6282 (N_6282,N_6176,N_6194);
nor U6283 (N_6283,N_6163,N_6199);
or U6284 (N_6284,N_6189,N_6107);
nor U6285 (N_6285,N_6138,N_6188);
and U6286 (N_6286,N_6196,N_6123);
nor U6287 (N_6287,N_6118,N_6166);
nand U6288 (N_6288,N_6150,N_6166);
and U6289 (N_6289,N_6170,N_6187);
nand U6290 (N_6290,N_6144,N_6101);
nor U6291 (N_6291,N_6125,N_6159);
xnor U6292 (N_6292,N_6150,N_6181);
nor U6293 (N_6293,N_6166,N_6186);
and U6294 (N_6294,N_6179,N_6178);
or U6295 (N_6295,N_6195,N_6134);
xor U6296 (N_6296,N_6139,N_6112);
xnor U6297 (N_6297,N_6100,N_6182);
nand U6298 (N_6298,N_6179,N_6171);
nand U6299 (N_6299,N_6122,N_6168);
nor U6300 (N_6300,N_6267,N_6215);
and U6301 (N_6301,N_6296,N_6221);
or U6302 (N_6302,N_6273,N_6277);
or U6303 (N_6303,N_6269,N_6278);
nand U6304 (N_6304,N_6294,N_6263);
nand U6305 (N_6305,N_6257,N_6229);
or U6306 (N_6306,N_6259,N_6291);
and U6307 (N_6307,N_6247,N_6239);
or U6308 (N_6308,N_6283,N_6209);
or U6309 (N_6309,N_6226,N_6266);
or U6310 (N_6310,N_6210,N_6293);
and U6311 (N_6311,N_6299,N_6252);
nand U6312 (N_6312,N_6279,N_6281);
and U6313 (N_6313,N_6204,N_6289);
xnor U6314 (N_6314,N_6206,N_6200);
nand U6315 (N_6315,N_6213,N_6225);
nor U6316 (N_6316,N_6249,N_6250);
xnor U6317 (N_6317,N_6260,N_6203);
nand U6318 (N_6318,N_6287,N_6231);
xnor U6319 (N_6319,N_6224,N_6286);
nand U6320 (N_6320,N_6248,N_6272);
and U6321 (N_6321,N_6265,N_6245);
or U6322 (N_6322,N_6297,N_6292);
and U6323 (N_6323,N_6246,N_6230);
nand U6324 (N_6324,N_6243,N_6241);
xor U6325 (N_6325,N_6220,N_6275);
and U6326 (N_6326,N_6216,N_6211);
and U6327 (N_6327,N_6240,N_6271);
or U6328 (N_6328,N_6280,N_6258);
or U6329 (N_6329,N_6201,N_6232);
nand U6330 (N_6330,N_6282,N_6274);
and U6331 (N_6331,N_6264,N_6270);
nand U6332 (N_6332,N_6285,N_6254);
nor U6333 (N_6333,N_6234,N_6290);
nor U6334 (N_6334,N_6244,N_6227);
or U6335 (N_6335,N_6202,N_6298);
or U6336 (N_6336,N_6217,N_6235);
and U6337 (N_6337,N_6251,N_6253);
nand U6338 (N_6338,N_6205,N_6268);
nor U6339 (N_6339,N_6214,N_6222);
nor U6340 (N_6340,N_6223,N_6284);
or U6341 (N_6341,N_6236,N_6255);
or U6342 (N_6342,N_6288,N_6238);
and U6343 (N_6343,N_6242,N_6219);
and U6344 (N_6344,N_6207,N_6218);
nand U6345 (N_6345,N_6261,N_6276);
nor U6346 (N_6346,N_6228,N_6256);
or U6347 (N_6347,N_6295,N_6233);
nand U6348 (N_6348,N_6208,N_6262);
nand U6349 (N_6349,N_6237,N_6212);
nand U6350 (N_6350,N_6205,N_6201);
or U6351 (N_6351,N_6206,N_6229);
nor U6352 (N_6352,N_6287,N_6243);
or U6353 (N_6353,N_6201,N_6256);
or U6354 (N_6354,N_6285,N_6262);
nor U6355 (N_6355,N_6244,N_6242);
and U6356 (N_6356,N_6200,N_6235);
and U6357 (N_6357,N_6239,N_6229);
or U6358 (N_6358,N_6290,N_6218);
nor U6359 (N_6359,N_6218,N_6214);
or U6360 (N_6360,N_6289,N_6290);
nor U6361 (N_6361,N_6238,N_6216);
nor U6362 (N_6362,N_6284,N_6274);
and U6363 (N_6363,N_6220,N_6273);
xnor U6364 (N_6364,N_6295,N_6218);
and U6365 (N_6365,N_6250,N_6242);
or U6366 (N_6366,N_6203,N_6270);
and U6367 (N_6367,N_6234,N_6298);
nor U6368 (N_6368,N_6204,N_6213);
nor U6369 (N_6369,N_6230,N_6292);
and U6370 (N_6370,N_6297,N_6222);
nand U6371 (N_6371,N_6265,N_6286);
and U6372 (N_6372,N_6261,N_6263);
nor U6373 (N_6373,N_6229,N_6283);
and U6374 (N_6374,N_6260,N_6219);
or U6375 (N_6375,N_6297,N_6256);
or U6376 (N_6376,N_6273,N_6242);
nor U6377 (N_6377,N_6272,N_6249);
and U6378 (N_6378,N_6292,N_6204);
nor U6379 (N_6379,N_6233,N_6217);
nand U6380 (N_6380,N_6265,N_6294);
and U6381 (N_6381,N_6232,N_6258);
and U6382 (N_6382,N_6295,N_6236);
or U6383 (N_6383,N_6276,N_6216);
nand U6384 (N_6384,N_6209,N_6257);
nor U6385 (N_6385,N_6286,N_6255);
nor U6386 (N_6386,N_6232,N_6221);
or U6387 (N_6387,N_6284,N_6277);
or U6388 (N_6388,N_6286,N_6271);
nor U6389 (N_6389,N_6293,N_6209);
and U6390 (N_6390,N_6247,N_6212);
nor U6391 (N_6391,N_6207,N_6238);
nor U6392 (N_6392,N_6248,N_6285);
nand U6393 (N_6393,N_6226,N_6202);
and U6394 (N_6394,N_6298,N_6223);
xor U6395 (N_6395,N_6285,N_6294);
or U6396 (N_6396,N_6265,N_6212);
xnor U6397 (N_6397,N_6263,N_6254);
xor U6398 (N_6398,N_6270,N_6215);
nand U6399 (N_6399,N_6257,N_6272);
nor U6400 (N_6400,N_6334,N_6356);
or U6401 (N_6401,N_6377,N_6354);
nor U6402 (N_6402,N_6389,N_6391);
nand U6403 (N_6403,N_6379,N_6396);
or U6404 (N_6404,N_6370,N_6358);
xnor U6405 (N_6405,N_6372,N_6364);
nand U6406 (N_6406,N_6371,N_6309);
xnor U6407 (N_6407,N_6340,N_6344);
or U6408 (N_6408,N_6302,N_6329);
and U6409 (N_6409,N_6382,N_6307);
or U6410 (N_6410,N_6349,N_6357);
xor U6411 (N_6411,N_6332,N_6326);
or U6412 (N_6412,N_6331,N_6342);
and U6413 (N_6413,N_6322,N_6373);
nor U6414 (N_6414,N_6386,N_6355);
xor U6415 (N_6415,N_6353,N_6368);
or U6416 (N_6416,N_6392,N_6327);
and U6417 (N_6417,N_6375,N_6335);
xor U6418 (N_6418,N_6378,N_6347);
nor U6419 (N_6419,N_6336,N_6328);
nand U6420 (N_6420,N_6395,N_6385);
or U6421 (N_6421,N_6330,N_6394);
nor U6422 (N_6422,N_6305,N_6321);
nor U6423 (N_6423,N_6313,N_6315);
nor U6424 (N_6424,N_6306,N_6325);
nand U6425 (N_6425,N_6333,N_6388);
and U6426 (N_6426,N_6352,N_6343);
nand U6427 (N_6427,N_6320,N_6324);
nor U6428 (N_6428,N_6317,N_6381);
or U6429 (N_6429,N_6308,N_6338);
nand U6430 (N_6430,N_6397,N_6316);
nand U6431 (N_6431,N_6318,N_6360);
and U6432 (N_6432,N_6399,N_6339);
nand U6433 (N_6433,N_6384,N_6311);
nand U6434 (N_6434,N_6390,N_6348);
or U6435 (N_6435,N_6383,N_6363);
or U6436 (N_6436,N_6314,N_6369);
nor U6437 (N_6437,N_6351,N_6345);
or U6438 (N_6438,N_6310,N_6301);
xnor U6439 (N_6439,N_6319,N_6393);
and U6440 (N_6440,N_6361,N_6374);
xnor U6441 (N_6441,N_6398,N_6323);
and U6442 (N_6442,N_6359,N_6346);
nand U6443 (N_6443,N_6376,N_6362);
or U6444 (N_6444,N_6341,N_6304);
nor U6445 (N_6445,N_6303,N_6300);
or U6446 (N_6446,N_6337,N_6365);
or U6447 (N_6447,N_6387,N_6380);
or U6448 (N_6448,N_6312,N_6367);
nor U6449 (N_6449,N_6366,N_6350);
xor U6450 (N_6450,N_6375,N_6361);
nor U6451 (N_6451,N_6345,N_6316);
and U6452 (N_6452,N_6391,N_6393);
or U6453 (N_6453,N_6302,N_6337);
nor U6454 (N_6454,N_6371,N_6335);
or U6455 (N_6455,N_6334,N_6309);
nand U6456 (N_6456,N_6301,N_6393);
or U6457 (N_6457,N_6380,N_6359);
nor U6458 (N_6458,N_6316,N_6349);
nor U6459 (N_6459,N_6323,N_6316);
nor U6460 (N_6460,N_6345,N_6306);
xnor U6461 (N_6461,N_6347,N_6377);
and U6462 (N_6462,N_6389,N_6360);
nor U6463 (N_6463,N_6339,N_6393);
and U6464 (N_6464,N_6354,N_6328);
and U6465 (N_6465,N_6313,N_6396);
or U6466 (N_6466,N_6351,N_6309);
and U6467 (N_6467,N_6363,N_6300);
nand U6468 (N_6468,N_6346,N_6302);
nand U6469 (N_6469,N_6340,N_6352);
nand U6470 (N_6470,N_6379,N_6371);
nand U6471 (N_6471,N_6381,N_6306);
and U6472 (N_6472,N_6388,N_6369);
or U6473 (N_6473,N_6357,N_6399);
xor U6474 (N_6474,N_6344,N_6356);
and U6475 (N_6475,N_6398,N_6349);
nand U6476 (N_6476,N_6368,N_6392);
or U6477 (N_6477,N_6364,N_6310);
nand U6478 (N_6478,N_6323,N_6339);
or U6479 (N_6479,N_6387,N_6381);
nor U6480 (N_6480,N_6366,N_6301);
or U6481 (N_6481,N_6326,N_6308);
and U6482 (N_6482,N_6337,N_6346);
nand U6483 (N_6483,N_6303,N_6348);
and U6484 (N_6484,N_6362,N_6397);
nand U6485 (N_6485,N_6366,N_6384);
and U6486 (N_6486,N_6351,N_6352);
or U6487 (N_6487,N_6319,N_6359);
and U6488 (N_6488,N_6332,N_6301);
xnor U6489 (N_6489,N_6348,N_6353);
xnor U6490 (N_6490,N_6345,N_6367);
nand U6491 (N_6491,N_6374,N_6313);
nand U6492 (N_6492,N_6374,N_6335);
and U6493 (N_6493,N_6347,N_6313);
nand U6494 (N_6494,N_6369,N_6337);
xnor U6495 (N_6495,N_6379,N_6344);
nand U6496 (N_6496,N_6368,N_6345);
or U6497 (N_6497,N_6354,N_6342);
nor U6498 (N_6498,N_6373,N_6305);
xnor U6499 (N_6499,N_6367,N_6361);
nand U6500 (N_6500,N_6448,N_6441);
and U6501 (N_6501,N_6488,N_6457);
nand U6502 (N_6502,N_6463,N_6421);
nand U6503 (N_6503,N_6458,N_6445);
and U6504 (N_6504,N_6444,N_6454);
nand U6505 (N_6505,N_6479,N_6450);
or U6506 (N_6506,N_6486,N_6483);
xor U6507 (N_6507,N_6415,N_6434);
or U6508 (N_6508,N_6404,N_6420);
nor U6509 (N_6509,N_6411,N_6409);
nor U6510 (N_6510,N_6433,N_6427);
nor U6511 (N_6511,N_6431,N_6453);
nor U6512 (N_6512,N_6456,N_6447);
xnor U6513 (N_6513,N_6497,N_6451);
nand U6514 (N_6514,N_6405,N_6464);
nand U6515 (N_6515,N_6452,N_6435);
nor U6516 (N_6516,N_6495,N_6496);
nor U6517 (N_6517,N_6416,N_6425);
nor U6518 (N_6518,N_6417,N_6439);
or U6519 (N_6519,N_6436,N_6482);
nor U6520 (N_6520,N_6466,N_6429);
or U6521 (N_6521,N_6493,N_6459);
or U6522 (N_6522,N_6424,N_6480);
nor U6523 (N_6523,N_6402,N_6449);
nor U6524 (N_6524,N_6494,N_6406);
and U6525 (N_6525,N_6422,N_6462);
or U6526 (N_6526,N_6442,N_6407);
xor U6527 (N_6527,N_6498,N_6461);
nor U6528 (N_6528,N_6410,N_6426);
or U6529 (N_6529,N_6440,N_6477);
and U6530 (N_6530,N_6473,N_6485);
or U6531 (N_6531,N_6472,N_6484);
and U6532 (N_6532,N_6487,N_6470);
nor U6533 (N_6533,N_6490,N_6475);
nand U6534 (N_6534,N_6481,N_6491);
or U6535 (N_6535,N_6428,N_6437);
nor U6536 (N_6536,N_6413,N_6432);
and U6537 (N_6537,N_6460,N_6455);
and U6538 (N_6538,N_6492,N_6474);
nor U6539 (N_6539,N_6469,N_6468);
nor U6540 (N_6540,N_6478,N_6489);
and U6541 (N_6541,N_6408,N_6446);
nor U6542 (N_6542,N_6423,N_6438);
xor U6543 (N_6543,N_6430,N_6476);
or U6544 (N_6544,N_6419,N_6465);
nand U6545 (N_6545,N_6418,N_6401);
and U6546 (N_6546,N_6499,N_6467);
and U6547 (N_6547,N_6412,N_6471);
and U6548 (N_6548,N_6414,N_6443);
nor U6549 (N_6549,N_6403,N_6400);
nand U6550 (N_6550,N_6423,N_6446);
and U6551 (N_6551,N_6438,N_6416);
and U6552 (N_6552,N_6499,N_6428);
nand U6553 (N_6553,N_6450,N_6486);
xor U6554 (N_6554,N_6408,N_6489);
nand U6555 (N_6555,N_6409,N_6487);
nand U6556 (N_6556,N_6448,N_6492);
or U6557 (N_6557,N_6468,N_6445);
and U6558 (N_6558,N_6432,N_6446);
and U6559 (N_6559,N_6485,N_6451);
nand U6560 (N_6560,N_6488,N_6489);
nand U6561 (N_6561,N_6483,N_6460);
or U6562 (N_6562,N_6431,N_6428);
or U6563 (N_6563,N_6465,N_6442);
nor U6564 (N_6564,N_6407,N_6463);
and U6565 (N_6565,N_6413,N_6457);
and U6566 (N_6566,N_6474,N_6403);
nand U6567 (N_6567,N_6413,N_6422);
and U6568 (N_6568,N_6407,N_6476);
nor U6569 (N_6569,N_6461,N_6404);
or U6570 (N_6570,N_6466,N_6494);
nand U6571 (N_6571,N_6496,N_6481);
nor U6572 (N_6572,N_6408,N_6481);
nand U6573 (N_6573,N_6417,N_6406);
nand U6574 (N_6574,N_6460,N_6453);
or U6575 (N_6575,N_6407,N_6466);
and U6576 (N_6576,N_6414,N_6473);
nand U6577 (N_6577,N_6455,N_6490);
or U6578 (N_6578,N_6444,N_6404);
or U6579 (N_6579,N_6441,N_6412);
nand U6580 (N_6580,N_6426,N_6420);
or U6581 (N_6581,N_6473,N_6420);
and U6582 (N_6582,N_6459,N_6418);
and U6583 (N_6583,N_6402,N_6465);
and U6584 (N_6584,N_6422,N_6428);
nor U6585 (N_6585,N_6488,N_6494);
or U6586 (N_6586,N_6464,N_6450);
and U6587 (N_6587,N_6478,N_6456);
and U6588 (N_6588,N_6442,N_6497);
nand U6589 (N_6589,N_6425,N_6412);
nand U6590 (N_6590,N_6440,N_6429);
nand U6591 (N_6591,N_6485,N_6404);
nand U6592 (N_6592,N_6407,N_6410);
nand U6593 (N_6593,N_6412,N_6491);
nand U6594 (N_6594,N_6467,N_6419);
or U6595 (N_6595,N_6460,N_6405);
or U6596 (N_6596,N_6421,N_6454);
nor U6597 (N_6597,N_6493,N_6466);
or U6598 (N_6598,N_6477,N_6454);
nor U6599 (N_6599,N_6488,N_6493);
nand U6600 (N_6600,N_6515,N_6503);
xnor U6601 (N_6601,N_6550,N_6552);
and U6602 (N_6602,N_6583,N_6561);
nor U6603 (N_6603,N_6522,N_6540);
nand U6604 (N_6604,N_6524,N_6571);
or U6605 (N_6605,N_6534,N_6501);
xnor U6606 (N_6606,N_6508,N_6548);
and U6607 (N_6607,N_6512,N_6595);
and U6608 (N_6608,N_6566,N_6505);
or U6609 (N_6609,N_6560,N_6536);
nor U6610 (N_6610,N_6516,N_6581);
or U6611 (N_6611,N_6530,N_6535);
nand U6612 (N_6612,N_6596,N_6549);
or U6613 (N_6613,N_6500,N_6528);
or U6614 (N_6614,N_6504,N_6576);
nor U6615 (N_6615,N_6562,N_6599);
nand U6616 (N_6616,N_6597,N_6554);
nor U6617 (N_6617,N_6509,N_6506);
and U6618 (N_6618,N_6578,N_6539);
or U6619 (N_6619,N_6513,N_6538);
and U6620 (N_6620,N_6568,N_6587);
and U6621 (N_6621,N_6502,N_6558);
nand U6622 (N_6622,N_6559,N_6545);
xnor U6623 (N_6623,N_6525,N_6572);
nor U6624 (N_6624,N_6531,N_6553);
or U6625 (N_6625,N_6589,N_6537);
nand U6626 (N_6626,N_6523,N_6579);
nor U6627 (N_6627,N_6555,N_6591);
or U6628 (N_6628,N_6517,N_6541);
xor U6629 (N_6629,N_6577,N_6570);
and U6630 (N_6630,N_6582,N_6592);
and U6631 (N_6631,N_6526,N_6544);
and U6632 (N_6632,N_6563,N_6547);
nand U6633 (N_6633,N_6546,N_6569);
nand U6634 (N_6634,N_6567,N_6580);
nor U6635 (N_6635,N_6543,N_6510);
and U6636 (N_6636,N_6575,N_6529);
and U6637 (N_6637,N_6518,N_6527);
and U6638 (N_6638,N_6533,N_6574);
or U6639 (N_6639,N_6590,N_6584);
nand U6640 (N_6640,N_6542,N_6598);
nand U6641 (N_6641,N_6556,N_6588);
nor U6642 (N_6642,N_6593,N_6564);
nand U6643 (N_6643,N_6573,N_6521);
nand U6644 (N_6644,N_6514,N_6520);
nor U6645 (N_6645,N_6557,N_6532);
nand U6646 (N_6646,N_6585,N_6511);
xnor U6647 (N_6647,N_6519,N_6565);
or U6648 (N_6648,N_6551,N_6586);
nand U6649 (N_6649,N_6594,N_6507);
xor U6650 (N_6650,N_6590,N_6568);
or U6651 (N_6651,N_6524,N_6553);
and U6652 (N_6652,N_6541,N_6555);
or U6653 (N_6653,N_6585,N_6574);
or U6654 (N_6654,N_6576,N_6524);
and U6655 (N_6655,N_6501,N_6527);
and U6656 (N_6656,N_6543,N_6540);
and U6657 (N_6657,N_6519,N_6525);
nor U6658 (N_6658,N_6593,N_6540);
and U6659 (N_6659,N_6510,N_6548);
nor U6660 (N_6660,N_6551,N_6589);
or U6661 (N_6661,N_6580,N_6568);
nand U6662 (N_6662,N_6525,N_6506);
or U6663 (N_6663,N_6584,N_6524);
nor U6664 (N_6664,N_6545,N_6516);
and U6665 (N_6665,N_6583,N_6553);
nand U6666 (N_6666,N_6569,N_6529);
nand U6667 (N_6667,N_6585,N_6592);
nor U6668 (N_6668,N_6586,N_6560);
or U6669 (N_6669,N_6566,N_6578);
nand U6670 (N_6670,N_6536,N_6521);
xor U6671 (N_6671,N_6586,N_6532);
or U6672 (N_6672,N_6564,N_6555);
nor U6673 (N_6673,N_6531,N_6543);
nand U6674 (N_6674,N_6534,N_6586);
and U6675 (N_6675,N_6507,N_6533);
nor U6676 (N_6676,N_6560,N_6535);
nand U6677 (N_6677,N_6597,N_6534);
nand U6678 (N_6678,N_6560,N_6585);
xor U6679 (N_6679,N_6571,N_6586);
nand U6680 (N_6680,N_6500,N_6532);
nand U6681 (N_6681,N_6599,N_6534);
and U6682 (N_6682,N_6500,N_6540);
nor U6683 (N_6683,N_6538,N_6572);
nand U6684 (N_6684,N_6578,N_6564);
and U6685 (N_6685,N_6577,N_6579);
and U6686 (N_6686,N_6529,N_6519);
nand U6687 (N_6687,N_6560,N_6540);
and U6688 (N_6688,N_6526,N_6598);
or U6689 (N_6689,N_6552,N_6504);
or U6690 (N_6690,N_6517,N_6581);
xor U6691 (N_6691,N_6543,N_6583);
nand U6692 (N_6692,N_6504,N_6547);
and U6693 (N_6693,N_6507,N_6573);
xnor U6694 (N_6694,N_6581,N_6549);
or U6695 (N_6695,N_6516,N_6583);
or U6696 (N_6696,N_6539,N_6552);
xor U6697 (N_6697,N_6502,N_6549);
and U6698 (N_6698,N_6530,N_6575);
nand U6699 (N_6699,N_6557,N_6535);
or U6700 (N_6700,N_6631,N_6676);
and U6701 (N_6701,N_6616,N_6633);
or U6702 (N_6702,N_6655,N_6638);
and U6703 (N_6703,N_6628,N_6609);
or U6704 (N_6704,N_6639,N_6694);
nand U6705 (N_6705,N_6672,N_6627);
and U6706 (N_6706,N_6660,N_6626);
and U6707 (N_6707,N_6654,N_6662);
nor U6708 (N_6708,N_6643,N_6647);
nor U6709 (N_6709,N_6648,N_6663);
and U6710 (N_6710,N_6683,N_6612);
and U6711 (N_6711,N_6688,N_6611);
nand U6712 (N_6712,N_6677,N_6636);
and U6713 (N_6713,N_6601,N_6691);
and U6714 (N_6714,N_6669,N_6698);
nand U6715 (N_6715,N_6674,N_6614);
nor U6716 (N_6716,N_6652,N_6665);
nor U6717 (N_6717,N_6646,N_6685);
and U6718 (N_6718,N_6666,N_6644);
and U6719 (N_6719,N_6696,N_6608);
and U6720 (N_6720,N_6692,N_6617);
nor U6721 (N_6721,N_6645,N_6630);
and U6722 (N_6722,N_6659,N_6632);
nand U6723 (N_6723,N_6678,N_6687);
or U6724 (N_6724,N_6673,N_6610);
and U6725 (N_6725,N_6668,N_6681);
nor U6726 (N_6726,N_6656,N_6629);
or U6727 (N_6727,N_6620,N_6641);
or U6728 (N_6728,N_6623,N_6670);
nand U6729 (N_6729,N_6602,N_6640);
nand U6730 (N_6730,N_6686,N_6695);
nand U6731 (N_6731,N_6682,N_6605);
or U6732 (N_6732,N_6689,N_6618);
nand U6733 (N_6733,N_6684,N_6690);
nor U6734 (N_6734,N_6615,N_6624);
and U6735 (N_6735,N_6699,N_6671);
nand U6736 (N_6736,N_6622,N_6649);
nand U6737 (N_6737,N_6667,N_6653);
nor U6738 (N_6738,N_6650,N_6651);
or U6739 (N_6739,N_6675,N_6604);
nor U6740 (N_6740,N_6603,N_6634);
and U6741 (N_6741,N_6661,N_6607);
and U6742 (N_6742,N_6606,N_6693);
nand U6743 (N_6743,N_6657,N_6642);
nor U6744 (N_6744,N_6637,N_6635);
and U6745 (N_6745,N_6600,N_6697);
nor U6746 (N_6746,N_6625,N_6658);
nand U6747 (N_6747,N_6664,N_6679);
and U6748 (N_6748,N_6680,N_6621);
nor U6749 (N_6749,N_6613,N_6619);
or U6750 (N_6750,N_6621,N_6652);
nor U6751 (N_6751,N_6686,N_6674);
and U6752 (N_6752,N_6690,N_6608);
nand U6753 (N_6753,N_6699,N_6652);
or U6754 (N_6754,N_6614,N_6637);
or U6755 (N_6755,N_6672,N_6671);
and U6756 (N_6756,N_6680,N_6610);
and U6757 (N_6757,N_6611,N_6604);
or U6758 (N_6758,N_6672,N_6629);
and U6759 (N_6759,N_6620,N_6660);
nand U6760 (N_6760,N_6612,N_6605);
and U6761 (N_6761,N_6639,N_6610);
nand U6762 (N_6762,N_6680,N_6653);
nand U6763 (N_6763,N_6646,N_6641);
and U6764 (N_6764,N_6621,N_6642);
or U6765 (N_6765,N_6686,N_6623);
nand U6766 (N_6766,N_6653,N_6630);
and U6767 (N_6767,N_6612,N_6684);
nor U6768 (N_6768,N_6600,N_6615);
nand U6769 (N_6769,N_6632,N_6640);
nor U6770 (N_6770,N_6602,N_6656);
nand U6771 (N_6771,N_6697,N_6648);
nor U6772 (N_6772,N_6657,N_6692);
xnor U6773 (N_6773,N_6652,N_6630);
and U6774 (N_6774,N_6693,N_6639);
or U6775 (N_6775,N_6655,N_6653);
nand U6776 (N_6776,N_6608,N_6625);
nor U6777 (N_6777,N_6612,N_6631);
and U6778 (N_6778,N_6685,N_6624);
nor U6779 (N_6779,N_6698,N_6672);
nor U6780 (N_6780,N_6600,N_6640);
nand U6781 (N_6781,N_6606,N_6616);
nand U6782 (N_6782,N_6648,N_6656);
nor U6783 (N_6783,N_6644,N_6634);
and U6784 (N_6784,N_6632,N_6626);
and U6785 (N_6785,N_6654,N_6667);
or U6786 (N_6786,N_6602,N_6675);
and U6787 (N_6787,N_6661,N_6657);
nand U6788 (N_6788,N_6616,N_6628);
nand U6789 (N_6789,N_6668,N_6657);
nor U6790 (N_6790,N_6677,N_6604);
or U6791 (N_6791,N_6683,N_6655);
and U6792 (N_6792,N_6655,N_6692);
or U6793 (N_6793,N_6635,N_6655);
nor U6794 (N_6794,N_6639,N_6631);
nor U6795 (N_6795,N_6691,N_6677);
nand U6796 (N_6796,N_6621,N_6622);
nor U6797 (N_6797,N_6648,N_6653);
and U6798 (N_6798,N_6655,N_6619);
and U6799 (N_6799,N_6610,N_6617);
nand U6800 (N_6800,N_6795,N_6789);
nand U6801 (N_6801,N_6785,N_6702);
or U6802 (N_6802,N_6779,N_6723);
or U6803 (N_6803,N_6759,N_6700);
and U6804 (N_6804,N_6742,N_6713);
nor U6805 (N_6805,N_6765,N_6725);
and U6806 (N_6806,N_6740,N_6791);
nand U6807 (N_6807,N_6735,N_6708);
nor U6808 (N_6808,N_6732,N_6780);
nand U6809 (N_6809,N_6710,N_6790);
nor U6810 (N_6810,N_6752,N_6736);
nand U6811 (N_6811,N_6706,N_6764);
nand U6812 (N_6812,N_6777,N_6738);
and U6813 (N_6813,N_6786,N_6754);
nand U6814 (N_6814,N_6749,N_6734);
and U6815 (N_6815,N_6748,N_6761);
or U6816 (N_6816,N_6712,N_6719);
nand U6817 (N_6817,N_6727,N_6792);
and U6818 (N_6818,N_6720,N_6701);
or U6819 (N_6819,N_6793,N_6770);
or U6820 (N_6820,N_6782,N_6787);
and U6821 (N_6821,N_6709,N_6772);
nor U6822 (N_6822,N_6774,N_6788);
nand U6823 (N_6823,N_6760,N_6784);
and U6824 (N_6824,N_6717,N_6762);
nor U6825 (N_6825,N_6730,N_6796);
nand U6826 (N_6826,N_6704,N_6737);
xor U6827 (N_6827,N_6766,N_6743);
and U6828 (N_6828,N_6745,N_6726);
and U6829 (N_6829,N_6771,N_6707);
nand U6830 (N_6830,N_6799,N_6729);
and U6831 (N_6831,N_6773,N_6715);
or U6832 (N_6832,N_6705,N_6741);
nand U6833 (N_6833,N_6731,N_6721);
nand U6834 (N_6834,N_6714,N_6755);
nand U6835 (N_6835,N_6751,N_6767);
nor U6836 (N_6836,N_6794,N_6718);
nand U6837 (N_6837,N_6724,N_6758);
or U6838 (N_6838,N_6746,N_6739);
nor U6839 (N_6839,N_6722,N_6776);
and U6840 (N_6840,N_6797,N_6716);
xor U6841 (N_6841,N_6728,N_6768);
and U6842 (N_6842,N_6703,N_6757);
nand U6843 (N_6843,N_6763,N_6781);
nand U6844 (N_6844,N_6756,N_6733);
or U6845 (N_6845,N_6744,N_6711);
or U6846 (N_6846,N_6775,N_6750);
or U6847 (N_6847,N_6798,N_6769);
nand U6848 (N_6848,N_6747,N_6753);
nand U6849 (N_6849,N_6783,N_6778);
nor U6850 (N_6850,N_6733,N_6725);
and U6851 (N_6851,N_6734,N_6798);
and U6852 (N_6852,N_6781,N_6766);
and U6853 (N_6853,N_6752,N_6793);
nor U6854 (N_6854,N_6723,N_6785);
nor U6855 (N_6855,N_6778,N_6786);
nor U6856 (N_6856,N_6750,N_6759);
nand U6857 (N_6857,N_6716,N_6768);
nor U6858 (N_6858,N_6742,N_6753);
nor U6859 (N_6859,N_6768,N_6776);
nand U6860 (N_6860,N_6759,N_6761);
or U6861 (N_6861,N_6767,N_6743);
nand U6862 (N_6862,N_6725,N_6741);
and U6863 (N_6863,N_6742,N_6778);
nand U6864 (N_6864,N_6793,N_6723);
or U6865 (N_6865,N_6739,N_6733);
xor U6866 (N_6866,N_6775,N_6711);
nand U6867 (N_6867,N_6731,N_6764);
and U6868 (N_6868,N_6793,N_6703);
xor U6869 (N_6869,N_6773,N_6752);
and U6870 (N_6870,N_6779,N_6719);
or U6871 (N_6871,N_6777,N_6752);
nor U6872 (N_6872,N_6744,N_6787);
nand U6873 (N_6873,N_6726,N_6798);
or U6874 (N_6874,N_6731,N_6717);
nand U6875 (N_6875,N_6701,N_6711);
nor U6876 (N_6876,N_6704,N_6733);
nand U6877 (N_6877,N_6730,N_6744);
or U6878 (N_6878,N_6703,N_6782);
nor U6879 (N_6879,N_6702,N_6796);
nand U6880 (N_6880,N_6754,N_6762);
nor U6881 (N_6881,N_6702,N_6768);
nand U6882 (N_6882,N_6782,N_6741);
and U6883 (N_6883,N_6733,N_6763);
nand U6884 (N_6884,N_6766,N_6773);
or U6885 (N_6885,N_6782,N_6729);
nor U6886 (N_6886,N_6792,N_6748);
nor U6887 (N_6887,N_6771,N_6748);
and U6888 (N_6888,N_6711,N_6760);
and U6889 (N_6889,N_6740,N_6701);
and U6890 (N_6890,N_6728,N_6798);
nor U6891 (N_6891,N_6798,N_6705);
nor U6892 (N_6892,N_6725,N_6793);
nand U6893 (N_6893,N_6777,N_6768);
and U6894 (N_6894,N_6788,N_6737);
xor U6895 (N_6895,N_6793,N_6738);
nand U6896 (N_6896,N_6722,N_6745);
or U6897 (N_6897,N_6776,N_6700);
and U6898 (N_6898,N_6785,N_6775);
and U6899 (N_6899,N_6719,N_6752);
and U6900 (N_6900,N_6847,N_6811);
xnor U6901 (N_6901,N_6857,N_6873);
or U6902 (N_6902,N_6886,N_6868);
or U6903 (N_6903,N_6887,N_6899);
nand U6904 (N_6904,N_6876,N_6879);
or U6905 (N_6905,N_6878,N_6865);
nor U6906 (N_6906,N_6894,N_6875);
xor U6907 (N_6907,N_6898,N_6801);
and U6908 (N_6908,N_6816,N_6800);
or U6909 (N_6909,N_6867,N_6812);
and U6910 (N_6910,N_6822,N_6892);
and U6911 (N_6911,N_6863,N_6828);
nand U6912 (N_6912,N_6820,N_6860);
and U6913 (N_6913,N_6856,N_6835);
nor U6914 (N_6914,N_6819,N_6836);
nand U6915 (N_6915,N_6840,N_6818);
or U6916 (N_6916,N_6869,N_6884);
nand U6917 (N_6917,N_6831,N_6853);
or U6918 (N_6918,N_6842,N_6814);
nor U6919 (N_6919,N_6804,N_6897);
xor U6920 (N_6920,N_6837,N_6885);
and U6921 (N_6921,N_6852,N_6846);
nand U6922 (N_6922,N_6877,N_6824);
and U6923 (N_6923,N_6866,N_6803);
or U6924 (N_6924,N_6854,N_6808);
xor U6925 (N_6925,N_6838,N_6859);
and U6926 (N_6926,N_6815,N_6806);
nor U6927 (N_6927,N_6882,N_6883);
nor U6928 (N_6928,N_6844,N_6832);
or U6929 (N_6929,N_6872,N_6829);
and U6930 (N_6930,N_6809,N_6807);
nor U6931 (N_6931,N_6889,N_6896);
nor U6932 (N_6932,N_6849,N_6864);
nor U6933 (N_6933,N_6862,N_6880);
or U6934 (N_6934,N_6839,N_6891);
or U6935 (N_6935,N_6810,N_6848);
nand U6936 (N_6936,N_6843,N_6817);
nor U6937 (N_6937,N_6870,N_6813);
nand U6938 (N_6938,N_6827,N_6895);
or U6939 (N_6939,N_6851,N_6841);
and U6940 (N_6940,N_6871,N_6802);
and U6941 (N_6941,N_6823,N_6845);
nor U6942 (N_6942,N_6834,N_6881);
nor U6943 (N_6943,N_6893,N_6858);
xor U6944 (N_6944,N_6855,N_6825);
and U6945 (N_6945,N_6890,N_6888);
nor U6946 (N_6946,N_6874,N_6861);
or U6947 (N_6947,N_6821,N_6826);
and U6948 (N_6948,N_6805,N_6830);
xor U6949 (N_6949,N_6850,N_6833);
nor U6950 (N_6950,N_6825,N_6847);
or U6951 (N_6951,N_6883,N_6833);
and U6952 (N_6952,N_6864,N_6834);
nand U6953 (N_6953,N_6855,N_6808);
and U6954 (N_6954,N_6800,N_6868);
or U6955 (N_6955,N_6898,N_6836);
or U6956 (N_6956,N_6835,N_6867);
and U6957 (N_6957,N_6831,N_6895);
xnor U6958 (N_6958,N_6821,N_6804);
nor U6959 (N_6959,N_6856,N_6898);
or U6960 (N_6960,N_6884,N_6859);
and U6961 (N_6961,N_6895,N_6839);
and U6962 (N_6962,N_6831,N_6861);
nand U6963 (N_6963,N_6839,N_6893);
nand U6964 (N_6964,N_6850,N_6887);
nor U6965 (N_6965,N_6835,N_6875);
and U6966 (N_6966,N_6823,N_6884);
or U6967 (N_6967,N_6868,N_6808);
and U6968 (N_6968,N_6812,N_6821);
and U6969 (N_6969,N_6802,N_6881);
nor U6970 (N_6970,N_6804,N_6838);
or U6971 (N_6971,N_6863,N_6827);
nor U6972 (N_6972,N_6881,N_6838);
nand U6973 (N_6973,N_6858,N_6813);
and U6974 (N_6974,N_6812,N_6873);
nor U6975 (N_6975,N_6891,N_6830);
or U6976 (N_6976,N_6838,N_6837);
and U6977 (N_6977,N_6890,N_6851);
nor U6978 (N_6978,N_6832,N_6838);
xor U6979 (N_6979,N_6876,N_6825);
nand U6980 (N_6980,N_6854,N_6852);
and U6981 (N_6981,N_6872,N_6852);
xor U6982 (N_6982,N_6872,N_6806);
and U6983 (N_6983,N_6856,N_6870);
nand U6984 (N_6984,N_6885,N_6877);
nand U6985 (N_6985,N_6856,N_6820);
nor U6986 (N_6986,N_6879,N_6875);
nor U6987 (N_6987,N_6846,N_6842);
nor U6988 (N_6988,N_6875,N_6814);
nor U6989 (N_6989,N_6846,N_6894);
or U6990 (N_6990,N_6870,N_6859);
and U6991 (N_6991,N_6819,N_6858);
nor U6992 (N_6992,N_6832,N_6816);
xor U6993 (N_6993,N_6856,N_6893);
nor U6994 (N_6994,N_6847,N_6868);
and U6995 (N_6995,N_6862,N_6839);
nand U6996 (N_6996,N_6896,N_6872);
nand U6997 (N_6997,N_6850,N_6892);
nand U6998 (N_6998,N_6869,N_6854);
or U6999 (N_6999,N_6857,N_6803);
nand U7000 (N_7000,N_6985,N_6957);
nand U7001 (N_7001,N_6917,N_6982);
nand U7002 (N_7002,N_6915,N_6989);
xnor U7003 (N_7003,N_6963,N_6959);
and U7004 (N_7004,N_6969,N_6958);
nor U7005 (N_7005,N_6981,N_6964);
or U7006 (N_7006,N_6975,N_6935);
and U7007 (N_7007,N_6903,N_6955);
and U7008 (N_7008,N_6939,N_6900);
nor U7009 (N_7009,N_6972,N_6909);
nand U7010 (N_7010,N_6943,N_6991);
nor U7011 (N_7011,N_6911,N_6914);
nor U7012 (N_7012,N_6987,N_6921);
nor U7013 (N_7013,N_6931,N_6908);
and U7014 (N_7014,N_6983,N_6998);
and U7015 (N_7015,N_6924,N_6960);
nand U7016 (N_7016,N_6910,N_6956);
nor U7017 (N_7017,N_6942,N_6974);
or U7018 (N_7018,N_6999,N_6904);
and U7019 (N_7019,N_6961,N_6949);
xnor U7020 (N_7020,N_6926,N_6925);
or U7021 (N_7021,N_6994,N_6944);
nand U7022 (N_7022,N_6940,N_6967);
nor U7023 (N_7023,N_6937,N_6945);
nor U7024 (N_7024,N_6979,N_6912);
nor U7025 (N_7025,N_6934,N_6919);
and U7026 (N_7026,N_6907,N_6901);
nand U7027 (N_7027,N_6986,N_6966);
nor U7028 (N_7028,N_6922,N_6946);
and U7029 (N_7029,N_6950,N_6953);
nor U7030 (N_7030,N_6948,N_6984);
or U7031 (N_7031,N_6970,N_6918);
nor U7032 (N_7032,N_6930,N_6929);
nand U7033 (N_7033,N_6905,N_6990);
xor U7034 (N_7034,N_6962,N_6938);
nor U7035 (N_7035,N_6997,N_6977);
or U7036 (N_7036,N_6902,N_6920);
nand U7037 (N_7037,N_6988,N_6978);
nor U7038 (N_7038,N_6992,N_6951);
or U7039 (N_7039,N_6995,N_6996);
and U7040 (N_7040,N_6976,N_6980);
nor U7041 (N_7041,N_6932,N_6954);
or U7042 (N_7042,N_6933,N_6952);
or U7043 (N_7043,N_6913,N_6936);
or U7044 (N_7044,N_6968,N_6927);
nor U7045 (N_7045,N_6965,N_6973);
nor U7046 (N_7046,N_6941,N_6928);
or U7047 (N_7047,N_6923,N_6993);
nor U7048 (N_7048,N_6971,N_6947);
nor U7049 (N_7049,N_6916,N_6906);
nor U7050 (N_7050,N_6988,N_6906);
or U7051 (N_7051,N_6968,N_6973);
nand U7052 (N_7052,N_6965,N_6999);
or U7053 (N_7053,N_6955,N_6943);
nor U7054 (N_7054,N_6943,N_6930);
or U7055 (N_7055,N_6950,N_6977);
nor U7056 (N_7056,N_6951,N_6949);
and U7057 (N_7057,N_6960,N_6919);
or U7058 (N_7058,N_6913,N_6926);
nor U7059 (N_7059,N_6993,N_6969);
nor U7060 (N_7060,N_6902,N_6903);
nor U7061 (N_7061,N_6947,N_6922);
nand U7062 (N_7062,N_6967,N_6972);
or U7063 (N_7063,N_6903,N_6934);
nand U7064 (N_7064,N_6982,N_6944);
nand U7065 (N_7065,N_6959,N_6922);
nand U7066 (N_7066,N_6924,N_6978);
nand U7067 (N_7067,N_6936,N_6996);
and U7068 (N_7068,N_6918,N_6919);
nor U7069 (N_7069,N_6986,N_6951);
and U7070 (N_7070,N_6970,N_6921);
xor U7071 (N_7071,N_6947,N_6973);
xor U7072 (N_7072,N_6905,N_6985);
nor U7073 (N_7073,N_6923,N_6968);
nand U7074 (N_7074,N_6900,N_6992);
or U7075 (N_7075,N_6955,N_6915);
xnor U7076 (N_7076,N_6996,N_6935);
or U7077 (N_7077,N_6990,N_6932);
nand U7078 (N_7078,N_6926,N_6946);
xnor U7079 (N_7079,N_6930,N_6957);
and U7080 (N_7080,N_6973,N_6934);
or U7081 (N_7081,N_6994,N_6990);
nor U7082 (N_7082,N_6918,N_6939);
nand U7083 (N_7083,N_6996,N_6920);
and U7084 (N_7084,N_6977,N_6999);
xnor U7085 (N_7085,N_6931,N_6904);
or U7086 (N_7086,N_6908,N_6987);
and U7087 (N_7087,N_6909,N_6912);
nor U7088 (N_7088,N_6998,N_6973);
and U7089 (N_7089,N_6908,N_6974);
nor U7090 (N_7090,N_6982,N_6956);
and U7091 (N_7091,N_6919,N_6942);
xnor U7092 (N_7092,N_6915,N_6975);
nand U7093 (N_7093,N_6915,N_6947);
nor U7094 (N_7094,N_6929,N_6995);
or U7095 (N_7095,N_6919,N_6991);
nor U7096 (N_7096,N_6998,N_6971);
or U7097 (N_7097,N_6917,N_6901);
nor U7098 (N_7098,N_6982,N_6936);
or U7099 (N_7099,N_6911,N_6962);
and U7100 (N_7100,N_7095,N_7014);
nor U7101 (N_7101,N_7088,N_7041);
or U7102 (N_7102,N_7044,N_7052);
or U7103 (N_7103,N_7069,N_7032);
nand U7104 (N_7104,N_7079,N_7023);
and U7105 (N_7105,N_7046,N_7073);
or U7106 (N_7106,N_7086,N_7051);
nand U7107 (N_7107,N_7028,N_7059);
and U7108 (N_7108,N_7090,N_7003);
and U7109 (N_7109,N_7020,N_7066);
nor U7110 (N_7110,N_7050,N_7061);
nand U7111 (N_7111,N_7084,N_7037);
and U7112 (N_7112,N_7060,N_7043);
xnor U7113 (N_7113,N_7033,N_7006);
nand U7114 (N_7114,N_7005,N_7057);
or U7115 (N_7115,N_7010,N_7089);
xnor U7116 (N_7116,N_7013,N_7072);
nor U7117 (N_7117,N_7036,N_7012);
xnor U7118 (N_7118,N_7029,N_7025);
xor U7119 (N_7119,N_7064,N_7015);
nand U7120 (N_7120,N_7031,N_7035);
and U7121 (N_7121,N_7001,N_7008);
and U7122 (N_7122,N_7002,N_7007);
or U7123 (N_7123,N_7000,N_7063);
xnor U7124 (N_7124,N_7017,N_7068);
nor U7125 (N_7125,N_7076,N_7009);
or U7126 (N_7126,N_7042,N_7087);
nor U7127 (N_7127,N_7056,N_7016);
or U7128 (N_7128,N_7094,N_7022);
nor U7129 (N_7129,N_7070,N_7099);
nor U7130 (N_7130,N_7034,N_7078);
or U7131 (N_7131,N_7047,N_7049);
or U7132 (N_7132,N_7075,N_7054);
nand U7133 (N_7133,N_7080,N_7018);
nand U7134 (N_7134,N_7045,N_7067);
nor U7135 (N_7135,N_7081,N_7096);
or U7136 (N_7136,N_7004,N_7021);
or U7137 (N_7137,N_7024,N_7055);
xnor U7138 (N_7138,N_7071,N_7077);
nand U7139 (N_7139,N_7062,N_7019);
or U7140 (N_7140,N_7026,N_7065);
nand U7141 (N_7141,N_7091,N_7098);
xnor U7142 (N_7142,N_7038,N_7030);
xor U7143 (N_7143,N_7027,N_7082);
or U7144 (N_7144,N_7040,N_7011);
or U7145 (N_7145,N_7053,N_7083);
or U7146 (N_7146,N_7048,N_7058);
nand U7147 (N_7147,N_7097,N_7039);
nand U7148 (N_7148,N_7093,N_7085);
and U7149 (N_7149,N_7092,N_7074);
nand U7150 (N_7150,N_7021,N_7027);
nor U7151 (N_7151,N_7078,N_7087);
nor U7152 (N_7152,N_7030,N_7007);
or U7153 (N_7153,N_7031,N_7034);
and U7154 (N_7154,N_7059,N_7084);
or U7155 (N_7155,N_7068,N_7006);
or U7156 (N_7156,N_7061,N_7046);
and U7157 (N_7157,N_7035,N_7042);
nor U7158 (N_7158,N_7038,N_7035);
xor U7159 (N_7159,N_7071,N_7006);
and U7160 (N_7160,N_7011,N_7027);
and U7161 (N_7161,N_7086,N_7002);
nor U7162 (N_7162,N_7039,N_7005);
and U7163 (N_7163,N_7028,N_7067);
nor U7164 (N_7164,N_7065,N_7016);
nand U7165 (N_7165,N_7019,N_7024);
or U7166 (N_7166,N_7066,N_7058);
nor U7167 (N_7167,N_7014,N_7017);
or U7168 (N_7168,N_7085,N_7007);
nor U7169 (N_7169,N_7040,N_7023);
nand U7170 (N_7170,N_7050,N_7001);
or U7171 (N_7171,N_7063,N_7073);
and U7172 (N_7172,N_7099,N_7033);
nor U7173 (N_7173,N_7087,N_7025);
nor U7174 (N_7174,N_7012,N_7002);
nand U7175 (N_7175,N_7004,N_7041);
or U7176 (N_7176,N_7087,N_7050);
xor U7177 (N_7177,N_7088,N_7062);
or U7178 (N_7178,N_7086,N_7029);
nand U7179 (N_7179,N_7064,N_7024);
nor U7180 (N_7180,N_7029,N_7069);
xor U7181 (N_7181,N_7003,N_7046);
nor U7182 (N_7182,N_7052,N_7000);
nor U7183 (N_7183,N_7026,N_7084);
nand U7184 (N_7184,N_7041,N_7006);
or U7185 (N_7185,N_7019,N_7079);
and U7186 (N_7186,N_7023,N_7067);
or U7187 (N_7187,N_7033,N_7044);
nand U7188 (N_7188,N_7043,N_7031);
or U7189 (N_7189,N_7027,N_7064);
or U7190 (N_7190,N_7011,N_7088);
nand U7191 (N_7191,N_7018,N_7088);
or U7192 (N_7192,N_7075,N_7097);
xor U7193 (N_7193,N_7017,N_7029);
nor U7194 (N_7194,N_7077,N_7027);
nor U7195 (N_7195,N_7070,N_7008);
and U7196 (N_7196,N_7027,N_7083);
and U7197 (N_7197,N_7088,N_7060);
and U7198 (N_7198,N_7098,N_7076);
nor U7199 (N_7199,N_7004,N_7025);
nand U7200 (N_7200,N_7196,N_7120);
and U7201 (N_7201,N_7189,N_7147);
or U7202 (N_7202,N_7158,N_7171);
or U7203 (N_7203,N_7168,N_7125);
xnor U7204 (N_7204,N_7128,N_7179);
xor U7205 (N_7205,N_7155,N_7102);
nor U7206 (N_7206,N_7118,N_7129);
nand U7207 (N_7207,N_7113,N_7138);
and U7208 (N_7208,N_7153,N_7123);
and U7209 (N_7209,N_7174,N_7104);
and U7210 (N_7210,N_7109,N_7176);
xnor U7211 (N_7211,N_7115,N_7173);
nand U7212 (N_7212,N_7130,N_7170);
or U7213 (N_7213,N_7101,N_7165);
or U7214 (N_7214,N_7142,N_7137);
or U7215 (N_7215,N_7197,N_7167);
and U7216 (N_7216,N_7181,N_7185);
xnor U7217 (N_7217,N_7166,N_7103);
nor U7218 (N_7218,N_7157,N_7161);
nor U7219 (N_7219,N_7111,N_7164);
nor U7220 (N_7220,N_7154,N_7116);
xor U7221 (N_7221,N_7124,N_7183);
nor U7222 (N_7222,N_7134,N_7190);
nor U7223 (N_7223,N_7106,N_7136);
nor U7224 (N_7224,N_7140,N_7107);
nand U7225 (N_7225,N_7177,N_7192);
nor U7226 (N_7226,N_7121,N_7198);
nor U7227 (N_7227,N_7114,N_7160);
and U7228 (N_7228,N_7139,N_7122);
nor U7229 (N_7229,N_7193,N_7105);
xor U7230 (N_7230,N_7143,N_7163);
nand U7231 (N_7231,N_7133,N_7152);
nand U7232 (N_7232,N_7187,N_7117);
nor U7233 (N_7233,N_7199,N_7188);
nor U7234 (N_7234,N_7150,N_7175);
nor U7235 (N_7235,N_7159,N_7151);
nand U7236 (N_7236,N_7194,N_7186);
nand U7237 (N_7237,N_7144,N_7148);
or U7238 (N_7238,N_7156,N_7135);
and U7239 (N_7239,N_7131,N_7149);
nand U7240 (N_7240,N_7178,N_7162);
and U7241 (N_7241,N_7119,N_7182);
nand U7242 (N_7242,N_7146,N_7108);
or U7243 (N_7243,N_7112,N_7195);
nor U7244 (N_7244,N_7100,N_7127);
xnor U7245 (N_7245,N_7141,N_7169);
and U7246 (N_7246,N_7184,N_7110);
or U7247 (N_7247,N_7132,N_7191);
or U7248 (N_7248,N_7145,N_7180);
xnor U7249 (N_7249,N_7126,N_7172);
nand U7250 (N_7250,N_7179,N_7198);
and U7251 (N_7251,N_7162,N_7187);
or U7252 (N_7252,N_7140,N_7130);
nor U7253 (N_7253,N_7137,N_7162);
and U7254 (N_7254,N_7112,N_7191);
and U7255 (N_7255,N_7199,N_7138);
xor U7256 (N_7256,N_7103,N_7154);
and U7257 (N_7257,N_7147,N_7128);
nand U7258 (N_7258,N_7154,N_7183);
and U7259 (N_7259,N_7171,N_7198);
nor U7260 (N_7260,N_7166,N_7177);
and U7261 (N_7261,N_7146,N_7151);
nor U7262 (N_7262,N_7195,N_7148);
nand U7263 (N_7263,N_7148,N_7177);
or U7264 (N_7264,N_7130,N_7141);
nand U7265 (N_7265,N_7139,N_7149);
nand U7266 (N_7266,N_7141,N_7135);
or U7267 (N_7267,N_7102,N_7189);
nor U7268 (N_7268,N_7148,N_7131);
and U7269 (N_7269,N_7143,N_7135);
nand U7270 (N_7270,N_7189,N_7132);
nor U7271 (N_7271,N_7107,N_7192);
or U7272 (N_7272,N_7145,N_7132);
and U7273 (N_7273,N_7113,N_7143);
nand U7274 (N_7274,N_7126,N_7134);
xnor U7275 (N_7275,N_7140,N_7149);
or U7276 (N_7276,N_7169,N_7170);
nor U7277 (N_7277,N_7184,N_7103);
and U7278 (N_7278,N_7129,N_7131);
nand U7279 (N_7279,N_7119,N_7105);
or U7280 (N_7280,N_7179,N_7129);
or U7281 (N_7281,N_7109,N_7131);
nor U7282 (N_7282,N_7131,N_7181);
and U7283 (N_7283,N_7142,N_7144);
and U7284 (N_7284,N_7192,N_7155);
nor U7285 (N_7285,N_7156,N_7159);
nor U7286 (N_7286,N_7168,N_7175);
nand U7287 (N_7287,N_7111,N_7166);
nor U7288 (N_7288,N_7108,N_7145);
xnor U7289 (N_7289,N_7165,N_7172);
nor U7290 (N_7290,N_7158,N_7134);
or U7291 (N_7291,N_7139,N_7162);
or U7292 (N_7292,N_7197,N_7193);
nand U7293 (N_7293,N_7127,N_7142);
nand U7294 (N_7294,N_7173,N_7121);
or U7295 (N_7295,N_7113,N_7101);
and U7296 (N_7296,N_7127,N_7116);
or U7297 (N_7297,N_7179,N_7166);
nor U7298 (N_7298,N_7151,N_7190);
nand U7299 (N_7299,N_7104,N_7195);
nor U7300 (N_7300,N_7282,N_7221);
nand U7301 (N_7301,N_7239,N_7281);
nand U7302 (N_7302,N_7277,N_7276);
nor U7303 (N_7303,N_7238,N_7257);
or U7304 (N_7304,N_7285,N_7270);
nor U7305 (N_7305,N_7283,N_7228);
nor U7306 (N_7306,N_7268,N_7290);
nand U7307 (N_7307,N_7294,N_7229);
xnor U7308 (N_7308,N_7200,N_7253);
or U7309 (N_7309,N_7272,N_7234);
or U7310 (N_7310,N_7288,N_7237);
nor U7311 (N_7311,N_7224,N_7291);
or U7312 (N_7312,N_7211,N_7261);
or U7313 (N_7313,N_7254,N_7255);
nor U7314 (N_7314,N_7271,N_7274);
and U7315 (N_7315,N_7289,N_7226);
or U7316 (N_7316,N_7202,N_7215);
and U7317 (N_7317,N_7246,N_7292);
or U7318 (N_7318,N_7262,N_7293);
and U7319 (N_7319,N_7218,N_7236);
xnor U7320 (N_7320,N_7258,N_7233);
or U7321 (N_7321,N_7212,N_7230);
and U7322 (N_7322,N_7280,N_7204);
and U7323 (N_7323,N_7269,N_7278);
nor U7324 (N_7324,N_7243,N_7256);
and U7325 (N_7325,N_7273,N_7235);
or U7326 (N_7326,N_7264,N_7249);
nand U7327 (N_7327,N_7208,N_7203);
nand U7328 (N_7328,N_7297,N_7265);
or U7329 (N_7329,N_7263,N_7284);
or U7330 (N_7330,N_7286,N_7279);
xor U7331 (N_7331,N_7207,N_7259);
nor U7332 (N_7332,N_7251,N_7205);
nand U7333 (N_7333,N_7210,N_7247);
or U7334 (N_7334,N_7260,N_7244);
nor U7335 (N_7335,N_7223,N_7232);
nor U7336 (N_7336,N_7222,N_7298);
nor U7337 (N_7337,N_7241,N_7240);
or U7338 (N_7338,N_7213,N_7242);
and U7339 (N_7339,N_7296,N_7299);
or U7340 (N_7340,N_7245,N_7248);
nand U7341 (N_7341,N_7219,N_7227);
and U7342 (N_7342,N_7231,N_7209);
nor U7343 (N_7343,N_7217,N_7220);
or U7344 (N_7344,N_7225,N_7206);
or U7345 (N_7345,N_7250,N_7201);
or U7346 (N_7346,N_7252,N_7216);
and U7347 (N_7347,N_7214,N_7295);
or U7348 (N_7348,N_7287,N_7267);
nor U7349 (N_7349,N_7266,N_7275);
and U7350 (N_7350,N_7237,N_7274);
xnor U7351 (N_7351,N_7288,N_7286);
or U7352 (N_7352,N_7236,N_7231);
nand U7353 (N_7353,N_7243,N_7210);
and U7354 (N_7354,N_7222,N_7272);
nor U7355 (N_7355,N_7209,N_7295);
nor U7356 (N_7356,N_7273,N_7277);
xor U7357 (N_7357,N_7289,N_7275);
xnor U7358 (N_7358,N_7227,N_7257);
or U7359 (N_7359,N_7271,N_7262);
xnor U7360 (N_7360,N_7286,N_7248);
nor U7361 (N_7361,N_7232,N_7217);
nor U7362 (N_7362,N_7284,N_7274);
and U7363 (N_7363,N_7266,N_7276);
nor U7364 (N_7364,N_7256,N_7273);
nand U7365 (N_7365,N_7297,N_7206);
and U7366 (N_7366,N_7205,N_7214);
nand U7367 (N_7367,N_7273,N_7210);
nor U7368 (N_7368,N_7224,N_7217);
xnor U7369 (N_7369,N_7280,N_7212);
xor U7370 (N_7370,N_7293,N_7220);
xor U7371 (N_7371,N_7208,N_7239);
nand U7372 (N_7372,N_7297,N_7228);
xnor U7373 (N_7373,N_7212,N_7285);
nor U7374 (N_7374,N_7233,N_7209);
or U7375 (N_7375,N_7233,N_7257);
and U7376 (N_7376,N_7214,N_7252);
nor U7377 (N_7377,N_7222,N_7266);
or U7378 (N_7378,N_7202,N_7246);
and U7379 (N_7379,N_7269,N_7244);
nor U7380 (N_7380,N_7211,N_7254);
nor U7381 (N_7381,N_7236,N_7258);
and U7382 (N_7382,N_7237,N_7241);
xor U7383 (N_7383,N_7259,N_7213);
or U7384 (N_7384,N_7276,N_7297);
nor U7385 (N_7385,N_7278,N_7234);
nor U7386 (N_7386,N_7252,N_7226);
and U7387 (N_7387,N_7255,N_7273);
nor U7388 (N_7388,N_7279,N_7243);
or U7389 (N_7389,N_7274,N_7296);
and U7390 (N_7390,N_7245,N_7214);
xor U7391 (N_7391,N_7220,N_7249);
or U7392 (N_7392,N_7283,N_7282);
nor U7393 (N_7393,N_7282,N_7238);
and U7394 (N_7394,N_7201,N_7233);
and U7395 (N_7395,N_7296,N_7268);
or U7396 (N_7396,N_7277,N_7258);
and U7397 (N_7397,N_7273,N_7289);
nor U7398 (N_7398,N_7250,N_7212);
nor U7399 (N_7399,N_7294,N_7227);
xnor U7400 (N_7400,N_7377,N_7394);
and U7401 (N_7401,N_7326,N_7334);
nor U7402 (N_7402,N_7353,N_7389);
and U7403 (N_7403,N_7381,N_7384);
nor U7404 (N_7404,N_7305,N_7320);
and U7405 (N_7405,N_7312,N_7309);
or U7406 (N_7406,N_7348,N_7380);
nand U7407 (N_7407,N_7374,N_7361);
or U7408 (N_7408,N_7393,N_7330);
or U7409 (N_7409,N_7378,N_7335);
nor U7410 (N_7410,N_7338,N_7342);
nor U7411 (N_7411,N_7355,N_7316);
or U7412 (N_7412,N_7367,N_7368);
or U7413 (N_7413,N_7391,N_7302);
xor U7414 (N_7414,N_7336,N_7333);
xnor U7415 (N_7415,N_7369,N_7352);
nand U7416 (N_7416,N_7346,N_7351);
and U7417 (N_7417,N_7366,N_7313);
and U7418 (N_7418,N_7371,N_7379);
nand U7419 (N_7419,N_7318,N_7347);
or U7420 (N_7420,N_7360,N_7325);
nor U7421 (N_7421,N_7306,N_7395);
xor U7422 (N_7422,N_7388,N_7344);
and U7423 (N_7423,N_7300,N_7383);
and U7424 (N_7424,N_7373,N_7396);
or U7425 (N_7425,N_7328,N_7358);
xor U7426 (N_7426,N_7314,N_7362);
nor U7427 (N_7427,N_7324,N_7390);
or U7428 (N_7428,N_7340,N_7365);
and U7429 (N_7429,N_7304,N_7399);
or U7430 (N_7430,N_7331,N_7397);
nor U7431 (N_7431,N_7308,N_7341);
nor U7432 (N_7432,N_7339,N_7359);
or U7433 (N_7433,N_7376,N_7349);
xnor U7434 (N_7434,N_7322,N_7387);
or U7435 (N_7435,N_7321,N_7343);
nand U7436 (N_7436,N_7385,N_7317);
or U7437 (N_7437,N_7332,N_7363);
nor U7438 (N_7438,N_7370,N_7356);
nor U7439 (N_7439,N_7392,N_7327);
nor U7440 (N_7440,N_7301,N_7345);
nor U7441 (N_7441,N_7319,N_7307);
or U7442 (N_7442,N_7323,N_7303);
and U7443 (N_7443,N_7329,N_7382);
xor U7444 (N_7444,N_7364,N_7350);
and U7445 (N_7445,N_7315,N_7311);
or U7446 (N_7446,N_7398,N_7372);
and U7447 (N_7447,N_7337,N_7357);
and U7448 (N_7448,N_7354,N_7375);
or U7449 (N_7449,N_7386,N_7310);
nand U7450 (N_7450,N_7385,N_7387);
or U7451 (N_7451,N_7324,N_7380);
nor U7452 (N_7452,N_7387,N_7344);
nand U7453 (N_7453,N_7307,N_7380);
or U7454 (N_7454,N_7311,N_7380);
nand U7455 (N_7455,N_7390,N_7327);
and U7456 (N_7456,N_7369,N_7399);
and U7457 (N_7457,N_7361,N_7399);
or U7458 (N_7458,N_7316,N_7368);
nand U7459 (N_7459,N_7362,N_7337);
nor U7460 (N_7460,N_7391,N_7324);
or U7461 (N_7461,N_7380,N_7304);
nor U7462 (N_7462,N_7386,N_7349);
and U7463 (N_7463,N_7388,N_7315);
xor U7464 (N_7464,N_7325,N_7389);
or U7465 (N_7465,N_7307,N_7344);
and U7466 (N_7466,N_7313,N_7394);
or U7467 (N_7467,N_7337,N_7312);
nor U7468 (N_7468,N_7317,N_7316);
and U7469 (N_7469,N_7366,N_7385);
or U7470 (N_7470,N_7319,N_7370);
nand U7471 (N_7471,N_7370,N_7342);
nand U7472 (N_7472,N_7376,N_7387);
or U7473 (N_7473,N_7375,N_7391);
and U7474 (N_7474,N_7399,N_7345);
nand U7475 (N_7475,N_7322,N_7344);
nor U7476 (N_7476,N_7341,N_7357);
nor U7477 (N_7477,N_7339,N_7315);
and U7478 (N_7478,N_7391,N_7343);
and U7479 (N_7479,N_7312,N_7390);
nand U7480 (N_7480,N_7397,N_7330);
nor U7481 (N_7481,N_7372,N_7311);
xor U7482 (N_7482,N_7322,N_7305);
nor U7483 (N_7483,N_7388,N_7384);
and U7484 (N_7484,N_7351,N_7301);
or U7485 (N_7485,N_7398,N_7303);
nor U7486 (N_7486,N_7326,N_7384);
nor U7487 (N_7487,N_7321,N_7373);
nor U7488 (N_7488,N_7334,N_7395);
and U7489 (N_7489,N_7308,N_7356);
nand U7490 (N_7490,N_7377,N_7384);
or U7491 (N_7491,N_7384,N_7315);
xnor U7492 (N_7492,N_7351,N_7392);
nor U7493 (N_7493,N_7330,N_7372);
or U7494 (N_7494,N_7305,N_7369);
or U7495 (N_7495,N_7379,N_7390);
nor U7496 (N_7496,N_7384,N_7312);
nand U7497 (N_7497,N_7362,N_7325);
nand U7498 (N_7498,N_7335,N_7334);
nand U7499 (N_7499,N_7333,N_7359);
and U7500 (N_7500,N_7450,N_7479);
nand U7501 (N_7501,N_7417,N_7432);
nor U7502 (N_7502,N_7464,N_7428);
and U7503 (N_7503,N_7433,N_7494);
nand U7504 (N_7504,N_7405,N_7459);
or U7505 (N_7505,N_7408,N_7401);
nand U7506 (N_7506,N_7430,N_7447);
nor U7507 (N_7507,N_7483,N_7423);
nor U7508 (N_7508,N_7468,N_7434);
nand U7509 (N_7509,N_7467,N_7498);
or U7510 (N_7510,N_7427,N_7488);
or U7511 (N_7511,N_7424,N_7478);
nor U7512 (N_7512,N_7403,N_7462);
nand U7513 (N_7513,N_7416,N_7487);
nor U7514 (N_7514,N_7465,N_7490);
nor U7515 (N_7515,N_7407,N_7472);
nand U7516 (N_7516,N_7446,N_7457);
xnor U7517 (N_7517,N_7481,N_7466);
nor U7518 (N_7518,N_7497,N_7471);
nand U7519 (N_7519,N_7449,N_7480);
nor U7520 (N_7520,N_7435,N_7469);
nor U7521 (N_7521,N_7422,N_7413);
or U7522 (N_7522,N_7489,N_7453);
and U7523 (N_7523,N_7456,N_7414);
and U7524 (N_7524,N_7444,N_7418);
and U7525 (N_7525,N_7491,N_7460);
and U7526 (N_7526,N_7470,N_7426);
and U7527 (N_7527,N_7402,N_7440);
nand U7528 (N_7528,N_7454,N_7441);
and U7529 (N_7529,N_7419,N_7429);
nand U7530 (N_7530,N_7437,N_7486);
nand U7531 (N_7531,N_7448,N_7421);
nor U7532 (N_7532,N_7476,N_7436);
nand U7533 (N_7533,N_7425,N_7482);
nand U7534 (N_7534,N_7431,N_7493);
or U7535 (N_7535,N_7475,N_7499);
and U7536 (N_7536,N_7410,N_7461);
and U7537 (N_7537,N_7477,N_7443);
nand U7538 (N_7538,N_7484,N_7406);
nand U7539 (N_7539,N_7445,N_7451);
and U7540 (N_7540,N_7442,N_7412);
nand U7541 (N_7541,N_7485,N_7474);
nor U7542 (N_7542,N_7411,N_7415);
nand U7543 (N_7543,N_7495,N_7458);
xor U7544 (N_7544,N_7404,N_7439);
and U7545 (N_7545,N_7452,N_7492);
nor U7546 (N_7546,N_7473,N_7455);
or U7547 (N_7547,N_7420,N_7438);
nor U7548 (N_7548,N_7409,N_7496);
nor U7549 (N_7549,N_7463,N_7400);
or U7550 (N_7550,N_7403,N_7425);
or U7551 (N_7551,N_7425,N_7454);
nand U7552 (N_7552,N_7498,N_7409);
or U7553 (N_7553,N_7429,N_7495);
nand U7554 (N_7554,N_7416,N_7420);
or U7555 (N_7555,N_7483,N_7435);
and U7556 (N_7556,N_7444,N_7429);
xnor U7557 (N_7557,N_7400,N_7495);
xor U7558 (N_7558,N_7406,N_7481);
and U7559 (N_7559,N_7419,N_7405);
and U7560 (N_7560,N_7408,N_7451);
or U7561 (N_7561,N_7416,N_7451);
nor U7562 (N_7562,N_7416,N_7462);
nor U7563 (N_7563,N_7468,N_7447);
xor U7564 (N_7564,N_7450,N_7480);
or U7565 (N_7565,N_7415,N_7449);
xnor U7566 (N_7566,N_7454,N_7424);
or U7567 (N_7567,N_7499,N_7470);
nor U7568 (N_7568,N_7483,N_7448);
nand U7569 (N_7569,N_7418,N_7487);
or U7570 (N_7570,N_7467,N_7487);
nand U7571 (N_7571,N_7448,N_7462);
nand U7572 (N_7572,N_7435,N_7499);
and U7573 (N_7573,N_7418,N_7428);
nand U7574 (N_7574,N_7440,N_7437);
and U7575 (N_7575,N_7458,N_7423);
xor U7576 (N_7576,N_7474,N_7460);
nor U7577 (N_7577,N_7436,N_7427);
and U7578 (N_7578,N_7417,N_7468);
xnor U7579 (N_7579,N_7489,N_7495);
or U7580 (N_7580,N_7417,N_7496);
or U7581 (N_7581,N_7453,N_7497);
nor U7582 (N_7582,N_7462,N_7434);
nand U7583 (N_7583,N_7415,N_7412);
or U7584 (N_7584,N_7474,N_7495);
nor U7585 (N_7585,N_7421,N_7411);
nor U7586 (N_7586,N_7490,N_7443);
nand U7587 (N_7587,N_7438,N_7492);
or U7588 (N_7588,N_7490,N_7453);
nand U7589 (N_7589,N_7423,N_7401);
and U7590 (N_7590,N_7449,N_7437);
xor U7591 (N_7591,N_7475,N_7439);
or U7592 (N_7592,N_7462,N_7457);
and U7593 (N_7593,N_7400,N_7484);
or U7594 (N_7594,N_7492,N_7499);
xnor U7595 (N_7595,N_7408,N_7404);
and U7596 (N_7596,N_7405,N_7490);
or U7597 (N_7597,N_7458,N_7468);
and U7598 (N_7598,N_7406,N_7492);
and U7599 (N_7599,N_7460,N_7479);
nor U7600 (N_7600,N_7566,N_7551);
nor U7601 (N_7601,N_7582,N_7570);
and U7602 (N_7602,N_7517,N_7554);
nand U7603 (N_7603,N_7539,N_7526);
nand U7604 (N_7604,N_7536,N_7553);
nand U7605 (N_7605,N_7543,N_7569);
and U7606 (N_7606,N_7579,N_7572);
xnor U7607 (N_7607,N_7559,N_7556);
nor U7608 (N_7608,N_7525,N_7518);
nand U7609 (N_7609,N_7509,N_7515);
nor U7610 (N_7610,N_7585,N_7513);
nand U7611 (N_7611,N_7593,N_7598);
xnor U7612 (N_7612,N_7578,N_7519);
or U7613 (N_7613,N_7502,N_7520);
and U7614 (N_7614,N_7589,N_7521);
nor U7615 (N_7615,N_7534,N_7583);
and U7616 (N_7616,N_7562,N_7549);
nor U7617 (N_7617,N_7573,N_7512);
nand U7618 (N_7618,N_7586,N_7596);
or U7619 (N_7619,N_7577,N_7524);
and U7620 (N_7620,N_7587,N_7575);
nor U7621 (N_7621,N_7529,N_7552);
nor U7622 (N_7622,N_7599,N_7584);
and U7623 (N_7623,N_7540,N_7538);
or U7624 (N_7624,N_7581,N_7547);
nand U7625 (N_7625,N_7532,N_7588);
or U7626 (N_7626,N_7507,N_7560);
or U7627 (N_7627,N_7563,N_7537);
or U7628 (N_7628,N_7516,N_7576);
nand U7629 (N_7629,N_7533,N_7503);
nor U7630 (N_7630,N_7592,N_7597);
or U7631 (N_7631,N_7523,N_7541);
and U7632 (N_7632,N_7545,N_7558);
or U7633 (N_7633,N_7506,N_7550);
nor U7634 (N_7634,N_7574,N_7567);
nand U7635 (N_7635,N_7505,N_7564);
or U7636 (N_7636,N_7555,N_7568);
nand U7637 (N_7637,N_7590,N_7528);
nand U7638 (N_7638,N_7527,N_7511);
and U7639 (N_7639,N_7500,N_7514);
and U7640 (N_7640,N_7504,N_7508);
nor U7641 (N_7641,N_7510,N_7571);
xnor U7642 (N_7642,N_7501,N_7594);
or U7643 (N_7643,N_7530,N_7522);
nor U7644 (N_7644,N_7557,N_7542);
or U7645 (N_7645,N_7548,N_7531);
nand U7646 (N_7646,N_7591,N_7595);
and U7647 (N_7647,N_7561,N_7535);
xnor U7648 (N_7648,N_7544,N_7565);
or U7649 (N_7649,N_7580,N_7546);
and U7650 (N_7650,N_7578,N_7557);
xor U7651 (N_7651,N_7523,N_7573);
and U7652 (N_7652,N_7517,N_7511);
or U7653 (N_7653,N_7534,N_7579);
xnor U7654 (N_7654,N_7505,N_7502);
nand U7655 (N_7655,N_7580,N_7570);
and U7656 (N_7656,N_7538,N_7566);
nor U7657 (N_7657,N_7532,N_7515);
or U7658 (N_7658,N_7596,N_7588);
nor U7659 (N_7659,N_7587,N_7516);
and U7660 (N_7660,N_7501,N_7505);
and U7661 (N_7661,N_7520,N_7500);
and U7662 (N_7662,N_7595,N_7507);
nand U7663 (N_7663,N_7592,N_7551);
nand U7664 (N_7664,N_7511,N_7572);
nand U7665 (N_7665,N_7533,N_7516);
and U7666 (N_7666,N_7541,N_7543);
nor U7667 (N_7667,N_7557,N_7500);
and U7668 (N_7668,N_7584,N_7559);
or U7669 (N_7669,N_7533,N_7562);
xor U7670 (N_7670,N_7573,N_7511);
nor U7671 (N_7671,N_7569,N_7532);
xnor U7672 (N_7672,N_7511,N_7509);
or U7673 (N_7673,N_7597,N_7586);
nand U7674 (N_7674,N_7539,N_7561);
and U7675 (N_7675,N_7541,N_7594);
xor U7676 (N_7676,N_7588,N_7526);
and U7677 (N_7677,N_7576,N_7599);
and U7678 (N_7678,N_7581,N_7517);
or U7679 (N_7679,N_7570,N_7577);
and U7680 (N_7680,N_7550,N_7518);
and U7681 (N_7681,N_7569,N_7508);
nor U7682 (N_7682,N_7582,N_7579);
nand U7683 (N_7683,N_7555,N_7515);
nor U7684 (N_7684,N_7558,N_7567);
nand U7685 (N_7685,N_7533,N_7578);
nand U7686 (N_7686,N_7597,N_7588);
or U7687 (N_7687,N_7543,N_7581);
or U7688 (N_7688,N_7503,N_7588);
nand U7689 (N_7689,N_7573,N_7584);
nor U7690 (N_7690,N_7568,N_7515);
or U7691 (N_7691,N_7569,N_7519);
and U7692 (N_7692,N_7590,N_7506);
and U7693 (N_7693,N_7589,N_7550);
nand U7694 (N_7694,N_7583,N_7573);
xor U7695 (N_7695,N_7591,N_7554);
nand U7696 (N_7696,N_7586,N_7508);
nor U7697 (N_7697,N_7581,N_7520);
or U7698 (N_7698,N_7553,N_7567);
nand U7699 (N_7699,N_7520,N_7588);
nand U7700 (N_7700,N_7604,N_7639);
nor U7701 (N_7701,N_7697,N_7682);
and U7702 (N_7702,N_7642,N_7654);
nor U7703 (N_7703,N_7641,N_7626);
nand U7704 (N_7704,N_7600,N_7645);
xor U7705 (N_7705,N_7629,N_7653);
and U7706 (N_7706,N_7649,N_7655);
nor U7707 (N_7707,N_7662,N_7637);
and U7708 (N_7708,N_7620,N_7610);
nor U7709 (N_7709,N_7699,N_7606);
and U7710 (N_7710,N_7621,N_7613);
and U7711 (N_7711,N_7681,N_7677);
and U7712 (N_7712,N_7686,N_7674);
nand U7713 (N_7713,N_7638,N_7602);
nor U7714 (N_7714,N_7651,N_7625);
or U7715 (N_7715,N_7663,N_7688);
nand U7716 (N_7716,N_7648,N_7694);
or U7717 (N_7717,N_7658,N_7672);
and U7718 (N_7718,N_7650,N_7673);
nand U7719 (N_7719,N_7670,N_7640);
or U7720 (N_7720,N_7630,N_7689);
or U7721 (N_7721,N_7687,N_7634);
or U7722 (N_7722,N_7685,N_7601);
nand U7723 (N_7723,N_7636,N_7633);
nand U7724 (N_7724,N_7628,N_7659);
nor U7725 (N_7725,N_7647,N_7614);
and U7726 (N_7726,N_7603,N_7656);
nand U7727 (N_7727,N_7657,N_7676);
xor U7728 (N_7728,N_7627,N_7691);
and U7729 (N_7729,N_7679,N_7669);
nand U7730 (N_7730,N_7684,N_7668);
and U7731 (N_7731,N_7615,N_7612);
or U7732 (N_7732,N_7607,N_7632);
or U7733 (N_7733,N_7609,N_7611);
nor U7734 (N_7734,N_7666,N_7678);
xor U7735 (N_7735,N_7665,N_7646);
and U7736 (N_7736,N_7661,N_7692);
or U7737 (N_7737,N_7690,N_7683);
nand U7738 (N_7738,N_7605,N_7631);
and U7739 (N_7739,N_7617,N_7618);
and U7740 (N_7740,N_7644,N_7680);
or U7741 (N_7741,N_7698,N_7695);
nand U7742 (N_7742,N_7693,N_7608);
nand U7743 (N_7743,N_7624,N_7623);
and U7744 (N_7744,N_7619,N_7664);
and U7745 (N_7745,N_7675,N_7616);
nand U7746 (N_7746,N_7652,N_7696);
nand U7747 (N_7747,N_7660,N_7622);
nand U7748 (N_7748,N_7667,N_7643);
nor U7749 (N_7749,N_7671,N_7635);
nand U7750 (N_7750,N_7669,N_7622);
or U7751 (N_7751,N_7630,N_7602);
nor U7752 (N_7752,N_7655,N_7604);
nor U7753 (N_7753,N_7633,N_7655);
nor U7754 (N_7754,N_7612,N_7657);
xnor U7755 (N_7755,N_7655,N_7644);
nor U7756 (N_7756,N_7678,N_7637);
and U7757 (N_7757,N_7689,N_7685);
and U7758 (N_7758,N_7666,N_7671);
nand U7759 (N_7759,N_7684,N_7603);
and U7760 (N_7760,N_7613,N_7697);
or U7761 (N_7761,N_7662,N_7638);
and U7762 (N_7762,N_7658,N_7660);
nand U7763 (N_7763,N_7659,N_7682);
nand U7764 (N_7764,N_7614,N_7621);
nor U7765 (N_7765,N_7620,N_7654);
xnor U7766 (N_7766,N_7682,N_7621);
or U7767 (N_7767,N_7607,N_7613);
nor U7768 (N_7768,N_7691,N_7609);
xor U7769 (N_7769,N_7690,N_7621);
or U7770 (N_7770,N_7653,N_7660);
or U7771 (N_7771,N_7635,N_7616);
nand U7772 (N_7772,N_7640,N_7673);
xnor U7773 (N_7773,N_7635,N_7623);
nand U7774 (N_7774,N_7645,N_7699);
or U7775 (N_7775,N_7621,N_7657);
and U7776 (N_7776,N_7668,N_7699);
nand U7777 (N_7777,N_7649,N_7676);
or U7778 (N_7778,N_7673,N_7652);
nand U7779 (N_7779,N_7649,N_7669);
and U7780 (N_7780,N_7621,N_7600);
nand U7781 (N_7781,N_7666,N_7698);
or U7782 (N_7782,N_7685,N_7686);
or U7783 (N_7783,N_7695,N_7655);
or U7784 (N_7784,N_7669,N_7626);
and U7785 (N_7785,N_7612,N_7617);
or U7786 (N_7786,N_7685,N_7634);
or U7787 (N_7787,N_7611,N_7605);
or U7788 (N_7788,N_7673,N_7632);
or U7789 (N_7789,N_7605,N_7625);
and U7790 (N_7790,N_7643,N_7618);
nand U7791 (N_7791,N_7617,N_7608);
nor U7792 (N_7792,N_7678,N_7665);
or U7793 (N_7793,N_7616,N_7699);
xnor U7794 (N_7794,N_7661,N_7651);
and U7795 (N_7795,N_7615,N_7653);
nand U7796 (N_7796,N_7676,N_7626);
or U7797 (N_7797,N_7670,N_7625);
and U7798 (N_7798,N_7653,N_7684);
and U7799 (N_7799,N_7608,N_7648);
nand U7800 (N_7800,N_7788,N_7757);
xor U7801 (N_7801,N_7716,N_7797);
and U7802 (N_7802,N_7764,N_7735);
nor U7803 (N_7803,N_7765,N_7751);
nor U7804 (N_7804,N_7710,N_7772);
and U7805 (N_7805,N_7776,N_7793);
or U7806 (N_7806,N_7774,N_7719);
xor U7807 (N_7807,N_7707,N_7726);
nor U7808 (N_7808,N_7727,N_7705);
nor U7809 (N_7809,N_7742,N_7703);
and U7810 (N_7810,N_7766,N_7701);
and U7811 (N_7811,N_7775,N_7796);
and U7812 (N_7812,N_7739,N_7784);
nor U7813 (N_7813,N_7773,N_7744);
nor U7814 (N_7814,N_7768,N_7758);
nor U7815 (N_7815,N_7732,N_7760);
xor U7816 (N_7816,N_7740,N_7791);
or U7817 (N_7817,N_7771,N_7725);
or U7818 (N_7818,N_7749,N_7741);
and U7819 (N_7819,N_7702,N_7754);
nor U7820 (N_7820,N_7730,N_7779);
or U7821 (N_7821,N_7728,N_7763);
nor U7822 (N_7822,N_7718,N_7745);
or U7823 (N_7823,N_7715,N_7746);
nand U7824 (N_7824,N_7790,N_7706);
nor U7825 (N_7825,N_7756,N_7700);
nand U7826 (N_7826,N_7759,N_7798);
or U7827 (N_7827,N_7787,N_7712);
or U7828 (N_7828,N_7792,N_7781);
or U7829 (N_7829,N_7769,N_7777);
nor U7830 (N_7830,N_7795,N_7722);
xnor U7831 (N_7831,N_7720,N_7724);
nand U7832 (N_7832,N_7721,N_7729);
or U7833 (N_7833,N_7780,N_7708);
nor U7834 (N_7834,N_7783,N_7753);
or U7835 (N_7835,N_7737,N_7778);
or U7836 (N_7836,N_7755,N_7717);
or U7837 (N_7837,N_7709,N_7734);
nor U7838 (N_7838,N_7711,N_7733);
nand U7839 (N_7839,N_7767,N_7785);
nand U7840 (N_7840,N_7743,N_7752);
nor U7841 (N_7841,N_7786,N_7799);
xnor U7842 (N_7842,N_7714,N_7736);
and U7843 (N_7843,N_7748,N_7713);
or U7844 (N_7844,N_7794,N_7762);
or U7845 (N_7845,N_7723,N_7750);
nor U7846 (N_7846,N_7782,N_7738);
or U7847 (N_7847,N_7731,N_7761);
nor U7848 (N_7848,N_7747,N_7789);
and U7849 (N_7849,N_7770,N_7704);
nor U7850 (N_7850,N_7778,N_7712);
nand U7851 (N_7851,N_7749,N_7733);
or U7852 (N_7852,N_7796,N_7784);
nor U7853 (N_7853,N_7770,N_7782);
and U7854 (N_7854,N_7779,N_7796);
nand U7855 (N_7855,N_7768,N_7708);
xnor U7856 (N_7856,N_7743,N_7793);
nor U7857 (N_7857,N_7775,N_7724);
and U7858 (N_7858,N_7713,N_7740);
or U7859 (N_7859,N_7719,N_7738);
and U7860 (N_7860,N_7722,N_7744);
nor U7861 (N_7861,N_7752,N_7737);
nand U7862 (N_7862,N_7791,N_7796);
or U7863 (N_7863,N_7753,N_7775);
nor U7864 (N_7864,N_7758,N_7780);
nor U7865 (N_7865,N_7776,N_7782);
and U7866 (N_7866,N_7741,N_7791);
and U7867 (N_7867,N_7739,N_7707);
nand U7868 (N_7868,N_7789,N_7783);
or U7869 (N_7869,N_7735,N_7778);
or U7870 (N_7870,N_7760,N_7765);
and U7871 (N_7871,N_7786,N_7773);
nor U7872 (N_7872,N_7736,N_7775);
or U7873 (N_7873,N_7745,N_7734);
nand U7874 (N_7874,N_7736,N_7783);
xnor U7875 (N_7875,N_7755,N_7785);
or U7876 (N_7876,N_7754,N_7705);
nor U7877 (N_7877,N_7751,N_7717);
and U7878 (N_7878,N_7759,N_7732);
nand U7879 (N_7879,N_7737,N_7749);
nor U7880 (N_7880,N_7721,N_7740);
or U7881 (N_7881,N_7753,N_7747);
nand U7882 (N_7882,N_7784,N_7705);
or U7883 (N_7883,N_7783,N_7786);
and U7884 (N_7884,N_7742,N_7792);
nand U7885 (N_7885,N_7777,N_7733);
nand U7886 (N_7886,N_7725,N_7739);
nand U7887 (N_7887,N_7734,N_7756);
and U7888 (N_7888,N_7743,N_7745);
or U7889 (N_7889,N_7763,N_7714);
and U7890 (N_7890,N_7763,N_7756);
or U7891 (N_7891,N_7776,N_7735);
nand U7892 (N_7892,N_7724,N_7735);
nand U7893 (N_7893,N_7728,N_7726);
or U7894 (N_7894,N_7714,N_7790);
nand U7895 (N_7895,N_7786,N_7792);
or U7896 (N_7896,N_7734,N_7771);
nor U7897 (N_7897,N_7723,N_7720);
nor U7898 (N_7898,N_7754,N_7796);
or U7899 (N_7899,N_7726,N_7779);
nand U7900 (N_7900,N_7860,N_7833);
nor U7901 (N_7901,N_7864,N_7850);
and U7902 (N_7902,N_7802,N_7861);
and U7903 (N_7903,N_7865,N_7818);
nand U7904 (N_7904,N_7893,N_7846);
nand U7905 (N_7905,N_7877,N_7896);
nand U7906 (N_7906,N_7817,N_7819);
nand U7907 (N_7907,N_7862,N_7807);
nor U7908 (N_7908,N_7886,N_7863);
nor U7909 (N_7909,N_7898,N_7866);
and U7910 (N_7910,N_7825,N_7822);
and U7911 (N_7911,N_7867,N_7851);
xor U7912 (N_7912,N_7872,N_7858);
or U7913 (N_7913,N_7838,N_7823);
or U7914 (N_7914,N_7891,N_7880);
nor U7915 (N_7915,N_7837,N_7852);
or U7916 (N_7916,N_7814,N_7804);
xnor U7917 (N_7917,N_7813,N_7868);
and U7918 (N_7918,N_7879,N_7839);
or U7919 (N_7919,N_7841,N_7847);
or U7920 (N_7920,N_7812,N_7844);
nor U7921 (N_7921,N_7845,N_7894);
and U7922 (N_7922,N_7800,N_7801);
or U7923 (N_7923,N_7897,N_7869);
or U7924 (N_7924,N_7826,N_7855);
nand U7925 (N_7925,N_7840,N_7854);
nor U7926 (N_7926,N_7848,N_7883);
and U7927 (N_7927,N_7889,N_7873);
nor U7928 (N_7928,N_7824,N_7871);
and U7929 (N_7929,N_7853,N_7878);
or U7930 (N_7930,N_7842,N_7816);
or U7931 (N_7931,N_7820,N_7810);
and U7932 (N_7932,N_7888,N_7887);
and U7933 (N_7933,N_7890,N_7835);
or U7934 (N_7934,N_7827,N_7808);
nand U7935 (N_7935,N_7834,N_7859);
nand U7936 (N_7936,N_7806,N_7831);
and U7937 (N_7937,N_7885,N_7805);
or U7938 (N_7938,N_7815,N_7836);
nor U7939 (N_7939,N_7803,N_7828);
xor U7940 (N_7940,N_7899,N_7875);
or U7941 (N_7941,N_7870,N_7809);
nand U7942 (N_7942,N_7843,N_7881);
or U7943 (N_7943,N_7876,N_7882);
nand U7944 (N_7944,N_7849,N_7884);
nor U7945 (N_7945,N_7892,N_7821);
nor U7946 (N_7946,N_7895,N_7829);
or U7947 (N_7947,N_7811,N_7832);
or U7948 (N_7948,N_7856,N_7830);
or U7949 (N_7949,N_7857,N_7874);
nand U7950 (N_7950,N_7872,N_7845);
or U7951 (N_7951,N_7844,N_7855);
xor U7952 (N_7952,N_7894,N_7841);
nor U7953 (N_7953,N_7894,N_7898);
or U7954 (N_7954,N_7813,N_7821);
nor U7955 (N_7955,N_7855,N_7843);
nor U7956 (N_7956,N_7831,N_7807);
and U7957 (N_7957,N_7886,N_7888);
or U7958 (N_7958,N_7892,N_7802);
and U7959 (N_7959,N_7881,N_7850);
xnor U7960 (N_7960,N_7808,N_7872);
xnor U7961 (N_7961,N_7898,N_7825);
nor U7962 (N_7962,N_7855,N_7813);
and U7963 (N_7963,N_7874,N_7822);
or U7964 (N_7964,N_7880,N_7830);
xor U7965 (N_7965,N_7801,N_7896);
and U7966 (N_7966,N_7864,N_7808);
xor U7967 (N_7967,N_7829,N_7821);
or U7968 (N_7968,N_7877,N_7881);
nand U7969 (N_7969,N_7897,N_7867);
or U7970 (N_7970,N_7890,N_7801);
or U7971 (N_7971,N_7894,N_7850);
nor U7972 (N_7972,N_7838,N_7895);
nor U7973 (N_7973,N_7829,N_7834);
nand U7974 (N_7974,N_7840,N_7891);
or U7975 (N_7975,N_7878,N_7891);
or U7976 (N_7976,N_7824,N_7886);
nor U7977 (N_7977,N_7807,N_7876);
nand U7978 (N_7978,N_7893,N_7844);
nand U7979 (N_7979,N_7898,N_7821);
nand U7980 (N_7980,N_7889,N_7822);
and U7981 (N_7981,N_7879,N_7885);
nand U7982 (N_7982,N_7835,N_7848);
and U7983 (N_7983,N_7870,N_7817);
nor U7984 (N_7984,N_7881,N_7815);
nor U7985 (N_7985,N_7851,N_7844);
or U7986 (N_7986,N_7895,N_7817);
xnor U7987 (N_7987,N_7813,N_7895);
or U7988 (N_7988,N_7826,N_7880);
nand U7989 (N_7989,N_7838,N_7858);
or U7990 (N_7990,N_7817,N_7844);
xor U7991 (N_7991,N_7898,N_7802);
nor U7992 (N_7992,N_7883,N_7863);
or U7993 (N_7993,N_7853,N_7805);
xnor U7994 (N_7994,N_7894,N_7804);
nand U7995 (N_7995,N_7824,N_7817);
nand U7996 (N_7996,N_7864,N_7812);
nand U7997 (N_7997,N_7848,N_7849);
and U7998 (N_7998,N_7806,N_7896);
and U7999 (N_7999,N_7877,N_7883);
and U8000 (N_8000,N_7924,N_7974);
nor U8001 (N_8001,N_7953,N_7968);
and U8002 (N_8002,N_7929,N_7905);
nor U8003 (N_8003,N_7933,N_7981);
xor U8004 (N_8004,N_7900,N_7993);
or U8005 (N_8005,N_7962,N_7951);
or U8006 (N_8006,N_7944,N_7921);
and U8007 (N_8007,N_7927,N_7932);
or U8008 (N_8008,N_7918,N_7965);
or U8009 (N_8009,N_7903,N_7961);
xnor U8010 (N_8010,N_7997,N_7907);
nor U8011 (N_8011,N_7941,N_7922);
and U8012 (N_8012,N_7919,N_7948);
and U8013 (N_8013,N_7958,N_7998);
nor U8014 (N_8014,N_7980,N_7964);
nor U8015 (N_8015,N_7988,N_7901);
and U8016 (N_8016,N_7970,N_7912);
nand U8017 (N_8017,N_7963,N_7913);
nand U8018 (N_8018,N_7934,N_7954);
and U8019 (N_8019,N_7943,N_7979);
or U8020 (N_8020,N_7952,N_7940);
or U8021 (N_8021,N_7914,N_7978);
nor U8022 (N_8022,N_7936,N_7931);
nand U8023 (N_8023,N_7902,N_7917);
nor U8024 (N_8024,N_7908,N_7996);
and U8025 (N_8025,N_7925,N_7976);
nand U8026 (N_8026,N_7911,N_7960);
nand U8027 (N_8027,N_7949,N_7984);
nand U8028 (N_8028,N_7906,N_7969);
xnor U8029 (N_8029,N_7938,N_7910);
or U8030 (N_8030,N_7977,N_7947);
nor U8031 (N_8031,N_7937,N_7994);
and U8032 (N_8032,N_7930,N_7923);
and U8033 (N_8033,N_7942,N_7975);
nor U8034 (N_8034,N_7946,N_7986);
nand U8035 (N_8035,N_7928,N_7985);
or U8036 (N_8036,N_7973,N_7916);
nor U8037 (N_8037,N_7956,N_7955);
xnor U8038 (N_8038,N_7959,N_7983);
nor U8039 (N_8039,N_7909,N_7999);
nor U8040 (N_8040,N_7967,N_7915);
nand U8041 (N_8041,N_7995,N_7992);
xor U8042 (N_8042,N_7939,N_7966);
and U8043 (N_8043,N_7971,N_7920);
nand U8044 (N_8044,N_7989,N_7904);
nand U8045 (N_8045,N_7990,N_7987);
or U8046 (N_8046,N_7935,N_7945);
or U8047 (N_8047,N_7950,N_7972);
or U8048 (N_8048,N_7957,N_7991);
and U8049 (N_8049,N_7982,N_7926);
nor U8050 (N_8050,N_7989,N_7930);
nand U8051 (N_8051,N_7967,N_7994);
nand U8052 (N_8052,N_7944,N_7949);
nand U8053 (N_8053,N_7958,N_7971);
nand U8054 (N_8054,N_7935,N_7911);
and U8055 (N_8055,N_7927,N_7962);
and U8056 (N_8056,N_7999,N_7978);
xor U8057 (N_8057,N_7978,N_7991);
or U8058 (N_8058,N_7906,N_7988);
and U8059 (N_8059,N_7958,N_7985);
nor U8060 (N_8060,N_7921,N_7906);
nor U8061 (N_8061,N_7961,N_7965);
xor U8062 (N_8062,N_7961,N_7900);
and U8063 (N_8063,N_7941,N_7919);
nand U8064 (N_8064,N_7958,N_7959);
and U8065 (N_8065,N_7906,N_7930);
or U8066 (N_8066,N_7928,N_7907);
nand U8067 (N_8067,N_7952,N_7992);
nor U8068 (N_8068,N_7998,N_7995);
or U8069 (N_8069,N_7955,N_7949);
or U8070 (N_8070,N_7933,N_7958);
or U8071 (N_8071,N_7946,N_7955);
or U8072 (N_8072,N_7912,N_7979);
or U8073 (N_8073,N_7985,N_7954);
nor U8074 (N_8074,N_7986,N_7943);
nand U8075 (N_8075,N_7934,N_7949);
and U8076 (N_8076,N_7944,N_7990);
nand U8077 (N_8077,N_7991,N_7910);
and U8078 (N_8078,N_7934,N_7999);
xnor U8079 (N_8079,N_7981,N_7998);
nand U8080 (N_8080,N_7983,N_7997);
nor U8081 (N_8081,N_7959,N_7925);
xnor U8082 (N_8082,N_7974,N_7906);
nor U8083 (N_8083,N_7917,N_7920);
nand U8084 (N_8084,N_7942,N_7928);
nor U8085 (N_8085,N_7980,N_7931);
or U8086 (N_8086,N_7943,N_7997);
or U8087 (N_8087,N_7959,N_7987);
nand U8088 (N_8088,N_7982,N_7921);
and U8089 (N_8089,N_7975,N_7993);
nand U8090 (N_8090,N_7972,N_7981);
nand U8091 (N_8091,N_7935,N_7902);
xnor U8092 (N_8092,N_7966,N_7985);
nor U8093 (N_8093,N_7920,N_7949);
nand U8094 (N_8094,N_7947,N_7916);
nand U8095 (N_8095,N_7959,N_7970);
nor U8096 (N_8096,N_7980,N_7934);
nor U8097 (N_8097,N_7919,N_7949);
nor U8098 (N_8098,N_7939,N_7901);
or U8099 (N_8099,N_7986,N_7944);
nor U8100 (N_8100,N_8067,N_8099);
and U8101 (N_8101,N_8020,N_8062);
xor U8102 (N_8102,N_8043,N_8077);
and U8103 (N_8103,N_8078,N_8048);
nand U8104 (N_8104,N_8071,N_8083);
nor U8105 (N_8105,N_8065,N_8028);
nor U8106 (N_8106,N_8091,N_8021);
xor U8107 (N_8107,N_8079,N_8055);
nand U8108 (N_8108,N_8014,N_8096);
and U8109 (N_8109,N_8093,N_8089);
and U8110 (N_8110,N_8076,N_8004);
nor U8111 (N_8111,N_8049,N_8030);
nand U8112 (N_8112,N_8003,N_8002);
nand U8113 (N_8113,N_8059,N_8061);
nand U8114 (N_8114,N_8086,N_8066);
nor U8115 (N_8115,N_8058,N_8007);
and U8116 (N_8116,N_8025,N_8044);
or U8117 (N_8117,N_8075,N_8070);
and U8118 (N_8118,N_8027,N_8087);
nor U8119 (N_8119,N_8019,N_8050);
nand U8120 (N_8120,N_8045,N_8041);
nand U8121 (N_8121,N_8063,N_8037);
or U8122 (N_8122,N_8094,N_8012);
nand U8123 (N_8123,N_8047,N_8052);
and U8124 (N_8124,N_8046,N_8085);
nor U8125 (N_8125,N_8035,N_8024);
nor U8126 (N_8126,N_8001,N_8064);
nand U8127 (N_8127,N_8074,N_8068);
and U8128 (N_8128,N_8011,N_8092);
nand U8129 (N_8129,N_8010,N_8098);
and U8130 (N_8130,N_8023,N_8097);
xor U8131 (N_8131,N_8032,N_8060);
or U8132 (N_8132,N_8006,N_8081);
and U8133 (N_8133,N_8038,N_8036);
or U8134 (N_8134,N_8082,N_8095);
and U8135 (N_8135,N_8053,N_8031);
xor U8136 (N_8136,N_8051,N_8016);
and U8137 (N_8137,N_8042,N_8017);
nor U8138 (N_8138,N_8073,N_8040);
nand U8139 (N_8139,N_8084,N_8057);
nand U8140 (N_8140,N_8034,N_8039);
nor U8141 (N_8141,N_8015,N_8008);
and U8142 (N_8142,N_8080,N_8009);
or U8143 (N_8143,N_8056,N_8022);
or U8144 (N_8144,N_8026,N_8069);
or U8145 (N_8145,N_8013,N_8088);
or U8146 (N_8146,N_8005,N_8090);
or U8147 (N_8147,N_8054,N_8033);
nor U8148 (N_8148,N_8018,N_8072);
nor U8149 (N_8149,N_8029,N_8000);
and U8150 (N_8150,N_8098,N_8024);
nor U8151 (N_8151,N_8071,N_8027);
and U8152 (N_8152,N_8045,N_8064);
nor U8153 (N_8153,N_8029,N_8016);
nor U8154 (N_8154,N_8063,N_8075);
nor U8155 (N_8155,N_8077,N_8067);
nor U8156 (N_8156,N_8000,N_8048);
or U8157 (N_8157,N_8019,N_8022);
and U8158 (N_8158,N_8005,N_8007);
nand U8159 (N_8159,N_8028,N_8071);
and U8160 (N_8160,N_8051,N_8083);
nor U8161 (N_8161,N_8048,N_8049);
and U8162 (N_8162,N_8019,N_8023);
and U8163 (N_8163,N_8096,N_8077);
and U8164 (N_8164,N_8058,N_8092);
and U8165 (N_8165,N_8062,N_8097);
nand U8166 (N_8166,N_8084,N_8070);
nor U8167 (N_8167,N_8078,N_8068);
or U8168 (N_8168,N_8054,N_8007);
nand U8169 (N_8169,N_8013,N_8007);
nand U8170 (N_8170,N_8072,N_8032);
nor U8171 (N_8171,N_8022,N_8033);
or U8172 (N_8172,N_8023,N_8051);
nand U8173 (N_8173,N_8010,N_8049);
nand U8174 (N_8174,N_8030,N_8007);
nand U8175 (N_8175,N_8030,N_8008);
and U8176 (N_8176,N_8026,N_8092);
or U8177 (N_8177,N_8016,N_8000);
or U8178 (N_8178,N_8076,N_8096);
xnor U8179 (N_8179,N_8013,N_8034);
nor U8180 (N_8180,N_8099,N_8061);
nor U8181 (N_8181,N_8048,N_8093);
or U8182 (N_8182,N_8075,N_8023);
nor U8183 (N_8183,N_8048,N_8001);
or U8184 (N_8184,N_8006,N_8074);
nand U8185 (N_8185,N_8061,N_8006);
and U8186 (N_8186,N_8039,N_8050);
nor U8187 (N_8187,N_8073,N_8045);
nand U8188 (N_8188,N_8092,N_8056);
nor U8189 (N_8189,N_8064,N_8071);
and U8190 (N_8190,N_8037,N_8009);
or U8191 (N_8191,N_8093,N_8017);
xnor U8192 (N_8192,N_8017,N_8085);
and U8193 (N_8193,N_8053,N_8040);
or U8194 (N_8194,N_8090,N_8050);
or U8195 (N_8195,N_8086,N_8035);
or U8196 (N_8196,N_8071,N_8053);
nor U8197 (N_8197,N_8016,N_8086);
xor U8198 (N_8198,N_8075,N_8053);
nor U8199 (N_8199,N_8093,N_8056);
or U8200 (N_8200,N_8158,N_8108);
nor U8201 (N_8201,N_8109,N_8107);
nor U8202 (N_8202,N_8176,N_8140);
nand U8203 (N_8203,N_8187,N_8147);
nand U8204 (N_8204,N_8177,N_8191);
or U8205 (N_8205,N_8123,N_8124);
xnor U8206 (N_8206,N_8153,N_8180);
nor U8207 (N_8207,N_8197,N_8169);
and U8208 (N_8208,N_8145,N_8133);
or U8209 (N_8209,N_8142,N_8154);
or U8210 (N_8210,N_8194,N_8198);
or U8211 (N_8211,N_8164,N_8185);
or U8212 (N_8212,N_8172,N_8183);
nor U8213 (N_8213,N_8152,N_8104);
and U8214 (N_8214,N_8125,N_8193);
and U8215 (N_8215,N_8132,N_8121);
nand U8216 (N_8216,N_8174,N_8114);
nor U8217 (N_8217,N_8106,N_8192);
nor U8218 (N_8218,N_8163,N_8165);
and U8219 (N_8219,N_8186,N_8160);
or U8220 (N_8220,N_8156,N_8157);
and U8221 (N_8221,N_8103,N_8111);
and U8222 (N_8222,N_8162,N_8146);
nor U8223 (N_8223,N_8148,N_8115);
or U8224 (N_8224,N_8127,N_8196);
or U8225 (N_8225,N_8100,N_8113);
nor U8226 (N_8226,N_8155,N_8173);
xor U8227 (N_8227,N_8110,N_8178);
nor U8228 (N_8228,N_8101,N_8116);
and U8229 (N_8229,N_8117,N_8112);
nand U8230 (N_8230,N_8195,N_8167);
nand U8231 (N_8231,N_8141,N_8150);
or U8232 (N_8232,N_8105,N_8134);
nand U8233 (N_8233,N_8199,N_8143);
nand U8234 (N_8234,N_8168,N_8161);
nor U8235 (N_8235,N_8182,N_8138);
or U8236 (N_8236,N_8166,N_8136);
or U8237 (N_8237,N_8189,N_8139);
and U8238 (N_8238,N_8119,N_8122);
nor U8239 (N_8239,N_8144,N_8181);
and U8240 (N_8240,N_8171,N_8149);
nor U8241 (N_8241,N_8175,N_8129);
and U8242 (N_8242,N_8118,N_8184);
xor U8243 (N_8243,N_8137,N_8102);
or U8244 (N_8244,N_8170,N_8130);
and U8245 (N_8245,N_8120,N_8131);
nand U8246 (N_8246,N_8135,N_8128);
and U8247 (N_8247,N_8179,N_8159);
nand U8248 (N_8248,N_8151,N_8126);
nand U8249 (N_8249,N_8190,N_8188);
nor U8250 (N_8250,N_8133,N_8180);
and U8251 (N_8251,N_8140,N_8103);
or U8252 (N_8252,N_8198,N_8151);
nor U8253 (N_8253,N_8154,N_8194);
nor U8254 (N_8254,N_8139,N_8176);
or U8255 (N_8255,N_8197,N_8187);
nand U8256 (N_8256,N_8164,N_8186);
or U8257 (N_8257,N_8149,N_8143);
nand U8258 (N_8258,N_8173,N_8106);
and U8259 (N_8259,N_8108,N_8101);
and U8260 (N_8260,N_8131,N_8154);
or U8261 (N_8261,N_8166,N_8110);
nor U8262 (N_8262,N_8199,N_8145);
xnor U8263 (N_8263,N_8176,N_8187);
or U8264 (N_8264,N_8187,N_8180);
or U8265 (N_8265,N_8189,N_8148);
nand U8266 (N_8266,N_8137,N_8195);
and U8267 (N_8267,N_8178,N_8199);
nor U8268 (N_8268,N_8196,N_8192);
xnor U8269 (N_8269,N_8194,N_8143);
or U8270 (N_8270,N_8164,N_8112);
or U8271 (N_8271,N_8134,N_8139);
and U8272 (N_8272,N_8138,N_8163);
or U8273 (N_8273,N_8111,N_8199);
and U8274 (N_8274,N_8152,N_8101);
xnor U8275 (N_8275,N_8174,N_8117);
nand U8276 (N_8276,N_8128,N_8181);
nand U8277 (N_8277,N_8132,N_8170);
nand U8278 (N_8278,N_8156,N_8102);
nand U8279 (N_8279,N_8148,N_8152);
nand U8280 (N_8280,N_8141,N_8184);
or U8281 (N_8281,N_8150,N_8170);
nand U8282 (N_8282,N_8100,N_8193);
nor U8283 (N_8283,N_8174,N_8198);
nand U8284 (N_8284,N_8122,N_8167);
nand U8285 (N_8285,N_8145,N_8148);
nand U8286 (N_8286,N_8167,N_8197);
xor U8287 (N_8287,N_8182,N_8136);
nor U8288 (N_8288,N_8143,N_8123);
nand U8289 (N_8289,N_8104,N_8140);
and U8290 (N_8290,N_8110,N_8126);
and U8291 (N_8291,N_8199,N_8183);
or U8292 (N_8292,N_8128,N_8173);
and U8293 (N_8293,N_8144,N_8101);
nor U8294 (N_8294,N_8153,N_8145);
nor U8295 (N_8295,N_8149,N_8122);
or U8296 (N_8296,N_8188,N_8101);
or U8297 (N_8297,N_8102,N_8119);
nor U8298 (N_8298,N_8192,N_8163);
or U8299 (N_8299,N_8129,N_8109);
nand U8300 (N_8300,N_8264,N_8230);
xor U8301 (N_8301,N_8266,N_8209);
xnor U8302 (N_8302,N_8261,N_8220);
nand U8303 (N_8303,N_8252,N_8204);
nand U8304 (N_8304,N_8289,N_8295);
nand U8305 (N_8305,N_8211,N_8257);
or U8306 (N_8306,N_8219,N_8288);
nor U8307 (N_8307,N_8286,N_8271);
and U8308 (N_8308,N_8223,N_8297);
and U8309 (N_8309,N_8270,N_8242);
xnor U8310 (N_8310,N_8221,N_8240);
nor U8311 (N_8311,N_8207,N_8299);
or U8312 (N_8312,N_8202,N_8283);
or U8313 (N_8313,N_8238,N_8285);
nand U8314 (N_8314,N_8250,N_8290);
or U8315 (N_8315,N_8235,N_8262);
nor U8316 (N_8316,N_8229,N_8215);
nor U8317 (N_8317,N_8253,N_8217);
xnor U8318 (N_8318,N_8210,N_8277);
or U8319 (N_8319,N_8296,N_8281);
nor U8320 (N_8320,N_8224,N_8214);
or U8321 (N_8321,N_8222,N_8276);
xnor U8322 (N_8322,N_8228,N_8244);
or U8323 (N_8323,N_8218,N_8231);
and U8324 (N_8324,N_8241,N_8298);
and U8325 (N_8325,N_8227,N_8200);
and U8326 (N_8326,N_8284,N_8208);
and U8327 (N_8327,N_8212,N_8275);
and U8328 (N_8328,N_8272,N_8259);
or U8329 (N_8329,N_8258,N_8282);
nand U8330 (N_8330,N_8274,N_8249);
and U8331 (N_8331,N_8216,N_8247);
or U8332 (N_8332,N_8251,N_8293);
nor U8333 (N_8333,N_8263,N_8232);
or U8334 (N_8334,N_8291,N_8287);
or U8335 (N_8335,N_8265,N_8237);
nand U8336 (N_8336,N_8248,N_8294);
nor U8337 (N_8337,N_8225,N_8255);
xor U8338 (N_8338,N_8268,N_8233);
and U8339 (N_8339,N_8205,N_8292);
nor U8340 (N_8340,N_8201,N_8273);
and U8341 (N_8341,N_8206,N_8226);
or U8342 (N_8342,N_8236,N_8203);
or U8343 (N_8343,N_8256,N_8243);
or U8344 (N_8344,N_8280,N_8278);
xor U8345 (N_8345,N_8245,N_8267);
nor U8346 (N_8346,N_8246,N_8269);
and U8347 (N_8347,N_8279,N_8254);
nor U8348 (N_8348,N_8213,N_8234);
or U8349 (N_8349,N_8260,N_8239);
or U8350 (N_8350,N_8208,N_8261);
and U8351 (N_8351,N_8244,N_8298);
xnor U8352 (N_8352,N_8292,N_8219);
nand U8353 (N_8353,N_8256,N_8269);
xor U8354 (N_8354,N_8266,N_8286);
and U8355 (N_8355,N_8294,N_8257);
and U8356 (N_8356,N_8265,N_8200);
or U8357 (N_8357,N_8228,N_8282);
nand U8358 (N_8358,N_8260,N_8227);
nand U8359 (N_8359,N_8207,N_8290);
and U8360 (N_8360,N_8275,N_8255);
nand U8361 (N_8361,N_8266,N_8210);
xor U8362 (N_8362,N_8242,N_8279);
nand U8363 (N_8363,N_8297,N_8253);
and U8364 (N_8364,N_8232,N_8288);
or U8365 (N_8365,N_8240,N_8212);
nand U8366 (N_8366,N_8216,N_8204);
nor U8367 (N_8367,N_8209,N_8201);
and U8368 (N_8368,N_8281,N_8265);
nand U8369 (N_8369,N_8256,N_8226);
and U8370 (N_8370,N_8247,N_8211);
nor U8371 (N_8371,N_8292,N_8248);
and U8372 (N_8372,N_8210,N_8242);
or U8373 (N_8373,N_8239,N_8277);
or U8374 (N_8374,N_8230,N_8278);
nand U8375 (N_8375,N_8269,N_8234);
xor U8376 (N_8376,N_8293,N_8244);
xor U8377 (N_8377,N_8264,N_8280);
nand U8378 (N_8378,N_8298,N_8254);
nand U8379 (N_8379,N_8253,N_8227);
and U8380 (N_8380,N_8200,N_8276);
nor U8381 (N_8381,N_8246,N_8284);
nor U8382 (N_8382,N_8254,N_8292);
nor U8383 (N_8383,N_8215,N_8218);
xor U8384 (N_8384,N_8291,N_8259);
nand U8385 (N_8385,N_8219,N_8252);
or U8386 (N_8386,N_8284,N_8288);
nor U8387 (N_8387,N_8287,N_8202);
or U8388 (N_8388,N_8264,N_8235);
or U8389 (N_8389,N_8269,N_8293);
nor U8390 (N_8390,N_8282,N_8232);
nor U8391 (N_8391,N_8223,N_8205);
or U8392 (N_8392,N_8233,N_8282);
or U8393 (N_8393,N_8254,N_8257);
and U8394 (N_8394,N_8238,N_8261);
nand U8395 (N_8395,N_8248,N_8275);
nand U8396 (N_8396,N_8213,N_8252);
and U8397 (N_8397,N_8273,N_8232);
nor U8398 (N_8398,N_8268,N_8222);
nand U8399 (N_8399,N_8230,N_8214);
and U8400 (N_8400,N_8328,N_8354);
nor U8401 (N_8401,N_8350,N_8338);
or U8402 (N_8402,N_8313,N_8331);
or U8403 (N_8403,N_8321,N_8366);
nor U8404 (N_8404,N_8320,N_8317);
nand U8405 (N_8405,N_8335,N_8364);
and U8406 (N_8406,N_8310,N_8303);
nand U8407 (N_8407,N_8373,N_8399);
or U8408 (N_8408,N_8300,N_8325);
nor U8409 (N_8409,N_8304,N_8347);
or U8410 (N_8410,N_8371,N_8352);
nor U8411 (N_8411,N_8375,N_8311);
nor U8412 (N_8412,N_8360,N_8365);
or U8413 (N_8413,N_8339,N_8356);
nor U8414 (N_8414,N_8305,N_8374);
and U8415 (N_8415,N_8397,N_8315);
xor U8416 (N_8416,N_8342,N_8308);
nand U8417 (N_8417,N_8353,N_8378);
nand U8418 (N_8418,N_8392,N_8359);
nand U8419 (N_8419,N_8391,N_8377);
nor U8420 (N_8420,N_8396,N_8324);
and U8421 (N_8421,N_8367,N_8312);
nand U8422 (N_8422,N_8340,N_8319);
nand U8423 (N_8423,N_8330,N_8314);
nor U8424 (N_8424,N_8388,N_8393);
nor U8425 (N_8425,N_8384,N_8345);
nor U8426 (N_8426,N_8334,N_8357);
or U8427 (N_8427,N_8346,N_8398);
and U8428 (N_8428,N_8362,N_8327);
and U8429 (N_8429,N_8368,N_8376);
xor U8430 (N_8430,N_8361,N_8329);
nand U8431 (N_8431,N_8323,N_8386);
nor U8432 (N_8432,N_8316,N_8318);
nor U8433 (N_8433,N_8383,N_8336);
and U8434 (N_8434,N_8379,N_8332);
or U8435 (N_8435,N_8326,N_8348);
nand U8436 (N_8436,N_8382,N_8341);
nor U8437 (N_8437,N_8381,N_8306);
and U8438 (N_8438,N_8349,N_8387);
or U8439 (N_8439,N_8351,N_8343);
or U8440 (N_8440,N_8370,N_8302);
or U8441 (N_8441,N_8337,N_8389);
nand U8442 (N_8442,N_8385,N_8358);
or U8443 (N_8443,N_8380,N_8355);
or U8444 (N_8444,N_8309,N_8390);
xnor U8445 (N_8445,N_8363,N_8333);
nor U8446 (N_8446,N_8344,N_8395);
or U8447 (N_8447,N_8322,N_8394);
and U8448 (N_8448,N_8301,N_8372);
nand U8449 (N_8449,N_8369,N_8307);
or U8450 (N_8450,N_8368,N_8362);
or U8451 (N_8451,N_8300,N_8328);
xor U8452 (N_8452,N_8392,N_8346);
nor U8453 (N_8453,N_8328,N_8380);
nand U8454 (N_8454,N_8395,N_8368);
or U8455 (N_8455,N_8330,N_8367);
nor U8456 (N_8456,N_8353,N_8361);
and U8457 (N_8457,N_8354,N_8357);
and U8458 (N_8458,N_8385,N_8329);
nor U8459 (N_8459,N_8349,N_8348);
xnor U8460 (N_8460,N_8360,N_8364);
nor U8461 (N_8461,N_8368,N_8361);
nor U8462 (N_8462,N_8389,N_8399);
and U8463 (N_8463,N_8323,N_8343);
nand U8464 (N_8464,N_8341,N_8363);
xor U8465 (N_8465,N_8376,N_8323);
nor U8466 (N_8466,N_8312,N_8364);
nand U8467 (N_8467,N_8359,N_8361);
and U8468 (N_8468,N_8317,N_8308);
xor U8469 (N_8469,N_8343,N_8370);
nand U8470 (N_8470,N_8320,N_8316);
nand U8471 (N_8471,N_8375,N_8368);
or U8472 (N_8472,N_8346,N_8333);
nand U8473 (N_8473,N_8309,N_8364);
and U8474 (N_8474,N_8339,N_8374);
or U8475 (N_8475,N_8354,N_8378);
nor U8476 (N_8476,N_8302,N_8331);
or U8477 (N_8477,N_8384,N_8321);
or U8478 (N_8478,N_8335,N_8333);
or U8479 (N_8479,N_8339,N_8306);
or U8480 (N_8480,N_8394,N_8331);
nand U8481 (N_8481,N_8378,N_8345);
nor U8482 (N_8482,N_8330,N_8301);
or U8483 (N_8483,N_8357,N_8384);
and U8484 (N_8484,N_8340,N_8339);
xnor U8485 (N_8485,N_8301,N_8346);
and U8486 (N_8486,N_8388,N_8357);
nor U8487 (N_8487,N_8311,N_8359);
nand U8488 (N_8488,N_8353,N_8334);
or U8489 (N_8489,N_8311,N_8383);
nand U8490 (N_8490,N_8311,N_8313);
or U8491 (N_8491,N_8301,N_8356);
nand U8492 (N_8492,N_8328,N_8306);
nor U8493 (N_8493,N_8316,N_8356);
or U8494 (N_8494,N_8331,N_8382);
and U8495 (N_8495,N_8364,N_8350);
and U8496 (N_8496,N_8393,N_8331);
nand U8497 (N_8497,N_8303,N_8390);
and U8498 (N_8498,N_8346,N_8309);
or U8499 (N_8499,N_8359,N_8308);
nor U8500 (N_8500,N_8441,N_8407);
nor U8501 (N_8501,N_8425,N_8465);
or U8502 (N_8502,N_8486,N_8433);
nand U8503 (N_8503,N_8489,N_8482);
nor U8504 (N_8504,N_8475,N_8402);
or U8505 (N_8505,N_8472,N_8413);
and U8506 (N_8506,N_8462,N_8435);
nor U8507 (N_8507,N_8458,N_8491);
or U8508 (N_8508,N_8446,N_8403);
nor U8509 (N_8509,N_8490,N_8427);
nand U8510 (N_8510,N_8404,N_8459);
xor U8511 (N_8511,N_8400,N_8426);
and U8512 (N_8512,N_8422,N_8498);
nand U8513 (N_8513,N_8438,N_8453);
or U8514 (N_8514,N_8409,N_8431);
or U8515 (N_8515,N_8421,N_8449);
or U8516 (N_8516,N_8473,N_8414);
xor U8517 (N_8517,N_8424,N_8460);
nor U8518 (N_8518,N_8432,N_8437);
and U8519 (N_8519,N_8463,N_8452);
or U8520 (N_8520,N_8405,N_8470);
and U8521 (N_8521,N_8496,N_8484);
or U8522 (N_8522,N_8478,N_8485);
nand U8523 (N_8523,N_8466,N_8456);
and U8524 (N_8524,N_8418,N_8447);
nor U8525 (N_8525,N_8467,N_8443);
nand U8526 (N_8526,N_8428,N_8434);
nand U8527 (N_8527,N_8445,N_8448);
or U8528 (N_8528,N_8483,N_8479);
nor U8529 (N_8529,N_8487,N_8492);
xnor U8530 (N_8530,N_8451,N_8440);
nor U8531 (N_8531,N_8429,N_8450);
or U8532 (N_8532,N_8406,N_8455);
nand U8533 (N_8533,N_8444,N_8442);
and U8534 (N_8534,N_8476,N_8439);
xor U8535 (N_8535,N_8497,N_8493);
and U8536 (N_8536,N_8420,N_8430);
or U8537 (N_8537,N_8464,N_8477);
and U8538 (N_8538,N_8474,N_8469);
xnor U8539 (N_8539,N_8454,N_8457);
or U8540 (N_8540,N_8494,N_8408);
xor U8541 (N_8541,N_8415,N_8412);
nand U8542 (N_8542,N_8481,N_8471);
and U8543 (N_8543,N_8436,N_8480);
or U8544 (N_8544,N_8495,N_8461);
or U8545 (N_8545,N_8423,N_8410);
and U8546 (N_8546,N_8468,N_8401);
nand U8547 (N_8547,N_8499,N_8419);
nor U8548 (N_8548,N_8411,N_8488);
and U8549 (N_8549,N_8416,N_8417);
nand U8550 (N_8550,N_8447,N_8483);
or U8551 (N_8551,N_8441,N_8465);
nand U8552 (N_8552,N_8422,N_8449);
nor U8553 (N_8553,N_8496,N_8478);
and U8554 (N_8554,N_8446,N_8450);
nand U8555 (N_8555,N_8481,N_8409);
nor U8556 (N_8556,N_8454,N_8442);
and U8557 (N_8557,N_8400,N_8440);
and U8558 (N_8558,N_8420,N_8431);
nor U8559 (N_8559,N_8427,N_8412);
nor U8560 (N_8560,N_8445,N_8479);
and U8561 (N_8561,N_8431,N_8460);
nor U8562 (N_8562,N_8478,N_8495);
or U8563 (N_8563,N_8472,N_8461);
and U8564 (N_8564,N_8465,N_8405);
or U8565 (N_8565,N_8425,N_8478);
or U8566 (N_8566,N_8444,N_8465);
or U8567 (N_8567,N_8487,N_8482);
nand U8568 (N_8568,N_8451,N_8400);
xor U8569 (N_8569,N_8479,N_8448);
xnor U8570 (N_8570,N_8484,N_8400);
or U8571 (N_8571,N_8490,N_8471);
xnor U8572 (N_8572,N_8415,N_8406);
nand U8573 (N_8573,N_8403,N_8469);
or U8574 (N_8574,N_8495,N_8407);
and U8575 (N_8575,N_8403,N_8454);
xor U8576 (N_8576,N_8428,N_8415);
and U8577 (N_8577,N_8463,N_8409);
xnor U8578 (N_8578,N_8434,N_8443);
or U8579 (N_8579,N_8456,N_8433);
nand U8580 (N_8580,N_8472,N_8444);
nand U8581 (N_8581,N_8478,N_8418);
nor U8582 (N_8582,N_8420,N_8458);
nor U8583 (N_8583,N_8468,N_8425);
xor U8584 (N_8584,N_8419,N_8496);
and U8585 (N_8585,N_8484,N_8421);
and U8586 (N_8586,N_8433,N_8408);
or U8587 (N_8587,N_8456,N_8406);
and U8588 (N_8588,N_8496,N_8413);
and U8589 (N_8589,N_8467,N_8439);
nand U8590 (N_8590,N_8477,N_8482);
xnor U8591 (N_8591,N_8407,N_8474);
and U8592 (N_8592,N_8443,N_8473);
and U8593 (N_8593,N_8462,N_8403);
xor U8594 (N_8594,N_8467,N_8402);
or U8595 (N_8595,N_8479,N_8449);
or U8596 (N_8596,N_8408,N_8479);
or U8597 (N_8597,N_8471,N_8435);
and U8598 (N_8598,N_8467,N_8450);
nor U8599 (N_8599,N_8403,N_8476);
nor U8600 (N_8600,N_8583,N_8535);
nand U8601 (N_8601,N_8529,N_8541);
nor U8602 (N_8602,N_8558,N_8544);
and U8603 (N_8603,N_8500,N_8520);
nor U8604 (N_8604,N_8561,N_8568);
nor U8605 (N_8605,N_8540,N_8590);
or U8606 (N_8606,N_8508,N_8557);
nand U8607 (N_8607,N_8543,N_8512);
nor U8608 (N_8608,N_8591,N_8570);
nor U8609 (N_8609,N_8507,N_8553);
nand U8610 (N_8610,N_8572,N_8552);
and U8611 (N_8611,N_8514,N_8503);
or U8612 (N_8612,N_8587,N_8515);
nor U8613 (N_8613,N_8519,N_8582);
nor U8614 (N_8614,N_8509,N_8564);
nand U8615 (N_8615,N_8589,N_8581);
nor U8616 (N_8616,N_8598,N_8545);
and U8617 (N_8617,N_8530,N_8586);
or U8618 (N_8618,N_8521,N_8518);
nand U8619 (N_8619,N_8556,N_8516);
nand U8620 (N_8620,N_8562,N_8560);
nand U8621 (N_8621,N_8592,N_8538);
and U8622 (N_8622,N_8549,N_8580);
and U8623 (N_8623,N_8511,N_8547);
xnor U8624 (N_8624,N_8506,N_8517);
or U8625 (N_8625,N_8523,N_8597);
nand U8626 (N_8626,N_8536,N_8588);
nor U8627 (N_8627,N_8528,N_8524);
xnor U8628 (N_8628,N_8584,N_8525);
nor U8629 (N_8629,N_8596,N_8579);
nand U8630 (N_8630,N_8571,N_8526);
or U8631 (N_8631,N_8563,N_8504);
or U8632 (N_8632,N_8559,N_8565);
and U8633 (N_8633,N_8578,N_8585);
or U8634 (N_8634,N_8546,N_8542);
nand U8635 (N_8635,N_8505,N_8522);
nor U8636 (N_8636,N_8532,N_8510);
and U8637 (N_8637,N_8575,N_8502);
nand U8638 (N_8638,N_8599,N_8574);
xor U8639 (N_8639,N_8548,N_8573);
or U8640 (N_8640,N_8554,N_8527);
nor U8641 (N_8641,N_8567,N_8550);
or U8642 (N_8642,N_8569,N_8513);
nand U8643 (N_8643,N_8537,N_8534);
or U8644 (N_8644,N_8501,N_8595);
xnor U8645 (N_8645,N_8551,N_8539);
and U8646 (N_8646,N_8593,N_8566);
nor U8647 (N_8647,N_8555,N_8577);
nand U8648 (N_8648,N_8533,N_8576);
xor U8649 (N_8649,N_8594,N_8531);
and U8650 (N_8650,N_8502,N_8565);
nor U8651 (N_8651,N_8585,N_8529);
nand U8652 (N_8652,N_8531,N_8540);
nand U8653 (N_8653,N_8530,N_8585);
or U8654 (N_8654,N_8586,N_8511);
or U8655 (N_8655,N_8501,N_8567);
nand U8656 (N_8656,N_8583,N_8502);
nand U8657 (N_8657,N_8567,N_8510);
and U8658 (N_8658,N_8559,N_8573);
or U8659 (N_8659,N_8507,N_8513);
nor U8660 (N_8660,N_8592,N_8543);
or U8661 (N_8661,N_8573,N_8519);
or U8662 (N_8662,N_8558,N_8562);
and U8663 (N_8663,N_8504,N_8549);
or U8664 (N_8664,N_8593,N_8540);
and U8665 (N_8665,N_8569,N_8582);
xnor U8666 (N_8666,N_8504,N_8519);
or U8667 (N_8667,N_8574,N_8568);
and U8668 (N_8668,N_8516,N_8563);
or U8669 (N_8669,N_8589,N_8504);
xnor U8670 (N_8670,N_8522,N_8541);
nor U8671 (N_8671,N_8563,N_8501);
and U8672 (N_8672,N_8597,N_8542);
xor U8673 (N_8673,N_8555,N_8507);
and U8674 (N_8674,N_8570,N_8521);
xnor U8675 (N_8675,N_8533,N_8592);
nor U8676 (N_8676,N_8522,N_8577);
nand U8677 (N_8677,N_8556,N_8527);
nand U8678 (N_8678,N_8547,N_8516);
nand U8679 (N_8679,N_8585,N_8575);
or U8680 (N_8680,N_8545,N_8593);
or U8681 (N_8681,N_8506,N_8590);
and U8682 (N_8682,N_8539,N_8540);
nand U8683 (N_8683,N_8505,N_8576);
nor U8684 (N_8684,N_8546,N_8554);
nor U8685 (N_8685,N_8527,N_8565);
and U8686 (N_8686,N_8566,N_8561);
nand U8687 (N_8687,N_8552,N_8558);
nand U8688 (N_8688,N_8576,N_8563);
nor U8689 (N_8689,N_8578,N_8598);
and U8690 (N_8690,N_8549,N_8543);
or U8691 (N_8691,N_8583,N_8599);
nor U8692 (N_8692,N_8556,N_8599);
or U8693 (N_8693,N_8596,N_8541);
or U8694 (N_8694,N_8536,N_8508);
and U8695 (N_8695,N_8528,N_8578);
nor U8696 (N_8696,N_8532,N_8549);
and U8697 (N_8697,N_8545,N_8564);
nand U8698 (N_8698,N_8550,N_8511);
nor U8699 (N_8699,N_8546,N_8535);
xnor U8700 (N_8700,N_8656,N_8612);
or U8701 (N_8701,N_8676,N_8652);
nand U8702 (N_8702,N_8680,N_8677);
nand U8703 (N_8703,N_8674,N_8681);
or U8704 (N_8704,N_8602,N_8617);
and U8705 (N_8705,N_8630,N_8641);
nor U8706 (N_8706,N_8622,N_8627);
nor U8707 (N_8707,N_8606,N_8692);
or U8708 (N_8708,N_8649,N_8693);
or U8709 (N_8709,N_8666,N_8631);
and U8710 (N_8710,N_8644,N_8615);
and U8711 (N_8711,N_8699,N_8614);
nor U8712 (N_8712,N_8646,N_8663);
or U8713 (N_8713,N_8648,N_8690);
nor U8714 (N_8714,N_8611,N_8657);
nor U8715 (N_8715,N_8691,N_8618);
nand U8716 (N_8716,N_8673,N_8620);
nor U8717 (N_8717,N_8636,N_8642);
xnor U8718 (N_8718,N_8623,N_8682);
or U8719 (N_8719,N_8601,N_8607);
and U8720 (N_8720,N_8668,N_8616);
and U8721 (N_8721,N_8610,N_8665);
and U8722 (N_8722,N_8619,N_8686);
and U8723 (N_8723,N_8629,N_8667);
nand U8724 (N_8724,N_8679,N_8655);
nor U8725 (N_8725,N_8639,N_8637);
nand U8726 (N_8726,N_8695,N_8604);
nand U8727 (N_8727,N_8633,N_8647);
or U8728 (N_8728,N_8628,N_8659);
or U8729 (N_8729,N_8638,N_8624);
nor U8730 (N_8730,N_8605,N_8609);
and U8731 (N_8731,N_8650,N_8689);
or U8732 (N_8732,N_8600,N_8603);
nor U8733 (N_8733,N_8696,N_8621);
and U8734 (N_8734,N_8653,N_8669);
nor U8735 (N_8735,N_8640,N_8664);
and U8736 (N_8736,N_8654,N_8688);
nand U8737 (N_8737,N_8698,N_8672);
and U8738 (N_8738,N_8684,N_8651);
xnor U8739 (N_8739,N_8675,N_8626);
nor U8740 (N_8740,N_8661,N_8635);
or U8741 (N_8741,N_8643,N_8685);
xor U8742 (N_8742,N_8660,N_8662);
and U8743 (N_8743,N_8678,N_8683);
xnor U8744 (N_8744,N_8625,N_8634);
and U8745 (N_8745,N_8687,N_8632);
nand U8746 (N_8746,N_8671,N_8608);
or U8747 (N_8747,N_8670,N_8694);
nand U8748 (N_8748,N_8645,N_8697);
nor U8749 (N_8749,N_8658,N_8613);
or U8750 (N_8750,N_8687,N_8673);
nor U8751 (N_8751,N_8651,N_8669);
xnor U8752 (N_8752,N_8684,N_8658);
or U8753 (N_8753,N_8669,N_8622);
xor U8754 (N_8754,N_8694,N_8612);
nand U8755 (N_8755,N_8640,N_8650);
or U8756 (N_8756,N_8604,N_8608);
or U8757 (N_8757,N_8684,N_8637);
nand U8758 (N_8758,N_8612,N_8642);
nand U8759 (N_8759,N_8608,N_8651);
nand U8760 (N_8760,N_8650,N_8692);
and U8761 (N_8761,N_8676,N_8677);
nor U8762 (N_8762,N_8602,N_8656);
or U8763 (N_8763,N_8659,N_8644);
nand U8764 (N_8764,N_8608,N_8642);
and U8765 (N_8765,N_8671,N_8685);
or U8766 (N_8766,N_8695,N_8617);
xnor U8767 (N_8767,N_8663,N_8667);
xor U8768 (N_8768,N_8618,N_8608);
xor U8769 (N_8769,N_8639,N_8658);
and U8770 (N_8770,N_8650,N_8609);
and U8771 (N_8771,N_8677,N_8639);
xor U8772 (N_8772,N_8600,N_8694);
nand U8773 (N_8773,N_8651,N_8672);
nor U8774 (N_8774,N_8674,N_8630);
nor U8775 (N_8775,N_8654,N_8689);
or U8776 (N_8776,N_8693,N_8679);
nand U8777 (N_8777,N_8615,N_8611);
nand U8778 (N_8778,N_8644,N_8654);
nand U8779 (N_8779,N_8686,N_8661);
nor U8780 (N_8780,N_8679,N_8622);
or U8781 (N_8781,N_8697,N_8626);
nor U8782 (N_8782,N_8667,N_8631);
nor U8783 (N_8783,N_8664,N_8684);
nor U8784 (N_8784,N_8661,N_8688);
and U8785 (N_8785,N_8626,N_8663);
nand U8786 (N_8786,N_8634,N_8678);
nor U8787 (N_8787,N_8641,N_8607);
and U8788 (N_8788,N_8686,N_8683);
xor U8789 (N_8789,N_8632,N_8626);
or U8790 (N_8790,N_8654,N_8685);
or U8791 (N_8791,N_8626,N_8617);
xor U8792 (N_8792,N_8676,N_8606);
nor U8793 (N_8793,N_8603,N_8616);
nand U8794 (N_8794,N_8630,N_8620);
and U8795 (N_8795,N_8679,N_8669);
and U8796 (N_8796,N_8614,N_8654);
or U8797 (N_8797,N_8648,N_8615);
nor U8798 (N_8798,N_8626,N_8652);
nor U8799 (N_8799,N_8676,N_8649);
or U8800 (N_8800,N_8779,N_8761);
nor U8801 (N_8801,N_8771,N_8716);
or U8802 (N_8802,N_8750,N_8702);
nand U8803 (N_8803,N_8714,N_8703);
nand U8804 (N_8804,N_8722,N_8740);
xnor U8805 (N_8805,N_8757,N_8741);
or U8806 (N_8806,N_8799,N_8751);
or U8807 (N_8807,N_8798,N_8735);
or U8808 (N_8808,N_8775,N_8758);
nand U8809 (N_8809,N_8795,N_8712);
nor U8810 (N_8810,N_8724,N_8759);
and U8811 (N_8811,N_8743,N_8753);
nand U8812 (N_8812,N_8774,N_8768);
and U8813 (N_8813,N_8762,N_8739);
and U8814 (N_8814,N_8785,N_8731);
nand U8815 (N_8815,N_8730,N_8780);
and U8816 (N_8816,N_8752,N_8770);
xnor U8817 (N_8817,N_8700,N_8786);
nand U8818 (N_8818,N_8733,N_8710);
nand U8819 (N_8819,N_8718,N_8755);
or U8820 (N_8820,N_8732,N_8749);
nor U8821 (N_8821,N_8707,N_8742);
nand U8822 (N_8822,N_8734,N_8704);
and U8823 (N_8823,N_8717,N_8769);
nor U8824 (N_8824,N_8788,N_8723);
nand U8825 (N_8825,N_8747,N_8789);
nand U8826 (N_8826,N_8781,N_8721);
nand U8827 (N_8827,N_8778,N_8760);
and U8828 (N_8828,N_8766,N_8772);
xor U8829 (N_8829,N_8792,N_8797);
or U8830 (N_8830,N_8782,N_8745);
nor U8831 (N_8831,N_8736,N_8738);
or U8832 (N_8832,N_8713,N_8725);
and U8833 (N_8833,N_8727,N_8705);
or U8834 (N_8834,N_8708,N_8754);
nor U8835 (N_8835,N_8701,N_8787);
and U8836 (N_8836,N_8726,N_8784);
nor U8837 (N_8837,N_8783,N_8711);
and U8838 (N_8838,N_8709,N_8790);
and U8839 (N_8839,N_8729,N_8756);
and U8840 (N_8840,N_8744,N_8794);
or U8841 (N_8841,N_8777,N_8728);
nor U8842 (N_8842,N_8793,N_8706);
or U8843 (N_8843,N_8796,N_8776);
or U8844 (N_8844,N_8765,N_8748);
or U8845 (N_8845,N_8715,N_8719);
nor U8846 (N_8846,N_8720,N_8791);
nor U8847 (N_8847,N_8737,N_8763);
nor U8848 (N_8848,N_8746,N_8773);
nand U8849 (N_8849,N_8767,N_8764);
xor U8850 (N_8850,N_8720,N_8795);
nor U8851 (N_8851,N_8732,N_8783);
or U8852 (N_8852,N_8754,N_8751);
or U8853 (N_8853,N_8761,N_8778);
xnor U8854 (N_8854,N_8705,N_8774);
and U8855 (N_8855,N_8702,N_8754);
nand U8856 (N_8856,N_8754,N_8759);
or U8857 (N_8857,N_8773,N_8713);
nand U8858 (N_8858,N_8700,N_8730);
nand U8859 (N_8859,N_8785,N_8737);
xor U8860 (N_8860,N_8779,N_8724);
nor U8861 (N_8861,N_8791,N_8727);
and U8862 (N_8862,N_8722,N_8728);
nand U8863 (N_8863,N_8760,N_8797);
or U8864 (N_8864,N_8701,N_8767);
nand U8865 (N_8865,N_8711,N_8760);
xor U8866 (N_8866,N_8783,N_8702);
or U8867 (N_8867,N_8744,N_8723);
xnor U8868 (N_8868,N_8756,N_8767);
nand U8869 (N_8869,N_8742,N_8712);
xor U8870 (N_8870,N_8739,N_8744);
xor U8871 (N_8871,N_8712,N_8784);
and U8872 (N_8872,N_8795,N_8767);
and U8873 (N_8873,N_8752,N_8722);
xnor U8874 (N_8874,N_8726,N_8728);
or U8875 (N_8875,N_8784,N_8749);
or U8876 (N_8876,N_8715,N_8720);
nor U8877 (N_8877,N_8730,N_8704);
and U8878 (N_8878,N_8797,N_8734);
nor U8879 (N_8879,N_8721,N_8738);
nand U8880 (N_8880,N_8753,N_8725);
nor U8881 (N_8881,N_8784,N_8783);
and U8882 (N_8882,N_8703,N_8754);
nand U8883 (N_8883,N_8753,N_8755);
or U8884 (N_8884,N_8786,N_8736);
or U8885 (N_8885,N_8777,N_8796);
nand U8886 (N_8886,N_8754,N_8764);
or U8887 (N_8887,N_8752,N_8783);
nor U8888 (N_8888,N_8733,N_8742);
or U8889 (N_8889,N_8776,N_8766);
nor U8890 (N_8890,N_8793,N_8787);
nor U8891 (N_8891,N_8775,N_8764);
nand U8892 (N_8892,N_8796,N_8743);
or U8893 (N_8893,N_8721,N_8740);
and U8894 (N_8894,N_8773,N_8730);
nand U8895 (N_8895,N_8790,N_8798);
nor U8896 (N_8896,N_8759,N_8743);
nand U8897 (N_8897,N_8725,N_8701);
and U8898 (N_8898,N_8782,N_8792);
nand U8899 (N_8899,N_8703,N_8701);
nor U8900 (N_8900,N_8860,N_8816);
and U8901 (N_8901,N_8854,N_8813);
nor U8902 (N_8902,N_8871,N_8822);
xor U8903 (N_8903,N_8817,N_8885);
and U8904 (N_8904,N_8857,N_8892);
nor U8905 (N_8905,N_8888,N_8838);
and U8906 (N_8906,N_8826,N_8837);
xor U8907 (N_8907,N_8839,N_8821);
and U8908 (N_8908,N_8848,N_8835);
and U8909 (N_8909,N_8894,N_8846);
and U8910 (N_8910,N_8895,N_8870);
and U8911 (N_8911,N_8829,N_8882);
or U8912 (N_8912,N_8884,N_8898);
nand U8913 (N_8913,N_8862,N_8859);
or U8914 (N_8914,N_8867,N_8881);
nor U8915 (N_8915,N_8861,N_8863);
and U8916 (N_8916,N_8880,N_8856);
nor U8917 (N_8917,N_8858,N_8875);
xor U8918 (N_8918,N_8810,N_8823);
nand U8919 (N_8919,N_8844,N_8847);
and U8920 (N_8920,N_8864,N_8872);
nor U8921 (N_8921,N_8819,N_8874);
nor U8922 (N_8922,N_8831,N_8834);
xnor U8923 (N_8923,N_8840,N_8805);
nand U8924 (N_8924,N_8889,N_8824);
and U8925 (N_8925,N_8841,N_8836);
xor U8926 (N_8926,N_8877,N_8845);
or U8927 (N_8927,N_8825,N_8808);
or U8928 (N_8928,N_8827,N_8899);
and U8929 (N_8929,N_8806,N_8801);
nand U8930 (N_8930,N_8866,N_8830);
xor U8931 (N_8931,N_8893,N_8832);
nor U8932 (N_8932,N_8812,N_8833);
nor U8933 (N_8933,N_8809,N_8883);
xnor U8934 (N_8934,N_8887,N_8891);
or U8935 (N_8935,N_8815,N_8868);
nand U8936 (N_8936,N_8849,N_8814);
or U8937 (N_8937,N_8842,N_8855);
nand U8938 (N_8938,N_8802,N_8803);
nand U8939 (N_8939,N_8853,N_8890);
or U8940 (N_8940,N_8804,N_8878);
nor U8941 (N_8941,N_8865,N_8873);
xor U8942 (N_8942,N_8896,N_8807);
xnor U8943 (N_8943,N_8828,N_8800);
nor U8944 (N_8944,N_8852,N_8818);
nand U8945 (N_8945,N_8843,N_8897);
nor U8946 (N_8946,N_8820,N_8811);
nor U8947 (N_8947,N_8886,N_8876);
nor U8948 (N_8948,N_8879,N_8850);
and U8949 (N_8949,N_8851,N_8869);
and U8950 (N_8950,N_8845,N_8885);
nor U8951 (N_8951,N_8807,N_8878);
nor U8952 (N_8952,N_8840,N_8882);
or U8953 (N_8953,N_8880,N_8812);
or U8954 (N_8954,N_8879,N_8865);
and U8955 (N_8955,N_8890,N_8815);
xor U8956 (N_8956,N_8898,N_8827);
nor U8957 (N_8957,N_8843,N_8888);
or U8958 (N_8958,N_8891,N_8839);
xor U8959 (N_8959,N_8836,N_8884);
xnor U8960 (N_8960,N_8893,N_8813);
xnor U8961 (N_8961,N_8861,N_8872);
nand U8962 (N_8962,N_8813,N_8886);
or U8963 (N_8963,N_8862,N_8888);
and U8964 (N_8964,N_8819,N_8861);
nor U8965 (N_8965,N_8838,N_8881);
xor U8966 (N_8966,N_8820,N_8877);
or U8967 (N_8967,N_8828,N_8823);
and U8968 (N_8968,N_8849,N_8886);
xnor U8969 (N_8969,N_8855,N_8809);
nor U8970 (N_8970,N_8857,N_8865);
nand U8971 (N_8971,N_8808,N_8822);
and U8972 (N_8972,N_8828,N_8895);
and U8973 (N_8973,N_8889,N_8894);
nand U8974 (N_8974,N_8864,N_8811);
or U8975 (N_8975,N_8859,N_8825);
nor U8976 (N_8976,N_8838,N_8811);
nor U8977 (N_8977,N_8835,N_8885);
nand U8978 (N_8978,N_8847,N_8882);
and U8979 (N_8979,N_8848,N_8814);
nor U8980 (N_8980,N_8873,N_8875);
or U8981 (N_8981,N_8884,N_8813);
nor U8982 (N_8982,N_8873,N_8822);
nand U8983 (N_8983,N_8874,N_8873);
nor U8984 (N_8984,N_8865,N_8825);
xor U8985 (N_8985,N_8849,N_8810);
or U8986 (N_8986,N_8813,N_8835);
or U8987 (N_8987,N_8851,N_8854);
and U8988 (N_8988,N_8834,N_8828);
nand U8989 (N_8989,N_8895,N_8820);
and U8990 (N_8990,N_8820,N_8851);
nand U8991 (N_8991,N_8849,N_8853);
nand U8992 (N_8992,N_8886,N_8892);
nor U8993 (N_8993,N_8891,N_8826);
or U8994 (N_8994,N_8879,N_8813);
and U8995 (N_8995,N_8842,N_8866);
nor U8996 (N_8996,N_8828,N_8866);
xor U8997 (N_8997,N_8847,N_8894);
xor U8998 (N_8998,N_8829,N_8889);
nor U8999 (N_8999,N_8839,N_8883);
xnor U9000 (N_9000,N_8992,N_8920);
nand U9001 (N_9001,N_8980,N_8949);
or U9002 (N_9002,N_8971,N_8914);
or U9003 (N_9003,N_8982,N_8944);
and U9004 (N_9004,N_8942,N_8931);
and U9005 (N_9005,N_8932,N_8943);
xnor U9006 (N_9006,N_8998,N_8917);
nor U9007 (N_9007,N_8977,N_8981);
or U9008 (N_9008,N_8908,N_8975);
nor U9009 (N_9009,N_8916,N_8902);
or U9010 (N_9010,N_8991,N_8987);
and U9011 (N_9011,N_8924,N_8933);
nand U9012 (N_9012,N_8994,N_8926);
or U9013 (N_9013,N_8940,N_8978);
nand U9014 (N_9014,N_8960,N_8997);
xor U9015 (N_9015,N_8906,N_8969);
nor U9016 (N_9016,N_8915,N_8937);
and U9017 (N_9017,N_8946,N_8905);
and U9018 (N_9018,N_8922,N_8907);
or U9019 (N_9019,N_8951,N_8972);
or U9020 (N_9020,N_8956,N_8930);
or U9021 (N_9021,N_8918,N_8970);
nor U9022 (N_9022,N_8963,N_8995);
and U9023 (N_9023,N_8983,N_8945);
nor U9024 (N_9024,N_8954,N_8959);
nand U9025 (N_9025,N_8996,N_8900);
and U9026 (N_9026,N_8929,N_8911);
and U9027 (N_9027,N_8938,N_8953);
nor U9028 (N_9028,N_8989,N_8979);
or U9029 (N_9029,N_8988,N_8990);
nor U9030 (N_9030,N_8984,N_8973);
nand U9031 (N_9031,N_8925,N_8965);
or U9032 (N_9032,N_8913,N_8928);
and U9033 (N_9033,N_8934,N_8903);
nor U9034 (N_9034,N_8993,N_8986);
nand U9035 (N_9035,N_8999,N_8909);
xnor U9036 (N_9036,N_8927,N_8901);
or U9037 (N_9037,N_8912,N_8958);
nor U9038 (N_9038,N_8957,N_8910);
xor U9039 (N_9039,N_8921,N_8936);
or U9040 (N_9040,N_8904,N_8950);
nor U9041 (N_9041,N_8947,N_8962);
xnor U9042 (N_9042,N_8939,N_8919);
nor U9043 (N_9043,N_8941,N_8964);
nor U9044 (N_9044,N_8976,N_8974);
or U9045 (N_9045,N_8985,N_8935);
nand U9046 (N_9046,N_8968,N_8967);
xnor U9047 (N_9047,N_8955,N_8948);
and U9048 (N_9048,N_8923,N_8966);
or U9049 (N_9049,N_8952,N_8961);
and U9050 (N_9050,N_8920,N_8973);
and U9051 (N_9051,N_8931,N_8981);
and U9052 (N_9052,N_8926,N_8930);
nand U9053 (N_9053,N_8999,N_8973);
or U9054 (N_9054,N_8924,N_8985);
and U9055 (N_9055,N_8902,N_8941);
nand U9056 (N_9056,N_8906,N_8991);
nor U9057 (N_9057,N_8978,N_8914);
nand U9058 (N_9058,N_8945,N_8969);
nor U9059 (N_9059,N_8970,N_8949);
nand U9060 (N_9060,N_8919,N_8977);
or U9061 (N_9061,N_8933,N_8987);
and U9062 (N_9062,N_8902,N_8992);
and U9063 (N_9063,N_8909,N_8967);
nor U9064 (N_9064,N_8945,N_8976);
nor U9065 (N_9065,N_8953,N_8972);
and U9066 (N_9066,N_8971,N_8909);
or U9067 (N_9067,N_8905,N_8959);
nand U9068 (N_9068,N_8964,N_8989);
or U9069 (N_9069,N_8970,N_8984);
or U9070 (N_9070,N_8963,N_8951);
xor U9071 (N_9071,N_8959,N_8949);
xnor U9072 (N_9072,N_8925,N_8932);
xor U9073 (N_9073,N_8960,N_8942);
nor U9074 (N_9074,N_8902,N_8950);
nor U9075 (N_9075,N_8978,N_8980);
nor U9076 (N_9076,N_8949,N_8939);
nand U9077 (N_9077,N_8982,N_8977);
and U9078 (N_9078,N_8942,N_8903);
and U9079 (N_9079,N_8952,N_8931);
or U9080 (N_9080,N_8956,N_8970);
and U9081 (N_9081,N_8964,N_8950);
and U9082 (N_9082,N_8966,N_8952);
or U9083 (N_9083,N_8920,N_8975);
xnor U9084 (N_9084,N_8916,N_8963);
nand U9085 (N_9085,N_8991,N_8936);
nor U9086 (N_9086,N_8925,N_8966);
nand U9087 (N_9087,N_8923,N_8916);
or U9088 (N_9088,N_8973,N_8955);
nand U9089 (N_9089,N_8963,N_8911);
or U9090 (N_9090,N_8996,N_8998);
nor U9091 (N_9091,N_8997,N_8966);
nor U9092 (N_9092,N_8979,N_8965);
nand U9093 (N_9093,N_8919,N_8941);
nand U9094 (N_9094,N_8934,N_8968);
and U9095 (N_9095,N_8937,N_8942);
and U9096 (N_9096,N_8965,N_8937);
nor U9097 (N_9097,N_8969,N_8981);
nand U9098 (N_9098,N_8922,N_8913);
and U9099 (N_9099,N_8929,N_8932);
nor U9100 (N_9100,N_9018,N_9011);
and U9101 (N_9101,N_9024,N_9089);
and U9102 (N_9102,N_9010,N_9060);
xnor U9103 (N_9103,N_9016,N_9071);
nand U9104 (N_9104,N_9004,N_9052);
nor U9105 (N_9105,N_9008,N_9015);
or U9106 (N_9106,N_9023,N_9003);
or U9107 (N_9107,N_9045,N_9055);
or U9108 (N_9108,N_9041,N_9050);
nor U9109 (N_9109,N_9049,N_9035);
nor U9110 (N_9110,N_9062,N_9005);
or U9111 (N_9111,N_9085,N_9088);
and U9112 (N_9112,N_9067,N_9036);
and U9113 (N_9113,N_9043,N_9019);
or U9114 (N_9114,N_9087,N_9044);
or U9115 (N_9115,N_9078,N_9031);
and U9116 (N_9116,N_9021,N_9007);
nand U9117 (N_9117,N_9000,N_9006);
or U9118 (N_9118,N_9068,N_9064);
xnor U9119 (N_9119,N_9001,N_9038);
nand U9120 (N_9120,N_9075,N_9027);
xnor U9121 (N_9121,N_9066,N_9028);
nand U9122 (N_9122,N_9095,N_9074);
or U9123 (N_9123,N_9020,N_9084);
and U9124 (N_9124,N_9090,N_9073);
or U9125 (N_9125,N_9042,N_9069);
or U9126 (N_9126,N_9091,N_9029);
nor U9127 (N_9127,N_9079,N_9034);
nor U9128 (N_9128,N_9092,N_9048);
nor U9129 (N_9129,N_9022,N_9081);
nor U9130 (N_9130,N_9080,N_9013);
and U9131 (N_9131,N_9026,N_9054);
nor U9132 (N_9132,N_9032,N_9025);
xor U9133 (N_9133,N_9059,N_9098);
nor U9134 (N_9134,N_9040,N_9061);
nor U9135 (N_9135,N_9002,N_9014);
and U9136 (N_9136,N_9070,N_9065);
and U9137 (N_9137,N_9009,N_9033);
nand U9138 (N_9138,N_9094,N_9097);
nand U9139 (N_9139,N_9099,N_9047);
nor U9140 (N_9140,N_9076,N_9057);
nand U9141 (N_9141,N_9093,N_9037);
nor U9142 (N_9142,N_9053,N_9030);
nor U9143 (N_9143,N_9096,N_9083);
or U9144 (N_9144,N_9082,N_9039);
xnor U9145 (N_9145,N_9058,N_9072);
and U9146 (N_9146,N_9012,N_9086);
and U9147 (N_9147,N_9051,N_9063);
nand U9148 (N_9148,N_9017,N_9046);
nand U9149 (N_9149,N_9077,N_9056);
or U9150 (N_9150,N_9017,N_9086);
nand U9151 (N_9151,N_9083,N_9093);
and U9152 (N_9152,N_9018,N_9070);
nor U9153 (N_9153,N_9071,N_9073);
nand U9154 (N_9154,N_9074,N_9040);
xor U9155 (N_9155,N_9062,N_9047);
nor U9156 (N_9156,N_9077,N_9036);
nor U9157 (N_9157,N_9015,N_9092);
nand U9158 (N_9158,N_9079,N_9001);
or U9159 (N_9159,N_9001,N_9042);
and U9160 (N_9160,N_9044,N_9042);
or U9161 (N_9161,N_9020,N_9014);
or U9162 (N_9162,N_9032,N_9054);
and U9163 (N_9163,N_9084,N_9027);
and U9164 (N_9164,N_9028,N_9059);
xor U9165 (N_9165,N_9093,N_9039);
and U9166 (N_9166,N_9018,N_9076);
nand U9167 (N_9167,N_9049,N_9067);
nor U9168 (N_9168,N_9073,N_9054);
nor U9169 (N_9169,N_9021,N_9082);
nand U9170 (N_9170,N_9084,N_9045);
nand U9171 (N_9171,N_9095,N_9062);
nor U9172 (N_9172,N_9055,N_9083);
and U9173 (N_9173,N_9012,N_9022);
nor U9174 (N_9174,N_9040,N_9080);
nor U9175 (N_9175,N_9014,N_9045);
and U9176 (N_9176,N_9061,N_9026);
and U9177 (N_9177,N_9025,N_9083);
and U9178 (N_9178,N_9047,N_9077);
nand U9179 (N_9179,N_9081,N_9094);
nor U9180 (N_9180,N_9055,N_9084);
and U9181 (N_9181,N_9078,N_9083);
nand U9182 (N_9182,N_9056,N_9007);
and U9183 (N_9183,N_9063,N_9011);
xor U9184 (N_9184,N_9073,N_9037);
xor U9185 (N_9185,N_9095,N_9098);
xnor U9186 (N_9186,N_9067,N_9034);
and U9187 (N_9187,N_9025,N_9005);
nand U9188 (N_9188,N_9023,N_9035);
nor U9189 (N_9189,N_9040,N_9065);
xor U9190 (N_9190,N_9061,N_9033);
and U9191 (N_9191,N_9086,N_9029);
and U9192 (N_9192,N_9049,N_9098);
nor U9193 (N_9193,N_9047,N_9024);
or U9194 (N_9194,N_9017,N_9073);
and U9195 (N_9195,N_9034,N_9045);
and U9196 (N_9196,N_9028,N_9023);
nand U9197 (N_9197,N_9017,N_9018);
nand U9198 (N_9198,N_9024,N_9068);
and U9199 (N_9199,N_9050,N_9062);
nor U9200 (N_9200,N_9192,N_9168);
nand U9201 (N_9201,N_9193,N_9107);
nor U9202 (N_9202,N_9157,N_9105);
and U9203 (N_9203,N_9182,N_9123);
nor U9204 (N_9204,N_9172,N_9141);
nor U9205 (N_9205,N_9116,N_9163);
and U9206 (N_9206,N_9101,N_9135);
and U9207 (N_9207,N_9130,N_9176);
nand U9208 (N_9208,N_9185,N_9184);
and U9209 (N_9209,N_9125,N_9146);
nand U9210 (N_9210,N_9162,N_9165);
nor U9211 (N_9211,N_9199,N_9147);
nand U9212 (N_9212,N_9197,N_9100);
nand U9213 (N_9213,N_9189,N_9171);
and U9214 (N_9214,N_9113,N_9183);
nor U9215 (N_9215,N_9102,N_9117);
or U9216 (N_9216,N_9198,N_9140);
xor U9217 (N_9217,N_9177,N_9187);
xnor U9218 (N_9218,N_9128,N_9188);
nor U9219 (N_9219,N_9196,N_9155);
and U9220 (N_9220,N_9137,N_9112);
or U9221 (N_9221,N_9148,N_9114);
nor U9222 (N_9222,N_9153,N_9110);
and U9223 (N_9223,N_9122,N_9191);
nor U9224 (N_9224,N_9111,N_9195);
and U9225 (N_9225,N_9156,N_9170);
nor U9226 (N_9226,N_9138,N_9154);
or U9227 (N_9227,N_9190,N_9144);
or U9228 (N_9228,N_9134,N_9126);
or U9229 (N_9229,N_9103,N_9180);
nand U9230 (N_9230,N_9127,N_9106);
and U9231 (N_9231,N_9139,N_9159);
nand U9232 (N_9232,N_9150,N_9119);
or U9233 (N_9233,N_9121,N_9152);
or U9234 (N_9234,N_9186,N_9151);
nor U9235 (N_9235,N_9118,N_9108);
xnor U9236 (N_9236,N_9179,N_9115);
or U9237 (N_9237,N_9161,N_9129);
nor U9238 (N_9238,N_9149,N_9104);
nor U9239 (N_9239,N_9109,N_9132);
nor U9240 (N_9240,N_9181,N_9167);
nand U9241 (N_9241,N_9194,N_9120);
or U9242 (N_9242,N_9174,N_9169);
nand U9243 (N_9243,N_9131,N_9136);
nor U9244 (N_9244,N_9173,N_9158);
xnor U9245 (N_9245,N_9166,N_9178);
nor U9246 (N_9246,N_9145,N_9175);
or U9247 (N_9247,N_9164,N_9142);
or U9248 (N_9248,N_9133,N_9160);
nor U9249 (N_9249,N_9124,N_9143);
or U9250 (N_9250,N_9129,N_9142);
and U9251 (N_9251,N_9141,N_9126);
or U9252 (N_9252,N_9198,N_9165);
or U9253 (N_9253,N_9120,N_9184);
or U9254 (N_9254,N_9113,N_9102);
or U9255 (N_9255,N_9103,N_9115);
or U9256 (N_9256,N_9169,N_9186);
or U9257 (N_9257,N_9173,N_9147);
nor U9258 (N_9258,N_9152,N_9151);
nand U9259 (N_9259,N_9117,N_9168);
and U9260 (N_9260,N_9107,N_9125);
nor U9261 (N_9261,N_9104,N_9131);
nand U9262 (N_9262,N_9154,N_9118);
nand U9263 (N_9263,N_9199,N_9124);
and U9264 (N_9264,N_9145,N_9162);
and U9265 (N_9265,N_9165,N_9166);
nand U9266 (N_9266,N_9155,N_9145);
and U9267 (N_9267,N_9193,N_9139);
nand U9268 (N_9268,N_9170,N_9106);
or U9269 (N_9269,N_9117,N_9149);
or U9270 (N_9270,N_9168,N_9140);
or U9271 (N_9271,N_9194,N_9125);
nor U9272 (N_9272,N_9153,N_9108);
nor U9273 (N_9273,N_9196,N_9108);
nor U9274 (N_9274,N_9198,N_9183);
nand U9275 (N_9275,N_9126,N_9117);
nand U9276 (N_9276,N_9131,N_9185);
or U9277 (N_9277,N_9169,N_9185);
nor U9278 (N_9278,N_9184,N_9193);
or U9279 (N_9279,N_9156,N_9141);
or U9280 (N_9280,N_9193,N_9131);
nand U9281 (N_9281,N_9188,N_9122);
nand U9282 (N_9282,N_9109,N_9145);
nand U9283 (N_9283,N_9167,N_9182);
or U9284 (N_9284,N_9140,N_9154);
or U9285 (N_9285,N_9102,N_9142);
nand U9286 (N_9286,N_9187,N_9182);
nand U9287 (N_9287,N_9162,N_9154);
or U9288 (N_9288,N_9174,N_9128);
nor U9289 (N_9289,N_9163,N_9140);
and U9290 (N_9290,N_9133,N_9169);
nand U9291 (N_9291,N_9186,N_9103);
or U9292 (N_9292,N_9130,N_9194);
nor U9293 (N_9293,N_9166,N_9122);
xor U9294 (N_9294,N_9108,N_9160);
xor U9295 (N_9295,N_9153,N_9182);
nor U9296 (N_9296,N_9128,N_9119);
nand U9297 (N_9297,N_9175,N_9165);
nand U9298 (N_9298,N_9143,N_9136);
or U9299 (N_9299,N_9126,N_9190);
nor U9300 (N_9300,N_9225,N_9257);
or U9301 (N_9301,N_9217,N_9218);
and U9302 (N_9302,N_9285,N_9263);
xor U9303 (N_9303,N_9210,N_9233);
and U9304 (N_9304,N_9236,N_9216);
or U9305 (N_9305,N_9221,N_9267);
nand U9306 (N_9306,N_9245,N_9275);
or U9307 (N_9307,N_9202,N_9255);
xor U9308 (N_9308,N_9239,N_9244);
nor U9309 (N_9309,N_9259,N_9270);
nor U9310 (N_9310,N_9232,N_9208);
or U9311 (N_9311,N_9246,N_9268);
nor U9312 (N_9312,N_9213,N_9269);
nor U9313 (N_9313,N_9278,N_9280);
nor U9314 (N_9314,N_9237,N_9274);
nand U9315 (N_9315,N_9207,N_9238);
or U9316 (N_9316,N_9228,N_9283);
and U9317 (N_9317,N_9206,N_9250);
nand U9318 (N_9318,N_9289,N_9201);
or U9319 (N_9319,N_9209,N_9200);
or U9320 (N_9320,N_9288,N_9264);
or U9321 (N_9321,N_9277,N_9212);
and U9322 (N_9322,N_9214,N_9254);
xor U9323 (N_9323,N_9235,N_9215);
and U9324 (N_9324,N_9220,N_9260);
or U9325 (N_9325,N_9203,N_9295);
nand U9326 (N_9326,N_9234,N_9296);
or U9327 (N_9327,N_9284,N_9227);
xor U9328 (N_9328,N_9222,N_9229);
nor U9329 (N_9329,N_9298,N_9282);
and U9330 (N_9330,N_9299,N_9291);
xnor U9331 (N_9331,N_9262,N_9211);
and U9332 (N_9332,N_9243,N_9294);
or U9333 (N_9333,N_9223,N_9293);
nand U9334 (N_9334,N_9266,N_9204);
nand U9335 (N_9335,N_9226,N_9272);
nor U9336 (N_9336,N_9292,N_9251);
and U9337 (N_9337,N_9290,N_9241);
and U9338 (N_9338,N_9279,N_9265);
nor U9339 (N_9339,N_9271,N_9240);
or U9340 (N_9340,N_9205,N_9258);
xnor U9341 (N_9341,N_9252,N_9249);
and U9342 (N_9342,N_9276,N_9231);
and U9343 (N_9343,N_9287,N_9253);
and U9344 (N_9344,N_9219,N_9261);
nand U9345 (N_9345,N_9256,N_9247);
or U9346 (N_9346,N_9248,N_9224);
nor U9347 (N_9347,N_9242,N_9230);
nand U9348 (N_9348,N_9286,N_9297);
or U9349 (N_9349,N_9273,N_9281);
or U9350 (N_9350,N_9219,N_9241);
and U9351 (N_9351,N_9217,N_9288);
nand U9352 (N_9352,N_9212,N_9217);
xnor U9353 (N_9353,N_9238,N_9266);
nand U9354 (N_9354,N_9215,N_9271);
and U9355 (N_9355,N_9220,N_9270);
and U9356 (N_9356,N_9273,N_9235);
nand U9357 (N_9357,N_9231,N_9247);
nor U9358 (N_9358,N_9271,N_9226);
xnor U9359 (N_9359,N_9282,N_9234);
xnor U9360 (N_9360,N_9288,N_9246);
xnor U9361 (N_9361,N_9289,N_9238);
nand U9362 (N_9362,N_9295,N_9254);
and U9363 (N_9363,N_9260,N_9286);
or U9364 (N_9364,N_9296,N_9215);
nor U9365 (N_9365,N_9293,N_9284);
and U9366 (N_9366,N_9207,N_9273);
xnor U9367 (N_9367,N_9202,N_9285);
and U9368 (N_9368,N_9260,N_9285);
nand U9369 (N_9369,N_9298,N_9295);
nand U9370 (N_9370,N_9288,N_9247);
nor U9371 (N_9371,N_9268,N_9206);
nor U9372 (N_9372,N_9287,N_9219);
and U9373 (N_9373,N_9237,N_9245);
or U9374 (N_9374,N_9270,N_9223);
nand U9375 (N_9375,N_9211,N_9276);
and U9376 (N_9376,N_9234,N_9242);
and U9377 (N_9377,N_9207,N_9279);
nand U9378 (N_9378,N_9210,N_9232);
and U9379 (N_9379,N_9274,N_9236);
and U9380 (N_9380,N_9256,N_9232);
and U9381 (N_9381,N_9217,N_9241);
nor U9382 (N_9382,N_9294,N_9204);
nand U9383 (N_9383,N_9273,N_9253);
xnor U9384 (N_9384,N_9274,N_9228);
and U9385 (N_9385,N_9265,N_9207);
and U9386 (N_9386,N_9264,N_9271);
or U9387 (N_9387,N_9284,N_9299);
nor U9388 (N_9388,N_9290,N_9204);
or U9389 (N_9389,N_9275,N_9211);
or U9390 (N_9390,N_9286,N_9275);
and U9391 (N_9391,N_9218,N_9262);
or U9392 (N_9392,N_9279,N_9272);
nor U9393 (N_9393,N_9264,N_9259);
and U9394 (N_9394,N_9293,N_9217);
and U9395 (N_9395,N_9251,N_9208);
and U9396 (N_9396,N_9227,N_9291);
xor U9397 (N_9397,N_9225,N_9272);
xor U9398 (N_9398,N_9292,N_9211);
nand U9399 (N_9399,N_9294,N_9262);
or U9400 (N_9400,N_9307,N_9359);
or U9401 (N_9401,N_9375,N_9394);
xnor U9402 (N_9402,N_9308,N_9348);
nor U9403 (N_9403,N_9340,N_9392);
or U9404 (N_9404,N_9391,N_9335);
nor U9405 (N_9405,N_9326,N_9365);
and U9406 (N_9406,N_9373,N_9379);
nand U9407 (N_9407,N_9396,N_9321);
xnor U9408 (N_9408,N_9311,N_9351);
and U9409 (N_9409,N_9328,N_9344);
nand U9410 (N_9410,N_9312,N_9360);
or U9411 (N_9411,N_9370,N_9347);
nand U9412 (N_9412,N_9361,N_9342);
and U9413 (N_9413,N_9304,N_9313);
and U9414 (N_9414,N_9387,N_9358);
or U9415 (N_9415,N_9323,N_9355);
xor U9416 (N_9416,N_9329,N_9374);
nor U9417 (N_9417,N_9363,N_9318);
nand U9418 (N_9418,N_9366,N_9397);
nand U9419 (N_9419,N_9369,N_9305);
or U9420 (N_9420,N_9332,N_9345);
and U9421 (N_9421,N_9325,N_9368);
nor U9422 (N_9422,N_9386,N_9381);
or U9423 (N_9423,N_9362,N_9330);
nand U9424 (N_9424,N_9324,N_9300);
nand U9425 (N_9425,N_9382,N_9364);
or U9426 (N_9426,N_9395,N_9314);
and U9427 (N_9427,N_9333,N_9393);
xor U9428 (N_9428,N_9357,N_9367);
and U9429 (N_9429,N_9320,N_9316);
nand U9430 (N_9430,N_9322,N_9354);
and U9431 (N_9431,N_9377,N_9331);
and U9432 (N_9432,N_9346,N_9327);
nand U9433 (N_9433,N_9385,N_9303);
or U9434 (N_9434,N_9306,N_9352);
xnor U9435 (N_9435,N_9383,N_9302);
nor U9436 (N_9436,N_9398,N_9390);
or U9437 (N_9437,N_9349,N_9336);
nand U9438 (N_9438,N_9317,N_9353);
nand U9439 (N_9439,N_9310,N_9309);
nand U9440 (N_9440,N_9384,N_9301);
nand U9441 (N_9441,N_9350,N_9376);
nand U9442 (N_9442,N_9343,N_9319);
and U9443 (N_9443,N_9399,N_9378);
nor U9444 (N_9444,N_9356,N_9372);
nor U9445 (N_9445,N_9334,N_9338);
xnor U9446 (N_9446,N_9371,N_9339);
xor U9447 (N_9447,N_9337,N_9388);
or U9448 (N_9448,N_9389,N_9341);
and U9449 (N_9449,N_9315,N_9380);
xor U9450 (N_9450,N_9340,N_9323);
nor U9451 (N_9451,N_9337,N_9390);
nor U9452 (N_9452,N_9383,N_9319);
and U9453 (N_9453,N_9353,N_9371);
nand U9454 (N_9454,N_9371,N_9382);
and U9455 (N_9455,N_9385,N_9358);
or U9456 (N_9456,N_9310,N_9336);
nand U9457 (N_9457,N_9359,N_9370);
or U9458 (N_9458,N_9372,N_9364);
nand U9459 (N_9459,N_9324,N_9343);
nand U9460 (N_9460,N_9396,N_9375);
nand U9461 (N_9461,N_9317,N_9327);
or U9462 (N_9462,N_9312,N_9380);
nand U9463 (N_9463,N_9329,N_9315);
nor U9464 (N_9464,N_9382,N_9376);
nor U9465 (N_9465,N_9365,N_9388);
nor U9466 (N_9466,N_9384,N_9307);
nand U9467 (N_9467,N_9319,N_9389);
nor U9468 (N_9468,N_9341,N_9307);
nand U9469 (N_9469,N_9358,N_9381);
nor U9470 (N_9470,N_9355,N_9366);
nand U9471 (N_9471,N_9389,N_9398);
and U9472 (N_9472,N_9352,N_9367);
and U9473 (N_9473,N_9367,N_9355);
nand U9474 (N_9474,N_9317,N_9320);
xor U9475 (N_9475,N_9339,N_9386);
and U9476 (N_9476,N_9396,N_9355);
nor U9477 (N_9477,N_9324,N_9321);
nor U9478 (N_9478,N_9303,N_9379);
nand U9479 (N_9479,N_9360,N_9392);
xnor U9480 (N_9480,N_9328,N_9350);
nor U9481 (N_9481,N_9343,N_9303);
or U9482 (N_9482,N_9393,N_9348);
and U9483 (N_9483,N_9395,N_9341);
nor U9484 (N_9484,N_9334,N_9370);
and U9485 (N_9485,N_9338,N_9377);
nand U9486 (N_9486,N_9335,N_9330);
nor U9487 (N_9487,N_9318,N_9380);
xnor U9488 (N_9488,N_9398,N_9358);
and U9489 (N_9489,N_9307,N_9387);
or U9490 (N_9490,N_9321,N_9331);
or U9491 (N_9491,N_9352,N_9371);
and U9492 (N_9492,N_9375,N_9351);
and U9493 (N_9493,N_9386,N_9354);
nor U9494 (N_9494,N_9302,N_9323);
nand U9495 (N_9495,N_9366,N_9327);
nor U9496 (N_9496,N_9365,N_9313);
nor U9497 (N_9497,N_9334,N_9343);
xor U9498 (N_9498,N_9335,N_9342);
and U9499 (N_9499,N_9361,N_9360);
and U9500 (N_9500,N_9479,N_9427);
nand U9501 (N_9501,N_9469,N_9497);
nor U9502 (N_9502,N_9420,N_9467);
and U9503 (N_9503,N_9453,N_9465);
xor U9504 (N_9504,N_9408,N_9489);
nand U9505 (N_9505,N_9457,N_9448);
nor U9506 (N_9506,N_9422,N_9468);
or U9507 (N_9507,N_9405,N_9404);
nand U9508 (N_9508,N_9402,N_9439);
nor U9509 (N_9509,N_9424,N_9452);
and U9510 (N_9510,N_9435,N_9407);
nand U9511 (N_9511,N_9464,N_9476);
nor U9512 (N_9512,N_9494,N_9414);
or U9513 (N_9513,N_9425,N_9441);
or U9514 (N_9514,N_9460,N_9406);
nor U9515 (N_9515,N_9477,N_9437);
and U9516 (N_9516,N_9472,N_9456);
or U9517 (N_9517,N_9423,N_9495);
nand U9518 (N_9518,N_9418,N_9438);
nand U9519 (N_9519,N_9454,N_9412);
or U9520 (N_9520,N_9403,N_9411);
nand U9521 (N_9521,N_9442,N_9483);
nand U9522 (N_9522,N_9419,N_9466);
nand U9523 (N_9523,N_9417,N_9447);
nor U9524 (N_9524,N_9455,N_9482);
or U9525 (N_9525,N_9426,N_9491);
or U9526 (N_9526,N_9462,N_9496);
or U9527 (N_9527,N_9400,N_9401);
nor U9528 (N_9528,N_9485,N_9444);
xnor U9529 (N_9529,N_9463,N_9492);
nor U9530 (N_9530,N_9440,N_9471);
xor U9531 (N_9531,N_9487,N_9409);
and U9532 (N_9532,N_9413,N_9474);
nand U9533 (N_9533,N_9436,N_9450);
or U9534 (N_9534,N_9484,N_9459);
nor U9535 (N_9535,N_9416,N_9431);
and U9536 (N_9536,N_9493,N_9430);
nor U9537 (N_9537,N_9488,N_9486);
or U9538 (N_9538,N_9458,N_9499);
and U9539 (N_9539,N_9481,N_9445);
or U9540 (N_9540,N_9478,N_9451);
or U9541 (N_9541,N_9449,N_9410);
or U9542 (N_9542,N_9434,N_9446);
nand U9543 (N_9543,N_9461,N_9473);
or U9544 (N_9544,N_9470,N_9433);
and U9545 (N_9545,N_9490,N_9432);
and U9546 (N_9546,N_9498,N_9428);
nor U9547 (N_9547,N_9429,N_9475);
nand U9548 (N_9548,N_9443,N_9415);
nor U9549 (N_9549,N_9421,N_9480);
and U9550 (N_9550,N_9494,N_9446);
nor U9551 (N_9551,N_9442,N_9485);
and U9552 (N_9552,N_9482,N_9479);
and U9553 (N_9553,N_9416,N_9442);
or U9554 (N_9554,N_9467,N_9490);
nand U9555 (N_9555,N_9489,N_9499);
and U9556 (N_9556,N_9456,N_9487);
nor U9557 (N_9557,N_9449,N_9418);
or U9558 (N_9558,N_9420,N_9474);
nor U9559 (N_9559,N_9485,N_9464);
nand U9560 (N_9560,N_9468,N_9434);
nand U9561 (N_9561,N_9415,N_9425);
nor U9562 (N_9562,N_9441,N_9483);
or U9563 (N_9563,N_9477,N_9480);
or U9564 (N_9564,N_9446,N_9403);
xnor U9565 (N_9565,N_9491,N_9474);
nor U9566 (N_9566,N_9427,N_9490);
nand U9567 (N_9567,N_9467,N_9483);
and U9568 (N_9568,N_9428,N_9405);
xor U9569 (N_9569,N_9413,N_9427);
and U9570 (N_9570,N_9490,N_9451);
or U9571 (N_9571,N_9460,N_9420);
and U9572 (N_9572,N_9423,N_9451);
or U9573 (N_9573,N_9468,N_9461);
or U9574 (N_9574,N_9491,N_9417);
nand U9575 (N_9575,N_9431,N_9460);
xnor U9576 (N_9576,N_9461,N_9432);
nand U9577 (N_9577,N_9492,N_9451);
and U9578 (N_9578,N_9403,N_9469);
nand U9579 (N_9579,N_9444,N_9479);
nor U9580 (N_9580,N_9499,N_9429);
and U9581 (N_9581,N_9431,N_9468);
nand U9582 (N_9582,N_9427,N_9423);
or U9583 (N_9583,N_9486,N_9481);
nor U9584 (N_9584,N_9404,N_9402);
xnor U9585 (N_9585,N_9491,N_9497);
nor U9586 (N_9586,N_9480,N_9420);
nor U9587 (N_9587,N_9459,N_9432);
nor U9588 (N_9588,N_9482,N_9438);
nand U9589 (N_9589,N_9467,N_9435);
nor U9590 (N_9590,N_9490,N_9422);
nor U9591 (N_9591,N_9486,N_9469);
and U9592 (N_9592,N_9463,N_9440);
or U9593 (N_9593,N_9498,N_9454);
nor U9594 (N_9594,N_9476,N_9467);
and U9595 (N_9595,N_9406,N_9462);
xor U9596 (N_9596,N_9475,N_9421);
nor U9597 (N_9597,N_9481,N_9413);
nand U9598 (N_9598,N_9469,N_9402);
nand U9599 (N_9599,N_9414,N_9404);
nor U9600 (N_9600,N_9576,N_9525);
nor U9601 (N_9601,N_9583,N_9500);
and U9602 (N_9602,N_9567,N_9516);
or U9603 (N_9603,N_9529,N_9526);
or U9604 (N_9604,N_9573,N_9505);
or U9605 (N_9605,N_9569,N_9511);
xor U9606 (N_9606,N_9544,N_9589);
and U9607 (N_9607,N_9534,N_9515);
nand U9608 (N_9608,N_9575,N_9501);
or U9609 (N_9609,N_9545,N_9561);
nor U9610 (N_9610,N_9597,N_9558);
and U9611 (N_9611,N_9565,N_9587);
or U9612 (N_9612,N_9527,N_9586);
and U9613 (N_9613,N_9564,N_9510);
nor U9614 (N_9614,N_9508,N_9572);
nand U9615 (N_9615,N_9532,N_9530);
or U9616 (N_9616,N_9533,N_9518);
and U9617 (N_9617,N_9522,N_9524);
and U9618 (N_9618,N_9568,N_9531);
or U9619 (N_9619,N_9549,N_9566);
and U9620 (N_9620,N_9560,N_9584);
nand U9621 (N_9621,N_9588,N_9535);
and U9622 (N_9622,N_9595,N_9563);
nand U9623 (N_9623,N_9541,N_9581);
or U9624 (N_9624,N_9578,N_9593);
or U9625 (N_9625,N_9553,N_9542);
nand U9626 (N_9626,N_9521,N_9536);
and U9627 (N_9627,N_9571,N_9552);
or U9628 (N_9628,N_9537,N_9598);
or U9629 (N_9629,N_9538,N_9596);
nand U9630 (N_9630,N_9543,N_9546);
and U9631 (N_9631,N_9513,N_9502);
or U9632 (N_9632,N_9550,N_9555);
or U9633 (N_9633,N_9574,N_9539);
nor U9634 (N_9634,N_9519,N_9556);
nor U9635 (N_9635,N_9557,N_9523);
nand U9636 (N_9636,N_9594,N_9590);
and U9637 (N_9637,N_9599,N_9514);
or U9638 (N_9638,N_9580,N_9582);
or U9639 (N_9639,N_9548,N_9509);
or U9640 (N_9640,N_9528,N_9503);
or U9641 (N_9641,N_9547,N_9559);
or U9642 (N_9642,N_9551,N_9562);
and U9643 (N_9643,N_9506,N_9577);
or U9644 (N_9644,N_9504,N_9554);
or U9645 (N_9645,N_9570,N_9520);
nor U9646 (N_9646,N_9591,N_9540);
nor U9647 (N_9647,N_9507,N_9512);
or U9648 (N_9648,N_9517,N_9592);
nor U9649 (N_9649,N_9579,N_9585);
nand U9650 (N_9650,N_9550,N_9542);
nor U9651 (N_9651,N_9503,N_9599);
nor U9652 (N_9652,N_9512,N_9550);
nor U9653 (N_9653,N_9511,N_9526);
nor U9654 (N_9654,N_9598,N_9527);
or U9655 (N_9655,N_9524,N_9514);
nor U9656 (N_9656,N_9510,N_9591);
nor U9657 (N_9657,N_9570,N_9569);
xnor U9658 (N_9658,N_9525,N_9575);
xnor U9659 (N_9659,N_9527,N_9504);
nor U9660 (N_9660,N_9537,N_9505);
nand U9661 (N_9661,N_9556,N_9547);
nand U9662 (N_9662,N_9527,N_9570);
xor U9663 (N_9663,N_9501,N_9596);
and U9664 (N_9664,N_9596,N_9565);
nor U9665 (N_9665,N_9560,N_9517);
or U9666 (N_9666,N_9597,N_9514);
nand U9667 (N_9667,N_9561,N_9569);
nand U9668 (N_9668,N_9508,N_9595);
nand U9669 (N_9669,N_9567,N_9566);
and U9670 (N_9670,N_9549,N_9507);
xnor U9671 (N_9671,N_9567,N_9545);
nor U9672 (N_9672,N_9537,N_9570);
nand U9673 (N_9673,N_9588,N_9562);
nand U9674 (N_9674,N_9530,N_9515);
nand U9675 (N_9675,N_9508,N_9560);
nor U9676 (N_9676,N_9551,N_9578);
and U9677 (N_9677,N_9506,N_9553);
or U9678 (N_9678,N_9536,N_9533);
nand U9679 (N_9679,N_9550,N_9526);
xor U9680 (N_9680,N_9548,N_9502);
nand U9681 (N_9681,N_9587,N_9568);
nand U9682 (N_9682,N_9566,N_9598);
or U9683 (N_9683,N_9593,N_9568);
or U9684 (N_9684,N_9521,N_9522);
or U9685 (N_9685,N_9523,N_9508);
nor U9686 (N_9686,N_9516,N_9507);
or U9687 (N_9687,N_9582,N_9534);
nor U9688 (N_9688,N_9589,N_9542);
nand U9689 (N_9689,N_9529,N_9519);
nand U9690 (N_9690,N_9587,N_9529);
nor U9691 (N_9691,N_9504,N_9545);
or U9692 (N_9692,N_9585,N_9506);
nor U9693 (N_9693,N_9511,N_9576);
and U9694 (N_9694,N_9559,N_9549);
or U9695 (N_9695,N_9520,N_9551);
xor U9696 (N_9696,N_9585,N_9550);
and U9697 (N_9697,N_9586,N_9579);
nor U9698 (N_9698,N_9577,N_9595);
xnor U9699 (N_9699,N_9544,N_9550);
nand U9700 (N_9700,N_9691,N_9604);
and U9701 (N_9701,N_9678,N_9603);
and U9702 (N_9702,N_9682,N_9653);
nor U9703 (N_9703,N_9624,N_9660);
and U9704 (N_9704,N_9622,N_9621);
or U9705 (N_9705,N_9607,N_9662);
or U9706 (N_9706,N_9698,N_9601);
xnor U9707 (N_9707,N_9658,N_9697);
nor U9708 (N_9708,N_9666,N_9618);
nor U9709 (N_9709,N_9628,N_9664);
and U9710 (N_9710,N_9668,N_9687);
and U9711 (N_9711,N_9656,N_9629);
and U9712 (N_9712,N_9611,N_9659);
nand U9713 (N_9713,N_9692,N_9644);
and U9714 (N_9714,N_9630,N_9600);
nor U9715 (N_9715,N_9674,N_9670);
or U9716 (N_9716,N_9680,N_9615);
nand U9717 (N_9717,N_9688,N_9679);
nand U9718 (N_9718,N_9627,N_9602);
and U9719 (N_9719,N_9635,N_9665);
nor U9720 (N_9720,N_9681,N_9605);
and U9721 (N_9721,N_9652,N_9673);
nor U9722 (N_9722,N_9677,N_9657);
nor U9723 (N_9723,N_9610,N_9609);
or U9724 (N_9724,N_9672,N_9650);
and U9725 (N_9725,N_9619,N_9649);
nand U9726 (N_9726,N_9631,N_9651);
nand U9727 (N_9727,N_9616,N_9689);
nor U9728 (N_9728,N_9683,N_9648);
and U9729 (N_9729,N_9647,N_9620);
nand U9730 (N_9730,N_9633,N_9641);
or U9731 (N_9731,N_9695,N_9661);
or U9732 (N_9732,N_9634,N_9671);
and U9733 (N_9733,N_9699,N_9623);
xor U9734 (N_9734,N_9636,N_9694);
nor U9735 (N_9735,N_9608,N_9626);
xor U9736 (N_9736,N_9646,N_9613);
xor U9737 (N_9737,N_9638,N_9676);
or U9738 (N_9738,N_9642,N_9663);
and U9739 (N_9739,N_9617,N_9612);
nor U9740 (N_9740,N_9640,N_9696);
nand U9741 (N_9741,N_9690,N_9675);
and U9742 (N_9742,N_9684,N_9632);
nand U9743 (N_9743,N_9645,N_9639);
and U9744 (N_9744,N_9625,N_9686);
nand U9745 (N_9745,N_9685,N_9614);
and U9746 (N_9746,N_9654,N_9669);
and U9747 (N_9747,N_9693,N_9637);
and U9748 (N_9748,N_9606,N_9655);
and U9749 (N_9749,N_9643,N_9667);
nand U9750 (N_9750,N_9684,N_9660);
and U9751 (N_9751,N_9643,N_9655);
nor U9752 (N_9752,N_9654,N_9648);
xor U9753 (N_9753,N_9645,N_9650);
nor U9754 (N_9754,N_9688,N_9603);
or U9755 (N_9755,N_9669,N_9615);
nor U9756 (N_9756,N_9657,N_9610);
xnor U9757 (N_9757,N_9620,N_9638);
or U9758 (N_9758,N_9630,N_9623);
nor U9759 (N_9759,N_9680,N_9665);
nand U9760 (N_9760,N_9607,N_9601);
nor U9761 (N_9761,N_9660,N_9669);
nor U9762 (N_9762,N_9663,N_9622);
nand U9763 (N_9763,N_9636,N_9642);
nor U9764 (N_9764,N_9642,N_9620);
or U9765 (N_9765,N_9682,N_9650);
and U9766 (N_9766,N_9633,N_9639);
nand U9767 (N_9767,N_9618,N_9622);
and U9768 (N_9768,N_9603,N_9616);
nor U9769 (N_9769,N_9609,N_9667);
nor U9770 (N_9770,N_9615,N_9668);
nand U9771 (N_9771,N_9605,N_9619);
or U9772 (N_9772,N_9607,N_9617);
nand U9773 (N_9773,N_9622,N_9628);
nor U9774 (N_9774,N_9665,N_9676);
nand U9775 (N_9775,N_9635,N_9689);
or U9776 (N_9776,N_9693,N_9682);
nand U9777 (N_9777,N_9646,N_9653);
nand U9778 (N_9778,N_9690,N_9689);
nor U9779 (N_9779,N_9606,N_9699);
nor U9780 (N_9780,N_9626,N_9623);
and U9781 (N_9781,N_9672,N_9640);
nor U9782 (N_9782,N_9626,N_9655);
and U9783 (N_9783,N_9693,N_9647);
and U9784 (N_9784,N_9677,N_9621);
xor U9785 (N_9785,N_9602,N_9617);
or U9786 (N_9786,N_9618,N_9652);
and U9787 (N_9787,N_9681,N_9630);
nand U9788 (N_9788,N_9661,N_9693);
xor U9789 (N_9789,N_9655,N_9693);
and U9790 (N_9790,N_9603,N_9686);
and U9791 (N_9791,N_9615,N_9692);
nor U9792 (N_9792,N_9683,N_9646);
or U9793 (N_9793,N_9654,N_9684);
or U9794 (N_9794,N_9635,N_9632);
nand U9795 (N_9795,N_9629,N_9678);
or U9796 (N_9796,N_9677,N_9688);
or U9797 (N_9797,N_9638,N_9692);
or U9798 (N_9798,N_9620,N_9665);
nor U9799 (N_9799,N_9643,N_9621);
nor U9800 (N_9800,N_9716,N_9737);
and U9801 (N_9801,N_9776,N_9787);
nor U9802 (N_9802,N_9745,N_9798);
or U9803 (N_9803,N_9765,N_9789);
and U9804 (N_9804,N_9780,N_9781);
nor U9805 (N_9805,N_9788,N_9760);
or U9806 (N_9806,N_9772,N_9700);
nor U9807 (N_9807,N_9732,N_9771);
and U9808 (N_9808,N_9755,N_9719);
nand U9809 (N_9809,N_9785,N_9795);
nor U9810 (N_9810,N_9769,N_9726);
or U9811 (N_9811,N_9753,N_9724);
or U9812 (N_9812,N_9773,N_9704);
nand U9813 (N_9813,N_9757,N_9743);
nor U9814 (N_9814,N_9761,N_9746);
xnor U9815 (N_9815,N_9793,N_9767);
xor U9816 (N_9816,N_9763,N_9723);
or U9817 (N_9817,N_9703,N_9791);
xnor U9818 (N_9818,N_9779,N_9735);
nand U9819 (N_9819,N_9749,N_9750);
xor U9820 (N_9820,N_9775,N_9734);
nor U9821 (N_9821,N_9748,N_9701);
nand U9822 (N_9822,N_9786,N_9783);
and U9823 (N_9823,N_9728,N_9758);
or U9824 (N_9824,N_9764,N_9727);
or U9825 (N_9825,N_9790,N_9722);
xor U9826 (N_9826,N_9740,N_9706);
xor U9827 (N_9827,N_9709,N_9762);
xnor U9828 (N_9828,N_9799,N_9797);
xor U9829 (N_9829,N_9759,N_9739);
nor U9830 (N_9830,N_9707,N_9730);
or U9831 (N_9831,N_9725,N_9796);
xnor U9832 (N_9832,N_9784,N_9733);
and U9833 (N_9833,N_9747,N_9756);
nor U9834 (N_9834,N_9778,N_9768);
xnor U9835 (N_9835,N_9744,N_9782);
and U9836 (N_9836,N_9794,N_9754);
nor U9837 (N_9837,N_9741,N_9792);
nand U9838 (N_9838,N_9711,N_9717);
or U9839 (N_9839,N_9742,N_9715);
and U9840 (N_9840,N_9736,N_9713);
or U9841 (N_9841,N_9752,N_9721);
xnor U9842 (N_9842,N_9718,N_9702);
nor U9843 (N_9843,N_9710,N_9708);
or U9844 (N_9844,N_9766,N_9705);
or U9845 (N_9845,N_9720,N_9714);
or U9846 (N_9846,N_9774,N_9751);
nor U9847 (N_9847,N_9770,N_9729);
xor U9848 (N_9848,N_9777,N_9712);
nor U9849 (N_9849,N_9738,N_9731);
xnor U9850 (N_9850,N_9797,N_9700);
or U9851 (N_9851,N_9750,N_9737);
or U9852 (N_9852,N_9712,N_9775);
nand U9853 (N_9853,N_9793,N_9762);
nand U9854 (N_9854,N_9702,N_9761);
or U9855 (N_9855,N_9770,N_9741);
xnor U9856 (N_9856,N_9792,N_9729);
nor U9857 (N_9857,N_9778,N_9799);
and U9858 (N_9858,N_9778,N_9786);
nor U9859 (N_9859,N_9773,N_9754);
and U9860 (N_9860,N_9762,N_9765);
or U9861 (N_9861,N_9793,N_9755);
nor U9862 (N_9862,N_9705,N_9796);
nor U9863 (N_9863,N_9747,N_9787);
nor U9864 (N_9864,N_9720,N_9779);
or U9865 (N_9865,N_9712,N_9747);
and U9866 (N_9866,N_9783,N_9707);
nand U9867 (N_9867,N_9784,N_9712);
or U9868 (N_9868,N_9777,N_9734);
nor U9869 (N_9869,N_9714,N_9778);
nor U9870 (N_9870,N_9733,N_9757);
nand U9871 (N_9871,N_9796,N_9745);
nand U9872 (N_9872,N_9739,N_9783);
nand U9873 (N_9873,N_9727,N_9706);
xnor U9874 (N_9874,N_9721,N_9753);
xor U9875 (N_9875,N_9715,N_9727);
and U9876 (N_9876,N_9704,N_9729);
or U9877 (N_9877,N_9767,N_9781);
nor U9878 (N_9878,N_9731,N_9742);
nor U9879 (N_9879,N_9797,N_9751);
nand U9880 (N_9880,N_9713,N_9776);
or U9881 (N_9881,N_9773,N_9718);
nand U9882 (N_9882,N_9792,N_9705);
nand U9883 (N_9883,N_9705,N_9725);
nand U9884 (N_9884,N_9717,N_9762);
nand U9885 (N_9885,N_9780,N_9796);
or U9886 (N_9886,N_9746,N_9716);
nand U9887 (N_9887,N_9797,N_9779);
and U9888 (N_9888,N_9791,N_9770);
or U9889 (N_9889,N_9764,N_9784);
or U9890 (N_9890,N_9724,N_9719);
and U9891 (N_9891,N_9792,N_9731);
nor U9892 (N_9892,N_9761,N_9731);
xor U9893 (N_9893,N_9745,N_9794);
nor U9894 (N_9894,N_9752,N_9753);
and U9895 (N_9895,N_9795,N_9736);
or U9896 (N_9896,N_9762,N_9760);
and U9897 (N_9897,N_9721,N_9756);
or U9898 (N_9898,N_9782,N_9748);
nand U9899 (N_9899,N_9709,N_9703);
nand U9900 (N_9900,N_9879,N_9871);
nand U9901 (N_9901,N_9856,N_9852);
nor U9902 (N_9902,N_9876,N_9839);
xor U9903 (N_9903,N_9866,N_9834);
or U9904 (N_9904,N_9802,N_9803);
and U9905 (N_9905,N_9867,N_9804);
or U9906 (N_9906,N_9831,N_9877);
nor U9907 (N_9907,N_9864,N_9884);
or U9908 (N_9908,N_9848,N_9891);
and U9909 (N_9909,N_9892,N_9813);
nor U9910 (N_9910,N_9816,N_9889);
and U9911 (N_9911,N_9821,N_9888);
nor U9912 (N_9912,N_9832,N_9808);
or U9913 (N_9913,N_9815,N_9847);
nand U9914 (N_9914,N_9833,N_9817);
nand U9915 (N_9915,N_9878,N_9811);
or U9916 (N_9916,N_9875,N_9827);
nor U9917 (N_9917,N_9899,N_9860);
xor U9918 (N_9918,N_9826,N_9896);
or U9919 (N_9919,N_9828,N_9897);
or U9920 (N_9920,N_9810,N_9812);
nand U9921 (N_9921,N_9806,N_9825);
nand U9922 (N_9922,N_9845,N_9869);
and U9923 (N_9923,N_9873,N_9870);
or U9924 (N_9924,N_9843,N_9880);
nand U9925 (N_9925,N_9820,N_9865);
and U9926 (N_9926,N_9849,N_9835);
nor U9927 (N_9927,N_9838,N_9822);
xor U9928 (N_9928,N_9801,N_9814);
nand U9929 (N_9929,N_9872,N_9885);
nand U9930 (N_9930,N_9824,N_9861);
and U9931 (N_9931,N_9823,N_9800);
and U9932 (N_9932,N_9818,N_9836);
nand U9933 (N_9933,N_9819,N_9853);
nor U9934 (N_9934,N_9851,N_9883);
nand U9935 (N_9935,N_9855,N_9807);
and U9936 (N_9936,N_9841,N_9858);
and U9937 (N_9937,N_9863,N_9882);
xnor U9938 (N_9938,N_9805,N_9859);
nor U9939 (N_9939,N_9857,N_9850);
and U9940 (N_9940,N_9844,N_9840);
or U9941 (N_9941,N_9829,N_9842);
xnor U9942 (N_9942,N_9890,N_9837);
nor U9943 (N_9943,N_9893,N_9830);
nand U9944 (N_9944,N_9874,N_9881);
xnor U9945 (N_9945,N_9862,N_9898);
nor U9946 (N_9946,N_9894,N_9895);
or U9947 (N_9947,N_9846,N_9854);
and U9948 (N_9948,N_9887,N_9809);
and U9949 (N_9949,N_9868,N_9886);
nor U9950 (N_9950,N_9858,N_9899);
nand U9951 (N_9951,N_9892,N_9829);
nand U9952 (N_9952,N_9883,N_9817);
and U9953 (N_9953,N_9827,N_9890);
nor U9954 (N_9954,N_9860,N_9873);
and U9955 (N_9955,N_9889,N_9896);
nand U9956 (N_9956,N_9843,N_9847);
and U9957 (N_9957,N_9826,N_9899);
or U9958 (N_9958,N_9872,N_9894);
and U9959 (N_9959,N_9826,N_9820);
nor U9960 (N_9960,N_9896,N_9867);
or U9961 (N_9961,N_9853,N_9860);
and U9962 (N_9962,N_9893,N_9878);
and U9963 (N_9963,N_9885,N_9893);
nand U9964 (N_9964,N_9804,N_9830);
nor U9965 (N_9965,N_9890,N_9839);
nor U9966 (N_9966,N_9863,N_9867);
and U9967 (N_9967,N_9840,N_9819);
nand U9968 (N_9968,N_9832,N_9825);
nor U9969 (N_9969,N_9867,N_9888);
nor U9970 (N_9970,N_9809,N_9862);
xor U9971 (N_9971,N_9838,N_9836);
nand U9972 (N_9972,N_9856,N_9892);
or U9973 (N_9973,N_9884,N_9803);
and U9974 (N_9974,N_9827,N_9803);
or U9975 (N_9975,N_9896,N_9817);
or U9976 (N_9976,N_9882,N_9816);
or U9977 (N_9977,N_9886,N_9882);
nor U9978 (N_9978,N_9803,N_9887);
nand U9979 (N_9979,N_9800,N_9897);
and U9980 (N_9980,N_9825,N_9834);
xnor U9981 (N_9981,N_9874,N_9855);
or U9982 (N_9982,N_9891,N_9858);
xnor U9983 (N_9983,N_9848,N_9874);
or U9984 (N_9984,N_9814,N_9886);
nor U9985 (N_9985,N_9838,N_9872);
or U9986 (N_9986,N_9822,N_9862);
nor U9987 (N_9987,N_9887,N_9847);
nor U9988 (N_9988,N_9899,N_9846);
and U9989 (N_9989,N_9895,N_9882);
nand U9990 (N_9990,N_9840,N_9866);
nor U9991 (N_9991,N_9820,N_9834);
nor U9992 (N_9992,N_9836,N_9850);
nand U9993 (N_9993,N_9804,N_9868);
nor U9994 (N_9994,N_9835,N_9831);
and U9995 (N_9995,N_9872,N_9876);
nand U9996 (N_9996,N_9850,N_9899);
nor U9997 (N_9997,N_9849,N_9825);
nand U9998 (N_9998,N_9882,N_9832);
and U9999 (N_9999,N_9861,N_9821);
xor UO_0 (O_0,N_9961,N_9973);
xnor UO_1 (O_1,N_9984,N_9918);
xnor UO_2 (O_2,N_9944,N_9996);
nand UO_3 (O_3,N_9939,N_9903);
or UO_4 (O_4,N_9920,N_9953);
nor UO_5 (O_5,N_9974,N_9945);
or UO_6 (O_6,N_9959,N_9917);
nand UO_7 (O_7,N_9949,N_9999);
or UO_8 (O_8,N_9993,N_9971);
or UO_9 (O_9,N_9985,N_9938);
nand UO_10 (O_10,N_9929,N_9921);
xor UO_11 (O_11,N_9976,N_9955);
nand UO_12 (O_12,N_9979,N_9924);
or UO_13 (O_13,N_9947,N_9987);
nand UO_14 (O_14,N_9998,N_9957);
and UO_15 (O_15,N_9995,N_9923);
nor UO_16 (O_16,N_9925,N_9915);
or UO_17 (O_17,N_9963,N_9982);
xor UO_18 (O_18,N_9966,N_9960);
or UO_19 (O_19,N_9919,N_9901);
nor UO_20 (O_20,N_9900,N_9911);
or UO_21 (O_21,N_9986,N_9977);
or UO_22 (O_22,N_9978,N_9990);
nand UO_23 (O_23,N_9934,N_9981);
xnor UO_24 (O_24,N_9926,N_9950);
or UO_25 (O_25,N_9922,N_9935);
nor UO_26 (O_26,N_9928,N_9933);
nor UO_27 (O_27,N_9954,N_9969);
or UO_28 (O_28,N_9983,N_9989);
and UO_29 (O_29,N_9916,N_9940);
nand UO_30 (O_30,N_9946,N_9906);
xnor UO_31 (O_31,N_9997,N_9937);
or UO_32 (O_32,N_9942,N_9904);
or UO_33 (O_33,N_9936,N_9948);
or UO_34 (O_34,N_9902,N_9980);
or UO_35 (O_35,N_9913,N_9943);
nor UO_36 (O_36,N_9962,N_9912);
or UO_37 (O_37,N_9908,N_9931);
nand UO_38 (O_38,N_9970,N_9909);
and UO_39 (O_39,N_9992,N_9968);
nor UO_40 (O_40,N_9965,N_9907);
and UO_41 (O_41,N_9975,N_9956);
or UO_42 (O_42,N_9958,N_9927);
or UO_43 (O_43,N_9952,N_9932);
xor UO_44 (O_44,N_9905,N_9914);
xnor UO_45 (O_45,N_9930,N_9910);
nand UO_46 (O_46,N_9964,N_9951);
and UO_47 (O_47,N_9941,N_9988);
and UO_48 (O_48,N_9967,N_9991);
and UO_49 (O_49,N_9994,N_9972);
xnor UO_50 (O_50,N_9972,N_9909);
nor UO_51 (O_51,N_9930,N_9933);
and UO_52 (O_52,N_9945,N_9997);
or UO_53 (O_53,N_9970,N_9966);
and UO_54 (O_54,N_9910,N_9916);
nand UO_55 (O_55,N_9936,N_9956);
nor UO_56 (O_56,N_9976,N_9950);
nor UO_57 (O_57,N_9938,N_9920);
or UO_58 (O_58,N_9992,N_9902);
nor UO_59 (O_59,N_9930,N_9966);
or UO_60 (O_60,N_9922,N_9907);
nand UO_61 (O_61,N_9956,N_9989);
nand UO_62 (O_62,N_9950,N_9943);
or UO_63 (O_63,N_9981,N_9918);
nand UO_64 (O_64,N_9961,N_9929);
nand UO_65 (O_65,N_9921,N_9956);
nor UO_66 (O_66,N_9909,N_9968);
or UO_67 (O_67,N_9940,N_9956);
and UO_68 (O_68,N_9909,N_9984);
nand UO_69 (O_69,N_9907,N_9947);
and UO_70 (O_70,N_9939,N_9966);
or UO_71 (O_71,N_9915,N_9960);
nor UO_72 (O_72,N_9990,N_9912);
or UO_73 (O_73,N_9987,N_9996);
and UO_74 (O_74,N_9966,N_9928);
and UO_75 (O_75,N_9983,N_9971);
xor UO_76 (O_76,N_9949,N_9978);
nor UO_77 (O_77,N_9986,N_9939);
nand UO_78 (O_78,N_9936,N_9930);
nor UO_79 (O_79,N_9962,N_9956);
and UO_80 (O_80,N_9954,N_9931);
and UO_81 (O_81,N_9928,N_9957);
nand UO_82 (O_82,N_9978,N_9943);
or UO_83 (O_83,N_9979,N_9953);
nand UO_84 (O_84,N_9998,N_9982);
or UO_85 (O_85,N_9918,N_9906);
or UO_86 (O_86,N_9923,N_9999);
nor UO_87 (O_87,N_9950,N_9958);
nand UO_88 (O_88,N_9944,N_9902);
nand UO_89 (O_89,N_9944,N_9920);
nor UO_90 (O_90,N_9963,N_9987);
nor UO_91 (O_91,N_9919,N_9900);
nand UO_92 (O_92,N_9968,N_9953);
nand UO_93 (O_93,N_9938,N_9974);
and UO_94 (O_94,N_9919,N_9958);
or UO_95 (O_95,N_9900,N_9915);
or UO_96 (O_96,N_9991,N_9936);
or UO_97 (O_97,N_9994,N_9933);
or UO_98 (O_98,N_9913,N_9904);
nor UO_99 (O_99,N_9982,N_9947);
nor UO_100 (O_100,N_9902,N_9918);
nor UO_101 (O_101,N_9981,N_9920);
or UO_102 (O_102,N_9998,N_9979);
xnor UO_103 (O_103,N_9972,N_9970);
and UO_104 (O_104,N_9930,N_9924);
nor UO_105 (O_105,N_9916,N_9995);
and UO_106 (O_106,N_9961,N_9994);
and UO_107 (O_107,N_9994,N_9913);
and UO_108 (O_108,N_9934,N_9922);
nor UO_109 (O_109,N_9939,N_9959);
nor UO_110 (O_110,N_9997,N_9990);
nand UO_111 (O_111,N_9911,N_9913);
and UO_112 (O_112,N_9999,N_9910);
and UO_113 (O_113,N_9946,N_9954);
or UO_114 (O_114,N_9903,N_9953);
nand UO_115 (O_115,N_9937,N_9931);
and UO_116 (O_116,N_9925,N_9985);
nand UO_117 (O_117,N_9906,N_9964);
nand UO_118 (O_118,N_9914,N_9979);
nand UO_119 (O_119,N_9995,N_9924);
and UO_120 (O_120,N_9930,N_9976);
or UO_121 (O_121,N_9947,N_9967);
nand UO_122 (O_122,N_9916,N_9941);
and UO_123 (O_123,N_9944,N_9979);
and UO_124 (O_124,N_9915,N_9957);
nand UO_125 (O_125,N_9910,N_9996);
nor UO_126 (O_126,N_9955,N_9927);
or UO_127 (O_127,N_9905,N_9929);
and UO_128 (O_128,N_9911,N_9979);
or UO_129 (O_129,N_9929,N_9983);
or UO_130 (O_130,N_9997,N_9909);
and UO_131 (O_131,N_9935,N_9966);
and UO_132 (O_132,N_9998,N_9976);
nor UO_133 (O_133,N_9963,N_9995);
or UO_134 (O_134,N_9922,N_9906);
nor UO_135 (O_135,N_9909,N_9994);
or UO_136 (O_136,N_9985,N_9902);
nand UO_137 (O_137,N_9989,N_9972);
nand UO_138 (O_138,N_9938,N_9940);
nand UO_139 (O_139,N_9945,N_9988);
nand UO_140 (O_140,N_9991,N_9903);
nand UO_141 (O_141,N_9963,N_9935);
xnor UO_142 (O_142,N_9995,N_9977);
nor UO_143 (O_143,N_9950,N_9928);
nand UO_144 (O_144,N_9937,N_9939);
nand UO_145 (O_145,N_9964,N_9935);
or UO_146 (O_146,N_9962,N_9982);
and UO_147 (O_147,N_9903,N_9960);
nor UO_148 (O_148,N_9939,N_9953);
or UO_149 (O_149,N_9931,N_9929);
and UO_150 (O_150,N_9965,N_9993);
and UO_151 (O_151,N_9916,N_9966);
nor UO_152 (O_152,N_9928,N_9905);
and UO_153 (O_153,N_9900,N_9962);
nand UO_154 (O_154,N_9906,N_9993);
xor UO_155 (O_155,N_9949,N_9967);
or UO_156 (O_156,N_9994,N_9935);
nor UO_157 (O_157,N_9993,N_9969);
nor UO_158 (O_158,N_9975,N_9922);
and UO_159 (O_159,N_9995,N_9908);
nand UO_160 (O_160,N_9943,N_9988);
and UO_161 (O_161,N_9973,N_9987);
xor UO_162 (O_162,N_9983,N_9935);
nor UO_163 (O_163,N_9901,N_9914);
or UO_164 (O_164,N_9981,N_9969);
nor UO_165 (O_165,N_9967,N_9994);
xor UO_166 (O_166,N_9939,N_9987);
xnor UO_167 (O_167,N_9971,N_9906);
and UO_168 (O_168,N_9991,N_9921);
or UO_169 (O_169,N_9951,N_9940);
nor UO_170 (O_170,N_9942,N_9966);
and UO_171 (O_171,N_9956,N_9964);
nor UO_172 (O_172,N_9972,N_9936);
or UO_173 (O_173,N_9932,N_9981);
nor UO_174 (O_174,N_9913,N_9917);
nand UO_175 (O_175,N_9911,N_9925);
and UO_176 (O_176,N_9994,N_9965);
or UO_177 (O_177,N_9949,N_9931);
and UO_178 (O_178,N_9931,N_9989);
xnor UO_179 (O_179,N_9923,N_9905);
nor UO_180 (O_180,N_9902,N_9997);
nand UO_181 (O_181,N_9918,N_9943);
xor UO_182 (O_182,N_9930,N_9991);
nand UO_183 (O_183,N_9913,N_9959);
nand UO_184 (O_184,N_9909,N_9963);
and UO_185 (O_185,N_9994,N_9927);
nand UO_186 (O_186,N_9976,N_9905);
and UO_187 (O_187,N_9938,N_9934);
and UO_188 (O_188,N_9951,N_9966);
nand UO_189 (O_189,N_9976,N_9940);
xor UO_190 (O_190,N_9961,N_9916);
nand UO_191 (O_191,N_9937,N_9930);
and UO_192 (O_192,N_9992,N_9987);
nor UO_193 (O_193,N_9947,N_9985);
nor UO_194 (O_194,N_9978,N_9997);
xnor UO_195 (O_195,N_9962,N_9907);
nor UO_196 (O_196,N_9984,N_9962);
nand UO_197 (O_197,N_9949,N_9922);
or UO_198 (O_198,N_9963,N_9925);
xnor UO_199 (O_199,N_9937,N_9909);
nor UO_200 (O_200,N_9995,N_9994);
nor UO_201 (O_201,N_9923,N_9954);
nand UO_202 (O_202,N_9947,N_9936);
or UO_203 (O_203,N_9906,N_9975);
or UO_204 (O_204,N_9927,N_9980);
and UO_205 (O_205,N_9907,N_9918);
nor UO_206 (O_206,N_9993,N_9951);
nor UO_207 (O_207,N_9991,N_9979);
and UO_208 (O_208,N_9961,N_9984);
and UO_209 (O_209,N_9923,N_9974);
nand UO_210 (O_210,N_9977,N_9997);
and UO_211 (O_211,N_9979,N_9907);
nand UO_212 (O_212,N_9987,N_9967);
nand UO_213 (O_213,N_9984,N_9957);
nand UO_214 (O_214,N_9947,N_9939);
or UO_215 (O_215,N_9987,N_9927);
nand UO_216 (O_216,N_9989,N_9906);
or UO_217 (O_217,N_9906,N_9904);
xor UO_218 (O_218,N_9906,N_9996);
nor UO_219 (O_219,N_9999,N_9976);
nand UO_220 (O_220,N_9973,N_9918);
or UO_221 (O_221,N_9913,N_9970);
nor UO_222 (O_222,N_9906,N_9924);
nor UO_223 (O_223,N_9982,N_9931);
xnor UO_224 (O_224,N_9992,N_9927);
nand UO_225 (O_225,N_9941,N_9954);
and UO_226 (O_226,N_9979,N_9994);
nand UO_227 (O_227,N_9916,N_9920);
and UO_228 (O_228,N_9967,N_9997);
xor UO_229 (O_229,N_9940,N_9994);
and UO_230 (O_230,N_9994,N_9942);
or UO_231 (O_231,N_9927,N_9938);
nand UO_232 (O_232,N_9912,N_9964);
nor UO_233 (O_233,N_9908,N_9982);
or UO_234 (O_234,N_9994,N_9989);
and UO_235 (O_235,N_9983,N_9960);
and UO_236 (O_236,N_9925,N_9931);
nand UO_237 (O_237,N_9926,N_9933);
or UO_238 (O_238,N_9964,N_9966);
xnor UO_239 (O_239,N_9982,N_9923);
nand UO_240 (O_240,N_9955,N_9998);
nor UO_241 (O_241,N_9962,N_9901);
or UO_242 (O_242,N_9999,N_9952);
and UO_243 (O_243,N_9913,N_9995);
nor UO_244 (O_244,N_9951,N_9906);
or UO_245 (O_245,N_9903,N_9925);
nor UO_246 (O_246,N_9917,N_9915);
nor UO_247 (O_247,N_9928,N_9911);
and UO_248 (O_248,N_9914,N_9974);
nand UO_249 (O_249,N_9918,N_9945);
nor UO_250 (O_250,N_9925,N_9904);
xnor UO_251 (O_251,N_9972,N_9944);
and UO_252 (O_252,N_9909,N_9985);
or UO_253 (O_253,N_9907,N_9946);
nand UO_254 (O_254,N_9942,N_9938);
or UO_255 (O_255,N_9968,N_9930);
or UO_256 (O_256,N_9966,N_9994);
and UO_257 (O_257,N_9981,N_9974);
and UO_258 (O_258,N_9914,N_9989);
nor UO_259 (O_259,N_9905,N_9913);
and UO_260 (O_260,N_9914,N_9913);
nand UO_261 (O_261,N_9991,N_9942);
and UO_262 (O_262,N_9954,N_9936);
nor UO_263 (O_263,N_9975,N_9919);
and UO_264 (O_264,N_9907,N_9908);
nor UO_265 (O_265,N_9940,N_9919);
xor UO_266 (O_266,N_9942,N_9931);
nand UO_267 (O_267,N_9955,N_9910);
and UO_268 (O_268,N_9938,N_9994);
nand UO_269 (O_269,N_9977,N_9901);
nor UO_270 (O_270,N_9985,N_9914);
xor UO_271 (O_271,N_9964,N_9955);
nand UO_272 (O_272,N_9923,N_9996);
and UO_273 (O_273,N_9919,N_9961);
and UO_274 (O_274,N_9952,N_9939);
nor UO_275 (O_275,N_9918,N_9916);
xor UO_276 (O_276,N_9929,N_9976);
or UO_277 (O_277,N_9972,N_9955);
xnor UO_278 (O_278,N_9935,N_9929);
nand UO_279 (O_279,N_9989,N_9961);
nor UO_280 (O_280,N_9997,N_9938);
or UO_281 (O_281,N_9972,N_9927);
or UO_282 (O_282,N_9912,N_9999);
and UO_283 (O_283,N_9919,N_9947);
and UO_284 (O_284,N_9987,N_9999);
nand UO_285 (O_285,N_9983,N_9968);
nand UO_286 (O_286,N_9999,N_9963);
nor UO_287 (O_287,N_9986,N_9968);
and UO_288 (O_288,N_9914,N_9955);
nor UO_289 (O_289,N_9924,N_9937);
and UO_290 (O_290,N_9959,N_9979);
nand UO_291 (O_291,N_9902,N_9935);
and UO_292 (O_292,N_9971,N_9922);
or UO_293 (O_293,N_9912,N_9932);
xnor UO_294 (O_294,N_9958,N_9936);
nand UO_295 (O_295,N_9951,N_9978);
xor UO_296 (O_296,N_9942,N_9998);
or UO_297 (O_297,N_9949,N_9986);
nand UO_298 (O_298,N_9941,N_9925);
nor UO_299 (O_299,N_9908,N_9989);
nor UO_300 (O_300,N_9932,N_9972);
nor UO_301 (O_301,N_9939,N_9922);
or UO_302 (O_302,N_9986,N_9988);
nand UO_303 (O_303,N_9951,N_9971);
and UO_304 (O_304,N_9956,N_9945);
and UO_305 (O_305,N_9966,N_9985);
nor UO_306 (O_306,N_9916,N_9954);
nand UO_307 (O_307,N_9946,N_9914);
nor UO_308 (O_308,N_9937,N_9902);
and UO_309 (O_309,N_9908,N_9956);
or UO_310 (O_310,N_9969,N_9974);
nor UO_311 (O_311,N_9903,N_9974);
nor UO_312 (O_312,N_9977,N_9990);
and UO_313 (O_313,N_9990,N_9966);
nor UO_314 (O_314,N_9969,N_9949);
or UO_315 (O_315,N_9953,N_9934);
nand UO_316 (O_316,N_9945,N_9998);
nor UO_317 (O_317,N_9916,N_9923);
nor UO_318 (O_318,N_9923,N_9930);
nand UO_319 (O_319,N_9917,N_9920);
nor UO_320 (O_320,N_9996,N_9973);
or UO_321 (O_321,N_9924,N_9902);
nand UO_322 (O_322,N_9955,N_9909);
and UO_323 (O_323,N_9988,N_9987);
nand UO_324 (O_324,N_9962,N_9980);
nand UO_325 (O_325,N_9986,N_9904);
or UO_326 (O_326,N_9937,N_9913);
or UO_327 (O_327,N_9950,N_9979);
or UO_328 (O_328,N_9951,N_9910);
nor UO_329 (O_329,N_9961,N_9948);
or UO_330 (O_330,N_9980,N_9923);
and UO_331 (O_331,N_9936,N_9911);
and UO_332 (O_332,N_9993,N_9931);
nand UO_333 (O_333,N_9976,N_9958);
nand UO_334 (O_334,N_9963,N_9913);
and UO_335 (O_335,N_9958,N_9907);
nand UO_336 (O_336,N_9977,N_9966);
and UO_337 (O_337,N_9970,N_9901);
nand UO_338 (O_338,N_9954,N_9968);
or UO_339 (O_339,N_9987,N_9950);
nor UO_340 (O_340,N_9968,N_9920);
and UO_341 (O_341,N_9969,N_9970);
nand UO_342 (O_342,N_9988,N_9962);
nor UO_343 (O_343,N_9950,N_9980);
xnor UO_344 (O_344,N_9978,N_9940);
xnor UO_345 (O_345,N_9923,N_9941);
xor UO_346 (O_346,N_9975,N_9962);
nor UO_347 (O_347,N_9906,N_9981);
nor UO_348 (O_348,N_9915,N_9901);
nand UO_349 (O_349,N_9987,N_9923);
xnor UO_350 (O_350,N_9999,N_9989);
or UO_351 (O_351,N_9952,N_9955);
nand UO_352 (O_352,N_9964,N_9983);
and UO_353 (O_353,N_9980,N_9987);
and UO_354 (O_354,N_9994,N_9920);
xor UO_355 (O_355,N_9948,N_9969);
and UO_356 (O_356,N_9919,N_9906);
and UO_357 (O_357,N_9998,N_9930);
and UO_358 (O_358,N_9997,N_9915);
and UO_359 (O_359,N_9966,N_9962);
nor UO_360 (O_360,N_9965,N_9984);
and UO_361 (O_361,N_9926,N_9954);
or UO_362 (O_362,N_9927,N_9921);
nand UO_363 (O_363,N_9961,N_9953);
nand UO_364 (O_364,N_9952,N_9922);
nand UO_365 (O_365,N_9950,N_9969);
or UO_366 (O_366,N_9977,N_9938);
and UO_367 (O_367,N_9982,N_9924);
nor UO_368 (O_368,N_9972,N_9938);
nand UO_369 (O_369,N_9920,N_9954);
xor UO_370 (O_370,N_9907,N_9934);
nand UO_371 (O_371,N_9948,N_9968);
nand UO_372 (O_372,N_9931,N_9985);
nand UO_373 (O_373,N_9966,N_9993);
nand UO_374 (O_374,N_9974,N_9927);
nor UO_375 (O_375,N_9900,N_9961);
xnor UO_376 (O_376,N_9932,N_9926);
and UO_377 (O_377,N_9902,N_9989);
and UO_378 (O_378,N_9900,N_9957);
and UO_379 (O_379,N_9916,N_9974);
nor UO_380 (O_380,N_9935,N_9949);
nand UO_381 (O_381,N_9937,N_9975);
xor UO_382 (O_382,N_9942,N_9969);
nor UO_383 (O_383,N_9989,N_9957);
nand UO_384 (O_384,N_9901,N_9936);
nand UO_385 (O_385,N_9979,N_9996);
or UO_386 (O_386,N_9904,N_9993);
or UO_387 (O_387,N_9926,N_9994);
or UO_388 (O_388,N_9924,N_9988);
nand UO_389 (O_389,N_9994,N_9964);
nor UO_390 (O_390,N_9908,N_9996);
or UO_391 (O_391,N_9906,N_9907);
nor UO_392 (O_392,N_9994,N_9932);
nand UO_393 (O_393,N_9936,N_9950);
or UO_394 (O_394,N_9959,N_9952);
nand UO_395 (O_395,N_9925,N_9980);
and UO_396 (O_396,N_9935,N_9930);
nor UO_397 (O_397,N_9928,N_9945);
or UO_398 (O_398,N_9961,N_9917);
nor UO_399 (O_399,N_9944,N_9984);
nor UO_400 (O_400,N_9922,N_9962);
nand UO_401 (O_401,N_9956,N_9935);
and UO_402 (O_402,N_9912,N_9973);
xnor UO_403 (O_403,N_9920,N_9923);
or UO_404 (O_404,N_9901,N_9994);
nor UO_405 (O_405,N_9935,N_9968);
nand UO_406 (O_406,N_9981,N_9948);
nor UO_407 (O_407,N_9956,N_9944);
nor UO_408 (O_408,N_9997,N_9950);
or UO_409 (O_409,N_9950,N_9934);
nor UO_410 (O_410,N_9908,N_9998);
or UO_411 (O_411,N_9980,N_9969);
nand UO_412 (O_412,N_9929,N_9964);
nor UO_413 (O_413,N_9911,N_9944);
or UO_414 (O_414,N_9990,N_9911);
nor UO_415 (O_415,N_9976,N_9924);
xnor UO_416 (O_416,N_9928,N_9997);
and UO_417 (O_417,N_9969,N_9994);
or UO_418 (O_418,N_9935,N_9967);
or UO_419 (O_419,N_9949,N_9917);
nand UO_420 (O_420,N_9952,N_9954);
nor UO_421 (O_421,N_9942,N_9993);
nand UO_422 (O_422,N_9973,N_9977);
nand UO_423 (O_423,N_9999,N_9927);
and UO_424 (O_424,N_9987,N_9919);
or UO_425 (O_425,N_9976,N_9935);
or UO_426 (O_426,N_9999,N_9957);
nand UO_427 (O_427,N_9950,N_9935);
or UO_428 (O_428,N_9995,N_9999);
nor UO_429 (O_429,N_9905,N_9996);
xor UO_430 (O_430,N_9969,N_9911);
nor UO_431 (O_431,N_9968,N_9961);
nor UO_432 (O_432,N_9924,N_9955);
and UO_433 (O_433,N_9992,N_9913);
nand UO_434 (O_434,N_9971,N_9973);
nor UO_435 (O_435,N_9953,N_9996);
or UO_436 (O_436,N_9927,N_9966);
and UO_437 (O_437,N_9940,N_9922);
nand UO_438 (O_438,N_9946,N_9972);
xnor UO_439 (O_439,N_9995,N_9944);
and UO_440 (O_440,N_9906,N_9987);
nand UO_441 (O_441,N_9966,N_9963);
nand UO_442 (O_442,N_9990,N_9949);
and UO_443 (O_443,N_9979,N_9999);
and UO_444 (O_444,N_9917,N_9946);
nor UO_445 (O_445,N_9951,N_9925);
and UO_446 (O_446,N_9932,N_9931);
or UO_447 (O_447,N_9919,N_9979);
nor UO_448 (O_448,N_9929,N_9984);
xnor UO_449 (O_449,N_9945,N_9977);
nand UO_450 (O_450,N_9920,N_9905);
or UO_451 (O_451,N_9980,N_9910);
and UO_452 (O_452,N_9954,N_9908);
or UO_453 (O_453,N_9950,N_9971);
or UO_454 (O_454,N_9963,N_9964);
nand UO_455 (O_455,N_9984,N_9986);
and UO_456 (O_456,N_9938,N_9915);
or UO_457 (O_457,N_9943,N_9912);
xnor UO_458 (O_458,N_9970,N_9953);
xnor UO_459 (O_459,N_9929,N_9994);
nor UO_460 (O_460,N_9989,N_9928);
xnor UO_461 (O_461,N_9971,N_9938);
nor UO_462 (O_462,N_9999,N_9911);
or UO_463 (O_463,N_9961,N_9954);
and UO_464 (O_464,N_9919,N_9950);
nand UO_465 (O_465,N_9967,N_9934);
nand UO_466 (O_466,N_9934,N_9964);
nor UO_467 (O_467,N_9990,N_9972);
and UO_468 (O_468,N_9999,N_9905);
nand UO_469 (O_469,N_9949,N_9918);
or UO_470 (O_470,N_9985,N_9957);
nor UO_471 (O_471,N_9973,N_9950);
nor UO_472 (O_472,N_9957,N_9921);
nand UO_473 (O_473,N_9938,N_9999);
nand UO_474 (O_474,N_9910,N_9944);
nor UO_475 (O_475,N_9936,N_9934);
and UO_476 (O_476,N_9901,N_9944);
nand UO_477 (O_477,N_9935,N_9900);
and UO_478 (O_478,N_9935,N_9957);
nand UO_479 (O_479,N_9993,N_9974);
or UO_480 (O_480,N_9936,N_9937);
and UO_481 (O_481,N_9938,N_9949);
or UO_482 (O_482,N_9900,N_9970);
xor UO_483 (O_483,N_9947,N_9912);
nand UO_484 (O_484,N_9970,N_9911);
nand UO_485 (O_485,N_9935,N_9928);
and UO_486 (O_486,N_9995,N_9967);
and UO_487 (O_487,N_9958,N_9966);
nor UO_488 (O_488,N_9928,N_9944);
nor UO_489 (O_489,N_9965,N_9980);
or UO_490 (O_490,N_9958,N_9948);
and UO_491 (O_491,N_9946,N_9921);
xor UO_492 (O_492,N_9954,N_9921);
nor UO_493 (O_493,N_9901,N_9964);
and UO_494 (O_494,N_9959,N_9931);
and UO_495 (O_495,N_9923,N_9971);
or UO_496 (O_496,N_9923,N_9925);
nand UO_497 (O_497,N_9909,N_9946);
and UO_498 (O_498,N_9976,N_9961);
and UO_499 (O_499,N_9910,N_9978);
nand UO_500 (O_500,N_9929,N_9907);
and UO_501 (O_501,N_9926,N_9906);
or UO_502 (O_502,N_9979,N_9932);
nand UO_503 (O_503,N_9945,N_9903);
and UO_504 (O_504,N_9902,N_9927);
nand UO_505 (O_505,N_9963,N_9947);
xnor UO_506 (O_506,N_9998,N_9975);
nor UO_507 (O_507,N_9956,N_9909);
nand UO_508 (O_508,N_9943,N_9975);
and UO_509 (O_509,N_9981,N_9965);
nand UO_510 (O_510,N_9949,N_9906);
or UO_511 (O_511,N_9919,N_9993);
or UO_512 (O_512,N_9913,N_9996);
xor UO_513 (O_513,N_9947,N_9998);
and UO_514 (O_514,N_9982,N_9900);
and UO_515 (O_515,N_9967,N_9960);
nor UO_516 (O_516,N_9965,N_9986);
or UO_517 (O_517,N_9951,N_9924);
nand UO_518 (O_518,N_9906,N_9914);
nand UO_519 (O_519,N_9917,N_9978);
and UO_520 (O_520,N_9911,N_9916);
nor UO_521 (O_521,N_9992,N_9993);
xnor UO_522 (O_522,N_9954,N_9963);
nand UO_523 (O_523,N_9912,N_9966);
nand UO_524 (O_524,N_9936,N_9978);
and UO_525 (O_525,N_9905,N_9991);
and UO_526 (O_526,N_9931,N_9958);
nand UO_527 (O_527,N_9932,N_9951);
xor UO_528 (O_528,N_9934,N_9941);
or UO_529 (O_529,N_9978,N_9987);
or UO_530 (O_530,N_9901,N_9931);
or UO_531 (O_531,N_9962,N_9973);
and UO_532 (O_532,N_9963,N_9952);
xnor UO_533 (O_533,N_9950,N_9930);
and UO_534 (O_534,N_9958,N_9994);
nand UO_535 (O_535,N_9993,N_9988);
or UO_536 (O_536,N_9994,N_9952);
nor UO_537 (O_537,N_9922,N_9913);
nor UO_538 (O_538,N_9949,N_9958);
and UO_539 (O_539,N_9909,N_9969);
nor UO_540 (O_540,N_9943,N_9906);
nand UO_541 (O_541,N_9957,N_9918);
or UO_542 (O_542,N_9981,N_9995);
xor UO_543 (O_543,N_9962,N_9993);
nor UO_544 (O_544,N_9939,N_9925);
and UO_545 (O_545,N_9918,N_9910);
nor UO_546 (O_546,N_9981,N_9977);
or UO_547 (O_547,N_9938,N_9903);
and UO_548 (O_548,N_9992,N_9963);
nor UO_549 (O_549,N_9999,N_9903);
or UO_550 (O_550,N_9930,N_9909);
and UO_551 (O_551,N_9933,N_9973);
or UO_552 (O_552,N_9998,N_9915);
or UO_553 (O_553,N_9969,N_9985);
nand UO_554 (O_554,N_9951,N_9992);
or UO_555 (O_555,N_9933,N_9916);
nor UO_556 (O_556,N_9971,N_9911);
or UO_557 (O_557,N_9939,N_9975);
nor UO_558 (O_558,N_9977,N_9996);
xor UO_559 (O_559,N_9974,N_9954);
nand UO_560 (O_560,N_9970,N_9991);
nor UO_561 (O_561,N_9996,N_9949);
or UO_562 (O_562,N_9985,N_9903);
nand UO_563 (O_563,N_9934,N_9956);
nor UO_564 (O_564,N_9976,N_9926);
or UO_565 (O_565,N_9997,N_9907);
nand UO_566 (O_566,N_9901,N_9933);
or UO_567 (O_567,N_9981,N_9983);
and UO_568 (O_568,N_9976,N_9903);
and UO_569 (O_569,N_9941,N_9939);
or UO_570 (O_570,N_9932,N_9988);
nor UO_571 (O_571,N_9997,N_9974);
or UO_572 (O_572,N_9944,N_9932);
nand UO_573 (O_573,N_9910,N_9990);
and UO_574 (O_574,N_9965,N_9937);
nor UO_575 (O_575,N_9961,N_9921);
nand UO_576 (O_576,N_9990,N_9930);
nor UO_577 (O_577,N_9905,N_9933);
nand UO_578 (O_578,N_9910,N_9957);
or UO_579 (O_579,N_9990,N_9901);
nand UO_580 (O_580,N_9973,N_9908);
nand UO_581 (O_581,N_9916,N_9906);
nand UO_582 (O_582,N_9979,N_9986);
nor UO_583 (O_583,N_9932,N_9953);
nor UO_584 (O_584,N_9940,N_9948);
or UO_585 (O_585,N_9901,N_9991);
nor UO_586 (O_586,N_9950,N_9981);
nand UO_587 (O_587,N_9986,N_9912);
nand UO_588 (O_588,N_9900,N_9943);
nand UO_589 (O_589,N_9930,N_9949);
and UO_590 (O_590,N_9902,N_9969);
or UO_591 (O_591,N_9915,N_9933);
or UO_592 (O_592,N_9948,N_9943);
and UO_593 (O_593,N_9945,N_9985);
and UO_594 (O_594,N_9981,N_9962);
or UO_595 (O_595,N_9933,N_9922);
and UO_596 (O_596,N_9943,N_9905);
or UO_597 (O_597,N_9903,N_9930);
and UO_598 (O_598,N_9985,N_9995);
nand UO_599 (O_599,N_9920,N_9980);
nand UO_600 (O_600,N_9902,N_9982);
and UO_601 (O_601,N_9980,N_9932);
and UO_602 (O_602,N_9914,N_9952);
and UO_603 (O_603,N_9968,N_9913);
nor UO_604 (O_604,N_9912,N_9951);
or UO_605 (O_605,N_9905,N_9941);
or UO_606 (O_606,N_9921,N_9958);
or UO_607 (O_607,N_9996,N_9924);
xnor UO_608 (O_608,N_9968,N_9990);
or UO_609 (O_609,N_9913,N_9961);
and UO_610 (O_610,N_9946,N_9916);
and UO_611 (O_611,N_9952,N_9996);
or UO_612 (O_612,N_9925,N_9944);
nor UO_613 (O_613,N_9945,N_9952);
nor UO_614 (O_614,N_9957,N_9942);
xor UO_615 (O_615,N_9989,N_9965);
nand UO_616 (O_616,N_9955,N_9987);
and UO_617 (O_617,N_9930,N_9948);
nand UO_618 (O_618,N_9967,N_9912);
nor UO_619 (O_619,N_9968,N_9982);
and UO_620 (O_620,N_9940,N_9993);
nand UO_621 (O_621,N_9976,N_9947);
nor UO_622 (O_622,N_9906,N_9958);
xnor UO_623 (O_623,N_9969,N_9957);
nor UO_624 (O_624,N_9902,N_9911);
nor UO_625 (O_625,N_9948,N_9956);
and UO_626 (O_626,N_9953,N_9999);
or UO_627 (O_627,N_9923,N_9959);
nor UO_628 (O_628,N_9989,N_9919);
and UO_629 (O_629,N_9921,N_9917);
nor UO_630 (O_630,N_9977,N_9947);
nor UO_631 (O_631,N_9963,N_9958);
or UO_632 (O_632,N_9970,N_9915);
xor UO_633 (O_633,N_9934,N_9900);
nor UO_634 (O_634,N_9925,N_9979);
xnor UO_635 (O_635,N_9946,N_9955);
nor UO_636 (O_636,N_9954,N_9995);
xor UO_637 (O_637,N_9981,N_9970);
nand UO_638 (O_638,N_9945,N_9936);
nor UO_639 (O_639,N_9989,N_9955);
or UO_640 (O_640,N_9924,N_9978);
and UO_641 (O_641,N_9986,N_9962);
or UO_642 (O_642,N_9994,N_9907);
nor UO_643 (O_643,N_9943,N_9901);
or UO_644 (O_644,N_9910,N_9942);
nor UO_645 (O_645,N_9984,N_9937);
xor UO_646 (O_646,N_9955,N_9968);
or UO_647 (O_647,N_9996,N_9985);
nand UO_648 (O_648,N_9958,N_9988);
nand UO_649 (O_649,N_9924,N_9935);
and UO_650 (O_650,N_9982,N_9945);
nand UO_651 (O_651,N_9946,N_9977);
or UO_652 (O_652,N_9974,N_9940);
or UO_653 (O_653,N_9915,N_9995);
xnor UO_654 (O_654,N_9932,N_9995);
xnor UO_655 (O_655,N_9941,N_9995);
and UO_656 (O_656,N_9948,N_9944);
xor UO_657 (O_657,N_9907,N_9973);
or UO_658 (O_658,N_9986,N_9956);
nor UO_659 (O_659,N_9931,N_9976);
nor UO_660 (O_660,N_9991,N_9963);
nand UO_661 (O_661,N_9982,N_9929);
or UO_662 (O_662,N_9910,N_9983);
xor UO_663 (O_663,N_9982,N_9961);
nand UO_664 (O_664,N_9923,N_9965);
xor UO_665 (O_665,N_9972,N_9949);
nand UO_666 (O_666,N_9989,N_9938);
or UO_667 (O_667,N_9986,N_9995);
nor UO_668 (O_668,N_9965,N_9954);
nor UO_669 (O_669,N_9911,N_9905);
nand UO_670 (O_670,N_9947,N_9983);
nor UO_671 (O_671,N_9905,N_9987);
and UO_672 (O_672,N_9948,N_9910);
nor UO_673 (O_673,N_9936,N_9914);
and UO_674 (O_674,N_9914,N_9995);
or UO_675 (O_675,N_9980,N_9947);
nor UO_676 (O_676,N_9986,N_9911);
nor UO_677 (O_677,N_9934,N_9966);
and UO_678 (O_678,N_9984,N_9933);
and UO_679 (O_679,N_9907,N_9959);
and UO_680 (O_680,N_9991,N_9949);
nor UO_681 (O_681,N_9978,N_9999);
or UO_682 (O_682,N_9965,N_9946);
and UO_683 (O_683,N_9941,N_9967);
and UO_684 (O_684,N_9959,N_9992);
or UO_685 (O_685,N_9996,N_9955);
nor UO_686 (O_686,N_9901,N_9948);
or UO_687 (O_687,N_9984,N_9953);
nand UO_688 (O_688,N_9961,N_9947);
or UO_689 (O_689,N_9908,N_9922);
nand UO_690 (O_690,N_9922,N_9996);
and UO_691 (O_691,N_9992,N_9938);
and UO_692 (O_692,N_9948,N_9904);
or UO_693 (O_693,N_9987,N_9903);
nand UO_694 (O_694,N_9914,N_9986);
nor UO_695 (O_695,N_9931,N_9909);
or UO_696 (O_696,N_9934,N_9960);
and UO_697 (O_697,N_9930,N_9938);
or UO_698 (O_698,N_9952,N_9923);
nor UO_699 (O_699,N_9997,N_9996);
nand UO_700 (O_700,N_9943,N_9953);
nand UO_701 (O_701,N_9936,N_9995);
or UO_702 (O_702,N_9960,N_9918);
and UO_703 (O_703,N_9918,N_9970);
nor UO_704 (O_704,N_9962,N_9947);
xnor UO_705 (O_705,N_9930,N_9957);
nor UO_706 (O_706,N_9941,N_9957);
nand UO_707 (O_707,N_9951,N_9973);
nand UO_708 (O_708,N_9943,N_9982);
nor UO_709 (O_709,N_9977,N_9962);
xor UO_710 (O_710,N_9958,N_9964);
nand UO_711 (O_711,N_9922,N_9993);
and UO_712 (O_712,N_9925,N_9918);
or UO_713 (O_713,N_9985,N_9924);
xnor UO_714 (O_714,N_9963,N_9957);
or UO_715 (O_715,N_9965,N_9903);
nand UO_716 (O_716,N_9914,N_9950);
or UO_717 (O_717,N_9963,N_9974);
or UO_718 (O_718,N_9971,N_9926);
nor UO_719 (O_719,N_9917,N_9957);
xnor UO_720 (O_720,N_9917,N_9922);
or UO_721 (O_721,N_9902,N_9936);
nand UO_722 (O_722,N_9910,N_9915);
nor UO_723 (O_723,N_9984,N_9945);
nor UO_724 (O_724,N_9982,N_9999);
nor UO_725 (O_725,N_9934,N_9984);
nand UO_726 (O_726,N_9967,N_9940);
nor UO_727 (O_727,N_9900,N_9921);
nor UO_728 (O_728,N_9998,N_9963);
or UO_729 (O_729,N_9950,N_9975);
and UO_730 (O_730,N_9959,N_9918);
nand UO_731 (O_731,N_9986,N_9916);
nand UO_732 (O_732,N_9962,N_9939);
or UO_733 (O_733,N_9968,N_9985);
nor UO_734 (O_734,N_9917,N_9934);
and UO_735 (O_735,N_9993,N_9990);
nand UO_736 (O_736,N_9912,N_9992);
xnor UO_737 (O_737,N_9956,N_9919);
or UO_738 (O_738,N_9954,N_9992);
and UO_739 (O_739,N_9983,N_9980);
or UO_740 (O_740,N_9915,N_9937);
nand UO_741 (O_741,N_9920,N_9930);
or UO_742 (O_742,N_9929,N_9942);
nor UO_743 (O_743,N_9979,N_9931);
and UO_744 (O_744,N_9947,N_9975);
and UO_745 (O_745,N_9933,N_9978);
nor UO_746 (O_746,N_9964,N_9974);
nand UO_747 (O_747,N_9975,N_9993);
nor UO_748 (O_748,N_9974,N_9956);
and UO_749 (O_749,N_9918,N_9963);
xor UO_750 (O_750,N_9912,N_9900);
or UO_751 (O_751,N_9938,N_9924);
xor UO_752 (O_752,N_9928,N_9979);
nand UO_753 (O_753,N_9937,N_9953);
nor UO_754 (O_754,N_9928,N_9947);
and UO_755 (O_755,N_9961,N_9995);
nor UO_756 (O_756,N_9990,N_9970);
nand UO_757 (O_757,N_9951,N_9975);
and UO_758 (O_758,N_9944,N_9974);
and UO_759 (O_759,N_9982,N_9930);
nand UO_760 (O_760,N_9940,N_9952);
xnor UO_761 (O_761,N_9910,N_9977);
nand UO_762 (O_762,N_9939,N_9936);
nand UO_763 (O_763,N_9933,N_9925);
nand UO_764 (O_764,N_9948,N_9962);
and UO_765 (O_765,N_9981,N_9980);
or UO_766 (O_766,N_9918,N_9952);
nand UO_767 (O_767,N_9965,N_9901);
or UO_768 (O_768,N_9986,N_9940);
xnor UO_769 (O_769,N_9904,N_9950);
or UO_770 (O_770,N_9932,N_9908);
nor UO_771 (O_771,N_9945,N_9989);
nor UO_772 (O_772,N_9908,N_9993);
nor UO_773 (O_773,N_9912,N_9946);
and UO_774 (O_774,N_9942,N_9971);
or UO_775 (O_775,N_9917,N_9955);
nor UO_776 (O_776,N_9903,N_9919);
and UO_777 (O_777,N_9924,N_9986);
nand UO_778 (O_778,N_9918,N_9922);
nand UO_779 (O_779,N_9980,N_9978);
nand UO_780 (O_780,N_9989,N_9909);
or UO_781 (O_781,N_9911,N_9972);
and UO_782 (O_782,N_9939,N_9993);
or UO_783 (O_783,N_9923,N_9940);
nor UO_784 (O_784,N_9973,N_9988);
nand UO_785 (O_785,N_9983,N_9998);
xnor UO_786 (O_786,N_9993,N_9915);
nor UO_787 (O_787,N_9937,N_9903);
nand UO_788 (O_788,N_9980,N_9913);
or UO_789 (O_789,N_9956,N_9926);
nor UO_790 (O_790,N_9954,N_9944);
and UO_791 (O_791,N_9995,N_9980);
xor UO_792 (O_792,N_9932,N_9903);
nor UO_793 (O_793,N_9997,N_9929);
and UO_794 (O_794,N_9945,N_9931);
and UO_795 (O_795,N_9932,N_9990);
nand UO_796 (O_796,N_9944,N_9964);
and UO_797 (O_797,N_9963,N_9904);
or UO_798 (O_798,N_9966,N_9979);
nand UO_799 (O_799,N_9979,N_9935);
nand UO_800 (O_800,N_9902,N_9999);
nor UO_801 (O_801,N_9911,N_9904);
nand UO_802 (O_802,N_9984,N_9995);
and UO_803 (O_803,N_9923,N_9948);
or UO_804 (O_804,N_9916,N_9928);
nand UO_805 (O_805,N_9909,N_9959);
nor UO_806 (O_806,N_9913,N_9990);
nor UO_807 (O_807,N_9949,N_9961);
and UO_808 (O_808,N_9947,N_9941);
nor UO_809 (O_809,N_9911,N_9996);
xor UO_810 (O_810,N_9977,N_9937);
and UO_811 (O_811,N_9945,N_9909);
nor UO_812 (O_812,N_9957,N_9920);
or UO_813 (O_813,N_9999,N_9935);
nor UO_814 (O_814,N_9944,N_9946);
nand UO_815 (O_815,N_9930,N_9940);
nand UO_816 (O_816,N_9913,N_9966);
nor UO_817 (O_817,N_9947,N_9913);
nor UO_818 (O_818,N_9987,N_9998);
and UO_819 (O_819,N_9935,N_9943);
nand UO_820 (O_820,N_9925,N_9968);
or UO_821 (O_821,N_9965,N_9935);
or UO_822 (O_822,N_9949,N_9989);
or UO_823 (O_823,N_9952,N_9978);
xor UO_824 (O_824,N_9902,N_9930);
xor UO_825 (O_825,N_9993,N_9946);
or UO_826 (O_826,N_9984,N_9927);
and UO_827 (O_827,N_9945,N_9972);
nor UO_828 (O_828,N_9991,N_9980);
and UO_829 (O_829,N_9996,N_9970);
or UO_830 (O_830,N_9918,N_9912);
xnor UO_831 (O_831,N_9947,N_9927);
xnor UO_832 (O_832,N_9903,N_9936);
or UO_833 (O_833,N_9948,N_9977);
nor UO_834 (O_834,N_9951,N_9915);
or UO_835 (O_835,N_9912,N_9976);
nand UO_836 (O_836,N_9987,N_9929);
nor UO_837 (O_837,N_9945,N_9924);
or UO_838 (O_838,N_9912,N_9944);
or UO_839 (O_839,N_9906,N_9913);
xnor UO_840 (O_840,N_9926,N_9931);
or UO_841 (O_841,N_9957,N_9927);
and UO_842 (O_842,N_9941,N_9951);
nor UO_843 (O_843,N_9978,N_9944);
nor UO_844 (O_844,N_9952,N_9927);
or UO_845 (O_845,N_9977,N_9915);
nor UO_846 (O_846,N_9914,N_9983);
and UO_847 (O_847,N_9960,N_9901);
nor UO_848 (O_848,N_9901,N_9951);
nand UO_849 (O_849,N_9982,N_9910);
and UO_850 (O_850,N_9921,N_9959);
and UO_851 (O_851,N_9933,N_9985);
and UO_852 (O_852,N_9956,N_9950);
xnor UO_853 (O_853,N_9998,N_9938);
xnor UO_854 (O_854,N_9928,N_9982);
and UO_855 (O_855,N_9914,N_9941);
nor UO_856 (O_856,N_9938,N_9964);
xnor UO_857 (O_857,N_9914,N_9971);
nand UO_858 (O_858,N_9947,N_9953);
nor UO_859 (O_859,N_9995,N_9949);
nor UO_860 (O_860,N_9921,N_9964);
or UO_861 (O_861,N_9914,N_9978);
nand UO_862 (O_862,N_9976,N_9979);
or UO_863 (O_863,N_9965,N_9969);
or UO_864 (O_864,N_9997,N_9941);
nand UO_865 (O_865,N_9974,N_9902);
and UO_866 (O_866,N_9904,N_9981);
nand UO_867 (O_867,N_9901,N_9918);
or UO_868 (O_868,N_9918,N_9936);
nor UO_869 (O_869,N_9990,N_9919);
and UO_870 (O_870,N_9984,N_9960);
and UO_871 (O_871,N_9913,N_9939);
or UO_872 (O_872,N_9977,N_9942);
xor UO_873 (O_873,N_9938,N_9995);
nor UO_874 (O_874,N_9915,N_9979);
and UO_875 (O_875,N_9950,N_9932);
xor UO_876 (O_876,N_9949,N_9981);
nor UO_877 (O_877,N_9954,N_9909);
and UO_878 (O_878,N_9944,N_9933);
nand UO_879 (O_879,N_9912,N_9911);
nand UO_880 (O_880,N_9954,N_9989);
xor UO_881 (O_881,N_9992,N_9945);
or UO_882 (O_882,N_9959,N_9953);
xor UO_883 (O_883,N_9976,N_9970);
xor UO_884 (O_884,N_9983,N_9937);
xor UO_885 (O_885,N_9968,N_9997);
xor UO_886 (O_886,N_9961,N_9992);
nor UO_887 (O_887,N_9936,N_9916);
nor UO_888 (O_888,N_9959,N_9956);
nand UO_889 (O_889,N_9986,N_9985);
and UO_890 (O_890,N_9980,N_9976);
or UO_891 (O_891,N_9976,N_9953);
nand UO_892 (O_892,N_9932,N_9966);
and UO_893 (O_893,N_9940,N_9911);
nand UO_894 (O_894,N_9938,N_9929);
nor UO_895 (O_895,N_9989,N_9930);
and UO_896 (O_896,N_9904,N_9987);
nand UO_897 (O_897,N_9943,N_9916);
and UO_898 (O_898,N_9916,N_9989);
nor UO_899 (O_899,N_9991,N_9912);
nand UO_900 (O_900,N_9927,N_9916);
or UO_901 (O_901,N_9976,N_9919);
nand UO_902 (O_902,N_9909,N_9953);
nor UO_903 (O_903,N_9972,N_9979);
or UO_904 (O_904,N_9918,N_9958);
or UO_905 (O_905,N_9962,N_9946);
or UO_906 (O_906,N_9917,N_9966);
nor UO_907 (O_907,N_9959,N_9943);
or UO_908 (O_908,N_9961,N_9941);
or UO_909 (O_909,N_9961,N_9971);
and UO_910 (O_910,N_9927,N_9943);
nand UO_911 (O_911,N_9942,N_9924);
nand UO_912 (O_912,N_9930,N_9942);
nand UO_913 (O_913,N_9902,N_9962);
nand UO_914 (O_914,N_9926,N_9999);
nor UO_915 (O_915,N_9922,N_9970);
nor UO_916 (O_916,N_9986,N_9957);
nor UO_917 (O_917,N_9905,N_9960);
nor UO_918 (O_918,N_9936,N_9953);
xnor UO_919 (O_919,N_9904,N_9951);
and UO_920 (O_920,N_9925,N_9942);
or UO_921 (O_921,N_9975,N_9989);
and UO_922 (O_922,N_9911,N_9963);
nand UO_923 (O_923,N_9995,N_9973);
nand UO_924 (O_924,N_9958,N_9939);
nor UO_925 (O_925,N_9997,N_9906);
or UO_926 (O_926,N_9935,N_9948);
and UO_927 (O_927,N_9973,N_9989);
or UO_928 (O_928,N_9934,N_9992);
or UO_929 (O_929,N_9942,N_9939);
and UO_930 (O_930,N_9952,N_9936);
xnor UO_931 (O_931,N_9997,N_9924);
nor UO_932 (O_932,N_9981,N_9914);
nor UO_933 (O_933,N_9913,N_9940);
nand UO_934 (O_934,N_9942,N_9956);
nand UO_935 (O_935,N_9944,N_9962);
and UO_936 (O_936,N_9997,N_9954);
and UO_937 (O_937,N_9991,N_9931);
or UO_938 (O_938,N_9992,N_9928);
nor UO_939 (O_939,N_9968,N_9906);
or UO_940 (O_940,N_9961,N_9940);
xor UO_941 (O_941,N_9939,N_9902);
or UO_942 (O_942,N_9933,N_9920);
nor UO_943 (O_943,N_9968,N_9950);
or UO_944 (O_944,N_9911,N_9973);
nand UO_945 (O_945,N_9933,N_9940);
and UO_946 (O_946,N_9975,N_9954);
nand UO_947 (O_947,N_9941,N_9919);
nor UO_948 (O_948,N_9923,N_9985);
nand UO_949 (O_949,N_9929,N_9992);
and UO_950 (O_950,N_9937,N_9963);
or UO_951 (O_951,N_9921,N_9968);
nand UO_952 (O_952,N_9988,N_9997);
xnor UO_953 (O_953,N_9942,N_9944);
xor UO_954 (O_954,N_9967,N_9933);
xor UO_955 (O_955,N_9920,N_9999);
and UO_956 (O_956,N_9960,N_9956);
nand UO_957 (O_957,N_9955,N_9941);
nor UO_958 (O_958,N_9935,N_9981);
or UO_959 (O_959,N_9971,N_9972);
nand UO_960 (O_960,N_9967,N_9919);
nand UO_961 (O_961,N_9988,N_9916);
nor UO_962 (O_962,N_9998,N_9924);
or UO_963 (O_963,N_9953,N_9956);
and UO_964 (O_964,N_9940,N_9920);
or UO_965 (O_965,N_9907,N_9913);
and UO_966 (O_966,N_9908,N_9947);
nor UO_967 (O_967,N_9987,N_9991);
nor UO_968 (O_968,N_9982,N_9976);
or UO_969 (O_969,N_9965,N_9999);
or UO_970 (O_970,N_9966,N_9936);
nor UO_971 (O_971,N_9903,N_9915);
nor UO_972 (O_972,N_9911,N_9954);
or UO_973 (O_973,N_9915,N_9963);
nand UO_974 (O_974,N_9904,N_9974);
and UO_975 (O_975,N_9903,N_9969);
nand UO_976 (O_976,N_9998,N_9990);
and UO_977 (O_977,N_9941,N_9980);
nand UO_978 (O_978,N_9937,N_9970);
xnor UO_979 (O_979,N_9972,N_9900);
or UO_980 (O_980,N_9910,N_9956);
or UO_981 (O_981,N_9960,N_9972);
nand UO_982 (O_982,N_9922,N_9953);
and UO_983 (O_983,N_9983,N_9955);
nand UO_984 (O_984,N_9904,N_9936);
xor UO_985 (O_985,N_9944,N_9998);
nor UO_986 (O_986,N_9985,N_9951);
and UO_987 (O_987,N_9968,N_9933);
and UO_988 (O_988,N_9925,N_9922);
nand UO_989 (O_989,N_9981,N_9900);
nor UO_990 (O_990,N_9928,N_9912);
nand UO_991 (O_991,N_9918,N_9990);
and UO_992 (O_992,N_9922,N_9986);
xor UO_993 (O_993,N_9995,N_9917);
or UO_994 (O_994,N_9939,N_9932);
nor UO_995 (O_995,N_9970,N_9968);
or UO_996 (O_996,N_9929,N_9963);
and UO_997 (O_997,N_9955,N_9923);
xor UO_998 (O_998,N_9955,N_9936);
nor UO_999 (O_999,N_9923,N_9968);
or UO_1000 (O_1000,N_9991,N_9951);
and UO_1001 (O_1001,N_9999,N_9934);
and UO_1002 (O_1002,N_9957,N_9973);
or UO_1003 (O_1003,N_9978,N_9911);
nand UO_1004 (O_1004,N_9963,N_9980);
and UO_1005 (O_1005,N_9925,N_9900);
nand UO_1006 (O_1006,N_9992,N_9903);
xor UO_1007 (O_1007,N_9972,N_9976);
xor UO_1008 (O_1008,N_9918,N_9947);
nand UO_1009 (O_1009,N_9996,N_9900);
nor UO_1010 (O_1010,N_9960,N_9958);
nor UO_1011 (O_1011,N_9916,N_9967);
and UO_1012 (O_1012,N_9935,N_9927);
or UO_1013 (O_1013,N_9948,N_9949);
nand UO_1014 (O_1014,N_9984,N_9926);
nand UO_1015 (O_1015,N_9940,N_9907);
nand UO_1016 (O_1016,N_9933,N_9995);
nor UO_1017 (O_1017,N_9932,N_9918);
nor UO_1018 (O_1018,N_9934,N_9976);
and UO_1019 (O_1019,N_9996,N_9927);
or UO_1020 (O_1020,N_9901,N_9980);
nor UO_1021 (O_1021,N_9996,N_9989);
and UO_1022 (O_1022,N_9941,N_9999);
nor UO_1023 (O_1023,N_9917,N_9902);
xnor UO_1024 (O_1024,N_9943,N_9964);
nor UO_1025 (O_1025,N_9977,N_9905);
and UO_1026 (O_1026,N_9920,N_9901);
and UO_1027 (O_1027,N_9976,N_9913);
or UO_1028 (O_1028,N_9988,N_9904);
nand UO_1029 (O_1029,N_9999,N_9969);
nand UO_1030 (O_1030,N_9904,N_9908);
and UO_1031 (O_1031,N_9936,N_9985);
xnor UO_1032 (O_1032,N_9997,N_9927);
nand UO_1033 (O_1033,N_9989,N_9907);
and UO_1034 (O_1034,N_9912,N_9923);
or UO_1035 (O_1035,N_9923,N_9947);
xnor UO_1036 (O_1036,N_9988,N_9990);
and UO_1037 (O_1037,N_9913,N_9945);
and UO_1038 (O_1038,N_9977,N_9908);
or UO_1039 (O_1039,N_9911,N_9985);
and UO_1040 (O_1040,N_9947,N_9935);
and UO_1041 (O_1041,N_9905,N_9955);
and UO_1042 (O_1042,N_9946,N_9959);
nand UO_1043 (O_1043,N_9999,N_9925);
or UO_1044 (O_1044,N_9961,N_9986);
or UO_1045 (O_1045,N_9984,N_9908);
nand UO_1046 (O_1046,N_9983,N_9958);
nand UO_1047 (O_1047,N_9973,N_9924);
xor UO_1048 (O_1048,N_9915,N_9956);
or UO_1049 (O_1049,N_9939,N_9948);
and UO_1050 (O_1050,N_9962,N_9919);
or UO_1051 (O_1051,N_9906,N_9920);
and UO_1052 (O_1052,N_9995,N_9953);
and UO_1053 (O_1053,N_9982,N_9942);
nand UO_1054 (O_1054,N_9910,N_9988);
nand UO_1055 (O_1055,N_9931,N_9922);
nand UO_1056 (O_1056,N_9984,N_9956);
and UO_1057 (O_1057,N_9911,N_9995);
and UO_1058 (O_1058,N_9934,N_9998);
xor UO_1059 (O_1059,N_9989,N_9962);
nor UO_1060 (O_1060,N_9936,N_9989);
or UO_1061 (O_1061,N_9972,N_9977);
nor UO_1062 (O_1062,N_9933,N_9954);
or UO_1063 (O_1063,N_9950,N_9986);
or UO_1064 (O_1064,N_9936,N_9997);
nor UO_1065 (O_1065,N_9977,N_9944);
nor UO_1066 (O_1066,N_9958,N_9957);
xor UO_1067 (O_1067,N_9954,N_9918);
nand UO_1068 (O_1068,N_9997,N_9955);
and UO_1069 (O_1069,N_9931,N_9907);
and UO_1070 (O_1070,N_9945,N_9957);
nand UO_1071 (O_1071,N_9979,N_9968);
nand UO_1072 (O_1072,N_9900,N_9954);
nor UO_1073 (O_1073,N_9979,N_9963);
and UO_1074 (O_1074,N_9942,N_9972);
and UO_1075 (O_1075,N_9950,N_9953);
nor UO_1076 (O_1076,N_9989,N_9951);
or UO_1077 (O_1077,N_9991,N_9947);
and UO_1078 (O_1078,N_9910,N_9920);
nand UO_1079 (O_1079,N_9910,N_9929);
nor UO_1080 (O_1080,N_9908,N_9945);
or UO_1081 (O_1081,N_9948,N_9926);
and UO_1082 (O_1082,N_9948,N_9953);
or UO_1083 (O_1083,N_9913,N_9929);
nand UO_1084 (O_1084,N_9900,N_9907);
and UO_1085 (O_1085,N_9996,N_9974);
nand UO_1086 (O_1086,N_9949,N_9905);
and UO_1087 (O_1087,N_9958,N_9974);
or UO_1088 (O_1088,N_9961,N_9907);
nor UO_1089 (O_1089,N_9997,N_9916);
nor UO_1090 (O_1090,N_9982,N_9997);
nor UO_1091 (O_1091,N_9993,N_9910);
xnor UO_1092 (O_1092,N_9934,N_9982);
nand UO_1093 (O_1093,N_9982,N_9925);
xor UO_1094 (O_1094,N_9932,N_9920);
and UO_1095 (O_1095,N_9988,N_9991);
or UO_1096 (O_1096,N_9957,N_9994);
or UO_1097 (O_1097,N_9990,N_9992);
nand UO_1098 (O_1098,N_9901,N_9952);
nand UO_1099 (O_1099,N_9967,N_9996);
and UO_1100 (O_1100,N_9906,N_9900);
nand UO_1101 (O_1101,N_9998,N_9928);
or UO_1102 (O_1102,N_9925,N_9908);
nand UO_1103 (O_1103,N_9973,N_9940);
or UO_1104 (O_1104,N_9981,N_9945);
nor UO_1105 (O_1105,N_9958,N_9923);
xnor UO_1106 (O_1106,N_9963,N_9928);
nand UO_1107 (O_1107,N_9907,N_9920);
and UO_1108 (O_1108,N_9901,N_9958);
nand UO_1109 (O_1109,N_9958,N_9975);
or UO_1110 (O_1110,N_9973,N_9960);
nand UO_1111 (O_1111,N_9995,N_9972);
nor UO_1112 (O_1112,N_9947,N_9925);
nor UO_1113 (O_1113,N_9907,N_9971);
nor UO_1114 (O_1114,N_9948,N_9945);
nand UO_1115 (O_1115,N_9946,N_9929);
or UO_1116 (O_1116,N_9962,N_9983);
nor UO_1117 (O_1117,N_9964,N_9926);
nor UO_1118 (O_1118,N_9992,N_9947);
xor UO_1119 (O_1119,N_9943,N_9951);
or UO_1120 (O_1120,N_9956,N_9980);
or UO_1121 (O_1121,N_9998,N_9909);
nand UO_1122 (O_1122,N_9986,N_9900);
nand UO_1123 (O_1123,N_9971,N_9917);
xnor UO_1124 (O_1124,N_9976,N_9945);
nor UO_1125 (O_1125,N_9969,N_9916);
nand UO_1126 (O_1126,N_9901,N_9930);
nor UO_1127 (O_1127,N_9970,N_9955);
and UO_1128 (O_1128,N_9983,N_9936);
and UO_1129 (O_1129,N_9993,N_9977);
xor UO_1130 (O_1130,N_9964,N_9945);
xor UO_1131 (O_1131,N_9960,N_9953);
or UO_1132 (O_1132,N_9933,N_9908);
nor UO_1133 (O_1133,N_9909,N_9965);
xor UO_1134 (O_1134,N_9956,N_9946);
xnor UO_1135 (O_1135,N_9951,N_9967);
nor UO_1136 (O_1136,N_9957,N_9906);
or UO_1137 (O_1137,N_9942,N_9927);
nor UO_1138 (O_1138,N_9928,N_9953);
or UO_1139 (O_1139,N_9933,N_9986);
and UO_1140 (O_1140,N_9908,N_9926);
nor UO_1141 (O_1141,N_9989,N_9934);
nor UO_1142 (O_1142,N_9926,N_9995);
xor UO_1143 (O_1143,N_9909,N_9996);
nand UO_1144 (O_1144,N_9927,N_9910);
nor UO_1145 (O_1145,N_9954,N_9993);
or UO_1146 (O_1146,N_9930,N_9969);
or UO_1147 (O_1147,N_9997,N_9980);
nor UO_1148 (O_1148,N_9927,N_9995);
or UO_1149 (O_1149,N_9938,N_9965);
nand UO_1150 (O_1150,N_9979,N_9985);
nor UO_1151 (O_1151,N_9906,N_9911);
xnor UO_1152 (O_1152,N_9928,N_9917);
nand UO_1153 (O_1153,N_9966,N_9902);
nor UO_1154 (O_1154,N_9973,N_9984);
xor UO_1155 (O_1155,N_9988,N_9960);
nor UO_1156 (O_1156,N_9952,N_9942);
nand UO_1157 (O_1157,N_9965,N_9905);
or UO_1158 (O_1158,N_9989,N_9988);
and UO_1159 (O_1159,N_9963,N_9990);
nor UO_1160 (O_1160,N_9948,N_9983);
or UO_1161 (O_1161,N_9984,N_9913);
and UO_1162 (O_1162,N_9961,N_9980);
nor UO_1163 (O_1163,N_9998,N_9984);
or UO_1164 (O_1164,N_9959,N_9969);
xnor UO_1165 (O_1165,N_9937,N_9987);
and UO_1166 (O_1166,N_9977,N_9936);
or UO_1167 (O_1167,N_9933,N_9975);
or UO_1168 (O_1168,N_9940,N_9954);
and UO_1169 (O_1169,N_9903,N_9995);
or UO_1170 (O_1170,N_9991,N_9998);
nand UO_1171 (O_1171,N_9980,N_9959);
nor UO_1172 (O_1172,N_9937,N_9946);
nand UO_1173 (O_1173,N_9929,N_9916);
nor UO_1174 (O_1174,N_9952,N_9935);
nor UO_1175 (O_1175,N_9978,N_9985);
nand UO_1176 (O_1176,N_9978,N_9919);
nand UO_1177 (O_1177,N_9913,N_9971);
nor UO_1178 (O_1178,N_9934,N_9952);
nand UO_1179 (O_1179,N_9980,N_9919);
and UO_1180 (O_1180,N_9970,N_9954);
nand UO_1181 (O_1181,N_9980,N_9993);
nor UO_1182 (O_1182,N_9995,N_9955);
nor UO_1183 (O_1183,N_9931,N_9972);
and UO_1184 (O_1184,N_9942,N_9907);
xnor UO_1185 (O_1185,N_9929,N_9936);
nor UO_1186 (O_1186,N_9954,N_9904);
xnor UO_1187 (O_1187,N_9950,N_9918);
xor UO_1188 (O_1188,N_9980,N_9912);
xor UO_1189 (O_1189,N_9990,N_9905);
or UO_1190 (O_1190,N_9944,N_9907);
or UO_1191 (O_1191,N_9926,N_9904);
or UO_1192 (O_1192,N_9942,N_9958);
and UO_1193 (O_1193,N_9929,N_9917);
xor UO_1194 (O_1194,N_9980,N_9905);
and UO_1195 (O_1195,N_9950,N_9992);
and UO_1196 (O_1196,N_9909,N_9907);
nand UO_1197 (O_1197,N_9988,N_9921);
and UO_1198 (O_1198,N_9900,N_9923);
xor UO_1199 (O_1199,N_9945,N_9959);
and UO_1200 (O_1200,N_9980,N_9931);
nand UO_1201 (O_1201,N_9954,N_9917);
and UO_1202 (O_1202,N_9972,N_9919);
and UO_1203 (O_1203,N_9957,N_9983);
nor UO_1204 (O_1204,N_9983,N_9900);
xor UO_1205 (O_1205,N_9916,N_9972);
nand UO_1206 (O_1206,N_9968,N_9972);
and UO_1207 (O_1207,N_9934,N_9979);
xor UO_1208 (O_1208,N_9974,N_9994);
nand UO_1209 (O_1209,N_9983,N_9949);
nand UO_1210 (O_1210,N_9967,N_9902);
and UO_1211 (O_1211,N_9911,N_9938);
nor UO_1212 (O_1212,N_9964,N_9970);
nor UO_1213 (O_1213,N_9926,N_9921);
nor UO_1214 (O_1214,N_9967,N_9986);
and UO_1215 (O_1215,N_9918,N_9971);
or UO_1216 (O_1216,N_9982,N_9980);
or UO_1217 (O_1217,N_9946,N_9984);
nand UO_1218 (O_1218,N_9911,N_9956);
xor UO_1219 (O_1219,N_9911,N_9945);
nor UO_1220 (O_1220,N_9972,N_9961);
nand UO_1221 (O_1221,N_9941,N_9937);
nand UO_1222 (O_1222,N_9911,N_9920);
and UO_1223 (O_1223,N_9975,N_9908);
and UO_1224 (O_1224,N_9933,N_9917);
nor UO_1225 (O_1225,N_9964,N_9911);
or UO_1226 (O_1226,N_9923,N_9926);
or UO_1227 (O_1227,N_9914,N_9993);
nand UO_1228 (O_1228,N_9938,N_9910);
nor UO_1229 (O_1229,N_9984,N_9997);
xnor UO_1230 (O_1230,N_9991,N_9977);
nor UO_1231 (O_1231,N_9962,N_9955);
nor UO_1232 (O_1232,N_9992,N_9994);
nor UO_1233 (O_1233,N_9959,N_9973);
or UO_1234 (O_1234,N_9902,N_9915);
nand UO_1235 (O_1235,N_9911,N_9977);
and UO_1236 (O_1236,N_9901,N_9966);
and UO_1237 (O_1237,N_9902,N_9928);
nor UO_1238 (O_1238,N_9993,N_9978);
nor UO_1239 (O_1239,N_9924,N_9964);
nor UO_1240 (O_1240,N_9930,N_9988);
xor UO_1241 (O_1241,N_9962,N_9985);
or UO_1242 (O_1242,N_9919,N_9998);
nand UO_1243 (O_1243,N_9987,N_9976);
and UO_1244 (O_1244,N_9919,N_9921);
nand UO_1245 (O_1245,N_9943,N_9987);
or UO_1246 (O_1246,N_9946,N_9952);
nand UO_1247 (O_1247,N_9933,N_9976);
nand UO_1248 (O_1248,N_9976,N_9911);
nor UO_1249 (O_1249,N_9931,N_9938);
nand UO_1250 (O_1250,N_9978,N_9959);
nand UO_1251 (O_1251,N_9989,N_9974);
nand UO_1252 (O_1252,N_9998,N_9911);
nor UO_1253 (O_1253,N_9928,N_9981);
nand UO_1254 (O_1254,N_9993,N_9999);
xnor UO_1255 (O_1255,N_9954,N_9913);
or UO_1256 (O_1256,N_9913,N_9978);
or UO_1257 (O_1257,N_9964,N_9922);
nor UO_1258 (O_1258,N_9910,N_9968);
and UO_1259 (O_1259,N_9972,N_9978);
or UO_1260 (O_1260,N_9915,N_9944);
and UO_1261 (O_1261,N_9952,N_9930);
or UO_1262 (O_1262,N_9947,N_9905);
or UO_1263 (O_1263,N_9995,N_9990);
or UO_1264 (O_1264,N_9911,N_9941);
nor UO_1265 (O_1265,N_9973,N_9953);
or UO_1266 (O_1266,N_9951,N_9981);
and UO_1267 (O_1267,N_9943,N_9904);
nand UO_1268 (O_1268,N_9988,N_9953);
and UO_1269 (O_1269,N_9919,N_9982);
nor UO_1270 (O_1270,N_9932,N_9902);
and UO_1271 (O_1271,N_9985,N_9997);
and UO_1272 (O_1272,N_9908,N_9959);
or UO_1273 (O_1273,N_9934,N_9957);
nor UO_1274 (O_1274,N_9937,N_9951);
nor UO_1275 (O_1275,N_9948,N_9970);
or UO_1276 (O_1276,N_9995,N_9987);
and UO_1277 (O_1277,N_9973,N_9919);
nand UO_1278 (O_1278,N_9969,N_9912);
nand UO_1279 (O_1279,N_9949,N_9940);
nand UO_1280 (O_1280,N_9981,N_9926);
and UO_1281 (O_1281,N_9986,N_9974);
nand UO_1282 (O_1282,N_9956,N_9923);
nand UO_1283 (O_1283,N_9958,N_9981);
nand UO_1284 (O_1284,N_9904,N_9999);
and UO_1285 (O_1285,N_9979,N_9970);
nor UO_1286 (O_1286,N_9972,N_9914);
and UO_1287 (O_1287,N_9967,N_9956);
xor UO_1288 (O_1288,N_9963,N_9942);
and UO_1289 (O_1289,N_9950,N_9945);
and UO_1290 (O_1290,N_9948,N_9906);
or UO_1291 (O_1291,N_9993,N_9934);
and UO_1292 (O_1292,N_9947,N_9917);
or UO_1293 (O_1293,N_9965,N_9983);
nand UO_1294 (O_1294,N_9914,N_9937);
and UO_1295 (O_1295,N_9909,N_9918);
or UO_1296 (O_1296,N_9988,N_9999);
nor UO_1297 (O_1297,N_9992,N_9966);
and UO_1298 (O_1298,N_9981,N_9964);
nor UO_1299 (O_1299,N_9933,N_9961);
and UO_1300 (O_1300,N_9909,N_9967);
or UO_1301 (O_1301,N_9968,N_9934);
and UO_1302 (O_1302,N_9995,N_9919);
or UO_1303 (O_1303,N_9910,N_9995);
or UO_1304 (O_1304,N_9913,N_9952);
or UO_1305 (O_1305,N_9948,N_9931);
or UO_1306 (O_1306,N_9947,N_9920);
nand UO_1307 (O_1307,N_9958,N_9909);
nand UO_1308 (O_1308,N_9959,N_9942);
nor UO_1309 (O_1309,N_9947,N_9901);
nand UO_1310 (O_1310,N_9963,N_9989);
or UO_1311 (O_1311,N_9997,N_9989);
nor UO_1312 (O_1312,N_9969,N_9973);
nand UO_1313 (O_1313,N_9916,N_9992);
nor UO_1314 (O_1314,N_9994,N_9955);
and UO_1315 (O_1315,N_9958,N_9945);
nor UO_1316 (O_1316,N_9981,N_9979);
nor UO_1317 (O_1317,N_9946,N_9983);
and UO_1318 (O_1318,N_9964,N_9933);
nand UO_1319 (O_1319,N_9964,N_9976);
nor UO_1320 (O_1320,N_9992,N_9955);
nor UO_1321 (O_1321,N_9979,N_9948);
or UO_1322 (O_1322,N_9901,N_9923);
and UO_1323 (O_1323,N_9963,N_9968);
nor UO_1324 (O_1324,N_9960,N_9945);
and UO_1325 (O_1325,N_9978,N_9927);
and UO_1326 (O_1326,N_9956,N_9969);
nand UO_1327 (O_1327,N_9900,N_9992);
and UO_1328 (O_1328,N_9940,N_9950);
nor UO_1329 (O_1329,N_9962,N_9936);
nor UO_1330 (O_1330,N_9971,N_9955);
and UO_1331 (O_1331,N_9973,N_9915);
or UO_1332 (O_1332,N_9926,N_9936);
nand UO_1333 (O_1333,N_9953,N_9958);
nand UO_1334 (O_1334,N_9993,N_9944);
nor UO_1335 (O_1335,N_9970,N_9932);
and UO_1336 (O_1336,N_9909,N_9960);
or UO_1337 (O_1337,N_9901,N_9984);
nand UO_1338 (O_1338,N_9902,N_9975);
or UO_1339 (O_1339,N_9995,N_9921);
xor UO_1340 (O_1340,N_9947,N_9921);
and UO_1341 (O_1341,N_9902,N_9933);
nand UO_1342 (O_1342,N_9913,N_9967);
nor UO_1343 (O_1343,N_9979,N_9992);
nor UO_1344 (O_1344,N_9904,N_9939);
nand UO_1345 (O_1345,N_9948,N_9963);
nand UO_1346 (O_1346,N_9960,N_9998);
nand UO_1347 (O_1347,N_9970,N_9994);
xor UO_1348 (O_1348,N_9971,N_9943);
nand UO_1349 (O_1349,N_9934,N_9997);
or UO_1350 (O_1350,N_9944,N_9917);
or UO_1351 (O_1351,N_9950,N_9957);
xnor UO_1352 (O_1352,N_9933,N_9942);
nor UO_1353 (O_1353,N_9941,N_9926);
xor UO_1354 (O_1354,N_9922,N_9915);
and UO_1355 (O_1355,N_9955,N_9954);
nor UO_1356 (O_1356,N_9942,N_9981);
nor UO_1357 (O_1357,N_9982,N_9904);
nor UO_1358 (O_1358,N_9920,N_9979);
nand UO_1359 (O_1359,N_9928,N_9930);
xnor UO_1360 (O_1360,N_9942,N_9936);
and UO_1361 (O_1361,N_9906,N_9923);
nor UO_1362 (O_1362,N_9918,N_9941);
nand UO_1363 (O_1363,N_9951,N_9999);
and UO_1364 (O_1364,N_9986,N_9913);
or UO_1365 (O_1365,N_9947,N_9943);
or UO_1366 (O_1366,N_9944,N_9999);
nor UO_1367 (O_1367,N_9923,N_9932);
or UO_1368 (O_1368,N_9995,N_9940);
nor UO_1369 (O_1369,N_9936,N_9974);
nand UO_1370 (O_1370,N_9965,N_9975);
xnor UO_1371 (O_1371,N_9962,N_9933);
or UO_1372 (O_1372,N_9968,N_9911);
nand UO_1373 (O_1373,N_9980,N_9974);
nor UO_1374 (O_1374,N_9942,N_9950);
or UO_1375 (O_1375,N_9945,N_9954);
nand UO_1376 (O_1376,N_9946,N_9918);
nor UO_1377 (O_1377,N_9965,N_9934);
nor UO_1378 (O_1378,N_9946,N_9903);
and UO_1379 (O_1379,N_9998,N_9972);
nand UO_1380 (O_1380,N_9900,N_9971);
and UO_1381 (O_1381,N_9978,N_9904);
and UO_1382 (O_1382,N_9919,N_9997);
and UO_1383 (O_1383,N_9929,N_9939);
and UO_1384 (O_1384,N_9984,N_9975);
nand UO_1385 (O_1385,N_9906,N_9955);
nand UO_1386 (O_1386,N_9995,N_9957);
and UO_1387 (O_1387,N_9925,N_9962);
nor UO_1388 (O_1388,N_9901,N_9989);
nand UO_1389 (O_1389,N_9927,N_9948);
nor UO_1390 (O_1390,N_9982,N_9909);
nor UO_1391 (O_1391,N_9940,N_9958);
nand UO_1392 (O_1392,N_9927,N_9977);
nor UO_1393 (O_1393,N_9962,N_9951);
and UO_1394 (O_1394,N_9940,N_9925);
or UO_1395 (O_1395,N_9962,N_9916);
or UO_1396 (O_1396,N_9973,N_9949);
nor UO_1397 (O_1397,N_9931,N_9992);
and UO_1398 (O_1398,N_9999,N_9980);
nor UO_1399 (O_1399,N_9980,N_9936);
nor UO_1400 (O_1400,N_9922,N_9904);
and UO_1401 (O_1401,N_9996,N_9959);
nor UO_1402 (O_1402,N_9969,N_9984);
xnor UO_1403 (O_1403,N_9957,N_9981);
nand UO_1404 (O_1404,N_9937,N_9929);
nor UO_1405 (O_1405,N_9960,N_9991);
and UO_1406 (O_1406,N_9993,N_9981);
nand UO_1407 (O_1407,N_9914,N_9938);
and UO_1408 (O_1408,N_9935,N_9908);
or UO_1409 (O_1409,N_9980,N_9975);
and UO_1410 (O_1410,N_9912,N_9934);
nand UO_1411 (O_1411,N_9914,N_9956);
nor UO_1412 (O_1412,N_9979,N_9973);
nand UO_1413 (O_1413,N_9920,N_9921);
nor UO_1414 (O_1414,N_9913,N_9949);
nor UO_1415 (O_1415,N_9957,N_9959);
nand UO_1416 (O_1416,N_9927,N_9922);
or UO_1417 (O_1417,N_9994,N_9959);
nand UO_1418 (O_1418,N_9955,N_9982);
and UO_1419 (O_1419,N_9916,N_9922);
nor UO_1420 (O_1420,N_9901,N_9985);
and UO_1421 (O_1421,N_9923,N_9989);
nor UO_1422 (O_1422,N_9906,N_9972);
xnor UO_1423 (O_1423,N_9935,N_9989);
nor UO_1424 (O_1424,N_9934,N_9963);
nor UO_1425 (O_1425,N_9974,N_9951);
or UO_1426 (O_1426,N_9985,N_9939);
nand UO_1427 (O_1427,N_9999,N_9967);
nor UO_1428 (O_1428,N_9926,N_9957);
and UO_1429 (O_1429,N_9997,N_9992);
nor UO_1430 (O_1430,N_9933,N_9938);
xnor UO_1431 (O_1431,N_9966,N_9923);
or UO_1432 (O_1432,N_9964,N_9985);
nand UO_1433 (O_1433,N_9943,N_9926);
or UO_1434 (O_1434,N_9933,N_9991);
and UO_1435 (O_1435,N_9943,N_9937);
nor UO_1436 (O_1436,N_9953,N_9992);
or UO_1437 (O_1437,N_9985,N_9934);
or UO_1438 (O_1438,N_9913,N_9985);
xor UO_1439 (O_1439,N_9974,N_9943);
nor UO_1440 (O_1440,N_9909,N_9999);
or UO_1441 (O_1441,N_9994,N_9912);
nand UO_1442 (O_1442,N_9908,N_9997);
nand UO_1443 (O_1443,N_9956,N_9952);
nand UO_1444 (O_1444,N_9953,N_9926);
nor UO_1445 (O_1445,N_9973,N_9932);
nor UO_1446 (O_1446,N_9963,N_9961);
nor UO_1447 (O_1447,N_9952,N_9970);
nor UO_1448 (O_1448,N_9937,N_9912);
nor UO_1449 (O_1449,N_9986,N_9982);
or UO_1450 (O_1450,N_9921,N_9913);
xnor UO_1451 (O_1451,N_9914,N_9918);
and UO_1452 (O_1452,N_9953,N_9954);
nor UO_1453 (O_1453,N_9929,N_9947);
and UO_1454 (O_1454,N_9998,N_9952);
nand UO_1455 (O_1455,N_9901,N_9998);
and UO_1456 (O_1456,N_9902,N_9943);
xnor UO_1457 (O_1457,N_9944,N_9961);
nand UO_1458 (O_1458,N_9943,N_9928);
nor UO_1459 (O_1459,N_9961,N_9983);
nand UO_1460 (O_1460,N_9988,N_9956);
nand UO_1461 (O_1461,N_9929,N_9980);
and UO_1462 (O_1462,N_9927,N_9949);
nand UO_1463 (O_1463,N_9901,N_9909);
and UO_1464 (O_1464,N_9905,N_9981);
and UO_1465 (O_1465,N_9991,N_9928);
or UO_1466 (O_1466,N_9986,N_9963);
nand UO_1467 (O_1467,N_9961,N_9959);
or UO_1468 (O_1468,N_9906,N_9934);
and UO_1469 (O_1469,N_9901,N_9908);
nand UO_1470 (O_1470,N_9975,N_9924);
and UO_1471 (O_1471,N_9914,N_9990);
or UO_1472 (O_1472,N_9935,N_9998);
nand UO_1473 (O_1473,N_9909,N_9987);
nand UO_1474 (O_1474,N_9994,N_9924);
and UO_1475 (O_1475,N_9918,N_9917);
or UO_1476 (O_1476,N_9978,N_9902);
and UO_1477 (O_1477,N_9985,N_9967);
nand UO_1478 (O_1478,N_9907,N_9950);
nand UO_1479 (O_1479,N_9906,N_9915);
xnor UO_1480 (O_1480,N_9984,N_9955);
nand UO_1481 (O_1481,N_9941,N_9978);
or UO_1482 (O_1482,N_9967,N_9925);
and UO_1483 (O_1483,N_9902,N_9986);
and UO_1484 (O_1484,N_9927,N_9907);
or UO_1485 (O_1485,N_9936,N_9943);
nand UO_1486 (O_1486,N_9959,N_9901);
nor UO_1487 (O_1487,N_9902,N_9952);
or UO_1488 (O_1488,N_9964,N_9984);
nand UO_1489 (O_1489,N_9986,N_9907);
and UO_1490 (O_1490,N_9953,N_9907);
or UO_1491 (O_1491,N_9982,N_9991);
xor UO_1492 (O_1492,N_9957,N_9904);
and UO_1493 (O_1493,N_9982,N_9958);
xor UO_1494 (O_1494,N_9965,N_9957);
nand UO_1495 (O_1495,N_9922,N_9969);
xnor UO_1496 (O_1496,N_9957,N_9947);
or UO_1497 (O_1497,N_9945,N_9906);
nand UO_1498 (O_1498,N_9925,N_9905);
or UO_1499 (O_1499,N_9959,N_9968);
endmodule