module basic_1500_15000_2000_3_levels_1xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10003,N_10004,N_10005,N_10007,N_10008,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10018,N_10019,N_10020,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10030,N_10031,N_10033,N_10035,N_10037,N_10039,N_10040,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10050,N_10052,N_10053,N_10055,N_10056,N_10059,N_10060,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10082,N_10083,N_10085,N_10086,N_10087,N_10088,N_10089,N_10091,N_10093,N_10094,N_10095,N_10096,N_10097,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10108,N_10109,N_10110,N_10111,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10137,N_10138,N_10139,N_10140,N_10142,N_10143,N_10144,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10161,N_10162,N_10163,N_10168,N_10169,N_10171,N_10172,N_10174,N_10175,N_10176,N_10177,N_10179,N_10180,N_10181,N_10182,N_10183,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10207,N_10208,N_10209,N_10210,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10219,N_10220,N_10222,N_10224,N_10225,N_10226,N_10228,N_10229,N_10231,N_10232,N_10233,N_10234,N_10235,N_10237,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10249,N_10252,N_10253,N_10254,N_10255,N_10256,N_10258,N_10259,N_10260,N_10262,N_10263,N_10265,N_10266,N_10268,N_10269,N_10270,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10279,N_10280,N_10281,N_10282,N_10284,N_10285,N_10286,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10299,N_10300,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10311,N_10312,N_10313,N_10314,N_10316,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10341,N_10342,N_10346,N_10347,N_10349,N_10350,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10383,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10394,N_10395,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10438,N_10440,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10459,N_10460,N_10461,N_10462,N_10463,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10476,N_10477,N_10478,N_10479,N_10480,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10490,N_10492,N_10494,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10554,N_10556,N_10557,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10576,N_10577,N_10578,N_10579,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10594,N_10595,N_10596,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10617,N_10619,N_10621,N_10622,N_10623,N_10624,N_10626,N_10627,N_10628,N_10629,N_10630,N_10632,N_10634,N_10635,N_10636,N_10638,N_10639,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10649,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10663,N_10664,N_10665,N_10667,N_10668,N_10669,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10691,N_10692,N_10696,N_10697,N_10698,N_10699,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10720,N_10723,N_10725,N_10726,N_10727,N_10728,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10738,N_10739,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10793,N_10794,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10837,N_10838,N_10839,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10849,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10859,N_10860,N_10861,N_10863,N_10864,N_10866,N_10867,N_10868,N_10869,N_10871,N_10872,N_10873,N_10875,N_10876,N_10877,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10931,N_10932,N_10933,N_10934,N_10935,N_10938,N_10940,N_10941,N_10942,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10958,N_10959,N_10960,N_10962,N_10963,N_10964,N_10966,N_10967,N_10968,N_10970,N_10972,N_10974,N_10975,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11016,N_11018,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11041,N_11043,N_11044,N_11045,N_11046,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11055,N_11056,N_11057,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11099,N_11100,N_11101,N_11102,N_11103,N_11105,N_11106,N_11107,N_11108,N_11109,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11122,N_11125,N_11126,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11138,N_11139,N_11140,N_11142,N_11143,N_11144,N_11148,N_11149,N_11150,N_11151,N_11152,N_11154,N_11155,N_11157,N_11158,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11167,N_11168,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11185,N_11186,N_11187,N_11189,N_11190,N_11191,N_11192,N_11194,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11209,N_11212,N_11213,N_11214,N_11215,N_11216,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11275,N_11276,N_11277,N_11279,N_11280,N_11281,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11364,N_11365,N_11367,N_11368,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11384,N_11385,N_11386,N_11387,N_11388,N_11390,N_11392,N_11393,N_11394,N_11395,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11405,N_11407,N_11408,N_11409,N_11411,N_11412,N_11413,N_11414,N_11415,N_11417,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11427,N_11428,N_11429,N_11430,N_11431,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11445,N_11446,N_11447,N_11448,N_11449,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11459,N_11460,N_11462,N_11463,N_11464,N_11465,N_11468,N_11469,N_11470,N_11471,N_11472,N_11474,N_11476,N_11477,N_11478,N_11479,N_11480,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11497,N_11498,N_11500,N_11503,N_11504,N_11505,N_11509,N_11510,N_11512,N_11513,N_11514,N_11515,N_11520,N_11521,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11542,N_11543,N_11544,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11559,N_11560,N_11561,N_11562,N_11564,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11577,N_11578,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11592,N_11593,N_11594,N_11595,N_11596,N_11599,N_11600,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11611,N_11615,N_11616,N_11617,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11627,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11651,N_11652,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11678,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11689,N_11690,N_11691,N_11692,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11713,N_11715,N_11717,N_11718,N_11721,N_11723,N_11725,N_11726,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11749,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11761,N_11762,N_11763,N_11764,N_11766,N_11768,N_11769,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11779,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11798,N_11799,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11821,N_11822,N_11824,N_11826,N_11827,N_11828,N_11829,N_11830,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11853,N_11855,N_11857,N_11858,N_11859,N_11860,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11872,N_11873,N_11878,N_11879,N_11881,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11918,N_11919,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11932,N_11933,N_11934,N_11936,N_11937,N_11938,N_11940,N_11941,N_11942,N_11943,N_11944,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11958,N_11959,N_11961,N_11962,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11973,N_11974,N_11976,N_11977,N_11978,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11987,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11996,N_11997,N_11999,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12033,N_12034,N_12035,N_12037,N_12038,N_12039,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12050,N_12051,N_12054,N_12055,N_12056,N_12058,N_12059,N_12060,N_12061,N_12062,N_12065,N_12066,N_12068,N_12069,N_12070,N_12072,N_12073,N_12074,N_12075,N_12077,N_12080,N_12081,N_12083,N_12086,N_12087,N_12088,N_12090,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12099,N_12100,N_12101,N_12102,N_12105,N_12106,N_12108,N_12109,N_12110,N_12112,N_12113,N_12114,N_12116,N_12117,N_12119,N_12120,N_12121,N_12123,N_12124,N_12125,N_12126,N_12129,N_12132,N_12133,N_12136,N_12137,N_12138,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12151,N_12153,N_12154,N_12155,N_12157,N_12158,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12170,N_12171,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12187,N_12188,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12203,N_12204,N_12207,N_12208,N_12209,N_12210,N_12211,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12226,N_12227,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12251,N_12252,N_12253,N_12254,N_12255,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12295,N_12297,N_12301,N_12302,N_12305,N_12306,N_12307,N_12308,N_12309,N_12311,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12323,N_12324,N_12327,N_12328,N_12330,N_12331,N_12332,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12355,N_12356,N_12357,N_12358,N_12359,N_12361,N_12362,N_12363,N_12365,N_12366,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12400,N_12401,N_12402,N_12404,N_12405,N_12407,N_12408,N_12409,N_12410,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12421,N_12422,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12440,N_12441,N_12442,N_12443,N_12445,N_12448,N_12449,N_12450,N_12451,N_12452,N_12454,N_12456,N_12457,N_12458,N_12459,N_12461,N_12462,N_12463,N_12464,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12481,N_12482,N_12484,N_12487,N_12488,N_12489,N_12490,N_12491,N_12493,N_12494,N_12496,N_12498,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12512,N_12513,N_12514,N_12516,N_12517,N_12518,N_12519,N_12521,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12531,N_12532,N_12534,N_12536,N_12540,N_12541,N_12542,N_12544,N_12545,N_12548,N_12549,N_12551,N_12552,N_12553,N_12556,N_12558,N_12559,N_12561,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12578,N_12579,N_12580,N_12582,N_12583,N_12584,N_12585,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12595,N_12596,N_12597,N_12598,N_12599,N_12602,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12612,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12621,N_12622,N_12624,N_12625,N_12626,N_12627,N_12629,N_12630,N_12631,N_12632,N_12633,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12649,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12705,N_12706,N_12707,N_12708,N_12710,N_12711,N_12712,N_12714,N_12715,N_12717,N_12718,N_12719,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12730,N_12731,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12765,N_12768,N_12769,N_12770,N_12771,N_12772,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12796,N_12797,N_12798,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12817,N_12818,N_12820,N_12821,N_12823,N_12824,N_12825,N_12827,N_12828,N_12829,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12841,N_12842,N_12843,N_12846,N_12848,N_12849,N_12850,N_12852,N_12853,N_12854,N_12855,N_12856,N_12858,N_12859,N_12861,N_12862,N_12863,N_12864,N_12866,N_12869,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12892,N_12894,N_12895,N_12897,N_12898,N_12899,N_12900,N_12901,N_12903,N_12904,N_12905,N_12906,N_12907,N_12909,N_12911,N_12913,N_12914,N_12916,N_12917,N_12918,N_12919,N_12920,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12937,N_12941,N_12942,N_12943,N_12944,N_12946,N_12948,N_12950,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12965,N_12966,N_12967,N_12968,N_12970,N_12971,N_12972,N_12973,N_12974,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12994,N_12995,N_12996,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13006,N_13007,N_13008,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13021,N_13022,N_13023,N_13025,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13036,N_13037,N_13039,N_13040,N_13041,N_13043,N_13044,N_13045,N_13047,N_13049,N_13051,N_13052,N_13053,N_13055,N_13056,N_13057,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13070,N_13071,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13081,N_13082,N_13083,N_13084,N_13085,N_13087,N_13089,N_13090,N_13091,N_13093,N_13095,N_13096,N_13097,N_13098,N_13100,N_13101,N_13103,N_13104,N_13105,N_13109,N_13111,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13147,N_13152,N_13154,N_13156,N_13157,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13172,N_13173,N_13174,N_13175,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13187,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13201,N_13202,N_13203,N_13204,N_13207,N_13209,N_13210,N_13211,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13231,N_13232,N_13233,N_13234,N_13235,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13244,N_13245,N_13246,N_13247,N_13248,N_13250,N_13251,N_13252,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13271,N_13272,N_13273,N_13274,N_13275,N_13277,N_13278,N_13279,N_13280,N_13281,N_13284,N_13285,N_13286,N_13287,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13297,N_13301,N_13304,N_13305,N_13306,N_13307,N_13308,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13317,N_13319,N_13320,N_13321,N_13322,N_13323,N_13325,N_13326,N_13327,N_13329,N_13330,N_13332,N_13333,N_13336,N_13339,N_13341,N_13343,N_13344,N_13345,N_13348,N_13350,N_13351,N_13352,N_13353,N_13354,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13388,N_13389,N_13390,N_13392,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13403,N_13404,N_13406,N_13407,N_13408,N_13409,N_13411,N_13412,N_13413,N_13414,N_13416,N_13417,N_13418,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13430,N_13431,N_13432,N_13433,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13450,N_13451,N_13453,N_13454,N_13455,N_13456,N_13458,N_13459,N_13460,N_13462,N_13463,N_13464,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13473,N_13474,N_13475,N_13476,N_13477,N_13479,N_13480,N_13482,N_13484,N_13485,N_13486,N_13487,N_13488,N_13490,N_13492,N_13493,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13514,N_13516,N_13517,N_13518,N_13519,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13542,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13564,N_13565,N_13566,N_13568,N_13570,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13579,N_13580,N_13582,N_13583,N_13584,N_13585,N_13586,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13598,N_13600,N_13601,N_13602,N_13604,N_13607,N_13608,N_13609,N_13610,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13628,N_13630,N_13632,N_13633,N_13634,N_13635,N_13636,N_13638,N_13640,N_13641,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13669,N_13671,N_13672,N_13673,N_13674,N_13676,N_13677,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13697,N_13699,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13713,N_13714,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13738,N_13739,N_13740,N_13741,N_13742,N_13745,N_13746,N_13748,N_13749,N_13750,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13784,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13801,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13828,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13840,N_13841,N_13843,N_13845,N_13846,N_13847,N_13848,N_13850,N_13851,N_13853,N_13854,N_13856,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13870,N_13871,N_13872,N_13873,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13882,N_13883,N_13884,N_13885,N_13887,N_13888,N_13889,N_13890,N_13891,N_13893,N_13894,N_13895,N_13896,N_13898,N_13899,N_13900,N_13901,N_13903,N_13904,N_13906,N_13907,N_13908,N_13909,N_13911,N_13914,N_13915,N_13916,N_13917,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13927,N_13928,N_13929,N_13930,N_13931,N_13933,N_13934,N_13936,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13947,N_13948,N_13949,N_13950,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14005,N_14006,N_14007,N_14008,N_14010,N_14011,N_14012,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14023,N_14024,N_14025,N_14026,N_14028,N_14029,N_14030,N_14032,N_14034,N_14035,N_14036,N_14037,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14060,N_14061,N_14062,N_14063,N_14064,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14077,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14086,N_14087,N_14088,N_14089,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14110,N_14112,N_14113,N_14114,N_14115,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14128,N_14129,N_14132,N_14134,N_14135,N_14137,N_14140,N_14142,N_14143,N_14144,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14176,N_14179,N_14180,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14198,N_14199,N_14200,N_14201,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14213,N_14214,N_14215,N_14216,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14227,N_14228,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14248,N_14249,N_14250,N_14251,N_14252,N_14254,N_14255,N_14256,N_14258,N_14260,N_14261,N_14262,N_14264,N_14265,N_14266,N_14267,N_14268,N_14270,N_14271,N_14272,N_14274,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14306,N_14307,N_14308,N_14309,N_14312,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14322,N_14323,N_14326,N_14327,N_14328,N_14330,N_14332,N_14333,N_14334,N_14335,N_14336,N_14338,N_14339,N_14340,N_14342,N_14343,N_14344,N_14347,N_14349,N_14350,N_14351,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14361,N_14362,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14372,N_14373,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14395,N_14397,N_14398,N_14400,N_14402,N_14403,N_14404,N_14405,N_14407,N_14411,N_14412,N_14413,N_14414,N_14417,N_14419,N_14420,N_14421,N_14423,N_14424,N_14425,N_14426,N_14428,N_14429,N_14430,N_14432,N_14433,N_14434,N_14435,N_14436,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14450,N_14451,N_14452,N_14453,N_14454,N_14456,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14470,N_14471,N_14472,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14484,N_14485,N_14487,N_14488,N_14491,N_14492,N_14493,N_14494,N_14496,N_14497,N_14498,N_14500,N_14501,N_14502,N_14505,N_14506,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14517,N_14518,N_14520,N_14521,N_14524,N_14525,N_14526,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14539,N_14540,N_14541,N_14542,N_14543,N_14546,N_14547,N_14548,N_14549,N_14551,N_14553,N_14554,N_14556,N_14557,N_14558,N_14560,N_14561,N_14562,N_14565,N_14567,N_14568,N_14569,N_14570,N_14572,N_14573,N_14574,N_14576,N_14579,N_14580,N_14581,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14590,N_14591,N_14594,N_14595,N_14596,N_14598,N_14599,N_14600,N_14602,N_14603,N_14604,N_14605,N_14607,N_14609,N_14611,N_14612,N_14615,N_14617,N_14618,N_14619,N_14620,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14632,N_14633,N_14635,N_14636,N_14637,N_14639,N_14640,N_14641,N_14643,N_14644,N_14645,N_14646,N_14648,N_14650,N_14651,N_14652,N_14653,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14662,N_14663,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14673,N_14674,N_14675,N_14676,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14689,N_14690,N_14691,N_14692,N_14693,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14721,N_14722,N_14723,N_14724,N_14725,N_14728,N_14729,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14762,N_14763,N_14764,N_14766,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14787,N_14788,N_14789,N_14790,N_14791,N_14793,N_14794,N_14795,N_14796,N_14798,N_14799,N_14800,N_14802,N_14803,N_14804,N_14805,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14827,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14837,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14849,N_14850,N_14851,N_14852,N_14853,N_14855,N_14856,N_14857,N_14858,N_14859,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14868,N_14869,N_14870,N_14872,N_14874,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14894,N_14895,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14914,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14933,N_14934,N_14935,N_14937,N_14938,N_14939,N_14942,N_14943,N_14944,N_14945,N_14947,N_14948,N_14950,N_14951,N_14952,N_14953,N_14954,N_14958,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14980,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14995,N_14996,N_14997,N_14998,N_14999;
nor U0 (N_0,In_1325,In_1292);
and U1 (N_1,In_61,In_1084);
or U2 (N_2,In_178,In_1195);
nand U3 (N_3,In_782,In_21);
nand U4 (N_4,In_759,In_675);
nor U5 (N_5,In_558,In_854);
xnor U6 (N_6,In_983,In_1434);
and U7 (N_7,In_663,In_415);
nor U8 (N_8,In_1426,In_630);
xnor U9 (N_9,In_476,In_343);
and U10 (N_10,In_609,In_708);
or U11 (N_11,In_511,In_1435);
or U12 (N_12,In_1384,In_769);
or U13 (N_13,In_765,In_90);
and U14 (N_14,In_1481,In_193);
nand U15 (N_15,In_1309,In_816);
nand U16 (N_16,In_1457,In_205);
or U17 (N_17,In_74,In_705);
nand U18 (N_18,In_1326,In_1028);
nor U19 (N_19,In_573,In_299);
or U20 (N_20,In_865,In_192);
and U21 (N_21,In_402,In_1089);
nor U22 (N_22,In_410,In_652);
nand U23 (N_23,In_625,In_820);
nor U24 (N_24,In_1013,In_365);
nor U25 (N_25,In_166,In_1188);
and U26 (N_26,In_408,In_662);
and U27 (N_27,In_901,In_751);
and U28 (N_28,In_1494,In_985);
nor U29 (N_29,In_849,In_232);
and U30 (N_30,In_256,In_230);
or U31 (N_31,In_34,In_517);
or U32 (N_32,In_453,In_744);
nor U33 (N_33,In_1454,In_151);
nand U34 (N_34,In_520,In_1035);
and U35 (N_35,In_199,In_799);
or U36 (N_36,In_1160,In_633);
and U37 (N_37,In_946,In_1213);
and U38 (N_38,In_73,In_784);
and U39 (N_39,In_1016,In_1189);
or U40 (N_40,In_1327,In_806);
nor U41 (N_41,In_1487,In_876);
nand U42 (N_42,In_1461,In_309);
and U43 (N_43,In_468,In_1424);
or U44 (N_44,In_1377,In_1446);
nor U45 (N_45,In_145,In_658);
nand U46 (N_46,In_1097,In_804);
and U47 (N_47,In_338,In_302);
and U48 (N_48,In_1268,In_363);
or U49 (N_49,In_459,In_1193);
and U50 (N_50,In_1087,In_1129);
nand U51 (N_51,In_323,In_1092);
and U52 (N_52,In_893,In_1318);
nand U53 (N_53,In_1418,In_959);
nand U54 (N_54,In_1364,In_605);
or U55 (N_55,In_933,In_726);
and U56 (N_56,In_670,In_1447);
and U57 (N_57,In_251,In_108);
and U58 (N_58,In_417,In_1080);
nor U59 (N_59,In_1007,In_1140);
and U60 (N_60,In_262,In_738);
or U61 (N_61,In_164,In_548);
and U62 (N_62,In_1190,In_1333);
or U63 (N_63,In_988,In_604);
or U64 (N_64,In_1230,In_183);
or U65 (N_65,In_106,In_1187);
nor U66 (N_66,In_1275,In_297);
nand U67 (N_67,In_1085,In_1395);
nor U68 (N_68,In_135,In_237);
and U69 (N_69,In_1430,In_949);
nor U70 (N_70,In_1284,In_858);
nor U71 (N_71,In_36,In_936);
nand U72 (N_72,In_269,In_794);
or U73 (N_73,In_430,In_177);
or U74 (N_74,In_1200,In_919);
and U75 (N_75,In_275,In_450);
or U76 (N_76,In_1210,In_614);
nor U77 (N_77,In_838,In_1228);
nand U78 (N_78,In_303,In_600);
nor U79 (N_79,In_119,In_247);
and U80 (N_80,In_886,In_288);
and U81 (N_81,In_219,In_1495);
nor U82 (N_82,In_481,In_1043);
nand U83 (N_83,In_954,In_1308);
and U84 (N_84,In_1038,In_149);
nand U85 (N_85,In_1340,In_968);
or U86 (N_86,In_137,In_1478);
nor U87 (N_87,In_24,In_215);
nand U88 (N_88,In_728,In_622);
nand U89 (N_89,In_1104,In_734);
and U90 (N_90,In_1030,In_562);
nand U91 (N_91,In_889,In_740);
and U92 (N_92,In_655,In_747);
nor U93 (N_93,In_317,In_357);
and U94 (N_94,In_1352,In_653);
nand U95 (N_95,In_1154,In_235);
nor U96 (N_96,In_130,In_1482);
nand U97 (N_97,In_1471,In_117);
and U98 (N_98,In_1264,In_465);
or U99 (N_99,In_138,In_1397);
and U100 (N_100,In_1003,In_576);
nor U101 (N_101,In_383,In_525);
nand U102 (N_102,In_348,In_371);
nand U103 (N_103,In_236,In_85);
nand U104 (N_104,In_25,In_987);
or U105 (N_105,In_732,In_411);
nor U106 (N_106,In_290,In_115);
or U107 (N_107,In_579,In_438);
and U108 (N_108,In_482,In_1438);
nor U109 (N_109,In_1412,In_861);
nand U110 (N_110,In_326,In_829);
or U111 (N_111,In_697,In_1433);
nand U112 (N_112,In_603,In_792);
nand U113 (N_113,In_758,In_100);
nor U114 (N_114,In_40,In_577);
or U115 (N_115,In_755,In_714);
nor U116 (N_116,In_1484,In_360);
or U117 (N_117,In_754,In_346);
nor U118 (N_118,In_686,In_1209);
nor U119 (N_119,In_1253,In_1000);
and U120 (N_120,In_696,In_429);
nor U121 (N_121,In_776,In_150);
or U122 (N_122,In_559,In_1081);
and U123 (N_123,In_1105,In_1354);
or U124 (N_124,In_185,In_1226);
or U125 (N_125,In_1423,In_679);
or U126 (N_126,In_294,In_1199);
nand U127 (N_127,In_599,In_1);
nor U128 (N_128,In_356,In_502);
or U129 (N_129,In_229,In_1436);
nor U130 (N_130,In_496,In_370);
nand U131 (N_131,In_1071,In_173);
nor U132 (N_132,In_1464,In_1068);
nor U133 (N_133,In_478,In_1116);
nor U134 (N_134,In_394,In_890);
and U135 (N_135,In_1148,In_1274);
and U136 (N_136,In_1450,In_1054);
or U137 (N_137,In_56,In_101);
nand U138 (N_138,In_82,In_97);
nand U139 (N_139,In_1192,In_1335);
and U140 (N_140,In_1019,In_165);
nor U141 (N_141,In_684,In_1021);
or U142 (N_142,In_116,In_657);
or U143 (N_143,In_241,In_195);
and U144 (N_144,In_1048,In_989);
nand U145 (N_145,In_1330,In_915);
nand U146 (N_146,In_10,In_1291);
nor U147 (N_147,In_1262,In_547);
or U148 (N_148,In_1197,In_211);
and U149 (N_149,In_872,In_171);
nor U150 (N_150,In_86,In_956);
nand U151 (N_151,In_1133,In_95);
nor U152 (N_152,In_479,In_953);
or U153 (N_153,In_1329,In_174);
nand U154 (N_154,In_339,In_584);
nand U155 (N_155,In_176,In_524);
nand U156 (N_156,In_322,In_197);
or U157 (N_157,In_632,In_623);
and U158 (N_158,In_1220,In_843);
or U159 (N_159,In_292,In_445);
nand U160 (N_160,In_1298,In_980);
nand U161 (N_161,In_1132,In_648);
nor U162 (N_162,In_1234,In_282);
and U163 (N_163,In_1248,In_353);
nor U164 (N_164,In_1166,In_369);
nor U165 (N_165,In_220,In_4);
nor U166 (N_166,In_291,In_713);
nand U167 (N_167,In_1491,In_159);
and U168 (N_168,In_773,In_301);
nor U169 (N_169,In_1496,In_32);
nor U170 (N_170,In_1285,In_1117);
or U171 (N_171,In_1277,In_1444);
nor U172 (N_172,In_198,In_939);
xor U173 (N_173,In_66,In_1211);
and U174 (N_174,In_1305,In_464);
nand U175 (N_175,In_1128,In_1208);
nor U176 (N_176,In_1075,In_332);
or U177 (N_177,In_659,In_763);
nand U178 (N_178,In_422,In_488);
and U179 (N_179,In_700,In_1079);
and U180 (N_180,In_362,In_568);
nor U181 (N_181,In_1360,In_606);
nor U182 (N_182,In_725,In_818);
nor U183 (N_183,In_1257,In_1029);
and U184 (N_184,In_498,In_1316);
nor U185 (N_185,In_227,In_1205);
and U186 (N_186,In_539,In_413);
nor U187 (N_187,In_1022,In_1405);
nand U188 (N_188,In_1100,In_1259);
and U189 (N_189,In_515,In_333);
and U190 (N_190,In_389,In_358);
and U191 (N_191,In_231,In_567);
nor U192 (N_192,In_1366,In_80);
or U193 (N_193,In_293,In_830);
or U194 (N_194,In_639,In_162);
or U195 (N_195,In_678,In_1247);
and U196 (N_196,In_17,In_337);
nor U197 (N_197,In_1051,In_1281);
nand U198 (N_198,In_1474,In_1065);
or U199 (N_199,In_973,In_15);
nand U200 (N_200,In_1147,In_400);
or U201 (N_201,In_129,In_248);
and U202 (N_202,In_393,In_898);
nand U203 (N_203,In_1175,In_1098);
or U204 (N_204,In_349,In_268);
and U205 (N_205,In_273,In_947);
and U206 (N_206,In_503,In_991);
nand U207 (N_207,In_418,In_1015);
nand U208 (N_208,In_813,In_1347);
and U209 (N_209,In_312,In_1388);
nand U210 (N_210,In_1296,In_955);
nand U211 (N_211,In_1427,In_118);
nor U212 (N_212,In_1207,In_878);
nor U213 (N_213,In_190,In_1243);
or U214 (N_214,In_480,In_1490);
nor U215 (N_215,In_233,In_1153);
nand U216 (N_216,In_1074,In_771);
nor U217 (N_217,In_1458,In_1251);
nand U218 (N_218,In_1311,In_1044);
or U219 (N_219,In_1402,In_692);
nor U220 (N_220,In_376,In_801);
and U221 (N_221,In_1314,In_902);
and U222 (N_222,In_557,In_132);
or U223 (N_223,In_996,In_3);
or U224 (N_224,In_404,In_142);
and U225 (N_225,In_967,In_749);
or U226 (N_226,In_373,In_699);
nor U227 (N_227,In_263,In_140);
and U228 (N_228,In_1428,In_327);
nor U229 (N_229,In_1224,In_777);
and U230 (N_230,In_1096,In_1497);
and U231 (N_231,In_1178,In_1313);
or U232 (N_232,In_1486,In_1113);
nand U233 (N_233,In_267,In_1398);
or U234 (N_234,In_797,In_407);
and U235 (N_235,In_531,In_258);
and U236 (N_236,In_922,In_1045);
and U237 (N_237,In_463,In_1467);
or U238 (N_238,In_242,In_1103);
nor U239 (N_239,In_743,In_501);
nand U240 (N_240,In_1331,In_542);
and U241 (N_241,In_352,In_1244);
or U242 (N_242,In_1181,In_1472);
nand U243 (N_243,In_375,In_810);
or U244 (N_244,In_1173,In_181);
or U245 (N_245,In_1265,In_828);
or U246 (N_246,In_1269,In_457);
nor U247 (N_247,In_172,In_672);
nor U248 (N_248,In_1076,In_855);
nor U249 (N_249,In_228,In_611);
nor U250 (N_250,In_1499,In_455);
nand U251 (N_251,In_433,In_272);
and U252 (N_252,In_1287,In_673);
or U253 (N_253,In_1368,In_970);
nand U254 (N_254,In_588,In_128);
or U255 (N_255,In_1004,In_504);
and U256 (N_256,In_1442,In_497);
and U257 (N_257,In_803,In_184);
and U258 (N_258,In_124,In_102);
xor U259 (N_259,In_1312,In_826);
and U260 (N_260,In_1455,In_1037);
and U261 (N_261,In_1083,In_239);
nand U262 (N_262,In_1252,In_264);
nand U263 (N_263,In_681,In_308);
nand U264 (N_264,In_880,In_1214);
and U265 (N_265,In_683,In_1168);
nand U266 (N_266,In_1349,In_216);
nand U267 (N_267,In_134,In_721);
nand U268 (N_268,In_1407,In_79);
nand U269 (N_269,In_189,In_1169);
nand U270 (N_270,In_1151,In_638);
nand U271 (N_271,In_602,In_521);
nand U272 (N_272,In_597,In_1249);
nand U273 (N_273,In_39,In_156);
and U274 (N_274,In_1498,In_1115);
nand U275 (N_275,In_23,In_368);
nor U276 (N_276,In_1218,In_432);
and U277 (N_277,In_381,In_1334);
nand U278 (N_278,In_847,In_607);
or U279 (N_279,In_957,In_1439);
nor U280 (N_280,In_1245,In_549);
or U281 (N_281,In_105,In_1167);
or U282 (N_282,In_1231,In_1399);
nor U283 (N_283,In_753,In_1417);
nor U284 (N_284,In_296,In_981);
and U285 (N_285,In_836,In_83);
and U286 (N_286,In_409,In_330);
nor U287 (N_287,In_179,In_664);
nand U288 (N_288,In_601,In_1282);
nor U289 (N_289,In_440,In_27);
nand U290 (N_290,In_772,In_221);
and U291 (N_291,In_1172,In_578);
or U292 (N_292,In_716,In_1093);
or U293 (N_293,In_1196,In_656);
or U294 (N_294,In_1440,In_1090);
nor U295 (N_295,In_1124,In_234);
or U296 (N_296,In_737,In_712);
xor U297 (N_297,In_729,In_359);
and U298 (N_298,In_431,In_152);
nor U299 (N_299,In_477,In_103);
and U300 (N_300,In_1062,In_839);
nor U301 (N_301,In_693,In_201);
nand U302 (N_302,In_1363,In_703);
or U303 (N_303,In_852,In_690);
nor U304 (N_304,In_971,In_1483);
and U305 (N_305,In_666,In_89);
nor U306 (N_306,In_88,In_127);
or U307 (N_307,In_1369,In_840);
or U308 (N_308,In_627,In_123);
nand U309 (N_309,In_419,In_718);
nor U310 (N_310,In_978,In_1343);
and U311 (N_311,In_821,In_770);
nor U312 (N_312,In_64,In_68);
or U313 (N_313,In_1039,In_487);
nor U314 (N_314,In_731,In_1355);
or U315 (N_315,In_1002,In_437);
and U316 (N_316,In_928,In_1415);
or U317 (N_317,In_781,In_489);
and U318 (N_318,In_768,In_321);
nor U319 (N_319,In_1164,In_1088);
nand U320 (N_320,In_120,In_706);
or U321 (N_321,In_18,In_815);
nand U322 (N_322,In_448,In_555);
nand U323 (N_323,In_715,In_780);
and U324 (N_324,In_1221,In_1473);
nand U325 (N_325,In_1232,In_191);
nor U326 (N_326,In_154,In_590);
or U327 (N_327,In_110,In_845);
or U328 (N_328,In_81,In_287);
nand U329 (N_329,In_1323,In_1256);
nand U330 (N_330,In_1158,In_976);
and U331 (N_331,In_385,In_874);
nand U332 (N_332,In_1437,In_764);
nand U333 (N_333,In_424,In_904);
or U334 (N_334,In_518,In_879);
or U335 (N_335,In_952,In_1025);
nor U336 (N_336,In_563,In_461);
nor U337 (N_337,In_319,In_667);
nand U338 (N_338,In_551,In_921);
nor U339 (N_339,In_680,In_109);
nor U340 (N_340,In_748,In_942);
nor U341 (N_341,In_733,In_1459);
nand U342 (N_342,In_730,In_1141);
xnor U343 (N_343,In_669,In_943);
and U344 (N_344,In_1293,In_51);
and U345 (N_345,In_833,In_1320);
nor U346 (N_346,In_711,In_1149);
or U347 (N_347,In_1034,In_1390);
or U348 (N_348,In_428,In_336);
nand U349 (N_349,In_1082,In_1111);
and U350 (N_350,In_1014,In_997);
xnor U351 (N_351,In_938,In_194);
and U352 (N_352,In_899,In_449);
nor U353 (N_353,In_351,In_1136);
or U354 (N_354,In_649,In_380);
or U355 (N_355,In_929,In_1371);
nor U356 (N_356,In_14,In_1338);
or U357 (N_357,In_1219,In_122);
or U358 (N_358,In_366,In_798);
and U359 (N_359,In_1049,In_1258);
or U360 (N_360,In_661,In_552);
or U361 (N_361,In_1008,In_945);
and U362 (N_362,In_701,In_687);
nand U363 (N_363,In_155,In_253);
nand U364 (N_364,In_1317,In_1392);
nand U365 (N_365,In_1493,In_580);
and U366 (N_366,In_289,In_722);
or U367 (N_367,In_1449,In_1488);
nand U368 (N_368,In_841,In_1063);
nor U369 (N_369,In_6,In_903);
nor U370 (N_370,In_441,In_592);
nand U371 (N_371,In_529,In_628);
and U372 (N_372,In_742,In_779);
nor U373 (N_373,In_1260,In_77);
nor U374 (N_374,In_1078,In_811);
nand U375 (N_375,In_819,In_1011);
nand U376 (N_376,In_1070,In_1416);
nor U377 (N_377,In_250,In_1010);
or U378 (N_378,In_483,In_33);
nand U379 (N_379,In_1046,In_196);
nand U380 (N_380,In_677,In_367);
and U381 (N_381,In_1394,In_175);
and U382 (N_382,In_1289,In_1303);
or U383 (N_383,In_500,In_761);
or U384 (N_384,In_354,In_1067);
and U385 (N_385,In_254,In_388);
nand U386 (N_386,In_442,In_1077);
or U387 (N_387,In_470,In_284);
nor U388 (N_388,In_544,In_1072);
nor U389 (N_389,In_361,In_1227);
or U390 (N_390,In_894,In_1099);
or U391 (N_391,In_1123,In_1223);
or U392 (N_392,In_45,In_1386);
or U393 (N_393,In_1047,In_530);
xnor U394 (N_394,In_634,In_534);
and U395 (N_395,In_1194,In_374);
and U396 (N_396,In_643,In_918);
nor U397 (N_397,In_1475,In_186);
nand U398 (N_398,In_1485,In_993);
nor U399 (N_399,In_925,In_28);
and U400 (N_400,In_707,In_923);
nor U401 (N_401,In_435,In_1137);
nor U402 (N_402,In_618,In_695);
and U403 (N_403,In_8,In_111);
nand U404 (N_404,In_995,In_519);
nand U405 (N_405,In_416,In_1413);
and U406 (N_406,In_222,In_931);
nand U407 (N_407,In_741,In_1212);
or U408 (N_408,In_596,In_49);
and U409 (N_409,In_924,In_1299);
nor U410 (N_410,In_546,In_1406);
nor U411 (N_411,In_310,In_63);
and U412 (N_412,In_848,In_1066);
or U413 (N_413,In_279,In_1120);
nor U414 (N_414,In_856,In_286);
and U415 (N_415,In_585,In_565);
nand U416 (N_416,In_1382,In_905);
or U417 (N_417,In_1315,In_1201);
nor U418 (N_418,In_1185,In_161);
and U419 (N_419,In_144,In_613);
nand U420 (N_420,In_493,In_60);
and U421 (N_421,In_1143,In_1060);
nor U422 (N_422,In_57,In_1182);
nor U423 (N_423,In_1225,In_1381);
nor U424 (N_424,In_1135,In_864);
and U425 (N_425,In_1286,In_543);
nor U426 (N_426,In_2,In_1112);
nand U427 (N_427,In_589,In_1403);
nand U428 (N_428,In_1448,In_1018);
nor U429 (N_429,In_871,In_1091);
or U430 (N_430,In_554,In_1353);
and U431 (N_431,In_1242,In_1463);
and U432 (N_432,In_527,In_514);
nand U433 (N_433,In_1250,In_626);
or U434 (N_434,In_1465,In_762);
nor U435 (N_435,In_927,In_390);
nor U436 (N_436,In_932,In_456);
nor U437 (N_437,In_1306,In_1180);
nand U438 (N_438,In_240,In_11);
nor U439 (N_439,In_1184,In_671);
and U440 (N_440,In_93,In_1300);
and U441 (N_441,In_746,In_1036);
and U442 (N_442,In_491,In_1126);
or U443 (N_443,In_1122,In_454);
nand U444 (N_444,In_566,In_281);
and U445 (N_445,In_1393,In_1337);
nand U446 (N_446,In_1283,In_735);
and U447 (N_447,In_1146,In_966);
nor U448 (N_448,In_1276,In_1050);
and U449 (N_449,In_1064,In_1336);
and U450 (N_450,In_846,In_646);
and U451 (N_451,In_1237,In_1342);
or U452 (N_452,In_160,In_492);
or U453 (N_453,In_775,In_574);
nor U454 (N_454,In_331,In_884);
or U455 (N_455,In_1239,In_572);
nor U456 (N_456,In_1156,In_556);
nor U457 (N_457,In_969,In_636);
nor U458 (N_458,In_148,In_398);
nand U459 (N_459,In_7,In_277);
nor U460 (N_460,In_1152,In_796);
nand U461 (N_461,In_1443,In_355);
nand U462 (N_462,In_1150,In_877);
nor U463 (N_463,In_209,In_1053);
or U464 (N_464,In_169,In_98);
and U465 (N_465,In_76,In_965);
and U466 (N_466,In_788,In_9);
xnor U467 (N_467,In_13,In_342);
or U468 (N_468,In_270,In_126);
and U469 (N_469,In_736,In_202);
nor U470 (N_470,In_484,In_121);
nor U471 (N_471,In_842,In_787);
or U472 (N_472,In_46,In_506);
or U473 (N_473,In_674,In_87);
and U474 (N_474,In_1310,In_96);
or U475 (N_475,In_1125,In_665);
or U476 (N_476,In_1346,In_1032);
and U477 (N_477,In_125,In_507);
nor U478 (N_478,In_598,In_1452);
and U479 (N_479,In_245,In_1420);
nand U480 (N_480,In_1139,In_1453);
nand U481 (N_481,In_1468,In_1006);
and U482 (N_482,In_617,In_575);
nor U483 (N_483,In_537,In_425);
nor U484 (N_484,In_1059,In_187);
nand U485 (N_485,In_844,In_906);
nor U486 (N_486,In_789,In_1408);
or U487 (N_487,In_399,In_1101);
and U488 (N_488,In_682,In_345);
or U489 (N_489,In_1378,In_909);
or U490 (N_490,In_1365,In_641);
nand U491 (N_491,In_569,In_960);
and U492 (N_492,In_823,In_1422);
and U493 (N_493,In_467,In_964);
nor U494 (N_494,In_944,In_1055);
and U495 (N_495,In_1206,In_1052);
nand U496 (N_496,In_1142,In_986);
and U497 (N_497,In_570,In_52);
or U498 (N_498,In_1261,In_203);
nand U499 (N_499,In_571,In_1020);
and U500 (N_500,In_131,In_139);
nand U501 (N_501,In_631,In_283);
or U502 (N_502,In_912,In_1263);
and U503 (N_503,In_513,In_720);
and U504 (N_504,In_44,In_200);
or U505 (N_505,In_1107,In_421);
and U506 (N_506,In_466,In_512);
or U507 (N_507,In_974,In_582);
or U508 (N_508,In_1134,In_850);
or U509 (N_509,In_892,In_1138);
nor U510 (N_510,In_1216,In_1217);
nand U511 (N_511,In_414,In_188);
nand U512 (N_512,In_1387,In_1373);
and U513 (N_513,In_167,In_94);
nor U514 (N_514,In_560,In_54);
nor U515 (N_515,In_474,In_862);
and U516 (N_516,In_940,In_397);
nor U517 (N_517,In_1033,In_107);
nor U518 (N_518,In_913,In_1280);
nand U519 (N_519,In_50,In_553);
nor U520 (N_520,In_612,In_1255);
nor U521 (N_521,In_43,In_444);
nand U522 (N_522,In_1238,In_69);
or U523 (N_523,In_564,In_1307);
or U524 (N_524,In_561,In_55);
nor U525 (N_525,In_212,In_37);
and U526 (N_526,In_897,In_727);
and U527 (N_527,In_1241,In_315);
nor U528 (N_528,In_757,In_832);
nand U529 (N_529,In_1400,In_328);
nand U530 (N_530,In_387,In_1328);
or U531 (N_531,In_647,In_451);
and U532 (N_532,In_1414,In_70);
and U533 (N_533,In_535,In_1295);
nand U534 (N_534,In_1106,In_752);
nand U535 (N_535,In_1012,In_688);
nor U536 (N_536,In_637,In_750);
and U537 (N_537,In_594,In_91);
nor U538 (N_538,In_875,In_490);
or U539 (N_539,In_340,In_1380);
nor U540 (N_540,In_868,In_528);
or U541 (N_541,In_1367,In_392);
nand U542 (N_542,In_831,In_1339);
or U543 (N_543,In_395,In_208);
or U544 (N_544,In_382,In_972);
or U545 (N_545,In_807,In_249);
nand U546 (N_546,In_710,In_0);
nor U547 (N_547,In_694,In_1095);
and U548 (N_548,In_213,In_460);
nor U549 (N_549,In_1351,In_824);
or U550 (N_550,In_888,In_1023);
or U551 (N_551,In_951,In_1419);
or U552 (N_552,In_226,In_1345);
and U553 (N_553,In_379,In_257);
nor U554 (N_554,In_469,In_885);
and U555 (N_555,In_217,In_462);
nor U556 (N_556,In_1376,In_1042);
nor U557 (N_557,In_1177,In_1094);
or U558 (N_558,In_278,In_1161);
or U559 (N_559,In_1058,In_907);
nand U560 (N_560,In_896,In_1017);
nand U561 (N_561,In_963,In_1396);
nand U562 (N_562,In_859,In_795);
nand U563 (N_563,In_1170,In_1466);
nor U564 (N_564,In_538,In_958);
or U565 (N_565,In_869,In_541);
and U566 (N_566,In_1026,In_802);
nor U567 (N_567,In_790,In_1429);
nor U568 (N_568,In_274,In_992);
nor U569 (N_569,In_295,In_1456);
or U570 (N_570,In_778,In_1374);
and U571 (N_571,In_163,In_1479);
or U572 (N_572,In_42,In_934);
or U573 (N_573,In_1031,In_808);
nand U574 (N_574,In_298,In_654);
nor U575 (N_575,In_406,In_853);
and U576 (N_576,In_1073,In_522);
nor U577 (N_577,In_591,In_774);
or U578 (N_578,In_396,In_516);
nor U579 (N_579,In_48,In_1476);
or U580 (N_580,In_1451,In_1421);
nand U581 (N_581,In_72,In_1357);
nor U582 (N_582,In_157,In_12);
nor U583 (N_583,In_717,In_1040);
nand U584 (N_584,In_59,In_311);
nand U585 (N_585,In_114,In_1183);
and U586 (N_586,In_1155,In_1041);
nand U587 (N_587,In_324,In_1270);
nand U588 (N_588,In_22,In_1469);
and U589 (N_589,In_329,In_1401);
and U590 (N_590,In_472,In_113);
nor U591 (N_591,In_1431,In_756);
nor U592 (N_592,In_1131,In_147);
nor U593 (N_593,In_252,In_914);
nor U594 (N_594,In_1273,In_533);
and U595 (N_595,In_1359,In_67);
or U596 (N_596,In_1024,In_473);
nand U597 (N_597,In_900,In_545);
or U598 (N_598,In_53,In_452);
or U599 (N_599,In_908,In_1198);
nor U600 (N_600,In_238,In_508);
nand U601 (N_601,In_31,In_485);
or U602 (N_602,In_881,In_146);
xnor U603 (N_603,In_887,In_583);
nand U604 (N_604,In_1163,In_1383);
and U605 (N_605,In_1278,In_926);
or U606 (N_606,In_509,In_1385);
nor U607 (N_607,In_793,In_41);
and U608 (N_608,In_1361,In_265);
and U609 (N_609,In_35,In_526);
or U610 (N_610,In_505,In_891);
and U611 (N_611,In_1157,In_20);
or U612 (N_612,In_835,In_1267);
or U613 (N_613,In_1409,In_608);
or U614 (N_614,In_739,In_1341);
and U615 (N_615,In_224,In_917);
and U616 (N_616,In_30,In_204);
nor U617 (N_617,In_158,In_447);
nand U618 (N_618,In_1358,In_259);
nand U619 (N_619,In_1191,In_1302);
and U620 (N_620,In_975,In_434);
nand U621 (N_621,In_1057,In_1171);
nor U622 (N_622,In_1119,In_168);
or U623 (N_623,In_883,In_1379);
nand U624 (N_624,In_47,In_1441);
nor U625 (N_625,In_350,In_948);
nand U626 (N_626,In_1324,In_1165);
nor U627 (N_627,In_471,In_1372);
and U628 (N_628,In_620,In_1061);
and U629 (N_629,In_827,In_260);
nand U630 (N_630,In_1240,In_619);
nand U631 (N_631,In_911,In_979);
or U632 (N_632,In_882,In_1301);
nand U633 (N_633,In_994,In_1288);
and U634 (N_634,In_378,In_99);
and U635 (N_635,In_1179,In_1272);
and U636 (N_636,In_1222,In_523);
nor U637 (N_637,In_225,In_593);
nand U638 (N_638,In_1056,In_261);
and U639 (N_639,In_391,In_624);
nor U640 (N_640,In_935,In_685);
and U641 (N_641,In_1102,In_180);
and U642 (N_642,In_709,In_29);
nor U643 (N_643,In_1114,In_1233);
nor U644 (N_644,In_704,In_316);
nand U645 (N_645,In_660,In_676);
and U646 (N_646,In_1144,In_962);
xor U647 (N_647,In_494,In_635);
nand U648 (N_648,In_920,In_1246);
nor U649 (N_649,In_423,In_313);
nor U650 (N_650,In_305,In_344);
nor U651 (N_651,In_645,In_1389);
nand U652 (N_652,In_1477,In_1229);
or U653 (N_653,In_214,In_1145);
or U654 (N_654,In_71,In_805);
nor U655 (N_655,In_486,In_961);
nor U656 (N_656,In_285,In_937);
and U657 (N_657,In_439,In_1322);
nor U658 (N_658,In_499,In_766);
nor U659 (N_659,In_1069,In_1356);
nand U660 (N_660,In_866,In_58);
nand U661 (N_661,In_640,In_1344);
and U662 (N_662,In_1086,In_817);
and U663 (N_663,In_1462,In_170);
or U664 (N_664,In_1266,In_420);
nor U665 (N_665,In_1162,In_384);
and U666 (N_666,In_999,In_1294);
nor U667 (N_667,In_1290,In_785);
nor U668 (N_668,In_16,In_1271);
or U669 (N_669,In_112,In_495);
nand U670 (N_670,In_244,In_1470);
nor U671 (N_671,In_341,In_304);
nor U672 (N_672,In_38,In_133);
nor U673 (N_673,In_1391,In_401);
or U674 (N_674,In_1279,In_1321);
nand U675 (N_675,In_1186,In_314);
nand U676 (N_676,In_825,In_143);
nor U677 (N_677,In_1118,In_1489);
or U678 (N_678,In_702,In_458);
and U679 (N_679,In_998,In_1110);
nor U680 (N_680,In_1425,In_307);
and U681 (N_681,In_510,In_650);
nand U682 (N_682,In_62,In_280);
and U683 (N_683,In_536,In_540);
and U684 (N_684,In_837,In_698);
and U685 (N_685,In_1445,In_412);
or U686 (N_686,In_1410,In_550);
and U687 (N_687,In_136,In_691);
nor U688 (N_688,In_1370,In_916);
and U689 (N_689,In_719,In_860);
or U690 (N_690,In_724,In_218);
nand U691 (N_691,In_642,In_223);
or U692 (N_692,In_786,In_403);
nor U693 (N_693,In_1375,In_910);
nand U694 (N_694,In_182,In_153);
nor U695 (N_695,In_1254,In_246);
nor U696 (N_696,In_206,In_65);
and U697 (N_697,In_1492,In_532);
nor U698 (N_698,In_982,In_1404);
nor U699 (N_699,In_1174,In_405);
and U700 (N_700,In_1027,In_1001);
nand U701 (N_701,In_1348,In_1121);
nor U702 (N_702,In_386,In_1480);
and U703 (N_703,In_629,In_851);
and U704 (N_704,In_347,In_791);
and U705 (N_705,In_1202,In_800);
or U706 (N_706,In_1235,In_1332);
nand U707 (N_707,In_595,In_92);
or U708 (N_708,In_723,In_320);
or U709 (N_709,In_446,In_581);
or U710 (N_710,In_5,In_783);
nor U711 (N_711,In_857,In_616);
and U712 (N_712,In_334,In_372);
or U713 (N_713,In_941,In_950);
nor U714 (N_714,In_1432,In_930);
nor U715 (N_715,In_689,In_436);
nand U716 (N_716,In_1005,In_1460);
and U717 (N_717,In_1304,In_812);
nand U718 (N_718,In_271,In_814);
and U719 (N_719,In_610,In_1203);
nor U720 (N_720,In_873,In_325);
or U721 (N_721,In_1109,In_207);
nor U722 (N_722,In_977,In_1130);
nor U723 (N_723,In_276,In_377);
and U724 (N_724,In_615,In_1362);
nand U725 (N_725,In_651,In_895);
nor U726 (N_726,In_26,In_1159);
nor U727 (N_727,In_870,In_587);
nor U728 (N_728,In_19,In_1009);
or U729 (N_729,In_1204,In_1108);
nand U730 (N_730,In_104,In_243);
xor U731 (N_731,In_1236,In_586);
xor U732 (N_732,In_990,In_443);
or U733 (N_733,In_767,In_745);
and U734 (N_734,In_1319,In_809);
and U735 (N_735,In_335,In_78);
nor U736 (N_736,In_426,In_1127);
nand U737 (N_737,In_984,In_141);
nor U738 (N_738,In_75,In_863);
nand U739 (N_739,In_1176,In_668);
nand U740 (N_740,In_318,In_210);
nor U741 (N_741,In_300,In_1411);
or U742 (N_742,In_1297,In_364);
nand U743 (N_743,In_1215,In_621);
nor U744 (N_744,In_306,In_822);
nor U745 (N_745,In_834,In_475);
nor U746 (N_746,In_1350,In_760);
and U747 (N_747,In_867,In_255);
or U748 (N_748,In_644,In_427);
or U749 (N_749,In_84,In_266);
nor U750 (N_750,In_722,In_1338);
nor U751 (N_751,In_328,In_1431);
nor U752 (N_752,In_1470,In_974);
and U753 (N_753,In_43,In_647);
and U754 (N_754,In_869,In_892);
nand U755 (N_755,In_891,In_83);
nor U756 (N_756,In_1307,In_244);
nor U757 (N_757,In_1415,In_1264);
nand U758 (N_758,In_641,In_464);
or U759 (N_759,In_1190,In_555);
and U760 (N_760,In_900,In_1022);
or U761 (N_761,In_1229,In_904);
and U762 (N_762,In_1059,In_1172);
nor U763 (N_763,In_233,In_3);
nand U764 (N_764,In_683,In_542);
nand U765 (N_765,In_1227,In_666);
nor U766 (N_766,In_877,In_101);
and U767 (N_767,In_484,In_123);
or U768 (N_768,In_1243,In_998);
nand U769 (N_769,In_330,In_1372);
and U770 (N_770,In_334,In_1139);
or U771 (N_771,In_780,In_1259);
and U772 (N_772,In_291,In_401);
and U773 (N_773,In_549,In_29);
or U774 (N_774,In_1320,In_917);
nand U775 (N_775,In_1499,In_432);
or U776 (N_776,In_1165,In_1147);
or U777 (N_777,In_1170,In_1241);
and U778 (N_778,In_922,In_602);
or U779 (N_779,In_17,In_935);
nor U780 (N_780,In_1069,In_282);
or U781 (N_781,In_443,In_1219);
or U782 (N_782,In_96,In_308);
nand U783 (N_783,In_517,In_143);
xor U784 (N_784,In_75,In_725);
nor U785 (N_785,In_1046,In_243);
and U786 (N_786,In_440,In_1081);
nor U787 (N_787,In_1056,In_1205);
nor U788 (N_788,In_548,In_454);
nor U789 (N_789,In_1410,In_544);
or U790 (N_790,In_166,In_1396);
nor U791 (N_791,In_101,In_1055);
or U792 (N_792,In_345,In_561);
or U793 (N_793,In_1229,In_687);
or U794 (N_794,In_579,In_1352);
nor U795 (N_795,In_722,In_282);
and U796 (N_796,In_1430,In_526);
nor U797 (N_797,In_164,In_495);
nand U798 (N_798,In_714,In_12);
nor U799 (N_799,In_683,In_1042);
or U800 (N_800,In_241,In_950);
nand U801 (N_801,In_1485,In_1050);
nand U802 (N_802,In_1171,In_484);
or U803 (N_803,In_1023,In_1229);
nand U804 (N_804,In_1448,In_341);
nor U805 (N_805,In_1248,In_494);
nor U806 (N_806,In_796,In_1438);
nor U807 (N_807,In_757,In_1108);
nor U808 (N_808,In_659,In_18);
nor U809 (N_809,In_29,In_150);
nor U810 (N_810,In_1072,In_1207);
nor U811 (N_811,In_727,In_1241);
or U812 (N_812,In_858,In_1278);
and U813 (N_813,In_403,In_1078);
nor U814 (N_814,In_1381,In_1181);
nor U815 (N_815,In_208,In_1410);
and U816 (N_816,In_1325,In_80);
or U817 (N_817,In_1205,In_966);
or U818 (N_818,In_96,In_847);
or U819 (N_819,In_766,In_681);
nor U820 (N_820,In_1384,In_121);
nand U821 (N_821,In_864,In_1348);
and U822 (N_822,In_152,In_71);
nand U823 (N_823,In_313,In_1432);
nor U824 (N_824,In_509,In_1245);
and U825 (N_825,In_1260,In_347);
and U826 (N_826,In_1348,In_683);
nand U827 (N_827,In_1121,In_513);
or U828 (N_828,In_121,In_1398);
and U829 (N_829,In_1129,In_1193);
or U830 (N_830,In_694,In_985);
or U831 (N_831,In_570,In_408);
nor U832 (N_832,In_1374,In_267);
nand U833 (N_833,In_1343,In_160);
and U834 (N_834,In_883,In_1427);
or U835 (N_835,In_1336,In_1031);
or U836 (N_836,In_371,In_210);
nand U837 (N_837,In_552,In_821);
nor U838 (N_838,In_433,In_588);
and U839 (N_839,In_967,In_1484);
nor U840 (N_840,In_183,In_795);
or U841 (N_841,In_1292,In_282);
nor U842 (N_842,In_771,In_1060);
nor U843 (N_843,In_324,In_940);
and U844 (N_844,In_1420,In_727);
and U845 (N_845,In_223,In_235);
or U846 (N_846,In_1251,In_146);
or U847 (N_847,In_1058,In_287);
nand U848 (N_848,In_1290,In_242);
nor U849 (N_849,In_105,In_1128);
and U850 (N_850,In_1030,In_1133);
and U851 (N_851,In_304,In_748);
nor U852 (N_852,In_726,In_1078);
or U853 (N_853,In_1196,In_1269);
and U854 (N_854,In_1281,In_160);
nand U855 (N_855,In_1443,In_859);
nor U856 (N_856,In_478,In_1062);
and U857 (N_857,In_630,In_497);
or U858 (N_858,In_1117,In_202);
nand U859 (N_859,In_270,In_5);
nor U860 (N_860,In_489,In_421);
nor U861 (N_861,In_1386,In_249);
or U862 (N_862,In_1105,In_1192);
or U863 (N_863,In_111,In_1480);
nand U864 (N_864,In_790,In_948);
xor U865 (N_865,In_1435,In_39);
or U866 (N_866,In_939,In_112);
and U867 (N_867,In_557,In_709);
nand U868 (N_868,In_221,In_842);
nor U869 (N_869,In_863,In_659);
and U870 (N_870,In_187,In_260);
nor U871 (N_871,In_1481,In_571);
xnor U872 (N_872,In_822,In_265);
nand U873 (N_873,In_1305,In_407);
or U874 (N_874,In_86,In_121);
nand U875 (N_875,In_840,In_1154);
nor U876 (N_876,In_69,In_1389);
or U877 (N_877,In_279,In_715);
nand U878 (N_878,In_1155,In_1081);
nand U879 (N_879,In_1186,In_1407);
nand U880 (N_880,In_295,In_397);
nand U881 (N_881,In_672,In_212);
or U882 (N_882,In_847,In_616);
and U883 (N_883,In_324,In_1456);
nand U884 (N_884,In_330,In_802);
and U885 (N_885,In_641,In_730);
or U886 (N_886,In_798,In_216);
or U887 (N_887,In_460,In_913);
nand U888 (N_888,In_1215,In_595);
nor U889 (N_889,In_1068,In_752);
nand U890 (N_890,In_975,In_63);
or U891 (N_891,In_426,In_192);
or U892 (N_892,In_173,In_517);
and U893 (N_893,In_295,In_1221);
nand U894 (N_894,In_68,In_1272);
and U895 (N_895,In_1073,In_1420);
nand U896 (N_896,In_1377,In_946);
or U897 (N_897,In_754,In_168);
nand U898 (N_898,In_139,In_378);
nor U899 (N_899,In_1287,In_1012);
and U900 (N_900,In_1171,In_1049);
and U901 (N_901,In_1370,In_467);
and U902 (N_902,In_992,In_425);
and U903 (N_903,In_1393,In_854);
and U904 (N_904,In_1393,In_990);
nor U905 (N_905,In_1369,In_95);
and U906 (N_906,In_909,In_1396);
and U907 (N_907,In_288,In_1200);
nand U908 (N_908,In_1294,In_412);
nand U909 (N_909,In_431,In_348);
xnor U910 (N_910,In_621,In_530);
nor U911 (N_911,In_1399,In_249);
and U912 (N_912,In_968,In_80);
or U913 (N_913,In_1358,In_881);
nor U914 (N_914,In_512,In_514);
nand U915 (N_915,In_141,In_1087);
and U916 (N_916,In_1160,In_675);
or U917 (N_917,In_495,In_1310);
nand U918 (N_918,In_528,In_121);
or U919 (N_919,In_854,In_786);
and U920 (N_920,In_1030,In_981);
or U921 (N_921,In_536,In_447);
and U922 (N_922,In_475,In_1197);
or U923 (N_923,In_252,In_1096);
or U924 (N_924,In_176,In_1021);
and U925 (N_925,In_142,In_1426);
and U926 (N_926,In_174,In_438);
nor U927 (N_927,In_259,In_584);
nand U928 (N_928,In_841,In_392);
nor U929 (N_929,In_311,In_701);
or U930 (N_930,In_1144,In_1181);
and U931 (N_931,In_259,In_1077);
or U932 (N_932,In_1219,In_1484);
and U933 (N_933,In_1244,In_1287);
and U934 (N_934,In_555,In_681);
nand U935 (N_935,In_648,In_563);
nand U936 (N_936,In_1417,In_423);
or U937 (N_937,In_76,In_1034);
and U938 (N_938,In_1213,In_762);
and U939 (N_939,In_897,In_729);
nand U940 (N_940,In_348,In_535);
or U941 (N_941,In_1048,In_298);
nor U942 (N_942,In_1161,In_353);
or U943 (N_943,In_631,In_919);
and U944 (N_944,In_496,In_737);
nand U945 (N_945,In_1006,In_1170);
nor U946 (N_946,In_447,In_445);
and U947 (N_947,In_549,In_493);
nor U948 (N_948,In_90,In_717);
nand U949 (N_949,In_1427,In_1375);
nand U950 (N_950,In_469,In_385);
or U951 (N_951,In_537,In_1349);
nor U952 (N_952,In_669,In_316);
or U953 (N_953,In_122,In_653);
and U954 (N_954,In_908,In_257);
or U955 (N_955,In_350,In_472);
and U956 (N_956,In_5,In_1301);
nor U957 (N_957,In_910,In_788);
and U958 (N_958,In_561,In_1214);
nor U959 (N_959,In_1255,In_1315);
nor U960 (N_960,In_1153,In_572);
and U961 (N_961,In_1373,In_1178);
nand U962 (N_962,In_998,In_657);
nand U963 (N_963,In_1398,In_201);
or U964 (N_964,In_1394,In_1147);
and U965 (N_965,In_54,In_1192);
nor U966 (N_966,In_1453,In_321);
nand U967 (N_967,In_320,In_1002);
nand U968 (N_968,In_543,In_1005);
nand U969 (N_969,In_751,In_947);
nand U970 (N_970,In_1326,In_547);
and U971 (N_971,In_113,In_409);
or U972 (N_972,In_668,In_364);
nand U973 (N_973,In_509,In_1204);
or U974 (N_974,In_590,In_1293);
nor U975 (N_975,In_1147,In_1142);
or U976 (N_976,In_1249,In_1423);
nand U977 (N_977,In_154,In_257);
and U978 (N_978,In_215,In_1212);
nor U979 (N_979,In_1245,In_1492);
nor U980 (N_980,In_890,In_196);
nand U981 (N_981,In_204,In_408);
nand U982 (N_982,In_783,In_415);
and U983 (N_983,In_1441,In_1100);
and U984 (N_984,In_820,In_677);
nand U985 (N_985,In_1312,In_1230);
or U986 (N_986,In_1369,In_656);
or U987 (N_987,In_794,In_1183);
or U988 (N_988,In_772,In_481);
nand U989 (N_989,In_247,In_709);
nand U990 (N_990,In_748,In_1098);
nor U991 (N_991,In_987,In_408);
and U992 (N_992,In_758,In_1488);
or U993 (N_993,In_203,In_1416);
or U994 (N_994,In_1419,In_9);
or U995 (N_995,In_1082,In_1063);
or U996 (N_996,In_1146,In_920);
nor U997 (N_997,In_186,In_938);
nand U998 (N_998,In_439,In_1028);
nand U999 (N_999,In_181,In_1198);
or U1000 (N_1000,In_68,In_1093);
nor U1001 (N_1001,In_98,In_1290);
and U1002 (N_1002,In_73,In_835);
nand U1003 (N_1003,In_147,In_13);
and U1004 (N_1004,In_897,In_1368);
or U1005 (N_1005,In_549,In_1156);
nand U1006 (N_1006,In_778,In_1313);
nand U1007 (N_1007,In_1166,In_13);
nor U1008 (N_1008,In_491,In_1116);
nor U1009 (N_1009,In_695,In_57);
nand U1010 (N_1010,In_925,In_770);
nand U1011 (N_1011,In_765,In_1022);
nand U1012 (N_1012,In_1491,In_554);
nand U1013 (N_1013,In_611,In_1170);
nand U1014 (N_1014,In_872,In_89);
nor U1015 (N_1015,In_227,In_336);
nor U1016 (N_1016,In_698,In_1217);
nand U1017 (N_1017,In_785,In_168);
or U1018 (N_1018,In_683,In_90);
or U1019 (N_1019,In_108,In_601);
nor U1020 (N_1020,In_1045,In_785);
nor U1021 (N_1021,In_1144,In_539);
nand U1022 (N_1022,In_680,In_604);
or U1023 (N_1023,In_437,In_616);
nand U1024 (N_1024,In_646,In_825);
nand U1025 (N_1025,In_607,In_741);
or U1026 (N_1026,In_1177,In_285);
nor U1027 (N_1027,In_1140,In_21);
and U1028 (N_1028,In_458,In_857);
nor U1029 (N_1029,In_766,In_88);
or U1030 (N_1030,In_825,In_954);
or U1031 (N_1031,In_539,In_1125);
or U1032 (N_1032,In_868,In_359);
or U1033 (N_1033,In_403,In_1486);
and U1034 (N_1034,In_641,In_903);
nand U1035 (N_1035,In_499,In_1078);
nand U1036 (N_1036,In_154,In_741);
nor U1037 (N_1037,In_399,In_43);
or U1038 (N_1038,In_1188,In_468);
and U1039 (N_1039,In_31,In_349);
nand U1040 (N_1040,In_369,In_1158);
or U1041 (N_1041,In_213,In_612);
nand U1042 (N_1042,In_558,In_301);
nand U1043 (N_1043,In_536,In_1499);
or U1044 (N_1044,In_263,In_1239);
or U1045 (N_1045,In_72,In_829);
nand U1046 (N_1046,In_1288,In_723);
and U1047 (N_1047,In_737,In_306);
nand U1048 (N_1048,In_839,In_492);
or U1049 (N_1049,In_1150,In_53);
or U1050 (N_1050,In_370,In_940);
or U1051 (N_1051,In_1470,In_74);
and U1052 (N_1052,In_1191,In_581);
or U1053 (N_1053,In_1124,In_1437);
nor U1054 (N_1054,In_1302,In_1461);
nor U1055 (N_1055,In_156,In_673);
and U1056 (N_1056,In_1207,In_612);
nand U1057 (N_1057,In_813,In_520);
nor U1058 (N_1058,In_424,In_847);
nor U1059 (N_1059,In_1129,In_1481);
or U1060 (N_1060,In_72,In_1076);
or U1061 (N_1061,In_991,In_1150);
or U1062 (N_1062,In_16,In_1366);
nor U1063 (N_1063,In_338,In_574);
nand U1064 (N_1064,In_231,In_1073);
or U1065 (N_1065,In_299,In_951);
and U1066 (N_1066,In_518,In_358);
and U1067 (N_1067,In_438,In_11);
or U1068 (N_1068,In_1459,In_1158);
and U1069 (N_1069,In_446,In_803);
or U1070 (N_1070,In_672,In_779);
nand U1071 (N_1071,In_104,In_1404);
nor U1072 (N_1072,In_514,In_861);
nand U1073 (N_1073,In_1165,In_515);
nand U1074 (N_1074,In_1186,In_93);
or U1075 (N_1075,In_392,In_1491);
nand U1076 (N_1076,In_374,In_1048);
nand U1077 (N_1077,In_727,In_1368);
nor U1078 (N_1078,In_437,In_290);
or U1079 (N_1079,In_1485,In_534);
or U1080 (N_1080,In_237,In_1409);
or U1081 (N_1081,In_177,In_744);
nand U1082 (N_1082,In_195,In_757);
or U1083 (N_1083,In_139,In_841);
and U1084 (N_1084,In_1389,In_1299);
or U1085 (N_1085,In_147,In_958);
nor U1086 (N_1086,In_404,In_152);
xnor U1087 (N_1087,In_119,In_686);
or U1088 (N_1088,In_1064,In_1257);
xor U1089 (N_1089,In_1369,In_1016);
nand U1090 (N_1090,In_748,In_1163);
or U1091 (N_1091,In_11,In_1302);
and U1092 (N_1092,In_249,In_1044);
and U1093 (N_1093,In_1417,In_381);
or U1094 (N_1094,In_423,In_1211);
nor U1095 (N_1095,In_331,In_1142);
or U1096 (N_1096,In_203,In_374);
or U1097 (N_1097,In_1433,In_1298);
and U1098 (N_1098,In_1459,In_470);
and U1099 (N_1099,In_585,In_680);
nor U1100 (N_1100,In_862,In_538);
nor U1101 (N_1101,In_916,In_390);
nor U1102 (N_1102,In_1013,In_1250);
or U1103 (N_1103,In_1270,In_1273);
nor U1104 (N_1104,In_539,In_935);
nand U1105 (N_1105,In_1393,In_1124);
nor U1106 (N_1106,In_283,In_442);
or U1107 (N_1107,In_979,In_380);
or U1108 (N_1108,In_643,In_156);
or U1109 (N_1109,In_1330,In_1023);
and U1110 (N_1110,In_1305,In_1066);
and U1111 (N_1111,In_500,In_310);
nand U1112 (N_1112,In_154,In_79);
nand U1113 (N_1113,In_1121,In_1054);
and U1114 (N_1114,In_856,In_1309);
nand U1115 (N_1115,In_1403,In_1358);
nand U1116 (N_1116,In_632,In_1201);
or U1117 (N_1117,In_521,In_469);
nand U1118 (N_1118,In_1080,In_534);
and U1119 (N_1119,In_1177,In_1128);
nor U1120 (N_1120,In_533,In_982);
and U1121 (N_1121,In_1374,In_36);
or U1122 (N_1122,In_931,In_848);
and U1123 (N_1123,In_1173,In_1267);
xnor U1124 (N_1124,In_757,In_1064);
nand U1125 (N_1125,In_913,In_103);
nand U1126 (N_1126,In_818,In_826);
or U1127 (N_1127,In_1456,In_539);
nor U1128 (N_1128,In_1077,In_179);
nand U1129 (N_1129,In_1101,In_563);
nor U1130 (N_1130,In_1019,In_364);
or U1131 (N_1131,In_178,In_1427);
nor U1132 (N_1132,In_167,In_1436);
nor U1133 (N_1133,In_1441,In_970);
nand U1134 (N_1134,In_109,In_990);
or U1135 (N_1135,In_169,In_444);
nand U1136 (N_1136,In_462,In_39);
or U1137 (N_1137,In_922,In_195);
and U1138 (N_1138,In_933,In_1355);
nand U1139 (N_1139,In_484,In_189);
nor U1140 (N_1140,In_1312,In_657);
and U1141 (N_1141,In_1355,In_1094);
and U1142 (N_1142,In_1034,In_1171);
nand U1143 (N_1143,In_578,In_748);
or U1144 (N_1144,In_779,In_224);
nor U1145 (N_1145,In_819,In_585);
or U1146 (N_1146,In_175,In_1041);
or U1147 (N_1147,In_241,In_1140);
or U1148 (N_1148,In_358,In_82);
nand U1149 (N_1149,In_164,In_99);
and U1150 (N_1150,In_756,In_740);
and U1151 (N_1151,In_1200,In_85);
nand U1152 (N_1152,In_1301,In_368);
nor U1153 (N_1153,In_157,In_359);
and U1154 (N_1154,In_106,In_1131);
nor U1155 (N_1155,In_1255,In_110);
or U1156 (N_1156,In_340,In_354);
and U1157 (N_1157,In_361,In_98);
nor U1158 (N_1158,In_444,In_1077);
or U1159 (N_1159,In_487,In_145);
nor U1160 (N_1160,In_204,In_1142);
nand U1161 (N_1161,In_797,In_984);
nor U1162 (N_1162,In_688,In_300);
nand U1163 (N_1163,In_701,In_626);
nor U1164 (N_1164,In_1363,In_1312);
nand U1165 (N_1165,In_1081,In_1097);
nand U1166 (N_1166,In_596,In_390);
nand U1167 (N_1167,In_421,In_335);
and U1168 (N_1168,In_994,In_1055);
or U1169 (N_1169,In_1052,In_653);
nor U1170 (N_1170,In_245,In_574);
and U1171 (N_1171,In_598,In_466);
and U1172 (N_1172,In_5,In_940);
nor U1173 (N_1173,In_657,In_1369);
and U1174 (N_1174,In_258,In_69);
and U1175 (N_1175,In_1218,In_225);
and U1176 (N_1176,In_1029,In_729);
nor U1177 (N_1177,In_1425,In_301);
nor U1178 (N_1178,In_1468,In_397);
nand U1179 (N_1179,In_279,In_1280);
nor U1180 (N_1180,In_898,In_674);
or U1181 (N_1181,In_1434,In_291);
and U1182 (N_1182,In_454,In_574);
or U1183 (N_1183,In_38,In_104);
nand U1184 (N_1184,In_1159,In_1384);
nor U1185 (N_1185,In_1010,In_1412);
and U1186 (N_1186,In_1484,In_1453);
or U1187 (N_1187,In_1154,In_16);
and U1188 (N_1188,In_542,In_1356);
nor U1189 (N_1189,In_401,In_816);
or U1190 (N_1190,In_895,In_1208);
or U1191 (N_1191,In_1496,In_1473);
or U1192 (N_1192,In_16,In_1051);
nor U1193 (N_1193,In_233,In_568);
and U1194 (N_1194,In_1216,In_1215);
nor U1195 (N_1195,In_509,In_437);
or U1196 (N_1196,In_312,In_95);
nor U1197 (N_1197,In_99,In_230);
nand U1198 (N_1198,In_260,In_212);
and U1199 (N_1199,In_483,In_945);
nand U1200 (N_1200,In_398,In_528);
or U1201 (N_1201,In_1266,In_831);
and U1202 (N_1202,In_985,In_469);
and U1203 (N_1203,In_1122,In_1473);
nor U1204 (N_1204,In_444,In_952);
nand U1205 (N_1205,In_369,In_241);
or U1206 (N_1206,In_1433,In_424);
and U1207 (N_1207,In_343,In_270);
nand U1208 (N_1208,In_1200,In_673);
nand U1209 (N_1209,In_1322,In_722);
or U1210 (N_1210,In_539,In_859);
or U1211 (N_1211,In_1289,In_1120);
and U1212 (N_1212,In_351,In_1257);
and U1213 (N_1213,In_1087,In_1376);
nor U1214 (N_1214,In_347,In_1257);
or U1215 (N_1215,In_860,In_652);
nor U1216 (N_1216,In_645,In_1191);
xor U1217 (N_1217,In_1417,In_462);
or U1218 (N_1218,In_786,In_546);
nor U1219 (N_1219,In_952,In_860);
nand U1220 (N_1220,In_714,In_800);
nand U1221 (N_1221,In_816,In_395);
nand U1222 (N_1222,In_527,In_1020);
nand U1223 (N_1223,In_1203,In_547);
nor U1224 (N_1224,In_1101,In_20);
nor U1225 (N_1225,In_582,In_735);
nand U1226 (N_1226,In_944,In_1277);
and U1227 (N_1227,In_289,In_1073);
nor U1228 (N_1228,In_114,In_1179);
or U1229 (N_1229,In_421,In_1488);
nand U1230 (N_1230,In_926,In_891);
and U1231 (N_1231,In_483,In_1126);
nand U1232 (N_1232,In_144,In_793);
nor U1233 (N_1233,In_1258,In_568);
nand U1234 (N_1234,In_52,In_1011);
nand U1235 (N_1235,In_1434,In_1000);
or U1236 (N_1236,In_643,In_300);
nor U1237 (N_1237,In_1287,In_190);
nor U1238 (N_1238,In_700,In_381);
or U1239 (N_1239,In_512,In_573);
or U1240 (N_1240,In_231,In_338);
nand U1241 (N_1241,In_130,In_243);
and U1242 (N_1242,In_486,In_204);
and U1243 (N_1243,In_1253,In_732);
and U1244 (N_1244,In_1152,In_857);
nor U1245 (N_1245,In_314,In_1449);
or U1246 (N_1246,In_371,In_953);
and U1247 (N_1247,In_695,In_1277);
nand U1248 (N_1248,In_501,In_895);
nor U1249 (N_1249,In_434,In_1015);
nand U1250 (N_1250,In_1409,In_724);
or U1251 (N_1251,In_1038,In_855);
and U1252 (N_1252,In_1476,In_207);
or U1253 (N_1253,In_1187,In_1341);
nand U1254 (N_1254,In_652,In_839);
nand U1255 (N_1255,In_140,In_1491);
or U1256 (N_1256,In_1220,In_162);
nand U1257 (N_1257,In_979,In_1096);
nand U1258 (N_1258,In_1077,In_341);
nand U1259 (N_1259,In_1380,In_1030);
nor U1260 (N_1260,In_649,In_203);
nand U1261 (N_1261,In_615,In_736);
nand U1262 (N_1262,In_1285,In_513);
and U1263 (N_1263,In_1137,In_891);
nand U1264 (N_1264,In_1234,In_983);
nor U1265 (N_1265,In_579,In_864);
nand U1266 (N_1266,In_1438,In_465);
or U1267 (N_1267,In_1181,In_1212);
nand U1268 (N_1268,In_675,In_670);
nor U1269 (N_1269,In_1325,In_31);
or U1270 (N_1270,In_1136,In_984);
and U1271 (N_1271,In_24,In_1205);
and U1272 (N_1272,In_575,In_365);
nor U1273 (N_1273,In_1125,In_1182);
and U1274 (N_1274,In_202,In_119);
nand U1275 (N_1275,In_1085,In_1043);
and U1276 (N_1276,In_1148,In_1203);
nor U1277 (N_1277,In_1475,In_476);
and U1278 (N_1278,In_232,In_822);
nand U1279 (N_1279,In_333,In_1457);
xor U1280 (N_1280,In_505,In_243);
and U1281 (N_1281,In_270,In_793);
or U1282 (N_1282,In_1023,In_140);
or U1283 (N_1283,In_67,In_1045);
or U1284 (N_1284,In_1075,In_1104);
nor U1285 (N_1285,In_1488,In_392);
or U1286 (N_1286,In_562,In_1443);
nand U1287 (N_1287,In_983,In_462);
and U1288 (N_1288,In_519,In_1343);
nor U1289 (N_1289,In_706,In_1157);
or U1290 (N_1290,In_906,In_97);
nor U1291 (N_1291,In_1134,In_275);
and U1292 (N_1292,In_14,In_1013);
or U1293 (N_1293,In_587,In_350);
or U1294 (N_1294,In_465,In_1243);
or U1295 (N_1295,In_1332,In_1033);
nor U1296 (N_1296,In_582,In_1438);
or U1297 (N_1297,In_1237,In_1229);
and U1298 (N_1298,In_304,In_909);
and U1299 (N_1299,In_222,In_941);
or U1300 (N_1300,In_1444,In_1119);
nand U1301 (N_1301,In_240,In_1473);
nor U1302 (N_1302,In_1114,In_696);
nand U1303 (N_1303,In_837,In_221);
or U1304 (N_1304,In_1177,In_272);
nand U1305 (N_1305,In_603,In_1450);
nand U1306 (N_1306,In_475,In_548);
xnor U1307 (N_1307,In_1043,In_14);
nand U1308 (N_1308,In_238,In_1394);
nor U1309 (N_1309,In_298,In_785);
nand U1310 (N_1310,In_1195,In_1086);
nor U1311 (N_1311,In_807,In_1454);
or U1312 (N_1312,In_209,In_697);
nor U1313 (N_1313,In_220,In_336);
nand U1314 (N_1314,In_1380,In_399);
nor U1315 (N_1315,In_113,In_163);
nor U1316 (N_1316,In_169,In_782);
or U1317 (N_1317,In_348,In_582);
nor U1318 (N_1318,In_605,In_465);
nor U1319 (N_1319,In_1079,In_524);
or U1320 (N_1320,In_832,In_1475);
and U1321 (N_1321,In_1312,In_802);
and U1322 (N_1322,In_814,In_788);
or U1323 (N_1323,In_563,In_21);
nand U1324 (N_1324,In_419,In_1228);
nand U1325 (N_1325,In_1270,In_264);
nand U1326 (N_1326,In_47,In_824);
and U1327 (N_1327,In_670,In_1335);
nand U1328 (N_1328,In_1427,In_478);
nand U1329 (N_1329,In_1182,In_163);
nand U1330 (N_1330,In_55,In_816);
nand U1331 (N_1331,In_113,In_623);
nor U1332 (N_1332,In_719,In_872);
nor U1333 (N_1333,In_244,In_1009);
and U1334 (N_1334,In_1346,In_33);
nand U1335 (N_1335,In_18,In_327);
or U1336 (N_1336,In_538,In_1238);
nor U1337 (N_1337,In_1460,In_299);
and U1338 (N_1338,In_491,In_387);
and U1339 (N_1339,In_218,In_564);
or U1340 (N_1340,In_638,In_1390);
or U1341 (N_1341,In_423,In_133);
or U1342 (N_1342,In_495,In_772);
and U1343 (N_1343,In_749,In_558);
nand U1344 (N_1344,In_717,In_857);
nor U1345 (N_1345,In_52,In_314);
and U1346 (N_1346,In_161,In_1242);
and U1347 (N_1347,In_479,In_816);
and U1348 (N_1348,In_1204,In_742);
or U1349 (N_1349,In_537,In_639);
and U1350 (N_1350,In_215,In_356);
and U1351 (N_1351,In_1466,In_534);
nor U1352 (N_1352,In_564,In_529);
and U1353 (N_1353,In_369,In_267);
or U1354 (N_1354,In_110,In_1060);
or U1355 (N_1355,In_163,In_1227);
or U1356 (N_1356,In_1290,In_1431);
or U1357 (N_1357,In_1217,In_409);
and U1358 (N_1358,In_1363,In_943);
nand U1359 (N_1359,In_133,In_305);
nand U1360 (N_1360,In_1396,In_875);
or U1361 (N_1361,In_1073,In_511);
nand U1362 (N_1362,In_1169,In_1376);
nand U1363 (N_1363,In_232,In_372);
and U1364 (N_1364,In_827,In_703);
or U1365 (N_1365,In_1271,In_623);
nor U1366 (N_1366,In_928,In_1365);
and U1367 (N_1367,In_1397,In_565);
and U1368 (N_1368,In_609,In_284);
and U1369 (N_1369,In_538,In_867);
and U1370 (N_1370,In_949,In_584);
nor U1371 (N_1371,In_82,In_1001);
and U1372 (N_1372,In_1,In_514);
or U1373 (N_1373,In_39,In_459);
and U1374 (N_1374,In_1202,In_595);
or U1375 (N_1375,In_835,In_157);
or U1376 (N_1376,In_1378,In_426);
nor U1377 (N_1377,In_1358,In_857);
nand U1378 (N_1378,In_514,In_200);
nand U1379 (N_1379,In_118,In_1295);
and U1380 (N_1380,In_1206,In_269);
and U1381 (N_1381,In_29,In_798);
and U1382 (N_1382,In_965,In_861);
or U1383 (N_1383,In_79,In_1197);
or U1384 (N_1384,In_489,In_326);
or U1385 (N_1385,In_1334,In_120);
or U1386 (N_1386,In_352,In_456);
nor U1387 (N_1387,In_69,In_475);
nand U1388 (N_1388,In_75,In_785);
and U1389 (N_1389,In_1159,In_793);
nand U1390 (N_1390,In_1353,In_580);
nor U1391 (N_1391,In_152,In_183);
or U1392 (N_1392,In_379,In_456);
and U1393 (N_1393,In_984,In_1483);
and U1394 (N_1394,In_823,In_341);
or U1395 (N_1395,In_1096,In_1039);
and U1396 (N_1396,In_47,In_217);
and U1397 (N_1397,In_1135,In_1272);
nor U1398 (N_1398,In_1095,In_1194);
and U1399 (N_1399,In_105,In_77);
or U1400 (N_1400,In_742,In_738);
and U1401 (N_1401,In_229,In_322);
nor U1402 (N_1402,In_499,In_1458);
or U1403 (N_1403,In_406,In_1014);
nor U1404 (N_1404,In_664,In_1417);
nand U1405 (N_1405,In_959,In_818);
nor U1406 (N_1406,In_1055,In_1121);
and U1407 (N_1407,In_301,In_1245);
and U1408 (N_1408,In_715,In_1160);
nor U1409 (N_1409,In_1214,In_7);
nor U1410 (N_1410,In_1210,In_1411);
nor U1411 (N_1411,In_1414,In_817);
nand U1412 (N_1412,In_188,In_196);
or U1413 (N_1413,In_745,In_495);
nor U1414 (N_1414,In_341,In_952);
nand U1415 (N_1415,In_241,In_1245);
nor U1416 (N_1416,In_485,In_452);
and U1417 (N_1417,In_1477,In_788);
nor U1418 (N_1418,In_485,In_803);
or U1419 (N_1419,In_678,In_1307);
or U1420 (N_1420,In_1,In_1455);
nand U1421 (N_1421,In_416,In_845);
or U1422 (N_1422,In_627,In_949);
and U1423 (N_1423,In_803,In_1341);
nor U1424 (N_1424,In_1170,In_409);
nand U1425 (N_1425,In_95,In_755);
nand U1426 (N_1426,In_558,In_856);
nand U1427 (N_1427,In_581,In_251);
nand U1428 (N_1428,In_260,In_850);
nor U1429 (N_1429,In_462,In_246);
nand U1430 (N_1430,In_542,In_785);
nor U1431 (N_1431,In_902,In_935);
and U1432 (N_1432,In_594,In_1391);
or U1433 (N_1433,In_322,In_738);
nor U1434 (N_1434,In_1492,In_970);
and U1435 (N_1435,In_741,In_66);
nand U1436 (N_1436,In_810,In_305);
nand U1437 (N_1437,In_1261,In_695);
nand U1438 (N_1438,In_1032,In_789);
nand U1439 (N_1439,In_1295,In_751);
xor U1440 (N_1440,In_928,In_1366);
or U1441 (N_1441,In_1422,In_418);
and U1442 (N_1442,In_154,In_1050);
nand U1443 (N_1443,In_1040,In_798);
and U1444 (N_1444,In_373,In_1004);
nor U1445 (N_1445,In_359,In_9);
nand U1446 (N_1446,In_1237,In_1186);
nand U1447 (N_1447,In_97,In_353);
or U1448 (N_1448,In_868,In_1272);
nor U1449 (N_1449,In_249,In_1456);
and U1450 (N_1450,In_189,In_1082);
nand U1451 (N_1451,In_646,In_1340);
nand U1452 (N_1452,In_1358,In_796);
and U1453 (N_1453,In_249,In_210);
nand U1454 (N_1454,In_1346,In_490);
nor U1455 (N_1455,In_876,In_100);
nand U1456 (N_1456,In_540,In_1263);
nor U1457 (N_1457,In_754,In_1398);
nand U1458 (N_1458,In_1169,In_1232);
and U1459 (N_1459,In_113,In_1069);
or U1460 (N_1460,In_80,In_877);
and U1461 (N_1461,In_127,In_8);
nor U1462 (N_1462,In_40,In_324);
and U1463 (N_1463,In_867,In_943);
or U1464 (N_1464,In_778,In_916);
nor U1465 (N_1465,In_205,In_677);
nand U1466 (N_1466,In_1265,In_815);
nor U1467 (N_1467,In_284,In_1456);
nand U1468 (N_1468,In_528,In_356);
and U1469 (N_1469,In_1151,In_1022);
or U1470 (N_1470,In_1208,In_1131);
and U1471 (N_1471,In_1204,In_1081);
nor U1472 (N_1472,In_949,In_702);
and U1473 (N_1473,In_115,In_206);
nand U1474 (N_1474,In_1128,In_463);
nand U1475 (N_1475,In_866,In_1054);
and U1476 (N_1476,In_554,In_930);
nand U1477 (N_1477,In_62,In_1310);
nand U1478 (N_1478,In_1393,In_39);
nor U1479 (N_1479,In_73,In_1253);
or U1480 (N_1480,In_904,In_1216);
and U1481 (N_1481,In_1211,In_59);
nand U1482 (N_1482,In_1012,In_128);
nor U1483 (N_1483,In_617,In_761);
and U1484 (N_1484,In_282,In_66);
and U1485 (N_1485,In_590,In_661);
and U1486 (N_1486,In_649,In_1228);
and U1487 (N_1487,In_423,In_387);
nand U1488 (N_1488,In_278,In_1393);
nand U1489 (N_1489,In_908,In_445);
nor U1490 (N_1490,In_246,In_696);
nor U1491 (N_1491,In_1325,In_125);
nor U1492 (N_1492,In_1416,In_822);
nand U1493 (N_1493,In_794,In_640);
and U1494 (N_1494,In_625,In_580);
nor U1495 (N_1495,In_1072,In_205);
and U1496 (N_1496,In_899,In_671);
nand U1497 (N_1497,In_905,In_239);
or U1498 (N_1498,In_1433,In_874);
nand U1499 (N_1499,In_458,In_912);
or U1500 (N_1500,In_1015,In_643);
nand U1501 (N_1501,In_1257,In_217);
and U1502 (N_1502,In_509,In_901);
nand U1503 (N_1503,In_1015,In_1331);
or U1504 (N_1504,In_1374,In_37);
nand U1505 (N_1505,In_1000,In_22);
nor U1506 (N_1506,In_684,In_771);
nor U1507 (N_1507,In_1407,In_426);
nand U1508 (N_1508,In_252,In_774);
nand U1509 (N_1509,In_698,In_583);
nor U1510 (N_1510,In_1169,In_633);
nand U1511 (N_1511,In_1375,In_994);
or U1512 (N_1512,In_1130,In_868);
nand U1513 (N_1513,In_858,In_394);
or U1514 (N_1514,In_839,In_184);
nand U1515 (N_1515,In_1088,In_670);
or U1516 (N_1516,In_640,In_689);
and U1517 (N_1517,In_246,In_190);
nor U1518 (N_1518,In_1141,In_743);
and U1519 (N_1519,In_1382,In_945);
and U1520 (N_1520,In_944,In_866);
or U1521 (N_1521,In_1434,In_54);
nor U1522 (N_1522,In_749,In_813);
and U1523 (N_1523,In_733,In_661);
and U1524 (N_1524,In_1324,In_891);
nand U1525 (N_1525,In_1347,In_397);
and U1526 (N_1526,In_603,In_1195);
nor U1527 (N_1527,In_714,In_1345);
or U1528 (N_1528,In_404,In_44);
nand U1529 (N_1529,In_1237,In_1145);
nand U1530 (N_1530,In_1123,In_911);
and U1531 (N_1531,In_178,In_856);
and U1532 (N_1532,In_1388,In_387);
nor U1533 (N_1533,In_1290,In_1259);
nor U1534 (N_1534,In_1198,In_781);
and U1535 (N_1535,In_1467,In_916);
nor U1536 (N_1536,In_939,In_1103);
and U1537 (N_1537,In_209,In_221);
and U1538 (N_1538,In_980,In_743);
and U1539 (N_1539,In_1111,In_1332);
and U1540 (N_1540,In_1498,In_1364);
nand U1541 (N_1541,In_1358,In_409);
nor U1542 (N_1542,In_1162,In_1144);
or U1543 (N_1543,In_1039,In_1183);
or U1544 (N_1544,In_661,In_770);
nand U1545 (N_1545,In_452,In_898);
nor U1546 (N_1546,In_1073,In_1483);
and U1547 (N_1547,In_651,In_252);
nand U1548 (N_1548,In_74,In_1336);
or U1549 (N_1549,In_400,In_1215);
and U1550 (N_1550,In_1333,In_673);
nand U1551 (N_1551,In_480,In_1281);
nor U1552 (N_1552,In_1391,In_609);
and U1553 (N_1553,In_34,In_704);
nand U1554 (N_1554,In_576,In_969);
or U1555 (N_1555,In_476,In_1432);
or U1556 (N_1556,In_997,In_97);
nand U1557 (N_1557,In_957,In_387);
or U1558 (N_1558,In_185,In_1466);
and U1559 (N_1559,In_1439,In_619);
nand U1560 (N_1560,In_8,In_311);
or U1561 (N_1561,In_393,In_62);
and U1562 (N_1562,In_902,In_1333);
nor U1563 (N_1563,In_1079,In_1046);
nor U1564 (N_1564,In_389,In_299);
nor U1565 (N_1565,In_1044,In_657);
and U1566 (N_1566,In_977,In_329);
nand U1567 (N_1567,In_840,In_741);
and U1568 (N_1568,In_538,In_486);
nor U1569 (N_1569,In_736,In_715);
nor U1570 (N_1570,In_909,In_1026);
nor U1571 (N_1571,In_711,In_971);
nor U1572 (N_1572,In_1383,In_391);
and U1573 (N_1573,In_843,In_600);
xnor U1574 (N_1574,In_1434,In_644);
and U1575 (N_1575,In_736,In_604);
nand U1576 (N_1576,In_1209,In_1082);
nor U1577 (N_1577,In_124,In_259);
nand U1578 (N_1578,In_1021,In_776);
or U1579 (N_1579,In_942,In_967);
and U1580 (N_1580,In_208,In_1226);
or U1581 (N_1581,In_514,In_826);
nand U1582 (N_1582,In_98,In_1105);
nor U1583 (N_1583,In_1126,In_123);
nand U1584 (N_1584,In_535,In_787);
nor U1585 (N_1585,In_1383,In_1089);
nor U1586 (N_1586,In_700,In_37);
nor U1587 (N_1587,In_1319,In_772);
nand U1588 (N_1588,In_282,In_1386);
and U1589 (N_1589,In_247,In_1436);
nor U1590 (N_1590,In_971,In_312);
nand U1591 (N_1591,In_1144,In_1209);
nand U1592 (N_1592,In_534,In_424);
nor U1593 (N_1593,In_304,In_67);
nand U1594 (N_1594,In_33,In_1245);
nand U1595 (N_1595,In_969,In_1489);
nand U1596 (N_1596,In_64,In_411);
nor U1597 (N_1597,In_1367,In_278);
or U1598 (N_1598,In_1287,In_138);
nand U1599 (N_1599,In_564,In_611);
nor U1600 (N_1600,In_166,In_1024);
nand U1601 (N_1601,In_76,In_298);
xnor U1602 (N_1602,In_1199,In_919);
nand U1603 (N_1603,In_500,In_544);
or U1604 (N_1604,In_635,In_146);
and U1605 (N_1605,In_1124,In_1295);
nand U1606 (N_1606,In_877,In_692);
or U1607 (N_1607,In_855,In_1027);
or U1608 (N_1608,In_1282,In_442);
nand U1609 (N_1609,In_1077,In_1471);
nand U1610 (N_1610,In_138,In_297);
and U1611 (N_1611,In_475,In_729);
nand U1612 (N_1612,In_960,In_1159);
and U1613 (N_1613,In_288,In_1255);
and U1614 (N_1614,In_844,In_71);
nor U1615 (N_1615,In_57,In_711);
nor U1616 (N_1616,In_1464,In_734);
nand U1617 (N_1617,In_1375,In_93);
or U1618 (N_1618,In_593,In_1355);
nor U1619 (N_1619,In_803,In_732);
or U1620 (N_1620,In_374,In_1160);
and U1621 (N_1621,In_695,In_1310);
or U1622 (N_1622,In_1253,In_926);
or U1623 (N_1623,In_1391,In_1226);
nand U1624 (N_1624,In_1120,In_1216);
nor U1625 (N_1625,In_687,In_163);
or U1626 (N_1626,In_161,In_995);
and U1627 (N_1627,In_737,In_215);
nand U1628 (N_1628,In_862,In_1252);
or U1629 (N_1629,In_852,In_1487);
nor U1630 (N_1630,In_1463,In_1488);
nand U1631 (N_1631,In_1420,In_1431);
nand U1632 (N_1632,In_983,In_1163);
nor U1633 (N_1633,In_315,In_6);
nand U1634 (N_1634,In_11,In_1036);
nand U1635 (N_1635,In_121,In_12);
or U1636 (N_1636,In_500,In_743);
or U1637 (N_1637,In_1487,In_277);
or U1638 (N_1638,In_1037,In_887);
nand U1639 (N_1639,In_1130,In_1496);
or U1640 (N_1640,In_800,In_156);
nor U1641 (N_1641,In_610,In_807);
nor U1642 (N_1642,In_1360,In_872);
nor U1643 (N_1643,In_1419,In_914);
and U1644 (N_1644,In_753,In_494);
xnor U1645 (N_1645,In_440,In_1400);
or U1646 (N_1646,In_1072,In_1036);
and U1647 (N_1647,In_281,In_935);
and U1648 (N_1648,In_1268,In_31);
and U1649 (N_1649,In_1286,In_23);
and U1650 (N_1650,In_1495,In_1228);
nand U1651 (N_1651,In_62,In_1132);
nor U1652 (N_1652,In_643,In_532);
nand U1653 (N_1653,In_1454,In_869);
or U1654 (N_1654,In_968,In_786);
or U1655 (N_1655,In_43,In_889);
and U1656 (N_1656,In_630,In_581);
nor U1657 (N_1657,In_1156,In_727);
or U1658 (N_1658,In_600,In_573);
nand U1659 (N_1659,In_1058,In_1208);
nand U1660 (N_1660,In_449,In_642);
and U1661 (N_1661,In_324,In_79);
nor U1662 (N_1662,In_1103,In_1182);
and U1663 (N_1663,In_552,In_1278);
nor U1664 (N_1664,In_659,In_334);
or U1665 (N_1665,In_11,In_53);
nor U1666 (N_1666,In_926,In_1200);
xnor U1667 (N_1667,In_568,In_746);
or U1668 (N_1668,In_1247,In_595);
nor U1669 (N_1669,In_1155,In_290);
or U1670 (N_1670,In_903,In_524);
nand U1671 (N_1671,In_860,In_93);
nor U1672 (N_1672,In_1402,In_276);
nor U1673 (N_1673,In_1196,In_549);
nand U1674 (N_1674,In_184,In_446);
nand U1675 (N_1675,In_480,In_441);
or U1676 (N_1676,In_220,In_75);
or U1677 (N_1677,In_1077,In_573);
or U1678 (N_1678,In_1159,In_1493);
and U1679 (N_1679,In_1388,In_209);
nor U1680 (N_1680,In_1214,In_579);
nor U1681 (N_1681,In_1346,In_403);
nor U1682 (N_1682,In_194,In_1017);
nand U1683 (N_1683,In_911,In_1363);
nand U1684 (N_1684,In_127,In_943);
xnor U1685 (N_1685,In_220,In_1254);
or U1686 (N_1686,In_392,In_633);
or U1687 (N_1687,In_1081,In_958);
or U1688 (N_1688,In_754,In_1409);
or U1689 (N_1689,In_1412,In_169);
or U1690 (N_1690,In_627,In_1205);
nand U1691 (N_1691,In_1293,In_1043);
nor U1692 (N_1692,In_186,In_204);
and U1693 (N_1693,In_493,In_135);
nand U1694 (N_1694,In_834,In_605);
nor U1695 (N_1695,In_1160,In_480);
and U1696 (N_1696,In_453,In_315);
nand U1697 (N_1697,In_814,In_924);
nor U1698 (N_1698,In_328,In_332);
and U1699 (N_1699,In_507,In_315);
nor U1700 (N_1700,In_332,In_62);
nor U1701 (N_1701,In_110,In_999);
nand U1702 (N_1702,In_630,In_895);
nand U1703 (N_1703,In_315,In_178);
nand U1704 (N_1704,In_217,In_277);
and U1705 (N_1705,In_122,In_639);
nor U1706 (N_1706,In_676,In_371);
nand U1707 (N_1707,In_148,In_401);
nor U1708 (N_1708,In_161,In_275);
and U1709 (N_1709,In_747,In_552);
nand U1710 (N_1710,In_746,In_396);
nor U1711 (N_1711,In_1264,In_653);
or U1712 (N_1712,In_278,In_1072);
or U1713 (N_1713,In_1257,In_514);
nor U1714 (N_1714,In_120,In_783);
nor U1715 (N_1715,In_569,In_920);
nand U1716 (N_1716,In_884,In_777);
nor U1717 (N_1717,In_148,In_1135);
and U1718 (N_1718,In_1127,In_480);
nor U1719 (N_1719,In_1347,In_186);
nand U1720 (N_1720,In_688,In_714);
nand U1721 (N_1721,In_44,In_12);
nor U1722 (N_1722,In_196,In_98);
nor U1723 (N_1723,In_1187,In_1034);
xor U1724 (N_1724,In_919,In_542);
and U1725 (N_1725,In_602,In_1372);
and U1726 (N_1726,In_997,In_249);
and U1727 (N_1727,In_1455,In_713);
or U1728 (N_1728,In_689,In_1362);
nor U1729 (N_1729,In_1084,In_237);
nand U1730 (N_1730,In_301,In_165);
nor U1731 (N_1731,In_1018,In_1064);
or U1732 (N_1732,In_1163,In_1398);
nor U1733 (N_1733,In_745,In_1470);
nor U1734 (N_1734,In_235,In_67);
or U1735 (N_1735,In_965,In_1372);
or U1736 (N_1736,In_1056,In_77);
or U1737 (N_1737,In_1413,In_1497);
nor U1738 (N_1738,In_1392,In_524);
and U1739 (N_1739,In_1075,In_445);
and U1740 (N_1740,In_679,In_1471);
nor U1741 (N_1741,In_700,In_335);
or U1742 (N_1742,In_1103,In_1227);
nor U1743 (N_1743,In_250,In_1136);
and U1744 (N_1744,In_383,In_66);
or U1745 (N_1745,In_1381,In_550);
and U1746 (N_1746,In_1326,In_188);
nor U1747 (N_1747,In_752,In_172);
nand U1748 (N_1748,In_116,In_883);
or U1749 (N_1749,In_1108,In_1429);
or U1750 (N_1750,In_784,In_409);
or U1751 (N_1751,In_1026,In_351);
nor U1752 (N_1752,In_18,In_1479);
nor U1753 (N_1753,In_1055,In_111);
or U1754 (N_1754,In_31,In_1443);
or U1755 (N_1755,In_1118,In_1420);
nor U1756 (N_1756,In_251,In_933);
or U1757 (N_1757,In_1497,In_1315);
nor U1758 (N_1758,In_58,In_950);
nand U1759 (N_1759,In_934,In_553);
and U1760 (N_1760,In_1475,In_569);
and U1761 (N_1761,In_331,In_1354);
nand U1762 (N_1762,In_310,In_215);
nand U1763 (N_1763,In_469,In_1094);
nor U1764 (N_1764,In_82,In_858);
nand U1765 (N_1765,In_790,In_511);
nand U1766 (N_1766,In_354,In_1065);
nand U1767 (N_1767,In_707,In_1380);
or U1768 (N_1768,In_654,In_235);
or U1769 (N_1769,In_1369,In_1199);
nor U1770 (N_1770,In_843,In_1429);
or U1771 (N_1771,In_551,In_740);
and U1772 (N_1772,In_273,In_432);
and U1773 (N_1773,In_22,In_723);
nor U1774 (N_1774,In_67,In_123);
and U1775 (N_1775,In_562,In_873);
and U1776 (N_1776,In_573,In_787);
nor U1777 (N_1777,In_798,In_26);
and U1778 (N_1778,In_466,In_980);
or U1779 (N_1779,In_1493,In_1439);
nor U1780 (N_1780,In_627,In_732);
and U1781 (N_1781,In_1406,In_483);
nor U1782 (N_1782,In_115,In_956);
nor U1783 (N_1783,In_933,In_245);
nand U1784 (N_1784,In_1257,In_1399);
nor U1785 (N_1785,In_476,In_710);
or U1786 (N_1786,In_371,In_1190);
or U1787 (N_1787,In_1286,In_117);
nor U1788 (N_1788,In_38,In_177);
nor U1789 (N_1789,In_796,In_1136);
nand U1790 (N_1790,In_673,In_60);
and U1791 (N_1791,In_748,In_175);
xnor U1792 (N_1792,In_528,In_1378);
nand U1793 (N_1793,In_1202,In_458);
or U1794 (N_1794,In_997,In_402);
or U1795 (N_1795,In_21,In_268);
nor U1796 (N_1796,In_1172,In_667);
nand U1797 (N_1797,In_1437,In_1432);
and U1798 (N_1798,In_1390,In_1053);
nand U1799 (N_1799,In_875,In_1262);
and U1800 (N_1800,In_537,In_1333);
nor U1801 (N_1801,In_505,In_751);
nor U1802 (N_1802,In_1212,In_657);
or U1803 (N_1803,In_295,In_13);
nor U1804 (N_1804,In_907,In_1008);
nand U1805 (N_1805,In_769,In_396);
and U1806 (N_1806,In_684,In_811);
nor U1807 (N_1807,In_166,In_46);
nand U1808 (N_1808,In_373,In_1059);
nand U1809 (N_1809,In_482,In_1132);
and U1810 (N_1810,In_929,In_856);
nand U1811 (N_1811,In_319,In_391);
or U1812 (N_1812,In_104,In_1415);
or U1813 (N_1813,In_728,In_1353);
nor U1814 (N_1814,In_94,In_1071);
nor U1815 (N_1815,In_979,In_1181);
and U1816 (N_1816,In_92,In_1002);
nor U1817 (N_1817,In_808,In_410);
nor U1818 (N_1818,In_78,In_1333);
or U1819 (N_1819,In_848,In_1055);
nor U1820 (N_1820,In_1175,In_830);
nand U1821 (N_1821,In_685,In_734);
nand U1822 (N_1822,In_408,In_1175);
nor U1823 (N_1823,In_968,In_35);
nand U1824 (N_1824,In_301,In_1124);
nor U1825 (N_1825,In_295,In_1347);
nor U1826 (N_1826,In_83,In_1402);
or U1827 (N_1827,In_1158,In_1429);
or U1828 (N_1828,In_825,In_1264);
nor U1829 (N_1829,In_812,In_299);
or U1830 (N_1830,In_149,In_16);
or U1831 (N_1831,In_1027,In_716);
nand U1832 (N_1832,In_321,In_827);
and U1833 (N_1833,In_955,In_1028);
nand U1834 (N_1834,In_831,In_373);
nor U1835 (N_1835,In_670,In_632);
nand U1836 (N_1836,In_199,In_1410);
nor U1837 (N_1837,In_261,In_700);
and U1838 (N_1838,In_335,In_946);
and U1839 (N_1839,In_512,In_741);
or U1840 (N_1840,In_793,In_604);
or U1841 (N_1841,In_123,In_1086);
or U1842 (N_1842,In_1275,In_1260);
nand U1843 (N_1843,In_176,In_279);
nor U1844 (N_1844,In_721,In_716);
nor U1845 (N_1845,In_1153,In_940);
nor U1846 (N_1846,In_1210,In_1218);
or U1847 (N_1847,In_1151,In_1227);
or U1848 (N_1848,In_1492,In_849);
and U1849 (N_1849,In_1101,In_781);
and U1850 (N_1850,In_25,In_1310);
nor U1851 (N_1851,In_58,In_212);
and U1852 (N_1852,In_1314,In_82);
or U1853 (N_1853,In_399,In_553);
nand U1854 (N_1854,In_199,In_641);
nand U1855 (N_1855,In_603,In_870);
nand U1856 (N_1856,In_191,In_1244);
and U1857 (N_1857,In_384,In_391);
or U1858 (N_1858,In_52,In_1158);
nor U1859 (N_1859,In_859,In_1486);
nand U1860 (N_1860,In_544,In_1212);
nor U1861 (N_1861,In_1364,In_727);
nor U1862 (N_1862,In_72,In_239);
or U1863 (N_1863,In_848,In_837);
nor U1864 (N_1864,In_1019,In_1441);
nand U1865 (N_1865,In_1465,In_805);
nor U1866 (N_1866,In_118,In_817);
nor U1867 (N_1867,In_987,In_9);
or U1868 (N_1868,In_680,In_15);
or U1869 (N_1869,In_1090,In_1162);
nor U1870 (N_1870,In_310,In_423);
or U1871 (N_1871,In_648,In_1261);
and U1872 (N_1872,In_1427,In_1152);
or U1873 (N_1873,In_620,In_843);
or U1874 (N_1874,In_141,In_1478);
and U1875 (N_1875,In_1129,In_1488);
nand U1876 (N_1876,In_669,In_261);
and U1877 (N_1877,In_1041,In_1274);
or U1878 (N_1878,In_186,In_106);
or U1879 (N_1879,In_819,In_106);
nand U1880 (N_1880,In_1352,In_1446);
or U1881 (N_1881,In_1262,In_1210);
and U1882 (N_1882,In_38,In_1343);
nor U1883 (N_1883,In_814,In_761);
and U1884 (N_1884,In_784,In_870);
and U1885 (N_1885,In_1390,In_1153);
or U1886 (N_1886,In_179,In_695);
or U1887 (N_1887,In_250,In_88);
or U1888 (N_1888,In_765,In_1322);
nand U1889 (N_1889,In_289,In_1075);
nor U1890 (N_1890,In_900,In_1257);
and U1891 (N_1891,In_588,In_149);
and U1892 (N_1892,In_979,In_1375);
nand U1893 (N_1893,In_1424,In_1250);
nor U1894 (N_1894,In_1415,In_792);
and U1895 (N_1895,In_1335,In_477);
nor U1896 (N_1896,In_1350,In_258);
nand U1897 (N_1897,In_101,In_634);
and U1898 (N_1898,In_448,In_1083);
nand U1899 (N_1899,In_26,In_590);
nor U1900 (N_1900,In_887,In_1381);
nand U1901 (N_1901,In_1357,In_618);
nand U1902 (N_1902,In_121,In_1095);
nand U1903 (N_1903,In_724,In_792);
nor U1904 (N_1904,In_410,In_338);
nand U1905 (N_1905,In_646,In_1141);
and U1906 (N_1906,In_171,In_691);
and U1907 (N_1907,In_131,In_127);
and U1908 (N_1908,In_469,In_495);
nand U1909 (N_1909,In_984,In_669);
nor U1910 (N_1910,In_222,In_108);
and U1911 (N_1911,In_1144,In_246);
nand U1912 (N_1912,In_1487,In_667);
nand U1913 (N_1913,In_505,In_941);
nand U1914 (N_1914,In_45,In_269);
and U1915 (N_1915,In_869,In_140);
nor U1916 (N_1916,In_979,In_304);
and U1917 (N_1917,In_1032,In_981);
or U1918 (N_1918,In_285,In_414);
nor U1919 (N_1919,In_558,In_1068);
and U1920 (N_1920,In_948,In_364);
or U1921 (N_1921,In_39,In_1256);
and U1922 (N_1922,In_964,In_1308);
nand U1923 (N_1923,In_86,In_38);
nor U1924 (N_1924,In_1185,In_852);
nor U1925 (N_1925,In_606,In_721);
nand U1926 (N_1926,In_1116,In_307);
nand U1927 (N_1927,In_439,In_19);
nor U1928 (N_1928,In_1325,In_1168);
nand U1929 (N_1929,In_1142,In_739);
or U1930 (N_1930,In_159,In_95);
or U1931 (N_1931,In_166,In_367);
nor U1932 (N_1932,In_1453,In_866);
nor U1933 (N_1933,In_435,In_966);
or U1934 (N_1934,In_843,In_1490);
nand U1935 (N_1935,In_330,In_779);
nor U1936 (N_1936,In_88,In_447);
nand U1937 (N_1937,In_81,In_1045);
nand U1938 (N_1938,In_102,In_433);
and U1939 (N_1939,In_865,In_1066);
and U1940 (N_1940,In_918,In_1204);
and U1941 (N_1941,In_1293,In_370);
and U1942 (N_1942,In_433,In_18);
nand U1943 (N_1943,In_1187,In_843);
nor U1944 (N_1944,In_429,In_296);
nor U1945 (N_1945,In_818,In_528);
xnor U1946 (N_1946,In_217,In_896);
or U1947 (N_1947,In_245,In_1183);
or U1948 (N_1948,In_579,In_716);
or U1949 (N_1949,In_412,In_115);
or U1950 (N_1950,In_942,In_74);
or U1951 (N_1951,In_1211,In_35);
nor U1952 (N_1952,In_1268,In_22);
or U1953 (N_1953,In_791,In_1224);
and U1954 (N_1954,In_251,In_556);
and U1955 (N_1955,In_844,In_1444);
nor U1956 (N_1956,In_329,In_1385);
nor U1957 (N_1957,In_901,In_465);
nor U1958 (N_1958,In_696,In_582);
nand U1959 (N_1959,In_220,In_912);
and U1960 (N_1960,In_1336,In_22);
nor U1961 (N_1961,In_1409,In_758);
nor U1962 (N_1962,In_119,In_848);
nand U1963 (N_1963,In_401,In_952);
nor U1964 (N_1964,In_678,In_967);
and U1965 (N_1965,In_5,In_482);
nor U1966 (N_1966,In_1181,In_876);
or U1967 (N_1967,In_1412,In_1003);
or U1968 (N_1968,In_1159,In_1360);
or U1969 (N_1969,In_161,In_392);
nand U1970 (N_1970,In_960,In_269);
nand U1971 (N_1971,In_1234,In_1034);
nor U1972 (N_1972,In_1059,In_998);
or U1973 (N_1973,In_677,In_380);
nand U1974 (N_1974,In_496,In_470);
or U1975 (N_1975,In_136,In_1224);
and U1976 (N_1976,In_1330,In_674);
and U1977 (N_1977,In_1450,In_35);
nor U1978 (N_1978,In_626,In_85);
nor U1979 (N_1979,In_142,In_1284);
or U1980 (N_1980,In_608,In_243);
and U1981 (N_1981,In_344,In_618);
nand U1982 (N_1982,In_852,In_1311);
or U1983 (N_1983,In_1104,In_7);
and U1984 (N_1984,In_105,In_686);
nand U1985 (N_1985,In_1158,In_457);
nor U1986 (N_1986,In_1035,In_152);
nor U1987 (N_1987,In_1162,In_392);
nand U1988 (N_1988,In_20,In_356);
and U1989 (N_1989,In_60,In_823);
nor U1990 (N_1990,In_1374,In_454);
nor U1991 (N_1991,In_883,In_560);
or U1992 (N_1992,In_1368,In_585);
nand U1993 (N_1993,In_1386,In_929);
or U1994 (N_1994,In_1362,In_987);
or U1995 (N_1995,In_793,In_1096);
and U1996 (N_1996,In_93,In_1453);
or U1997 (N_1997,In_677,In_1151);
and U1998 (N_1998,In_824,In_847);
and U1999 (N_1999,In_666,In_1126);
or U2000 (N_2000,In_646,In_1403);
nand U2001 (N_2001,In_1000,In_163);
nand U2002 (N_2002,In_1349,In_509);
nor U2003 (N_2003,In_318,In_812);
nor U2004 (N_2004,In_795,In_259);
and U2005 (N_2005,In_957,In_866);
nor U2006 (N_2006,In_124,In_1451);
nor U2007 (N_2007,In_1398,In_1381);
or U2008 (N_2008,In_932,In_1064);
and U2009 (N_2009,In_1144,In_296);
xor U2010 (N_2010,In_1091,In_1086);
nor U2011 (N_2011,In_972,In_1179);
nor U2012 (N_2012,In_279,In_1061);
nor U2013 (N_2013,In_825,In_1185);
nand U2014 (N_2014,In_1249,In_1364);
nor U2015 (N_2015,In_1325,In_612);
or U2016 (N_2016,In_1091,In_560);
and U2017 (N_2017,In_671,In_461);
and U2018 (N_2018,In_128,In_1499);
or U2019 (N_2019,In_921,In_531);
and U2020 (N_2020,In_1050,In_1041);
and U2021 (N_2021,In_376,In_475);
nand U2022 (N_2022,In_1006,In_1202);
nand U2023 (N_2023,In_1201,In_46);
nor U2024 (N_2024,In_543,In_333);
or U2025 (N_2025,In_607,In_1138);
and U2026 (N_2026,In_1422,In_484);
or U2027 (N_2027,In_516,In_709);
and U2028 (N_2028,In_984,In_425);
and U2029 (N_2029,In_1236,In_423);
or U2030 (N_2030,In_297,In_82);
and U2031 (N_2031,In_509,In_1454);
nor U2032 (N_2032,In_910,In_290);
or U2033 (N_2033,In_422,In_413);
or U2034 (N_2034,In_118,In_1467);
nor U2035 (N_2035,In_262,In_1088);
and U2036 (N_2036,In_1278,In_502);
and U2037 (N_2037,In_235,In_498);
or U2038 (N_2038,In_636,In_1136);
nand U2039 (N_2039,In_1458,In_721);
and U2040 (N_2040,In_280,In_1117);
nand U2041 (N_2041,In_464,In_274);
and U2042 (N_2042,In_1126,In_379);
nor U2043 (N_2043,In_844,In_63);
nand U2044 (N_2044,In_348,In_152);
or U2045 (N_2045,In_1355,In_1436);
and U2046 (N_2046,In_548,In_544);
xor U2047 (N_2047,In_442,In_407);
or U2048 (N_2048,In_562,In_86);
and U2049 (N_2049,In_1033,In_415);
nand U2050 (N_2050,In_777,In_1162);
and U2051 (N_2051,In_952,In_405);
nor U2052 (N_2052,In_50,In_767);
nand U2053 (N_2053,In_1044,In_214);
or U2054 (N_2054,In_1489,In_1479);
and U2055 (N_2055,In_1482,In_1213);
or U2056 (N_2056,In_466,In_366);
or U2057 (N_2057,In_1189,In_1486);
or U2058 (N_2058,In_1065,In_718);
nor U2059 (N_2059,In_1440,In_938);
nor U2060 (N_2060,In_1273,In_996);
nand U2061 (N_2061,In_1453,In_1023);
and U2062 (N_2062,In_348,In_1006);
or U2063 (N_2063,In_1093,In_626);
nor U2064 (N_2064,In_992,In_404);
nor U2065 (N_2065,In_739,In_1310);
or U2066 (N_2066,In_933,In_735);
nand U2067 (N_2067,In_678,In_227);
or U2068 (N_2068,In_136,In_394);
nor U2069 (N_2069,In_216,In_61);
nand U2070 (N_2070,In_1268,In_74);
or U2071 (N_2071,In_212,In_736);
xor U2072 (N_2072,In_478,In_992);
nor U2073 (N_2073,In_113,In_450);
and U2074 (N_2074,In_1350,In_1269);
nor U2075 (N_2075,In_444,In_1400);
or U2076 (N_2076,In_404,In_758);
or U2077 (N_2077,In_358,In_1279);
or U2078 (N_2078,In_998,In_542);
nand U2079 (N_2079,In_935,In_473);
nand U2080 (N_2080,In_367,In_978);
or U2081 (N_2081,In_716,In_797);
or U2082 (N_2082,In_1436,In_679);
and U2083 (N_2083,In_1384,In_57);
and U2084 (N_2084,In_44,In_243);
nor U2085 (N_2085,In_1041,In_178);
nor U2086 (N_2086,In_679,In_1001);
nand U2087 (N_2087,In_900,In_1311);
and U2088 (N_2088,In_90,In_555);
nor U2089 (N_2089,In_918,In_1284);
nand U2090 (N_2090,In_298,In_1049);
nor U2091 (N_2091,In_166,In_451);
and U2092 (N_2092,In_342,In_321);
nor U2093 (N_2093,In_351,In_1074);
nand U2094 (N_2094,In_55,In_1300);
and U2095 (N_2095,In_931,In_206);
nor U2096 (N_2096,In_1206,In_1241);
nor U2097 (N_2097,In_1494,In_1085);
or U2098 (N_2098,In_607,In_688);
nand U2099 (N_2099,In_937,In_635);
or U2100 (N_2100,In_246,In_785);
or U2101 (N_2101,In_1297,In_1188);
or U2102 (N_2102,In_240,In_207);
nand U2103 (N_2103,In_235,In_804);
or U2104 (N_2104,In_688,In_549);
or U2105 (N_2105,In_251,In_1276);
and U2106 (N_2106,In_818,In_157);
nand U2107 (N_2107,In_340,In_85);
and U2108 (N_2108,In_1088,In_672);
nor U2109 (N_2109,In_1005,In_1453);
or U2110 (N_2110,In_64,In_646);
nor U2111 (N_2111,In_5,In_393);
nand U2112 (N_2112,In_485,In_1098);
or U2113 (N_2113,In_1269,In_203);
nor U2114 (N_2114,In_1493,In_1019);
and U2115 (N_2115,In_1275,In_973);
or U2116 (N_2116,In_864,In_110);
or U2117 (N_2117,In_1239,In_124);
nor U2118 (N_2118,In_641,In_4);
and U2119 (N_2119,In_1301,In_473);
or U2120 (N_2120,In_1075,In_926);
nor U2121 (N_2121,In_218,In_999);
nor U2122 (N_2122,In_1400,In_195);
nand U2123 (N_2123,In_272,In_815);
and U2124 (N_2124,In_1397,In_312);
or U2125 (N_2125,In_1051,In_800);
nor U2126 (N_2126,In_1433,In_195);
and U2127 (N_2127,In_756,In_470);
nor U2128 (N_2128,In_1172,In_387);
and U2129 (N_2129,In_394,In_1353);
nand U2130 (N_2130,In_982,In_861);
or U2131 (N_2131,In_899,In_1230);
nor U2132 (N_2132,In_505,In_348);
nand U2133 (N_2133,In_1302,In_930);
and U2134 (N_2134,In_1184,In_222);
and U2135 (N_2135,In_1030,In_1251);
xor U2136 (N_2136,In_1101,In_1463);
and U2137 (N_2137,In_320,In_1085);
or U2138 (N_2138,In_44,In_1181);
nor U2139 (N_2139,In_734,In_451);
nand U2140 (N_2140,In_387,In_1382);
or U2141 (N_2141,In_1444,In_389);
and U2142 (N_2142,In_472,In_55);
nand U2143 (N_2143,In_918,In_970);
xnor U2144 (N_2144,In_501,In_632);
or U2145 (N_2145,In_1270,In_479);
nand U2146 (N_2146,In_1015,In_195);
and U2147 (N_2147,In_1216,In_196);
and U2148 (N_2148,In_1247,In_1046);
nand U2149 (N_2149,In_793,In_161);
nand U2150 (N_2150,In_110,In_10);
or U2151 (N_2151,In_183,In_776);
nor U2152 (N_2152,In_583,In_403);
and U2153 (N_2153,In_1119,In_586);
nand U2154 (N_2154,In_529,In_825);
or U2155 (N_2155,In_259,In_377);
and U2156 (N_2156,In_514,In_547);
or U2157 (N_2157,In_510,In_809);
and U2158 (N_2158,In_735,In_1320);
or U2159 (N_2159,In_266,In_1240);
nand U2160 (N_2160,In_628,In_736);
nand U2161 (N_2161,In_843,In_195);
and U2162 (N_2162,In_618,In_605);
nand U2163 (N_2163,In_277,In_352);
nor U2164 (N_2164,In_61,In_1107);
and U2165 (N_2165,In_604,In_524);
nand U2166 (N_2166,In_168,In_1218);
and U2167 (N_2167,In_118,In_1479);
nand U2168 (N_2168,In_224,In_90);
and U2169 (N_2169,In_421,In_808);
and U2170 (N_2170,In_824,In_845);
or U2171 (N_2171,In_1024,In_201);
or U2172 (N_2172,In_826,In_441);
or U2173 (N_2173,In_749,In_922);
or U2174 (N_2174,In_1294,In_1048);
or U2175 (N_2175,In_810,In_597);
nand U2176 (N_2176,In_693,In_950);
or U2177 (N_2177,In_256,In_132);
nand U2178 (N_2178,In_646,In_1465);
nor U2179 (N_2179,In_1331,In_450);
nand U2180 (N_2180,In_1298,In_806);
nand U2181 (N_2181,In_1401,In_551);
nand U2182 (N_2182,In_1195,In_639);
or U2183 (N_2183,In_526,In_635);
nand U2184 (N_2184,In_1398,In_540);
or U2185 (N_2185,In_1185,In_233);
and U2186 (N_2186,In_429,In_200);
or U2187 (N_2187,In_105,In_388);
or U2188 (N_2188,In_1272,In_138);
nor U2189 (N_2189,In_290,In_346);
or U2190 (N_2190,In_1289,In_261);
nor U2191 (N_2191,In_667,In_76);
and U2192 (N_2192,In_732,In_562);
and U2193 (N_2193,In_729,In_1055);
or U2194 (N_2194,In_225,In_102);
or U2195 (N_2195,In_164,In_1028);
or U2196 (N_2196,In_1225,In_1086);
and U2197 (N_2197,In_857,In_247);
nand U2198 (N_2198,In_1276,In_1044);
and U2199 (N_2199,In_68,In_412);
nor U2200 (N_2200,In_322,In_1310);
nand U2201 (N_2201,In_555,In_1286);
nor U2202 (N_2202,In_1037,In_714);
nor U2203 (N_2203,In_548,In_543);
and U2204 (N_2204,In_684,In_6);
nand U2205 (N_2205,In_888,In_1498);
and U2206 (N_2206,In_477,In_102);
or U2207 (N_2207,In_501,In_1478);
nand U2208 (N_2208,In_639,In_808);
or U2209 (N_2209,In_86,In_1288);
or U2210 (N_2210,In_118,In_1033);
nor U2211 (N_2211,In_159,In_761);
nor U2212 (N_2212,In_643,In_228);
or U2213 (N_2213,In_1028,In_1220);
or U2214 (N_2214,In_549,In_488);
nand U2215 (N_2215,In_1337,In_1246);
or U2216 (N_2216,In_928,In_497);
nor U2217 (N_2217,In_909,In_1212);
or U2218 (N_2218,In_1223,In_196);
nor U2219 (N_2219,In_309,In_390);
nand U2220 (N_2220,In_282,In_335);
nor U2221 (N_2221,In_1174,In_1314);
nor U2222 (N_2222,In_721,In_264);
or U2223 (N_2223,In_1016,In_508);
and U2224 (N_2224,In_1042,In_1073);
nor U2225 (N_2225,In_1294,In_637);
and U2226 (N_2226,In_555,In_369);
or U2227 (N_2227,In_792,In_1330);
and U2228 (N_2228,In_250,In_1418);
nand U2229 (N_2229,In_323,In_251);
or U2230 (N_2230,In_537,In_1296);
nand U2231 (N_2231,In_1162,In_1410);
nand U2232 (N_2232,In_299,In_1158);
nand U2233 (N_2233,In_949,In_1065);
and U2234 (N_2234,In_837,In_1329);
nor U2235 (N_2235,In_899,In_916);
nand U2236 (N_2236,In_661,In_454);
and U2237 (N_2237,In_1208,In_20);
or U2238 (N_2238,In_1118,In_114);
or U2239 (N_2239,In_1049,In_747);
and U2240 (N_2240,In_659,In_1);
and U2241 (N_2241,In_1484,In_1166);
and U2242 (N_2242,In_1017,In_854);
nand U2243 (N_2243,In_869,In_1489);
nand U2244 (N_2244,In_1413,In_1012);
and U2245 (N_2245,In_481,In_444);
nand U2246 (N_2246,In_700,In_1283);
or U2247 (N_2247,In_379,In_742);
or U2248 (N_2248,In_1091,In_1253);
and U2249 (N_2249,In_686,In_1496);
and U2250 (N_2250,In_1060,In_610);
or U2251 (N_2251,In_732,In_77);
xor U2252 (N_2252,In_1275,In_931);
nor U2253 (N_2253,In_298,In_577);
nor U2254 (N_2254,In_499,In_1105);
or U2255 (N_2255,In_1142,In_268);
or U2256 (N_2256,In_697,In_376);
xnor U2257 (N_2257,In_150,In_701);
and U2258 (N_2258,In_1082,In_153);
or U2259 (N_2259,In_303,In_452);
nand U2260 (N_2260,In_917,In_1134);
and U2261 (N_2261,In_75,In_873);
nand U2262 (N_2262,In_1476,In_472);
and U2263 (N_2263,In_1023,In_896);
or U2264 (N_2264,In_1454,In_239);
or U2265 (N_2265,In_981,In_1058);
and U2266 (N_2266,In_951,In_664);
and U2267 (N_2267,In_1371,In_51);
nor U2268 (N_2268,In_1104,In_668);
nor U2269 (N_2269,In_275,In_765);
or U2270 (N_2270,In_1360,In_814);
or U2271 (N_2271,In_1220,In_305);
and U2272 (N_2272,In_1147,In_875);
and U2273 (N_2273,In_624,In_1235);
and U2274 (N_2274,In_1291,In_810);
nand U2275 (N_2275,In_314,In_946);
nand U2276 (N_2276,In_153,In_814);
nor U2277 (N_2277,In_114,In_1120);
and U2278 (N_2278,In_1366,In_248);
xor U2279 (N_2279,In_876,In_520);
and U2280 (N_2280,In_926,In_1488);
nand U2281 (N_2281,In_961,In_1063);
nand U2282 (N_2282,In_382,In_1261);
nand U2283 (N_2283,In_1223,In_1018);
and U2284 (N_2284,In_691,In_1083);
or U2285 (N_2285,In_730,In_1431);
nand U2286 (N_2286,In_1388,In_1420);
or U2287 (N_2287,In_356,In_1498);
and U2288 (N_2288,In_1414,In_820);
or U2289 (N_2289,In_378,In_242);
and U2290 (N_2290,In_1463,In_1467);
xor U2291 (N_2291,In_35,In_1015);
nor U2292 (N_2292,In_1117,In_289);
or U2293 (N_2293,In_462,In_1044);
nor U2294 (N_2294,In_780,In_702);
and U2295 (N_2295,In_1392,In_395);
and U2296 (N_2296,In_864,In_253);
or U2297 (N_2297,In_840,In_137);
nand U2298 (N_2298,In_520,In_206);
nor U2299 (N_2299,In_1198,In_1025);
or U2300 (N_2300,In_438,In_945);
nand U2301 (N_2301,In_1457,In_350);
or U2302 (N_2302,In_585,In_1312);
nor U2303 (N_2303,In_856,In_301);
nand U2304 (N_2304,In_202,In_1418);
and U2305 (N_2305,In_335,In_542);
or U2306 (N_2306,In_918,In_446);
or U2307 (N_2307,In_1009,In_1088);
or U2308 (N_2308,In_284,In_1370);
and U2309 (N_2309,In_306,In_675);
nand U2310 (N_2310,In_39,In_1333);
and U2311 (N_2311,In_605,In_507);
and U2312 (N_2312,In_1211,In_873);
nand U2313 (N_2313,In_1277,In_945);
nor U2314 (N_2314,In_1064,In_901);
nand U2315 (N_2315,In_171,In_1291);
nand U2316 (N_2316,In_1479,In_144);
and U2317 (N_2317,In_853,In_968);
and U2318 (N_2318,In_634,In_123);
nand U2319 (N_2319,In_536,In_688);
and U2320 (N_2320,In_330,In_974);
or U2321 (N_2321,In_563,In_174);
or U2322 (N_2322,In_576,In_1431);
nor U2323 (N_2323,In_862,In_525);
nand U2324 (N_2324,In_1144,In_368);
or U2325 (N_2325,In_440,In_485);
nor U2326 (N_2326,In_1190,In_1083);
or U2327 (N_2327,In_1076,In_211);
or U2328 (N_2328,In_797,In_413);
nand U2329 (N_2329,In_231,In_1182);
nor U2330 (N_2330,In_256,In_1465);
and U2331 (N_2331,In_592,In_1305);
nand U2332 (N_2332,In_43,In_165);
or U2333 (N_2333,In_591,In_1041);
and U2334 (N_2334,In_132,In_1187);
nor U2335 (N_2335,In_125,In_804);
and U2336 (N_2336,In_254,In_127);
and U2337 (N_2337,In_1050,In_113);
nand U2338 (N_2338,In_1405,In_1173);
and U2339 (N_2339,In_903,In_1028);
or U2340 (N_2340,In_940,In_1126);
and U2341 (N_2341,In_350,In_51);
nor U2342 (N_2342,In_1448,In_1102);
and U2343 (N_2343,In_489,In_1091);
or U2344 (N_2344,In_779,In_544);
nor U2345 (N_2345,In_1422,In_590);
and U2346 (N_2346,In_1301,In_1149);
and U2347 (N_2347,In_490,In_1138);
nor U2348 (N_2348,In_973,In_398);
nor U2349 (N_2349,In_115,In_24);
and U2350 (N_2350,In_1220,In_582);
nor U2351 (N_2351,In_177,In_1355);
and U2352 (N_2352,In_1013,In_1128);
nor U2353 (N_2353,In_227,In_7);
nor U2354 (N_2354,In_643,In_346);
nand U2355 (N_2355,In_599,In_1034);
nor U2356 (N_2356,In_524,In_1140);
nand U2357 (N_2357,In_760,In_318);
nand U2358 (N_2358,In_744,In_847);
or U2359 (N_2359,In_785,In_42);
or U2360 (N_2360,In_1409,In_1074);
or U2361 (N_2361,In_555,In_732);
and U2362 (N_2362,In_80,In_299);
nand U2363 (N_2363,In_1321,In_1152);
and U2364 (N_2364,In_467,In_1051);
nor U2365 (N_2365,In_899,In_1497);
or U2366 (N_2366,In_438,In_801);
and U2367 (N_2367,In_415,In_696);
nor U2368 (N_2368,In_926,In_1330);
nor U2369 (N_2369,In_510,In_604);
and U2370 (N_2370,In_1085,In_1301);
and U2371 (N_2371,In_781,In_330);
xnor U2372 (N_2372,In_570,In_1392);
nor U2373 (N_2373,In_477,In_949);
nand U2374 (N_2374,In_1445,In_1060);
and U2375 (N_2375,In_277,In_372);
nor U2376 (N_2376,In_468,In_229);
and U2377 (N_2377,In_516,In_1066);
or U2378 (N_2378,In_561,In_1136);
or U2379 (N_2379,In_338,In_663);
nand U2380 (N_2380,In_71,In_1079);
nand U2381 (N_2381,In_362,In_1010);
or U2382 (N_2382,In_438,In_838);
and U2383 (N_2383,In_1169,In_987);
and U2384 (N_2384,In_277,In_1410);
nand U2385 (N_2385,In_890,In_708);
and U2386 (N_2386,In_1280,In_512);
nand U2387 (N_2387,In_73,In_928);
or U2388 (N_2388,In_626,In_565);
nor U2389 (N_2389,In_585,In_1478);
nand U2390 (N_2390,In_440,In_628);
or U2391 (N_2391,In_1490,In_853);
and U2392 (N_2392,In_1353,In_1295);
or U2393 (N_2393,In_759,In_553);
and U2394 (N_2394,In_30,In_401);
nor U2395 (N_2395,In_1497,In_274);
and U2396 (N_2396,In_1337,In_680);
nor U2397 (N_2397,In_260,In_1086);
or U2398 (N_2398,In_1183,In_213);
and U2399 (N_2399,In_1045,In_1001);
and U2400 (N_2400,In_459,In_920);
nand U2401 (N_2401,In_712,In_1168);
nand U2402 (N_2402,In_556,In_1199);
nor U2403 (N_2403,In_182,In_1396);
nand U2404 (N_2404,In_852,In_183);
nor U2405 (N_2405,In_1338,In_592);
nor U2406 (N_2406,In_11,In_316);
and U2407 (N_2407,In_1046,In_631);
nand U2408 (N_2408,In_76,In_1326);
or U2409 (N_2409,In_340,In_54);
nand U2410 (N_2410,In_449,In_715);
or U2411 (N_2411,In_1116,In_347);
or U2412 (N_2412,In_1497,In_1083);
or U2413 (N_2413,In_1281,In_136);
or U2414 (N_2414,In_794,In_775);
nand U2415 (N_2415,In_689,In_30);
nand U2416 (N_2416,In_740,In_695);
or U2417 (N_2417,In_36,In_1294);
nor U2418 (N_2418,In_510,In_1329);
or U2419 (N_2419,In_1410,In_1011);
or U2420 (N_2420,In_834,In_1187);
nand U2421 (N_2421,In_1158,In_527);
nand U2422 (N_2422,In_833,In_1039);
nand U2423 (N_2423,In_382,In_712);
nand U2424 (N_2424,In_288,In_275);
or U2425 (N_2425,In_693,In_229);
nand U2426 (N_2426,In_1371,In_281);
nor U2427 (N_2427,In_1065,In_89);
nand U2428 (N_2428,In_1193,In_170);
nand U2429 (N_2429,In_256,In_1089);
and U2430 (N_2430,In_1090,In_1460);
and U2431 (N_2431,In_7,In_254);
or U2432 (N_2432,In_1277,In_63);
or U2433 (N_2433,In_40,In_56);
nor U2434 (N_2434,In_851,In_1025);
or U2435 (N_2435,In_717,In_654);
nor U2436 (N_2436,In_1155,In_977);
nand U2437 (N_2437,In_1385,In_1211);
and U2438 (N_2438,In_514,In_1274);
or U2439 (N_2439,In_1191,In_821);
nor U2440 (N_2440,In_1308,In_1066);
or U2441 (N_2441,In_1035,In_505);
nor U2442 (N_2442,In_1403,In_738);
and U2443 (N_2443,In_1029,In_329);
and U2444 (N_2444,In_1012,In_352);
nand U2445 (N_2445,In_256,In_1313);
nor U2446 (N_2446,In_1327,In_1060);
nor U2447 (N_2447,In_430,In_907);
or U2448 (N_2448,In_527,In_851);
and U2449 (N_2449,In_48,In_1388);
nand U2450 (N_2450,In_58,In_1216);
nor U2451 (N_2451,In_178,In_416);
nor U2452 (N_2452,In_66,In_455);
nand U2453 (N_2453,In_1370,In_1428);
or U2454 (N_2454,In_459,In_1318);
or U2455 (N_2455,In_1417,In_774);
and U2456 (N_2456,In_700,In_592);
or U2457 (N_2457,In_393,In_674);
nor U2458 (N_2458,In_489,In_1462);
or U2459 (N_2459,In_1074,In_829);
or U2460 (N_2460,In_1293,In_1448);
or U2461 (N_2461,In_833,In_1473);
nor U2462 (N_2462,In_478,In_599);
or U2463 (N_2463,In_745,In_318);
or U2464 (N_2464,In_457,In_1313);
nor U2465 (N_2465,In_282,In_887);
nand U2466 (N_2466,In_584,In_525);
or U2467 (N_2467,In_1255,In_1262);
and U2468 (N_2468,In_1210,In_858);
and U2469 (N_2469,In_1453,In_1477);
nor U2470 (N_2470,In_348,In_1482);
and U2471 (N_2471,In_974,In_610);
or U2472 (N_2472,In_1277,In_1149);
or U2473 (N_2473,In_1387,In_99);
and U2474 (N_2474,In_248,In_1141);
nor U2475 (N_2475,In_17,In_824);
or U2476 (N_2476,In_1035,In_517);
and U2477 (N_2477,In_1432,In_909);
or U2478 (N_2478,In_107,In_737);
and U2479 (N_2479,In_1304,In_1000);
nor U2480 (N_2480,In_277,In_291);
or U2481 (N_2481,In_383,In_1232);
and U2482 (N_2482,In_1325,In_1076);
or U2483 (N_2483,In_614,In_60);
and U2484 (N_2484,In_360,In_285);
nor U2485 (N_2485,In_1030,In_45);
nand U2486 (N_2486,In_689,In_669);
nand U2487 (N_2487,In_442,In_1066);
or U2488 (N_2488,In_1070,In_319);
and U2489 (N_2489,In_951,In_33);
nor U2490 (N_2490,In_1423,In_284);
nand U2491 (N_2491,In_783,In_1034);
and U2492 (N_2492,In_900,In_1120);
or U2493 (N_2493,In_66,In_149);
or U2494 (N_2494,In_803,In_276);
nor U2495 (N_2495,In_359,In_222);
nor U2496 (N_2496,In_378,In_673);
or U2497 (N_2497,In_116,In_1291);
nand U2498 (N_2498,In_1290,In_266);
or U2499 (N_2499,In_323,In_200);
or U2500 (N_2500,In_1208,In_1292);
or U2501 (N_2501,In_572,In_463);
nand U2502 (N_2502,In_895,In_1396);
nand U2503 (N_2503,In_373,In_1092);
nand U2504 (N_2504,In_129,In_116);
or U2505 (N_2505,In_764,In_174);
nor U2506 (N_2506,In_1214,In_600);
or U2507 (N_2507,In_335,In_1171);
nand U2508 (N_2508,In_1235,In_798);
nand U2509 (N_2509,In_596,In_1261);
and U2510 (N_2510,In_661,In_136);
nand U2511 (N_2511,In_1383,In_700);
nor U2512 (N_2512,In_1323,In_1244);
nand U2513 (N_2513,In_618,In_1363);
nand U2514 (N_2514,In_814,In_275);
nor U2515 (N_2515,In_1044,In_1434);
or U2516 (N_2516,In_111,In_445);
nor U2517 (N_2517,In_1449,In_1274);
and U2518 (N_2518,In_1438,In_894);
nand U2519 (N_2519,In_835,In_1184);
or U2520 (N_2520,In_482,In_1461);
nor U2521 (N_2521,In_569,In_548);
and U2522 (N_2522,In_166,In_507);
or U2523 (N_2523,In_374,In_1002);
nor U2524 (N_2524,In_1257,In_1154);
nor U2525 (N_2525,In_60,In_631);
nor U2526 (N_2526,In_995,In_989);
or U2527 (N_2527,In_72,In_713);
nor U2528 (N_2528,In_43,In_698);
nor U2529 (N_2529,In_961,In_772);
and U2530 (N_2530,In_1283,In_701);
nor U2531 (N_2531,In_783,In_1242);
and U2532 (N_2532,In_816,In_1049);
or U2533 (N_2533,In_700,In_1379);
or U2534 (N_2534,In_1360,In_925);
nor U2535 (N_2535,In_1177,In_901);
or U2536 (N_2536,In_266,In_1188);
nand U2537 (N_2537,In_1370,In_136);
and U2538 (N_2538,In_858,In_1171);
and U2539 (N_2539,In_1318,In_913);
nor U2540 (N_2540,In_50,In_910);
or U2541 (N_2541,In_399,In_1480);
or U2542 (N_2542,In_585,In_239);
or U2543 (N_2543,In_793,In_900);
and U2544 (N_2544,In_749,In_1424);
nor U2545 (N_2545,In_1491,In_1035);
nand U2546 (N_2546,In_1000,In_1232);
nand U2547 (N_2547,In_1132,In_195);
nor U2548 (N_2548,In_862,In_213);
nand U2549 (N_2549,In_1452,In_864);
or U2550 (N_2550,In_400,In_1227);
or U2551 (N_2551,In_814,In_682);
or U2552 (N_2552,In_1072,In_505);
nor U2553 (N_2553,In_1062,In_295);
and U2554 (N_2554,In_38,In_845);
or U2555 (N_2555,In_995,In_819);
and U2556 (N_2556,In_211,In_868);
nand U2557 (N_2557,In_33,In_286);
nor U2558 (N_2558,In_1084,In_1451);
or U2559 (N_2559,In_481,In_1280);
nand U2560 (N_2560,In_790,In_209);
nand U2561 (N_2561,In_940,In_1194);
xor U2562 (N_2562,In_965,In_238);
xor U2563 (N_2563,In_962,In_991);
nand U2564 (N_2564,In_741,In_7);
or U2565 (N_2565,In_1089,In_1407);
nor U2566 (N_2566,In_1290,In_1245);
or U2567 (N_2567,In_319,In_786);
and U2568 (N_2568,In_860,In_1064);
nor U2569 (N_2569,In_1178,In_1336);
or U2570 (N_2570,In_1417,In_32);
nand U2571 (N_2571,In_798,In_1372);
nand U2572 (N_2572,In_954,In_115);
nor U2573 (N_2573,In_532,In_401);
and U2574 (N_2574,In_393,In_1422);
and U2575 (N_2575,In_356,In_1201);
nand U2576 (N_2576,In_1426,In_400);
and U2577 (N_2577,In_1161,In_191);
or U2578 (N_2578,In_18,In_25);
and U2579 (N_2579,In_1494,In_175);
or U2580 (N_2580,In_786,In_1105);
nor U2581 (N_2581,In_1192,In_1488);
or U2582 (N_2582,In_1238,In_823);
nand U2583 (N_2583,In_866,In_1192);
nor U2584 (N_2584,In_1092,In_172);
and U2585 (N_2585,In_1081,In_1289);
and U2586 (N_2586,In_1035,In_358);
xor U2587 (N_2587,In_395,In_385);
or U2588 (N_2588,In_481,In_361);
nor U2589 (N_2589,In_1406,In_578);
nand U2590 (N_2590,In_452,In_656);
or U2591 (N_2591,In_1261,In_522);
or U2592 (N_2592,In_1374,In_171);
nand U2593 (N_2593,In_619,In_498);
nor U2594 (N_2594,In_26,In_1062);
nor U2595 (N_2595,In_1175,In_1210);
and U2596 (N_2596,In_1439,In_463);
nor U2597 (N_2597,In_246,In_991);
nor U2598 (N_2598,In_599,In_1465);
and U2599 (N_2599,In_114,In_1071);
or U2600 (N_2600,In_1499,In_1255);
nor U2601 (N_2601,In_695,In_800);
nand U2602 (N_2602,In_1089,In_816);
nand U2603 (N_2603,In_1443,In_596);
or U2604 (N_2604,In_1370,In_849);
and U2605 (N_2605,In_51,In_377);
and U2606 (N_2606,In_613,In_332);
nand U2607 (N_2607,In_1197,In_130);
nand U2608 (N_2608,In_396,In_268);
nand U2609 (N_2609,In_141,In_88);
or U2610 (N_2610,In_1164,In_762);
and U2611 (N_2611,In_970,In_1386);
or U2612 (N_2612,In_1250,In_1349);
and U2613 (N_2613,In_713,In_577);
and U2614 (N_2614,In_855,In_1018);
and U2615 (N_2615,In_35,In_1436);
and U2616 (N_2616,In_300,In_1067);
and U2617 (N_2617,In_1254,In_1498);
and U2618 (N_2618,In_1368,In_839);
or U2619 (N_2619,In_1099,In_993);
nor U2620 (N_2620,In_1459,In_782);
nand U2621 (N_2621,In_424,In_773);
nor U2622 (N_2622,In_234,In_32);
nor U2623 (N_2623,In_548,In_349);
and U2624 (N_2624,In_1404,In_1245);
nand U2625 (N_2625,In_557,In_422);
nor U2626 (N_2626,In_234,In_1199);
nor U2627 (N_2627,In_7,In_35);
or U2628 (N_2628,In_700,In_954);
nand U2629 (N_2629,In_739,In_1170);
xor U2630 (N_2630,In_1033,In_222);
nand U2631 (N_2631,In_599,In_1331);
and U2632 (N_2632,In_515,In_260);
nor U2633 (N_2633,In_641,In_377);
or U2634 (N_2634,In_269,In_474);
nor U2635 (N_2635,In_749,In_780);
or U2636 (N_2636,In_1279,In_1286);
or U2637 (N_2637,In_1470,In_1022);
and U2638 (N_2638,In_614,In_673);
or U2639 (N_2639,In_1197,In_231);
and U2640 (N_2640,In_542,In_1432);
nor U2641 (N_2641,In_514,In_1128);
or U2642 (N_2642,In_843,In_802);
and U2643 (N_2643,In_1444,In_566);
nand U2644 (N_2644,In_598,In_943);
nand U2645 (N_2645,In_429,In_1136);
nor U2646 (N_2646,In_1284,In_1414);
and U2647 (N_2647,In_740,In_778);
nand U2648 (N_2648,In_969,In_1402);
nand U2649 (N_2649,In_94,In_95);
nand U2650 (N_2650,In_710,In_1099);
and U2651 (N_2651,In_350,In_983);
or U2652 (N_2652,In_1150,In_853);
nor U2653 (N_2653,In_593,In_1010);
nor U2654 (N_2654,In_124,In_496);
or U2655 (N_2655,In_918,In_721);
nand U2656 (N_2656,In_1399,In_1042);
and U2657 (N_2657,In_869,In_1440);
or U2658 (N_2658,In_1179,In_8);
and U2659 (N_2659,In_693,In_87);
nor U2660 (N_2660,In_694,In_1463);
nor U2661 (N_2661,In_375,In_155);
nor U2662 (N_2662,In_926,In_728);
nor U2663 (N_2663,In_438,In_1463);
or U2664 (N_2664,In_1008,In_1177);
and U2665 (N_2665,In_938,In_117);
xor U2666 (N_2666,In_1199,In_917);
or U2667 (N_2667,In_482,In_467);
and U2668 (N_2668,In_1423,In_1452);
or U2669 (N_2669,In_1498,In_55);
nand U2670 (N_2670,In_452,In_1484);
and U2671 (N_2671,In_161,In_244);
nor U2672 (N_2672,In_1400,In_483);
and U2673 (N_2673,In_166,In_762);
nor U2674 (N_2674,In_885,In_477);
nand U2675 (N_2675,In_366,In_1475);
nand U2676 (N_2676,In_155,In_588);
nor U2677 (N_2677,In_62,In_73);
nand U2678 (N_2678,In_95,In_1422);
or U2679 (N_2679,In_1082,In_453);
nor U2680 (N_2680,In_1401,In_861);
nand U2681 (N_2681,In_679,In_693);
or U2682 (N_2682,In_443,In_1449);
nand U2683 (N_2683,In_190,In_191);
or U2684 (N_2684,In_775,In_538);
nand U2685 (N_2685,In_1376,In_666);
and U2686 (N_2686,In_832,In_85);
nand U2687 (N_2687,In_892,In_1383);
nand U2688 (N_2688,In_1274,In_1153);
nor U2689 (N_2689,In_451,In_1124);
nor U2690 (N_2690,In_1136,In_1176);
nand U2691 (N_2691,In_1195,In_706);
or U2692 (N_2692,In_1320,In_1272);
nand U2693 (N_2693,In_984,In_833);
and U2694 (N_2694,In_30,In_863);
or U2695 (N_2695,In_747,In_249);
and U2696 (N_2696,In_1302,In_786);
nand U2697 (N_2697,In_686,In_296);
nand U2698 (N_2698,In_806,In_1195);
nand U2699 (N_2699,In_378,In_626);
nand U2700 (N_2700,In_1097,In_710);
nand U2701 (N_2701,In_341,In_1160);
nor U2702 (N_2702,In_679,In_821);
and U2703 (N_2703,In_150,In_1109);
nor U2704 (N_2704,In_554,In_1272);
or U2705 (N_2705,In_167,In_472);
and U2706 (N_2706,In_223,In_77);
or U2707 (N_2707,In_654,In_634);
or U2708 (N_2708,In_1200,In_437);
and U2709 (N_2709,In_996,In_247);
nor U2710 (N_2710,In_222,In_497);
and U2711 (N_2711,In_654,In_887);
or U2712 (N_2712,In_190,In_882);
xnor U2713 (N_2713,In_1475,In_548);
nor U2714 (N_2714,In_719,In_98);
or U2715 (N_2715,In_976,In_347);
and U2716 (N_2716,In_254,In_345);
nor U2717 (N_2717,In_396,In_616);
or U2718 (N_2718,In_1463,In_254);
nand U2719 (N_2719,In_1407,In_95);
and U2720 (N_2720,In_912,In_949);
or U2721 (N_2721,In_1296,In_253);
nor U2722 (N_2722,In_41,In_429);
and U2723 (N_2723,In_809,In_1371);
nand U2724 (N_2724,In_1044,In_721);
nor U2725 (N_2725,In_627,In_93);
nor U2726 (N_2726,In_1238,In_555);
nor U2727 (N_2727,In_549,In_256);
nor U2728 (N_2728,In_680,In_1363);
and U2729 (N_2729,In_437,In_1376);
xnor U2730 (N_2730,In_892,In_476);
or U2731 (N_2731,In_394,In_222);
or U2732 (N_2732,In_219,In_1384);
nor U2733 (N_2733,In_967,In_520);
or U2734 (N_2734,In_138,In_377);
nor U2735 (N_2735,In_964,In_1363);
nor U2736 (N_2736,In_469,In_939);
nand U2737 (N_2737,In_344,In_1364);
or U2738 (N_2738,In_471,In_304);
and U2739 (N_2739,In_1480,In_1360);
nand U2740 (N_2740,In_1160,In_230);
nand U2741 (N_2741,In_773,In_474);
nand U2742 (N_2742,In_712,In_90);
nand U2743 (N_2743,In_670,In_247);
nand U2744 (N_2744,In_417,In_1146);
nand U2745 (N_2745,In_258,In_749);
and U2746 (N_2746,In_283,In_1107);
or U2747 (N_2747,In_1296,In_518);
nor U2748 (N_2748,In_520,In_86);
and U2749 (N_2749,In_259,In_1301);
nor U2750 (N_2750,In_1125,In_392);
and U2751 (N_2751,In_175,In_185);
or U2752 (N_2752,In_708,In_568);
and U2753 (N_2753,In_1218,In_20);
or U2754 (N_2754,In_698,In_767);
or U2755 (N_2755,In_9,In_316);
nand U2756 (N_2756,In_720,In_163);
or U2757 (N_2757,In_388,In_936);
or U2758 (N_2758,In_141,In_960);
or U2759 (N_2759,In_489,In_154);
nand U2760 (N_2760,In_1306,In_638);
or U2761 (N_2761,In_1037,In_1439);
nor U2762 (N_2762,In_791,In_509);
nor U2763 (N_2763,In_184,In_1171);
nor U2764 (N_2764,In_75,In_718);
or U2765 (N_2765,In_1268,In_96);
and U2766 (N_2766,In_1420,In_1405);
xor U2767 (N_2767,In_86,In_585);
nand U2768 (N_2768,In_1468,In_1097);
and U2769 (N_2769,In_1029,In_38);
nand U2770 (N_2770,In_1011,In_1211);
nor U2771 (N_2771,In_784,In_320);
nand U2772 (N_2772,In_733,In_934);
and U2773 (N_2773,In_636,In_142);
nand U2774 (N_2774,In_1002,In_144);
or U2775 (N_2775,In_784,In_1245);
nor U2776 (N_2776,In_560,In_599);
and U2777 (N_2777,In_1043,In_1317);
nand U2778 (N_2778,In_490,In_464);
and U2779 (N_2779,In_1461,In_1120);
nor U2780 (N_2780,In_1027,In_596);
nor U2781 (N_2781,In_1110,In_1332);
nand U2782 (N_2782,In_426,In_17);
nand U2783 (N_2783,In_334,In_1484);
nor U2784 (N_2784,In_961,In_1051);
or U2785 (N_2785,In_313,In_588);
nor U2786 (N_2786,In_194,In_941);
and U2787 (N_2787,In_873,In_480);
nor U2788 (N_2788,In_321,In_340);
or U2789 (N_2789,In_748,In_1417);
nand U2790 (N_2790,In_411,In_686);
nand U2791 (N_2791,In_1082,In_465);
nor U2792 (N_2792,In_347,In_589);
nor U2793 (N_2793,In_492,In_1361);
and U2794 (N_2794,In_642,In_933);
nor U2795 (N_2795,In_644,In_328);
and U2796 (N_2796,In_6,In_791);
nand U2797 (N_2797,In_658,In_1013);
nand U2798 (N_2798,In_547,In_502);
or U2799 (N_2799,In_1050,In_1469);
nand U2800 (N_2800,In_472,In_619);
or U2801 (N_2801,In_280,In_1316);
and U2802 (N_2802,In_1186,In_279);
nand U2803 (N_2803,In_1059,In_789);
and U2804 (N_2804,In_290,In_102);
nand U2805 (N_2805,In_1188,In_109);
and U2806 (N_2806,In_562,In_1005);
or U2807 (N_2807,In_711,In_442);
and U2808 (N_2808,In_527,In_705);
nand U2809 (N_2809,In_384,In_448);
and U2810 (N_2810,In_852,In_1079);
and U2811 (N_2811,In_1214,In_171);
nor U2812 (N_2812,In_59,In_913);
and U2813 (N_2813,In_597,In_267);
nor U2814 (N_2814,In_652,In_85);
or U2815 (N_2815,In_198,In_265);
or U2816 (N_2816,In_67,In_252);
or U2817 (N_2817,In_1412,In_1488);
and U2818 (N_2818,In_833,In_499);
and U2819 (N_2819,In_368,In_1367);
nor U2820 (N_2820,In_1010,In_1228);
nor U2821 (N_2821,In_937,In_457);
nor U2822 (N_2822,In_220,In_479);
or U2823 (N_2823,In_941,In_136);
and U2824 (N_2824,In_251,In_1122);
nor U2825 (N_2825,In_608,In_68);
nand U2826 (N_2826,In_359,In_1241);
nor U2827 (N_2827,In_137,In_1349);
nand U2828 (N_2828,In_1049,In_1300);
nor U2829 (N_2829,In_1109,In_574);
or U2830 (N_2830,In_812,In_190);
and U2831 (N_2831,In_661,In_757);
and U2832 (N_2832,In_570,In_1268);
nand U2833 (N_2833,In_43,In_1458);
nand U2834 (N_2834,In_1198,In_189);
nand U2835 (N_2835,In_93,In_1095);
nor U2836 (N_2836,In_587,In_1107);
nor U2837 (N_2837,In_1272,In_799);
or U2838 (N_2838,In_648,In_1326);
and U2839 (N_2839,In_1409,In_1299);
or U2840 (N_2840,In_957,In_1464);
nand U2841 (N_2841,In_675,In_323);
nor U2842 (N_2842,In_982,In_1040);
nor U2843 (N_2843,In_274,In_847);
nor U2844 (N_2844,In_735,In_875);
nand U2845 (N_2845,In_1176,In_855);
or U2846 (N_2846,In_239,In_1261);
nor U2847 (N_2847,In_208,In_850);
nor U2848 (N_2848,In_1352,In_208);
or U2849 (N_2849,In_392,In_330);
and U2850 (N_2850,In_891,In_719);
and U2851 (N_2851,In_498,In_1361);
xnor U2852 (N_2852,In_1363,In_973);
nand U2853 (N_2853,In_21,In_599);
nor U2854 (N_2854,In_699,In_1381);
or U2855 (N_2855,In_973,In_1200);
and U2856 (N_2856,In_840,In_217);
and U2857 (N_2857,In_295,In_1319);
nor U2858 (N_2858,In_49,In_855);
nand U2859 (N_2859,In_165,In_1102);
and U2860 (N_2860,In_429,In_855);
nor U2861 (N_2861,In_1366,In_545);
or U2862 (N_2862,In_607,In_1068);
or U2863 (N_2863,In_952,In_593);
nand U2864 (N_2864,In_1431,In_485);
nor U2865 (N_2865,In_932,In_1298);
and U2866 (N_2866,In_1457,In_966);
and U2867 (N_2867,In_524,In_1349);
or U2868 (N_2868,In_1089,In_611);
nand U2869 (N_2869,In_333,In_246);
or U2870 (N_2870,In_440,In_663);
and U2871 (N_2871,In_1365,In_1136);
and U2872 (N_2872,In_77,In_115);
or U2873 (N_2873,In_941,In_750);
xnor U2874 (N_2874,In_424,In_973);
or U2875 (N_2875,In_29,In_827);
and U2876 (N_2876,In_162,In_241);
nor U2877 (N_2877,In_257,In_761);
nor U2878 (N_2878,In_842,In_400);
or U2879 (N_2879,In_1420,In_900);
nand U2880 (N_2880,In_1495,In_171);
nand U2881 (N_2881,In_884,In_1087);
or U2882 (N_2882,In_1116,In_677);
nor U2883 (N_2883,In_1264,In_1268);
nor U2884 (N_2884,In_235,In_974);
and U2885 (N_2885,In_1162,In_76);
nand U2886 (N_2886,In_111,In_399);
or U2887 (N_2887,In_1358,In_765);
and U2888 (N_2888,In_782,In_299);
and U2889 (N_2889,In_626,In_1064);
and U2890 (N_2890,In_275,In_60);
xor U2891 (N_2891,In_440,In_1384);
or U2892 (N_2892,In_1366,In_88);
or U2893 (N_2893,In_1469,In_630);
or U2894 (N_2894,In_376,In_1265);
and U2895 (N_2895,In_1120,In_732);
and U2896 (N_2896,In_393,In_1117);
and U2897 (N_2897,In_708,In_698);
and U2898 (N_2898,In_407,In_1426);
nand U2899 (N_2899,In_1061,In_1486);
and U2900 (N_2900,In_345,In_13);
nand U2901 (N_2901,In_1034,In_694);
and U2902 (N_2902,In_571,In_241);
nand U2903 (N_2903,In_96,In_888);
or U2904 (N_2904,In_444,In_1135);
nand U2905 (N_2905,In_678,In_649);
or U2906 (N_2906,In_431,In_818);
nor U2907 (N_2907,In_913,In_1425);
nand U2908 (N_2908,In_1119,In_1231);
nand U2909 (N_2909,In_1437,In_1160);
nand U2910 (N_2910,In_634,In_255);
and U2911 (N_2911,In_951,In_510);
nand U2912 (N_2912,In_1290,In_363);
and U2913 (N_2913,In_1388,In_1239);
nor U2914 (N_2914,In_216,In_561);
nand U2915 (N_2915,In_510,In_1407);
or U2916 (N_2916,In_300,In_340);
or U2917 (N_2917,In_185,In_753);
nand U2918 (N_2918,In_487,In_1308);
or U2919 (N_2919,In_341,In_806);
nand U2920 (N_2920,In_1217,In_1440);
or U2921 (N_2921,In_1112,In_1353);
nor U2922 (N_2922,In_1101,In_50);
nand U2923 (N_2923,In_186,In_1203);
nor U2924 (N_2924,In_990,In_434);
and U2925 (N_2925,In_1152,In_754);
nor U2926 (N_2926,In_486,In_1481);
nor U2927 (N_2927,In_1364,In_1102);
nor U2928 (N_2928,In_861,In_1044);
or U2929 (N_2929,In_168,In_524);
and U2930 (N_2930,In_336,In_180);
or U2931 (N_2931,In_901,In_1223);
and U2932 (N_2932,In_1021,In_987);
nand U2933 (N_2933,In_485,In_85);
and U2934 (N_2934,In_504,In_1132);
xnor U2935 (N_2935,In_1337,In_225);
and U2936 (N_2936,In_49,In_1284);
and U2937 (N_2937,In_204,In_281);
or U2938 (N_2938,In_62,In_1425);
or U2939 (N_2939,In_1496,In_391);
and U2940 (N_2940,In_495,In_667);
nand U2941 (N_2941,In_326,In_1272);
and U2942 (N_2942,In_911,In_360);
nand U2943 (N_2943,In_984,In_1365);
nand U2944 (N_2944,In_62,In_1328);
nand U2945 (N_2945,In_463,In_861);
nand U2946 (N_2946,In_1080,In_46);
nor U2947 (N_2947,In_1188,In_894);
nor U2948 (N_2948,In_431,In_1298);
and U2949 (N_2949,In_527,In_813);
or U2950 (N_2950,In_1336,In_1173);
and U2951 (N_2951,In_17,In_224);
nand U2952 (N_2952,In_1375,In_556);
or U2953 (N_2953,In_1186,In_978);
and U2954 (N_2954,In_210,In_403);
nand U2955 (N_2955,In_839,In_1310);
xnor U2956 (N_2956,In_1430,In_1160);
and U2957 (N_2957,In_1488,In_133);
or U2958 (N_2958,In_656,In_508);
nor U2959 (N_2959,In_198,In_1192);
and U2960 (N_2960,In_237,In_919);
or U2961 (N_2961,In_1051,In_808);
or U2962 (N_2962,In_942,In_305);
and U2963 (N_2963,In_61,In_693);
and U2964 (N_2964,In_406,In_62);
nand U2965 (N_2965,In_488,In_796);
or U2966 (N_2966,In_1435,In_1145);
nand U2967 (N_2967,In_585,In_1115);
and U2968 (N_2968,In_117,In_146);
or U2969 (N_2969,In_326,In_1013);
and U2970 (N_2970,In_665,In_1249);
nor U2971 (N_2971,In_679,In_1141);
and U2972 (N_2972,In_239,In_1444);
and U2973 (N_2973,In_1161,In_153);
and U2974 (N_2974,In_885,In_217);
or U2975 (N_2975,In_68,In_1463);
nor U2976 (N_2976,In_142,In_1424);
and U2977 (N_2977,In_959,In_548);
nor U2978 (N_2978,In_724,In_24);
nor U2979 (N_2979,In_1310,In_500);
nor U2980 (N_2980,In_46,In_725);
and U2981 (N_2981,In_939,In_666);
or U2982 (N_2982,In_1390,In_444);
or U2983 (N_2983,In_426,In_121);
and U2984 (N_2984,In_474,In_108);
or U2985 (N_2985,In_678,In_722);
and U2986 (N_2986,In_508,In_1206);
and U2987 (N_2987,In_1384,In_1359);
nand U2988 (N_2988,In_918,In_1471);
nor U2989 (N_2989,In_400,In_290);
nor U2990 (N_2990,In_942,In_1029);
or U2991 (N_2991,In_1366,In_1476);
and U2992 (N_2992,In_691,In_975);
and U2993 (N_2993,In_1131,In_1181);
nor U2994 (N_2994,In_651,In_526);
and U2995 (N_2995,In_1459,In_455);
nand U2996 (N_2996,In_306,In_253);
nor U2997 (N_2997,In_754,In_891);
or U2998 (N_2998,In_1269,In_48);
nor U2999 (N_2999,In_368,In_49);
and U3000 (N_3000,In_1340,In_771);
nand U3001 (N_3001,In_500,In_14);
nor U3002 (N_3002,In_1250,In_405);
or U3003 (N_3003,In_311,In_406);
nor U3004 (N_3004,In_544,In_4);
nand U3005 (N_3005,In_897,In_1413);
or U3006 (N_3006,In_1153,In_257);
and U3007 (N_3007,In_472,In_1078);
and U3008 (N_3008,In_1376,In_825);
or U3009 (N_3009,In_1020,In_975);
and U3010 (N_3010,In_1272,In_5);
nand U3011 (N_3011,In_457,In_248);
and U3012 (N_3012,In_760,In_316);
and U3013 (N_3013,In_244,In_396);
or U3014 (N_3014,In_489,In_1419);
nand U3015 (N_3015,In_1426,In_877);
nor U3016 (N_3016,In_1473,In_532);
nand U3017 (N_3017,In_1438,In_1019);
nor U3018 (N_3018,In_1322,In_1377);
nor U3019 (N_3019,In_1192,In_925);
nor U3020 (N_3020,In_647,In_47);
nand U3021 (N_3021,In_716,In_204);
nand U3022 (N_3022,In_1024,In_1301);
and U3023 (N_3023,In_645,In_883);
and U3024 (N_3024,In_1338,In_151);
nand U3025 (N_3025,In_1257,In_1413);
and U3026 (N_3026,In_1180,In_976);
nand U3027 (N_3027,In_141,In_815);
nand U3028 (N_3028,In_993,In_1063);
or U3029 (N_3029,In_802,In_859);
nor U3030 (N_3030,In_592,In_1027);
nor U3031 (N_3031,In_1154,In_308);
nand U3032 (N_3032,In_1003,In_1342);
or U3033 (N_3033,In_903,In_318);
nand U3034 (N_3034,In_1268,In_411);
nor U3035 (N_3035,In_957,In_569);
or U3036 (N_3036,In_1287,In_352);
or U3037 (N_3037,In_651,In_1034);
or U3038 (N_3038,In_654,In_3);
and U3039 (N_3039,In_1288,In_938);
nor U3040 (N_3040,In_912,In_126);
and U3041 (N_3041,In_1301,In_631);
nand U3042 (N_3042,In_655,In_1380);
or U3043 (N_3043,In_842,In_1391);
and U3044 (N_3044,In_1137,In_1043);
or U3045 (N_3045,In_99,In_16);
nand U3046 (N_3046,In_430,In_330);
nand U3047 (N_3047,In_239,In_1072);
or U3048 (N_3048,In_736,In_1250);
or U3049 (N_3049,In_600,In_521);
nand U3050 (N_3050,In_1419,In_1251);
nor U3051 (N_3051,In_1016,In_603);
nor U3052 (N_3052,In_1070,In_223);
and U3053 (N_3053,In_1433,In_710);
nand U3054 (N_3054,In_99,In_1058);
and U3055 (N_3055,In_356,In_1164);
nand U3056 (N_3056,In_323,In_278);
nor U3057 (N_3057,In_491,In_892);
or U3058 (N_3058,In_631,In_1466);
and U3059 (N_3059,In_947,In_158);
nand U3060 (N_3060,In_1348,In_1090);
nor U3061 (N_3061,In_1178,In_1097);
nor U3062 (N_3062,In_595,In_1434);
and U3063 (N_3063,In_770,In_1133);
or U3064 (N_3064,In_263,In_1333);
nor U3065 (N_3065,In_830,In_652);
nor U3066 (N_3066,In_1456,In_1465);
or U3067 (N_3067,In_494,In_342);
or U3068 (N_3068,In_284,In_726);
nand U3069 (N_3069,In_1271,In_536);
and U3070 (N_3070,In_813,In_1293);
or U3071 (N_3071,In_224,In_369);
nor U3072 (N_3072,In_450,In_328);
or U3073 (N_3073,In_907,In_972);
xor U3074 (N_3074,In_112,In_860);
nor U3075 (N_3075,In_274,In_1079);
or U3076 (N_3076,In_728,In_1266);
and U3077 (N_3077,In_899,In_466);
and U3078 (N_3078,In_956,In_434);
nand U3079 (N_3079,In_1252,In_1243);
and U3080 (N_3080,In_84,In_454);
and U3081 (N_3081,In_160,In_373);
nand U3082 (N_3082,In_874,In_197);
nor U3083 (N_3083,In_158,In_1439);
xnor U3084 (N_3084,In_920,In_356);
and U3085 (N_3085,In_627,In_882);
nand U3086 (N_3086,In_532,In_686);
or U3087 (N_3087,In_490,In_295);
nor U3088 (N_3088,In_293,In_689);
nand U3089 (N_3089,In_1341,In_273);
nor U3090 (N_3090,In_455,In_726);
or U3091 (N_3091,In_1324,In_207);
and U3092 (N_3092,In_47,In_357);
nor U3093 (N_3093,In_1284,In_215);
nand U3094 (N_3094,In_153,In_1332);
and U3095 (N_3095,In_974,In_535);
nand U3096 (N_3096,In_914,In_216);
or U3097 (N_3097,In_1006,In_106);
nand U3098 (N_3098,In_1408,In_1216);
nand U3099 (N_3099,In_103,In_886);
and U3100 (N_3100,In_62,In_81);
or U3101 (N_3101,In_1065,In_674);
or U3102 (N_3102,In_346,In_1378);
nand U3103 (N_3103,In_647,In_718);
and U3104 (N_3104,In_792,In_1173);
and U3105 (N_3105,In_1051,In_658);
or U3106 (N_3106,In_1134,In_1420);
nor U3107 (N_3107,In_935,In_525);
and U3108 (N_3108,In_522,In_280);
and U3109 (N_3109,In_1481,In_823);
or U3110 (N_3110,In_633,In_1161);
nand U3111 (N_3111,In_1142,In_448);
or U3112 (N_3112,In_751,In_1014);
nor U3113 (N_3113,In_1165,In_389);
nand U3114 (N_3114,In_825,In_1014);
nor U3115 (N_3115,In_176,In_1156);
nor U3116 (N_3116,In_448,In_1014);
or U3117 (N_3117,In_118,In_1436);
and U3118 (N_3118,In_8,In_480);
and U3119 (N_3119,In_907,In_13);
nor U3120 (N_3120,In_1326,In_765);
nor U3121 (N_3121,In_835,In_864);
and U3122 (N_3122,In_437,In_1232);
nor U3123 (N_3123,In_1407,In_107);
nor U3124 (N_3124,In_1374,In_384);
and U3125 (N_3125,In_343,In_1424);
nand U3126 (N_3126,In_843,In_1202);
nand U3127 (N_3127,In_224,In_1353);
nand U3128 (N_3128,In_924,In_848);
nor U3129 (N_3129,In_897,In_768);
nand U3130 (N_3130,In_927,In_118);
or U3131 (N_3131,In_1444,In_105);
nor U3132 (N_3132,In_869,In_1396);
or U3133 (N_3133,In_617,In_504);
nand U3134 (N_3134,In_450,In_634);
and U3135 (N_3135,In_1170,In_1336);
nor U3136 (N_3136,In_473,In_249);
and U3137 (N_3137,In_222,In_466);
nand U3138 (N_3138,In_1141,In_911);
and U3139 (N_3139,In_1469,In_709);
nand U3140 (N_3140,In_936,In_1240);
and U3141 (N_3141,In_1283,In_1449);
and U3142 (N_3142,In_264,In_999);
and U3143 (N_3143,In_601,In_667);
nand U3144 (N_3144,In_559,In_671);
or U3145 (N_3145,In_331,In_269);
or U3146 (N_3146,In_787,In_1088);
or U3147 (N_3147,In_1072,In_709);
nand U3148 (N_3148,In_1342,In_158);
nor U3149 (N_3149,In_616,In_1456);
and U3150 (N_3150,In_118,In_109);
and U3151 (N_3151,In_760,In_401);
nor U3152 (N_3152,In_808,In_1014);
nor U3153 (N_3153,In_1051,In_803);
or U3154 (N_3154,In_807,In_162);
xnor U3155 (N_3155,In_4,In_621);
nand U3156 (N_3156,In_412,In_146);
or U3157 (N_3157,In_1017,In_823);
or U3158 (N_3158,In_426,In_527);
or U3159 (N_3159,In_1195,In_1007);
or U3160 (N_3160,In_746,In_1339);
and U3161 (N_3161,In_919,In_148);
nor U3162 (N_3162,In_606,In_1027);
and U3163 (N_3163,In_1324,In_828);
and U3164 (N_3164,In_149,In_895);
and U3165 (N_3165,In_276,In_802);
and U3166 (N_3166,In_929,In_826);
nor U3167 (N_3167,In_132,In_824);
nor U3168 (N_3168,In_1156,In_797);
nor U3169 (N_3169,In_854,In_785);
or U3170 (N_3170,In_1136,In_179);
nor U3171 (N_3171,In_804,In_1289);
nand U3172 (N_3172,In_397,In_30);
or U3173 (N_3173,In_830,In_418);
and U3174 (N_3174,In_894,In_48);
and U3175 (N_3175,In_65,In_862);
nand U3176 (N_3176,In_500,In_1328);
and U3177 (N_3177,In_983,In_222);
or U3178 (N_3178,In_1068,In_839);
or U3179 (N_3179,In_1106,In_352);
nor U3180 (N_3180,In_899,In_850);
and U3181 (N_3181,In_387,In_1006);
and U3182 (N_3182,In_1199,In_1210);
nor U3183 (N_3183,In_578,In_429);
nor U3184 (N_3184,In_542,In_344);
nor U3185 (N_3185,In_145,In_1173);
nor U3186 (N_3186,In_732,In_254);
nand U3187 (N_3187,In_1155,In_118);
or U3188 (N_3188,In_782,In_513);
nor U3189 (N_3189,In_124,In_946);
nor U3190 (N_3190,In_852,In_1392);
and U3191 (N_3191,In_216,In_632);
and U3192 (N_3192,In_1363,In_979);
and U3193 (N_3193,In_760,In_411);
or U3194 (N_3194,In_372,In_1475);
nand U3195 (N_3195,In_1354,In_926);
and U3196 (N_3196,In_955,In_649);
nor U3197 (N_3197,In_974,In_495);
and U3198 (N_3198,In_791,In_69);
and U3199 (N_3199,In_698,In_533);
nor U3200 (N_3200,In_938,In_105);
nor U3201 (N_3201,In_716,In_693);
and U3202 (N_3202,In_1339,In_1110);
nand U3203 (N_3203,In_112,In_1205);
or U3204 (N_3204,In_1022,In_919);
nor U3205 (N_3205,In_591,In_515);
nor U3206 (N_3206,In_1421,In_1400);
nand U3207 (N_3207,In_909,In_1258);
and U3208 (N_3208,In_695,In_1392);
or U3209 (N_3209,In_1053,In_1231);
nor U3210 (N_3210,In_1450,In_661);
or U3211 (N_3211,In_1402,In_661);
and U3212 (N_3212,In_1043,In_957);
nand U3213 (N_3213,In_370,In_953);
nand U3214 (N_3214,In_425,In_721);
or U3215 (N_3215,In_1199,In_1415);
or U3216 (N_3216,In_589,In_1412);
or U3217 (N_3217,In_481,In_448);
nand U3218 (N_3218,In_123,In_1123);
nand U3219 (N_3219,In_272,In_1008);
or U3220 (N_3220,In_326,In_1111);
nor U3221 (N_3221,In_1389,In_625);
nor U3222 (N_3222,In_945,In_890);
and U3223 (N_3223,In_1414,In_206);
nor U3224 (N_3224,In_1229,In_61);
or U3225 (N_3225,In_489,In_532);
and U3226 (N_3226,In_1494,In_689);
or U3227 (N_3227,In_1260,In_145);
nand U3228 (N_3228,In_249,In_622);
nor U3229 (N_3229,In_274,In_1281);
nand U3230 (N_3230,In_560,In_239);
or U3231 (N_3231,In_444,In_413);
nand U3232 (N_3232,In_194,In_34);
nor U3233 (N_3233,In_893,In_1050);
nor U3234 (N_3234,In_369,In_39);
or U3235 (N_3235,In_1379,In_131);
or U3236 (N_3236,In_38,In_663);
nor U3237 (N_3237,In_1270,In_214);
and U3238 (N_3238,In_818,In_115);
or U3239 (N_3239,In_838,In_1200);
nand U3240 (N_3240,In_1489,In_804);
and U3241 (N_3241,In_50,In_1051);
and U3242 (N_3242,In_1404,In_818);
and U3243 (N_3243,In_150,In_7);
nand U3244 (N_3244,In_306,In_235);
nand U3245 (N_3245,In_1283,In_115);
and U3246 (N_3246,In_371,In_1412);
nor U3247 (N_3247,In_1127,In_670);
nor U3248 (N_3248,In_990,In_736);
nor U3249 (N_3249,In_583,In_624);
nand U3250 (N_3250,In_736,In_1076);
or U3251 (N_3251,In_917,In_519);
and U3252 (N_3252,In_261,In_404);
and U3253 (N_3253,In_416,In_487);
nand U3254 (N_3254,In_878,In_1047);
nor U3255 (N_3255,In_275,In_1059);
and U3256 (N_3256,In_627,In_1430);
nand U3257 (N_3257,In_1397,In_983);
nor U3258 (N_3258,In_1065,In_1475);
and U3259 (N_3259,In_993,In_1151);
nor U3260 (N_3260,In_533,In_68);
or U3261 (N_3261,In_403,In_118);
nor U3262 (N_3262,In_1234,In_1001);
nand U3263 (N_3263,In_1429,In_480);
or U3264 (N_3264,In_542,In_956);
and U3265 (N_3265,In_428,In_1082);
nor U3266 (N_3266,In_1050,In_66);
nand U3267 (N_3267,In_250,In_1026);
or U3268 (N_3268,In_1309,In_253);
nor U3269 (N_3269,In_819,In_37);
and U3270 (N_3270,In_793,In_1499);
nor U3271 (N_3271,In_977,In_614);
or U3272 (N_3272,In_412,In_338);
nand U3273 (N_3273,In_1171,In_572);
and U3274 (N_3274,In_810,In_1387);
nor U3275 (N_3275,In_829,In_16);
nor U3276 (N_3276,In_1330,In_911);
and U3277 (N_3277,In_967,In_838);
nor U3278 (N_3278,In_1333,In_713);
and U3279 (N_3279,In_327,In_1258);
or U3280 (N_3280,In_591,In_888);
nor U3281 (N_3281,In_474,In_794);
and U3282 (N_3282,In_536,In_703);
nand U3283 (N_3283,In_1450,In_40);
and U3284 (N_3284,In_738,In_1299);
and U3285 (N_3285,In_1244,In_845);
and U3286 (N_3286,In_299,In_823);
and U3287 (N_3287,In_680,In_356);
nand U3288 (N_3288,In_683,In_156);
and U3289 (N_3289,In_205,In_135);
nor U3290 (N_3290,In_1138,In_417);
or U3291 (N_3291,In_1170,In_1217);
nand U3292 (N_3292,In_295,In_429);
and U3293 (N_3293,In_194,In_835);
or U3294 (N_3294,In_503,In_1063);
nor U3295 (N_3295,In_293,In_283);
nor U3296 (N_3296,In_1106,In_638);
or U3297 (N_3297,In_872,In_994);
and U3298 (N_3298,In_318,In_467);
and U3299 (N_3299,In_61,In_844);
nor U3300 (N_3300,In_1447,In_419);
and U3301 (N_3301,In_571,In_587);
and U3302 (N_3302,In_382,In_1253);
nor U3303 (N_3303,In_826,In_222);
nor U3304 (N_3304,In_1371,In_1450);
or U3305 (N_3305,In_1258,In_520);
and U3306 (N_3306,In_437,In_760);
nand U3307 (N_3307,In_288,In_1326);
or U3308 (N_3308,In_892,In_1135);
or U3309 (N_3309,In_572,In_1140);
nor U3310 (N_3310,In_861,In_686);
nor U3311 (N_3311,In_993,In_976);
nor U3312 (N_3312,In_1321,In_1443);
and U3313 (N_3313,In_878,In_886);
nor U3314 (N_3314,In_1344,In_780);
nand U3315 (N_3315,In_542,In_566);
nand U3316 (N_3316,In_1046,In_604);
nand U3317 (N_3317,In_1233,In_570);
or U3318 (N_3318,In_541,In_952);
and U3319 (N_3319,In_624,In_989);
and U3320 (N_3320,In_455,In_152);
nor U3321 (N_3321,In_657,In_873);
and U3322 (N_3322,In_689,In_1013);
and U3323 (N_3323,In_762,In_114);
and U3324 (N_3324,In_182,In_543);
and U3325 (N_3325,In_1045,In_936);
nand U3326 (N_3326,In_706,In_532);
nand U3327 (N_3327,In_99,In_1087);
or U3328 (N_3328,In_889,In_565);
and U3329 (N_3329,In_966,In_789);
and U3330 (N_3330,In_1149,In_43);
and U3331 (N_3331,In_1006,In_201);
nor U3332 (N_3332,In_655,In_913);
and U3333 (N_3333,In_300,In_1128);
nor U3334 (N_3334,In_90,In_1136);
nor U3335 (N_3335,In_995,In_1122);
or U3336 (N_3336,In_667,In_826);
nor U3337 (N_3337,In_457,In_1007);
and U3338 (N_3338,In_932,In_1234);
or U3339 (N_3339,In_1187,In_1139);
nand U3340 (N_3340,In_1028,In_7);
nor U3341 (N_3341,In_1308,In_1051);
nand U3342 (N_3342,In_1162,In_817);
or U3343 (N_3343,In_84,In_1218);
nand U3344 (N_3344,In_714,In_112);
nor U3345 (N_3345,In_1183,In_814);
nand U3346 (N_3346,In_1093,In_1002);
or U3347 (N_3347,In_665,In_153);
and U3348 (N_3348,In_1273,In_289);
nor U3349 (N_3349,In_858,In_180);
or U3350 (N_3350,In_702,In_216);
and U3351 (N_3351,In_212,In_1406);
nor U3352 (N_3352,In_610,In_1230);
or U3353 (N_3353,In_1435,In_764);
nor U3354 (N_3354,In_347,In_1452);
nand U3355 (N_3355,In_1408,In_109);
and U3356 (N_3356,In_804,In_734);
or U3357 (N_3357,In_229,In_1048);
nand U3358 (N_3358,In_1377,In_976);
nor U3359 (N_3359,In_1208,In_764);
and U3360 (N_3360,In_782,In_66);
nand U3361 (N_3361,In_106,In_772);
nor U3362 (N_3362,In_1476,In_1315);
nor U3363 (N_3363,In_419,In_78);
nor U3364 (N_3364,In_273,In_439);
and U3365 (N_3365,In_1192,In_1021);
or U3366 (N_3366,In_1244,In_166);
nor U3367 (N_3367,In_1047,In_767);
nor U3368 (N_3368,In_80,In_1093);
and U3369 (N_3369,In_155,In_1421);
nor U3370 (N_3370,In_1249,In_141);
and U3371 (N_3371,In_1259,In_50);
and U3372 (N_3372,In_133,In_712);
and U3373 (N_3373,In_847,In_423);
or U3374 (N_3374,In_1017,In_1172);
and U3375 (N_3375,In_222,In_1420);
and U3376 (N_3376,In_1128,In_411);
nor U3377 (N_3377,In_976,In_1077);
nand U3378 (N_3378,In_415,In_1383);
nor U3379 (N_3379,In_767,In_661);
nor U3380 (N_3380,In_851,In_1231);
and U3381 (N_3381,In_1074,In_879);
nor U3382 (N_3382,In_122,In_388);
nor U3383 (N_3383,In_117,In_1118);
or U3384 (N_3384,In_136,In_1223);
and U3385 (N_3385,In_877,In_911);
or U3386 (N_3386,In_496,In_1207);
or U3387 (N_3387,In_923,In_825);
nor U3388 (N_3388,In_530,In_227);
and U3389 (N_3389,In_1007,In_1278);
or U3390 (N_3390,In_147,In_686);
nand U3391 (N_3391,In_712,In_319);
nor U3392 (N_3392,In_1092,In_489);
and U3393 (N_3393,In_582,In_1453);
nor U3394 (N_3394,In_170,In_1032);
nand U3395 (N_3395,In_848,In_995);
and U3396 (N_3396,In_970,In_175);
or U3397 (N_3397,In_548,In_1131);
or U3398 (N_3398,In_1053,In_830);
or U3399 (N_3399,In_711,In_836);
and U3400 (N_3400,In_1187,In_105);
or U3401 (N_3401,In_167,In_679);
and U3402 (N_3402,In_770,In_1058);
and U3403 (N_3403,In_400,In_524);
and U3404 (N_3404,In_1198,In_1461);
and U3405 (N_3405,In_574,In_131);
nand U3406 (N_3406,In_1052,In_1494);
nand U3407 (N_3407,In_1145,In_1077);
nand U3408 (N_3408,In_954,In_1078);
nor U3409 (N_3409,In_1075,In_907);
or U3410 (N_3410,In_436,In_1385);
and U3411 (N_3411,In_1388,In_785);
nand U3412 (N_3412,In_524,In_559);
nor U3413 (N_3413,In_762,In_1376);
nor U3414 (N_3414,In_678,In_249);
and U3415 (N_3415,In_858,In_853);
and U3416 (N_3416,In_609,In_778);
nand U3417 (N_3417,In_819,In_247);
nand U3418 (N_3418,In_1187,In_1249);
and U3419 (N_3419,In_702,In_883);
and U3420 (N_3420,In_1426,In_309);
and U3421 (N_3421,In_142,In_638);
nor U3422 (N_3422,In_310,In_748);
and U3423 (N_3423,In_1151,In_440);
and U3424 (N_3424,In_1444,In_1033);
or U3425 (N_3425,In_852,In_1002);
nor U3426 (N_3426,In_1498,In_366);
and U3427 (N_3427,In_834,In_501);
or U3428 (N_3428,In_133,In_1414);
nor U3429 (N_3429,In_1256,In_1346);
nor U3430 (N_3430,In_1309,In_905);
xor U3431 (N_3431,In_1391,In_1017);
or U3432 (N_3432,In_26,In_153);
or U3433 (N_3433,In_258,In_1375);
or U3434 (N_3434,In_1325,In_638);
or U3435 (N_3435,In_710,In_953);
or U3436 (N_3436,In_1466,In_1324);
nand U3437 (N_3437,In_700,In_1114);
nand U3438 (N_3438,In_687,In_441);
and U3439 (N_3439,In_1027,In_1400);
nand U3440 (N_3440,In_1310,In_109);
and U3441 (N_3441,In_1409,In_37);
and U3442 (N_3442,In_578,In_1349);
nor U3443 (N_3443,In_804,In_140);
or U3444 (N_3444,In_34,In_735);
nand U3445 (N_3445,In_515,In_1461);
nor U3446 (N_3446,In_1336,In_1054);
or U3447 (N_3447,In_637,In_173);
nand U3448 (N_3448,In_516,In_1491);
or U3449 (N_3449,In_244,In_939);
nor U3450 (N_3450,In_316,In_1065);
or U3451 (N_3451,In_347,In_282);
nor U3452 (N_3452,In_912,In_1362);
or U3453 (N_3453,In_1100,In_132);
and U3454 (N_3454,In_65,In_1467);
or U3455 (N_3455,In_139,In_31);
or U3456 (N_3456,In_1124,In_926);
nand U3457 (N_3457,In_1247,In_844);
or U3458 (N_3458,In_1158,In_1411);
or U3459 (N_3459,In_306,In_66);
or U3460 (N_3460,In_1211,In_760);
xnor U3461 (N_3461,In_930,In_1006);
nand U3462 (N_3462,In_273,In_96);
and U3463 (N_3463,In_41,In_152);
nor U3464 (N_3464,In_1057,In_390);
nand U3465 (N_3465,In_386,In_1144);
or U3466 (N_3466,In_333,In_1073);
and U3467 (N_3467,In_451,In_1173);
or U3468 (N_3468,In_855,In_1428);
nor U3469 (N_3469,In_274,In_1295);
nor U3470 (N_3470,In_908,In_1050);
or U3471 (N_3471,In_869,In_1171);
or U3472 (N_3472,In_175,In_1436);
nand U3473 (N_3473,In_1152,In_169);
and U3474 (N_3474,In_801,In_110);
nand U3475 (N_3475,In_1118,In_229);
nor U3476 (N_3476,In_1167,In_1366);
and U3477 (N_3477,In_317,In_87);
and U3478 (N_3478,In_114,In_731);
and U3479 (N_3479,In_1267,In_1402);
nor U3480 (N_3480,In_1443,In_574);
and U3481 (N_3481,In_343,In_468);
or U3482 (N_3482,In_1019,In_919);
and U3483 (N_3483,In_27,In_517);
nand U3484 (N_3484,In_590,In_779);
nor U3485 (N_3485,In_873,In_1439);
nor U3486 (N_3486,In_472,In_1317);
or U3487 (N_3487,In_243,In_476);
xnor U3488 (N_3488,In_406,In_1345);
or U3489 (N_3489,In_332,In_650);
nor U3490 (N_3490,In_1198,In_431);
and U3491 (N_3491,In_958,In_247);
nand U3492 (N_3492,In_892,In_563);
nand U3493 (N_3493,In_1396,In_1066);
and U3494 (N_3494,In_1108,In_1357);
nor U3495 (N_3495,In_1331,In_1124);
and U3496 (N_3496,In_1207,In_209);
nand U3497 (N_3497,In_68,In_991);
nor U3498 (N_3498,In_182,In_144);
nor U3499 (N_3499,In_68,In_824);
nand U3500 (N_3500,In_18,In_308);
nor U3501 (N_3501,In_978,In_1426);
and U3502 (N_3502,In_603,In_802);
nor U3503 (N_3503,In_874,In_1279);
nor U3504 (N_3504,In_930,In_1034);
nand U3505 (N_3505,In_414,In_671);
and U3506 (N_3506,In_1159,In_1016);
nor U3507 (N_3507,In_1354,In_1178);
or U3508 (N_3508,In_550,In_290);
and U3509 (N_3509,In_241,In_696);
nand U3510 (N_3510,In_651,In_770);
or U3511 (N_3511,In_62,In_13);
or U3512 (N_3512,In_473,In_891);
nor U3513 (N_3513,In_368,In_705);
and U3514 (N_3514,In_626,In_1348);
and U3515 (N_3515,In_963,In_306);
xor U3516 (N_3516,In_270,In_1320);
nor U3517 (N_3517,In_854,In_1109);
or U3518 (N_3518,In_1306,In_878);
nand U3519 (N_3519,In_1423,In_964);
nand U3520 (N_3520,In_422,In_753);
or U3521 (N_3521,In_958,In_1296);
nand U3522 (N_3522,In_1197,In_990);
or U3523 (N_3523,In_351,In_4);
or U3524 (N_3524,In_866,In_428);
or U3525 (N_3525,In_744,In_1143);
nand U3526 (N_3526,In_737,In_760);
or U3527 (N_3527,In_947,In_1321);
nand U3528 (N_3528,In_87,In_658);
or U3529 (N_3529,In_324,In_841);
nand U3530 (N_3530,In_23,In_1370);
nor U3531 (N_3531,In_584,In_705);
and U3532 (N_3532,In_643,In_454);
nand U3533 (N_3533,In_20,In_647);
or U3534 (N_3534,In_1029,In_837);
nor U3535 (N_3535,In_1227,In_509);
and U3536 (N_3536,In_667,In_1165);
nor U3537 (N_3537,In_1344,In_120);
and U3538 (N_3538,In_248,In_181);
nor U3539 (N_3539,In_395,In_366);
and U3540 (N_3540,In_1400,In_161);
and U3541 (N_3541,In_663,In_1303);
nor U3542 (N_3542,In_1371,In_1082);
and U3543 (N_3543,In_594,In_447);
nand U3544 (N_3544,In_564,In_1391);
or U3545 (N_3545,In_1232,In_560);
nand U3546 (N_3546,In_1017,In_383);
nand U3547 (N_3547,In_969,In_848);
nor U3548 (N_3548,In_205,In_1119);
nor U3549 (N_3549,In_853,In_1102);
nand U3550 (N_3550,In_1012,In_166);
nand U3551 (N_3551,In_264,In_67);
nand U3552 (N_3552,In_623,In_362);
and U3553 (N_3553,In_11,In_679);
nor U3554 (N_3554,In_1011,In_1470);
and U3555 (N_3555,In_453,In_378);
or U3556 (N_3556,In_375,In_402);
xnor U3557 (N_3557,In_35,In_396);
nand U3558 (N_3558,In_1145,In_1174);
nand U3559 (N_3559,In_1418,In_1235);
nand U3560 (N_3560,In_461,In_89);
or U3561 (N_3561,In_805,In_1341);
or U3562 (N_3562,In_1389,In_1489);
nand U3563 (N_3563,In_1017,In_662);
and U3564 (N_3564,In_87,In_1040);
and U3565 (N_3565,In_213,In_518);
nand U3566 (N_3566,In_1121,In_1030);
nand U3567 (N_3567,In_1148,In_96);
nand U3568 (N_3568,In_1085,In_1129);
or U3569 (N_3569,In_1384,In_207);
xnor U3570 (N_3570,In_682,In_88);
or U3571 (N_3571,In_1455,In_1109);
and U3572 (N_3572,In_307,In_792);
nand U3573 (N_3573,In_107,In_1499);
and U3574 (N_3574,In_805,In_1064);
and U3575 (N_3575,In_285,In_290);
nand U3576 (N_3576,In_978,In_1416);
nor U3577 (N_3577,In_1221,In_1191);
nand U3578 (N_3578,In_313,In_14);
or U3579 (N_3579,In_335,In_201);
or U3580 (N_3580,In_329,In_1300);
nor U3581 (N_3581,In_233,In_511);
nand U3582 (N_3582,In_57,In_820);
nor U3583 (N_3583,In_212,In_846);
and U3584 (N_3584,In_361,In_1427);
or U3585 (N_3585,In_489,In_1296);
nor U3586 (N_3586,In_302,In_1447);
and U3587 (N_3587,In_383,In_1263);
nor U3588 (N_3588,In_904,In_625);
nand U3589 (N_3589,In_435,In_923);
and U3590 (N_3590,In_1090,In_1157);
nor U3591 (N_3591,In_198,In_233);
nor U3592 (N_3592,In_84,In_1030);
and U3593 (N_3593,In_480,In_840);
or U3594 (N_3594,In_1478,In_1226);
nand U3595 (N_3595,In_913,In_152);
nor U3596 (N_3596,In_1214,In_70);
nand U3597 (N_3597,In_1350,In_79);
and U3598 (N_3598,In_1133,In_1273);
or U3599 (N_3599,In_1021,In_839);
or U3600 (N_3600,In_682,In_32);
or U3601 (N_3601,In_750,In_900);
nor U3602 (N_3602,In_130,In_28);
or U3603 (N_3603,In_600,In_794);
and U3604 (N_3604,In_778,In_502);
and U3605 (N_3605,In_684,In_138);
or U3606 (N_3606,In_412,In_534);
nor U3607 (N_3607,In_788,In_415);
and U3608 (N_3608,In_1388,In_423);
nand U3609 (N_3609,In_630,In_710);
nor U3610 (N_3610,In_741,In_1036);
nand U3611 (N_3611,In_65,In_1398);
nand U3612 (N_3612,In_1286,In_1009);
and U3613 (N_3613,In_1286,In_1195);
nand U3614 (N_3614,In_541,In_1026);
nor U3615 (N_3615,In_1223,In_95);
or U3616 (N_3616,In_239,In_951);
nor U3617 (N_3617,In_652,In_178);
nor U3618 (N_3618,In_805,In_300);
nor U3619 (N_3619,In_1258,In_1240);
nor U3620 (N_3620,In_307,In_1468);
xor U3621 (N_3621,In_961,In_982);
and U3622 (N_3622,In_1257,In_211);
xor U3623 (N_3623,In_398,In_237);
or U3624 (N_3624,In_1468,In_1244);
nor U3625 (N_3625,In_276,In_963);
nor U3626 (N_3626,In_966,In_387);
or U3627 (N_3627,In_866,In_275);
and U3628 (N_3628,In_1423,In_1334);
nor U3629 (N_3629,In_1031,In_106);
and U3630 (N_3630,In_394,In_848);
nor U3631 (N_3631,In_889,In_1460);
nor U3632 (N_3632,In_1230,In_322);
nand U3633 (N_3633,In_690,In_118);
xnor U3634 (N_3634,In_614,In_1091);
nor U3635 (N_3635,In_962,In_837);
and U3636 (N_3636,In_944,In_1492);
nor U3637 (N_3637,In_1072,In_651);
or U3638 (N_3638,In_248,In_237);
nor U3639 (N_3639,In_47,In_718);
or U3640 (N_3640,In_928,In_1062);
nand U3641 (N_3641,In_217,In_828);
or U3642 (N_3642,In_1119,In_848);
nand U3643 (N_3643,In_945,In_1402);
nor U3644 (N_3644,In_1351,In_621);
nor U3645 (N_3645,In_1349,In_223);
nand U3646 (N_3646,In_495,In_280);
and U3647 (N_3647,In_150,In_614);
nor U3648 (N_3648,In_867,In_766);
nand U3649 (N_3649,In_601,In_196);
or U3650 (N_3650,In_1020,In_746);
nand U3651 (N_3651,In_996,In_463);
or U3652 (N_3652,In_1195,In_910);
nor U3653 (N_3653,In_1215,In_997);
nand U3654 (N_3654,In_95,In_685);
or U3655 (N_3655,In_1485,In_1279);
and U3656 (N_3656,In_624,In_1418);
nand U3657 (N_3657,In_1078,In_1283);
and U3658 (N_3658,In_677,In_713);
nor U3659 (N_3659,In_87,In_98);
nor U3660 (N_3660,In_1064,In_1131);
or U3661 (N_3661,In_210,In_225);
nor U3662 (N_3662,In_709,In_571);
nand U3663 (N_3663,In_1140,In_707);
nor U3664 (N_3664,In_1068,In_510);
nor U3665 (N_3665,In_237,In_377);
nor U3666 (N_3666,In_567,In_849);
nor U3667 (N_3667,In_984,In_234);
and U3668 (N_3668,In_726,In_818);
or U3669 (N_3669,In_315,In_1389);
or U3670 (N_3670,In_344,In_252);
nand U3671 (N_3671,In_1059,In_1442);
or U3672 (N_3672,In_671,In_929);
nand U3673 (N_3673,In_184,In_1450);
nand U3674 (N_3674,In_607,In_1062);
nand U3675 (N_3675,In_1258,In_1232);
nor U3676 (N_3676,In_1168,In_1238);
nor U3677 (N_3677,In_297,In_790);
nor U3678 (N_3678,In_1258,In_1224);
and U3679 (N_3679,In_322,In_730);
and U3680 (N_3680,In_385,In_987);
nor U3681 (N_3681,In_765,In_1461);
and U3682 (N_3682,In_669,In_826);
nor U3683 (N_3683,In_21,In_1047);
or U3684 (N_3684,In_1003,In_244);
or U3685 (N_3685,In_78,In_228);
nor U3686 (N_3686,In_1178,In_528);
or U3687 (N_3687,In_1413,In_972);
nand U3688 (N_3688,In_408,In_1465);
nand U3689 (N_3689,In_1101,In_1461);
and U3690 (N_3690,In_963,In_911);
nand U3691 (N_3691,In_1331,In_650);
nand U3692 (N_3692,In_85,In_761);
or U3693 (N_3693,In_273,In_188);
and U3694 (N_3694,In_528,In_474);
or U3695 (N_3695,In_1430,In_922);
and U3696 (N_3696,In_264,In_525);
nor U3697 (N_3697,In_1320,In_325);
nand U3698 (N_3698,In_1185,In_938);
and U3699 (N_3699,In_13,In_1213);
and U3700 (N_3700,In_663,In_1453);
or U3701 (N_3701,In_1115,In_931);
nand U3702 (N_3702,In_684,In_562);
and U3703 (N_3703,In_51,In_414);
or U3704 (N_3704,In_116,In_328);
or U3705 (N_3705,In_1417,In_537);
nand U3706 (N_3706,In_1047,In_897);
or U3707 (N_3707,In_1115,In_111);
or U3708 (N_3708,In_528,In_420);
or U3709 (N_3709,In_455,In_1175);
nor U3710 (N_3710,In_756,In_141);
xor U3711 (N_3711,In_1434,In_296);
or U3712 (N_3712,In_397,In_787);
or U3713 (N_3713,In_1083,In_1164);
nor U3714 (N_3714,In_258,In_992);
or U3715 (N_3715,In_1452,In_1120);
and U3716 (N_3716,In_913,In_526);
nor U3717 (N_3717,In_1142,In_341);
and U3718 (N_3718,In_516,In_633);
nand U3719 (N_3719,In_684,In_25);
nand U3720 (N_3720,In_948,In_248);
nand U3721 (N_3721,In_1414,In_1145);
nand U3722 (N_3722,In_92,In_4);
nor U3723 (N_3723,In_1327,In_843);
nor U3724 (N_3724,In_1450,In_352);
nor U3725 (N_3725,In_537,In_693);
nor U3726 (N_3726,In_1470,In_1225);
nand U3727 (N_3727,In_811,In_782);
or U3728 (N_3728,In_875,In_503);
and U3729 (N_3729,In_87,In_324);
or U3730 (N_3730,In_1218,In_868);
and U3731 (N_3731,In_249,In_1326);
and U3732 (N_3732,In_712,In_25);
and U3733 (N_3733,In_815,In_741);
nor U3734 (N_3734,In_265,In_671);
nand U3735 (N_3735,In_353,In_817);
nor U3736 (N_3736,In_1029,In_515);
or U3737 (N_3737,In_127,In_342);
nand U3738 (N_3738,In_449,In_285);
nor U3739 (N_3739,In_1418,In_1240);
and U3740 (N_3740,In_192,In_790);
nor U3741 (N_3741,In_392,In_1320);
or U3742 (N_3742,In_431,In_1215);
and U3743 (N_3743,In_931,In_693);
or U3744 (N_3744,In_708,In_733);
nand U3745 (N_3745,In_408,In_975);
or U3746 (N_3746,In_1480,In_526);
or U3747 (N_3747,In_1366,In_844);
nand U3748 (N_3748,In_806,In_656);
nand U3749 (N_3749,In_942,In_1344);
nor U3750 (N_3750,In_175,In_1088);
nor U3751 (N_3751,In_14,In_1394);
nand U3752 (N_3752,In_1384,In_274);
nand U3753 (N_3753,In_1263,In_1357);
nor U3754 (N_3754,In_1000,In_926);
or U3755 (N_3755,In_1396,In_1174);
and U3756 (N_3756,In_495,In_602);
nand U3757 (N_3757,In_812,In_806);
nor U3758 (N_3758,In_1080,In_1141);
or U3759 (N_3759,In_138,In_1159);
or U3760 (N_3760,In_279,In_866);
or U3761 (N_3761,In_290,In_124);
nand U3762 (N_3762,In_855,In_410);
nor U3763 (N_3763,In_679,In_1094);
xor U3764 (N_3764,In_316,In_1267);
nor U3765 (N_3765,In_544,In_403);
or U3766 (N_3766,In_572,In_181);
or U3767 (N_3767,In_223,In_229);
and U3768 (N_3768,In_1298,In_1238);
nor U3769 (N_3769,In_1377,In_978);
or U3770 (N_3770,In_703,In_50);
and U3771 (N_3771,In_61,In_285);
and U3772 (N_3772,In_349,In_228);
and U3773 (N_3773,In_112,In_1264);
nor U3774 (N_3774,In_888,In_394);
or U3775 (N_3775,In_67,In_718);
xor U3776 (N_3776,In_1055,In_1460);
or U3777 (N_3777,In_727,In_570);
or U3778 (N_3778,In_1475,In_497);
and U3779 (N_3779,In_373,In_68);
nand U3780 (N_3780,In_1254,In_595);
nor U3781 (N_3781,In_664,In_227);
nor U3782 (N_3782,In_496,In_1338);
or U3783 (N_3783,In_1283,In_623);
or U3784 (N_3784,In_1495,In_1239);
and U3785 (N_3785,In_1139,In_984);
nor U3786 (N_3786,In_27,In_1260);
xor U3787 (N_3787,In_857,In_911);
and U3788 (N_3788,In_1087,In_1316);
nand U3789 (N_3789,In_708,In_328);
and U3790 (N_3790,In_735,In_327);
or U3791 (N_3791,In_53,In_1341);
xnor U3792 (N_3792,In_1295,In_595);
nor U3793 (N_3793,In_529,In_728);
nand U3794 (N_3794,In_1384,In_828);
or U3795 (N_3795,In_398,In_684);
or U3796 (N_3796,In_1155,In_659);
and U3797 (N_3797,In_471,In_1214);
and U3798 (N_3798,In_545,In_1180);
nor U3799 (N_3799,In_607,In_1199);
nor U3800 (N_3800,In_547,In_563);
or U3801 (N_3801,In_943,In_776);
nand U3802 (N_3802,In_157,In_495);
nand U3803 (N_3803,In_137,In_129);
or U3804 (N_3804,In_1436,In_1083);
nor U3805 (N_3805,In_779,In_767);
or U3806 (N_3806,In_1004,In_1190);
nor U3807 (N_3807,In_243,In_56);
and U3808 (N_3808,In_1295,In_679);
nor U3809 (N_3809,In_936,In_1025);
nor U3810 (N_3810,In_127,In_24);
nand U3811 (N_3811,In_638,In_361);
nor U3812 (N_3812,In_1164,In_1039);
and U3813 (N_3813,In_426,In_1085);
or U3814 (N_3814,In_1208,In_690);
nand U3815 (N_3815,In_1397,In_1181);
or U3816 (N_3816,In_1042,In_1165);
xor U3817 (N_3817,In_499,In_1260);
nor U3818 (N_3818,In_326,In_1465);
nand U3819 (N_3819,In_417,In_949);
or U3820 (N_3820,In_221,In_997);
and U3821 (N_3821,In_217,In_35);
nand U3822 (N_3822,In_556,In_560);
nor U3823 (N_3823,In_777,In_1370);
or U3824 (N_3824,In_1263,In_639);
nor U3825 (N_3825,In_1006,In_131);
and U3826 (N_3826,In_487,In_1262);
and U3827 (N_3827,In_198,In_1105);
xnor U3828 (N_3828,In_757,In_1008);
nand U3829 (N_3829,In_1423,In_621);
or U3830 (N_3830,In_1320,In_781);
and U3831 (N_3831,In_395,In_582);
nand U3832 (N_3832,In_21,In_352);
nor U3833 (N_3833,In_812,In_1202);
and U3834 (N_3834,In_855,In_452);
nand U3835 (N_3835,In_1167,In_1047);
nor U3836 (N_3836,In_903,In_403);
or U3837 (N_3837,In_939,In_247);
nand U3838 (N_3838,In_578,In_387);
or U3839 (N_3839,In_41,In_1030);
and U3840 (N_3840,In_440,In_1487);
xor U3841 (N_3841,In_535,In_117);
and U3842 (N_3842,In_1190,In_850);
nor U3843 (N_3843,In_1470,In_761);
and U3844 (N_3844,In_1289,In_1435);
nand U3845 (N_3845,In_910,In_753);
and U3846 (N_3846,In_2,In_291);
nor U3847 (N_3847,In_325,In_628);
and U3848 (N_3848,In_747,In_856);
and U3849 (N_3849,In_721,In_712);
nand U3850 (N_3850,In_452,In_211);
nor U3851 (N_3851,In_909,In_831);
and U3852 (N_3852,In_1307,In_86);
and U3853 (N_3853,In_1426,In_1061);
or U3854 (N_3854,In_176,In_277);
nand U3855 (N_3855,In_1052,In_1380);
nor U3856 (N_3856,In_253,In_455);
nand U3857 (N_3857,In_1261,In_143);
or U3858 (N_3858,In_472,In_367);
nand U3859 (N_3859,In_1057,In_156);
and U3860 (N_3860,In_1178,In_184);
nor U3861 (N_3861,In_333,In_306);
nor U3862 (N_3862,In_103,In_163);
nand U3863 (N_3863,In_43,In_530);
nand U3864 (N_3864,In_1417,In_957);
and U3865 (N_3865,In_524,In_573);
nand U3866 (N_3866,In_647,In_750);
or U3867 (N_3867,In_159,In_116);
or U3868 (N_3868,In_1018,In_1376);
nor U3869 (N_3869,In_719,In_290);
nor U3870 (N_3870,In_665,In_147);
or U3871 (N_3871,In_322,In_71);
nand U3872 (N_3872,In_323,In_10);
nor U3873 (N_3873,In_309,In_1408);
and U3874 (N_3874,In_831,In_1049);
nor U3875 (N_3875,In_639,In_635);
or U3876 (N_3876,In_464,In_514);
and U3877 (N_3877,In_34,In_1172);
and U3878 (N_3878,In_30,In_1278);
or U3879 (N_3879,In_1026,In_226);
nor U3880 (N_3880,In_916,In_333);
and U3881 (N_3881,In_349,In_1478);
nor U3882 (N_3882,In_1113,In_231);
or U3883 (N_3883,In_1489,In_1190);
nor U3884 (N_3884,In_69,In_731);
and U3885 (N_3885,In_1440,In_329);
or U3886 (N_3886,In_689,In_175);
and U3887 (N_3887,In_432,In_988);
nor U3888 (N_3888,In_199,In_549);
and U3889 (N_3889,In_1236,In_1138);
nand U3890 (N_3890,In_221,In_1007);
or U3891 (N_3891,In_294,In_1272);
and U3892 (N_3892,In_809,In_1027);
nor U3893 (N_3893,In_52,In_600);
nand U3894 (N_3894,In_1012,In_491);
or U3895 (N_3895,In_584,In_197);
nand U3896 (N_3896,In_800,In_233);
nor U3897 (N_3897,In_849,In_614);
and U3898 (N_3898,In_519,In_777);
or U3899 (N_3899,In_521,In_1476);
nand U3900 (N_3900,In_555,In_908);
nand U3901 (N_3901,In_287,In_96);
and U3902 (N_3902,In_87,In_578);
or U3903 (N_3903,In_1119,In_191);
nor U3904 (N_3904,In_944,In_553);
nand U3905 (N_3905,In_1347,In_1115);
or U3906 (N_3906,In_1200,In_1052);
or U3907 (N_3907,In_231,In_678);
nand U3908 (N_3908,In_275,In_1106);
or U3909 (N_3909,In_1164,In_360);
and U3910 (N_3910,In_1012,In_526);
nor U3911 (N_3911,In_1241,In_921);
nor U3912 (N_3912,In_1377,In_1293);
or U3913 (N_3913,In_1224,In_349);
or U3914 (N_3914,In_371,In_402);
or U3915 (N_3915,In_1346,In_674);
nand U3916 (N_3916,In_526,In_1120);
or U3917 (N_3917,In_1121,In_218);
nor U3918 (N_3918,In_1104,In_480);
or U3919 (N_3919,In_66,In_1053);
and U3920 (N_3920,In_939,In_454);
or U3921 (N_3921,In_1232,In_1349);
nand U3922 (N_3922,In_797,In_1390);
nand U3923 (N_3923,In_635,In_417);
nand U3924 (N_3924,In_820,In_1283);
nand U3925 (N_3925,In_1465,In_1492);
and U3926 (N_3926,In_911,In_1249);
nand U3927 (N_3927,In_155,In_1180);
and U3928 (N_3928,In_348,In_1342);
or U3929 (N_3929,In_1356,In_1404);
nand U3930 (N_3930,In_220,In_223);
or U3931 (N_3931,In_199,In_515);
or U3932 (N_3932,In_1296,In_803);
nor U3933 (N_3933,In_1338,In_858);
or U3934 (N_3934,In_538,In_838);
or U3935 (N_3935,In_172,In_1218);
nor U3936 (N_3936,In_273,In_1082);
or U3937 (N_3937,In_805,In_871);
or U3938 (N_3938,In_1404,In_1044);
and U3939 (N_3939,In_749,In_655);
nand U3940 (N_3940,In_745,In_1388);
and U3941 (N_3941,In_657,In_483);
or U3942 (N_3942,In_970,In_1423);
nor U3943 (N_3943,In_1320,In_683);
or U3944 (N_3944,In_1407,In_1055);
and U3945 (N_3945,In_257,In_968);
or U3946 (N_3946,In_1290,In_842);
or U3947 (N_3947,In_248,In_902);
nor U3948 (N_3948,In_251,In_1268);
nand U3949 (N_3949,In_1326,In_943);
or U3950 (N_3950,In_784,In_1443);
nor U3951 (N_3951,In_329,In_430);
and U3952 (N_3952,In_1124,In_1445);
and U3953 (N_3953,In_602,In_629);
nand U3954 (N_3954,In_634,In_855);
or U3955 (N_3955,In_1320,In_268);
xor U3956 (N_3956,In_697,In_834);
nor U3957 (N_3957,In_584,In_506);
nand U3958 (N_3958,In_1381,In_1305);
nand U3959 (N_3959,In_1036,In_61);
nand U3960 (N_3960,In_1426,In_64);
and U3961 (N_3961,In_987,In_1387);
nor U3962 (N_3962,In_1300,In_1422);
nand U3963 (N_3963,In_1176,In_334);
nand U3964 (N_3964,In_1291,In_359);
or U3965 (N_3965,In_465,In_1334);
or U3966 (N_3966,In_402,In_856);
or U3967 (N_3967,In_1041,In_51);
or U3968 (N_3968,In_397,In_317);
nand U3969 (N_3969,In_549,In_1185);
nand U3970 (N_3970,In_1002,In_1041);
and U3971 (N_3971,In_1289,In_831);
and U3972 (N_3972,In_510,In_496);
nor U3973 (N_3973,In_1314,In_98);
or U3974 (N_3974,In_542,In_1241);
nand U3975 (N_3975,In_778,In_459);
or U3976 (N_3976,In_286,In_783);
nand U3977 (N_3977,In_763,In_313);
or U3978 (N_3978,In_839,In_52);
nand U3979 (N_3979,In_43,In_1295);
or U3980 (N_3980,In_445,In_657);
nor U3981 (N_3981,In_697,In_630);
or U3982 (N_3982,In_568,In_1078);
or U3983 (N_3983,In_1346,In_1307);
nand U3984 (N_3984,In_51,In_358);
and U3985 (N_3985,In_974,In_322);
and U3986 (N_3986,In_804,In_1275);
and U3987 (N_3987,In_1485,In_1012);
nor U3988 (N_3988,In_801,In_1187);
nand U3989 (N_3989,In_1413,In_40);
nor U3990 (N_3990,In_863,In_27);
and U3991 (N_3991,In_315,In_1479);
xnor U3992 (N_3992,In_1331,In_76);
nand U3993 (N_3993,In_892,In_223);
nand U3994 (N_3994,In_1337,In_1280);
nor U3995 (N_3995,In_1498,In_376);
or U3996 (N_3996,In_880,In_1263);
or U3997 (N_3997,In_1045,In_1166);
nor U3998 (N_3998,In_352,In_61);
nor U3999 (N_3999,In_22,In_344);
nand U4000 (N_4000,In_433,In_1100);
and U4001 (N_4001,In_454,In_1487);
nor U4002 (N_4002,In_1182,In_1318);
or U4003 (N_4003,In_1439,In_1205);
and U4004 (N_4004,In_195,In_1428);
or U4005 (N_4005,In_1078,In_179);
and U4006 (N_4006,In_919,In_1071);
nand U4007 (N_4007,In_607,In_751);
nand U4008 (N_4008,In_1188,In_309);
and U4009 (N_4009,In_466,In_1171);
and U4010 (N_4010,In_652,In_1321);
or U4011 (N_4011,In_1323,In_868);
nand U4012 (N_4012,In_884,In_166);
and U4013 (N_4013,In_1133,In_467);
nor U4014 (N_4014,In_991,In_643);
or U4015 (N_4015,In_445,In_626);
and U4016 (N_4016,In_200,In_135);
nor U4017 (N_4017,In_204,In_242);
nor U4018 (N_4018,In_249,In_1498);
and U4019 (N_4019,In_1494,In_598);
nand U4020 (N_4020,In_319,In_927);
and U4021 (N_4021,In_1116,In_939);
nor U4022 (N_4022,In_1213,In_220);
nor U4023 (N_4023,In_809,In_832);
nor U4024 (N_4024,In_1222,In_849);
nand U4025 (N_4025,In_937,In_828);
nand U4026 (N_4026,In_133,In_188);
nand U4027 (N_4027,In_74,In_1449);
and U4028 (N_4028,In_1345,In_757);
nor U4029 (N_4029,In_62,In_321);
and U4030 (N_4030,In_1437,In_612);
or U4031 (N_4031,In_162,In_779);
and U4032 (N_4032,In_478,In_163);
or U4033 (N_4033,In_1405,In_931);
and U4034 (N_4034,In_401,In_179);
and U4035 (N_4035,In_658,In_250);
nand U4036 (N_4036,In_442,In_1252);
and U4037 (N_4037,In_1297,In_1348);
and U4038 (N_4038,In_448,In_764);
nand U4039 (N_4039,In_275,In_675);
nand U4040 (N_4040,In_252,In_320);
and U4041 (N_4041,In_915,In_953);
nor U4042 (N_4042,In_340,In_49);
nor U4043 (N_4043,In_1367,In_850);
nor U4044 (N_4044,In_817,In_401);
and U4045 (N_4045,In_998,In_36);
nor U4046 (N_4046,In_307,In_460);
or U4047 (N_4047,In_0,In_567);
nor U4048 (N_4048,In_1160,In_45);
nand U4049 (N_4049,In_932,In_1244);
nand U4050 (N_4050,In_1160,In_161);
or U4051 (N_4051,In_1253,In_305);
and U4052 (N_4052,In_1210,In_797);
and U4053 (N_4053,In_837,In_1103);
and U4054 (N_4054,In_622,In_130);
and U4055 (N_4055,In_482,In_754);
and U4056 (N_4056,In_908,In_835);
and U4057 (N_4057,In_453,In_877);
nand U4058 (N_4058,In_1236,In_728);
and U4059 (N_4059,In_504,In_54);
and U4060 (N_4060,In_737,In_682);
nand U4061 (N_4061,In_1111,In_1302);
and U4062 (N_4062,In_185,In_557);
nor U4063 (N_4063,In_179,In_1412);
xnor U4064 (N_4064,In_226,In_683);
and U4065 (N_4065,In_209,In_81);
or U4066 (N_4066,In_1333,In_722);
or U4067 (N_4067,In_532,In_891);
nor U4068 (N_4068,In_65,In_1296);
and U4069 (N_4069,In_1292,In_1017);
or U4070 (N_4070,In_1306,In_900);
and U4071 (N_4071,In_772,In_337);
nand U4072 (N_4072,In_699,In_1315);
nor U4073 (N_4073,In_1112,In_921);
nor U4074 (N_4074,In_102,In_1265);
or U4075 (N_4075,In_1055,In_881);
nand U4076 (N_4076,In_496,In_308);
and U4077 (N_4077,In_787,In_1310);
and U4078 (N_4078,In_907,In_1073);
nand U4079 (N_4079,In_717,In_1338);
nand U4080 (N_4080,In_1285,In_476);
nor U4081 (N_4081,In_308,In_1431);
or U4082 (N_4082,In_274,In_383);
and U4083 (N_4083,In_1246,In_1299);
or U4084 (N_4084,In_1086,In_1329);
and U4085 (N_4085,In_72,In_710);
or U4086 (N_4086,In_613,In_1009);
nor U4087 (N_4087,In_244,In_921);
and U4088 (N_4088,In_774,In_677);
and U4089 (N_4089,In_1085,In_940);
and U4090 (N_4090,In_1436,In_969);
nand U4091 (N_4091,In_1270,In_631);
and U4092 (N_4092,In_1360,In_437);
nor U4093 (N_4093,In_1141,In_870);
nor U4094 (N_4094,In_307,In_436);
or U4095 (N_4095,In_1427,In_1299);
or U4096 (N_4096,In_359,In_1018);
nor U4097 (N_4097,In_485,In_442);
nor U4098 (N_4098,In_633,In_1461);
nor U4099 (N_4099,In_27,In_1221);
or U4100 (N_4100,In_1361,In_144);
nor U4101 (N_4101,In_1064,In_1016);
or U4102 (N_4102,In_909,In_1023);
nand U4103 (N_4103,In_330,In_1375);
nor U4104 (N_4104,In_578,In_155);
nand U4105 (N_4105,In_800,In_1079);
and U4106 (N_4106,In_253,In_907);
or U4107 (N_4107,In_910,In_939);
xor U4108 (N_4108,In_1254,In_1103);
nor U4109 (N_4109,In_490,In_1048);
or U4110 (N_4110,In_61,In_1224);
or U4111 (N_4111,In_1355,In_38);
and U4112 (N_4112,In_432,In_313);
and U4113 (N_4113,In_813,In_589);
or U4114 (N_4114,In_1449,In_846);
nand U4115 (N_4115,In_1369,In_1115);
and U4116 (N_4116,In_650,In_499);
nor U4117 (N_4117,In_198,In_282);
nor U4118 (N_4118,In_1142,In_742);
and U4119 (N_4119,In_731,In_152);
or U4120 (N_4120,In_1241,In_381);
nand U4121 (N_4121,In_1288,In_778);
nor U4122 (N_4122,In_299,In_167);
or U4123 (N_4123,In_1484,In_1120);
or U4124 (N_4124,In_136,In_63);
and U4125 (N_4125,In_425,In_51);
and U4126 (N_4126,In_224,In_177);
or U4127 (N_4127,In_984,In_577);
nand U4128 (N_4128,In_1239,In_119);
and U4129 (N_4129,In_631,In_1102);
nand U4130 (N_4130,In_426,In_1108);
and U4131 (N_4131,In_870,In_116);
or U4132 (N_4132,In_791,In_1003);
and U4133 (N_4133,In_489,In_237);
or U4134 (N_4134,In_447,In_70);
or U4135 (N_4135,In_102,In_335);
nand U4136 (N_4136,In_689,In_311);
and U4137 (N_4137,In_1065,In_1064);
or U4138 (N_4138,In_206,In_1207);
nor U4139 (N_4139,In_436,In_754);
nor U4140 (N_4140,In_592,In_533);
or U4141 (N_4141,In_930,In_437);
and U4142 (N_4142,In_783,In_914);
xor U4143 (N_4143,In_81,In_580);
nand U4144 (N_4144,In_1044,In_315);
nand U4145 (N_4145,In_1187,In_279);
and U4146 (N_4146,In_803,In_1032);
nand U4147 (N_4147,In_609,In_338);
xnor U4148 (N_4148,In_655,In_458);
nand U4149 (N_4149,In_222,In_1215);
and U4150 (N_4150,In_1468,In_830);
nand U4151 (N_4151,In_1406,In_366);
nor U4152 (N_4152,In_1427,In_952);
nor U4153 (N_4153,In_926,In_1302);
or U4154 (N_4154,In_105,In_1125);
nand U4155 (N_4155,In_541,In_1116);
or U4156 (N_4156,In_606,In_1221);
nand U4157 (N_4157,In_1458,In_835);
nand U4158 (N_4158,In_424,In_340);
or U4159 (N_4159,In_1181,In_532);
nand U4160 (N_4160,In_247,In_246);
and U4161 (N_4161,In_1044,In_1378);
nor U4162 (N_4162,In_1308,In_554);
and U4163 (N_4163,In_1126,In_1084);
and U4164 (N_4164,In_345,In_383);
nor U4165 (N_4165,In_115,In_653);
nor U4166 (N_4166,In_535,In_826);
nand U4167 (N_4167,In_682,In_608);
or U4168 (N_4168,In_1079,In_167);
and U4169 (N_4169,In_1254,In_292);
and U4170 (N_4170,In_886,In_677);
nand U4171 (N_4171,In_992,In_486);
and U4172 (N_4172,In_1468,In_305);
or U4173 (N_4173,In_189,In_22);
nor U4174 (N_4174,In_1487,In_1254);
and U4175 (N_4175,In_93,In_1075);
or U4176 (N_4176,In_1487,In_1046);
and U4177 (N_4177,In_928,In_258);
or U4178 (N_4178,In_35,In_1272);
nor U4179 (N_4179,In_1030,In_1240);
and U4180 (N_4180,In_325,In_541);
nand U4181 (N_4181,In_1440,In_681);
nand U4182 (N_4182,In_140,In_354);
nor U4183 (N_4183,In_1270,In_459);
and U4184 (N_4184,In_1466,In_1197);
nand U4185 (N_4185,In_1400,In_701);
or U4186 (N_4186,In_78,In_560);
and U4187 (N_4187,In_675,In_1293);
nand U4188 (N_4188,In_617,In_386);
or U4189 (N_4189,In_648,In_454);
nand U4190 (N_4190,In_445,In_347);
nor U4191 (N_4191,In_592,In_1060);
or U4192 (N_4192,In_1477,In_902);
nand U4193 (N_4193,In_47,In_390);
nor U4194 (N_4194,In_1482,In_300);
or U4195 (N_4195,In_318,In_523);
nand U4196 (N_4196,In_81,In_74);
and U4197 (N_4197,In_1099,In_630);
and U4198 (N_4198,In_477,In_1444);
nor U4199 (N_4199,In_784,In_937);
nor U4200 (N_4200,In_709,In_126);
or U4201 (N_4201,In_1216,In_992);
nand U4202 (N_4202,In_38,In_937);
nand U4203 (N_4203,In_943,In_656);
nand U4204 (N_4204,In_876,In_863);
or U4205 (N_4205,In_32,In_114);
and U4206 (N_4206,In_719,In_1437);
nand U4207 (N_4207,In_1215,In_532);
nand U4208 (N_4208,In_1387,In_930);
and U4209 (N_4209,In_581,In_1406);
and U4210 (N_4210,In_643,In_662);
nand U4211 (N_4211,In_782,In_544);
nor U4212 (N_4212,In_1163,In_243);
and U4213 (N_4213,In_1470,In_1003);
nor U4214 (N_4214,In_638,In_1422);
and U4215 (N_4215,In_792,In_242);
or U4216 (N_4216,In_643,In_1154);
nand U4217 (N_4217,In_300,In_1080);
xnor U4218 (N_4218,In_707,In_781);
nor U4219 (N_4219,In_87,In_289);
or U4220 (N_4220,In_1175,In_354);
nand U4221 (N_4221,In_1349,In_815);
and U4222 (N_4222,In_1313,In_440);
nor U4223 (N_4223,In_865,In_204);
or U4224 (N_4224,In_453,In_1308);
and U4225 (N_4225,In_528,In_1431);
and U4226 (N_4226,In_432,In_1041);
nor U4227 (N_4227,In_498,In_91);
nand U4228 (N_4228,In_1049,In_1419);
nor U4229 (N_4229,In_1082,In_701);
nand U4230 (N_4230,In_680,In_871);
and U4231 (N_4231,In_575,In_154);
and U4232 (N_4232,In_718,In_664);
or U4233 (N_4233,In_1137,In_913);
nor U4234 (N_4234,In_528,In_1379);
and U4235 (N_4235,In_1023,In_445);
nand U4236 (N_4236,In_1364,In_1017);
nand U4237 (N_4237,In_113,In_1269);
and U4238 (N_4238,In_172,In_1235);
nand U4239 (N_4239,In_309,In_734);
nor U4240 (N_4240,In_435,In_712);
nand U4241 (N_4241,In_1415,In_1021);
nand U4242 (N_4242,In_670,In_1313);
and U4243 (N_4243,In_25,In_52);
or U4244 (N_4244,In_501,In_648);
or U4245 (N_4245,In_858,In_13);
or U4246 (N_4246,In_803,In_999);
or U4247 (N_4247,In_157,In_692);
nor U4248 (N_4248,In_708,In_794);
nand U4249 (N_4249,In_377,In_1277);
or U4250 (N_4250,In_660,In_176);
nand U4251 (N_4251,In_160,In_734);
nand U4252 (N_4252,In_1037,In_921);
nand U4253 (N_4253,In_1081,In_1044);
nand U4254 (N_4254,In_1240,In_122);
nor U4255 (N_4255,In_946,In_1374);
nor U4256 (N_4256,In_1189,In_76);
nor U4257 (N_4257,In_1251,In_705);
and U4258 (N_4258,In_150,In_1338);
or U4259 (N_4259,In_1345,In_97);
nor U4260 (N_4260,In_792,In_718);
nand U4261 (N_4261,In_981,In_1492);
and U4262 (N_4262,In_797,In_812);
and U4263 (N_4263,In_1325,In_1133);
nand U4264 (N_4264,In_927,In_819);
xnor U4265 (N_4265,In_434,In_287);
or U4266 (N_4266,In_486,In_1135);
or U4267 (N_4267,In_1391,In_661);
and U4268 (N_4268,In_1141,In_474);
or U4269 (N_4269,In_1292,In_1065);
nor U4270 (N_4270,In_907,In_504);
and U4271 (N_4271,In_194,In_1302);
or U4272 (N_4272,In_510,In_218);
and U4273 (N_4273,In_943,In_762);
nand U4274 (N_4274,In_410,In_449);
or U4275 (N_4275,In_982,In_423);
and U4276 (N_4276,In_765,In_345);
and U4277 (N_4277,In_699,In_497);
nand U4278 (N_4278,In_881,In_65);
and U4279 (N_4279,In_641,In_946);
nor U4280 (N_4280,In_1034,In_1068);
or U4281 (N_4281,In_834,In_178);
nand U4282 (N_4282,In_845,In_475);
and U4283 (N_4283,In_376,In_570);
nand U4284 (N_4284,In_734,In_863);
nor U4285 (N_4285,In_461,In_181);
or U4286 (N_4286,In_1280,In_67);
nor U4287 (N_4287,In_1086,In_216);
and U4288 (N_4288,In_356,In_82);
nand U4289 (N_4289,In_1322,In_1219);
nor U4290 (N_4290,In_428,In_398);
nor U4291 (N_4291,In_302,In_1450);
nor U4292 (N_4292,In_1489,In_475);
and U4293 (N_4293,In_857,In_1390);
nor U4294 (N_4294,In_1340,In_1353);
nor U4295 (N_4295,In_41,In_944);
and U4296 (N_4296,In_1214,In_71);
xnor U4297 (N_4297,In_576,In_763);
or U4298 (N_4298,In_1080,In_848);
or U4299 (N_4299,In_1142,In_176);
nor U4300 (N_4300,In_1216,In_614);
or U4301 (N_4301,In_1100,In_840);
nor U4302 (N_4302,In_874,In_1283);
nor U4303 (N_4303,In_898,In_1078);
or U4304 (N_4304,In_1341,In_1329);
or U4305 (N_4305,In_1241,In_761);
nor U4306 (N_4306,In_478,In_666);
and U4307 (N_4307,In_17,In_737);
nand U4308 (N_4308,In_1315,In_743);
nand U4309 (N_4309,In_671,In_1419);
or U4310 (N_4310,In_1407,In_798);
and U4311 (N_4311,In_24,In_1153);
nor U4312 (N_4312,In_54,In_320);
nand U4313 (N_4313,In_369,In_21);
or U4314 (N_4314,In_298,In_776);
or U4315 (N_4315,In_967,In_1045);
or U4316 (N_4316,In_1469,In_847);
and U4317 (N_4317,In_845,In_1103);
or U4318 (N_4318,In_1083,In_1397);
and U4319 (N_4319,In_305,In_415);
and U4320 (N_4320,In_101,In_937);
or U4321 (N_4321,In_742,In_579);
or U4322 (N_4322,In_320,In_1032);
nor U4323 (N_4323,In_1371,In_354);
and U4324 (N_4324,In_466,In_1416);
or U4325 (N_4325,In_495,In_1396);
nor U4326 (N_4326,In_134,In_533);
nand U4327 (N_4327,In_1402,In_17);
and U4328 (N_4328,In_544,In_88);
nand U4329 (N_4329,In_847,In_132);
or U4330 (N_4330,In_9,In_592);
xor U4331 (N_4331,In_905,In_1350);
nand U4332 (N_4332,In_743,In_112);
and U4333 (N_4333,In_150,In_440);
or U4334 (N_4334,In_739,In_1083);
or U4335 (N_4335,In_1138,In_634);
and U4336 (N_4336,In_111,In_385);
and U4337 (N_4337,In_1131,In_232);
nor U4338 (N_4338,In_200,In_83);
nand U4339 (N_4339,In_164,In_350);
and U4340 (N_4340,In_76,In_1219);
nor U4341 (N_4341,In_705,In_345);
or U4342 (N_4342,In_1198,In_1452);
xnor U4343 (N_4343,In_1012,In_710);
and U4344 (N_4344,In_1236,In_9);
and U4345 (N_4345,In_663,In_1002);
nor U4346 (N_4346,In_427,In_1442);
or U4347 (N_4347,In_1019,In_277);
nand U4348 (N_4348,In_589,In_757);
or U4349 (N_4349,In_71,In_219);
nand U4350 (N_4350,In_412,In_1090);
nor U4351 (N_4351,In_680,In_955);
or U4352 (N_4352,In_807,In_673);
and U4353 (N_4353,In_817,In_1427);
nand U4354 (N_4354,In_488,In_1322);
nor U4355 (N_4355,In_581,In_1347);
or U4356 (N_4356,In_1248,In_1030);
or U4357 (N_4357,In_1135,In_1145);
nor U4358 (N_4358,In_539,In_13);
and U4359 (N_4359,In_949,In_1094);
and U4360 (N_4360,In_1457,In_151);
nor U4361 (N_4361,In_388,In_1168);
nand U4362 (N_4362,In_1245,In_161);
nand U4363 (N_4363,In_100,In_1118);
and U4364 (N_4364,In_382,In_146);
nand U4365 (N_4365,In_1499,In_454);
nand U4366 (N_4366,In_958,In_1432);
nand U4367 (N_4367,In_1265,In_1450);
nand U4368 (N_4368,In_88,In_382);
nor U4369 (N_4369,In_844,In_361);
nand U4370 (N_4370,In_1326,In_1443);
or U4371 (N_4371,In_741,In_627);
nand U4372 (N_4372,In_377,In_1269);
or U4373 (N_4373,In_268,In_980);
nor U4374 (N_4374,In_1280,In_1013);
nor U4375 (N_4375,In_408,In_727);
or U4376 (N_4376,In_739,In_13);
nor U4377 (N_4377,In_1179,In_1037);
nor U4378 (N_4378,In_1353,In_18);
nand U4379 (N_4379,In_326,In_1412);
and U4380 (N_4380,In_425,In_912);
and U4381 (N_4381,In_836,In_77);
nand U4382 (N_4382,In_1054,In_732);
nor U4383 (N_4383,In_29,In_746);
and U4384 (N_4384,In_1430,In_54);
nor U4385 (N_4385,In_340,In_688);
or U4386 (N_4386,In_1225,In_1307);
nor U4387 (N_4387,In_331,In_1331);
nand U4388 (N_4388,In_298,In_977);
or U4389 (N_4389,In_1360,In_13);
nor U4390 (N_4390,In_1340,In_512);
nor U4391 (N_4391,In_1452,In_838);
nand U4392 (N_4392,In_748,In_1426);
or U4393 (N_4393,In_1194,In_799);
nor U4394 (N_4394,In_378,In_1402);
or U4395 (N_4395,In_468,In_302);
nand U4396 (N_4396,In_1084,In_865);
nand U4397 (N_4397,In_825,In_425);
nor U4398 (N_4398,In_217,In_615);
nand U4399 (N_4399,In_526,In_49);
nor U4400 (N_4400,In_919,In_1135);
xor U4401 (N_4401,In_561,In_196);
nor U4402 (N_4402,In_517,In_934);
nor U4403 (N_4403,In_174,In_523);
and U4404 (N_4404,In_625,In_499);
and U4405 (N_4405,In_39,In_321);
nand U4406 (N_4406,In_1427,In_54);
nand U4407 (N_4407,In_1180,In_1220);
or U4408 (N_4408,In_218,In_117);
and U4409 (N_4409,In_996,In_376);
nor U4410 (N_4410,In_1438,In_334);
and U4411 (N_4411,In_839,In_1142);
nand U4412 (N_4412,In_1444,In_716);
nor U4413 (N_4413,In_656,In_1380);
nor U4414 (N_4414,In_317,In_1418);
nor U4415 (N_4415,In_359,In_725);
nor U4416 (N_4416,In_66,In_195);
nand U4417 (N_4417,In_113,In_904);
nand U4418 (N_4418,In_475,In_1332);
nand U4419 (N_4419,In_1115,In_740);
nor U4420 (N_4420,In_620,In_1187);
or U4421 (N_4421,In_761,In_23);
nor U4422 (N_4422,In_605,In_437);
or U4423 (N_4423,In_233,In_481);
nand U4424 (N_4424,In_749,In_548);
and U4425 (N_4425,In_788,In_496);
and U4426 (N_4426,In_340,In_1074);
or U4427 (N_4427,In_639,In_336);
nand U4428 (N_4428,In_866,In_750);
nand U4429 (N_4429,In_287,In_607);
and U4430 (N_4430,In_722,In_325);
and U4431 (N_4431,In_948,In_374);
and U4432 (N_4432,In_861,In_819);
nor U4433 (N_4433,In_1329,In_1158);
and U4434 (N_4434,In_874,In_653);
nor U4435 (N_4435,In_1165,In_387);
nor U4436 (N_4436,In_824,In_334);
nand U4437 (N_4437,In_1325,In_1224);
and U4438 (N_4438,In_893,In_1349);
nor U4439 (N_4439,In_1252,In_672);
nand U4440 (N_4440,In_27,In_1405);
nor U4441 (N_4441,In_679,In_1209);
and U4442 (N_4442,In_532,In_621);
nor U4443 (N_4443,In_333,In_728);
and U4444 (N_4444,In_481,In_275);
and U4445 (N_4445,In_792,In_1288);
nand U4446 (N_4446,In_1128,In_1309);
nand U4447 (N_4447,In_716,In_911);
nor U4448 (N_4448,In_243,In_816);
and U4449 (N_4449,In_1478,In_797);
and U4450 (N_4450,In_1024,In_495);
nand U4451 (N_4451,In_136,In_535);
nand U4452 (N_4452,In_584,In_794);
nor U4453 (N_4453,In_867,In_1008);
or U4454 (N_4454,In_844,In_1085);
nand U4455 (N_4455,In_617,In_1214);
or U4456 (N_4456,In_832,In_1177);
or U4457 (N_4457,In_222,In_831);
or U4458 (N_4458,In_704,In_766);
and U4459 (N_4459,In_416,In_1351);
nand U4460 (N_4460,In_19,In_1263);
or U4461 (N_4461,In_69,In_154);
or U4462 (N_4462,In_1236,In_509);
nand U4463 (N_4463,In_1205,In_1172);
and U4464 (N_4464,In_885,In_750);
nor U4465 (N_4465,In_560,In_1379);
nand U4466 (N_4466,In_736,In_744);
or U4467 (N_4467,In_898,In_153);
or U4468 (N_4468,In_342,In_502);
or U4469 (N_4469,In_840,In_774);
and U4470 (N_4470,In_378,In_712);
and U4471 (N_4471,In_1253,In_197);
nand U4472 (N_4472,In_1419,In_909);
and U4473 (N_4473,In_684,In_105);
nor U4474 (N_4474,In_527,In_1402);
nor U4475 (N_4475,In_1159,In_1124);
nand U4476 (N_4476,In_1204,In_1193);
nand U4477 (N_4477,In_1345,In_567);
and U4478 (N_4478,In_422,In_309);
nand U4479 (N_4479,In_422,In_477);
nand U4480 (N_4480,In_1466,In_1031);
nor U4481 (N_4481,In_134,In_1487);
and U4482 (N_4482,In_1017,In_1019);
nand U4483 (N_4483,In_709,In_447);
or U4484 (N_4484,In_538,In_668);
nand U4485 (N_4485,In_927,In_601);
and U4486 (N_4486,In_1236,In_566);
and U4487 (N_4487,In_1489,In_1142);
nor U4488 (N_4488,In_760,In_1491);
or U4489 (N_4489,In_735,In_61);
nor U4490 (N_4490,In_318,In_370);
nor U4491 (N_4491,In_451,In_458);
nand U4492 (N_4492,In_141,In_966);
and U4493 (N_4493,In_980,In_832);
or U4494 (N_4494,In_121,In_622);
nor U4495 (N_4495,In_1324,In_586);
or U4496 (N_4496,In_239,In_785);
nor U4497 (N_4497,In_491,In_810);
nand U4498 (N_4498,In_633,In_864);
nand U4499 (N_4499,In_239,In_1116);
nor U4500 (N_4500,In_99,In_327);
nor U4501 (N_4501,In_1204,In_1071);
or U4502 (N_4502,In_216,In_323);
nand U4503 (N_4503,In_1053,In_306);
nand U4504 (N_4504,In_484,In_1003);
nor U4505 (N_4505,In_1207,In_737);
or U4506 (N_4506,In_74,In_1471);
nand U4507 (N_4507,In_1057,In_797);
nand U4508 (N_4508,In_38,In_619);
nor U4509 (N_4509,In_171,In_1444);
nor U4510 (N_4510,In_1109,In_580);
nor U4511 (N_4511,In_419,In_1086);
nor U4512 (N_4512,In_822,In_1402);
nand U4513 (N_4513,In_204,In_1346);
or U4514 (N_4514,In_1326,In_382);
and U4515 (N_4515,In_1163,In_570);
or U4516 (N_4516,In_926,In_77);
nand U4517 (N_4517,In_954,In_1250);
nor U4518 (N_4518,In_962,In_38);
nand U4519 (N_4519,In_1351,In_562);
nor U4520 (N_4520,In_114,In_301);
or U4521 (N_4521,In_458,In_1040);
and U4522 (N_4522,In_783,In_588);
and U4523 (N_4523,In_105,In_62);
or U4524 (N_4524,In_212,In_1090);
nor U4525 (N_4525,In_925,In_1106);
and U4526 (N_4526,In_226,In_1082);
or U4527 (N_4527,In_682,In_1456);
nor U4528 (N_4528,In_1149,In_388);
or U4529 (N_4529,In_1446,In_1157);
or U4530 (N_4530,In_498,In_127);
nor U4531 (N_4531,In_317,In_1107);
or U4532 (N_4532,In_502,In_1151);
nor U4533 (N_4533,In_19,In_6);
nand U4534 (N_4534,In_744,In_729);
nand U4535 (N_4535,In_1313,In_1383);
or U4536 (N_4536,In_173,In_512);
nor U4537 (N_4537,In_684,In_532);
and U4538 (N_4538,In_1304,In_864);
and U4539 (N_4539,In_335,In_215);
nor U4540 (N_4540,In_1303,In_70);
or U4541 (N_4541,In_873,In_1486);
nor U4542 (N_4542,In_1058,In_1165);
nand U4543 (N_4543,In_449,In_1372);
nor U4544 (N_4544,In_1079,In_1405);
or U4545 (N_4545,In_1242,In_21);
nor U4546 (N_4546,In_963,In_757);
or U4547 (N_4547,In_1491,In_214);
nor U4548 (N_4548,In_1128,In_128);
or U4549 (N_4549,In_672,In_1105);
nand U4550 (N_4550,In_534,In_913);
nand U4551 (N_4551,In_1248,In_559);
and U4552 (N_4552,In_685,In_213);
nor U4553 (N_4553,In_1302,In_1363);
or U4554 (N_4554,In_1269,In_1099);
nand U4555 (N_4555,In_168,In_890);
and U4556 (N_4556,In_1193,In_453);
nor U4557 (N_4557,In_1413,In_1410);
nor U4558 (N_4558,In_123,In_288);
nor U4559 (N_4559,In_321,In_245);
nand U4560 (N_4560,In_1114,In_392);
or U4561 (N_4561,In_479,In_1393);
and U4562 (N_4562,In_1277,In_1184);
and U4563 (N_4563,In_867,In_586);
or U4564 (N_4564,In_1477,In_546);
or U4565 (N_4565,In_298,In_629);
nand U4566 (N_4566,In_542,In_93);
or U4567 (N_4567,In_139,In_771);
or U4568 (N_4568,In_1067,In_1383);
nand U4569 (N_4569,In_1174,In_1022);
nor U4570 (N_4570,In_1352,In_891);
xnor U4571 (N_4571,In_1422,In_1322);
and U4572 (N_4572,In_1394,In_892);
nor U4573 (N_4573,In_1214,In_1068);
or U4574 (N_4574,In_647,In_1215);
or U4575 (N_4575,In_1410,In_162);
or U4576 (N_4576,In_241,In_670);
and U4577 (N_4577,In_602,In_898);
nand U4578 (N_4578,In_1141,In_1228);
or U4579 (N_4579,In_1017,In_920);
or U4580 (N_4580,In_444,In_924);
nand U4581 (N_4581,In_1425,In_1492);
nand U4582 (N_4582,In_706,In_12);
nor U4583 (N_4583,In_699,In_1475);
nor U4584 (N_4584,In_896,In_829);
nor U4585 (N_4585,In_631,In_516);
or U4586 (N_4586,In_1268,In_204);
or U4587 (N_4587,In_1312,In_672);
nor U4588 (N_4588,In_343,In_241);
nand U4589 (N_4589,In_512,In_704);
and U4590 (N_4590,In_1463,In_62);
nand U4591 (N_4591,In_334,In_690);
nand U4592 (N_4592,In_398,In_1452);
nand U4593 (N_4593,In_535,In_982);
and U4594 (N_4594,In_178,In_1028);
or U4595 (N_4595,In_63,In_319);
nand U4596 (N_4596,In_185,In_811);
nand U4597 (N_4597,In_531,In_498);
nor U4598 (N_4598,In_518,In_406);
nor U4599 (N_4599,In_836,In_1415);
or U4600 (N_4600,In_238,In_717);
nor U4601 (N_4601,In_674,In_832);
and U4602 (N_4602,In_1346,In_1405);
nor U4603 (N_4603,In_1343,In_299);
nand U4604 (N_4604,In_708,In_903);
nand U4605 (N_4605,In_908,In_1040);
nand U4606 (N_4606,In_1103,In_169);
nand U4607 (N_4607,In_356,In_224);
and U4608 (N_4608,In_243,In_528);
or U4609 (N_4609,In_948,In_908);
nor U4610 (N_4610,In_1395,In_302);
nor U4611 (N_4611,In_508,In_1248);
and U4612 (N_4612,In_1311,In_904);
nand U4613 (N_4613,In_1188,In_1178);
nor U4614 (N_4614,In_1155,In_534);
or U4615 (N_4615,In_169,In_139);
or U4616 (N_4616,In_46,In_783);
nor U4617 (N_4617,In_283,In_878);
nand U4618 (N_4618,In_55,In_995);
and U4619 (N_4619,In_1330,In_199);
nor U4620 (N_4620,In_33,In_832);
and U4621 (N_4621,In_2,In_584);
nand U4622 (N_4622,In_1400,In_1445);
and U4623 (N_4623,In_691,In_1039);
nand U4624 (N_4624,In_1132,In_409);
or U4625 (N_4625,In_645,In_1073);
nor U4626 (N_4626,In_528,In_363);
or U4627 (N_4627,In_679,In_747);
and U4628 (N_4628,In_1198,In_1280);
and U4629 (N_4629,In_123,In_23);
or U4630 (N_4630,In_554,In_546);
nand U4631 (N_4631,In_602,In_1247);
nor U4632 (N_4632,In_376,In_860);
nor U4633 (N_4633,In_1192,In_880);
nor U4634 (N_4634,In_95,In_1026);
and U4635 (N_4635,In_199,In_705);
or U4636 (N_4636,In_1354,In_231);
nor U4637 (N_4637,In_1138,In_731);
or U4638 (N_4638,In_47,In_321);
or U4639 (N_4639,In_1289,In_619);
nor U4640 (N_4640,In_1224,In_39);
nand U4641 (N_4641,In_736,In_83);
or U4642 (N_4642,In_1473,In_1178);
or U4643 (N_4643,In_1122,In_1144);
or U4644 (N_4644,In_639,In_85);
and U4645 (N_4645,In_1353,In_50);
nor U4646 (N_4646,In_443,In_1082);
and U4647 (N_4647,In_1082,In_499);
nor U4648 (N_4648,In_205,In_393);
nor U4649 (N_4649,In_623,In_1123);
and U4650 (N_4650,In_71,In_244);
nor U4651 (N_4651,In_104,In_412);
nand U4652 (N_4652,In_1257,In_992);
and U4653 (N_4653,In_818,In_1101);
or U4654 (N_4654,In_356,In_1412);
nor U4655 (N_4655,In_1189,In_1020);
nand U4656 (N_4656,In_1279,In_119);
nand U4657 (N_4657,In_1074,In_1125);
or U4658 (N_4658,In_656,In_639);
nor U4659 (N_4659,In_374,In_1165);
or U4660 (N_4660,In_1120,In_425);
nor U4661 (N_4661,In_1003,In_1077);
nand U4662 (N_4662,In_1438,In_953);
nand U4663 (N_4663,In_1383,In_207);
nor U4664 (N_4664,In_1210,In_320);
nor U4665 (N_4665,In_353,In_1285);
and U4666 (N_4666,In_1015,In_1118);
nor U4667 (N_4667,In_1118,In_59);
nand U4668 (N_4668,In_1442,In_181);
nor U4669 (N_4669,In_1340,In_1489);
nor U4670 (N_4670,In_413,In_1469);
or U4671 (N_4671,In_859,In_443);
and U4672 (N_4672,In_1274,In_1455);
or U4673 (N_4673,In_577,In_612);
and U4674 (N_4674,In_1386,In_496);
and U4675 (N_4675,In_296,In_785);
or U4676 (N_4676,In_1010,In_647);
nor U4677 (N_4677,In_724,In_950);
nand U4678 (N_4678,In_4,In_159);
or U4679 (N_4679,In_1025,In_513);
and U4680 (N_4680,In_327,In_660);
and U4681 (N_4681,In_1008,In_191);
nor U4682 (N_4682,In_285,In_62);
or U4683 (N_4683,In_267,In_1411);
nand U4684 (N_4684,In_1372,In_309);
nand U4685 (N_4685,In_921,In_669);
nor U4686 (N_4686,In_414,In_366);
and U4687 (N_4687,In_519,In_873);
nor U4688 (N_4688,In_1258,In_1460);
nor U4689 (N_4689,In_449,In_835);
nor U4690 (N_4690,In_612,In_65);
or U4691 (N_4691,In_1348,In_1057);
nand U4692 (N_4692,In_933,In_544);
nand U4693 (N_4693,In_772,In_917);
nand U4694 (N_4694,In_1449,In_159);
nand U4695 (N_4695,In_517,In_263);
or U4696 (N_4696,In_167,In_4);
xnor U4697 (N_4697,In_1292,In_63);
and U4698 (N_4698,In_1179,In_711);
or U4699 (N_4699,In_69,In_906);
nor U4700 (N_4700,In_258,In_1461);
nand U4701 (N_4701,In_1277,In_671);
or U4702 (N_4702,In_1061,In_637);
nor U4703 (N_4703,In_906,In_1101);
nand U4704 (N_4704,In_523,In_603);
and U4705 (N_4705,In_34,In_1075);
nand U4706 (N_4706,In_949,In_1028);
nand U4707 (N_4707,In_1339,In_495);
nor U4708 (N_4708,In_449,In_1086);
nand U4709 (N_4709,In_130,In_829);
nor U4710 (N_4710,In_81,In_1429);
and U4711 (N_4711,In_1388,In_53);
or U4712 (N_4712,In_1115,In_831);
or U4713 (N_4713,In_422,In_600);
or U4714 (N_4714,In_1368,In_196);
or U4715 (N_4715,In_1219,In_1382);
and U4716 (N_4716,In_885,In_150);
nand U4717 (N_4717,In_1333,In_376);
and U4718 (N_4718,In_365,In_206);
nand U4719 (N_4719,In_311,In_1046);
and U4720 (N_4720,In_842,In_576);
nand U4721 (N_4721,In_727,In_1322);
and U4722 (N_4722,In_375,In_22);
nor U4723 (N_4723,In_313,In_1386);
nor U4724 (N_4724,In_884,In_219);
or U4725 (N_4725,In_634,In_919);
and U4726 (N_4726,In_163,In_304);
nor U4727 (N_4727,In_370,In_716);
and U4728 (N_4728,In_812,In_731);
nor U4729 (N_4729,In_1123,In_1435);
nand U4730 (N_4730,In_130,In_792);
nor U4731 (N_4731,In_1201,In_940);
nor U4732 (N_4732,In_1451,In_396);
nand U4733 (N_4733,In_129,In_1314);
and U4734 (N_4734,In_511,In_94);
and U4735 (N_4735,In_1021,In_1282);
and U4736 (N_4736,In_593,In_1386);
nor U4737 (N_4737,In_1340,In_1449);
and U4738 (N_4738,In_833,In_1379);
nor U4739 (N_4739,In_541,In_1391);
nor U4740 (N_4740,In_258,In_1071);
nand U4741 (N_4741,In_320,In_996);
or U4742 (N_4742,In_1413,In_35);
and U4743 (N_4743,In_118,In_10);
or U4744 (N_4744,In_740,In_973);
nor U4745 (N_4745,In_898,In_1261);
or U4746 (N_4746,In_1445,In_846);
nor U4747 (N_4747,In_791,In_1168);
and U4748 (N_4748,In_131,In_1262);
nor U4749 (N_4749,In_739,In_2);
and U4750 (N_4750,In_506,In_440);
nand U4751 (N_4751,In_484,In_1);
nand U4752 (N_4752,In_709,In_1080);
nand U4753 (N_4753,In_1205,In_471);
nor U4754 (N_4754,In_466,In_1003);
and U4755 (N_4755,In_1393,In_874);
nand U4756 (N_4756,In_11,In_1289);
nand U4757 (N_4757,In_920,In_1358);
nand U4758 (N_4758,In_866,In_1040);
nand U4759 (N_4759,In_1110,In_172);
nand U4760 (N_4760,In_1280,In_379);
or U4761 (N_4761,In_937,In_1013);
nand U4762 (N_4762,In_668,In_1294);
and U4763 (N_4763,In_1092,In_1001);
and U4764 (N_4764,In_410,In_972);
or U4765 (N_4765,In_1355,In_572);
nor U4766 (N_4766,In_517,In_1353);
or U4767 (N_4767,In_1111,In_1184);
or U4768 (N_4768,In_1375,In_843);
nand U4769 (N_4769,In_1117,In_1006);
or U4770 (N_4770,In_1180,In_112);
nor U4771 (N_4771,In_355,In_1203);
or U4772 (N_4772,In_1479,In_954);
or U4773 (N_4773,In_6,In_1058);
nand U4774 (N_4774,In_335,In_110);
nor U4775 (N_4775,In_935,In_202);
nor U4776 (N_4776,In_857,In_1266);
nand U4777 (N_4777,In_124,In_89);
nor U4778 (N_4778,In_388,In_1170);
nand U4779 (N_4779,In_31,In_947);
nor U4780 (N_4780,In_1285,In_946);
nor U4781 (N_4781,In_785,In_920);
and U4782 (N_4782,In_1269,In_572);
and U4783 (N_4783,In_1286,In_1371);
or U4784 (N_4784,In_327,In_1433);
and U4785 (N_4785,In_348,In_478);
or U4786 (N_4786,In_929,In_729);
nor U4787 (N_4787,In_1305,In_206);
or U4788 (N_4788,In_1266,In_419);
nand U4789 (N_4789,In_314,In_388);
or U4790 (N_4790,In_797,In_171);
and U4791 (N_4791,In_1176,In_1281);
and U4792 (N_4792,In_550,In_429);
or U4793 (N_4793,In_0,In_1031);
or U4794 (N_4794,In_826,In_334);
nand U4795 (N_4795,In_1258,In_643);
nor U4796 (N_4796,In_188,In_263);
or U4797 (N_4797,In_1342,In_1380);
and U4798 (N_4798,In_1287,In_1165);
nand U4799 (N_4799,In_791,In_329);
or U4800 (N_4800,In_82,In_310);
nor U4801 (N_4801,In_395,In_709);
and U4802 (N_4802,In_884,In_843);
nand U4803 (N_4803,In_1009,In_305);
or U4804 (N_4804,In_533,In_735);
or U4805 (N_4805,In_342,In_914);
nor U4806 (N_4806,In_1427,In_921);
and U4807 (N_4807,In_699,In_770);
and U4808 (N_4808,In_999,In_909);
nand U4809 (N_4809,In_983,In_593);
nand U4810 (N_4810,In_1206,In_1264);
and U4811 (N_4811,In_856,In_481);
and U4812 (N_4812,In_334,In_353);
nand U4813 (N_4813,In_973,In_747);
xnor U4814 (N_4814,In_14,In_1321);
nand U4815 (N_4815,In_202,In_689);
nor U4816 (N_4816,In_673,In_698);
nand U4817 (N_4817,In_957,In_96);
and U4818 (N_4818,In_877,In_843);
or U4819 (N_4819,In_808,In_799);
and U4820 (N_4820,In_253,In_1173);
nor U4821 (N_4821,In_996,In_784);
nor U4822 (N_4822,In_101,In_400);
nand U4823 (N_4823,In_276,In_244);
nand U4824 (N_4824,In_1438,In_1223);
and U4825 (N_4825,In_262,In_1459);
nor U4826 (N_4826,In_662,In_1165);
or U4827 (N_4827,In_982,In_54);
nand U4828 (N_4828,In_493,In_137);
nand U4829 (N_4829,In_213,In_972);
and U4830 (N_4830,In_1480,In_500);
nor U4831 (N_4831,In_669,In_1265);
and U4832 (N_4832,In_1091,In_88);
or U4833 (N_4833,In_197,In_630);
or U4834 (N_4834,In_1303,In_852);
and U4835 (N_4835,In_1496,In_45);
nor U4836 (N_4836,In_1414,In_680);
or U4837 (N_4837,In_420,In_645);
and U4838 (N_4838,In_1140,In_506);
nor U4839 (N_4839,In_389,In_176);
nand U4840 (N_4840,In_950,In_1363);
nor U4841 (N_4841,In_1273,In_862);
nor U4842 (N_4842,In_484,In_1050);
nor U4843 (N_4843,In_1235,In_563);
and U4844 (N_4844,In_910,In_415);
nor U4845 (N_4845,In_1170,In_1381);
nor U4846 (N_4846,In_866,In_120);
nor U4847 (N_4847,In_932,In_1499);
and U4848 (N_4848,In_225,In_848);
and U4849 (N_4849,In_1363,In_1287);
nor U4850 (N_4850,In_940,In_1249);
nor U4851 (N_4851,In_573,In_1227);
and U4852 (N_4852,In_888,In_753);
or U4853 (N_4853,In_1445,In_1449);
nand U4854 (N_4854,In_927,In_1104);
nand U4855 (N_4855,In_296,In_53);
nand U4856 (N_4856,In_275,In_871);
and U4857 (N_4857,In_1232,In_867);
or U4858 (N_4858,In_272,In_362);
nand U4859 (N_4859,In_1073,In_574);
or U4860 (N_4860,In_1001,In_1464);
or U4861 (N_4861,In_81,In_1476);
or U4862 (N_4862,In_1187,In_1314);
nand U4863 (N_4863,In_104,In_1380);
or U4864 (N_4864,In_1175,In_261);
nand U4865 (N_4865,In_1189,In_727);
nor U4866 (N_4866,In_1003,In_507);
xnor U4867 (N_4867,In_926,In_656);
or U4868 (N_4868,In_784,In_549);
nor U4869 (N_4869,In_129,In_330);
and U4870 (N_4870,In_1473,In_1257);
and U4871 (N_4871,In_1180,In_1244);
or U4872 (N_4872,In_281,In_1026);
and U4873 (N_4873,In_1094,In_1347);
nor U4874 (N_4874,In_22,In_1475);
or U4875 (N_4875,In_541,In_191);
and U4876 (N_4876,In_1135,In_1329);
or U4877 (N_4877,In_228,In_237);
or U4878 (N_4878,In_297,In_570);
nand U4879 (N_4879,In_78,In_406);
or U4880 (N_4880,In_1286,In_1458);
nand U4881 (N_4881,In_1352,In_894);
or U4882 (N_4882,In_711,In_406);
nor U4883 (N_4883,In_372,In_1026);
or U4884 (N_4884,In_97,In_109);
nor U4885 (N_4885,In_1144,In_523);
nor U4886 (N_4886,In_615,In_728);
xor U4887 (N_4887,In_967,In_1137);
and U4888 (N_4888,In_428,In_525);
or U4889 (N_4889,In_1157,In_35);
or U4890 (N_4890,In_79,In_666);
and U4891 (N_4891,In_982,In_246);
nand U4892 (N_4892,In_731,In_1425);
or U4893 (N_4893,In_755,In_497);
and U4894 (N_4894,In_228,In_261);
nor U4895 (N_4895,In_1023,In_71);
nand U4896 (N_4896,In_406,In_1453);
nand U4897 (N_4897,In_1422,In_1230);
nor U4898 (N_4898,In_750,In_764);
nand U4899 (N_4899,In_1423,In_499);
and U4900 (N_4900,In_907,In_507);
and U4901 (N_4901,In_930,In_98);
or U4902 (N_4902,In_406,In_282);
nor U4903 (N_4903,In_47,In_817);
nand U4904 (N_4904,In_1454,In_413);
or U4905 (N_4905,In_1332,In_570);
nor U4906 (N_4906,In_60,In_208);
nor U4907 (N_4907,In_1000,In_40);
or U4908 (N_4908,In_868,In_1003);
and U4909 (N_4909,In_1160,In_968);
nand U4910 (N_4910,In_396,In_100);
or U4911 (N_4911,In_1031,In_969);
nand U4912 (N_4912,In_1317,In_299);
nor U4913 (N_4913,In_222,In_484);
or U4914 (N_4914,In_906,In_101);
nor U4915 (N_4915,In_820,In_1036);
or U4916 (N_4916,In_945,In_334);
or U4917 (N_4917,In_1318,In_1112);
nor U4918 (N_4918,In_771,In_248);
or U4919 (N_4919,In_1120,In_221);
nor U4920 (N_4920,In_945,In_172);
or U4921 (N_4921,In_289,In_406);
and U4922 (N_4922,In_983,In_1227);
nand U4923 (N_4923,In_303,In_562);
nor U4924 (N_4924,In_300,In_1443);
and U4925 (N_4925,In_1097,In_76);
or U4926 (N_4926,In_1104,In_1453);
or U4927 (N_4927,In_1212,In_972);
nand U4928 (N_4928,In_9,In_308);
and U4929 (N_4929,In_1084,In_1206);
nor U4930 (N_4930,In_1017,In_418);
nor U4931 (N_4931,In_592,In_577);
nor U4932 (N_4932,In_120,In_278);
or U4933 (N_4933,In_1327,In_345);
and U4934 (N_4934,In_847,In_750);
nand U4935 (N_4935,In_12,In_1307);
and U4936 (N_4936,In_982,In_773);
and U4937 (N_4937,In_500,In_180);
and U4938 (N_4938,In_1197,In_1429);
or U4939 (N_4939,In_800,In_202);
nor U4940 (N_4940,In_969,In_64);
and U4941 (N_4941,In_566,In_1142);
nand U4942 (N_4942,In_887,In_1230);
and U4943 (N_4943,In_519,In_634);
nor U4944 (N_4944,In_1089,In_267);
or U4945 (N_4945,In_1380,In_1096);
nor U4946 (N_4946,In_242,In_1157);
nor U4947 (N_4947,In_294,In_1482);
nand U4948 (N_4948,In_565,In_205);
nor U4949 (N_4949,In_1403,In_1194);
nor U4950 (N_4950,In_1312,In_812);
nand U4951 (N_4951,In_1230,In_1141);
or U4952 (N_4952,In_1006,In_947);
and U4953 (N_4953,In_655,In_754);
nor U4954 (N_4954,In_1054,In_1312);
and U4955 (N_4955,In_1375,In_589);
or U4956 (N_4956,In_1300,In_915);
and U4957 (N_4957,In_705,In_659);
or U4958 (N_4958,In_595,In_574);
nor U4959 (N_4959,In_969,In_782);
nor U4960 (N_4960,In_656,In_136);
nor U4961 (N_4961,In_572,In_1128);
and U4962 (N_4962,In_266,In_1379);
and U4963 (N_4963,In_1236,In_1230);
and U4964 (N_4964,In_988,In_570);
or U4965 (N_4965,In_235,In_859);
nor U4966 (N_4966,In_1028,In_604);
or U4967 (N_4967,In_261,In_970);
nand U4968 (N_4968,In_1389,In_702);
or U4969 (N_4969,In_702,In_1346);
and U4970 (N_4970,In_520,In_755);
nand U4971 (N_4971,In_1312,In_623);
and U4972 (N_4972,In_837,In_528);
nor U4973 (N_4973,In_316,In_551);
or U4974 (N_4974,In_703,In_685);
or U4975 (N_4975,In_647,In_76);
nor U4976 (N_4976,In_1227,In_1124);
and U4977 (N_4977,In_1260,In_255);
nor U4978 (N_4978,In_532,In_659);
and U4979 (N_4979,In_326,In_772);
nand U4980 (N_4980,In_78,In_1375);
and U4981 (N_4981,In_666,In_1380);
nor U4982 (N_4982,In_1425,In_447);
nand U4983 (N_4983,In_793,In_529);
nor U4984 (N_4984,In_1228,In_233);
nand U4985 (N_4985,In_469,In_920);
and U4986 (N_4986,In_359,In_515);
nor U4987 (N_4987,In_734,In_989);
nor U4988 (N_4988,In_1396,In_1029);
nor U4989 (N_4989,In_850,In_1461);
nor U4990 (N_4990,In_807,In_870);
nor U4991 (N_4991,In_1182,In_1444);
nor U4992 (N_4992,In_515,In_566);
nor U4993 (N_4993,In_809,In_480);
and U4994 (N_4994,In_808,In_820);
or U4995 (N_4995,In_509,In_474);
or U4996 (N_4996,In_935,In_867);
nor U4997 (N_4997,In_1421,In_107);
or U4998 (N_4998,In_1460,In_1308);
or U4999 (N_4999,In_297,In_304);
nor U5000 (N_5000,N_3857,N_2537);
or U5001 (N_5001,N_4811,N_3030);
nand U5002 (N_5002,N_1923,N_2526);
nor U5003 (N_5003,N_4425,N_735);
nand U5004 (N_5004,N_1289,N_3087);
or U5005 (N_5005,N_222,N_132);
nand U5006 (N_5006,N_960,N_4738);
and U5007 (N_5007,N_203,N_50);
and U5008 (N_5008,N_2734,N_3652);
or U5009 (N_5009,N_1027,N_4832);
or U5010 (N_5010,N_2903,N_4126);
nand U5011 (N_5011,N_3586,N_4391);
and U5012 (N_5012,N_335,N_4430);
nand U5013 (N_5013,N_4505,N_935);
and U5014 (N_5014,N_1160,N_1563);
nor U5015 (N_5015,N_4601,N_3106);
or U5016 (N_5016,N_612,N_556);
nor U5017 (N_5017,N_2943,N_1285);
nand U5018 (N_5018,N_2379,N_3972);
and U5019 (N_5019,N_2293,N_309);
nor U5020 (N_5020,N_3997,N_2969);
nand U5021 (N_5021,N_1817,N_3481);
or U5022 (N_5022,N_2487,N_3193);
nor U5023 (N_5023,N_421,N_3530);
nand U5024 (N_5024,N_312,N_413);
xor U5025 (N_5025,N_2535,N_1973);
or U5026 (N_5026,N_4997,N_4813);
nand U5027 (N_5027,N_3603,N_633);
nor U5028 (N_5028,N_2071,N_3460);
or U5029 (N_5029,N_3350,N_2182);
nand U5030 (N_5030,N_4135,N_1757);
and U5031 (N_5031,N_4572,N_455);
nor U5032 (N_5032,N_320,N_641);
or U5033 (N_5033,N_2138,N_2013);
nand U5034 (N_5034,N_727,N_2850);
nand U5035 (N_5035,N_4648,N_4259);
nor U5036 (N_5036,N_1975,N_4082);
xor U5037 (N_5037,N_315,N_3257);
or U5038 (N_5038,N_2172,N_3388);
nand U5039 (N_5039,N_3303,N_5);
nor U5040 (N_5040,N_851,N_3994);
and U5041 (N_5041,N_3579,N_2377);
nor U5042 (N_5042,N_1348,N_1768);
and U5043 (N_5043,N_2766,N_337);
nand U5044 (N_5044,N_4713,N_372);
nor U5045 (N_5045,N_1804,N_357);
nand U5046 (N_5046,N_4466,N_3915);
and U5047 (N_5047,N_2591,N_3041);
nand U5048 (N_5048,N_1476,N_2627);
and U5049 (N_5049,N_2163,N_2603);
nor U5050 (N_5050,N_2726,N_2883);
and U5051 (N_5051,N_2514,N_1577);
or U5052 (N_5052,N_3502,N_1152);
or U5053 (N_5053,N_4544,N_998);
or U5054 (N_5054,N_82,N_1257);
and U5055 (N_5055,N_2855,N_587);
nor U5056 (N_5056,N_1031,N_532);
nor U5057 (N_5057,N_278,N_338);
nand U5058 (N_5058,N_2137,N_2359);
nand U5059 (N_5059,N_1085,N_2911);
nor U5060 (N_5060,N_1049,N_2560);
and U5061 (N_5061,N_4957,N_940);
nand U5062 (N_5062,N_570,N_4991);
and U5063 (N_5063,N_4860,N_836);
or U5064 (N_5064,N_2236,N_2049);
or U5065 (N_5065,N_4881,N_1342);
and U5066 (N_5066,N_2081,N_2465);
nand U5067 (N_5067,N_3564,N_2544);
nor U5068 (N_5068,N_1738,N_1066);
or U5069 (N_5069,N_2792,N_508);
nor U5070 (N_5070,N_2130,N_872);
nor U5071 (N_5071,N_4041,N_1964);
or U5072 (N_5072,N_475,N_4439);
and U5073 (N_5073,N_1698,N_2413);
and U5074 (N_5074,N_2770,N_4543);
or U5075 (N_5075,N_3679,N_632);
nor U5076 (N_5076,N_3837,N_2993);
nor U5077 (N_5077,N_1167,N_1742);
nor U5078 (N_5078,N_4761,N_3540);
or U5079 (N_5079,N_2134,N_71);
nor U5080 (N_5080,N_4321,N_2853);
nor U5081 (N_5081,N_3080,N_3392);
nand U5082 (N_5082,N_4786,N_808);
or U5083 (N_5083,N_1276,N_2160);
nor U5084 (N_5084,N_4388,N_604);
nand U5085 (N_5085,N_1983,N_1337);
or U5086 (N_5086,N_885,N_2374);
or U5087 (N_5087,N_3656,N_3766);
nand U5088 (N_5088,N_3212,N_4229);
and U5089 (N_5089,N_3835,N_399);
or U5090 (N_5090,N_3071,N_1882);
or U5091 (N_5091,N_2292,N_1221);
nand U5092 (N_5092,N_2167,N_3744);
nand U5093 (N_5093,N_1314,N_299);
nor U5094 (N_5094,N_4252,N_3066);
or U5095 (N_5095,N_2011,N_4619);
and U5096 (N_5096,N_221,N_4281);
nor U5097 (N_5097,N_4473,N_3356);
or U5098 (N_5098,N_3498,N_2324);
or U5099 (N_5099,N_1640,N_683);
nor U5100 (N_5100,N_3861,N_4568);
nor U5101 (N_5101,N_3639,N_2450);
and U5102 (N_5102,N_3200,N_4093);
nor U5103 (N_5103,N_626,N_3007);
or U5104 (N_5104,N_4420,N_1797);
nor U5105 (N_5105,N_261,N_3364);
or U5106 (N_5106,N_4112,N_3209);
nand U5107 (N_5107,N_4682,N_3871);
nor U5108 (N_5108,N_4354,N_1562);
nor U5109 (N_5109,N_396,N_2237);
nor U5110 (N_5110,N_2382,N_2857);
or U5111 (N_5111,N_1029,N_4248);
nor U5112 (N_5112,N_2513,N_2610);
nor U5113 (N_5113,N_2987,N_692);
xor U5114 (N_5114,N_2454,N_3886);
nor U5115 (N_5115,N_2367,N_4254);
nor U5116 (N_5116,N_1790,N_582);
and U5117 (N_5117,N_4445,N_2039);
nand U5118 (N_5118,N_2538,N_311);
nand U5119 (N_5119,N_979,N_1542);
nand U5120 (N_5120,N_911,N_1649);
or U5121 (N_5121,N_2336,N_2949);
xnor U5122 (N_5122,N_3769,N_2676);
and U5123 (N_5123,N_680,N_4181);
or U5124 (N_5124,N_3346,N_3267);
or U5125 (N_5125,N_893,N_3841);
nand U5126 (N_5126,N_1767,N_964);
or U5127 (N_5127,N_1075,N_624);
and U5128 (N_5128,N_1264,N_2098);
nand U5129 (N_5129,N_2510,N_3668);
nand U5130 (N_5130,N_794,N_4821);
and U5131 (N_5131,N_4690,N_4455);
or U5132 (N_5132,N_1583,N_1635);
nor U5133 (N_5133,N_4605,N_4737);
nand U5134 (N_5134,N_2349,N_548);
or U5135 (N_5135,N_2278,N_3144);
nand U5136 (N_5136,N_2396,N_3555);
nor U5137 (N_5137,N_2418,N_1129);
and U5138 (N_5138,N_2781,N_1709);
or U5139 (N_5139,N_3607,N_4409);
or U5140 (N_5140,N_416,N_34);
xor U5141 (N_5141,N_1426,N_3439);
nand U5142 (N_5142,N_3796,N_620);
or U5143 (N_5143,N_3775,N_3486);
and U5144 (N_5144,N_4551,N_2147);
nor U5145 (N_5145,N_1752,N_3285);
nand U5146 (N_5146,N_3107,N_2555);
and U5147 (N_5147,N_4182,N_4674);
nor U5148 (N_5148,N_2506,N_3853);
nand U5149 (N_5149,N_4867,N_4747);
nand U5150 (N_5150,N_2588,N_3593);
nor U5151 (N_5151,N_2248,N_3405);
or U5152 (N_5152,N_4374,N_4644);
and U5153 (N_5153,N_4139,N_695);
nand U5154 (N_5154,N_287,N_3322);
or U5155 (N_5155,N_2372,N_317);
or U5156 (N_5156,N_816,N_3608);
xnor U5157 (N_5157,N_3811,N_3617);
and U5158 (N_5158,N_401,N_2932);
nor U5159 (N_5159,N_1101,N_371);
nand U5160 (N_5160,N_787,N_2233);
nand U5161 (N_5161,N_4693,N_1082);
and U5162 (N_5162,N_4552,N_186);
and U5163 (N_5163,N_4459,N_4197);
or U5164 (N_5164,N_168,N_833);
nand U5165 (N_5165,N_4649,N_671);
or U5166 (N_5166,N_4069,N_3123);
nand U5167 (N_5167,N_2635,N_1393);
or U5168 (N_5168,N_2992,N_2585);
nand U5169 (N_5169,N_4758,N_173);
nor U5170 (N_5170,N_3522,N_4148);
nor U5171 (N_5171,N_253,N_1070);
or U5172 (N_5172,N_3170,N_397);
nand U5173 (N_5173,N_1901,N_4107);
nand U5174 (N_5174,N_2780,N_1339);
or U5175 (N_5175,N_4656,N_656);
or U5176 (N_5176,N_453,N_557);
nor U5177 (N_5177,N_3445,N_2811);
and U5178 (N_5178,N_4958,N_1914);
or U5179 (N_5179,N_4576,N_3137);
nand U5180 (N_5180,N_4461,N_2456);
and U5181 (N_5181,N_1853,N_162);
and U5182 (N_5182,N_4438,N_1971);
nor U5183 (N_5183,N_3271,N_1412);
nand U5184 (N_5184,N_3753,N_2567);
or U5185 (N_5185,N_2773,N_1886);
or U5186 (N_5186,N_3273,N_730);
or U5187 (N_5187,N_2867,N_2864);
nand U5188 (N_5188,N_4683,N_646);
nor U5189 (N_5189,N_572,N_688);
nand U5190 (N_5190,N_1148,N_3951);
nor U5191 (N_5191,N_845,N_1364);
nand U5192 (N_5192,N_3810,N_1045);
or U5193 (N_5193,N_1730,N_3019);
nor U5194 (N_5194,N_2976,N_4011);
and U5195 (N_5195,N_3295,N_4634);
or U5196 (N_5196,N_1388,N_3403);
nand U5197 (N_5197,N_1528,N_1317);
nor U5198 (N_5198,N_625,N_163);
and U5199 (N_5199,N_3014,N_1127);
and U5200 (N_5200,N_2741,N_4852);
or U5201 (N_5201,N_1290,N_3044);
nor U5202 (N_5202,N_3677,N_2662);
and U5203 (N_5203,N_19,N_4650);
or U5204 (N_5204,N_677,N_2898);
nand U5205 (N_5205,N_2247,N_3021);
and U5206 (N_5206,N_2575,N_3050);
or U5207 (N_5207,N_481,N_3912);
nand U5208 (N_5208,N_3942,N_1704);
or U5209 (N_5209,N_1311,N_4978);
or U5210 (N_5210,N_3154,N_980);
nand U5211 (N_5211,N_1786,N_4692);
nor U5212 (N_5212,N_4386,N_4295);
nor U5213 (N_5213,N_342,N_4294);
or U5214 (N_5214,N_2159,N_4176);
nor U5215 (N_5215,N_159,N_1969);
or U5216 (N_5216,N_1865,N_4119);
nand U5217 (N_5217,N_4127,N_1042);
nor U5218 (N_5218,N_1970,N_2375);
nor U5219 (N_5219,N_3117,N_2965);
or U5220 (N_5220,N_1609,N_1193);
and U5221 (N_5221,N_3217,N_47);
nor U5222 (N_5222,N_202,N_2862);
nand U5223 (N_5223,N_2841,N_3230);
nand U5224 (N_5224,N_2542,N_2907);
nand U5225 (N_5225,N_2263,N_3268);
or U5226 (N_5226,N_4034,N_1647);
xor U5227 (N_5227,N_2649,N_1407);
nand U5228 (N_5228,N_4897,N_2813);
and U5229 (N_5229,N_3203,N_3497);
or U5230 (N_5230,N_1713,N_3110);
nor U5231 (N_5231,N_3449,N_1057);
nand U5232 (N_5232,N_2809,N_810);
nor U5233 (N_5233,N_1785,N_2938);
or U5234 (N_5234,N_757,N_900);
or U5235 (N_5235,N_2188,N_4444);
nor U5236 (N_5236,N_2577,N_2709);
and U5237 (N_5237,N_2045,N_3535);
or U5238 (N_5238,N_1479,N_4959);
nand U5239 (N_5239,N_2498,N_2020);
nand U5240 (N_5240,N_69,N_1215);
nand U5241 (N_5241,N_4789,N_4901);
nor U5242 (N_5242,N_4460,N_4186);
and U5243 (N_5243,N_4285,N_423);
or U5244 (N_5244,N_207,N_454);
and U5245 (N_5245,N_2435,N_3284);
and U5246 (N_5246,N_1714,N_4608);
nor U5247 (N_5247,N_855,N_1720);
or U5248 (N_5248,N_130,N_4701);
nor U5249 (N_5249,N_711,N_3708);
or U5250 (N_5250,N_3276,N_4952);
and U5251 (N_5251,N_1995,N_2275);
and U5252 (N_5252,N_92,N_4290);
nand U5253 (N_5253,N_4205,N_4984);
nor U5254 (N_5254,N_4508,N_4178);
or U5255 (N_5255,N_2810,N_1875);
and U5256 (N_5256,N_1623,N_3124);
or U5257 (N_5257,N_3638,N_4861);
and U5258 (N_5258,N_450,N_1416);
nand U5259 (N_5259,N_2330,N_725);
or U5260 (N_5260,N_3145,N_4055);
and U5261 (N_5261,N_2754,N_1222);
nand U5262 (N_5262,N_1778,N_4574);
nor U5263 (N_5263,N_3293,N_133);
or U5264 (N_5264,N_4160,N_3297);
and U5265 (N_5265,N_1135,N_1262);
or U5266 (N_5266,N_1324,N_3910);
nor U5267 (N_5267,N_2356,N_2141);
nand U5268 (N_5268,N_3888,N_2474);
nor U5269 (N_5269,N_3183,N_244);
and U5270 (N_5270,N_3771,N_4211);
nand U5271 (N_5271,N_555,N_594);
nand U5272 (N_5272,N_906,N_216);
nor U5273 (N_5273,N_4255,N_3770);
and U5274 (N_5274,N_1207,N_1689);
nor U5275 (N_5275,N_2623,N_3148);
nor U5276 (N_5276,N_3316,N_3527);
and U5277 (N_5277,N_2197,N_274);
nor U5278 (N_5278,N_1297,N_830);
nand U5279 (N_5279,N_942,N_1808);
nand U5280 (N_5280,N_4390,N_3948);
nand U5281 (N_5281,N_2281,N_3783);
nand U5282 (N_5282,N_2948,N_1253);
or U5283 (N_5283,N_4943,N_3214);
nand U5284 (N_5284,N_1958,N_4037);
nor U5285 (N_5285,N_1774,N_1715);
or U5286 (N_5286,N_4316,N_1077);
and U5287 (N_5287,N_689,N_3558);
nor U5288 (N_5288,N_3323,N_4021);
nor U5289 (N_5289,N_2040,N_3325);
nor U5290 (N_5290,N_3892,N_1357);
and U5291 (N_5291,N_1549,N_1770);
or U5292 (N_5292,N_2926,N_3611);
nand U5293 (N_5293,N_4450,N_2775);
nand U5294 (N_5294,N_1344,N_3831);
nor U5295 (N_5295,N_3626,N_1283);
and U5296 (N_5296,N_4829,N_543);
or U5297 (N_5297,N_1519,N_1481);
nor U5298 (N_5298,N_2398,N_1181);
and U5299 (N_5299,N_4724,N_180);
or U5300 (N_5300,N_869,N_779);
and U5301 (N_5301,N_2433,N_565);
and U5302 (N_5302,N_3950,N_2132);
and U5303 (N_5303,N_3778,N_4270);
or U5304 (N_5304,N_2845,N_2686);
nand U5305 (N_5305,N_1320,N_4537);
or U5306 (N_5306,N_4804,N_929);
or U5307 (N_5307,N_1304,N_1679);
nor U5308 (N_5308,N_3706,N_306);
and U5309 (N_5309,N_3413,N_4188);
nor U5310 (N_5310,N_3105,N_4357);
and U5311 (N_5311,N_369,N_1989);
nand U5312 (N_5312,N_3999,N_175);
nand U5313 (N_5313,N_440,N_431);
nand U5314 (N_5314,N_1932,N_694);
or U5315 (N_5315,N_4194,N_4451);
nand U5316 (N_5316,N_1722,N_3890);
or U5317 (N_5317,N_1037,N_3342);
and U5318 (N_5318,N_2713,N_1775);
and U5319 (N_5319,N_3559,N_3519);
nor U5320 (N_5320,N_3598,N_1369);
and U5321 (N_5321,N_662,N_2552);
nand U5322 (N_5322,N_789,N_2900);
and U5323 (N_5323,N_2699,N_1219);
nor U5324 (N_5324,N_404,N_4472);
or U5325 (N_5325,N_3962,N_1190);
or U5326 (N_5326,N_3795,N_831);
and U5327 (N_5327,N_3202,N_2483);
and U5328 (N_5328,N_430,N_266);
or U5329 (N_5329,N_4609,N_524);
nand U5330 (N_5330,N_1736,N_4371);
nor U5331 (N_5331,N_1558,N_1537);
xor U5332 (N_5332,N_3873,N_2540);
nand U5333 (N_5333,N_2208,N_922);
nor U5334 (N_5334,N_1773,N_284);
or U5335 (N_5335,N_2674,N_4585);
or U5336 (N_5336,N_2946,N_719);
and U5337 (N_5337,N_20,N_729);
or U5338 (N_5338,N_760,N_1180);
and U5339 (N_5339,N_2599,N_2164);
or U5340 (N_5340,N_4237,N_2616);
xnor U5341 (N_5341,N_3306,N_125);
and U5342 (N_5342,N_702,N_3340);
and U5343 (N_5343,N_2981,N_83);
or U5344 (N_5344,N_2534,N_4210);
nor U5345 (N_5345,N_4888,N_3520);
nor U5346 (N_5346,N_1404,N_1732);
or U5347 (N_5347,N_4129,N_4528);
nand U5348 (N_5348,N_3651,N_4350);
and U5349 (N_5349,N_3550,N_3554);
or U5350 (N_5350,N_21,N_255);
and U5351 (N_5351,N_2351,N_4571);
nand U5352 (N_5352,N_3462,N_3165);
nor U5353 (N_5353,N_4795,N_1899);
or U5354 (N_5354,N_3411,N_1483);
or U5355 (N_5355,N_3955,N_44);
nor U5356 (N_5356,N_923,N_2776);
nand U5357 (N_5357,N_4032,N_1579);
nor U5358 (N_5358,N_2466,N_4546);
or U5359 (N_5359,N_4039,N_3648);
nor U5360 (N_5360,N_2724,N_1918);
or U5361 (N_5361,N_2626,N_997);
nor U5362 (N_5362,N_31,N_275);
nand U5363 (N_5363,N_1189,N_4654);
nor U5364 (N_5364,N_1599,N_1735);
nor U5365 (N_5365,N_2690,N_3973);
and U5366 (N_5366,N_2111,N_2343);
nand U5367 (N_5367,N_1521,N_4727);
or U5368 (N_5368,N_2645,N_4926);
or U5369 (N_5369,N_746,N_2968);
nor U5370 (N_5370,N_682,N_4617);
nand U5371 (N_5371,N_4620,N_1218);
or U5372 (N_5372,N_4643,N_828);
nand U5373 (N_5373,N_788,N_2119);
or U5374 (N_5374,N_1398,N_290);
or U5375 (N_5375,N_1740,N_1420);
or U5376 (N_5376,N_2066,N_4723);
nor U5377 (N_5377,N_3553,N_4307);
nor U5378 (N_5378,N_2786,N_3157);
nand U5379 (N_5379,N_3664,N_3697);
or U5380 (N_5380,N_3587,N_2711);
nand U5381 (N_5381,N_4808,N_1118);
nor U5382 (N_5382,N_2607,N_3101);
or U5383 (N_5383,N_1503,N_4293);
and U5384 (N_5384,N_2858,N_4876);
or U5385 (N_5385,N_1810,N_1963);
nor U5386 (N_5386,N_4686,N_4048);
and U5387 (N_5387,N_884,N_4191);
or U5388 (N_5388,N_648,N_2608);
nor U5389 (N_5389,N_1150,N_1796);
nor U5390 (N_5390,N_4311,N_3485);
nand U5391 (N_5391,N_1897,N_4812);
or U5392 (N_5392,N_298,N_573);
or U5393 (N_5393,N_1798,N_4198);
and U5394 (N_5394,N_3365,N_151);
nor U5395 (N_5395,N_2458,N_4040);
nand U5396 (N_5396,N_3815,N_2403);
and U5397 (N_5397,N_1888,N_4224);
and U5398 (N_5398,N_1831,N_4873);
nor U5399 (N_5399,N_2999,N_2777);
or U5400 (N_5400,N_4655,N_1145);
or U5401 (N_5401,N_4116,N_4217);
nand U5402 (N_5402,N_3779,N_4763);
and U5403 (N_5403,N_3684,N_4028);
nor U5404 (N_5404,N_661,N_4563);
nor U5405 (N_5405,N_2918,N_1827);
nand U5406 (N_5406,N_1799,N_3000);
nor U5407 (N_5407,N_983,N_599);
and U5408 (N_5408,N_743,N_1096);
and U5409 (N_5409,N_4302,N_3072);
nor U5410 (N_5410,N_1915,N_1272);
or U5411 (N_5411,N_1889,N_2881);
and U5412 (N_5412,N_2428,N_4880);
nand U5413 (N_5413,N_2950,N_4657);
nand U5414 (N_5414,N_2913,N_4268);
nand U5415 (N_5415,N_2222,N_4060);
nor U5416 (N_5416,N_3175,N_3671);
or U5417 (N_5417,N_1660,N_4839);
xor U5418 (N_5418,N_3637,N_580);
nand U5419 (N_5419,N_2984,N_1325);
nor U5420 (N_5420,N_744,N_3862);
nand U5421 (N_5421,N_937,N_2235);
and U5422 (N_5422,N_3058,N_4258);
nor U5423 (N_5423,N_509,N_1992);
nand U5424 (N_5424,N_892,N_3454);
or U5425 (N_5425,N_1873,N_1541);
nand U5426 (N_5426,N_2667,N_478);
and U5427 (N_5427,N_2869,N_4320);
nor U5428 (N_5428,N_447,N_1333);
or U5429 (N_5429,N_1450,N_4338);
nor U5430 (N_5430,N_256,N_4018);
nand U5431 (N_5431,N_3623,N_4700);
or U5432 (N_5432,N_1004,N_4712);
and U5433 (N_5433,N_517,N_1198);
nand U5434 (N_5434,N_4641,N_1957);
nor U5435 (N_5435,N_1642,N_590);
nor U5436 (N_5436,N_2192,N_304);
xnor U5437 (N_5437,N_3083,N_4562);
or U5438 (N_5438,N_806,N_2824);
xor U5439 (N_5439,N_4714,N_3216);
and U5440 (N_5440,N_1507,N_56);
nand U5441 (N_5441,N_844,N_1972);
nor U5442 (N_5442,N_527,N_1216);
nor U5443 (N_5443,N_2847,N_419);
or U5444 (N_5444,N_992,N_3222);
and U5445 (N_5445,N_2389,N_4065);
nor U5446 (N_5446,N_1384,N_4798);
or U5447 (N_5447,N_3799,N_3560);
nand U5448 (N_5448,N_2405,N_3140);
and U5449 (N_5449,N_3930,N_2459);
nor U5450 (N_5450,N_1358,N_3224);
or U5451 (N_5451,N_316,N_2580);
nor U5452 (N_5452,N_2037,N_1377);
nand U5453 (N_5453,N_4257,N_1151);
nor U5454 (N_5454,N_1881,N_4553);
nor U5455 (N_5455,N_4499,N_2621);
nor U5456 (N_5456,N_4636,N_2395);
nand U5457 (N_5457,N_1811,N_1287);
or U5458 (N_5458,N_4587,N_2573);
nand U5459 (N_5459,N_1656,N_3337);
and U5460 (N_5460,N_4494,N_4317);
or U5461 (N_5461,N_4470,N_1254);
nand U5462 (N_5462,N_1187,N_4969);
nor U5463 (N_5463,N_1230,N_1690);
nor U5464 (N_5464,N_3855,N_1102);
or U5465 (N_5465,N_1605,N_3064);
or U5466 (N_5466,N_2095,N_90);
nand U5467 (N_5467,N_4043,N_373);
or U5468 (N_5468,N_2348,N_2022);
and U5469 (N_5469,N_387,N_2486);
nand U5470 (N_5470,N_1655,N_9);
nor U5471 (N_5471,N_2002,N_753);
or U5472 (N_5472,N_4569,N_2657);
xnor U5473 (N_5473,N_4748,N_1359);
and U5474 (N_5474,N_3479,N_801);
nand U5475 (N_5475,N_4331,N_3243);
and U5476 (N_5476,N_1636,N_2415);
nand U5477 (N_5477,N_4104,N_4687);
nand U5478 (N_5478,N_2682,N_668);
and U5479 (N_5479,N_1500,N_4756);
or U5480 (N_5480,N_4530,N_3722);
and U5481 (N_5481,N_3232,N_1097);
or U5482 (N_5482,N_3641,N_731);
or U5483 (N_5483,N_966,N_49);
or U5484 (N_5484,N_2581,N_1700);
and U5485 (N_5485,N_348,N_3009);
or U5486 (N_5486,N_2848,N_852);
nand U5487 (N_5487,N_2497,N_42);
and U5488 (N_5488,N_269,N_4419);
nor U5489 (N_5489,N_1858,N_3046);
nand U5490 (N_5490,N_4288,N_797);
or U5491 (N_5491,N_1301,N_3965);
or U5492 (N_5492,N_194,N_4796);
and U5493 (N_5493,N_3172,N_2205);
nand U5494 (N_5494,N_2963,N_4699);
nor U5495 (N_5495,N_4218,N_2661);
or U5496 (N_5496,N_1841,N_4545);
nor U5497 (N_5497,N_4326,N_3146);
nand U5498 (N_5498,N_4744,N_3191);
or U5499 (N_5499,N_3039,N_1456);
nand U5500 (N_5500,N_3678,N_2865);
nand U5501 (N_5501,N_879,N_696);
nor U5502 (N_5502,N_1249,N_2878);
or U5503 (N_5503,N_4204,N_4230);
or U5504 (N_5504,N_2658,N_4799);
nor U5505 (N_5505,N_4379,N_217);
nand U5506 (N_5506,N_2378,N_1361);
nand U5507 (N_5507,N_3451,N_907);
or U5508 (N_5508,N_972,N_4970);
nand U5509 (N_5509,N_3086,N_4790);
and U5510 (N_5510,N_2957,N_2408);
or U5511 (N_5511,N_1996,N_2624);
nand U5512 (N_5512,N_1133,N_1039);
nand U5513 (N_5513,N_874,N_3278);
nor U5514 (N_5514,N_3301,N_127);
or U5515 (N_5515,N_977,N_2902);
nor U5516 (N_5516,N_790,N_1073);
and U5517 (N_5517,N_4904,N_1560);
nor U5518 (N_5518,N_4823,N_4187);
and U5519 (N_5519,N_4730,N_3468);
and U5520 (N_5520,N_2305,N_1044);
or U5521 (N_5521,N_4029,N_25);
or U5522 (N_5522,N_301,N_364);
or U5523 (N_5523,N_1782,N_2082);
and U5524 (N_5524,N_3991,N_2301);
and U5525 (N_5525,N_4355,N_1179);
nand U5526 (N_5526,N_4785,N_3343);
nor U5527 (N_5527,N_1123,N_3528);
nand U5528 (N_5528,N_2941,N_4073);
and U5529 (N_5529,N_2669,N_2106);
or U5530 (N_5530,N_1863,N_3731);
nand U5531 (N_5531,N_2333,N_3493);
or U5532 (N_5532,N_2671,N_927);
nand U5533 (N_5533,N_2894,N_4076);
or U5534 (N_5534,N_2750,N_307);
nor U5535 (N_5535,N_4673,N_2196);
or U5536 (N_5536,N_2590,N_1243);
and U5537 (N_5537,N_2030,N_1203);
and U5538 (N_5538,N_1171,N_469);
nand U5539 (N_5539,N_409,N_2572);
nand U5540 (N_5540,N_1511,N_3488);
nor U5541 (N_5541,N_2551,N_826);
nand U5542 (N_5542,N_1210,N_1505);
nor U5543 (N_5543,N_2480,N_2710);
nand U5544 (N_5544,N_4953,N_411);
or U5545 (N_5545,N_4577,N_2150);
or U5546 (N_5546,N_4359,N_29);
nor U5547 (N_5547,N_4990,N_1725);
nor U5548 (N_5548,N_1,N_2527);
or U5549 (N_5549,N_1451,N_994);
nor U5550 (N_5550,N_4579,N_1229);
and U5551 (N_5551,N_3317,N_4754);
or U5552 (N_5552,N_4023,N_2730);
nor U5553 (N_5553,N_2092,N_1170);
or U5554 (N_5554,N_856,N_3534);
or U5555 (N_5555,N_3457,N_468);
nand U5556 (N_5556,N_282,N_205);
nand U5557 (N_5557,N_1463,N_3859);
and U5558 (N_5558,N_947,N_827);
and U5559 (N_5559,N_2118,N_4529);
nand U5560 (N_5560,N_2241,N_2287);
nor U5561 (N_5561,N_1477,N_2121);
nor U5562 (N_5562,N_3218,N_982);
and U5563 (N_5563,N_3151,N_35);
nand U5564 (N_5564,N_4309,N_40);
or U5565 (N_5565,N_3673,N_45);
and U5566 (N_5566,N_3875,N_4342);
nand U5567 (N_5567,N_3932,N_499);
or U5568 (N_5568,N_8,N_3026);
nand U5569 (N_5569,N_4911,N_4598);
nand U5570 (N_5570,N_4866,N_538);
nor U5571 (N_5571,N_2371,N_2489);
nand U5572 (N_5572,N_358,N_1663);
xnor U5573 (N_5573,N_4006,N_4411);
and U5574 (N_5574,N_456,N_4105);
and U5575 (N_5575,N_1731,N_2908);
nand U5576 (N_5576,N_2899,N_3483);
or U5577 (N_5577,N_3945,N_4910);
and U5578 (N_5578,N_4675,N_4014);
nand U5579 (N_5579,N_800,N_1007);
or U5580 (N_5580,N_1631,N_3867);
and U5581 (N_5581,N_3287,N_798);
or U5582 (N_5582,N_3686,N_142);
and U5583 (N_5583,N_791,N_4109);
nor U5584 (N_5584,N_700,N_4540);
or U5585 (N_5585,N_3088,N_3081);
xnor U5586 (N_5586,N_3023,N_507);
or U5587 (N_5587,N_1898,N_1188);
or U5588 (N_5588,N_1685,N_1499);
nor U5589 (N_5589,N_1072,N_2617);
nand U5590 (N_5590,N_4130,N_1514);
or U5591 (N_5591,N_4865,N_3043);
nand U5592 (N_5592,N_1332,N_1495);
nor U5593 (N_5593,N_3984,N_4017);
nor U5594 (N_5594,N_4312,N_3128);
and U5595 (N_5595,N_13,N_1356);
nand U5596 (N_5596,N_4125,N_1502);
or U5597 (N_5597,N_2909,N_591);
and U5598 (N_5598,N_1403,N_4183);
nor U5599 (N_5599,N_4512,N_152);
and U5600 (N_5600,N_4117,N_4142);
nor U5601 (N_5601,N_1637,N_374);
and U5602 (N_5602,N_4304,N_2436);
nand U5603 (N_5603,N_750,N_3850);
nand U5604 (N_5604,N_2743,N_2229);
or U5605 (N_5605,N_1251,N_770);
nand U5606 (N_5606,N_4004,N_1803);
and U5607 (N_5607,N_2615,N_3767);
nand U5608 (N_5608,N_4986,N_1292);
nand U5609 (N_5609,N_3416,N_1658);
nand U5610 (N_5610,N_426,N_3180);
and U5611 (N_5611,N_1936,N_3756);
or U5612 (N_5612,N_3310,N_4265);
or U5613 (N_5613,N_3969,N_1509);
nor U5614 (N_5614,N_2860,N_3567);
or U5615 (N_5615,N_3448,N_3698);
and U5616 (N_5616,N_418,N_3688);
or U5617 (N_5617,N_1868,N_3477);
or U5618 (N_5618,N_4013,N_2288);
xor U5619 (N_5619,N_549,N_171);
and U5620 (N_5620,N_1061,N_2818);
nor U5621 (N_5621,N_3078,N_4835);
nand U5622 (N_5622,N_2888,N_3882);
and U5623 (N_5623,N_4378,N_3198);
and U5624 (N_5624,N_4666,N_184);
nor U5625 (N_5625,N_1506,N_1454);
nor U5626 (N_5626,N_2820,N_1184);
and U5627 (N_5627,N_368,N_3139);
and U5628 (N_5628,N_4633,N_601);
nand U5629 (N_5629,N_4877,N_4822);
nand U5630 (N_5630,N_2072,N_4516);
nand U5631 (N_5631,N_3463,N_3800);
nor U5632 (N_5632,N_2757,N_1680);
nand U5633 (N_5633,N_3329,N_1792);
and U5634 (N_5634,N_119,N_4846);
nor U5635 (N_5635,N_3309,N_2733);
and U5636 (N_5636,N_2499,N_684);
or U5637 (N_5637,N_3712,N_2554);
or U5638 (N_5638,N_3111,N_4679);
nand U5639 (N_5639,N_276,N_533);
and U5640 (N_5640,N_3279,N_4965);
nand U5641 (N_5641,N_460,N_488);
nor U5642 (N_5642,N_4456,N_752);
nand U5643 (N_5643,N_767,N_2720);
nand U5644 (N_5644,N_4383,N_1224);
and U5645 (N_5645,N_2975,N_782);
nor U5646 (N_5646,N_1026,N_1744);
and U5647 (N_5647,N_3065,N_1575);
and U5648 (N_5648,N_424,N_451);
and U5649 (N_5649,N_2019,N_3536);
nor U5650 (N_5650,N_2209,N_4502);
and U5651 (N_5651,N_4449,N_2655);
nor U5652 (N_5652,N_835,N_2634);
nor U5653 (N_5653,N_4361,N_987);
xor U5654 (N_5654,N_129,N_3647);
nand U5655 (N_5655,N_1413,N_390);
and U5656 (N_5656,N_4826,N_4898);
or U5657 (N_5657,N_4800,N_537);
or U5658 (N_5658,N_873,N_3851);
nand U5659 (N_5659,N_502,N_2728);
nand U5660 (N_5660,N_354,N_635);
or U5661 (N_5661,N_717,N_1529);
nor U5662 (N_5662,N_4567,N_969);
and U5663 (N_5663,N_1270,N_3791);
nand U5664 (N_5664,N_3314,N_2745);
nor U5665 (N_5665,N_2628,N_902);
nor U5666 (N_5666,N_3825,N_813);
and U5667 (N_5667,N_859,N_639);
nand U5668 (N_5668,N_3369,N_1269);
and U5669 (N_5669,N_1727,N_4066);
and U5670 (N_5670,N_3982,N_2831);
or U5671 (N_5671,N_286,N_3265);
xor U5672 (N_5672,N_39,N_3037);
nor U5673 (N_5673,N_3521,N_3153);
nand U5674 (N_5674,N_1789,N_3235);
nand U5675 (N_5675,N_1385,N_3619);
or U5676 (N_5676,N_531,N_3409);
nor U5677 (N_5677,N_3395,N_332);
nor U5678 (N_5678,N_675,N_4559);
and U5679 (N_5679,N_4190,N_64);
nor U5680 (N_5680,N_4720,N_3420);
or U5681 (N_5681,N_2226,N_2771);
nor U5682 (N_5682,N_3508,N_1427);
nand U5683 (N_5683,N_1830,N_3562);
nand U5684 (N_5684,N_3625,N_3348);
or U5685 (N_5685,N_3042,N_109);
nor U5686 (N_5686,N_4031,N_461);
nand U5687 (N_5687,N_3121,N_622);
or U5688 (N_5688,N_948,N_2493);
nor U5689 (N_5689,N_1567,N_4090);
nor U5690 (N_5690,N_2007,N_2856);
and U5691 (N_5691,N_406,N_512);
nor U5692 (N_5692,N_4964,N_3500);
and U5693 (N_5693,N_3162,N_4161);
nand U5694 (N_5694,N_408,N_2939);
and U5695 (N_5695,N_1445,N_1137);
nor U5696 (N_5696,N_4653,N_473);
nor U5697 (N_5697,N_4740,N_4356);
xor U5698 (N_5698,N_2595,N_2064);
and U5699 (N_5699,N_2816,N_636);
nand U5700 (N_5700,N_3277,N_4431);
and U5701 (N_5701,N_4858,N_4526);
or U5702 (N_5702,N_501,N_3570);
or U5703 (N_5703,N_1688,N_3242);
or U5704 (N_5704,N_2723,N_4110);
and U5705 (N_5705,N_1781,N_3824);
and U5706 (N_5706,N_4838,N_3926);
nor U5707 (N_5707,N_2562,N_1568);
nor U5708 (N_5708,N_4478,N_3548);
nand U5709 (N_5709,N_2310,N_825);
nand U5710 (N_5710,N_3970,N_4946);
and U5711 (N_5711,N_2169,N_3763);
or U5712 (N_5712,N_1316,N_2417);
xor U5713 (N_5713,N_181,N_3048);
nor U5714 (N_5714,N_4940,N_628);
or U5715 (N_5715,N_3379,N_3499);
or U5716 (N_5716,N_1443,N_1000);
nor U5717 (N_5717,N_1517,N_2206);
nand U5718 (N_5718,N_1092,N_2046);
nor U5719 (N_5719,N_1435,N_2755);
nand U5720 (N_5720,N_4195,N_1076);
or U5721 (N_5721,N_1728,N_1662);
or U5722 (N_5722,N_4751,N_4932);
nand U5723 (N_5723,N_2473,N_3115);
or U5724 (N_5724,N_3856,N_3130);
nand U5725 (N_5725,N_2947,N_3675);
nand U5726 (N_5726,N_3367,N_2133);
and U5727 (N_5727,N_263,N_3613);
and U5728 (N_5728,N_2265,N_3027);
xor U5729 (N_5729,N_3572,N_4413);
nand U5730 (N_5730,N_3734,N_452);
nor U5731 (N_5731,N_3354,N_3581);
nand U5732 (N_5732,N_1162,N_3906);
nand U5733 (N_5733,N_3254,N_3985);
nand U5734 (N_5734,N_849,N_2556);
and U5735 (N_5735,N_1233,N_2484);
nand U5736 (N_5736,N_2570,N_3787);
and U5737 (N_5737,N_1908,N_3432);
and U5738 (N_5738,N_237,N_1139);
xnor U5739 (N_5739,N_349,N_3474);
and U5740 (N_5740,N_4928,N_1331);
nor U5741 (N_5741,N_1465,N_1372);
and U5742 (N_5742,N_3788,N_803);
and U5743 (N_5743,N_1111,N_4177);
or U5744 (N_5744,N_2569,N_1997);
or U5745 (N_5745,N_3255,N_4707);
nand U5746 (N_5746,N_1273,N_1200);
or U5747 (N_5747,N_2479,N_3120);
nor U5748 (N_5748,N_3427,N_2221);
nor U5749 (N_5749,N_723,N_1191);
nand U5750 (N_5750,N_1832,N_3312);
nand U5751 (N_5751,N_3082,N_4582);
or U5752 (N_5752,N_2732,N_2673);
nand U5753 (N_5753,N_4418,N_2342);
or U5754 (N_5754,N_579,N_3236);
and U5755 (N_5755,N_4871,N_4328);
and U5756 (N_5756,N_4635,N_4847);
nor U5757 (N_5757,N_2619,N_560);
nor U5758 (N_5758,N_1462,N_3748);
nor U5759 (N_5759,N_3672,N_3126);
nor U5760 (N_5760,N_3693,N_3911);
nor U5761 (N_5761,N_2611,N_793);
and U5762 (N_5762,N_4251,N_773);
and U5763 (N_5763,N_498,N_1105);
nor U5764 (N_5764,N_4137,N_961);
and U5765 (N_5765,N_2689,N_2402);
or U5766 (N_5766,N_3011,N_4890);
nand U5767 (N_5767,N_759,N_3620);
nand U5768 (N_5768,N_3854,N_2763);
nand U5769 (N_5769,N_3434,N_1355);
nand U5770 (N_5770,N_4094,N_4005);
or U5771 (N_5771,N_70,N_4708);
nand U5772 (N_5772,N_4496,N_2298);
nor U5773 (N_5773,N_3685,N_3681);
nand U5774 (N_5774,N_3138,N_1981);
nor U5775 (N_5775,N_3506,N_4891);
nand U5776 (N_5776,N_4919,N_933);
or U5777 (N_5777,N_2691,N_2601);
or U5778 (N_5778,N_1482,N_3390);
nor U5779 (N_5779,N_1121,N_429);
or U5780 (N_5780,N_574,N_4733);
nand U5781 (N_5781,N_3661,N_2996);
and U5782 (N_5782,N_341,N_3702);
nor U5783 (N_5783,N_3935,N_3975);
nor U5784 (N_5784,N_1448,N_1192);
and U5785 (N_5785,N_3490,N_3341);
nor U5786 (N_5786,N_2681,N_755);
nand U5787 (N_5787,N_2680,N_520);
or U5788 (N_5788,N_4256,N_3933);
nor U5789 (N_5789,N_63,N_4671);
and U5790 (N_5790,N_655,N_3517);
nand U5791 (N_5791,N_2937,N_2803);
nand U5792 (N_5792,N_2024,N_3917);
nor U5793 (N_5793,N_1182,N_271);
nand U5794 (N_5794,N_1795,N_3399);
nor U5795 (N_5795,N_1467,N_4979);
and U5796 (N_5796,N_139,N_709);
nor U5797 (N_5797,N_2747,N_183);
nor U5798 (N_5798,N_3921,N_3262);
nand U5799 (N_5799,N_4096,N_2990);
nand U5800 (N_5800,N_909,N_2953);
nand U5801 (N_5801,N_4219,N_2067);
nand U5802 (N_5802,N_2496,N_1874);
and U5803 (N_5803,N_62,N_4400);
or U5804 (N_5804,N_443,N_384);
nand U5805 (N_5805,N_904,N_3624);
nor U5806 (N_5806,N_978,N_4141);
or U5807 (N_5807,N_4539,N_1919);
and U5808 (N_5808,N_3010,N_886);
and U5809 (N_5809,N_2276,N_1110);
nand U5810 (N_5810,N_2653,N_3429);
nor U5811 (N_5811,N_3036,N_563);
or U5812 (N_5812,N_4533,N_3876);
nor U5813 (N_5813,N_3832,N_3458);
and U5814 (N_5814,N_4053,N_1472);
and U5815 (N_5815,N_734,N_2231);
and U5816 (N_5816,N_386,N_4664);
nor U5817 (N_5817,N_1389,N_1048);
or U5818 (N_5818,N_1693,N_2912);
and U5819 (N_5819,N_4081,N_4353);
nor U5820 (N_5820,N_2602,N_365);
and U5821 (N_5821,N_2694,N_1158);
nand U5822 (N_5822,N_4166,N_722);
and U5823 (N_5823,N_229,N_3430);
nor U5824 (N_5824,N_500,N_1522);
nand U5825 (N_5825,N_4487,N_778);
nor U5826 (N_5826,N_1366,N_4676);
nor U5827 (N_5827,N_314,N_3571);
and U5828 (N_5828,N_1800,N_616);
nand U5829 (N_5829,N_4917,N_762);
nand U5830 (N_5830,N_2906,N_4063);
or U5831 (N_5831,N_1668,N_1933);
nor U5832 (N_5832,N_1006,N_12);
and U5833 (N_5833,N_4920,N_351);
nand U5834 (N_5834,N_3440,N_3400);
nand U5835 (N_5835,N_1539,N_1760);
and U5836 (N_5836,N_1571,N_2416);
or U5837 (N_5837,N_4044,N_1852);
or U5838 (N_5838,N_2814,N_4154);
or U5839 (N_5839,N_2721,N_3849);
or U5840 (N_5840,N_2260,N_1436);
nand U5841 (N_5841,N_3417,N_2337);
nand U5842 (N_5842,N_4098,N_2751);
or U5843 (N_5843,N_4403,N_4557);
or U5844 (N_5844,N_2054,N_4375);
or U5845 (N_5845,N_4101,N_113);
or U5846 (N_5846,N_2517,N_839);
nand U5847 (N_5847,N_3765,N_343);
or U5848 (N_5848,N_4067,N_24);
nand U5849 (N_5849,N_72,N_2446);
or U5850 (N_5850,N_3059,N_2297);
nand U5851 (N_5851,N_4351,N_3104);
and U5852 (N_5852,N_2835,N_3883);
nand U5853 (N_5853,N_2523,N_3270);
nand U5854 (N_5854,N_4232,N_4003);
nor U5855 (N_5855,N_2269,N_882);
or U5856 (N_5856,N_550,N_3239);
nand U5857 (N_5857,N_38,N_2700);
nand U5858 (N_5858,N_1588,N_3290);
nor U5859 (N_5859,N_2441,N_2335);
nand U5860 (N_5860,N_3455,N_3627);
or U5861 (N_5861,N_1323,N_2325);
nor U5862 (N_5862,N_2460,N_1570);
nand U5863 (N_5863,N_2284,N_3334);
and U5864 (N_5864,N_4108,N_80);
or U5865 (N_5865,N_4358,N_597);
nor U5866 (N_5866,N_4469,N_4234);
or U5867 (N_5867,N_2285,N_1673);
and U5868 (N_5868,N_11,N_2890);
or U5869 (N_5869,N_1982,N_3464);
or U5870 (N_5870,N_4074,N_3974);
nor U5871 (N_5871,N_1783,N_2528);
and U5872 (N_5872,N_1950,N_1589);
or U5873 (N_5873,N_3155,N_1909);
nand U5874 (N_5874,N_2419,N_190);
and U5875 (N_5875,N_1460,N_3067);
nor U5876 (N_5876,N_1845,N_2452);
nor U5877 (N_5877,N_17,N_672);
nand U5878 (N_5878,N_391,N_1153);
or U5879 (N_5879,N_67,N_4875);
or U5880 (N_5880,N_812,N_792);
or U5881 (N_5881,N_589,N_1433);
or U5882 (N_5882,N_3537,N_1769);
nand U5883 (N_5883,N_3809,N_1402);
nor U5884 (N_5884,N_676,N_4261);
nand U5885 (N_5885,N_2805,N_4291);
nor U5886 (N_5886,N_3299,N_603);
and U5887 (N_5887,N_3952,N_167);
and U5888 (N_5888,N_4276,N_4019);
and U5889 (N_5889,N_1611,N_2453);
nand U5890 (N_5890,N_593,N_2886);
nand U5891 (N_5891,N_4627,N_3908);
or U5892 (N_5892,N_1968,N_1653);
nand U5893 (N_5893,N_883,N_1846);
and U5894 (N_5894,N_4441,N_2181);
or U5895 (N_5895,N_3142,N_1392);
and U5896 (N_5896,N_596,N_4133);
nand U5897 (N_5897,N_973,N_4344);
nor U5898 (N_5898,N_3714,N_1205);
nor U5899 (N_5899,N_4764,N_710);
nand U5900 (N_5900,N_619,N_3251);
nor U5901 (N_5901,N_3786,N_4238);
nor U5902 (N_5902,N_3237,N_742);
and U5903 (N_5903,N_1354,N_2849);
and U5904 (N_5904,N_2885,N_4414);
nor U5905 (N_5905,N_3947,N_4807);
nand U5906 (N_5906,N_1527,N_1136);
nor U5907 (N_5907,N_2062,N_4404);
or U5908 (N_5908,N_3256,N_3738);
and U5909 (N_5909,N_3609,N_2074);
and U5910 (N_5910,N_1306,N_658);
and U5911 (N_5911,N_545,N_3670);
or U5912 (N_5912,N_2110,N_2744);
nand U5913 (N_5913,N_2982,N_4842);
nor U5914 (N_5914,N_1536,N_4089);
nor U5915 (N_5915,N_1629,N_4440);
and U5916 (N_5916,N_170,N_4365);
nor U5917 (N_5917,N_3382,N_3865);
nand U5918 (N_5918,N_2283,N_1703);
nor U5919 (N_5919,N_3531,N_3163);
and U5920 (N_5920,N_2195,N_4515);
nor U5921 (N_5921,N_3260,N_1754);
and U5922 (N_5922,N_1058,N_2704);
and U5923 (N_5923,N_2096,N_1286);
nand U5924 (N_5924,N_3781,N_741);
nand U5925 (N_5925,N_215,N_4239);
nor U5926 (N_5926,N_880,N_4925);
or U5927 (N_5927,N_1346,N_1002);
and U5928 (N_5928,N_1440,N_427);
nor U5929 (N_5929,N_4282,N_4850);
or U5930 (N_5930,N_2340,N_2268);
nor U5931 (N_5931,N_375,N_4841);
nor U5932 (N_5932,N_240,N_1924);
nor U5933 (N_5933,N_3879,N_1592);
nor U5934 (N_5934,N_123,N_4012);
nor U5935 (N_5935,N_2097,N_3507);
or U5936 (N_5936,N_1606,N_4169);
nor U5937 (N_5937,N_2184,N_3798);
nor U5938 (N_5938,N_2085,N_2327);
nand U5939 (N_5939,N_1144,N_330);
and U5940 (N_5940,N_323,N_2687);
nor U5941 (N_5941,N_3207,N_2175);
nand U5942 (N_5942,N_1766,N_4468);
nand U5943 (N_5943,N_2178,N_1177);
and U5944 (N_5944,N_4446,N_637);
or U5945 (N_5945,N_2495,N_3492);
nor U5946 (N_5946,N_1156,N_2316);
or U5947 (N_5947,N_615,N_2782);
nor U5948 (N_5948,N_2756,N_3713);
nand U5949 (N_5949,N_2749,N_712);
nor U5950 (N_5950,N_4595,N_1523);
or U5951 (N_5951,N_1422,N_2696);
nand U5952 (N_5952,N_748,N_2875);
or U5953 (N_5953,N_135,N_1296);
and U5954 (N_5954,N_3726,N_3355);
nor U5955 (N_5955,N_4646,N_2411);
and U5956 (N_5956,N_4336,N_595);
nor U5957 (N_5957,N_4271,N_2931);
or U5958 (N_5958,N_1459,N_1594);
nand U5959 (N_5959,N_820,N_1343);
xor U5960 (N_5960,N_1293,N_2431);
xor U5961 (N_5961,N_2334,N_1379);
and U5962 (N_5962,N_2594,N_1282);
nor U5963 (N_5963,N_1812,N_2300);
or U5964 (N_5964,N_2870,N_2804);
or U5965 (N_5965,N_1014,N_2978);
or U5966 (N_5966,N_728,N_1603);
or U5967 (N_5967,N_1471,N_2381);
nand U5968 (N_5968,N_3189,N_3653);
or U5969 (N_5969,N_2507,N_3660);
nand U5970 (N_5970,N_1993,N_4745);
or U5971 (N_5971,N_4463,N_1441);
and U5972 (N_5972,N_2187,N_2541);
nor U5973 (N_5973,N_310,N_536);
nor U5974 (N_5974,N_3085,N_2578);
nand U5975 (N_5975,N_4163,N_1475);
or U5976 (N_5976,N_4769,N_4193);
nor U5977 (N_5977,N_3079,N_2564);
and U5978 (N_5978,N_346,N_3227);
nor U5979 (N_5979,N_1326,N_1809);
nand U5980 (N_5980,N_1737,N_569);
nand U5981 (N_5981,N_1621,N_2469);
nor U5982 (N_5982,N_1093,N_985);
or U5983 (N_5983,N_3838,N_2942);
nor U5984 (N_5984,N_4289,N_272);
and U5985 (N_5985,N_850,N_1584);
nor U5986 (N_5986,N_4902,N_432);
nor U5987 (N_5987,N_4752,N_3169);
and U5988 (N_5988,N_2970,N_1408);
and U5989 (N_5989,N_1596,N_4367);
nor U5990 (N_5990,N_4532,N_585);
nand U5991 (N_5991,N_340,N_1305);
and U5992 (N_5992,N_2308,N_614);
nand U5993 (N_5993,N_2522,N_4848);
nand U5994 (N_5994,N_2212,N_3075);
or U5995 (N_5995,N_2960,N_4274);
nand U5996 (N_5996,N_3344,N_3219);
or U5997 (N_5997,N_1298,N_3667);
nand U5998 (N_5998,N_283,N_3176);
and U5999 (N_5999,N_4616,N_4330);
or U6000 (N_6000,N_1322,N_3053);
or U6001 (N_6001,N_4410,N_3363);
and U6002 (N_6002,N_2376,N_1235);
nor U6003 (N_6003,N_3074,N_4284);
or U6004 (N_6004,N_939,N_3665);
nor U6005 (N_6005,N_2463,N_436);
nor U6006 (N_6006,N_402,N_4201);
or U6007 (N_6007,N_4717,N_4721);
nor U6008 (N_6008,N_2394,N_2077);
and U6009 (N_6009,N_4849,N_4147);
and U6010 (N_6010,N_721,N_4206);
and U6011 (N_6011,N_3990,N_959);
or U6012 (N_6012,N_2306,N_1244);
nand U6013 (N_6013,N_4263,N_389);
and U6014 (N_6014,N_3473,N_2478);
or U6015 (N_6015,N_4437,N_949);
nor U6016 (N_6016,N_1266,N_1319);
nor U6017 (N_6017,N_4392,N_3511);
nor U6018 (N_6018,N_3378,N_3467);
nand U6019 (N_6019,N_1676,N_356);
nor U6020 (N_6020,N_4828,N_3264);
nor U6021 (N_6021,N_4642,N_4068);
and U6022 (N_6022,N_1033,N_3015);
and U6023 (N_6023,N_4493,N_176);
nor U6024 (N_6024,N_2105,N_4794);
nor U6025 (N_6025,N_1741,N_4554);
nor U6026 (N_6026,N_4915,N_575);
and U6027 (N_6027,N_1473,N_2261);
nor U6028 (N_6028,N_2242,N_417);
and U6029 (N_6029,N_318,N_3826);
nor U6030 (N_6030,N_2738,N_2023);
and U6031 (N_6031,N_3742,N_1213);
and U6032 (N_6032,N_2793,N_2027);
or U6033 (N_6033,N_3359,N_2998);
or U6034 (N_6034,N_4373,N_4615);
or U6035 (N_6035,N_3319,N_4347);
nor U6036 (N_6036,N_3289,N_740);
nand U6037 (N_6037,N_1163,N_2383);
or U6038 (N_6038,N_122,N_4924);
or U6039 (N_6039,N_2086,N_4672);
and U6040 (N_6040,N_3983,N_2044);
or U6041 (N_6041,N_4222,N_3149);
and U6042 (N_6042,N_1710,N_3171);
nand U6043 (N_6043,N_2083,N_3094);
nand U6044 (N_6044,N_2323,N_1911);
nand U6045 (N_6045,N_4960,N_3201);
nor U6046 (N_6046,N_4453,N_4146);
nor U6047 (N_6047,N_871,N_4504);
nand U6048 (N_6048,N_4909,N_1559);
nand U6049 (N_6049,N_1652,N_1634);
nand U6050 (N_6050,N_765,N_2967);
and U6051 (N_6051,N_2219,N_4912);
or U6052 (N_6052,N_3961,N_2220);
nor U6053 (N_6053,N_976,N_2951);
nor U6054 (N_6054,N_558,N_523);
or U6055 (N_6055,N_4010,N_3247);
or U6056 (N_6056,N_2807,N_1212);
nor U6057 (N_6057,N_4513,N_2505);
nand U6058 (N_6058,N_3398,N_1607);
and U6059 (N_6059,N_1194,N_4534);
nand U6060 (N_6060,N_3307,N_1258);
nand U6061 (N_6061,N_2329,N_4235);
and U6062 (N_6062,N_2830,N_4784);
nor U6063 (N_6063,N_761,N_3311);
and U6064 (N_6064,N_777,N_2515);
and U6065 (N_6065,N_425,N_2051);
nor U6066 (N_6066,N_1890,N_738);
nand U6067 (N_6067,N_3541,N_1423);
or U6068 (N_6068,N_4026,N_3631);
nor U6069 (N_6069,N_1894,N_2005);
nand U6070 (N_6070,N_1185,N_4519);
nand U6071 (N_6071,N_1234,N_465);
nand U6072 (N_6072,N_1387,N_2518);
nand U6073 (N_6073,N_4339,N_367);
and U6074 (N_6074,N_225,N_4333);
and U6075 (N_6075,N_2642,N_4592);
nor U6076 (N_6076,N_1532,N_4038);
nor U6077 (N_6077,N_4998,N_3489);
and U6078 (N_6078,N_1925,N_3730);
and U6079 (N_6079,N_2904,N_4522);
or U6080 (N_6080,N_2360,N_3895);
or U6081 (N_6081,N_1712,N_4827);
and U6082 (N_6082,N_4524,N_4085);
and U6083 (N_6083,N_3127,N_2656);
nand U6084 (N_6084,N_4308,N_1247);
nand U6085 (N_6085,N_1036,N_3335);
and U6086 (N_6086,N_2705,N_106);
and U6087 (N_6087,N_2238,N_497);
and U6088 (N_6088,N_4996,N_1554);
nand U6089 (N_6089,N_1368,N_3780);
nand U6090 (N_6090,N_3360,N_1892);
and U6091 (N_6091,N_4766,N_4227);
or U6092 (N_6092,N_3286,N_1374);
nor U6093 (N_6093,N_3470,N_2125);
nor U6094 (N_6094,N_3621,N_3655);
nand U6095 (N_6095,N_4366,N_124);
or U6096 (N_6096,N_1161,N_3391);
or U6097 (N_6097,N_4243,N_353);
and U6098 (N_6098,N_496,N_3056);
nand U6099 (N_6099,N_1094,N_3001);
and U6100 (N_6100,N_3112,N_4640);
nand U6101 (N_6101,N_3784,N_3816);
nand U6102 (N_6102,N_30,N_1818);
or U6103 (N_6103,N_2618,N_3339);
nand U6104 (N_6104,N_3676,N_4879);
nor U6105 (N_6105,N_196,N_2409);
or U6106 (N_6106,N_3633,N_1217);
and U6107 (N_6107,N_3351,N_472);
nand U6108 (N_6108,N_3496,N_4610);
and U6109 (N_6109,N_3551,N_4782);
or U6110 (N_6110,N_265,N_3931);
or U6111 (N_6111,N_3749,N_1484);
and U6112 (N_6112,N_780,N_4088);
nor U6113 (N_6113,N_4523,N_1686);
nor U6114 (N_6114,N_3381,N_4868);
nor U6115 (N_6115,N_4853,N_4059);
and U6116 (N_6116,N_2587,N_3476);
nand U6117 (N_6117,N_2769,N_1501);
nor U6118 (N_6118,N_2146,N_3320);
or U6119 (N_6119,N_2001,N_1871);
or U6120 (N_6120,N_4626,N_1526);
nor U6121 (N_6121,N_1370,N_1492);
and U6122 (N_6122,N_4296,N_4025);
and U6123 (N_6123,N_4240,N_4002);
and U6124 (N_6124,N_1197,N_962);
nand U6125 (N_6125,N_2108,N_1428);
and U6126 (N_6126,N_347,N_3397);
nor U6127 (N_6127,N_1418,N_1081);
nor U6128 (N_6128,N_2041,N_2837);
or U6129 (N_6129,N_3663,N_1880);
or U6130 (N_6130,N_3909,N_617);
and U6131 (N_6131,N_3006,N_2016);
nor U6132 (N_6132,N_2277,N_564);
nand U6133 (N_6133,N_1828,N_1746);
or U6134 (N_6134,N_3711,N_1059);
nor U6135 (N_6135,N_1119,N_3135);
or U6136 (N_6136,N_2986,N_4988);
nand U6137 (N_6137,N_4612,N_2889);
or U6138 (N_6138,N_3588,N_2386);
nand U6139 (N_6139,N_3545,N_4994);
nand U6140 (N_6140,N_2317,N_3185);
or U6141 (N_6141,N_2252,N_2557);
nand U6142 (N_6142,N_4913,N_568);
or U6143 (N_6143,N_666,N_2451);
nand U6144 (N_6144,N_552,N_2109);
nor U6145 (N_6145,N_4573,N_2529);
or U6146 (N_6146,N_3737,N_4632);
or U6147 (N_6147,N_2613,N_4833);
nand U6148 (N_6148,N_506,N_2091);
and U6149 (N_6149,N_381,N_3283);
or U6150 (N_6150,N_150,N_783);
nand U6151 (N_6151,N_3844,N_1434);
or U6152 (N_6152,N_2641,N_2806);
or U6153 (N_6153,N_2739,N_2512);
nand U6154 (N_6154,N_2921,N_2093);
and U6155 (N_6155,N_3872,N_4008);
xnor U6156 (N_6156,N_1627,N_7);
or U6157 (N_6157,N_1242,N_2318);
or U6158 (N_6158,N_754,N_4697);
and U6159 (N_6159,N_3096,N_1951);
and U6160 (N_6160,N_4318,N_2761);
nand U6161 (N_6161,N_2832,N_2971);
nor U6162 (N_6162,N_187,N_1793);
nor U6163 (N_6163,N_470,N_1063);
nor U6164 (N_6164,N_4772,N_2742);
nand U6165 (N_6165,N_1705,N_3568);
and U6166 (N_6166,N_2475,N_4491);
and U6167 (N_6167,N_3801,N_2116);
and U6168 (N_6168,N_158,N_407);
and U6169 (N_6169,N_1930,N_3592);
and U6170 (N_6170,N_4405,N_4269);
nand U6171 (N_6171,N_3055,N_1816);
nand U6172 (N_6172,N_4164,N_2177);
or U6173 (N_6173,N_3885,N_598);
and U6174 (N_6174,N_3887,N_2663);
nor U6175 (N_6175,N_4278,N_3958);
nor U6176 (N_6176,N_2678,N_3184);
nor U6177 (N_6177,N_2922,N_784);
and U6178 (N_6178,N_2695,N_3328);
nand U6179 (N_6179,N_3658,N_4973);
and U6180 (N_6180,N_643,N_4578);
nor U6181 (N_6181,N_3968,N_4734);
or U6182 (N_6182,N_4287,N_1893);
or U6183 (N_6183,N_2715,N_1518);
or U6184 (N_6184,N_3258,N_3368);
and U6185 (N_6185,N_3407,N_248);
or U6186 (N_6186,N_3480,N_3772);
nand U6187 (N_6187,N_4120,N_1008);
or U6188 (N_6188,N_4180,N_4100);
nand U6189 (N_6189,N_3238,N_1718);
and U6190 (N_6190,N_613,N_273);
nand U6191 (N_6191,N_1616,N_3022);
nand U6192 (N_6192,N_618,N_4621);
or U6193 (N_6193,N_1531,N_4603);
nand U6194 (N_6194,N_1052,N_172);
or U6195 (N_6195,N_1921,N_654);
nand U6196 (N_6196,N_1650,N_2056);
nand U6197 (N_6197,N_954,N_936);
nor U6198 (N_6198,N_1256,N_3211);
nand U6199 (N_6199,N_1442,N_249);
nand U6200 (N_6200,N_2199,N_1580);
nand U6201 (N_6201,N_3747,N_1779);
or U6202 (N_6202,N_2014,N_3389);
nand U6203 (N_6203,N_1904,N_110);
or U6204 (N_6204,N_3966,N_3125);
or U6205 (N_6205,N_2256,N_4755);
and U6206 (N_6206,N_4977,N_3512);
or U6207 (N_6207,N_3246,N_2142);
and U6208 (N_6208,N_3063,N_345);
and U6209 (N_6209,N_503,N_3345);
and U6210 (N_6210,N_4757,N_1848);
nand U6211 (N_6211,N_1406,N_3482);
nor U6212 (N_6212,N_3031,N_66);
and U6213 (N_6213,N_1620,N_958);
or U6214 (N_6214,N_3582,N_4077);
nand U6215 (N_6215,N_491,N_4702);
nor U6216 (N_6216,N_1078,N_334);
or U6217 (N_6217,N_913,N_660);
or U6218 (N_6218,N_1857,N_2145);
nand U6219 (N_6219,N_4314,N_3585);
nand U6220 (N_6220,N_4668,N_1833);
or U6221 (N_6221,N_280,N_776);
nor U6222 (N_6222,N_3774,N_3443);
nand U6223 (N_6223,N_2315,N_2508);
or U6224 (N_6224,N_4020,N_84);
nor U6225 (N_6225,N_4503,N_4192);
and U6226 (N_6226,N_3739,N_308);
nand U6227 (N_6227,N_382,N_3804);
or U6228 (N_6228,N_291,N_1378);
nor U6229 (N_6229,N_1062,N_1421);
and U6230 (N_6230,N_2959,N_4771);
nor U6231 (N_6231,N_647,N_3404);
or U6232 (N_6232,N_2790,N_567);
nor U6233 (N_6233,N_3510,N_895);
nand U6234 (N_6234,N_3741,N_1265);
nand U6235 (N_6235,N_3423,N_504);
and U6236 (N_6236,N_1867,N_905);
and U6237 (N_6237,N_4625,N_2683);
or U6238 (N_6238,N_3563,N_1383);
or U6239 (N_6239,N_2115,N_292);
and U6240 (N_6240,N_3659,N_329);
nor U6241 (N_6241,N_128,N_294);
and U6242 (N_6242,N_4900,N_663);
or U6243 (N_6243,N_380,N_1664);
nor U6244 (N_6244,N_3141,N_3494);
or U6245 (N_6245,N_189,N_1879);
xnor U6246 (N_6246,N_3616,N_901);
or U6247 (N_6247,N_4706,N_1869);
and U6248 (N_6248,N_513,N_4443);
and U6249 (N_6249,N_4694,N_3760);
nor U6250 (N_6250,N_3891,N_4918);
nor U6251 (N_6251,N_2488,N_4922);
nand U6252 (N_6252,N_2622,N_1034);
nor U6253 (N_6253,N_3466,N_2797);
or U6254 (N_6254,N_476,N_3441);
nor U6255 (N_6255,N_474,N_2759);
or U6256 (N_6256,N_433,N_657);
or U6257 (N_6257,N_3281,N_2789);
and U6258 (N_6258,N_4681,N_3724);
and U6259 (N_6259,N_4903,N_1802);
or U6260 (N_6260,N_3197,N_2015);
or U6261 (N_6261,N_3136,N_2825);
nor U6262 (N_6262,N_2076,N_2914);
nor U6263 (N_6263,N_1086,N_3929);
and U6264 (N_6264,N_1159,N_3707);
nor U6265 (N_6265,N_344,N_3353);
nor U6266 (N_6266,N_4145,N_2010);
nor U6267 (N_6267,N_236,N_2068);
nor U6268 (N_6268,N_4001,N_4223);
or U6269 (N_6269,N_379,N_485);
nand U6270 (N_6270,N_4298,N_3033);
and U6271 (N_6271,N_1115,N_1360);
and U6272 (N_6272,N_745,N_3596);
nand U6273 (N_6273,N_4015,N_818);
and U6274 (N_6274,N_2101,N_1295);
nand U6275 (N_6275,N_4334,N_4981);
nor U6276 (N_6276,N_758,N_3386);
nor U6277 (N_6277,N_2006,N_1626);
nor U6278 (N_6278,N_2933,N_2800);
nor U6279 (N_6279,N_4250,N_193);
or U6280 (N_6280,N_1005,N_2155);
and U6281 (N_6281,N_786,N_118);
or U6282 (N_6282,N_3424,N_3505);
or U6283 (N_6283,N_2384,N_1409);
nand U6284 (N_6284,N_2179,N_2162);
nor U6285 (N_6285,N_321,N_3674);
nand U6286 (N_6286,N_1279,N_3098);
and U6287 (N_6287,N_1574,N_1255);
nor U6288 (N_6288,N_3370,N_4079);
or U6289 (N_6289,N_2029,N_3192);
and U6290 (N_6290,N_1328,N_4992);
and U6291 (N_6291,N_3099,N_2180);
nor U6292 (N_6292,N_3813,N_1849);
nand U6293 (N_6293,N_1395,N_3347);
and U6294 (N_6294,N_3987,N_3988);
and U6295 (N_6295,N_3182,N_945);
and U6296 (N_6296,N_3332,N_1260);
or U6297 (N_6297,N_4980,N_428);
and U6298 (N_6298,N_105,N_1748);
xnor U6299 (N_6299,N_3993,N_188);
and U6300 (N_6300,N_1405,N_3269);
and U6301 (N_6301,N_101,N_4927);
and U6302 (N_6302,N_3324,N_4072);
and U6303 (N_6303,N_3976,N_3539);
nand U6304 (N_6304,N_4623,N_143);
nand U6305 (N_6305,N_547,N_2701);
nor U6306 (N_6306,N_953,N_1474);
nor U6307 (N_6307,N_2217,N_1651);
nand U6308 (N_6308,N_1961,N_2157);
or U6309 (N_6309,N_4045,N_3881);
and U6310 (N_6310,N_1199,N_1478);
nand U6311 (N_6311,N_326,N_4102);
and U6312 (N_6312,N_2915,N_2198);
nand U6313 (N_6313,N_690,N_1883);
nor U6314 (N_6314,N_2974,N_4140);
nor U6315 (N_6315,N_1321,N_4983);
and U6316 (N_6316,N_1819,N_2373);
or U6317 (N_6317,N_1220,N_2251);
nand U6318 (N_6318,N_4422,N_995);
nor U6319 (N_6319,N_4507,N_3752);
nor U6320 (N_6320,N_121,N_4138);
nand U6321 (N_6321,N_1862,N_965);
or U6322 (N_6322,N_4486,N_924);
or U6323 (N_6323,N_2385,N_1496);
nand U6324 (N_6324,N_107,N_4770);
and U6325 (N_6325,N_1967,N_2414);
nand U6326 (N_6326,N_2207,N_3168);
or U6327 (N_6327,N_3913,N_809);
nand U6328 (N_6328,N_457,N_1906);
and U6329 (N_6329,N_3782,N_2928);
nor U6330 (N_6330,N_796,N_4599);
and U6331 (N_6331,N_2600,N_897);
and U6332 (N_6332,N_2255,N_4773);
nor U6333 (N_6333,N_3689,N_2788);
nand U6334 (N_6334,N_2122,N_4791);
nor U6335 (N_6335,N_1699,N_325);
and U6336 (N_6336,N_4199,N_1415);
and U6337 (N_6337,N_2834,N_4985);
or U6338 (N_6338,N_4963,N_1822);
and U6339 (N_6339,N_2230,N_4221);
nand U6340 (N_6340,N_2966,N_2200);
or U6341 (N_6341,N_4305,N_4225);
nand U6342 (N_6342,N_4246,N_4337);
or U6343 (N_6343,N_2822,N_829);
nor U6344 (N_6344,N_3946,N_4412);
and U6345 (N_6345,N_103,N_2203);
or U6346 (N_6346,N_4645,N_652);
or U6347 (N_6347,N_467,N_4124);
and U6348 (N_6348,N_212,N_1598);
nor U6349 (N_6349,N_1900,N_2640);
nor U6350 (N_6350,N_2731,N_3561);
nand U6351 (N_6351,N_1038,N_1843);
or U6352 (N_6352,N_1907,N_4762);
and U6353 (N_6353,N_4564,N_1669);
or U6354 (N_6354,N_930,N_3822);
nor U6355 (N_6355,N_4185,N_889);
and U6356 (N_6356,N_1856,N_1947);
and U6357 (N_6357,N_4325,N_3645);
nand U6358 (N_6358,N_4854,N_14);
nand U6359 (N_6359,N_1345,N_147);
or U6360 (N_6360,N_1237,N_732);
and U6361 (N_6361,N_4735,N_4492);
nor U6362 (N_6362,N_1941,N_2279);
and U6363 (N_6363,N_1087,N_3709);
and U6364 (N_6364,N_2516,N_2638);
nor U6365 (N_6365,N_775,N_2295);
nor U6366 (N_6366,N_4741,N_1683);
or U6367 (N_6367,N_4212,N_704);
and U6368 (N_6368,N_3839,N_3591);
or U6369 (N_6369,N_441,N_3435);
or U6370 (N_6370,N_1104,N_352);
nand U6371 (N_6371,N_2532,N_2539);
xor U6372 (N_6372,N_4729,N_3352);
and U6373 (N_6373,N_4972,N_2035);
nor U6374 (N_6374,N_1677,N_3957);
or U6375 (N_6375,N_993,N_2365);
or U6376 (N_6376,N_4931,N_4319);
nor U6377 (N_6377,N_1487,N_1485);
or U6378 (N_6378,N_2003,N_3234);
and U6379 (N_6379,N_3604,N_3259);
and U6380 (N_6380,N_3898,N_1252);
and U6381 (N_6381,N_4759,N_2455);
nor U6382 (N_6382,N_2060,N_117);
or U6383 (N_6383,N_3682,N_3574);
and U6384 (N_6384,N_4051,N_4556);
nor U6385 (N_6385,N_3691,N_1763);
nand U6386 (N_6386,N_1974,N_157);
nor U6387 (N_6387,N_516,N_1525);
and U6388 (N_6388,N_3077,N_2844);
nor U6389 (N_6389,N_4016,N_4179);
or U6390 (N_6390,N_459,N_2917);
nand U6391 (N_6391,N_769,N_4511);
or U6392 (N_6392,N_2684,N_3294);
or U6393 (N_6393,N_1917,N_383);
and U6394 (N_6394,N_843,N_3643);
or U6395 (N_6395,N_405,N_1916);
nand U6396 (N_6396,N_2407,N_2366);
or U6397 (N_6397,N_2063,N_2787);
and U6398 (N_6398,N_3143,N_4836);
or U6399 (N_6399,N_4315,N_4416);
or U6400 (N_6400,N_4372,N_444);
and U6401 (N_6401,N_2204,N_164);
or U6402 (N_6402,N_1859,N_4151);
and U6403 (N_6403,N_957,N_2243);
nor U6404 (N_6404,N_805,N_1064);
nor U6405 (N_6405,N_1610,N_1979);
nor U6406 (N_6406,N_679,N_3599);
nand U6407 (N_6407,N_819,N_1065);
nand U6408 (N_6408,N_2274,N_4007);
nor U6409 (N_6409,N_4541,N_3924);
or U6410 (N_6410,N_3275,N_57);
nor U6411 (N_6411,N_3878,N_297);
nand U6412 (N_6412,N_3715,N_4870);
or U6413 (N_6413,N_3916,N_4606);
or U6414 (N_6414,N_1100,N_2802);
nor U6415 (N_6415,N_138,N_1226);
nor U6416 (N_6416,N_1486,N_3630);
and U6417 (N_6417,N_1751,N_1966);
and U6418 (N_6418,N_2925,N_3812);
or U6419 (N_6419,N_1955,N_4777);
nor U6420 (N_6420,N_1556,N_4514);
nor U6421 (N_6421,N_140,N_4809);
and U6422 (N_6422,N_3272,N_2012);
nand U6423 (N_6423,N_815,N_4421);
and U6424 (N_6424,N_665,N_2977);
nor U6425 (N_6425,N_4266,N_1926);
nor U6426 (N_6426,N_2719,N_1011);
nor U6427 (N_6427,N_1430,N_2783);
or U6428 (N_6428,N_2549,N_2833);
or U6429 (N_6429,N_3375,N_2361);
and U6430 (N_6430,N_3907,N_3040);
nor U6431 (N_6431,N_1108,N_1855);
and U6432 (N_6432,N_860,N_2491);
or U6433 (N_6433,N_1447,N_3013);
and U6434 (N_6434,N_1399,N_4590);
and U6435 (N_6435,N_2568,N_2767);
and U6436 (N_6436,N_3808,N_1555);
or U6437 (N_6437,N_3501,N_795);
and U6438 (N_6438,N_3989,N_232);
and U6439 (N_6439,N_3828,N_211);
nand U6440 (N_6440,N_1548,N_2859);
and U6441 (N_6441,N_4042,N_1733);
nor U6442 (N_6442,N_919,N_2112);
nor U6443 (N_6443,N_1595,N_104);
or U6444 (N_6444,N_2930,N_4474);
or U6445 (N_6445,N_4942,N_4710);
or U6446 (N_6446,N_1854,N_2706);
and U6447 (N_6447,N_1363,N_3584);
nor U6448 (N_6448,N_888,N_4046);
and U6449 (N_6449,N_1338,N_4874);
or U6450 (N_6450,N_60,N_1807);
nand U6451 (N_6451,N_1581,N_1396);
and U6452 (N_6452,N_1759,N_667);
and U6453 (N_6453,N_3244,N_1134);
nand U6454 (N_6454,N_4857,N_4893);
nand U6455 (N_6455,N_1552,N_4159);
nand U6456 (N_6456,N_4696,N_3181);
or U6457 (N_6457,N_3187,N_3889);
nand U6458 (N_6458,N_1309,N_2154);
or U6459 (N_6459,N_1240,N_3544);
or U6460 (N_6460,N_2707,N_2500);
nand U6461 (N_6461,N_3903,N_3475);
xnor U6462 (N_6462,N_1468,N_2448);
nand U6463 (N_6463,N_2107,N_971);
and U6464 (N_6464,N_2103,N_3716);
and U6465 (N_6465,N_1672,N_1540);
and U6466 (N_6466,N_3794,N_1458);
or U6467 (N_6467,N_4155,N_362);
nand U6468 (N_6468,N_4099,N_3394);
or U6469 (N_6469,N_1861,N_706);
or U6470 (N_6470,N_908,N_4343);
nor U6471 (N_6471,N_4688,N_97);
nor U6472 (N_6472,N_2280,N_3594);
nand U6473 (N_6473,N_1001,N_2666);
or U6474 (N_6474,N_934,N_4622);
nand U6475 (N_6475,N_2735,N_1994);
nand U6476 (N_6476,N_1692,N_1391);
or U6477 (N_6477,N_1791,N_653);
xnor U6478 (N_6478,N_600,N_1125);
nand U6479 (N_6479,N_1446,N_1053);
nor U6480 (N_6480,N_1455,N_1706);
nand U6481 (N_6481,N_4095,N_3327);
nor U6482 (N_6482,N_4394,N_2357);
nor U6483 (N_6483,N_1721,N_2369);
and U6484 (N_6484,N_4153,N_3628);
nand U6485 (N_6485,N_3199,N_834);
nor U6486 (N_6486,N_4480,N_3421);
nor U6487 (N_6487,N_3024,N_3326);
or U6488 (N_6488,N_1608,N_4780);
and U6489 (N_6489,N_4731,N_4236);
or U6490 (N_6490,N_1183,N_4123);
or U6491 (N_6491,N_1587,N_2171);
or U6492 (N_6492,N_3410,N_1232);
and U6493 (N_6493,N_1223,N_3754);
xnor U6494 (N_6494,N_2173,N_3843);
and U6495 (N_6495,N_227,N_394);
and U6496 (N_6496,N_2183,N_4935);
or U6497 (N_6497,N_4549,N_41);
nor U6498 (N_6498,N_605,N_1619);
nand U6499 (N_6499,N_1214,N_771);
or U6500 (N_6500,N_1041,N_3605);
or U6501 (N_6501,N_3240,N_3231);
nand U6502 (N_6502,N_2482,N_1444);
nor U6503 (N_6503,N_448,N_1271);
nand U6504 (N_6504,N_1944,N_2387);
nor U6505 (N_6505,N_2502,N_2740);
or U6506 (N_6506,N_4956,N_1696);
or U6507 (N_6507,N_2430,N_606);
nand U6508 (N_6508,N_4510,N_116);
nor U6509 (N_6509,N_975,N_4856);
and U6510 (N_6510,N_3401,N_295);
nor U6511 (N_6511,N_988,N_238);
and U6512 (N_6512,N_1114,N_4638);
and U6513 (N_6513,N_4447,N_4739);
or U6514 (N_6514,N_0,N_489);
nor U6515 (N_6515,N_3967,N_4680);
or U6516 (N_6516,N_867,N_4889);
and U6517 (N_6517,N_3662,N_2794);
nor U6518 (N_6518,N_1533,N_2320);
nor U6519 (N_6519,N_4501,N_4728);
nand U6520 (N_6520,N_1836,N_2468);
and U6521 (N_6521,N_963,N_3692);
nor U6522 (N_6522,N_2079,N_1098);
and U6523 (N_6523,N_2785,N_4158);
nand U6524 (N_6524,N_4398,N_2791);
nand U6525 (N_6525,N_1512,N_4233);
nor U6526 (N_6526,N_697,N_4075);
or U6527 (N_6527,N_3649,N_2347);
nor U6528 (N_6528,N_1010,N_1397);
and U6529 (N_6529,N_925,N_2956);
and U6530 (N_6530,N_3830,N_2927);
nand U6531 (N_6531,N_1942,N_2470);
or U6532 (N_6532,N_2058,N_4950);
nand U6533 (N_6533,N_1015,N_3618);
and U6534 (N_6534,N_2228,N_1573);
or U6535 (N_6535,N_75,N_2910);
or U6536 (N_6536,N_991,N_1239);
or U6537 (N_6537,N_4387,N_1648);
nor U6538 (N_6538,N_952,N_156);
nor U6539 (N_6539,N_1962,N_2464);
or U6540 (N_6540,N_395,N_2048);
nand U6541 (N_6541,N_4264,N_1470);
nand U6542 (N_6542,N_4830,N_2302);
nand U6543 (N_6543,N_3415,N_2579);
and U6544 (N_6544,N_2973,N_3959);
nand U6545 (N_6545,N_1717,N_3266);
nor U6546 (N_6546,N_4705,N_1702);
and U6547 (N_6547,N_4482,N_1639);
or U6548 (N_6548,N_1277,N_916);
nand U6549 (N_6549,N_2423,N_1762);
and U6550 (N_6550,N_951,N_4767);
or U6551 (N_6551,N_511,N_3291);
or U6552 (N_6552,N_3814,N_1178);
nand U6553 (N_6553,N_4561,N_2380);
and U6554 (N_6554,N_621,N_3156);
and U6555 (N_6555,N_2936,N_4122);
and U6556 (N_6556,N_3789,N_1231);
nand U6557 (N_6557,N_2346,N_4433);
nor U6558 (N_6558,N_4086,N_1632);
and U6559 (N_6559,N_3870,N_3102);
or U6560 (N_6560,N_1659,N_4535);
nand U6561 (N_6561,N_3699,N_18);
nand U6562 (N_6562,N_1173,N_1248);
and U6563 (N_6563,N_3054,N_1489);
and U6564 (N_6564,N_4345,N_2444);
nor U6565 (N_6565,N_3858,N_2);
xor U6566 (N_6566,N_4377,N_571);
nor U6567 (N_6567,N_1887,N_146);
or U6568 (N_6568,N_1401,N_1241);
nor U6569 (N_6569,N_2882,N_578);
and U6570 (N_6570,N_4208,N_4944);
nand U6571 (N_6571,N_1390,N_638);
nand U6572 (N_6572,N_3817,N_1711);
nand U6573 (N_6573,N_1055,N_2397);
and U6574 (N_6574,N_1080,N_4384);
and U6575 (N_6575,N_3028,N_3717);
nor U6576 (N_6576,N_2632,N_247);
and U6577 (N_6577,N_2213,N_3208);
nor U6578 (N_6578,N_3109,N_3495);
nand U6579 (N_6579,N_1837,N_1109);
nand U6580 (N_6580,N_802,N_4247);
nor U6581 (N_6581,N_1835,N_1380);
or U6582 (N_6582,N_1771,N_2765);
nor U6583 (N_6583,N_3132,N_3758);
nor U6584 (N_6584,N_4716,N_1654);
nor U6585 (N_6585,N_4009,N_3385);
nor U6586 (N_6586,N_4078,N_3941);
nand U6587 (N_6587,N_4310,N_2303);
nor U6588 (N_6588,N_3821,N_581);
nor U6589 (N_6589,N_3114,N_2216);
and U6590 (N_6590,N_3590,N_1431);
nor U6591 (N_6591,N_4518,N_4196);
nand U6592 (N_6592,N_2872,N_363);
or U6593 (N_6593,N_3920,N_1801);
and U6594 (N_6594,N_288,N_1565);
or U6595 (N_6595,N_4584,N_2313);
and U6596 (N_6596,N_1870,N_3450);
nor U6597 (N_6597,N_3321,N_1050);
or U6598 (N_6598,N_3091,N_938);
and U6599 (N_6599,N_2017,N_1274);
xor U6600 (N_6600,N_1691,N_3971);
or U6601 (N_6601,N_81,N_3070);
nand U6602 (N_6602,N_1530,N_1697);
nand U6603 (N_6603,N_1977,N_2524);
xor U6604 (N_6604,N_865,N_1553);
nand U6605 (N_6605,N_2434,N_3047);
nand U6606 (N_6606,N_2929,N_2887);
and U6607 (N_6607,N_393,N_1820);
nor U6608 (N_6608,N_2412,N_2547);
and U6609 (N_6609,N_3188,N_2884);
and U6610 (N_6610,N_4277,N_4052);
and U6611 (N_6611,N_3904,N_3695);
nor U6612 (N_6612,N_3491,N_3928);
nand U6613 (N_6613,N_1597,N_234);
nor U6614 (N_6614,N_230,N_3740);
or U6615 (N_6615,N_4171,N_528);
and U6616 (N_6616,N_3615,N_1281);
nand U6617 (N_6617,N_259,N_4937);
nand U6618 (N_6618,N_764,N_3869);
nand U6619 (N_6619,N_588,N_1922);
and U6620 (N_6620,N_715,N_861);
and U6621 (N_6621,N_2840,N_285);
and U6622 (N_6622,N_1261,N_627);
or U6623 (N_6623,N_3728,N_2102);
and U6624 (N_6624,N_4818,N_3453);
and U6625 (N_6625,N_4157,N_1308);
or U6626 (N_6626,N_4558,N_392);
and U6627 (N_6627,N_2644,N_4272);
and U6628 (N_6628,N_3195,N_1787);
and U6629 (N_6629,N_169,N_27);
or U6630 (N_6630,N_984,N_4566);
and U6631 (N_6631,N_3565,N_1515);
nor U6632 (N_6632,N_529,N_4968);
nor U6633 (N_6633,N_3600,N_824);
nand U6634 (N_6634,N_2997,N_2267);
nor U6635 (N_6635,N_4570,N_1615);
nand U6636 (N_6636,N_1327,N_246);
nor U6637 (N_6637,N_53,N_3469);
and U6638 (N_6638,N_1168,N_2693);
nand U6639 (N_6639,N_1851,N_3785);
nor U6640 (N_6640,N_2503,N_3);
and U6641 (N_6641,N_4933,N_4509);
nand U6642 (N_6642,N_4607,N_1821);
and U6643 (N_6643,N_2437,N_4536);
nor U6644 (N_6644,N_2042,N_4691);
or U6645 (N_6645,N_2117,N_2920);
nor U6646 (N_6646,N_2457,N_3733);
nor U6647 (N_6647,N_1520,N_1166);
or U6648 (N_6648,N_4531,N_1928);
nand U6649 (N_6649,N_4774,N_4810);
or U6650 (N_6650,N_2191,N_1023);
or U6651 (N_6651,N_701,N_2868);
nor U6652 (N_6652,N_3953,N_4521);
nor U6653 (N_6653,N_2194,N_3308);
or U6654 (N_6654,N_2031,N_4143);
or U6655 (N_6655,N_1998,N_4131);
nor U6656 (N_6656,N_4583,N_3250);
and U6657 (N_6657,N_726,N_3371);
and U6658 (N_6658,N_1747,N_302);
and U6659 (N_6659,N_2879,N_1938);
or U6660 (N_6660,N_1927,N_2234);
and U6661 (N_6661,N_2406,N_678);
nor U6662 (N_6662,N_2940,N_2144);
and U6663 (N_6663,N_4630,N_2954);
nand U6664 (N_6664,N_1643,N_2801);
nor U6665 (N_6665,N_126,N_4709);
nand U6666 (N_6666,N_2633,N_4899);
or U6667 (N_6667,N_3612,N_1872);
nor U6668 (N_6668,N_200,N_3241);
nand U6669 (N_6669,N_2390,N_640);
or U6670 (N_6670,N_3636,N_1142);
nand U6671 (N_6671,N_2087,N_313);
and U6672 (N_6672,N_4370,N_2190);
and U6673 (N_6673,N_4961,N_4047);
nand U6674 (N_6674,N_521,N_4226);
or U6675 (N_6675,N_3732,N_2069);
and U6676 (N_6676,N_733,N_2664);
or U6677 (N_6677,N_2826,N_388);
nor U6678 (N_6678,N_2548,N_2670);
or U6679 (N_6679,N_2289,N_1910);
nand U6680 (N_6680,N_2559,N_4678);
or U6681 (N_6681,N_4173,N_2139);
or U6682 (N_6682,N_98,N_3580);
or U6683 (N_6683,N_766,N_96);
and U6684 (N_6684,N_2819,N_4936);
or U6685 (N_6685,N_3133,N_3103);
nand U6686 (N_6686,N_442,N_2565);
nand U6687 (N_6687,N_4884,N_3874);
xor U6688 (N_6688,N_493,N_898);
nand U6689 (N_6689,N_2852,N_1263);
nor U6690 (N_6690,N_137,N_4906);
nor U6691 (N_6691,N_1275,N_3762);
or U6692 (N_6692,N_3338,N_4152);
nand U6693 (N_6693,N_3504,N_2176);
and U6694 (N_6694,N_2736,N_804);
nand U6695 (N_6695,N_4149,N_1824);
nor U6696 (N_6696,N_208,N_289);
or U6697 (N_6697,N_2311,N_3513);
nand U6698 (N_6698,N_4588,N_3751);
nor U6699 (N_6699,N_896,N_77);
nand U6700 (N_6700,N_3412,N_918);
xnor U6701 (N_6701,N_823,N_1952);
nand U6702 (N_6702,N_4092,N_3790);
or U6703 (N_6703,N_3017,N_4207);
nor U6704 (N_6704,N_1375,N_2368);
nor U6705 (N_6705,N_807,N_2828);
and U6706 (N_6706,N_2223,N_2393);
and U6707 (N_6707,N_514,N_2531);
and U6708 (N_6708,N_2808,N_1195);
and U6709 (N_6709,N_3073,N_3298);
nor U6710 (N_6710,N_178,N_4778);
and U6711 (N_6711,N_4061,N_3300);
nand U6712 (N_6712,N_699,N_2426);
nor U6713 (N_6713,N_4262,N_1743);
nor U6714 (N_6714,N_55,N_2646);
nor U6715 (N_6715,N_920,N_2307);
and U6716 (N_6716,N_2135,N_4855);
nand U6717 (N_6717,N_2566,N_3755);
nand U6718 (N_6718,N_4362,N_4618);
nor U6719 (N_6719,N_3981,N_1978);
or U6720 (N_6720,N_2718,N_1018);
nor U6721 (N_6721,N_4883,N_2262);
or U6722 (N_6722,N_917,N_4951);
nand U6723 (N_6723,N_2328,N_322);
and U6724 (N_6724,N_4267,N_1866);
and U6725 (N_6725,N_3057,N_3601);
nand U6726 (N_6726,N_3842,N_3578);
or U6727 (N_6727,N_1755,N_838);
nand U6728 (N_6728,N_1480,N_703);
nand U6729 (N_6729,N_3745,N_2100);
and U6730 (N_6730,N_3866,N_4244);
nor U6731 (N_6731,N_2244,N_3635);
and U6732 (N_6732,N_3060,N_525);
and U6733 (N_6733,N_26,N_3122);
and U6734 (N_6734,N_2113,N_4802);
and U6735 (N_6735,N_3863,N_2589);
and U6736 (N_6736,N_4781,N_4442);
or U6737 (N_6737,N_912,N_2795);
nor U6738 (N_6738,N_1132,N_1494);
nand U6739 (N_6739,N_4022,N_2746);
or U6740 (N_6740,N_2073,N_1035);
nand U6741 (N_6741,N_3899,N_4035);
and U6742 (N_6742,N_4895,N_4967);
nor U6743 (N_6743,N_385,N_4776);
and U6744 (N_6744,N_1891,N_1112);
nor U6745 (N_6745,N_910,N_739);
or U6746 (N_6746,N_2593,N_1912);
nor U6747 (N_6747,N_2314,N_3012);
nand U6748 (N_6748,N_378,N_33);
nor U6749 (N_6749,N_2768,N_4803);
or U6750 (N_6750,N_3896,N_2421);
or U6751 (N_6751,N_4611,N_3134);
nor U6752 (N_6752,N_1934,N_3880);
nor U6753 (N_6753,N_4118,N_4929);
nor U6754 (N_6754,N_4214,N_1410);
nand U6755 (N_6755,N_3524,N_4805);
or U6756 (N_6756,N_4399,N_749);
and U6757 (N_6757,N_1943,N_3361);
nand U6758 (N_6758,N_220,N_1394);
and U6759 (N_6759,N_659,N_3936);
nor U6760 (N_6760,N_93,N_3186);
nand U6761 (N_6761,N_3438,N_915);
and U6762 (N_6762,N_518,N_4736);
or U6763 (N_6763,N_148,N_281);
nand U6764 (N_6764,N_631,N_3215);
or U6765 (N_6765,N_32,N_3288);
nor U6766 (N_6766,N_1734,N_204);
or U6767 (N_6767,N_3868,N_2185);
or U6768 (N_6768,N_3426,N_2677);
or U6769 (N_6769,N_3174,N_3549);
and U6770 (N_6770,N_3897,N_4548);
nand U6771 (N_6771,N_2440,N_1155);
or U6772 (N_6772,N_2660,N_3823);
nor U6773 (N_6773,N_2165,N_2059);
nor U6774 (N_6774,N_4887,N_4050);
nor U6775 (N_6775,N_3263,N_2821);
nor U6776 (N_6776,N_3084,N_1149);
nor U6777 (N_6777,N_4488,N_876);
and U6778 (N_6778,N_1545,N_3543);
nor U6779 (N_6779,N_1307,N_2224);
nand U6780 (N_6780,N_54,N_3776);
nor U6781 (N_6781,N_4286,N_4389);
and U6782 (N_6782,N_4036,N_4363);
nor U6783 (N_6783,N_1572,N_4200);
and U6784 (N_6784,N_3557,N_2123);
and U6785 (N_6785,N_4427,N_3226);
or U6786 (N_6786,N_3610,N_4454);
nor U6787 (N_6787,N_1429,N_16);
nand U6788 (N_6788,N_630,N_153);
nand U6789 (N_6789,N_2958,N_4896);
nor U6790 (N_6790,N_3377,N_846);
nand U6791 (N_6791,N_2708,N_4434);
nand U6792 (N_6792,N_1362,N_3248);
or U6793 (N_6793,N_3158,N_2571);
nor U6794 (N_6794,N_3422,N_3992);
nand U6795 (N_6795,N_2717,N_366);
and U6796 (N_6796,N_932,N_74);
nand U6797 (N_6797,N_4415,N_1457);
and U6798 (N_6798,N_4202,N_1090);
and U6799 (N_6799,N_4843,N_2606);
nor U6800 (N_6800,N_300,N_928);
nor U6801 (N_6801,N_403,N_1547);
or U6802 (N_6802,N_1140,N_2140);
nand U6803 (N_6803,N_2364,N_4279);
nand U6804 (N_6804,N_1544,N_3703);
or U6805 (N_6805,N_1074,N_705);
nor U6806 (N_6806,N_4624,N_2861);
and U6807 (N_6807,N_3573,N_2533);
or U6808 (N_6808,N_1674,N_3002);
nand U6809 (N_6809,N_319,N_1201);
and U6810 (N_6810,N_3803,N_4273);
or U6811 (N_6811,N_4429,N_3852);
nor U6812 (N_6812,N_3221,N_1984);
and U6813 (N_6813,N_2090,N_4346);
or U6814 (N_6814,N_3380,N_2519);
nor U6815 (N_6815,N_2410,N_2774);
nor U6816 (N_6816,N_1543,N_3161);
nand U6817 (N_6817,N_4923,N_1386);
nand U6818 (N_6818,N_870,N_4581);
and U6819 (N_6819,N_2391,N_268);
nand U6820 (N_6820,N_4292,N_1667);
nand U6821 (N_6821,N_28,N_2321);
and U6822 (N_6822,N_4203,N_3223);
or U6823 (N_6823,N_3632,N_4213);
and U6824 (N_6824,N_2136,N_4753);
nor U6825 (N_6825,N_561,N_1991);
or U6826 (N_6826,N_515,N_3414);
nor U6827 (N_6827,N_179,N_1131);
nand U6828 (N_6828,N_1582,N_3894);
nand U6829 (N_6829,N_43,N_862);
nor U6830 (N_6830,N_3431,N_3061);
nor U6831 (N_6831,N_3606,N_86);
and U6832 (N_6832,N_2866,N_1365);
nor U6833 (N_6833,N_479,N_1299);
and U6834 (N_6834,N_2891,N_1777);
nor U6835 (N_6835,N_4787,N_2322);
nor U6836 (N_6836,N_1116,N_4614);
and U6837 (N_6837,N_4560,N_3444);
nor U6838 (N_6838,N_3005,N_505);
or U6839 (N_6839,N_1088,N_2525);
nand U6840 (N_6840,N_2722,N_1056);
or U6841 (N_6841,N_4742,N_1765);
nand U6842 (N_6842,N_1047,N_2546);
and U6843 (N_6843,N_4797,N_4136);
nor U6844 (N_6844,N_3963,N_1141);
nor U6845 (N_6845,N_2392,N_3396);
and U6846 (N_6846,N_2760,N_1687);
nor U6847 (N_6847,N_277,N_3514);
or U6848 (N_6848,N_1823,N_887);
nor U6849 (N_6849,N_3980,N_1099);
or U6850 (N_6850,N_3383,N_182);
nand U6851 (N_6851,N_3718,N_4743);
nand U6852 (N_6852,N_4859,N_2550);
and U6853 (N_6853,N_422,N_4132);
or U6854 (N_6854,N_4517,N_4718);
and U6855 (N_6855,N_3049,N_4477);
or U6856 (N_6856,N_1103,N_1939);
nand U6857 (N_6857,N_3523,N_2592);
and U6858 (N_6858,N_583,N_3986);
or U6859 (N_6859,N_3940,N_36);
nand U6860 (N_6860,N_4024,N_2218);
nand U6861 (N_6861,N_853,N_2895);
nand U6862 (N_6862,N_1089,N_1113);
or U6863 (N_6863,N_2692,N_3818);
nand U6864 (N_6864,N_1032,N_4448);
and U6865 (N_6865,N_651,N_4156);
nand U6866 (N_6866,N_914,N_2363);
and U6867 (N_6867,N_1864,N_2404);
and U6868 (N_6868,N_4462,N_4580);
nor U6869 (N_6869,N_2873,N_155);
nor U6870 (N_6870,N_2659,N_670);
nor U6871 (N_6871,N_2388,N_4436);
nand U6872 (N_6872,N_4783,N_2089);
nor U6873 (N_6873,N_1376,N_233);
and U6874 (N_6874,N_3529,N_3696);
nand U6875 (N_6875,N_681,N_1624);
nand U6876 (N_6876,N_2065,N_4300);
nand U6877 (N_6877,N_2033,N_868);
and U6878 (N_6878,N_2679,N_2563);
or U6879 (N_6879,N_4698,N_3723);
nand U6880 (N_6880,N_1665,N_3433);
or U6881 (N_6881,N_1350,N_1877);
nand U6882 (N_6882,N_482,N_4381);
nand U6883 (N_6883,N_2319,N_439);
or U6884 (N_6884,N_223,N_713);
and U6885 (N_6885,N_480,N_4091);
and U6886 (N_6886,N_2598,N_4667);
and U6887 (N_6887,N_3008,N_1948);
or U6888 (N_6888,N_4083,N_4845);
or U6889 (N_6889,N_1945,N_774);
nor U6890 (N_6890,N_327,N_541);
and U6891 (N_6891,N_1666,N_361);
nand U6892 (N_6892,N_2764,N_4167);
nand U6893 (N_6893,N_946,N_1204);
and U6894 (N_6894,N_1980,N_1122);
or U6895 (N_6895,N_1432,N_751);
and U6896 (N_6896,N_4892,N_2685);
nand U6897 (N_6897,N_4485,N_2643);
or U6898 (N_6898,N_4837,N_3938);
and U6899 (N_6899,N_2294,N_1310);
nand U6900 (N_6900,N_629,N_2445);
and U6901 (N_6901,N_4908,N_3602);
nor U6902 (N_6902,N_4306,N_2259);
and U6903 (N_6903,N_2962,N_3204);
or U6904 (N_6904,N_2637,N_463);
nor U6905 (N_6905,N_198,N_76);
nand U6906 (N_6906,N_2326,N_3700);
nor U6907 (N_6907,N_3978,N_1335);
or U6908 (N_6908,N_88,N_3773);
nand U6909 (N_6909,N_3960,N_737);
nor U6910 (N_6910,N_3113,N_1202);
nor U6911 (N_6911,N_2075,N_2161);
nor U6912 (N_6912,N_1278,N_3998);
and U6913 (N_6913,N_4417,N_1228);
or U6914 (N_6914,N_2494,N_3964);
or U6915 (N_6915,N_4484,N_2239);
nor U6916 (N_6916,N_1935,N_2994);
and U6917 (N_6917,N_2714,N_1794);
and U6918 (N_6918,N_68,N_1937);
nor U6919 (N_6919,N_3847,N_3634);
nand U6920 (N_6920,N_2201,N_2471);
nand U6921 (N_6921,N_814,N_4765);
nor U6922 (N_6922,N_2047,N_3090);
and U6923 (N_6923,N_1060,N_3076);
and U6924 (N_6924,N_3666,N_3160);
and U6925 (N_6925,N_4825,N_2358);
nor U6926 (N_6926,N_2672,N_1294);
or U6927 (N_6927,N_4054,N_3119);
or U6928 (N_6928,N_2225,N_2153);
nor U6929 (N_6929,N_1154,N_23);
nor U6930 (N_6930,N_370,N_842);
and U6931 (N_6931,N_2309,N_2057);
nand U6932 (N_6932,N_141,N_2472);
and U6933 (N_6933,N_3669,N_4215);
nor U6934 (N_6934,N_3147,N_4111);
and U6935 (N_6935,N_4174,N_192);
and U6936 (N_6936,N_360,N_2355);
or U6937 (N_6937,N_4685,N_339);
nor U6938 (N_6938,N_2874,N_3194);
or U6939 (N_6939,N_262,N_1876);
nand U6940 (N_6940,N_4934,N_3472);
nor U6941 (N_6941,N_4820,N_530);
or U6942 (N_6942,N_970,N_2815);
nor U6943 (N_6943,N_1569,N_1825);
nand U6944 (N_6944,N_412,N_4475);
and U6945 (N_6945,N_95,N_3680);
nand U6946 (N_6946,N_2291,N_4216);
or U6947 (N_6947,N_2399,N_1756);
nand U6948 (N_6948,N_3358,N_2438);
xor U6949 (N_6949,N_1905,N_602);
and U6950 (N_6950,N_446,N_4360);
or U6951 (N_6951,N_3374,N_1903);
xnor U6952 (N_6952,N_359,N_4283);
nand U6953 (N_6953,N_2980,N_2501);
nand U6954 (N_6954,N_2282,N_3629);
nand U6955 (N_6955,N_1946,N_1206);
and U6956 (N_6956,N_1267,N_2877);
nor U6957 (N_6957,N_3032,N_2174);
or U6958 (N_6958,N_1622,N_943);
or U6959 (N_6959,N_1780,N_2214);
nand U6960 (N_6960,N_1022,N_1838);
or U6961 (N_6961,N_1840,N_4349);
and U6962 (N_6962,N_2584,N_3743);
nand U6963 (N_6963,N_4500,N_562);
and U6964 (N_6964,N_1303,N_410);
and U6965 (N_6965,N_59,N_1557);
xor U6966 (N_6966,N_4424,N_2842);
nor U6967 (N_6967,N_736,N_1017);
nor U6968 (N_6968,N_1227,N_3820);
nor U6969 (N_6969,N_1268,N_772);
nand U6970 (N_6970,N_3705,N_3280);
or U6971 (N_6971,N_2651,N_1046);
or U6972 (N_6972,N_4834,N_4596);
or U6973 (N_6973,N_1051,N_2271);
nand U6974 (N_6974,N_2227,N_785);
nor U6975 (N_6975,N_3914,N_2061);
nand U6976 (N_6976,N_4916,N_3729);
and U6977 (N_6977,N_2827,N_4840);
or U6978 (N_6978,N_2530,N_2270);
or U6979 (N_6979,N_1493,N_1949);
and U6980 (N_6980,N_2901,N_2851);
nand U6981 (N_6981,N_1028,N_4322);
and U6982 (N_6982,N_1815,N_1708);
or U6983 (N_6983,N_4775,N_2812);
and U6984 (N_6984,N_250,N_3918);
or U6985 (N_6985,N_1604,N_3349);
and U6986 (N_6986,N_4364,N_584);
and U6987 (N_6987,N_2266,N_144);
nand U6988 (N_6988,N_4746,N_576);
or U6989 (N_6989,N_3900,N_3546);
or U6990 (N_6990,N_1024,N_3051);
nand U6991 (N_6991,N_1211,N_245);
nand U6992 (N_6992,N_2186,N_2979);
and U6993 (N_6993,N_673,N_3331);
nand U6994 (N_6994,N_2630,N_4669);
and U6995 (N_6995,N_161,N_4749);
nand U6996 (N_6996,N_4407,N_649);
and U6997 (N_6997,N_2586,N_4995);
or U6998 (N_6998,N_4301,N_3330);
nor U6999 (N_6999,N_2652,N_254);
or U7000 (N_7000,N_4779,N_3927);
nor U7001 (N_7001,N_3547,N_3577);
and U7002 (N_7002,N_4550,N_4652);
nor U7003 (N_7003,N_2000,N_398);
nor U7004 (N_7004,N_15,N_714);
or U7005 (N_7005,N_2923,N_3944);
and U7006 (N_7006,N_944,N_2158);
or U7007 (N_7007,N_2905,N_708);
nand U7008 (N_7008,N_2614,N_4814);
and U7009 (N_7009,N_2668,N_1788);
nor U7010 (N_7010,N_458,N_3761);
nand U7011 (N_7011,N_4962,N_3196);
and U7012 (N_7012,N_1576,N_1842);
or U7013 (N_7013,N_3614,N_2520);
nor U7014 (N_7014,N_210,N_707);
nand U7015 (N_7015,N_3735,N_941);
or U7016 (N_7016,N_1284,N_445);
and U7017 (N_7017,N_1593,N_3229);
and U7018 (N_7018,N_4975,N_61);
nor U7019 (N_7019,N_1165,N_1776);
or U7020 (N_7020,N_2876,N_1954);
or U7021 (N_7021,N_89,N_4971);
or U7022 (N_7022,N_1367,N_2985);
nand U7023 (N_7023,N_2443,N_4280);
nand U7024 (N_7024,N_3069,N_716);
nand U7025 (N_7025,N_1990,N_4949);
nor U7026 (N_7026,N_2490,N_4476);
nor U7027 (N_7027,N_1641,N_4665);
nand U7028 (N_7028,N_494,N_1352);
or U7029 (N_7029,N_471,N_1612);
nor U7030 (N_7030,N_2675,N_3437);
nor U7031 (N_7031,N_3292,N_160);
or U7032 (N_7032,N_857,N_1083);
nand U7033 (N_7033,N_1411,N_487);
nor U7034 (N_7034,N_4426,N_303);
nor U7035 (N_7035,N_2509,N_1986);
nand U7036 (N_7036,N_214,N_3848);
and U7037 (N_7037,N_1829,N_3949);
nand U7038 (N_7038,N_2008,N_3020);
or U7039 (N_7039,N_4938,N_1351);
nor U7040 (N_7040,N_2189,N_3583);
and U7041 (N_7041,N_2104,N_3166);
nor U7042 (N_7042,N_4722,N_1929);
or U7043 (N_7043,N_3793,N_3305);
nand U7044 (N_7044,N_2596,N_4948);
and U7045 (N_7045,N_3152,N_3313);
or U7046 (N_7046,N_3484,N_1896);
nand U7047 (N_7047,N_955,N_4604);
or U7048 (N_7048,N_3683,N_1329);
nor U7049 (N_7049,N_490,N_2476);
nand U7050 (N_7050,N_3402,N_644);
or U7051 (N_7051,N_1417,N_1126);
and U7052 (N_7052,N_664,N_3116);
nand U7053 (N_7053,N_1671,N_2156);
or U7054 (N_7054,N_4408,N_1546);
nor U7055 (N_7055,N_1259,N_623);
or U7056 (N_7056,N_1054,N_799);
nor U7057 (N_7057,N_1753,N_279);
nor U7058 (N_7058,N_251,N_3282);
nor U7059 (N_7059,N_3376,N_2038);
nand U7060 (N_7060,N_1382,N_1313);
nor U7061 (N_7061,N_2620,N_2304);
nor U7062 (N_7062,N_3357,N_3108);
nor U7063 (N_7063,N_2148,N_242);
and U7064 (N_7064,N_1724,N_4575);
nand U7065 (N_7065,N_112,N_111);
nor U7066 (N_7066,N_3690,N_1625);
or U7067 (N_7067,N_3436,N_1196);
nand U7068 (N_7068,N_3977,N_2778);
nand U7069 (N_7069,N_4030,N_3694);
or U7070 (N_7070,N_1107,N_3526);
nand U7071 (N_7071,N_4732,N_2836);
nand U7072 (N_7072,N_858,N_956);
or U7073 (N_7073,N_4452,N_2698);
or U7074 (N_7074,N_4396,N_1895);
and U7075 (N_7075,N_1209,N_1461);
and U7076 (N_7076,N_1701,N_686);
and U7077 (N_7077,N_1644,N_2149);
or U7078 (N_7078,N_3442,N_4976);
and U7079 (N_7079,N_1030,N_2650);
and U7080 (N_7080,N_2043,N_3566);
nand U7081 (N_7081,N_3408,N_586);
nor U7082 (N_7082,N_1013,N_1225);
and U7083 (N_7083,N_3654,N_3834);
nand U7084 (N_7084,N_1513,N_674);
nand U7085 (N_7085,N_2688,N_2702);
and U7086 (N_7086,N_3487,N_3045);
and U7087 (N_7087,N_4056,N_1586);
nand U7088 (N_7088,N_4947,N_145);
or U7089 (N_7089,N_2264,N_4660);
nor U7090 (N_7090,N_4397,N_2245);
nor U7091 (N_7091,N_4231,N_2120);
and U7092 (N_7092,N_2989,N_257);
nor U7093 (N_7093,N_645,N_333);
nand U7094 (N_7094,N_2249,N_2880);
nand U7095 (N_7095,N_3934,N_1043);
and U7096 (N_7096,N_3471,N_2648);
nand U7097 (N_7097,N_3956,N_1147);
nor U7098 (N_7098,N_2258,N_4882);
nand U7099 (N_7099,N_4999,N_4869);
nor U7100 (N_7100,N_903,N_3954);
or U7101 (N_7101,N_1534,N_4189);
nor U7102 (N_7102,N_4520,N_2597);
nand U7103 (N_7103,N_134,N_553);
and U7104 (N_7104,N_4087,N_4458);
nand U7105 (N_7105,N_3092,N_1466);
or U7106 (N_7106,N_2210,N_206);
nand U7107 (N_7107,N_1020,N_3062);
and U7108 (N_7108,N_3253,N_3372);
or U7109 (N_7109,N_2246,N_2725);
and U7110 (N_7110,N_2422,N_293);
nor U7111 (N_7111,N_1124,N_4033);
nand U7112 (N_7112,N_376,N_1067);
nor U7113 (N_7113,N_718,N_3509);
nand U7114 (N_7114,N_1524,N_438);
nand U7115 (N_7115,N_4170,N_3937);
or U7116 (N_7116,N_305,N_4299);
nand U7117 (N_7117,N_2341,N_1646);
and U7118 (N_7118,N_166,N_239);
nor U7119 (N_7119,N_1613,N_4382);
nor U7120 (N_7120,N_3418,N_2250);
nor U7121 (N_7121,N_2429,N_3533);
or U7122 (N_7122,N_2796,N_1645);
and U7123 (N_7123,N_2050,N_1630);
or U7124 (N_7124,N_3845,N_2427);
nor U7125 (N_7125,N_1591,N_2576);
nor U7126 (N_7126,N_4954,N_400);
nand U7127 (N_7127,N_2370,N_3446);
and U7128 (N_7128,N_551,N_3118);
or U7129 (N_7129,N_4369,N_1238);
nand U7130 (N_7130,N_102,N_1491);
or U7131 (N_7131,N_1488,N_1452);
nand U7132 (N_7132,N_1508,N_1340);
or U7133 (N_7133,N_1618,N_2312);
nand U7134 (N_7134,N_2536,N_3642);
nand U7135 (N_7135,N_4115,N_4602);
nor U7136 (N_7136,N_4703,N_875);
or U7137 (N_7137,N_4402,N_4175);
nor U7138 (N_7138,N_2477,N_1716);
or U7139 (N_7139,N_1884,N_1959);
nor U7140 (N_7140,N_2896,N_3939);
or U7141 (N_7141,N_377,N_1860);
or U7142 (N_7142,N_2964,N_3428);
nor U7143 (N_7143,N_3979,N_1438);
nor U7144 (N_7144,N_999,N_608);
nor U7145 (N_7145,N_1550,N_4062);
or U7146 (N_7146,N_2991,N_4027);
and U7147 (N_7147,N_2127,N_4260);
or U7148 (N_7148,N_811,N_3727);
or U7149 (N_7149,N_1175,N_2114);
or U7150 (N_7150,N_149,N_3864);
nor U7151 (N_7151,N_3764,N_267);
and U7152 (N_7152,N_4057,N_4467);
xor U7153 (N_7153,N_3456,N_355);
nand U7154 (N_7154,N_1719,N_2829);
nand U7155 (N_7155,N_3833,N_3205);
and U7156 (N_7156,N_4498,N_4941);
or U7157 (N_7157,N_2697,N_191);
nand U7158 (N_7158,N_878,N_4150);
and U7159 (N_7159,N_4380,N_201);
or U7160 (N_7160,N_4851,N_4886);
or U7161 (N_7161,N_4162,N_1729);
nand U7162 (N_7162,N_2350,N_4815);
nor U7163 (N_7163,N_2028,N_4589);
nand U7164 (N_7164,N_4670,N_3710);
or U7165 (N_7165,N_1745,N_1551);
or U7166 (N_7166,N_3923,N_3905);
and U7167 (N_7167,N_3759,N_2286);
nand U7168 (N_7168,N_3097,N_2080);
nor U7169 (N_7169,N_2543,N_1469);
nor U7170 (N_7170,N_3213,N_4878);
nand U7171 (N_7171,N_2574,N_4049);
nor U7172 (N_7172,N_4393,N_4659);
or U7173 (N_7173,N_840,N_2094);
nor U7174 (N_7174,N_3190,N_2290);
nand U7175 (N_7175,N_4594,N_4974);
nand U7176 (N_7176,N_87,N_4241);
and U7177 (N_7177,N_4435,N_165);
and U7178 (N_7178,N_2070,N_3089);
and U7179 (N_7179,N_4831,N_1095);
nand U7180 (N_7180,N_4715,N_1302);
nand U7181 (N_7181,N_4819,N_252);
nor U7182 (N_7182,N_1826,N_219);
or U7183 (N_7183,N_3746,N_328);
or U7184 (N_7184,N_1424,N_3893);
and U7185 (N_7185,N_3220,N_51);
or U7186 (N_7186,N_3719,N_4348);
or U7187 (N_7187,N_2254,N_3025);
or U7188 (N_7188,N_3261,N_437);
or U7189 (N_7189,N_4070,N_4341);
nand U7190 (N_7190,N_2339,N_2561);
nor U7191 (N_7191,N_131,N_1805);
nand U7192 (N_7192,N_3846,N_3052);
nor U7193 (N_7193,N_3802,N_4000);
and U7194 (N_7194,N_1535,N_4376);
nand U7195 (N_7195,N_1585,N_1600);
nor U7196 (N_7196,N_79,N_4165);
and U7197 (N_7197,N_1504,N_4097);
nand U7198 (N_7198,N_477,N_747);
and U7199 (N_7199,N_3569,N_687);
or U7200 (N_7200,N_1164,N_1106);
nor U7201 (N_7201,N_4987,N_650);
and U7202 (N_7202,N_3315,N_228);
nor U7203 (N_7203,N_837,N_2168);
or U7204 (N_7204,N_2004,N_2647);
or U7205 (N_7205,N_1902,N_3589);
or U7206 (N_7206,N_1186,N_243);
and U7207 (N_7207,N_1341,N_4168);
nand U7208 (N_7208,N_763,N_2362);
nand U7209 (N_7209,N_415,N_2799);
xnor U7210 (N_7210,N_2924,N_1439);
nand U7211 (N_7211,N_4768,N_4864);
nor U7212 (N_7212,N_177,N_2639);
nor U7213 (N_7213,N_4639,N_2128);
nand U7214 (N_7214,N_540,N_1772);
nand U7215 (N_7215,N_2124,N_1976);
nor U7216 (N_7216,N_756,N_4184);
nor U7217 (N_7217,N_2084,N_950);
and U7218 (N_7218,N_526,N_3943);
or U7219 (N_7219,N_464,N_519);
or U7220 (N_7220,N_270,N_848);
nor U7221 (N_7221,N_996,N_1913);
and U7222 (N_7222,N_4121,N_4966);
or U7223 (N_7223,N_3035,N_1347);
nand U7224 (N_7224,N_4428,N_3750);
nor U7225 (N_7225,N_3925,N_4423);
nor U7226 (N_7226,N_2253,N_2558);
nor U7227 (N_7227,N_720,N_1464);
and U7228 (N_7228,N_3459,N_4457);
nand U7229 (N_7229,N_3516,N_724);
nor U7230 (N_7230,N_1953,N_2838);
nor U7231 (N_7231,N_1675,N_6);
and U7232 (N_7232,N_1084,N_2944);
nand U7233 (N_7233,N_264,N_2961);
nor U7234 (N_7234,N_4726,N_2945);
nand U7235 (N_7235,N_58,N_1117);
nand U7236 (N_7236,N_611,N_3333);
and U7237 (N_7237,N_539,N_4989);
nor U7238 (N_7238,N_3503,N_2055);
or U7239 (N_7239,N_3210,N_492);
and U7240 (N_7240,N_4323,N_2625);
nor U7241 (N_7241,N_3996,N_3552);
and U7242 (N_7242,N_2485,N_114);
or U7243 (N_7243,N_2420,N_2053);
nand U7244 (N_7244,N_3902,N_2521);
and U7245 (N_7245,N_3532,N_1723);
xor U7246 (N_7246,N_891,N_832);
or U7247 (N_7247,N_1300,N_3515);
or U7248 (N_7248,N_4113,N_350);
or U7249 (N_7249,N_1850,N_3720);
nand U7250 (N_7250,N_3425,N_968);
or U7251 (N_7251,N_2036,N_2442);
or U7252 (N_7252,N_4793,N_2758);
and U7253 (N_7253,N_2099,N_331);
or U7254 (N_7254,N_2352,N_768);
or U7255 (N_7255,N_1695,N_414);
or U7256 (N_7256,N_1349,N_2604);
and U7257 (N_7257,N_2400,N_2354);
nand U7258 (N_7258,N_4711,N_4862);
and U7259 (N_7259,N_2545,N_3836);
and U7260 (N_7260,N_231,N_1678);
nor U7261 (N_7261,N_4172,N_2129);
nor U7262 (N_7262,N_1590,N_4324);
and U7263 (N_7263,N_3827,N_3757);
or U7264 (N_7264,N_610,N_2863);
nand U7265 (N_7265,N_2052,N_1564);
and U7266 (N_7266,N_1498,N_1009);
nand U7267 (N_7267,N_559,N_1172);
nor U7268 (N_7268,N_894,N_99);
nor U7269 (N_7269,N_3178,N_1373);
nor U7270 (N_7270,N_1940,N_4275);
nand U7271 (N_7271,N_1834,N_4591);
nand U7272 (N_7272,N_3805,N_1661);
or U7273 (N_7273,N_4064,N_3004);
and U7274 (N_7274,N_4631,N_22);
or U7275 (N_7275,N_3177,N_4490);
nand U7276 (N_7276,N_4114,N_554);
and U7277 (N_7277,N_4071,N_3164);
or U7278 (N_7278,N_1538,N_2892);
and U7279 (N_7279,N_986,N_1617);
nor U7280 (N_7280,N_4939,N_1236);
or U7281 (N_7281,N_2151,N_4658);
nor U7282 (N_7282,N_3901,N_1334);
nand U7283 (N_7283,N_4662,N_1025);
nor U7284 (N_7284,N_546,N_2716);
nand U7285 (N_7285,N_3336,N_2504);
or U7286 (N_7286,N_3792,N_94);
nand U7287 (N_7287,N_136,N_3819);
and U7288 (N_7288,N_336,N_4401);
nor U7289 (N_7289,N_822,N_4750);
nor U7290 (N_7290,N_1739,N_2665);
or U7291 (N_7291,N_2034,N_3179);
nand U7292 (N_7292,N_4945,N_46);
nand U7293 (N_7293,N_863,N_4586);
and U7294 (N_7294,N_226,N_2215);
or U7295 (N_7295,N_1068,N_2345);
nor U7296 (N_7296,N_2026,N_1750);
and U7297 (N_7297,N_4313,N_3919);
and U7298 (N_7298,N_881,N_4080);
and U7299 (N_7299,N_2447,N_2553);
or U7300 (N_7300,N_1130,N_4329);
or U7301 (N_7301,N_3384,N_3736);
and U7302 (N_7302,N_1764,N_4677);
nor U7303 (N_7303,N_2897,N_2753);
nor U7304 (N_7304,N_1425,N_120);
or U7305 (N_7305,N_4332,N_199);
or U7306 (N_7306,N_4914,N_3644);
nand U7307 (N_7307,N_3167,N_2078);
or U7308 (N_7308,N_2609,N_2629);
nor U7309 (N_7309,N_981,N_2934);
nand U7310 (N_7310,N_1985,N_1657);
nand U7311 (N_7311,N_4907,N_3597);
or U7312 (N_7312,N_3701,N_3840);
or U7313 (N_7313,N_685,N_1561);
and U7314 (N_7314,N_1601,N_921);
nor U7315 (N_7315,N_1400,N_841);
or U7316 (N_7316,N_3447,N_37);
or U7317 (N_7317,N_2299,N_4249);
and U7318 (N_7318,N_4395,N_2823);
nor U7319 (N_7319,N_2893,N_4385);
and U7320 (N_7320,N_4,N_73);
and U7321 (N_7321,N_1602,N_258);
nor U7322 (N_7322,N_3877,N_1965);
nor U7323 (N_7323,N_1749,N_542);
and U7324 (N_7324,N_3995,N_185);
nor U7325 (N_7325,N_1999,N_4368);
nand U7326 (N_7326,N_2332,N_4863);
nand U7327 (N_7327,N_1371,N_4651);
nor U7328 (N_7328,N_2762,N_1449);
or U7329 (N_7329,N_1813,N_1318);
and U7330 (N_7330,N_4982,N_3452);
and U7331 (N_7331,N_2846,N_1694);
nand U7332 (N_7332,N_4106,N_235);
nor U7333 (N_7333,N_3807,N_3150);
and U7334 (N_7334,N_2202,N_3542);
or U7335 (N_7335,N_4497,N_1157);
nor U7336 (N_7336,N_821,N_1021);
nand U7337 (N_7337,N_2935,N_1960);
and U7338 (N_7338,N_2817,N_1146);
or U7339 (N_7339,N_3304,N_4335);
and U7340 (N_7340,N_296,N_866);
nor U7341 (N_7341,N_4816,N_4327);
and U7342 (N_7342,N_4801,N_4565);
and U7343 (N_7343,N_4885,N_535);
xor U7344 (N_7344,N_698,N_4538);
or U7345 (N_7345,N_3093,N_2995);
and U7346 (N_7346,N_224,N_1143);
or U7347 (N_7347,N_4684,N_52);
nand U7348 (N_7348,N_2152,N_2088);
nand U7349 (N_7349,N_899,N_4506);
or U7350 (N_7350,N_2843,N_3302);
nand U7351 (N_7351,N_483,N_3034);
nand U7352 (N_7352,N_1208,N_3173);
nor U7353 (N_7353,N_2232,N_2467);
nand U7354 (N_7354,N_4489,N_241);
or U7355 (N_7355,N_4613,N_1931);
nand U7356 (N_7356,N_2712,N_154);
nand U7357 (N_7357,N_967,N_1516);
and U7358 (N_7358,N_1128,N_4547);
nand U7359 (N_7359,N_4471,N_1176);
nand U7360 (N_7360,N_4245,N_4144);
and U7361 (N_7361,N_3387,N_434);
or U7362 (N_7362,N_1437,N_2798);
nand U7363 (N_7363,N_1280,N_4465);
nor U7364 (N_7364,N_218,N_91);
or U7365 (N_7365,N_4647,N_642);
or U7366 (N_7366,N_974,N_2972);
nor U7367 (N_7367,N_3884,N_3318);
nor U7368 (N_7368,N_781,N_4872);
nor U7369 (N_7369,N_4103,N_4495);
or U7370 (N_7370,N_1920,N_420);
nand U7371 (N_7371,N_4597,N_4483);
or U7372 (N_7372,N_4242,N_4527);
nand U7373 (N_7373,N_1246,N_2193);
nand U7374 (N_7374,N_3595,N_2779);
nor U7375 (N_7375,N_4479,N_1885);
nand U7376 (N_7376,N_2032,N_544);
or U7377 (N_7377,N_4628,N_1638);
nand U7378 (N_7378,N_3129,N_4930);
nor U7379 (N_7379,N_609,N_4340);
nor U7380 (N_7380,N_2401,N_2432);
or U7381 (N_7381,N_3650,N_3419);
nand U7382 (N_7382,N_1174,N_209);
and U7383 (N_7383,N_534,N_2839);
nand U7384 (N_7384,N_691,N_2131);
or U7385 (N_7385,N_1414,N_3159);
or U7386 (N_7386,N_4760,N_1138);
nand U7387 (N_7387,N_2983,N_1566);
nand U7388 (N_7388,N_2166,N_3829);
and U7389 (N_7389,N_2257,N_1839);
nand U7390 (N_7390,N_1684,N_3252);
nor U7391 (N_7391,N_4725,N_1315);
nand U7392 (N_7392,N_2737,N_1758);
nand U7393 (N_7393,N_4689,N_3233);
or U7394 (N_7394,N_1614,N_1878);
and U7395 (N_7395,N_669,N_3556);
or U7396 (N_7396,N_85,N_3068);
and U7397 (N_7397,N_854,N_693);
or U7398 (N_7398,N_2009,N_2462);
and U7399 (N_7399,N_2784,N_3003);
or U7400 (N_7400,N_2605,N_1761);
and U7401 (N_7401,N_2511,N_108);
and U7402 (N_7402,N_2919,N_3362);
nand U7403 (N_7403,N_1091,N_3622);
or U7404 (N_7404,N_3228,N_4704);
or U7405 (N_7405,N_1814,N_2439);
and U7406 (N_7406,N_484,N_324);
nand U7407 (N_7407,N_1040,N_2916);
nand U7408 (N_7408,N_2425,N_3016);
nand U7409 (N_7409,N_4481,N_990);
or U7410 (N_7410,N_4637,N_1497);
nor U7411 (N_7411,N_3538,N_1012);
nand U7412 (N_7412,N_4228,N_435);
nand U7413 (N_7413,N_1071,N_1291);
and U7414 (N_7414,N_4220,N_4663);
nor U7415 (N_7415,N_2021,N_4629);
and U7416 (N_7416,N_4134,N_2636);
or U7417 (N_7417,N_1353,N_3131);
and U7418 (N_7418,N_3038,N_3245);
or U7419 (N_7419,N_78,N_65);
or U7420 (N_7420,N_3274,N_4352);
nor U7421 (N_7421,N_4542,N_817);
and U7422 (N_7422,N_4894,N_2170);
nor U7423 (N_7423,N_2703,N_2772);
or U7424 (N_7424,N_2955,N_486);
or U7425 (N_7425,N_3725,N_2492);
nor U7426 (N_7426,N_890,N_1336);
nand U7427 (N_7427,N_989,N_3465);
nor U7428 (N_7428,N_3366,N_4844);
and U7429 (N_7429,N_864,N_1288);
or U7430 (N_7430,N_3721,N_4406);
nor U7431 (N_7431,N_3095,N_3018);
and U7432 (N_7432,N_1069,N_2240);
nand U7433 (N_7433,N_4955,N_1670);
or U7434 (N_7434,N_3768,N_4661);
and U7435 (N_7435,N_3922,N_4464);
nor U7436 (N_7436,N_3797,N_2025);
nor U7437 (N_7437,N_4084,N_495);
and U7438 (N_7438,N_4432,N_2449);
or U7439 (N_7439,N_1628,N_4253);
nand U7440 (N_7440,N_2273,N_1681);
and U7441 (N_7441,N_1003,N_2461);
nand U7442 (N_7442,N_2143,N_4806);
nand U7443 (N_7443,N_3575,N_3806);
nand U7444 (N_7444,N_3478,N_3461);
and U7445 (N_7445,N_4817,N_3029);
nor U7446 (N_7446,N_3406,N_1988);
nand U7447 (N_7447,N_1019,N_510);
or U7448 (N_7448,N_634,N_3296);
and U7449 (N_7449,N_3704,N_1079);
nand U7450 (N_7450,N_3100,N_174);
or U7451 (N_7451,N_4921,N_462);
nand U7452 (N_7452,N_2272,N_2871);
nand U7453 (N_7453,N_260,N_48);
or U7454 (N_7454,N_3249,N_1381);
and U7455 (N_7455,N_4993,N_3860);
and U7456 (N_7456,N_1682,N_2729);
and U7457 (N_7457,N_566,N_607);
and U7458 (N_7458,N_2344,N_2296);
or U7459 (N_7459,N_4128,N_3225);
nor U7460 (N_7460,N_1806,N_10);
nand U7461 (N_7461,N_2748,N_3576);
and U7462 (N_7462,N_3373,N_2582);
nor U7463 (N_7463,N_4525,N_1726);
nor U7464 (N_7464,N_4303,N_3518);
or U7465 (N_7465,N_449,N_2211);
or U7466 (N_7466,N_1633,N_4058);
nor U7467 (N_7467,N_577,N_100);
nand U7468 (N_7468,N_1419,N_931);
nor U7469 (N_7469,N_1250,N_3206);
nor U7470 (N_7470,N_1120,N_3646);
or U7471 (N_7471,N_1245,N_2018);
nand U7472 (N_7472,N_2612,N_197);
nor U7473 (N_7473,N_3393,N_3525);
nand U7474 (N_7474,N_213,N_1510);
nand U7475 (N_7475,N_2631,N_4593);
and U7476 (N_7476,N_2583,N_1578);
or U7477 (N_7477,N_115,N_4555);
nor U7478 (N_7478,N_1956,N_1312);
nor U7479 (N_7479,N_1330,N_1016);
nor U7480 (N_7480,N_2338,N_2331);
nand U7481 (N_7481,N_466,N_4824);
and U7482 (N_7482,N_847,N_4719);
or U7483 (N_7483,N_1844,N_926);
and U7484 (N_7484,N_592,N_1490);
and U7485 (N_7485,N_1169,N_3640);
nand U7486 (N_7486,N_4297,N_4695);
and U7487 (N_7487,N_2988,N_2952);
nor U7488 (N_7488,N_2481,N_4600);
or U7489 (N_7489,N_2752,N_877);
and U7490 (N_7490,N_4905,N_522);
and U7491 (N_7491,N_3777,N_1453);
or U7492 (N_7492,N_4209,N_4792);
nor U7493 (N_7493,N_1987,N_3687);
nor U7494 (N_7494,N_2126,N_3657);
nor U7495 (N_7495,N_4788,N_1784);
nand U7496 (N_7496,N_1707,N_1847);
or U7497 (N_7497,N_2854,N_2424);
nor U7498 (N_7498,N_2727,N_195);
or U7499 (N_7499,N_2353,N_2654);
and U7500 (N_7500,N_3827,N_158);
nor U7501 (N_7501,N_1591,N_4632);
nor U7502 (N_7502,N_4843,N_1526);
or U7503 (N_7503,N_3235,N_2703);
or U7504 (N_7504,N_380,N_4108);
and U7505 (N_7505,N_3337,N_3224);
nand U7506 (N_7506,N_3769,N_4615);
nor U7507 (N_7507,N_582,N_1018);
or U7508 (N_7508,N_2579,N_1274);
nor U7509 (N_7509,N_43,N_1745);
nor U7510 (N_7510,N_4198,N_4297);
nand U7511 (N_7511,N_3199,N_325);
nand U7512 (N_7512,N_1253,N_3202);
and U7513 (N_7513,N_4284,N_2213);
or U7514 (N_7514,N_3114,N_1702);
nand U7515 (N_7515,N_2144,N_4669);
nand U7516 (N_7516,N_2876,N_4501);
nor U7517 (N_7517,N_1397,N_3238);
or U7518 (N_7518,N_168,N_4024);
nor U7519 (N_7519,N_3687,N_4912);
nand U7520 (N_7520,N_1263,N_2598);
nand U7521 (N_7521,N_2866,N_3010);
nor U7522 (N_7522,N_1717,N_1841);
or U7523 (N_7523,N_2594,N_40);
or U7524 (N_7524,N_4316,N_82);
or U7525 (N_7525,N_1888,N_3440);
nor U7526 (N_7526,N_1039,N_4584);
and U7527 (N_7527,N_438,N_1437);
nor U7528 (N_7528,N_3285,N_4168);
nand U7529 (N_7529,N_4643,N_3625);
nand U7530 (N_7530,N_1137,N_2961);
and U7531 (N_7531,N_1281,N_488);
and U7532 (N_7532,N_2058,N_148);
and U7533 (N_7533,N_155,N_1498);
or U7534 (N_7534,N_1725,N_3776);
nand U7535 (N_7535,N_306,N_2969);
or U7536 (N_7536,N_3478,N_1594);
nand U7537 (N_7537,N_4440,N_1633);
and U7538 (N_7538,N_1131,N_4604);
nor U7539 (N_7539,N_657,N_1584);
or U7540 (N_7540,N_3005,N_884);
nor U7541 (N_7541,N_2232,N_4502);
nor U7542 (N_7542,N_3741,N_398);
nand U7543 (N_7543,N_2905,N_4852);
nor U7544 (N_7544,N_2621,N_2144);
nor U7545 (N_7545,N_2476,N_3385);
nor U7546 (N_7546,N_3548,N_3425);
nand U7547 (N_7547,N_3963,N_4180);
and U7548 (N_7548,N_4194,N_283);
nand U7549 (N_7549,N_121,N_4421);
nand U7550 (N_7550,N_1012,N_444);
and U7551 (N_7551,N_533,N_3342);
nor U7552 (N_7552,N_794,N_3315);
or U7553 (N_7553,N_2895,N_4699);
nor U7554 (N_7554,N_2943,N_2476);
nor U7555 (N_7555,N_4885,N_2682);
nand U7556 (N_7556,N_2237,N_3063);
or U7557 (N_7557,N_2141,N_2440);
nor U7558 (N_7558,N_4039,N_379);
or U7559 (N_7559,N_3978,N_2133);
and U7560 (N_7560,N_3286,N_2925);
and U7561 (N_7561,N_584,N_210);
or U7562 (N_7562,N_3578,N_3831);
nor U7563 (N_7563,N_4580,N_44);
or U7564 (N_7564,N_1780,N_247);
nor U7565 (N_7565,N_2892,N_3663);
nor U7566 (N_7566,N_269,N_2474);
nand U7567 (N_7567,N_1465,N_1827);
or U7568 (N_7568,N_170,N_1771);
nor U7569 (N_7569,N_4761,N_2339);
or U7570 (N_7570,N_3210,N_3316);
or U7571 (N_7571,N_2390,N_960);
and U7572 (N_7572,N_1235,N_1053);
nand U7573 (N_7573,N_4020,N_2299);
and U7574 (N_7574,N_1749,N_3433);
or U7575 (N_7575,N_1556,N_3313);
nor U7576 (N_7576,N_973,N_1296);
nand U7577 (N_7577,N_2381,N_137);
or U7578 (N_7578,N_4238,N_77);
nand U7579 (N_7579,N_2892,N_2033);
nor U7580 (N_7580,N_1587,N_2556);
and U7581 (N_7581,N_1359,N_4294);
and U7582 (N_7582,N_504,N_2241);
or U7583 (N_7583,N_4144,N_2091);
nor U7584 (N_7584,N_470,N_2154);
and U7585 (N_7585,N_793,N_3163);
nor U7586 (N_7586,N_424,N_993);
nand U7587 (N_7587,N_3116,N_4054);
nand U7588 (N_7588,N_311,N_2022);
nand U7589 (N_7589,N_553,N_2357);
and U7590 (N_7590,N_109,N_1132);
or U7591 (N_7591,N_381,N_3729);
xnor U7592 (N_7592,N_3404,N_2958);
and U7593 (N_7593,N_4035,N_2438);
or U7594 (N_7594,N_2553,N_1476);
nand U7595 (N_7595,N_2114,N_819);
and U7596 (N_7596,N_4462,N_3074);
or U7597 (N_7597,N_3491,N_2912);
nand U7598 (N_7598,N_3321,N_4053);
nand U7599 (N_7599,N_3575,N_1116);
or U7600 (N_7600,N_1137,N_3380);
xnor U7601 (N_7601,N_1531,N_3817);
or U7602 (N_7602,N_120,N_2215);
nand U7603 (N_7603,N_881,N_1773);
or U7604 (N_7604,N_852,N_2391);
or U7605 (N_7605,N_3768,N_1833);
nand U7606 (N_7606,N_2878,N_4665);
and U7607 (N_7607,N_1459,N_844);
nand U7608 (N_7608,N_4118,N_4622);
and U7609 (N_7609,N_1575,N_4743);
or U7610 (N_7610,N_4375,N_93);
nor U7611 (N_7611,N_3606,N_4606);
nor U7612 (N_7612,N_3336,N_4500);
nor U7613 (N_7613,N_4876,N_1247);
nor U7614 (N_7614,N_1028,N_2273);
nand U7615 (N_7615,N_1105,N_3721);
nor U7616 (N_7616,N_396,N_3951);
nand U7617 (N_7617,N_178,N_2701);
or U7618 (N_7618,N_3604,N_4629);
nor U7619 (N_7619,N_2703,N_4175);
and U7620 (N_7620,N_4962,N_2721);
and U7621 (N_7621,N_1605,N_1582);
and U7622 (N_7622,N_2731,N_258);
nand U7623 (N_7623,N_3685,N_2156);
nand U7624 (N_7624,N_1154,N_918);
or U7625 (N_7625,N_4218,N_4358);
nand U7626 (N_7626,N_2332,N_1329);
nor U7627 (N_7627,N_3521,N_4200);
or U7628 (N_7628,N_1883,N_797);
nand U7629 (N_7629,N_4713,N_2547);
and U7630 (N_7630,N_3455,N_514);
and U7631 (N_7631,N_1093,N_2514);
nand U7632 (N_7632,N_180,N_2970);
and U7633 (N_7633,N_3601,N_415);
nor U7634 (N_7634,N_1198,N_3170);
and U7635 (N_7635,N_2401,N_2624);
or U7636 (N_7636,N_3607,N_628);
nor U7637 (N_7637,N_25,N_1816);
and U7638 (N_7638,N_2702,N_2042);
nand U7639 (N_7639,N_136,N_2608);
nand U7640 (N_7640,N_1113,N_4500);
or U7641 (N_7641,N_4186,N_3644);
nand U7642 (N_7642,N_1511,N_1266);
nand U7643 (N_7643,N_4297,N_1833);
and U7644 (N_7644,N_3965,N_3721);
and U7645 (N_7645,N_1709,N_1719);
nand U7646 (N_7646,N_873,N_1816);
nand U7647 (N_7647,N_3098,N_725);
nand U7648 (N_7648,N_214,N_1985);
nand U7649 (N_7649,N_1074,N_4604);
nand U7650 (N_7650,N_878,N_4741);
nand U7651 (N_7651,N_2033,N_958);
nor U7652 (N_7652,N_414,N_3016);
nor U7653 (N_7653,N_657,N_3917);
nor U7654 (N_7654,N_3848,N_508);
and U7655 (N_7655,N_520,N_4927);
nand U7656 (N_7656,N_124,N_597);
or U7657 (N_7657,N_4900,N_4701);
and U7658 (N_7658,N_3028,N_2250);
or U7659 (N_7659,N_2592,N_149);
nor U7660 (N_7660,N_2271,N_4224);
nor U7661 (N_7661,N_1895,N_4640);
and U7662 (N_7662,N_1434,N_4910);
and U7663 (N_7663,N_3688,N_1124);
or U7664 (N_7664,N_1820,N_1431);
or U7665 (N_7665,N_4184,N_1767);
or U7666 (N_7666,N_1465,N_3067);
nand U7667 (N_7667,N_4879,N_2302);
or U7668 (N_7668,N_2121,N_237);
nand U7669 (N_7669,N_833,N_2479);
nor U7670 (N_7670,N_833,N_718);
or U7671 (N_7671,N_1022,N_4946);
nand U7672 (N_7672,N_4136,N_966);
and U7673 (N_7673,N_870,N_4590);
or U7674 (N_7674,N_597,N_4392);
or U7675 (N_7675,N_2179,N_939);
nand U7676 (N_7676,N_2825,N_1742);
nand U7677 (N_7677,N_3802,N_4129);
and U7678 (N_7678,N_895,N_4261);
and U7679 (N_7679,N_2863,N_3128);
nor U7680 (N_7680,N_1870,N_4419);
nand U7681 (N_7681,N_677,N_4905);
or U7682 (N_7682,N_4244,N_3372);
and U7683 (N_7683,N_1604,N_3187);
or U7684 (N_7684,N_1305,N_4223);
nor U7685 (N_7685,N_302,N_3793);
nor U7686 (N_7686,N_1863,N_4523);
or U7687 (N_7687,N_816,N_130);
nor U7688 (N_7688,N_2070,N_3621);
or U7689 (N_7689,N_2835,N_2526);
or U7690 (N_7690,N_4810,N_1075);
or U7691 (N_7691,N_2321,N_2026);
nor U7692 (N_7692,N_3024,N_862);
and U7693 (N_7693,N_2867,N_500);
nor U7694 (N_7694,N_1828,N_190);
nor U7695 (N_7695,N_1877,N_423);
and U7696 (N_7696,N_950,N_710);
and U7697 (N_7697,N_2664,N_3268);
and U7698 (N_7698,N_999,N_3341);
nor U7699 (N_7699,N_998,N_389);
and U7700 (N_7700,N_3008,N_316);
or U7701 (N_7701,N_2973,N_1501);
or U7702 (N_7702,N_1815,N_660);
and U7703 (N_7703,N_3064,N_4264);
nand U7704 (N_7704,N_3814,N_4377);
nor U7705 (N_7705,N_2193,N_2306);
nand U7706 (N_7706,N_3053,N_3067);
nand U7707 (N_7707,N_3316,N_3773);
nor U7708 (N_7708,N_2993,N_2805);
nand U7709 (N_7709,N_4519,N_4479);
nand U7710 (N_7710,N_1307,N_4323);
or U7711 (N_7711,N_1343,N_3618);
nand U7712 (N_7712,N_3804,N_2071);
or U7713 (N_7713,N_4438,N_3208);
nand U7714 (N_7714,N_4950,N_3067);
and U7715 (N_7715,N_2127,N_4066);
nor U7716 (N_7716,N_4143,N_3584);
nand U7717 (N_7717,N_873,N_1908);
nand U7718 (N_7718,N_845,N_4380);
nor U7719 (N_7719,N_3124,N_2304);
or U7720 (N_7720,N_3126,N_2502);
nand U7721 (N_7721,N_2460,N_3020);
and U7722 (N_7722,N_1155,N_512);
and U7723 (N_7723,N_898,N_1647);
nor U7724 (N_7724,N_3744,N_3069);
or U7725 (N_7725,N_1489,N_4852);
nand U7726 (N_7726,N_2103,N_772);
nor U7727 (N_7727,N_3190,N_3044);
nand U7728 (N_7728,N_285,N_933);
nand U7729 (N_7729,N_3579,N_2500);
nand U7730 (N_7730,N_161,N_4955);
nand U7731 (N_7731,N_2441,N_2689);
nand U7732 (N_7732,N_120,N_4943);
nand U7733 (N_7733,N_449,N_2077);
or U7734 (N_7734,N_3141,N_616);
nand U7735 (N_7735,N_4842,N_2584);
nor U7736 (N_7736,N_1784,N_4699);
nand U7737 (N_7737,N_3325,N_4248);
nand U7738 (N_7738,N_3846,N_4332);
nor U7739 (N_7739,N_4272,N_4079);
and U7740 (N_7740,N_1960,N_2860);
or U7741 (N_7741,N_1486,N_311);
and U7742 (N_7742,N_89,N_3242);
nor U7743 (N_7743,N_4048,N_3684);
nand U7744 (N_7744,N_2196,N_920);
or U7745 (N_7745,N_3124,N_2729);
nor U7746 (N_7746,N_3957,N_1982);
or U7747 (N_7747,N_567,N_4954);
nor U7748 (N_7748,N_1598,N_519);
nor U7749 (N_7749,N_136,N_3459);
nor U7750 (N_7750,N_593,N_855);
nand U7751 (N_7751,N_4664,N_4345);
nand U7752 (N_7752,N_4507,N_3052);
or U7753 (N_7753,N_3976,N_1348);
and U7754 (N_7754,N_1538,N_642);
nand U7755 (N_7755,N_792,N_4926);
and U7756 (N_7756,N_4714,N_2758);
or U7757 (N_7757,N_2239,N_658);
or U7758 (N_7758,N_3086,N_1606);
or U7759 (N_7759,N_687,N_976);
and U7760 (N_7760,N_2491,N_3541);
and U7761 (N_7761,N_4194,N_2404);
nand U7762 (N_7762,N_2252,N_2720);
or U7763 (N_7763,N_3289,N_2897);
or U7764 (N_7764,N_893,N_2444);
and U7765 (N_7765,N_1520,N_2443);
nor U7766 (N_7766,N_2384,N_3014);
or U7767 (N_7767,N_4345,N_4237);
nand U7768 (N_7768,N_4428,N_2002);
nand U7769 (N_7769,N_595,N_3318);
nand U7770 (N_7770,N_3143,N_1580);
nor U7771 (N_7771,N_3561,N_3210);
and U7772 (N_7772,N_4652,N_3598);
nand U7773 (N_7773,N_1627,N_4269);
or U7774 (N_7774,N_1279,N_3017);
and U7775 (N_7775,N_896,N_4188);
or U7776 (N_7776,N_34,N_4357);
nand U7777 (N_7777,N_3733,N_2724);
xnor U7778 (N_7778,N_1199,N_4023);
nand U7779 (N_7779,N_2142,N_3711);
nor U7780 (N_7780,N_2171,N_4422);
or U7781 (N_7781,N_28,N_4554);
nor U7782 (N_7782,N_2586,N_2140);
or U7783 (N_7783,N_436,N_1489);
or U7784 (N_7784,N_4716,N_2860);
and U7785 (N_7785,N_110,N_3652);
nor U7786 (N_7786,N_762,N_1856);
nand U7787 (N_7787,N_3182,N_1806);
nor U7788 (N_7788,N_1872,N_1880);
nor U7789 (N_7789,N_1896,N_2284);
nand U7790 (N_7790,N_3665,N_853);
and U7791 (N_7791,N_3047,N_448);
nand U7792 (N_7792,N_516,N_2860);
nor U7793 (N_7793,N_2852,N_2900);
or U7794 (N_7794,N_670,N_295);
or U7795 (N_7795,N_112,N_1904);
and U7796 (N_7796,N_4969,N_2858);
and U7797 (N_7797,N_1192,N_3796);
or U7798 (N_7798,N_2750,N_2999);
nor U7799 (N_7799,N_3731,N_156);
and U7800 (N_7800,N_3003,N_851);
and U7801 (N_7801,N_2401,N_3802);
or U7802 (N_7802,N_3138,N_1085);
and U7803 (N_7803,N_4907,N_624);
nand U7804 (N_7804,N_2610,N_367);
nand U7805 (N_7805,N_2624,N_794);
or U7806 (N_7806,N_91,N_1595);
and U7807 (N_7807,N_2006,N_3865);
and U7808 (N_7808,N_4757,N_1776);
or U7809 (N_7809,N_2965,N_119);
or U7810 (N_7810,N_3342,N_3650);
and U7811 (N_7811,N_3332,N_3076);
and U7812 (N_7812,N_2266,N_3062);
and U7813 (N_7813,N_2370,N_1503);
nor U7814 (N_7814,N_4993,N_2883);
or U7815 (N_7815,N_1132,N_2706);
or U7816 (N_7816,N_146,N_921);
or U7817 (N_7817,N_1352,N_1568);
nor U7818 (N_7818,N_1284,N_4135);
nor U7819 (N_7819,N_2727,N_2472);
nor U7820 (N_7820,N_277,N_4509);
nor U7821 (N_7821,N_2519,N_4203);
and U7822 (N_7822,N_3454,N_5);
nand U7823 (N_7823,N_1512,N_4088);
nand U7824 (N_7824,N_3167,N_2780);
nand U7825 (N_7825,N_300,N_3383);
nand U7826 (N_7826,N_1660,N_856);
nor U7827 (N_7827,N_3654,N_919);
and U7828 (N_7828,N_3360,N_660);
and U7829 (N_7829,N_3530,N_324);
or U7830 (N_7830,N_1616,N_2418);
nor U7831 (N_7831,N_2870,N_2737);
nand U7832 (N_7832,N_2668,N_645);
or U7833 (N_7833,N_4626,N_827);
nor U7834 (N_7834,N_4499,N_73);
nor U7835 (N_7835,N_3655,N_2707);
or U7836 (N_7836,N_1624,N_2467);
and U7837 (N_7837,N_3661,N_3104);
nor U7838 (N_7838,N_1593,N_182);
nor U7839 (N_7839,N_69,N_754);
or U7840 (N_7840,N_3045,N_3727);
or U7841 (N_7841,N_177,N_1649);
nand U7842 (N_7842,N_1354,N_4198);
nor U7843 (N_7843,N_4256,N_266);
or U7844 (N_7844,N_4852,N_3434);
nor U7845 (N_7845,N_4210,N_3161);
and U7846 (N_7846,N_3471,N_3);
or U7847 (N_7847,N_830,N_2500);
or U7848 (N_7848,N_1163,N_638);
and U7849 (N_7849,N_373,N_1464);
and U7850 (N_7850,N_2740,N_3344);
nand U7851 (N_7851,N_3139,N_1970);
or U7852 (N_7852,N_4927,N_2951);
or U7853 (N_7853,N_4993,N_3334);
and U7854 (N_7854,N_3496,N_4993);
nand U7855 (N_7855,N_3541,N_4812);
nand U7856 (N_7856,N_4833,N_4168);
and U7857 (N_7857,N_3918,N_4680);
or U7858 (N_7858,N_4952,N_4850);
or U7859 (N_7859,N_3559,N_2747);
nand U7860 (N_7860,N_838,N_4025);
and U7861 (N_7861,N_4057,N_2750);
and U7862 (N_7862,N_2524,N_4790);
nor U7863 (N_7863,N_1557,N_1347);
and U7864 (N_7864,N_3703,N_2971);
nor U7865 (N_7865,N_3935,N_2445);
nand U7866 (N_7866,N_1353,N_2488);
and U7867 (N_7867,N_3287,N_3156);
nor U7868 (N_7868,N_2942,N_3453);
nand U7869 (N_7869,N_4701,N_4751);
nand U7870 (N_7870,N_616,N_4972);
nand U7871 (N_7871,N_2699,N_4793);
or U7872 (N_7872,N_2360,N_3166);
nand U7873 (N_7873,N_653,N_4721);
nor U7874 (N_7874,N_968,N_1931);
nor U7875 (N_7875,N_967,N_271);
nand U7876 (N_7876,N_1361,N_1509);
nand U7877 (N_7877,N_442,N_1985);
nor U7878 (N_7878,N_3413,N_2014);
and U7879 (N_7879,N_3055,N_1189);
xnor U7880 (N_7880,N_2450,N_2004);
nor U7881 (N_7881,N_3955,N_3165);
nand U7882 (N_7882,N_1689,N_787);
or U7883 (N_7883,N_4242,N_2593);
and U7884 (N_7884,N_1921,N_1916);
or U7885 (N_7885,N_4556,N_2207);
and U7886 (N_7886,N_2268,N_762);
or U7887 (N_7887,N_463,N_4138);
and U7888 (N_7888,N_539,N_2804);
and U7889 (N_7889,N_321,N_1787);
nand U7890 (N_7890,N_3732,N_1576);
or U7891 (N_7891,N_236,N_4450);
and U7892 (N_7892,N_4916,N_2822);
or U7893 (N_7893,N_666,N_1809);
or U7894 (N_7894,N_3856,N_1004);
nor U7895 (N_7895,N_2279,N_3678);
or U7896 (N_7896,N_3005,N_435);
nor U7897 (N_7897,N_3091,N_2921);
xor U7898 (N_7898,N_2964,N_1181);
or U7899 (N_7899,N_2796,N_2347);
nand U7900 (N_7900,N_1665,N_481);
nand U7901 (N_7901,N_3040,N_1542);
nand U7902 (N_7902,N_4290,N_4577);
nand U7903 (N_7903,N_1621,N_4835);
or U7904 (N_7904,N_1033,N_1711);
nand U7905 (N_7905,N_4674,N_957);
nor U7906 (N_7906,N_4561,N_4307);
nor U7907 (N_7907,N_1611,N_2727);
or U7908 (N_7908,N_3903,N_1142);
and U7909 (N_7909,N_1089,N_2106);
and U7910 (N_7910,N_3943,N_2645);
or U7911 (N_7911,N_4690,N_3120);
nor U7912 (N_7912,N_2296,N_2774);
nor U7913 (N_7913,N_305,N_959);
or U7914 (N_7914,N_569,N_2008);
and U7915 (N_7915,N_942,N_4592);
or U7916 (N_7916,N_2460,N_1428);
and U7917 (N_7917,N_4248,N_696);
or U7918 (N_7918,N_63,N_1429);
and U7919 (N_7919,N_605,N_3930);
and U7920 (N_7920,N_4046,N_2862);
and U7921 (N_7921,N_402,N_3225);
nor U7922 (N_7922,N_800,N_4151);
nand U7923 (N_7923,N_2754,N_4350);
nor U7924 (N_7924,N_1895,N_3748);
or U7925 (N_7925,N_2273,N_4042);
nand U7926 (N_7926,N_2295,N_831);
nand U7927 (N_7927,N_3207,N_3650);
nor U7928 (N_7928,N_4565,N_2668);
or U7929 (N_7929,N_1721,N_169);
and U7930 (N_7930,N_2890,N_1426);
nand U7931 (N_7931,N_3127,N_3109);
or U7932 (N_7932,N_2005,N_2020);
nor U7933 (N_7933,N_838,N_3911);
nand U7934 (N_7934,N_2885,N_3463);
nand U7935 (N_7935,N_790,N_4938);
and U7936 (N_7936,N_4932,N_649);
or U7937 (N_7937,N_1669,N_2971);
nand U7938 (N_7938,N_2818,N_808);
or U7939 (N_7939,N_4497,N_1465);
nand U7940 (N_7940,N_1915,N_1941);
nor U7941 (N_7941,N_3332,N_148);
and U7942 (N_7942,N_1579,N_3496);
xnor U7943 (N_7943,N_2940,N_4063);
nand U7944 (N_7944,N_873,N_1864);
nor U7945 (N_7945,N_818,N_3458);
nor U7946 (N_7946,N_3405,N_555);
nand U7947 (N_7947,N_1405,N_4979);
and U7948 (N_7948,N_1081,N_3448);
nor U7949 (N_7949,N_3770,N_1497);
and U7950 (N_7950,N_2735,N_2505);
nor U7951 (N_7951,N_3109,N_1661);
and U7952 (N_7952,N_4173,N_240);
or U7953 (N_7953,N_776,N_1123);
nor U7954 (N_7954,N_1857,N_732);
nor U7955 (N_7955,N_4326,N_3902);
or U7956 (N_7956,N_3306,N_1463);
and U7957 (N_7957,N_3375,N_542);
or U7958 (N_7958,N_363,N_3426);
nor U7959 (N_7959,N_2881,N_838);
nand U7960 (N_7960,N_1705,N_977);
and U7961 (N_7961,N_4747,N_768);
nor U7962 (N_7962,N_1462,N_4446);
xor U7963 (N_7963,N_1025,N_2534);
xor U7964 (N_7964,N_993,N_2413);
nor U7965 (N_7965,N_2026,N_2953);
or U7966 (N_7966,N_3275,N_4585);
or U7967 (N_7967,N_4336,N_2217);
nand U7968 (N_7968,N_2473,N_4628);
and U7969 (N_7969,N_4760,N_4912);
nor U7970 (N_7970,N_925,N_1500);
nand U7971 (N_7971,N_4956,N_2980);
or U7972 (N_7972,N_876,N_1023);
nand U7973 (N_7973,N_3942,N_4852);
or U7974 (N_7974,N_1341,N_3918);
or U7975 (N_7975,N_1413,N_1086);
or U7976 (N_7976,N_773,N_3281);
nor U7977 (N_7977,N_2875,N_4503);
nor U7978 (N_7978,N_2803,N_2809);
and U7979 (N_7979,N_3236,N_1884);
nor U7980 (N_7980,N_4978,N_3502);
and U7981 (N_7981,N_4132,N_3015);
nor U7982 (N_7982,N_568,N_904);
and U7983 (N_7983,N_4031,N_3675);
or U7984 (N_7984,N_4973,N_1782);
nor U7985 (N_7985,N_1540,N_1520);
nand U7986 (N_7986,N_1197,N_2699);
nand U7987 (N_7987,N_3447,N_3143);
nand U7988 (N_7988,N_2965,N_3889);
nor U7989 (N_7989,N_3718,N_2409);
nor U7990 (N_7990,N_4168,N_4487);
and U7991 (N_7991,N_101,N_3734);
and U7992 (N_7992,N_2316,N_1039);
or U7993 (N_7993,N_609,N_1488);
nand U7994 (N_7994,N_3445,N_549);
and U7995 (N_7995,N_3645,N_588);
or U7996 (N_7996,N_4938,N_4082);
nor U7997 (N_7997,N_2589,N_2897);
and U7998 (N_7998,N_4592,N_3887);
nor U7999 (N_7999,N_2634,N_4752);
or U8000 (N_8000,N_2939,N_4956);
or U8001 (N_8001,N_4879,N_3975);
or U8002 (N_8002,N_3308,N_2623);
nand U8003 (N_8003,N_3567,N_3742);
nor U8004 (N_8004,N_2066,N_1362);
nor U8005 (N_8005,N_3803,N_3978);
or U8006 (N_8006,N_2748,N_651);
nor U8007 (N_8007,N_3619,N_189);
and U8008 (N_8008,N_441,N_4488);
or U8009 (N_8009,N_2126,N_684);
xor U8010 (N_8010,N_2324,N_2128);
and U8011 (N_8011,N_3159,N_3612);
xor U8012 (N_8012,N_2330,N_505);
or U8013 (N_8013,N_511,N_3947);
nor U8014 (N_8014,N_3076,N_3176);
nor U8015 (N_8015,N_3513,N_990);
nand U8016 (N_8016,N_2618,N_2437);
or U8017 (N_8017,N_3328,N_1113);
or U8018 (N_8018,N_2803,N_314);
and U8019 (N_8019,N_4540,N_3883);
xnor U8020 (N_8020,N_2166,N_3056);
nor U8021 (N_8021,N_2892,N_3195);
or U8022 (N_8022,N_3233,N_1491);
or U8023 (N_8023,N_2592,N_1487);
nor U8024 (N_8024,N_4503,N_1252);
or U8025 (N_8025,N_2755,N_359);
or U8026 (N_8026,N_3573,N_3269);
and U8027 (N_8027,N_2906,N_921);
and U8028 (N_8028,N_2559,N_3691);
nand U8029 (N_8029,N_847,N_135);
nor U8030 (N_8030,N_3720,N_2532);
and U8031 (N_8031,N_4723,N_4641);
or U8032 (N_8032,N_84,N_2680);
xor U8033 (N_8033,N_3056,N_4513);
and U8034 (N_8034,N_1901,N_69);
or U8035 (N_8035,N_445,N_3151);
and U8036 (N_8036,N_2608,N_4013);
nor U8037 (N_8037,N_616,N_4081);
nand U8038 (N_8038,N_2449,N_4208);
nand U8039 (N_8039,N_3157,N_4057);
and U8040 (N_8040,N_3628,N_575);
nor U8041 (N_8041,N_2616,N_3453);
or U8042 (N_8042,N_393,N_396);
or U8043 (N_8043,N_666,N_393);
and U8044 (N_8044,N_723,N_1653);
nor U8045 (N_8045,N_1711,N_480);
nor U8046 (N_8046,N_2900,N_3743);
and U8047 (N_8047,N_1782,N_697);
nor U8048 (N_8048,N_4263,N_1600);
nor U8049 (N_8049,N_4920,N_2116);
and U8050 (N_8050,N_3475,N_1346);
or U8051 (N_8051,N_4329,N_3163);
nand U8052 (N_8052,N_3209,N_1176);
or U8053 (N_8053,N_4215,N_1627);
or U8054 (N_8054,N_3931,N_2074);
nor U8055 (N_8055,N_2083,N_182);
xor U8056 (N_8056,N_2171,N_4549);
nor U8057 (N_8057,N_2979,N_1183);
and U8058 (N_8058,N_1143,N_3473);
and U8059 (N_8059,N_2496,N_2807);
or U8060 (N_8060,N_4204,N_3539);
or U8061 (N_8061,N_4667,N_414);
nor U8062 (N_8062,N_665,N_2732);
or U8063 (N_8063,N_3523,N_1938);
or U8064 (N_8064,N_2061,N_4335);
and U8065 (N_8065,N_490,N_2744);
nand U8066 (N_8066,N_1642,N_2698);
nand U8067 (N_8067,N_1597,N_361);
and U8068 (N_8068,N_1141,N_2806);
nand U8069 (N_8069,N_2334,N_2487);
and U8070 (N_8070,N_1662,N_1328);
and U8071 (N_8071,N_1767,N_3069);
nand U8072 (N_8072,N_3570,N_3833);
and U8073 (N_8073,N_2996,N_2587);
and U8074 (N_8074,N_2171,N_2487);
or U8075 (N_8075,N_886,N_4304);
nand U8076 (N_8076,N_2444,N_1309);
and U8077 (N_8077,N_1494,N_557);
nand U8078 (N_8078,N_4971,N_3245);
nor U8079 (N_8079,N_3108,N_2588);
nand U8080 (N_8080,N_2505,N_4983);
and U8081 (N_8081,N_3763,N_1139);
nor U8082 (N_8082,N_4030,N_2694);
nand U8083 (N_8083,N_967,N_3479);
and U8084 (N_8084,N_784,N_1135);
nor U8085 (N_8085,N_844,N_2605);
or U8086 (N_8086,N_2634,N_3980);
or U8087 (N_8087,N_2109,N_3384);
or U8088 (N_8088,N_9,N_3442);
or U8089 (N_8089,N_1692,N_4817);
nor U8090 (N_8090,N_2690,N_175);
nor U8091 (N_8091,N_2712,N_300);
nand U8092 (N_8092,N_1593,N_4966);
nor U8093 (N_8093,N_4967,N_87);
xnor U8094 (N_8094,N_1272,N_1819);
nand U8095 (N_8095,N_4326,N_2955);
and U8096 (N_8096,N_1677,N_3810);
and U8097 (N_8097,N_498,N_183);
and U8098 (N_8098,N_3509,N_327);
and U8099 (N_8099,N_3784,N_882);
and U8100 (N_8100,N_3768,N_4295);
and U8101 (N_8101,N_2150,N_4679);
or U8102 (N_8102,N_4556,N_2109);
xnor U8103 (N_8103,N_3557,N_496);
xnor U8104 (N_8104,N_2152,N_3446);
nand U8105 (N_8105,N_1191,N_4603);
nor U8106 (N_8106,N_921,N_110);
or U8107 (N_8107,N_798,N_4339);
or U8108 (N_8108,N_2338,N_1493);
and U8109 (N_8109,N_1802,N_3481);
or U8110 (N_8110,N_1994,N_355);
nor U8111 (N_8111,N_3473,N_3227);
or U8112 (N_8112,N_70,N_2727);
and U8113 (N_8113,N_2129,N_3504);
nand U8114 (N_8114,N_3820,N_2575);
or U8115 (N_8115,N_3202,N_1939);
and U8116 (N_8116,N_4202,N_3409);
nor U8117 (N_8117,N_20,N_4962);
and U8118 (N_8118,N_3,N_747);
or U8119 (N_8119,N_597,N_1821);
or U8120 (N_8120,N_3243,N_3655);
and U8121 (N_8121,N_1842,N_4285);
or U8122 (N_8122,N_3450,N_485);
and U8123 (N_8123,N_4167,N_3741);
or U8124 (N_8124,N_3600,N_2143);
or U8125 (N_8125,N_4070,N_2531);
or U8126 (N_8126,N_1017,N_3310);
and U8127 (N_8127,N_1452,N_2205);
nand U8128 (N_8128,N_1844,N_905);
nand U8129 (N_8129,N_3500,N_4387);
or U8130 (N_8130,N_1876,N_4723);
nor U8131 (N_8131,N_1577,N_3638);
or U8132 (N_8132,N_1020,N_2927);
or U8133 (N_8133,N_1528,N_4540);
or U8134 (N_8134,N_3128,N_4838);
or U8135 (N_8135,N_4531,N_4047);
and U8136 (N_8136,N_1779,N_4481);
and U8137 (N_8137,N_4037,N_4905);
or U8138 (N_8138,N_3293,N_4619);
or U8139 (N_8139,N_2938,N_4010);
or U8140 (N_8140,N_2923,N_1180);
nor U8141 (N_8141,N_3449,N_1782);
or U8142 (N_8142,N_3958,N_2829);
and U8143 (N_8143,N_2691,N_76);
or U8144 (N_8144,N_3982,N_3949);
or U8145 (N_8145,N_3021,N_4768);
nor U8146 (N_8146,N_4654,N_106);
nand U8147 (N_8147,N_4149,N_55);
nor U8148 (N_8148,N_2656,N_2892);
nor U8149 (N_8149,N_1175,N_2337);
nand U8150 (N_8150,N_286,N_2431);
and U8151 (N_8151,N_4180,N_4074);
nor U8152 (N_8152,N_4354,N_2695);
nand U8153 (N_8153,N_1638,N_2894);
nand U8154 (N_8154,N_2982,N_4212);
nor U8155 (N_8155,N_1162,N_4990);
nor U8156 (N_8156,N_3416,N_4973);
and U8157 (N_8157,N_2845,N_446);
nand U8158 (N_8158,N_4387,N_4385);
and U8159 (N_8159,N_467,N_1494);
and U8160 (N_8160,N_1358,N_4772);
and U8161 (N_8161,N_1967,N_2730);
or U8162 (N_8162,N_3053,N_513);
and U8163 (N_8163,N_1193,N_173);
nor U8164 (N_8164,N_2161,N_4067);
nor U8165 (N_8165,N_2065,N_4389);
nand U8166 (N_8166,N_4102,N_1915);
nor U8167 (N_8167,N_1107,N_3626);
nand U8168 (N_8168,N_1415,N_1018);
or U8169 (N_8169,N_2625,N_1720);
nand U8170 (N_8170,N_1660,N_327);
nand U8171 (N_8171,N_974,N_1759);
and U8172 (N_8172,N_1758,N_2079);
nor U8173 (N_8173,N_4212,N_1486);
and U8174 (N_8174,N_1147,N_2394);
and U8175 (N_8175,N_2606,N_4647);
nor U8176 (N_8176,N_4215,N_3531);
and U8177 (N_8177,N_4053,N_3194);
and U8178 (N_8178,N_1569,N_2902);
nor U8179 (N_8179,N_2171,N_3487);
nor U8180 (N_8180,N_952,N_4161);
xor U8181 (N_8181,N_4161,N_4078);
nor U8182 (N_8182,N_687,N_4245);
or U8183 (N_8183,N_3792,N_1061);
nand U8184 (N_8184,N_4774,N_4294);
and U8185 (N_8185,N_2366,N_4219);
and U8186 (N_8186,N_1814,N_2711);
nor U8187 (N_8187,N_18,N_762);
nand U8188 (N_8188,N_1333,N_2530);
nor U8189 (N_8189,N_257,N_1373);
and U8190 (N_8190,N_1859,N_1356);
or U8191 (N_8191,N_3053,N_54);
or U8192 (N_8192,N_4974,N_40);
nor U8193 (N_8193,N_4069,N_1006);
nor U8194 (N_8194,N_1025,N_959);
or U8195 (N_8195,N_1946,N_3594);
or U8196 (N_8196,N_2676,N_1718);
nor U8197 (N_8197,N_2364,N_1617);
xor U8198 (N_8198,N_4792,N_3142);
nand U8199 (N_8199,N_853,N_999);
nand U8200 (N_8200,N_3713,N_2785);
or U8201 (N_8201,N_4255,N_2484);
and U8202 (N_8202,N_3109,N_4061);
and U8203 (N_8203,N_404,N_4406);
and U8204 (N_8204,N_1021,N_1153);
and U8205 (N_8205,N_4216,N_859);
or U8206 (N_8206,N_76,N_4762);
nand U8207 (N_8207,N_3503,N_3242);
or U8208 (N_8208,N_2722,N_2132);
nand U8209 (N_8209,N_559,N_4502);
or U8210 (N_8210,N_4377,N_267);
nor U8211 (N_8211,N_3227,N_1928);
nand U8212 (N_8212,N_1867,N_3363);
or U8213 (N_8213,N_1631,N_1677);
and U8214 (N_8214,N_4016,N_2304);
nand U8215 (N_8215,N_608,N_1382);
and U8216 (N_8216,N_341,N_163);
and U8217 (N_8217,N_3971,N_2001);
nand U8218 (N_8218,N_460,N_267);
or U8219 (N_8219,N_2949,N_4509);
or U8220 (N_8220,N_150,N_1058);
nand U8221 (N_8221,N_3600,N_1986);
or U8222 (N_8222,N_1709,N_4567);
and U8223 (N_8223,N_3610,N_463);
or U8224 (N_8224,N_503,N_1550);
and U8225 (N_8225,N_1853,N_3914);
nand U8226 (N_8226,N_2039,N_1277);
nor U8227 (N_8227,N_461,N_2776);
and U8228 (N_8228,N_2976,N_1817);
and U8229 (N_8229,N_2341,N_639);
and U8230 (N_8230,N_665,N_743);
or U8231 (N_8231,N_4003,N_2295);
nor U8232 (N_8232,N_3115,N_4439);
or U8233 (N_8233,N_4163,N_1841);
nor U8234 (N_8234,N_496,N_4414);
nand U8235 (N_8235,N_848,N_3313);
or U8236 (N_8236,N_2141,N_2276);
nand U8237 (N_8237,N_1097,N_3541);
xor U8238 (N_8238,N_1381,N_271);
nor U8239 (N_8239,N_2886,N_1823);
nand U8240 (N_8240,N_869,N_289);
nand U8241 (N_8241,N_2441,N_821);
nand U8242 (N_8242,N_477,N_1757);
or U8243 (N_8243,N_4241,N_686);
nor U8244 (N_8244,N_1778,N_1735);
nor U8245 (N_8245,N_3214,N_4303);
or U8246 (N_8246,N_2764,N_1009);
nor U8247 (N_8247,N_567,N_3116);
or U8248 (N_8248,N_2098,N_4163);
or U8249 (N_8249,N_2337,N_4775);
nand U8250 (N_8250,N_3407,N_964);
nand U8251 (N_8251,N_4033,N_2025);
nand U8252 (N_8252,N_1384,N_2719);
nand U8253 (N_8253,N_2135,N_2882);
nand U8254 (N_8254,N_2331,N_166);
nor U8255 (N_8255,N_1113,N_774);
nand U8256 (N_8256,N_508,N_3044);
nand U8257 (N_8257,N_1044,N_2399);
nand U8258 (N_8258,N_2121,N_179);
nor U8259 (N_8259,N_3201,N_3661);
and U8260 (N_8260,N_4923,N_3276);
nand U8261 (N_8261,N_3304,N_2621);
nand U8262 (N_8262,N_458,N_605);
or U8263 (N_8263,N_2549,N_3475);
nand U8264 (N_8264,N_1718,N_4966);
nor U8265 (N_8265,N_3436,N_4143);
nand U8266 (N_8266,N_164,N_2205);
or U8267 (N_8267,N_552,N_2031);
or U8268 (N_8268,N_1257,N_4613);
or U8269 (N_8269,N_279,N_4031);
nand U8270 (N_8270,N_3411,N_2683);
and U8271 (N_8271,N_3124,N_1949);
nand U8272 (N_8272,N_1773,N_4612);
nor U8273 (N_8273,N_4661,N_3889);
nor U8274 (N_8274,N_3385,N_1107);
and U8275 (N_8275,N_77,N_1548);
nor U8276 (N_8276,N_2760,N_2284);
nand U8277 (N_8277,N_4090,N_4969);
and U8278 (N_8278,N_233,N_3663);
nor U8279 (N_8279,N_3253,N_1822);
nor U8280 (N_8280,N_2897,N_3352);
nor U8281 (N_8281,N_4828,N_1367);
or U8282 (N_8282,N_3255,N_3368);
nor U8283 (N_8283,N_1838,N_2218);
and U8284 (N_8284,N_2889,N_883);
xnor U8285 (N_8285,N_1628,N_3507);
and U8286 (N_8286,N_1365,N_3764);
and U8287 (N_8287,N_1319,N_4055);
and U8288 (N_8288,N_3507,N_1605);
or U8289 (N_8289,N_1578,N_2112);
or U8290 (N_8290,N_2835,N_3719);
and U8291 (N_8291,N_2860,N_3646);
and U8292 (N_8292,N_1830,N_1958);
nand U8293 (N_8293,N_956,N_2021);
or U8294 (N_8294,N_2687,N_2234);
nor U8295 (N_8295,N_601,N_964);
nand U8296 (N_8296,N_865,N_3476);
nor U8297 (N_8297,N_3929,N_2984);
and U8298 (N_8298,N_717,N_2405);
or U8299 (N_8299,N_726,N_1204);
or U8300 (N_8300,N_2930,N_3762);
nor U8301 (N_8301,N_2008,N_1281);
or U8302 (N_8302,N_4760,N_1739);
or U8303 (N_8303,N_3432,N_1562);
and U8304 (N_8304,N_3004,N_427);
nand U8305 (N_8305,N_4018,N_1872);
nand U8306 (N_8306,N_3111,N_3112);
and U8307 (N_8307,N_597,N_4410);
nand U8308 (N_8308,N_3812,N_4542);
nor U8309 (N_8309,N_3226,N_778);
nand U8310 (N_8310,N_1620,N_4263);
nand U8311 (N_8311,N_4864,N_3001);
nand U8312 (N_8312,N_2139,N_4130);
nor U8313 (N_8313,N_1648,N_2254);
and U8314 (N_8314,N_3475,N_1309);
nand U8315 (N_8315,N_1833,N_2280);
nor U8316 (N_8316,N_734,N_2737);
and U8317 (N_8317,N_3482,N_250);
or U8318 (N_8318,N_608,N_1738);
and U8319 (N_8319,N_1564,N_4710);
nand U8320 (N_8320,N_3299,N_2213);
or U8321 (N_8321,N_1533,N_4027);
nor U8322 (N_8322,N_2750,N_4281);
nor U8323 (N_8323,N_228,N_174);
nand U8324 (N_8324,N_2448,N_333);
xnor U8325 (N_8325,N_1893,N_1722);
or U8326 (N_8326,N_3408,N_801);
nor U8327 (N_8327,N_1860,N_4044);
or U8328 (N_8328,N_4050,N_709);
or U8329 (N_8329,N_1986,N_399);
or U8330 (N_8330,N_4546,N_2781);
or U8331 (N_8331,N_4356,N_1163);
nor U8332 (N_8332,N_4112,N_3474);
nor U8333 (N_8333,N_270,N_1220);
or U8334 (N_8334,N_420,N_1124);
xnor U8335 (N_8335,N_3733,N_978);
nor U8336 (N_8336,N_433,N_3772);
nor U8337 (N_8337,N_2560,N_1828);
or U8338 (N_8338,N_1018,N_356);
nor U8339 (N_8339,N_1375,N_3880);
nor U8340 (N_8340,N_3347,N_4007);
and U8341 (N_8341,N_2321,N_4891);
and U8342 (N_8342,N_451,N_2307);
xor U8343 (N_8343,N_515,N_1570);
or U8344 (N_8344,N_592,N_3048);
nand U8345 (N_8345,N_82,N_3810);
nor U8346 (N_8346,N_4591,N_3145);
or U8347 (N_8347,N_3351,N_163);
and U8348 (N_8348,N_1542,N_2795);
nor U8349 (N_8349,N_1797,N_1539);
nor U8350 (N_8350,N_2252,N_436);
nor U8351 (N_8351,N_4794,N_3144);
nor U8352 (N_8352,N_2863,N_1582);
and U8353 (N_8353,N_998,N_4481);
nor U8354 (N_8354,N_3036,N_4578);
nand U8355 (N_8355,N_325,N_399);
nand U8356 (N_8356,N_4845,N_91);
nor U8357 (N_8357,N_4662,N_541);
or U8358 (N_8358,N_1088,N_3631);
and U8359 (N_8359,N_2407,N_1402);
nor U8360 (N_8360,N_1067,N_1808);
and U8361 (N_8361,N_3624,N_2956);
or U8362 (N_8362,N_3050,N_4798);
nor U8363 (N_8363,N_4464,N_455);
and U8364 (N_8364,N_3105,N_4829);
or U8365 (N_8365,N_1497,N_1640);
nor U8366 (N_8366,N_3111,N_466);
and U8367 (N_8367,N_2981,N_1816);
nor U8368 (N_8368,N_1001,N_1813);
and U8369 (N_8369,N_4297,N_2625);
and U8370 (N_8370,N_2705,N_454);
and U8371 (N_8371,N_2029,N_3712);
or U8372 (N_8372,N_1573,N_1188);
or U8373 (N_8373,N_482,N_2822);
or U8374 (N_8374,N_3259,N_2959);
and U8375 (N_8375,N_4449,N_2367);
and U8376 (N_8376,N_1589,N_989);
or U8377 (N_8377,N_3212,N_4573);
nor U8378 (N_8378,N_3258,N_3833);
or U8379 (N_8379,N_4933,N_398);
xnor U8380 (N_8380,N_2431,N_4654);
nand U8381 (N_8381,N_4527,N_1151);
nor U8382 (N_8382,N_2832,N_4258);
nor U8383 (N_8383,N_2220,N_4205);
nand U8384 (N_8384,N_4466,N_3769);
and U8385 (N_8385,N_3395,N_1208);
nand U8386 (N_8386,N_3600,N_1980);
and U8387 (N_8387,N_3002,N_1620);
nor U8388 (N_8388,N_59,N_4372);
or U8389 (N_8389,N_544,N_2597);
or U8390 (N_8390,N_4260,N_2795);
and U8391 (N_8391,N_1410,N_1288);
nand U8392 (N_8392,N_1915,N_4691);
or U8393 (N_8393,N_109,N_4969);
and U8394 (N_8394,N_520,N_1680);
nor U8395 (N_8395,N_1602,N_3866);
and U8396 (N_8396,N_1795,N_3017);
or U8397 (N_8397,N_3583,N_3652);
and U8398 (N_8398,N_1963,N_2472);
nand U8399 (N_8399,N_3498,N_3419);
or U8400 (N_8400,N_1914,N_370);
nand U8401 (N_8401,N_4697,N_971);
nor U8402 (N_8402,N_3187,N_2401);
nor U8403 (N_8403,N_4443,N_74);
or U8404 (N_8404,N_4816,N_3691);
nand U8405 (N_8405,N_2990,N_3176);
nand U8406 (N_8406,N_1833,N_436);
and U8407 (N_8407,N_937,N_727);
nand U8408 (N_8408,N_524,N_1804);
or U8409 (N_8409,N_1527,N_1393);
and U8410 (N_8410,N_744,N_1884);
and U8411 (N_8411,N_4653,N_3178);
and U8412 (N_8412,N_3466,N_1065);
nor U8413 (N_8413,N_3317,N_3862);
nand U8414 (N_8414,N_2718,N_582);
nand U8415 (N_8415,N_1062,N_2880);
and U8416 (N_8416,N_3390,N_2205);
and U8417 (N_8417,N_1529,N_932);
nand U8418 (N_8418,N_4216,N_1115);
nand U8419 (N_8419,N_3664,N_4702);
nand U8420 (N_8420,N_1573,N_3619);
nor U8421 (N_8421,N_63,N_152);
and U8422 (N_8422,N_320,N_311);
nor U8423 (N_8423,N_4738,N_3957);
nand U8424 (N_8424,N_4289,N_2187);
nor U8425 (N_8425,N_2642,N_3057);
or U8426 (N_8426,N_3460,N_1191);
nor U8427 (N_8427,N_3054,N_3294);
and U8428 (N_8428,N_4846,N_4558);
or U8429 (N_8429,N_3782,N_2822);
nand U8430 (N_8430,N_2581,N_1322);
or U8431 (N_8431,N_1697,N_2941);
and U8432 (N_8432,N_1274,N_1561);
and U8433 (N_8433,N_3302,N_3939);
nand U8434 (N_8434,N_739,N_190);
nor U8435 (N_8435,N_1647,N_4147);
and U8436 (N_8436,N_2198,N_4718);
nand U8437 (N_8437,N_3115,N_1176);
and U8438 (N_8438,N_2837,N_4806);
and U8439 (N_8439,N_1683,N_4650);
or U8440 (N_8440,N_4601,N_331);
nand U8441 (N_8441,N_2594,N_69);
or U8442 (N_8442,N_3582,N_4629);
or U8443 (N_8443,N_1107,N_4247);
nor U8444 (N_8444,N_3430,N_2783);
and U8445 (N_8445,N_4218,N_4899);
and U8446 (N_8446,N_709,N_3607);
and U8447 (N_8447,N_4296,N_1171);
nand U8448 (N_8448,N_4275,N_295);
nand U8449 (N_8449,N_1070,N_3881);
or U8450 (N_8450,N_1910,N_3655);
nor U8451 (N_8451,N_1915,N_4601);
nand U8452 (N_8452,N_2277,N_845);
or U8453 (N_8453,N_1444,N_4051);
nand U8454 (N_8454,N_3879,N_1795);
nor U8455 (N_8455,N_1951,N_4622);
or U8456 (N_8456,N_634,N_1740);
or U8457 (N_8457,N_748,N_3475);
and U8458 (N_8458,N_3099,N_1261);
nor U8459 (N_8459,N_128,N_4244);
nand U8460 (N_8460,N_3666,N_3590);
and U8461 (N_8461,N_1230,N_3121);
nor U8462 (N_8462,N_3443,N_2759);
nor U8463 (N_8463,N_870,N_3171);
or U8464 (N_8464,N_2953,N_4706);
or U8465 (N_8465,N_2502,N_714);
or U8466 (N_8466,N_1451,N_3858);
or U8467 (N_8467,N_4737,N_2732);
and U8468 (N_8468,N_3799,N_519);
nand U8469 (N_8469,N_1150,N_4782);
or U8470 (N_8470,N_4021,N_2288);
and U8471 (N_8471,N_1084,N_2397);
nand U8472 (N_8472,N_4286,N_3089);
nor U8473 (N_8473,N_2146,N_1867);
and U8474 (N_8474,N_3848,N_2960);
and U8475 (N_8475,N_257,N_2557);
or U8476 (N_8476,N_0,N_1759);
and U8477 (N_8477,N_788,N_2314);
or U8478 (N_8478,N_1653,N_683);
nand U8479 (N_8479,N_1381,N_1555);
nor U8480 (N_8480,N_519,N_3930);
nand U8481 (N_8481,N_2012,N_3830);
and U8482 (N_8482,N_1580,N_1803);
or U8483 (N_8483,N_3891,N_768);
or U8484 (N_8484,N_50,N_4323);
or U8485 (N_8485,N_504,N_3083);
or U8486 (N_8486,N_2319,N_1502);
nand U8487 (N_8487,N_2007,N_4680);
or U8488 (N_8488,N_1529,N_44);
nor U8489 (N_8489,N_3953,N_4447);
and U8490 (N_8490,N_478,N_4221);
nor U8491 (N_8491,N_642,N_3240);
nor U8492 (N_8492,N_4373,N_3550);
and U8493 (N_8493,N_12,N_520);
nor U8494 (N_8494,N_2470,N_4453);
xor U8495 (N_8495,N_1956,N_3628);
or U8496 (N_8496,N_749,N_4715);
and U8497 (N_8497,N_726,N_2073);
nor U8498 (N_8498,N_4128,N_2562);
nand U8499 (N_8499,N_4127,N_522);
or U8500 (N_8500,N_3902,N_4877);
and U8501 (N_8501,N_4229,N_1176);
nand U8502 (N_8502,N_726,N_2938);
or U8503 (N_8503,N_2143,N_4883);
nand U8504 (N_8504,N_503,N_533);
or U8505 (N_8505,N_251,N_2437);
nor U8506 (N_8506,N_2973,N_2723);
or U8507 (N_8507,N_982,N_67);
nand U8508 (N_8508,N_1550,N_3345);
or U8509 (N_8509,N_3929,N_2381);
and U8510 (N_8510,N_2179,N_57);
nor U8511 (N_8511,N_2212,N_3919);
nor U8512 (N_8512,N_512,N_1691);
nand U8513 (N_8513,N_977,N_2954);
and U8514 (N_8514,N_806,N_3359);
nor U8515 (N_8515,N_642,N_2541);
nor U8516 (N_8516,N_3207,N_3508);
nand U8517 (N_8517,N_1076,N_3107);
or U8518 (N_8518,N_114,N_545);
or U8519 (N_8519,N_3098,N_4645);
nor U8520 (N_8520,N_764,N_3770);
nand U8521 (N_8521,N_1566,N_1405);
nand U8522 (N_8522,N_2296,N_4720);
nand U8523 (N_8523,N_747,N_4978);
or U8524 (N_8524,N_4804,N_1419);
and U8525 (N_8525,N_1073,N_1381);
nor U8526 (N_8526,N_1648,N_236);
nor U8527 (N_8527,N_1659,N_4714);
nand U8528 (N_8528,N_868,N_3061);
and U8529 (N_8529,N_4913,N_3786);
and U8530 (N_8530,N_4444,N_99);
or U8531 (N_8531,N_2428,N_1079);
or U8532 (N_8532,N_386,N_365);
nand U8533 (N_8533,N_2840,N_2241);
or U8534 (N_8534,N_4780,N_847);
nand U8535 (N_8535,N_2686,N_624);
and U8536 (N_8536,N_2520,N_4539);
and U8537 (N_8537,N_3603,N_3942);
and U8538 (N_8538,N_2135,N_2456);
nand U8539 (N_8539,N_1162,N_2845);
and U8540 (N_8540,N_1356,N_4497);
nor U8541 (N_8541,N_3270,N_2977);
nor U8542 (N_8542,N_1304,N_260);
and U8543 (N_8543,N_2853,N_1936);
or U8544 (N_8544,N_899,N_342);
nor U8545 (N_8545,N_4288,N_222);
nor U8546 (N_8546,N_519,N_843);
nor U8547 (N_8547,N_2076,N_258);
nand U8548 (N_8548,N_3833,N_299);
and U8549 (N_8549,N_1357,N_1583);
nand U8550 (N_8550,N_1831,N_2798);
and U8551 (N_8551,N_2258,N_4193);
nand U8552 (N_8552,N_2577,N_514);
and U8553 (N_8553,N_4584,N_4950);
and U8554 (N_8554,N_2681,N_3238);
or U8555 (N_8555,N_436,N_4083);
nand U8556 (N_8556,N_2545,N_4472);
or U8557 (N_8557,N_2236,N_1841);
nor U8558 (N_8558,N_570,N_1224);
or U8559 (N_8559,N_990,N_1634);
nand U8560 (N_8560,N_791,N_4382);
and U8561 (N_8561,N_2768,N_1021);
and U8562 (N_8562,N_527,N_953);
nand U8563 (N_8563,N_2345,N_3146);
nand U8564 (N_8564,N_1770,N_3460);
and U8565 (N_8565,N_4034,N_1068);
and U8566 (N_8566,N_2513,N_827);
or U8567 (N_8567,N_1389,N_3102);
nor U8568 (N_8568,N_2016,N_414);
nor U8569 (N_8569,N_309,N_3710);
or U8570 (N_8570,N_1391,N_3612);
and U8571 (N_8571,N_3566,N_2165);
or U8572 (N_8572,N_1977,N_1877);
and U8573 (N_8573,N_1280,N_3853);
nor U8574 (N_8574,N_554,N_4791);
and U8575 (N_8575,N_717,N_2513);
and U8576 (N_8576,N_4242,N_2628);
nor U8577 (N_8577,N_821,N_3391);
nor U8578 (N_8578,N_4267,N_2297);
nand U8579 (N_8579,N_817,N_1130);
and U8580 (N_8580,N_3039,N_3465);
or U8581 (N_8581,N_4457,N_1369);
and U8582 (N_8582,N_4104,N_1664);
or U8583 (N_8583,N_3908,N_1558);
and U8584 (N_8584,N_3652,N_4806);
or U8585 (N_8585,N_1711,N_4551);
nand U8586 (N_8586,N_4692,N_881);
or U8587 (N_8587,N_3894,N_3770);
nand U8588 (N_8588,N_3849,N_3062);
nor U8589 (N_8589,N_843,N_306);
nor U8590 (N_8590,N_1138,N_3594);
nand U8591 (N_8591,N_466,N_4097);
nor U8592 (N_8592,N_3519,N_1410);
nor U8593 (N_8593,N_626,N_2151);
and U8594 (N_8594,N_4985,N_868);
nand U8595 (N_8595,N_4971,N_263);
nor U8596 (N_8596,N_3818,N_242);
nand U8597 (N_8597,N_1124,N_465);
or U8598 (N_8598,N_325,N_3727);
or U8599 (N_8599,N_1491,N_3148);
or U8600 (N_8600,N_1862,N_135);
and U8601 (N_8601,N_2075,N_4648);
or U8602 (N_8602,N_205,N_4844);
nand U8603 (N_8603,N_4200,N_3757);
nand U8604 (N_8604,N_4936,N_4384);
nand U8605 (N_8605,N_4784,N_3269);
or U8606 (N_8606,N_1703,N_3036);
nor U8607 (N_8607,N_4714,N_3466);
and U8608 (N_8608,N_1718,N_833);
nand U8609 (N_8609,N_4142,N_4148);
and U8610 (N_8610,N_1824,N_3127);
or U8611 (N_8611,N_4114,N_4051);
nor U8612 (N_8612,N_885,N_614);
and U8613 (N_8613,N_2099,N_69);
and U8614 (N_8614,N_1425,N_308);
and U8615 (N_8615,N_477,N_4462);
and U8616 (N_8616,N_2209,N_3141);
or U8617 (N_8617,N_1421,N_3369);
and U8618 (N_8618,N_442,N_4267);
nand U8619 (N_8619,N_781,N_4087);
and U8620 (N_8620,N_1025,N_436);
and U8621 (N_8621,N_24,N_2797);
or U8622 (N_8622,N_2468,N_4921);
nand U8623 (N_8623,N_4402,N_2953);
nand U8624 (N_8624,N_3085,N_4982);
or U8625 (N_8625,N_3469,N_566);
or U8626 (N_8626,N_1214,N_3593);
or U8627 (N_8627,N_3914,N_3445);
and U8628 (N_8628,N_2174,N_124);
nor U8629 (N_8629,N_4371,N_2643);
nor U8630 (N_8630,N_3903,N_2669);
or U8631 (N_8631,N_4717,N_2642);
xor U8632 (N_8632,N_1875,N_3448);
or U8633 (N_8633,N_333,N_3912);
nand U8634 (N_8634,N_2859,N_3725);
or U8635 (N_8635,N_1787,N_4672);
and U8636 (N_8636,N_414,N_1059);
nand U8637 (N_8637,N_1423,N_3908);
nor U8638 (N_8638,N_1611,N_521);
nor U8639 (N_8639,N_1080,N_4875);
and U8640 (N_8640,N_2104,N_30);
and U8641 (N_8641,N_4611,N_1258);
nor U8642 (N_8642,N_4230,N_4565);
and U8643 (N_8643,N_4571,N_1439);
nor U8644 (N_8644,N_4241,N_4402);
and U8645 (N_8645,N_4836,N_522);
nor U8646 (N_8646,N_4074,N_2062);
nor U8647 (N_8647,N_3113,N_4663);
nand U8648 (N_8648,N_2955,N_3034);
and U8649 (N_8649,N_3829,N_2378);
nor U8650 (N_8650,N_163,N_1522);
nor U8651 (N_8651,N_3434,N_3950);
or U8652 (N_8652,N_1149,N_3164);
and U8653 (N_8653,N_1127,N_3582);
or U8654 (N_8654,N_2383,N_1251);
and U8655 (N_8655,N_4855,N_3928);
xnor U8656 (N_8656,N_1122,N_4206);
nor U8657 (N_8657,N_3760,N_2910);
nand U8658 (N_8658,N_3929,N_3453);
and U8659 (N_8659,N_3644,N_1628);
nor U8660 (N_8660,N_4256,N_4630);
and U8661 (N_8661,N_445,N_3514);
and U8662 (N_8662,N_3036,N_205);
or U8663 (N_8663,N_3705,N_1414);
nand U8664 (N_8664,N_3146,N_1076);
nor U8665 (N_8665,N_1544,N_4503);
and U8666 (N_8666,N_1245,N_1739);
and U8667 (N_8667,N_2024,N_1932);
nor U8668 (N_8668,N_3536,N_36);
and U8669 (N_8669,N_3255,N_2164);
and U8670 (N_8670,N_993,N_956);
nor U8671 (N_8671,N_830,N_2220);
nand U8672 (N_8672,N_4381,N_3725);
and U8673 (N_8673,N_1382,N_33);
nand U8674 (N_8674,N_1690,N_1464);
and U8675 (N_8675,N_737,N_1943);
nand U8676 (N_8676,N_1918,N_4451);
and U8677 (N_8677,N_1928,N_2141);
or U8678 (N_8678,N_2102,N_1072);
nand U8679 (N_8679,N_1088,N_1785);
nand U8680 (N_8680,N_688,N_3331);
or U8681 (N_8681,N_2101,N_1264);
and U8682 (N_8682,N_3645,N_4741);
nand U8683 (N_8683,N_3876,N_1518);
and U8684 (N_8684,N_1954,N_2850);
and U8685 (N_8685,N_3795,N_4527);
nand U8686 (N_8686,N_273,N_137);
and U8687 (N_8687,N_3221,N_1799);
nand U8688 (N_8688,N_3830,N_4155);
nand U8689 (N_8689,N_396,N_608);
or U8690 (N_8690,N_3454,N_3927);
nand U8691 (N_8691,N_4086,N_898);
and U8692 (N_8692,N_4262,N_1930);
nor U8693 (N_8693,N_4854,N_2650);
or U8694 (N_8694,N_4775,N_2482);
or U8695 (N_8695,N_2068,N_1999);
and U8696 (N_8696,N_4551,N_1824);
or U8697 (N_8697,N_3061,N_413);
nand U8698 (N_8698,N_2418,N_3027);
and U8699 (N_8699,N_3701,N_1886);
nand U8700 (N_8700,N_4607,N_1488);
nand U8701 (N_8701,N_1993,N_3096);
or U8702 (N_8702,N_1737,N_4358);
or U8703 (N_8703,N_1951,N_696);
nor U8704 (N_8704,N_795,N_1948);
or U8705 (N_8705,N_4401,N_1618);
nor U8706 (N_8706,N_4063,N_4556);
nor U8707 (N_8707,N_3832,N_476);
nand U8708 (N_8708,N_2956,N_385);
nor U8709 (N_8709,N_3254,N_776);
or U8710 (N_8710,N_1870,N_1359);
nor U8711 (N_8711,N_1025,N_2025);
and U8712 (N_8712,N_4436,N_1031);
and U8713 (N_8713,N_3454,N_3173);
or U8714 (N_8714,N_409,N_1271);
nor U8715 (N_8715,N_3197,N_1822);
nor U8716 (N_8716,N_2605,N_4022);
and U8717 (N_8717,N_28,N_3398);
or U8718 (N_8718,N_1640,N_1001);
nor U8719 (N_8719,N_4012,N_1129);
and U8720 (N_8720,N_3504,N_2310);
and U8721 (N_8721,N_746,N_4136);
or U8722 (N_8722,N_4836,N_1727);
nand U8723 (N_8723,N_4539,N_2990);
and U8724 (N_8724,N_3105,N_944);
nor U8725 (N_8725,N_3964,N_677);
nand U8726 (N_8726,N_2055,N_4993);
nor U8727 (N_8727,N_3405,N_1022);
nor U8728 (N_8728,N_3076,N_255);
and U8729 (N_8729,N_1921,N_716);
nand U8730 (N_8730,N_4860,N_354);
nor U8731 (N_8731,N_4067,N_296);
and U8732 (N_8732,N_1761,N_3505);
or U8733 (N_8733,N_908,N_2063);
nor U8734 (N_8734,N_2333,N_4608);
nor U8735 (N_8735,N_3276,N_626);
nand U8736 (N_8736,N_111,N_4705);
and U8737 (N_8737,N_2607,N_4477);
and U8738 (N_8738,N_4865,N_2580);
nand U8739 (N_8739,N_3964,N_562);
or U8740 (N_8740,N_2057,N_4340);
xor U8741 (N_8741,N_4284,N_1071);
or U8742 (N_8742,N_1691,N_1462);
nand U8743 (N_8743,N_3098,N_1824);
nor U8744 (N_8744,N_376,N_2965);
and U8745 (N_8745,N_1921,N_4537);
and U8746 (N_8746,N_228,N_4523);
and U8747 (N_8747,N_678,N_4782);
and U8748 (N_8748,N_4117,N_2427);
or U8749 (N_8749,N_4864,N_1819);
or U8750 (N_8750,N_1495,N_1487);
nor U8751 (N_8751,N_2259,N_4386);
and U8752 (N_8752,N_2548,N_4343);
and U8753 (N_8753,N_1759,N_4507);
and U8754 (N_8754,N_205,N_1233);
or U8755 (N_8755,N_1394,N_3323);
nand U8756 (N_8756,N_961,N_4592);
or U8757 (N_8757,N_3989,N_2323);
or U8758 (N_8758,N_2289,N_165);
and U8759 (N_8759,N_3368,N_3872);
and U8760 (N_8760,N_904,N_3617);
and U8761 (N_8761,N_4256,N_1700);
nand U8762 (N_8762,N_4200,N_305);
and U8763 (N_8763,N_2578,N_5);
or U8764 (N_8764,N_3492,N_4171);
or U8765 (N_8765,N_297,N_3551);
or U8766 (N_8766,N_3484,N_4471);
nor U8767 (N_8767,N_3873,N_1288);
nor U8768 (N_8768,N_1056,N_691);
and U8769 (N_8769,N_673,N_882);
or U8770 (N_8770,N_3462,N_2384);
nor U8771 (N_8771,N_1687,N_3764);
nand U8772 (N_8772,N_3763,N_1079);
or U8773 (N_8773,N_2874,N_4644);
nor U8774 (N_8774,N_4557,N_452);
nand U8775 (N_8775,N_2276,N_4160);
and U8776 (N_8776,N_4527,N_3825);
nand U8777 (N_8777,N_4226,N_3109);
and U8778 (N_8778,N_4203,N_1763);
nor U8779 (N_8779,N_1392,N_141);
or U8780 (N_8780,N_4991,N_448);
and U8781 (N_8781,N_72,N_2256);
or U8782 (N_8782,N_367,N_3763);
and U8783 (N_8783,N_4012,N_3154);
and U8784 (N_8784,N_3415,N_2599);
nand U8785 (N_8785,N_4653,N_4645);
nor U8786 (N_8786,N_1836,N_214);
or U8787 (N_8787,N_1107,N_4409);
and U8788 (N_8788,N_2156,N_3788);
nand U8789 (N_8789,N_2073,N_3778);
nand U8790 (N_8790,N_3333,N_1991);
nand U8791 (N_8791,N_2637,N_853);
or U8792 (N_8792,N_3247,N_2713);
nand U8793 (N_8793,N_2441,N_4616);
and U8794 (N_8794,N_4779,N_4243);
nand U8795 (N_8795,N_556,N_870);
or U8796 (N_8796,N_2397,N_4225);
nor U8797 (N_8797,N_138,N_2935);
nand U8798 (N_8798,N_2121,N_2784);
and U8799 (N_8799,N_2899,N_440);
and U8800 (N_8800,N_3651,N_2939);
or U8801 (N_8801,N_2610,N_2304);
nand U8802 (N_8802,N_1086,N_1514);
nand U8803 (N_8803,N_1453,N_1376);
and U8804 (N_8804,N_3566,N_3637);
nor U8805 (N_8805,N_3184,N_2297);
nor U8806 (N_8806,N_4647,N_4951);
and U8807 (N_8807,N_4009,N_4661);
nand U8808 (N_8808,N_3664,N_1795);
nor U8809 (N_8809,N_557,N_4870);
and U8810 (N_8810,N_3363,N_1742);
nand U8811 (N_8811,N_1971,N_1629);
or U8812 (N_8812,N_1641,N_3373);
nand U8813 (N_8813,N_1621,N_1075);
and U8814 (N_8814,N_3894,N_4641);
nand U8815 (N_8815,N_3170,N_3852);
nand U8816 (N_8816,N_3222,N_705);
nor U8817 (N_8817,N_519,N_4259);
nor U8818 (N_8818,N_1731,N_2176);
nand U8819 (N_8819,N_3075,N_3463);
nand U8820 (N_8820,N_4071,N_2309);
nand U8821 (N_8821,N_4228,N_2184);
and U8822 (N_8822,N_335,N_3076);
nand U8823 (N_8823,N_275,N_59);
and U8824 (N_8824,N_3178,N_1458);
nor U8825 (N_8825,N_3128,N_2199);
or U8826 (N_8826,N_1305,N_2741);
nand U8827 (N_8827,N_267,N_4424);
nor U8828 (N_8828,N_4781,N_3829);
nor U8829 (N_8829,N_1587,N_195);
or U8830 (N_8830,N_396,N_2269);
and U8831 (N_8831,N_3700,N_2914);
nor U8832 (N_8832,N_1361,N_303);
and U8833 (N_8833,N_1453,N_466);
nand U8834 (N_8834,N_1066,N_2806);
nor U8835 (N_8835,N_1621,N_3227);
nand U8836 (N_8836,N_1993,N_2230);
nor U8837 (N_8837,N_3767,N_4641);
nor U8838 (N_8838,N_6,N_2998);
nor U8839 (N_8839,N_537,N_125);
and U8840 (N_8840,N_2662,N_4092);
nand U8841 (N_8841,N_1145,N_842);
and U8842 (N_8842,N_2716,N_3664);
and U8843 (N_8843,N_4716,N_544);
and U8844 (N_8844,N_404,N_3586);
and U8845 (N_8845,N_2765,N_1818);
nor U8846 (N_8846,N_3753,N_1012);
or U8847 (N_8847,N_270,N_2843);
or U8848 (N_8848,N_3975,N_91);
nor U8849 (N_8849,N_791,N_3044);
and U8850 (N_8850,N_827,N_3133);
or U8851 (N_8851,N_1477,N_1371);
and U8852 (N_8852,N_1440,N_4112);
or U8853 (N_8853,N_1519,N_4250);
or U8854 (N_8854,N_3987,N_3637);
nor U8855 (N_8855,N_2416,N_179);
or U8856 (N_8856,N_925,N_2887);
nor U8857 (N_8857,N_4610,N_43);
or U8858 (N_8858,N_443,N_1505);
nor U8859 (N_8859,N_4239,N_3575);
nand U8860 (N_8860,N_3618,N_3841);
and U8861 (N_8861,N_2356,N_15);
nor U8862 (N_8862,N_1312,N_4277);
or U8863 (N_8863,N_4440,N_4632);
nand U8864 (N_8864,N_2205,N_383);
or U8865 (N_8865,N_1810,N_2644);
nand U8866 (N_8866,N_3553,N_40);
nor U8867 (N_8867,N_4885,N_1633);
nor U8868 (N_8868,N_2181,N_3305);
and U8869 (N_8869,N_4915,N_4795);
and U8870 (N_8870,N_18,N_1612);
nand U8871 (N_8871,N_3412,N_576);
nor U8872 (N_8872,N_2833,N_3043);
nor U8873 (N_8873,N_4893,N_4242);
and U8874 (N_8874,N_3248,N_3121);
or U8875 (N_8875,N_3986,N_1971);
and U8876 (N_8876,N_3280,N_642);
and U8877 (N_8877,N_4578,N_2717);
nand U8878 (N_8878,N_3108,N_1463);
or U8879 (N_8879,N_4835,N_2215);
or U8880 (N_8880,N_37,N_3161);
nor U8881 (N_8881,N_4635,N_4715);
xor U8882 (N_8882,N_4478,N_2542);
and U8883 (N_8883,N_3921,N_964);
and U8884 (N_8884,N_1928,N_859);
or U8885 (N_8885,N_2249,N_3389);
nor U8886 (N_8886,N_2367,N_3940);
nor U8887 (N_8887,N_1268,N_2001);
or U8888 (N_8888,N_4343,N_1275);
or U8889 (N_8889,N_3149,N_3713);
nand U8890 (N_8890,N_4596,N_1637);
or U8891 (N_8891,N_4999,N_4315);
or U8892 (N_8892,N_2250,N_2339);
nand U8893 (N_8893,N_2683,N_1223);
nand U8894 (N_8894,N_3249,N_1312);
nand U8895 (N_8895,N_4851,N_714);
nand U8896 (N_8896,N_1396,N_253);
nor U8897 (N_8897,N_456,N_1731);
or U8898 (N_8898,N_1396,N_1156);
xor U8899 (N_8899,N_3128,N_4133);
and U8900 (N_8900,N_4330,N_4086);
or U8901 (N_8901,N_4114,N_2294);
and U8902 (N_8902,N_2286,N_1570);
and U8903 (N_8903,N_2921,N_1968);
nor U8904 (N_8904,N_2730,N_632);
and U8905 (N_8905,N_4283,N_4435);
nand U8906 (N_8906,N_953,N_2731);
nor U8907 (N_8907,N_1025,N_2109);
and U8908 (N_8908,N_651,N_1756);
nand U8909 (N_8909,N_3913,N_2286);
xor U8910 (N_8910,N_4113,N_3314);
or U8911 (N_8911,N_592,N_2584);
nor U8912 (N_8912,N_3868,N_4586);
nor U8913 (N_8913,N_3245,N_4715);
nand U8914 (N_8914,N_4888,N_1967);
nor U8915 (N_8915,N_928,N_92);
or U8916 (N_8916,N_2573,N_1274);
nor U8917 (N_8917,N_2869,N_3913);
xor U8918 (N_8918,N_3593,N_4611);
or U8919 (N_8919,N_2299,N_815);
nor U8920 (N_8920,N_3935,N_1506);
nor U8921 (N_8921,N_4627,N_4882);
and U8922 (N_8922,N_3012,N_1542);
and U8923 (N_8923,N_1867,N_2703);
nor U8924 (N_8924,N_3449,N_4288);
nand U8925 (N_8925,N_569,N_1495);
or U8926 (N_8926,N_4755,N_2072);
nand U8927 (N_8927,N_3826,N_3841);
and U8928 (N_8928,N_4305,N_2279);
and U8929 (N_8929,N_4625,N_3218);
nor U8930 (N_8930,N_812,N_1160);
or U8931 (N_8931,N_2792,N_1988);
or U8932 (N_8932,N_4320,N_601);
or U8933 (N_8933,N_3457,N_4539);
and U8934 (N_8934,N_2938,N_27);
nand U8935 (N_8935,N_4925,N_606);
nand U8936 (N_8936,N_673,N_3092);
nor U8937 (N_8937,N_977,N_2120);
nand U8938 (N_8938,N_2292,N_3542);
nand U8939 (N_8939,N_3203,N_2973);
nand U8940 (N_8940,N_848,N_1852);
nand U8941 (N_8941,N_3027,N_2860);
or U8942 (N_8942,N_1773,N_2342);
and U8943 (N_8943,N_4802,N_2193);
nor U8944 (N_8944,N_1899,N_725);
and U8945 (N_8945,N_3786,N_4273);
and U8946 (N_8946,N_361,N_3539);
nor U8947 (N_8947,N_467,N_3000);
nor U8948 (N_8948,N_3070,N_2799);
and U8949 (N_8949,N_3910,N_1913);
nand U8950 (N_8950,N_1055,N_1281);
or U8951 (N_8951,N_3969,N_647);
nor U8952 (N_8952,N_1390,N_2945);
nand U8953 (N_8953,N_4378,N_4707);
nor U8954 (N_8954,N_2634,N_2764);
or U8955 (N_8955,N_1857,N_1313);
or U8956 (N_8956,N_1407,N_4679);
or U8957 (N_8957,N_1883,N_1201);
or U8958 (N_8958,N_2114,N_912);
nand U8959 (N_8959,N_1336,N_4195);
or U8960 (N_8960,N_4797,N_2743);
nor U8961 (N_8961,N_4634,N_160);
or U8962 (N_8962,N_3114,N_63);
nor U8963 (N_8963,N_2887,N_788);
or U8964 (N_8964,N_2348,N_4771);
nor U8965 (N_8965,N_1979,N_4104);
nand U8966 (N_8966,N_4643,N_172);
or U8967 (N_8967,N_743,N_3126);
nand U8968 (N_8968,N_2554,N_721);
nor U8969 (N_8969,N_2017,N_1670);
nor U8970 (N_8970,N_2360,N_2411);
and U8971 (N_8971,N_313,N_308);
and U8972 (N_8972,N_2566,N_3819);
and U8973 (N_8973,N_2026,N_3665);
and U8974 (N_8974,N_1556,N_4882);
nor U8975 (N_8975,N_4188,N_2700);
and U8976 (N_8976,N_2912,N_1272);
nand U8977 (N_8977,N_1809,N_3281);
and U8978 (N_8978,N_544,N_4801);
nor U8979 (N_8979,N_3535,N_970);
and U8980 (N_8980,N_627,N_2176);
or U8981 (N_8981,N_2619,N_4087);
nand U8982 (N_8982,N_4622,N_1251);
nor U8983 (N_8983,N_2034,N_3136);
or U8984 (N_8984,N_3026,N_4237);
nor U8985 (N_8985,N_2783,N_3511);
nor U8986 (N_8986,N_3192,N_3225);
xor U8987 (N_8987,N_1297,N_35);
and U8988 (N_8988,N_4269,N_897);
and U8989 (N_8989,N_606,N_364);
nor U8990 (N_8990,N_1212,N_1660);
or U8991 (N_8991,N_37,N_755);
nor U8992 (N_8992,N_1278,N_898);
or U8993 (N_8993,N_4641,N_2081);
nand U8994 (N_8994,N_4910,N_4543);
or U8995 (N_8995,N_4254,N_2346);
nor U8996 (N_8996,N_438,N_4556);
and U8997 (N_8997,N_1747,N_4219);
nand U8998 (N_8998,N_1915,N_2372);
or U8999 (N_8999,N_4565,N_2431);
and U9000 (N_9000,N_2207,N_2287);
nand U9001 (N_9001,N_2255,N_2976);
xnor U9002 (N_9002,N_4523,N_4495);
or U9003 (N_9003,N_4535,N_4912);
xnor U9004 (N_9004,N_1962,N_3204);
and U9005 (N_9005,N_2926,N_1813);
and U9006 (N_9006,N_2340,N_1597);
nor U9007 (N_9007,N_1218,N_4270);
or U9008 (N_9008,N_2780,N_2399);
or U9009 (N_9009,N_1787,N_49);
nor U9010 (N_9010,N_79,N_4332);
nand U9011 (N_9011,N_2342,N_352);
or U9012 (N_9012,N_4439,N_1745);
nor U9013 (N_9013,N_3903,N_102);
xnor U9014 (N_9014,N_27,N_1987);
and U9015 (N_9015,N_2728,N_4440);
or U9016 (N_9016,N_1070,N_1051);
or U9017 (N_9017,N_1085,N_4059);
or U9018 (N_9018,N_2625,N_2240);
or U9019 (N_9019,N_1987,N_4862);
nor U9020 (N_9020,N_3340,N_938);
or U9021 (N_9021,N_2568,N_4555);
and U9022 (N_9022,N_4151,N_942);
or U9023 (N_9023,N_774,N_1799);
nand U9024 (N_9024,N_1710,N_1311);
nor U9025 (N_9025,N_3652,N_841);
nand U9026 (N_9026,N_1211,N_1050);
and U9027 (N_9027,N_3760,N_4329);
or U9028 (N_9028,N_2608,N_4871);
nor U9029 (N_9029,N_3545,N_1312);
nand U9030 (N_9030,N_4621,N_2419);
and U9031 (N_9031,N_1140,N_3707);
nor U9032 (N_9032,N_3678,N_1761);
nor U9033 (N_9033,N_4903,N_2387);
nand U9034 (N_9034,N_4312,N_3660);
or U9035 (N_9035,N_353,N_3770);
or U9036 (N_9036,N_1022,N_4386);
nand U9037 (N_9037,N_1316,N_1421);
nor U9038 (N_9038,N_4256,N_3580);
nor U9039 (N_9039,N_270,N_2302);
nand U9040 (N_9040,N_2043,N_3643);
nor U9041 (N_9041,N_4455,N_1045);
or U9042 (N_9042,N_21,N_4965);
and U9043 (N_9043,N_3768,N_394);
and U9044 (N_9044,N_4886,N_741);
nor U9045 (N_9045,N_4118,N_3764);
nand U9046 (N_9046,N_4163,N_3014);
and U9047 (N_9047,N_230,N_1774);
nor U9048 (N_9048,N_4487,N_1736);
or U9049 (N_9049,N_4260,N_2635);
nand U9050 (N_9050,N_1427,N_624);
nor U9051 (N_9051,N_1111,N_4833);
nand U9052 (N_9052,N_2919,N_3887);
and U9053 (N_9053,N_3698,N_4952);
nand U9054 (N_9054,N_4337,N_2564);
nor U9055 (N_9055,N_1872,N_3664);
and U9056 (N_9056,N_761,N_3461);
nor U9057 (N_9057,N_4653,N_437);
or U9058 (N_9058,N_2956,N_310);
nand U9059 (N_9059,N_3013,N_1195);
or U9060 (N_9060,N_2999,N_2256);
nor U9061 (N_9061,N_4332,N_4010);
nor U9062 (N_9062,N_1350,N_4983);
nand U9063 (N_9063,N_3998,N_4972);
nor U9064 (N_9064,N_612,N_4211);
and U9065 (N_9065,N_3566,N_1167);
nand U9066 (N_9066,N_632,N_993);
nor U9067 (N_9067,N_4851,N_815);
nand U9068 (N_9068,N_4941,N_408);
or U9069 (N_9069,N_1347,N_1235);
and U9070 (N_9070,N_1481,N_4887);
nor U9071 (N_9071,N_2479,N_2726);
nor U9072 (N_9072,N_4693,N_2045);
nand U9073 (N_9073,N_838,N_4180);
or U9074 (N_9074,N_1092,N_4737);
nor U9075 (N_9075,N_3585,N_985);
and U9076 (N_9076,N_2985,N_2995);
nor U9077 (N_9077,N_3136,N_3013);
or U9078 (N_9078,N_4771,N_535);
nand U9079 (N_9079,N_2227,N_4296);
and U9080 (N_9080,N_1738,N_375);
and U9081 (N_9081,N_1175,N_3365);
and U9082 (N_9082,N_3615,N_1786);
nor U9083 (N_9083,N_462,N_3322);
and U9084 (N_9084,N_1659,N_2382);
or U9085 (N_9085,N_1951,N_4295);
nor U9086 (N_9086,N_1561,N_815);
nor U9087 (N_9087,N_2327,N_99);
or U9088 (N_9088,N_3295,N_1107);
or U9089 (N_9089,N_4736,N_2265);
nand U9090 (N_9090,N_1394,N_4888);
and U9091 (N_9091,N_4626,N_3561);
nor U9092 (N_9092,N_3263,N_3812);
nor U9093 (N_9093,N_3882,N_1105);
nor U9094 (N_9094,N_4810,N_3891);
nor U9095 (N_9095,N_4091,N_1943);
xnor U9096 (N_9096,N_4720,N_3877);
nand U9097 (N_9097,N_970,N_258);
and U9098 (N_9098,N_3295,N_469);
nand U9099 (N_9099,N_1717,N_2959);
nor U9100 (N_9100,N_2990,N_2694);
nor U9101 (N_9101,N_4845,N_4978);
nand U9102 (N_9102,N_4254,N_515);
and U9103 (N_9103,N_1492,N_3921);
and U9104 (N_9104,N_1720,N_2004);
nand U9105 (N_9105,N_1346,N_2237);
nand U9106 (N_9106,N_2249,N_4779);
and U9107 (N_9107,N_4667,N_3373);
and U9108 (N_9108,N_4888,N_2726);
nor U9109 (N_9109,N_3143,N_558);
or U9110 (N_9110,N_2697,N_398);
nor U9111 (N_9111,N_1221,N_3862);
and U9112 (N_9112,N_3467,N_3401);
and U9113 (N_9113,N_2948,N_273);
nand U9114 (N_9114,N_1612,N_3537);
or U9115 (N_9115,N_947,N_3589);
and U9116 (N_9116,N_4090,N_2390);
nand U9117 (N_9117,N_3941,N_3867);
and U9118 (N_9118,N_3022,N_2998);
or U9119 (N_9119,N_2722,N_2561);
or U9120 (N_9120,N_1306,N_3160);
or U9121 (N_9121,N_3830,N_4112);
nor U9122 (N_9122,N_3735,N_4187);
nand U9123 (N_9123,N_3671,N_2466);
and U9124 (N_9124,N_1957,N_2260);
or U9125 (N_9125,N_1790,N_3033);
nand U9126 (N_9126,N_1581,N_176);
nand U9127 (N_9127,N_2732,N_1120);
and U9128 (N_9128,N_477,N_4402);
nor U9129 (N_9129,N_2592,N_2360);
and U9130 (N_9130,N_4919,N_3003);
nand U9131 (N_9131,N_3268,N_3308);
nor U9132 (N_9132,N_687,N_864);
nor U9133 (N_9133,N_463,N_2998);
nand U9134 (N_9134,N_1181,N_2703);
nor U9135 (N_9135,N_4824,N_4980);
and U9136 (N_9136,N_4779,N_291);
nand U9137 (N_9137,N_2722,N_4424);
and U9138 (N_9138,N_3085,N_1758);
or U9139 (N_9139,N_4248,N_4020);
and U9140 (N_9140,N_3683,N_1067);
and U9141 (N_9141,N_4860,N_740);
or U9142 (N_9142,N_1141,N_2114);
nor U9143 (N_9143,N_489,N_3995);
or U9144 (N_9144,N_1117,N_1502);
nor U9145 (N_9145,N_439,N_3718);
or U9146 (N_9146,N_322,N_4317);
nor U9147 (N_9147,N_79,N_561);
nand U9148 (N_9148,N_2128,N_4726);
and U9149 (N_9149,N_1733,N_2439);
nand U9150 (N_9150,N_4265,N_1808);
nand U9151 (N_9151,N_3396,N_1566);
or U9152 (N_9152,N_3549,N_862);
nand U9153 (N_9153,N_3628,N_2680);
nand U9154 (N_9154,N_921,N_3548);
nor U9155 (N_9155,N_3666,N_2570);
nor U9156 (N_9156,N_211,N_3835);
and U9157 (N_9157,N_778,N_3989);
or U9158 (N_9158,N_3196,N_3966);
nor U9159 (N_9159,N_2877,N_1892);
nand U9160 (N_9160,N_1454,N_536);
nand U9161 (N_9161,N_1348,N_275);
nor U9162 (N_9162,N_4005,N_4272);
nand U9163 (N_9163,N_3303,N_2713);
nand U9164 (N_9164,N_3037,N_80);
nand U9165 (N_9165,N_4295,N_1096);
nand U9166 (N_9166,N_4382,N_1148);
nand U9167 (N_9167,N_2401,N_1146);
and U9168 (N_9168,N_4407,N_1696);
nand U9169 (N_9169,N_456,N_2885);
and U9170 (N_9170,N_3935,N_4065);
and U9171 (N_9171,N_2638,N_2978);
and U9172 (N_9172,N_2701,N_4509);
and U9173 (N_9173,N_1820,N_1413);
and U9174 (N_9174,N_2511,N_2313);
nor U9175 (N_9175,N_2209,N_998);
or U9176 (N_9176,N_357,N_3638);
or U9177 (N_9177,N_4589,N_590);
nand U9178 (N_9178,N_6,N_3008);
and U9179 (N_9179,N_3729,N_366);
and U9180 (N_9180,N_4174,N_2112);
or U9181 (N_9181,N_115,N_3042);
nor U9182 (N_9182,N_3628,N_3356);
or U9183 (N_9183,N_2660,N_4901);
nand U9184 (N_9184,N_3564,N_752);
and U9185 (N_9185,N_543,N_1467);
nor U9186 (N_9186,N_2041,N_1247);
or U9187 (N_9187,N_950,N_116);
nor U9188 (N_9188,N_3069,N_2797);
or U9189 (N_9189,N_4508,N_2261);
or U9190 (N_9190,N_3106,N_2028);
nor U9191 (N_9191,N_4555,N_3049);
or U9192 (N_9192,N_4657,N_4371);
or U9193 (N_9193,N_276,N_2750);
and U9194 (N_9194,N_1832,N_4439);
or U9195 (N_9195,N_3719,N_4949);
and U9196 (N_9196,N_3000,N_976);
and U9197 (N_9197,N_3944,N_2382);
nor U9198 (N_9198,N_169,N_4438);
nand U9199 (N_9199,N_3800,N_4060);
nor U9200 (N_9200,N_3868,N_3529);
nor U9201 (N_9201,N_305,N_3292);
nand U9202 (N_9202,N_1695,N_2788);
nand U9203 (N_9203,N_4419,N_4272);
nor U9204 (N_9204,N_710,N_977);
nand U9205 (N_9205,N_2708,N_161);
nand U9206 (N_9206,N_4925,N_1972);
nor U9207 (N_9207,N_3592,N_1741);
and U9208 (N_9208,N_1575,N_1457);
xnor U9209 (N_9209,N_2862,N_3185);
nand U9210 (N_9210,N_2357,N_3792);
nor U9211 (N_9211,N_4889,N_2006);
nand U9212 (N_9212,N_4243,N_2181);
and U9213 (N_9213,N_743,N_3349);
nor U9214 (N_9214,N_2624,N_2484);
nor U9215 (N_9215,N_696,N_2000);
and U9216 (N_9216,N_1220,N_3389);
nor U9217 (N_9217,N_488,N_907);
and U9218 (N_9218,N_3834,N_706);
nor U9219 (N_9219,N_1979,N_2539);
nor U9220 (N_9220,N_2565,N_3037);
and U9221 (N_9221,N_3193,N_3606);
and U9222 (N_9222,N_754,N_2247);
or U9223 (N_9223,N_976,N_2256);
or U9224 (N_9224,N_981,N_4876);
or U9225 (N_9225,N_4512,N_837);
nor U9226 (N_9226,N_3561,N_3228);
or U9227 (N_9227,N_4770,N_549);
nand U9228 (N_9228,N_2574,N_2151);
and U9229 (N_9229,N_4257,N_641);
and U9230 (N_9230,N_4006,N_4127);
or U9231 (N_9231,N_145,N_4414);
and U9232 (N_9232,N_2853,N_1086);
nor U9233 (N_9233,N_3850,N_619);
and U9234 (N_9234,N_269,N_4449);
and U9235 (N_9235,N_4449,N_4301);
and U9236 (N_9236,N_4181,N_4714);
or U9237 (N_9237,N_207,N_4432);
nand U9238 (N_9238,N_4739,N_2238);
nor U9239 (N_9239,N_4877,N_3386);
nor U9240 (N_9240,N_4371,N_2420);
nor U9241 (N_9241,N_1613,N_2807);
nand U9242 (N_9242,N_4456,N_3075);
and U9243 (N_9243,N_2897,N_2463);
nand U9244 (N_9244,N_1514,N_3127);
nor U9245 (N_9245,N_2582,N_1029);
nor U9246 (N_9246,N_3955,N_825);
or U9247 (N_9247,N_2850,N_1925);
nor U9248 (N_9248,N_1852,N_2411);
or U9249 (N_9249,N_3586,N_290);
and U9250 (N_9250,N_3612,N_484);
nand U9251 (N_9251,N_4744,N_3408);
or U9252 (N_9252,N_3204,N_4052);
or U9253 (N_9253,N_4086,N_3363);
or U9254 (N_9254,N_3835,N_1108);
nor U9255 (N_9255,N_1120,N_113);
and U9256 (N_9256,N_3022,N_2683);
and U9257 (N_9257,N_2922,N_2406);
nor U9258 (N_9258,N_1998,N_1139);
nand U9259 (N_9259,N_1801,N_3296);
and U9260 (N_9260,N_4041,N_161);
and U9261 (N_9261,N_768,N_2236);
or U9262 (N_9262,N_643,N_1710);
nand U9263 (N_9263,N_3472,N_357);
nor U9264 (N_9264,N_1890,N_1403);
nor U9265 (N_9265,N_3435,N_4315);
nand U9266 (N_9266,N_1899,N_71);
and U9267 (N_9267,N_4584,N_1083);
or U9268 (N_9268,N_805,N_3297);
and U9269 (N_9269,N_3137,N_859);
and U9270 (N_9270,N_4616,N_1191);
nand U9271 (N_9271,N_2418,N_53);
nor U9272 (N_9272,N_1878,N_570);
and U9273 (N_9273,N_2809,N_3862);
nor U9274 (N_9274,N_1009,N_871);
nor U9275 (N_9275,N_4740,N_4701);
nand U9276 (N_9276,N_153,N_2252);
nor U9277 (N_9277,N_1657,N_4388);
nand U9278 (N_9278,N_4875,N_1436);
and U9279 (N_9279,N_2787,N_1711);
or U9280 (N_9280,N_2623,N_4508);
and U9281 (N_9281,N_3294,N_1530);
and U9282 (N_9282,N_2848,N_4278);
nand U9283 (N_9283,N_1979,N_3986);
nand U9284 (N_9284,N_225,N_1771);
and U9285 (N_9285,N_285,N_2815);
and U9286 (N_9286,N_3872,N_2175);
nor U9287 (N_9287,N_1084,N_3590);
or U9288 (N_9288,N_1410,N_3042);
nand U9289 (N_9289,N_4208,N_4168);
nand U9290 (N_9290,N_173,N_4430);
or U9291 (N_9291,N_3709,N_2875);
and U9292 (N_9292,N_3921,N_1982);
nand U9293 (N_9293,N_3266,N_2120);
nor U9294 (N_9294,N_3622,N_1178);
and U9295 (N_9295,N_3731,N_4796);
nand U9296 (N_9296,N_1300,N_2950);
and U9297 (N_9297,N_4135,N_1456);
or U9298 (N_9298,N_2782,N_3443);
or U9299 (N_9299,N_2200,N_2030);
and U9300 (N_9300,N_1681,N_2431);
or U9301 (N_9301,N_3888,N_1574);
nor U9302 (N_9302,N_478,N_2923);
or U9303 (N_9303,N_1485,N_4314);
or U9304 (N_9304,N_1033,N_4816);
nor U9305 (N_9305,N_1512,N_4018);
and U9306 (N_9306,N_4641,N_2860);
nor U9307 (N_9307,N_2304,N_3469);
or U9308 (N_9308,N_2636,N_3087);
nor U9309 (N_9309,N_1611,N_3520);
and U9310 (N_9310,N_803,N_4752);
nor U9311 (N_9311,N_2051,N_2311);
or U9312 (N_9312,N_4394,N_3787);
nor U9313 (N_9313,N_4490,N_894);
nor U9314 (N_9314,N_1784,N_3053);
nand U9315 (N_9315,N_2640,N_9);
or U9316 (N_9316,N_1041,N_1078);
or U9317 (N_9317,N_3774,N_813);
or U9318 (N_9318,N_1382,N_1197);
and U9319 (N_9319,N_2591,N_2971);
or U9320 (N_9320,N_1877,N_1738);
nor U9321 (N_9321,N_4595,N_2226);
nand U9322 (N_9322,N_2344,N_3171);
nor U9323 (N_9323,N_4370,N_589);
and U9324 (N_9324,N_1759,N_3419);
or U9325 (N_9325,N_787,N_379);
nor U9326 (N_9326,N_1432,N_155);
nor U9327 (N_9327,N_1152,N_4592);
and U9328 (N_9328,N_1852,N_1185);
or U9329 (N_9329,N_4109,N_2392);
nand U9330 (N_9330,N_3640,N_2930);
or U9331 (N_9331,N_3260,N_4590);
nand U9332 (N_9332,N_1040,N_21);
nor U9333 (N_9333,N_4646,N_4393);
and U9334 (N_9334,N_3868,N_178);
nor U9335 (N_9335,N_368,N_4995);
or U9336 (N_9336,N_3843,N_1616);
nand U9337 (N_9337,N_3936,N_728);
and U9338 (N_9338,N_1543,N_3815);
or U9339 (N_9339,N_3800,N_930);
or U9340 (N_9340,N_2342,N_533);
nor U9341 (N_9341,N_666,N_4091);
or U9342 (N_9342,N_2249,N_4776);
nand U9343 (N_9343,N_2855,N_2086);
xnor U9344 (N_9344,N_4179,N_3044);
nand U9345 (N_9345,N_254,N_4066);
and U9346 (N_9346,N_3533,N_224);
or U9347 (N_9347,N_121,N_899);
nand U9348 (N_9348,N_3415,N_3201);
or U9349 (N_9349,N_4844,N_4091);
nand U9350 (N_9350,N_1295,N_389);
or U9351 (N_9351,N_1766,N_1618);
xor U9352 (N_9352,N_4278,N_1195);
and U9353 (N_9353,N_2655,N_1368);
or U9354 (N_9354,N_925,N_4853);
nor U9355 (N_9355,N_4762,N_3798);
and U9356 (N_9356,N_1318,N_43);
or U9357 (N_9357,N_1852,N_1466);
and U9358 (N_9358,N_2205,N_3872);
or U9359 (N_9359,N_1323,N_4069);
nor U9360 (N_9360,N_1778,N_363);
and U9361 (N_9361,N_3936,N_1428);
and U9362 (N_9362,N_584,N_1645);
nor U9363 (N_9363,N_2906,N_1910);
or U9364 (N_9364,N_4146,N_3829);
and U9365 (N_9365,N_3563,N_1488);
nor U9366 (N_9366,N_2049,N_79);
or U9367 (N_9367,N_223,N_2735);
and U9368 (N_9368,N_1539,N_452);
nor U9369 (N_9369,N_310,N_4173);
nor U9370 (N_9370,N_2783,N_1479);
or U9371 (N_9371,N_372,N_2039);
nand U9372 (N_9372,N_3762,N_3489);
or U9373 (N_9373,N_1343,N_4919);
nor U9374 (N_9374,N_704,N_107);
nor U9375 (N_9375,N_2055,N_2412);
and U9376 (N_9376,N_1506,N_2655);
and U9377 (N_9377,N_3793,N_942);
and U9378 (N_9378,N_3259,N_4126);
nor U9379 (N_9379,N_41,N_3516);
and U9380 (N_9380,N_244,N_233);
or U9381 (N_9381,N_1510,N_820);
nor U9382 (N_9382,N_1890,N_2941);
nand U9383 (N_9383,N_4003,N_1138);
nor U9384 (N_9384,N_3116,N_1424);
nand U9385 (N_9385,N_965,N_3825);
nor U9386 (N_9386,N_975,N_2489);
nand U9387 (N_9387,N_367,N_1259);
nand U9388 (N_9388,N_805,N_2760);
nand U9389 (N_9389,N_2904,N_427);
or U9390 (N_9390,N_4496,N_1586);
xor U9391 (N_9391,N_1129,N_3123);
nor U9392 (N_9392,N_3617,N_3369);
nand U9393 (N_9393,N_4594,N_1056);
nand U9394 (N_9394,N_4864,N_3847);
nand U9395 (N_9395,N_36,N_2784);
nand U9396 (N_9396,N_2269,N_2853);
nor U9397 (N_9397,N_4576,N_2042);
and U9398 (N_9398,N_1633,N_2589);
and U9399 (N_9399,N_4705,N_3110);
nand U9400 (N_9400,N_798,N_381);
xnor U9401 (N_9401,N_807,N_4696);
nand U9402 (N_9402,N_4281,N_861);
or U9403 (N_9403,N_2092,N_3630);
or U9404 (N_9404,N_2212,N_4012);
or U9405 (N_9405,N_3389,N_4115);
xnor U9406 (N_9406,N_366,N_3675);
nand U9407 (N_9407,N_2934,N_4851);
or U9408 (N_9408,N_4709,N_287);
nor U9409 (N_9409,N_2791,N_3308);
and U9410 (N_9410,N_2582,N_1099);
nand U9411 (N_9411,N_1321,N_4929);
and U9412 (N_9412,N_1201,N_2487);
or U9413 (N_9413,N_1546,N_2679);
nor U9414 (N_9414,N_3569,N_3648);
nor U9415 (N_9415,N_2372,N_2144);
and U9416 (N_9416,N_3054,N_3100);
and U9417 (N_9417,N_553,N_4917);
and U9418 (N_9418,N_100,N_3345);
and U9419 (N_9419,N_3988,N_2407);
nand U9420 (N_9420,N_4221,N_2737);
nor U9421 (N_9421,N_3038,N_3896);
or U9422 (N_9422,N_3875,N_1740);
nor U9423 (N_9423,N_1999,N_325);
and U9424 (N_9424,N_3934,N_4974);
nand U9425 (N_9425,N_2182,N_2161);
or U9426 (N_9426,N_3914,N_3942);
nor U9427 (N_9427,N_2307,N_4249);
nor U9428 (N_9428,N_306,N_3939);
and U9429 (N_9429,N_2390,N_2138);
and U9430 (N_9430,N_1236,N_84);
and U9431 (N_9431,N_272,N_1028);
or U9432 (N_9432,N_723,N_2803);
nand U9433 (N_9433,N_1114,N_4006);
nand U9434 (N_9434,N_4623,N_4583);
and U9435 (N_9435,N_1825,N_3814);
nand U9436 (N_9436,N_4874,N_1972);
nand U9437 (N_9437,N_2760,N_3592);
and U9438 (N_9438,N_2776,N_4521);
nor U9439 (N_9439,N_100,N_3654);
or U9440 (N_9440,N_2844,N_420);
nor U9441 (N_9441,N_4467,N_2216);
nand U9442 (N_9442,N_375,N_1005);
and U9443 (N_9443,N_985,N_4972);
or U9444 (N_9444,N_2210,N_3179);
nand U9445 (N_9445,N_583,N_4312);
nand U9446 (N_9446,N_3166,N_1321);
and U9447 (N_9447,N_483,N_772);
nand U9448 (N_9448,N_263,N_2814);
and U9449 (N_9449,N_3126,N_1197);
nand U9450 (N_9450,N_2531,N_2804);
and U9451 (N_9451,N_2434,N_3186);
or U9452 (N_9452,N_4030,N_4969);
or U9453 (N_9453,N_3952,N_599);
nand U9454 (N_9454,N_4955,N_864);
or U9455 (N_9455,N_2093,N_441);
or U9456 (N_9456,N_3834,N_458);
nor U9457 (N_9457,N_4662,N_4708);
and U9458 (N_9458,N_3905,N_920);
xnor U9459 (N_9459,N_1037,N_2159);
or U9460 (N_9460,N_2618,N_2175);
nor U9461 (N_9461,N_2894,N_2670);
and U9462 (N_9462,N_4237,N_1196);
nand U9463 (N_9463,N_2401,N_2778);
nor U9464 (N_9464,N_1231,N_1784);
or U9465 (N_9465,N_3618,N_3532);
nand U9466 (N_9466,N_46,N_655);
and U9467 (N_9467,N_1236,N_2571);
or U9468 (N_9468,N_151,N_2414);
nand U9469 (N_9469,N_224,N_2296);
and U9470 (N_9470,N_292,N_1711);
nand U9471 (N_9471,N_883,N_1393);
or U9472 (N_9472,N_2638,N_4008);
or U9473 (N_9473,N_1291,N_1155);
and U9474 (N_9474,N_2343,N_4697);
nand U9475 (N_9475,N_295,N_155);
or U9476 (N_9476,N_1597,N_2610);
and U9477 (N_9477,N_3164,N_1770);
or U9478 (N_9478,N_1181,N_3046);
nand U9479 (N_9479,N_3720,N_3686);
nand U9480 (N_9480,N_10,N_406);
nor U9481 (N_9481,N_1884,N_1413);
nand U9482 (N_9482,N_1897,N_3506);
and U9483 (N_9483,N_1467,N_2766);
nand U9484 (N_9484,N_3923,N_3374);
or U9485 (N_9485,N_788,N_4473);
nand U9486 (N_9486,N_3232,N_2651);
and U9487 (N_9487,N_3907,N_320);
nor U9488 (N_9488,N_992,N_1204);
or U9489 (N_9489,N_2661,N_2891);
nand U9490 (N_9490,N_11,N_4795);
nand U9491 (N_9491,N_4438,N_3214);
nor U9492 (N_9492,N_4685,N_648);
nand U9493 (N_9493,N_1737,N_2098);
or U9494 (N_9494,N_1,N_2585);
and U9495 (N_9495,N_1966,N_4031);
and U9496 (N_9496,N_2623,N_4606);
or U9497 (N_9497,N_2478,N_866);
nand U9498 (N_9498,N_703,N_4687);
nor U9499 (N_9499,N_1743,N_1411);
nand U9500 (N_9500,N_2032,N_119);
nor U9501 (N_9501,N_3630,N_3381);
and U9502 (N_9502,N_986,N_1623);
and U9503 (N_9503,N_2163,N_415);
and U9504 (N_9504,N_3456,N_2654);
and U9505 (N_9505,N_4893,N_4766);
nand U9506 (N_9506,N_2939,N_880);
or U9507 (N_9507,N_805,N_4643);
or U9508 (N_9508,N_897,N_401);
xnor U9509 (N_9509,N_1586,N_3962);
nor U9510 (N_9510,N_3879,N_673);
nand U9511 (N_9511,N_352,N_4294);
and U9512 (N_9512,N_177,N_623);
or U9513 (N_9513,N_122,N_2623);
nand U9514 (N_9514,N_3247,N_249);
or U9515 (N_9515,N_3268,N_2681);
nor U9516 (N_9516,N_8,N_3672);
nor U9517 (N_9517,N_3365,N_3357);
and U9518 (N_9518,N_2417,N_2246);
nand U9519 (N_9519,N_2275,N_1098);
nor U9520 (N_9520,N_2713,N_692);
nand U9521 (N_9521,N_167,N_928);
nor U9522 (N_9522,N_442,N_955);
nor U9523 (N_9523,N_4562,N_148);
nor U9524 (N_9524,N_1030,N_310);
nor U9525 (N_9525,N_3232,N_3895);
nand U9526 (N_9526,N_2523,N_4965);
nand U9527 (N_9527,N_3055,N_66);
nor U9528 (N_9528,N_135,N_4308);
nor U9529 (N_9529,N_3244,N_4128);
xor U9530 (N_9530,N_1807,N_1076);
and U9531 (N_9531,N_1093,N_972);
and U9532 (N_9532,N_3030,N_4539);
nor U9533 (N_9533,N_4117,N_1843);
nand U9534 (N_9534,N_3267,N_4699);
nand U9535 (N_9535,N_1801,N_1159);
nand U9536 (N_9536,N_4535,N_3399);
or U9537 (N_9537,N_3879,N_2220);
or U9538 (N_9538,N_514,N_2407);
or U9539 (N_9539,N_1431,N_4403);
and U9540 (N_9540,N_3978,N_539);
or U9541 (N_9541,N_3323,N_1665);
nor U9542 (N_9542,N_4201,N_1681);
nor U9543 (N_9543,N_4884,N_2955);
or U9544 (N_9544,N_3945,N_2598);
nand U9545 (N_9545,N_4610,N_1933);
nand U9546 (N_9546,N_817,N_4865);
nand U9547 (N_9547,N_1271,N_272);
or U9548 (N_9548,N_3344,N_4256);
and U9549 (N_9549,N_3189,N_2683);
nand U9550 (N_9550,N_147,N_2548);
or U9551 (N_9551,N_95,N_1569);
nor U9552 (N_9552,N_1098,N_3112);
nor U9553 (N_9553,N_657,N_3900);
nor U9554 (N_9554,N_2403,N_2);
and U9555 (N_9555,N_1791,N_4159);
nand U9556 (N_9556,N_3777,N_693);
nor U9557 (N_9557,N_2136,N_3799);
or U9558 (N_9558,N_3000,N_2263);
and U9559 (N_9559,N_42,N_819);
nor U9560 (N_9560,N_2412,N_2471);
nor U9561 (N_9561,N_4856,N_1949);
nand U9562 (N_9562,N_1113,N_3587);
and U9563 (N_9563,N_3731,N_1278);
and U9564 (N_9564,N_3215,N_1268);
and U9565 (N_9565,N_2168,N_576);
and U9566 (N_9566,N_871,N_1220);
nor U9567 (N_9567,N_878,N_2452);
nor U9568 (N_9568,N_3781,N_3670);
nand U9569 (N_9569,N_4968,N_2957);
or U9570 (N_9570,N_2177,N_997);
nand U9571 (N_9571,N_725,N_653);
nor U9572 (N_9572,N_592,N_4530);
nand U9573 (N_9573,N_535,N_3317);
and U9574 (N_9574,N_2475,N_4047);
or U9575 (N_9575,N_2967,N_4271);
and U9576 (N_9576,N_500,N_1266);
nor U9577 (N_9577,N_514,N_3316);
nand U9578 (N_9578,N_2933,N_3394);
and U9579 (N_9579,N_4870,N_2592);
nor U9580 (N_9580,N_1966,N_3209);
or U9581 (N_9581,N_681,N_298);
and U9582 (N_9582,N_1905,N_216);
or U9583 (N_9583,N_3366,N_3522);
nand U9584 (N_9584,N_1631,N_1562);
nand U9585 (N_9585,N_4132,N_1938);
and U9586 (N_9586,N_4159,N_2136);
or U9587 (N_9587,N_866,N_3805);
or U9588 (N_9588,N_2332,N_1362);
nand U9589 (N_9589,N_1016,N_4993);
nand U9590 (N_9590,N_4601,N_1036);
nand U9591 (N_9591,N_1819,N_3452);
and U9592 (N_9592,N_3517,N_2815);
nor U9593 (N_9593,N_4524,N_4555);
nand U9594 (N_9594,N_4859,N_933);
nor U9595 (N_9595,N_4634,N_1713);
or U9596 (N_9596,N_4308,N_1666);
nor U9597 (N_9597,N_2673,N_3983);
nand U9598 (N_9598,N_826,N_2531);
nor U9599 (N_9599,N_1423,N_1160);
nor U9600 (N_9600,N_3798,N_3162);
or U9601 (N_9601,N_2885,N_487);
and U9602 (N_9602,N_3304,N_640);
or U9603 (N_9603,N_1702,N_3184);
nor U9604 (N_9604,N_2856,N_2878);
or U9605 (N_9605,N_3034,N_2800);
or U9606 (N_9606,N_2399,N_4569);
nand U9607 (N_9607,N_1295,N_1588);
or U9608 (N_9608,N_4783,N_1292);
or U9609 (N_9609,N_3221,N_1059);
nor U9610 (N_9610,N_3788,N_2639);
and U9611 (N_9611,N_941,N_2724);
nor U9612 (N_9612,N_3278,N_2862);
nor U9613 (N_9613,N_3497,N_2184);
nand U9614 (N_9614,N_2208,N_3775);
nand U9615 (N_9615,N_1112,N_4207);
nand U9616 (N_9616,N_173,N_2099);
nand U9617 (N_9617,N_206,N_2398);
nand U9618 (N_9618,N_464,N_1154);
nor U9619 (N_9619,N_2638,N_3600);
nor U9620 (N_9620,N_1776,N_1875);
or U9621 (N_9621,N_104,N_4314);
or U9622 (N_9622,N_4291,N_3116);
nor U9623 (N_9623,N_2187,N_2306);
nor U9624 (N_9624,N_4974,N_2223);
and U9625 (N_9625,N_381,N_1818);
and U9626 (N_9626,N_3916,N_2329);
or U9627 (N_9627,N_3955,N_3281);
or U9628 (N_9628,N_1148,N_3138);
or U9629 (N_9629,N_3489,N_4290);
and U9630 (N_9630,N_4466,N_2780);
nor U9631 (N_9631,N_343,N_388);
nand U9632 (N_9632,N_2952,N_2050);
nand U9633 (N_9633,N_4206,N_2937);
and U9634 (N_9634,N_1689,N_1926);
and U9635 (N_9635,N_3902,N_4727);
and U9636 (N_9636,N_2376,N_2613);
and U9637 (N_9637,N_4024,N_3023);
or U9638 (N_9638,N_2132,N_4513);
nor U9639 (N_9639,N_701,N_939);
nor U9640 (N_9640,N_3933,N_2236);
nor U9641 (N_9641,N_3566,N_1371);
nor U9642 (N_9642,N_3062,N_3824);
nor U9643 (N_9643,N_4708,N_3700);
or U9644 (N_9644,N_121,N_2713);
nand U9645 (N_9645,N_4171,N_2134);
nand U9646 (N_9646,N_1756,N_1380);
and U9647 (N_9647,N_278,N_435);
and U9648 (N_9648,N_1991,N_1429);
or U9649 (N_9649,N_4306,N_866);
or U9650 (N_9650,N_4511,N_2470);
and U9651 (N_9651,N_2838,N_3995);
nand U9652 (N_9652,N_4186,N_2868);
or U9653 (N_9653,N_1291,N_1965);
nand U9654 (N_9654,N_2261,N_4181);
nor U9655 (N_9655,N_2923,N_411);
xor U9656 (N_9656,N_4748,N_1377);
nand U9657 (N_9657,N_2110,N_1581);
or U9658 (N_9658,N_39,N_3880);
and U9659 (N_9659,N_4913,N_918);
and U9660 (N_9660,N_2778,N_2174);
nand U9661 (N_9661,N_3708,N_2146);
and U9662 (N_9662,N_4434,N_914);
nor U9663 (N_9663,N_4789,N_4344);
or U9664 (N_9664,N_4225,N_2056);
or U9665 (N_9665,N_4079,N_3824);
nand U9666 (N_9666,N_1374,N_1538);
nand U9667 (N_9667,N_2501,N_805);
and U9668 (N_9668,N_1460,N_4795);
nand U9669 (N_9669,N_2631,N_4669);
or U9670 (N_9670,N_651,N_1610);
and U9671 (N_9671,N_4355,N_1026);
nand U9672 (N_9672,N_2034,N_669);
nand U9673 (N_9673,N_1486,N_62);
and U9674 (N_9674,N_1676,N_4334);
and U9675 (N_9675,N_630,N_4929);
or U9676 (N_9676,N_1159,N_3450);
nor U9677 (N_9677,N_350,N_4755);
nor U9678 (N_9678,N_3289,N_4870);
nand U9679 (N_9679,N_2252,N_2824);
nand U9680 (N_9680,N_1898,N_3489);
nor U9681 (N_9681,N_3147,N_734);
nor U9682 (N_9682,N_906,N_3914);
and U9683 (N_9683,N_1834,N_4434);
nand U9684 (N_9684,N_317,N_3867);
and U9685 (N_9685,N_3497,N_2276);
nand U9686 (N_9686,N_4404,N_342);
or U9687 (N_9687,N_4509,N_3273);
and U9688 (N_9688,N_3567,N_3806);
or U9689 (N_9689,N_3065,N_4927);
nor U9690 (N_9690,N_1949,N_4013);
nand U9691 (N_9691,N_3181,N_2563);
and U9692 (N_9692,N_3403,N_3954);
nand U9693 (N_9693,N_4853,N_2458);
nor U9694 (N_9694,N_2543,N_3473);
nor U9695 (N_9695,N_2977,N_4581);
or U9696 (N_9696,N_836,N_724);
nand U9697 (N_9697,N_2585,N_1110);
nor U9698 (N_9698,N_3940,N_3028);
and U9699 (N_9699,N_4569,N_1449);
or U9700 (N_9700,N_2856,N_1791);
and U9701 (N_9701,N_4081,N_2157);
nor U9702 (N_9702,N_3738,N_3071);
nand U9703 (N_9703,N_3320,N_4316);
nand U9704 (N_9704,N_2044,N_1411);
or U9705 (N_9705,N_2581,N_643);
and U9706 (N_9706,N_4228,N_1914);
nor U9707 (N_9707,N_4477,N_1749);
and U9708 (N_9708,N_3161,N_531);
nand U9709 (N_9709,N_2155,N_3119);
or U9710 (N_9710,N_4537,N_912);
and U9711 (N_9711,N_3254,N_4864);
nor U9712 (N_9712,N_3520,N_4819);
or U9713 (N_9713,N_4540,N_2463);
nor U9714 (N_9714,N_2041,N_3706);
or U9715 (N_9715,N_269,N_3410);
or U9716 (N_9716,N_534,N_884);
nand U9717 (N_9717,N_817,N_3602);
nor U9718 (N_9718,N_2614,N_1317);
and U9719 (N_9719,N_860,N_1703);
and U9720 (N_9720,N_867,N_4191);
or U9721 (N_9721,N_837,N_3062);
and U9722 (N_9722,N_4041,N_1738);
and U9723 (N_9723,N_2186,N_660);
and U9724 (N_9724,N_678,N_4101);
or U9725 (N_9725,N_4724,N_3114);
or U9726 (N_9726,N_2818,N_4967);
nor U9727 (N_9727,N_1214,N_4744);
and U9728 (N_9728,N_3688,N_2364);
nor U9729 (N_9729,N_358,N_4272);
nand U9730 (N_9730,N_4411,N_1857);
nor U9731 (N_9731,N_2166,N_154);
nor U9732 (N_9732,N_2856,N_1536);
and U9733 (N_9733,N_3089,N_2609);
or U9734 (N_9734,N_3839,N_4264);
or U9735 (N_9735,N_2154,N_4471);
and U9736 (N_9736,N_2257,N_2186);
nand U9737 (N_9737,N_1422,N_2647);
and U9738 (N_9738,N_210,N_3192);
and U9739 (N_9739,N_3014,N_3301);
nor U9740 (N_9740,N_4130,N_2837);
and U9741 (N_9741,N_4643,N_3795);
nor U9742 (N_9742,N_4056,N_2515);
nand U9743 (N_9743,N_3821,N_719);
or U9744 (N_9744,N_1422,N_1001);
nor U9745 (N_9745,N_4395,N_1863);
and U9746 (N_9746,N_4409,N_3929);
and U9747 (N_9747,N_617,N_2824);
or U9748 (N_9748,N_668,N_2853);
nand U9749 (N_9749,N_4835,N_2151);
nor U9750 (N_9750,N_3167,N_993);
nand U9751 (N_9751,N_169,N_4321);
or U9752 (N_9752,N_1347,N_3074);
nor U9753 (N_9753,N_3732,N_2830);
nor U9754 (N_9754,N_491,N_4611);
and U9755 (N_9755,N_1415,N_4597);
nand U9756 (N_9756,N_589,N_409);
nand U9757 (N_9757,N_3159,N_1391);
nand U9758 (N_9758,N_3547,N_2747);
or U9759 (N_9759,N_204,N_4563);
or U9760 (N_9760,N_920,N_2164);
and U9761 (N_9761,N_3311,N_1086);
or U9762 (N_9762,N_444,N_3906);
nor U9763 (N_9763,N_4398,N_3802);
or U9764 (N_9764,N_141,N_4615);
nor U9765 (N_9765,N_1553,N_1472);
nor U9766 (N_9766,N_1007,N_3558);
and U9767 (N_9767,N_3833,N_3933);
nor U9768 (N_9768,N_4408,N_3082);
nand U9769 (N_9769,N_4139,N_3573);
nor U9770 (N_9770,N_2216,N_1441);
or U9771 (N_9771,N_2675,N_4261);
nor U9772 (N_9772,N_2473,N_2020);
nor U9773 (N_9773,N_750,N_2238);
or U9774 (N_9774,N_2570,N_2555);
or U9775 (N_9775,N_3059,N_2403);
nor U9776 (N_9776,N_2520,N_3135);
nand U9777 (N_9777,N_74,N_1132);
nor U9778 (N_9778,N_2399,N_4077);
or U9779 (N_9779,N_386,N_1884);
or U9780 (N_9780,N_583,N_2722);
xor U9781 (N_9781,N_2452,N_3798);
nor U9782 (N_9782,N_1800,N_4306);
or U9783 (N_9783,N_405,N_3552);
nand U9784 (N_9784,N_3965,N_4904);
or U9785 (N_9785,N_403,N_405);
and U9786 (N_9786,N_2449,N_4007);
or U9787 (N_9787,N_2495,N_377);
nand U9788 (N_9788,N_4113,N_3212);
and U9789 (N_9789,N_471,N_3066);
nor U9790 (N_9790,N_110,N_2847);
and U9791 (N_9791,N_2772,N_2252);
and U9792 (N_9792,N_2061,N_2770);
nor U9793 (N_9793,N_3662,N_508);
nand U9794 (N_9794,N_1140,N_732);
nor U9795 (N_9795,N_3239,N_2077);
nor U9796 (N_9796,N_4665,N_4120);
nand U9797 (N_9797,N_4122,N_4991);
nor U9798 (N_9798,N_842,N_2893);
or U9799 (N_9799,N_3604,N_2681);
xor U9800 (N_9800,N_3597,N_2846);
nor U9801 (N_9801,N_4973,N_4440);
and U9802 (N_9802,N_4990,N_712);
or U9803 (N_9803,N_2143,N_507);
nand U9804 (N_9804,N_4134,N_421);
nand U9805 (N_9805,N_2445,N_3001);
nand U9806 (N_9806,N_20,N_3458);
or U9807 (N_9807,N_3842,N_4866);
and U9808 (N_9808,N_543,N_338);
and U9809 (N_9809,N_2425,N_1137);
or U9810 (N_9810,N_863,N_3556);
or U9811 (N_9811,N_1080,N_211);
and U9812 (N_9812,N_1334,N_2429);
and U9813 (N_9813,N_4843,N_758);
and U9814 (N_9814,N_4411,N_3231);
and U9815 (N_9815,N_4721,N_4867);
and U9816 (N_9816,N_2718,N_860);
nor U9817 (N_9817,N_1722,N_4866);
and U9818 (N_9818,N_4182,N_2899);
nor U9819 (N_9819,N_296,N_2963);
nor U9820 (N_9820,N_384,N_3749);
nand U9821 (N_9821,N_4785,N_1450);
nor U9822 (N_9822,N_3136,N_2381);
nor U9823 (N_9823,N_647,N_4567);
or U9824 (N_9824,N_230,N_2897);
nand U9825 (N_9825,N_1586,N_808);
or U9826 (N_9826,N_153,N_2545);
nor U9827 (N_9827,N_307,N_1533);
nand U9828 (N_9828,N_1992,N_50);
or U9829 (N_9829,N_71,N_4508);
nor U9830 (N_9830,N_4962,N_1749);
or U9831 (N_9831,N_1624,N_3413);
or U9832 (N_9832,N_2954,N_2888);
nand U9833 (N_9833,N_3232,N_1758);
or U9834 (N_9834,N_1110,N_1319);
or U9835 (N_9835,N_253,N_2304);
nand U9836 (N_9836,N_2545,N_4805);
nor U9837 (N_9837,N_386,N_726);
or U9838 (N_9838,N_4046,N_442);
or U9839 (N_9839,N_2401,N_3472);
or U9840 (N_9840,N_2329,N_703);
or U9841 (N_9841,N_547,N_1936);
and U9842 (N_9842,N_1665,N_4773);
nand U9843 (N_9843,N_2849,N_2682);
or U9844 (N_9844,N_455,N_4833);
nand U9845 (N_9845,N_2696,N_3320);
and U9846 (N_9846,N_1075,N_3181);
nor U9847 (N_9847,N_4851,N_4250);
nand U9848 (N_9848,N_1330,N_4011);
nand U9849 (N_9849,N_2538,N_4714);
nand U9850 (N_9850,N_1667,N_2947);
nor U9851 (N_9851,N_3964,N_4447);
and U9852 (N_9852,N_65,N_4634);
or U9853 (N_9853,N_325,N_2285);
or U9854 (N_9854,N_1391,N_460);
nor U9855 (N_9855,N_4878,N_3962);
nor U9856 (N_9856,N_3770,N_1969);
or U9857 (N_9857,N_4867,N_4941);
and U9858 (N_9858,N_2109,N_149);
or U9859 (N_9859,N_3667,N_3975);
nand U9860 (N_9860,N_3721,N_1064);
and U9861 (N_9861,N_174,N_1654);
nand U9862 (N_9862,N_2708,N_780);
or U9863 (N_9863,N_4978,N_2689);
nand U9864 (N_9864,N_3100,N_3319);
nor U9865 (N_9865,N_3626,N_1963);
and U9866 (N_9866,N_1189,N_2445);
and U9867 (N_9867,N_510,N_1263);
nor U9868 (N_9868,N_4713,N_3507);
and U9869 (N_9869,N_1051,N_1744);
nand U9870 (N_9870,N_1202,N_4687);
and U9871 (N_9871,N_2831,N_1451);
and U9872 (N_9872,N_4860,N_454);
nand U9873 (N_9873,N_2113,N_3821);
nand U9874 (N_9874,N_244,N_488);
and U9875 (N_9875,N_1458,N_3120);
nand U9876 (N_9876,N_943,N_2707);
and U9877 (N_9877,N_2998,N_3521);
nor U9878 (N_9878,N_2561,N_1585);
and U9879 (N_9879,N_2137,N_2555);
nor U9880 (N_9880,N_4915,N_2018);
and U9881 (N_9881,N_266,N_4088);
or U9882 (N_9882,N_246,N_2283);
and U9883 (N_9883,N_1444,N_4646);
or U9884 (N_9884,N_4828,N_4116);
and U9885 (N_9885,N_4708,N_1869);
and U9886 (N_9886,N_2948,N_3055);
and U9887 (N_9887,N_1164,N_3609);
or U9888 (N_9888,N_4307,N_2803);
nor U9889 (N_9889,N_39,N_4371);
nand U9890 (N_9890,N_775,N_761);
nor U9891 (N_9891,N_2490,N_3032);
nand U9892 (N_9892,N_1918,N_1748);
and U9893 (N_9893,N_2692,N_2759);
nor U9894 (N_9894,N_3684,N_4586);
nor U9895 (N_9895,N_1220,N_800);
nor U9896 (N_9896,N_2241,N_402);
or U9897 (N_9897,N_468,N_3980);
nand U9898 (N_9898,N_3170,N_1848);
nor U9899 (N_9899,N_3856,N_4392);
nand U9900 (N_9900,N_4209,N_3436);
nor U9901 (N_9901,N_710,N_3300);
or U9902 (N_9902,N_1420,N_928);
or U9903 (N_9903,N_3107,N_3203);
nand U9904 (N_9904,N_4771,N_2328);
nor U9905 (N_9905,N_4065,N_2775);
or U9906 (N_9906,N_1474,N_2303);
nor U9907 (N_9907,N_3875,N_555);
or U9908 (N_9908,N_2959,N_220);
and U9909 (N_9909,N_2006,N_4777);
nand U9910 (N_9910,N_2414,N_3524);
nor U9911 (N_9911,N_4217,N_3879);
and U9912 (N_9912,N_1268,N_3197);
nor U9913 (N_9913,N_3057,N_1447);
nor U9914 (N_9914,N_2514,N_2563);
and U9915 (N_9915,N_2874,N_1577);
and U9916 (N_9916,N_4885,N_2913);
nand U9917 (N_9917,N_383,N_4899);
and U9918 (N_9918,N_4212,N_4676);
or U9919 (N_9919,N_1192,N_3667);
or U9920 (N_9920,N_4531,N_940);
and U9921 (N_9921,N_1113,N_318);
or U9922 (N_9922,N_4270,N_3025);
or U9923 (N_9923,N_1571,N_523);
and U9924 (N_9924,N_227,N_2765);
nor U9925 (N_9925,N_2560,N_3843);
nand U9926 (N_9926,N_2757,N_4051);
nand U9927 (N_9927,N_3999,N_2062);
or U9928 (N_9928,N_3066,N_1333);
or U9929 (N_9929,N_1231,N_798);
nor U9930 (N_9930,N_4132,N_3049);
or U9931 (N_9931,N_4643,N_2965);
or U9932 (N_9932,N_1912,N_562);
or U9933 (N_9933,N_1373,N_3605);
nand U9934 (N_9934,N_4199,N_4844);
and U9935 (N_9935,N_2389,N_3506);
nor U9936 (N_9936,N_4889,N_2104);
or U9937 (N_9937,N_1038,N_1336);
or U9938 (N_9938,N_3969,N_2233);
or U9939 (N_9939,N_2106,N_356);
or U9940 (N_9940,N_3040,N_3920);
or U9941 (N_9941,N_1524,N_291);
and U9942 (N_9942,N_2697,N_3884);
and U9943 (N_9943,N_2286,N_2445);
and U9944 (N_9944,N_1838,N_3065);
and U9945 (N_9945,N_3113,N_1205);
nor U9946 (N_9946,N_1733,N_1415);
and U9947 (N_9947,N_925,N_3183);
nand U9948 (N_9948,N_114,N_900);
or U9949 (N_9949,N_4812,N_4315);
and U9950 (N_9950,N_667,N_916);
nand U9951 (N_9951,N_4104,N_483);
or U9952 (N_9952,N_567,N_3546);
nor U9953 (N_9953,N_931,N_2268);
or U9954 (N_9954,N_3502,N_2777);
xor U9955 (N_9955,N_1651,N_4645);
and U9956 (N_9956,N_1607,N_4677);
or U9957 (N_9957,N_156,N_230);
and U9958 (N_9958,N_4833,N_4399);
or U9959 (N_9959,N_3630,N_986);
nand U9960 (N_9960,N_3695,N_2189);
nor U9961 (N_9961,N_4269,N_776);
or U9962 (N_9962,N_4754,N_195);
or U9963 (N_9963,N_2238,N_3959);
and U9964 (N_9964,N_536,N_3139);
or U9965 (N_9965,N_3240,N_3365);
and U9966 (N_9966,N_67,N_1263);
nand U9967 (N_9967,N_4984,N_118);
nand U9968 (N_9968,N_1863,N_4739);
and U9969 (N_9969,N_4843,N_3279);
nor U9970 (N_9970,N_2567,N_1477);
nor U9971 (N_9971,N_3622,N_4883);
or U9972 (N_9972,N_4021,N_1267);
nand U9973 (N_9973,N_2558,N_2849);
nor U9974 (N_9974,N_964,N_1163);
or U9975 (N_9975,N_1777,N_1594);
xnor U9976 (N_9976,N_1933,N_1429);
nor U9977 (N_9977,N_3731,N_4587);
nand U9978 (N_9978,N_3162,N_579);
and U9979 (N_9979,N_3660,N_1228);
nand U9980 (N_9980,N_3037,N_1381);
nor U9981 (N_9981,N_3954,N_3278);
and U9982 (N_9982,N_634,N_4239);
nor U9983 (N_9983,N_3345,N_4936);
and U9984 (N_9984,N_4408,N_1083);
nand U9985 (N_9985,N_4278,N_3775);
nand U9986 (N_9986,N_3871,N_1538);
or U9987 (N_9987,N_3875,N_2205);
or U9988 (N_9988,N_1434,N_1700);
and U9989 (N_9989,N_519,N_119);
or U9990 (N_9990,N_2552,N_2252);
nor U9991 (N_9991,N_1269,N_2737);
or U9992 (N_9992,N_3921,N_4431);
nand U9993 (N_9993,N_4200,N_2645);
or U9994 (N_9994,N_3195,N_600);
and U9995 (N_9995,N_3711,N_4854);
nor U9996 (N_9996,N_1022,N_4155);
nand U9997 (N_9997,N_2861,N_3179);
or U9998 (N_9998,N_356,N_3088);
nand U9999 (N_9999,N_4856,N_3264);
or U10000 (N_10000,N_6874,N_9335);
or U10001 (N_10001,N_6099,N_7212);
nand U10002 (N_10002,N_9344,N_5473);
and U10003 (N_10003,N_5046,N_5674);
nor U10004 (N_10004,N_5508,N_9253);
and U10005 (N_10005,N_5227,N_8177);
nor U10006 (N_10006,N_6338,N_5908);
and U10007 (N_10007,N_9265,N_8641);
or U10008 (N_10008,N_7176,N_9180);
nor U10009 (N_10009,N_9321,N_5417);
or U10010 (N_10010,N_8821,N_6981);
and U10011 (N_10011,N_6899,N_6503);
and U10012 (N_10012,N_6204,N_7437);
or U10013 (N_10013,N_5540,N_7477);
nand U10014 (N_10014,N_6571,N_8661);
nor U10015 (N_10015,N_5468,N_7878);
or U10016 (N_10016,N_7162,N_9067);
nor U10017 (N_10017,N_7155,N_6404);
or U10018 (N_10018,N_5048,N_8590);
nor U10019 (N_10019,N_9743,N_7194);
and U10020 (N_10020,N_5056,N_6812);
nor U10021 (N_10021,N_6700,N_7684);
nand U10022 (N_10022,N_9858,N_7959);
nand U10023 (N_10023,N_8147,N_6027);
nor U10024 (N_10024,N_8395,N_5743);
and U10025 (N_10025,N_9832,N_8600);
nor U10026 (N_10026,N_5941,N_5856);
or U10027 (N_10027,N_6472,N_8095);
nor U10028 (N_10028,N_9699,N_7356);
nand U10029 (N_10029,N_5442,N_7998);
or U10030 (N_10030,N_7943,N_7106);
and U10031 (N_10031,N_6672,N_9276);
or U10032 (N_10032,N_5357,N_9234);
nand U10033 (N_10033,N_8328,N_7785);
or U10034 (N_10034,N_9838,N_7593);
nor U10035 (N_10035,N_7445,N_5556);
or U10036 (N_10036,N_6114,N_6478);
nor U10037 (N_10037,N_9856,N_6241);
nor U10038 (N_10038,N_8539,N_6973);
nor U10039 (N_10039,N_5455,N_6795);
and U10040 (N_10040,N_7016,N_7860);
nand U10041 (N_10041,N_5632,N_9592);
nand U10042 (N_10042,N_8794,N_9079);
nor U10043 (N_10043,N_9998,N_8749);
or U10044 (N_10044,N_8312,N_7283);
nor U10045 (N_10045,N_8933,N_8023);
and U10046 (N_10046,N_7449,N_6534);
or U10047 (N_10047,N_6658,N_5958);
and U10048 (N_10048,N_6090,N_5249);
or U10049 (N_10049,N_7496,N_8561);
nand U10050 (N_10050,N_7444,N_7701);
and U10051 (N_10051,N_5741,N_9806);
nand U10052 (N_10052,N_7110,N_5237);
and U10053 (N_10053,N_5122,N_8847);
and U10054 (N_10054,N_6011,N_8591);
nor U10055 (N_10055,N_8251,N_7281);
and U10056 (N_10056,N_9917,N_6751);
or U10057 (N_10057,N_9547,N_8596);
nand U10058 (N_10058,N_5800,N_5603);
and U10059 (N_10059,N_9720,N_7011);
nand U10060 (N_10060,N_6126,N_8027);
nor U10061 (N_10061,N_7493,N_9694);
or U10062 (N_10062,N_8293,N_9319);
or U10063 (N_10063,N_8717,N_6978);
nor U10064 (N_10064,N_9907,N_7778);
or U10065 (N_10065,N_8086,N_8508);
nand U10066 (N_10066,N_7656,N_7198);
nand U10067 (N_10067,N_6158,N_5796);
or U10068 (N_10068,N_5270,N_9380);
or U10069 (N_10069,N_6063,N_7555);
nand U10070 (N_10070,N_9016,N_6618);
nor U10071 (N_10071,N_6284,N_7976);
nand U10072 (N_10072,N_6036,N_6489);
and U10073 (N_10073,N_7374,N_9656);
nand U10074 (N_10074,N_5115,N_5678);
nor U10075 (N_10075,N_7763,N_9800);
nand U10076 (N_10076,N_9073,N_6287);
nor U10077 (N_10077,N_8343,N_5960);
nand U10078 (N_10078,N_9054,N_6359);
nor U10079 (N_10079,N_6373,N_9673);
and U10080 (N_10080,N_7983,N_5261);
nor U10081 (N_10081,N_5119,N_7648);
nand U10082 (N_10082,N_5204,N_6049);
or U10083 (N_10083,N_9453,N_9691);
or U10084 (N_10084,N_5505,N_5133);
nor U10085 (N_10085,N_5441,N_6021);
nand U10086 (N_10086,N_6444,N_7012);
nor U10087 (N_10087,N_5416,N_8030);
nor U10088 (N_10088,N_6463,N_5456);
nor U10089 (N_10089,N_5397,N_9870);
and U10090 (N_10090,N_9290,N_7719);
nand U10091 (N_10091,N_8684,N_8746);
or U10092 (N_10092,N_5266,N_6428);
and U10093 (N_10093,N_5512,N_8034);
nand U10094 (N_10094,N_9298,N_6593);
and U10095 (N_10095,N_6807,N_6647);
nor U10096 (N_10096,N_5054,N_6175);
and U10097 (N_10097,N_8434,N_9139);
and U10098 (N_10098,N_6977,N_7459);
nand U10099 (N_10099,N_6668,N_9063);
nand U10100 (N_10100,N_9764,N_8164);
nor U10101 (N_10101,N_8545,N_9881);
nand U10102 (N_10102,N_7050,N_9864);
and U10103 (N_10103,N_9920,N_6667);
or U10104 (N_10104,N_8321,N_8965);
and U10105 (N_10105,N_7175,N_6828);
nand U10106 (N_10106,N_8189,N_8056);
nor U10107 (N_10107,N_7148,N_7364);
nand U10108 (N_10108,N_6402,N_9065);
nand U10109 (N_10109,N_8697,N_9299);
nand U10110 (N_10110,N_7083,N_9495);
and U10111 (N_10111,N_7940,N_8142);
and U10112 (N_10112,N_7252,N_8808);
nor U10113 (N_10113,N_5689,N_6565);
nor U10114 (N_10114,N_6709,N_9947);
nand U10115 (N_10115,N_6414,N_5079);
and U10116 (N_10116,N_9215,N_8777);
or U10117 (N_10117,N_8390,N_6080);
and U10118 (N_10118,N_5475,N_9423);
or U10119 (N_10119,N_9786,N_5969);
nor U10120 (N_10120,N_7726,N_6198);
and U10121 (N_10121,N_6336,N_5268);
and U10122 (N_10122,N_8152,N_7655);
and U10123 (N_10123,N_9831,N_6420);
nand U10124 (N_10124,N_5345,N_6281);
and U10125 (N_10125,N_9991,N_7208);
or U10126 (N_10126,N_6216,N_6050);
nand U10127 (N_10127,N_8642,N_8000);
xor U10128 (N_10128,N_8995,N_8076);
or U10129 (N_10129,N_7897,N_6048);
or U10130 (N_10130,N_9436,N_8671);
nand U10131 (N_10131,N_5061,N_9373);
nor U10132 (N_10132,N_5434,N_9040);
nor U10133 (N_10133,N_6136,N_6413);
nor U10134 (N_10134,N_9899,N_9327);
or U10135 (N_10135,N_8410,N_9179);
nand U10136 (N_10136,N_7008,N_7560);
nor U10137 (N_10137,N_7948,N_8734);
or U10138 (N_10138,N_8331,N_7332);
or U10139 (N_10139,N_5067,N_7028);
nor U10140 (N_10140,N_5923,N_9150);
nand U10141 (N_10141,N_7325,N_9284);
and U10142 (N_10142,N_5229,N_9377);
or U10143 (N_10143,N_8703,N_9702);
nand U10144 (N_10144,N_7000,N_7779);
nand U10145 (N_10145,N_6217,N_6713);
and U10146 (N_10146,N_7287,N_5503);
nor U10147 (N_10147,N_9768,N_6346);
or U10148 (N_10148,N_7640,N_5953);
and U10149 (N_10149,N_5672,N_7305);
and U10150 (N_10150,N_8552,N_9445);
or U10151 (N_10151,N_8557,N_6151);
nand U10152 (N_10152,N_8565,N_8976);
and U10153 (N_10153,N_5590,N_8594);
nor U10154 (N_10154,N_8687,N_9523);
and U10155 (N_10155,N_9894,N_7740);
nand U10156 (N_10156,N_7461,N_9585);
and U10157 (N_10157,N_5636,N_6105);
and U10158 (N_10158,N_9697,N_9482);
and U10159 (N_10159,N_9905,N_5784);
and U10160 (N_10160,N_7264,N_7761);
nor U10161 (N_10161,N_8036,N_5722);
nor U10162 (N_10162,N_5879,N_8427);
nor U10163 (N_10163,N_7334,N_8806);
or U10164 (N_10164,N_9337,N_9071);
nand U10165 (N_10165,N_8825,N_9326);
nor U10166 (N_10166,N_6799,N_8253);
and U10167 (N_10167,N_9343,N_9074);
or U10168 (N_10168,N_9061,N_9834);
or U10169 (N_10169,N_5491,N_6846);
and U10170 (N_10170,N_7253,N_8722);
or U10171 (N_10171,N_9993,N_6741);
nor U10172 (N_10172,N_6317,N_7724);
or U10173 (N_10173,N_6590,N_6748);
or U10174 (N_10174,N_8582,N_9243);
nor U10175 (N_10175,N_7200,N_9840);
nor U10176 (N_10176,N_6675,N_7801);
or U10177 (N_10177,N_8329,N_8209);
nor U10178 (N_10178,N_5078,N_5364);
nor U10179 (N_10179,N_6429,N_7616);
and U10180 (N_10180,N_7346,N_6333);
nor U10181 (N_10181,N_9629,N_8573);
nand U10182 (N_10182,N_5607,N_6689);
xor U10183 (N_10183,N_9518,N_8327);
nand U10184 (N_10184,N_6766,N_5690);
nand U10185 (N_10185,N_5778,N_8021);
or U10186 (N_10186,N_7780,N_9900);
nor U10187 (N_10187,N_9526,N_8644);
nand U10188 (N_10188,N_7438,N_5549);
and U10189 (N_10189,N_6327,N_8396);
nor U10190 (N_10190,N_8219,N_8357);
or U10191 (N_10191,N_9604,N_6531);
and U10192 (N_10192,N_8917,N_8063);
and U10193 (N_10193,N_6696,N_6314);
and U10194 (N_10194,N_9506,N_6172);
nor U10195 (N_10195,N_6882,N_7034);
and U10196 (N_10196,N_8504,N_7864);
and U10197 (N_10197,N_6500,N_6165);
nor U10198 (N_10198,N_5637,N_8769);
nor U10199 (N_10199,N_7803,N_6178);
nand U10200 (N_10200,N_7085,N_5164);
or U10201 (N_10201,N_7368,N_6487);
or U10202 (N_10202,N_6409,N_8580);
nand U10203 (N_10203,N_5527,N_7971);
nand U10204 (N_10204,N_5428,N_7970);
or U10205 (N_10205,N_8955,N_5329);
xor U10206 (N_10206,N_8991,N_8583);
nand U10207 (N_10207,N_9739,N_8320);
or U10208 (N_10208,N_5410,N_8185);
and U10209 (N_10209,N_5658,N_5446);
and U10210 (N_10210,N_9589,N_5276);
and U10211 (N_10211,N_5724,N_8347);
nand U10212 (N_10212,N_6291,N_7105);
nor U10213 (N_10213,N_9573,N_9594);
and U10214 (N_10214,N_9317,N_6037);
and U10215 (N_10215,N_6827,N_5826);
or U10216 (N_10216,N_7394,N_9501);
nor U10217 (N_10217,N_6497,N_9636);
nor U10218 (N_10218,N_6499,N_9166);
and U10219 (N_10219,N_6613,N_6555);
and U10220 (N_10220,N_7172,N_6580);
nor U10221 (N_10221,N_7313,N_7343);
or U10222 (N_10222,N_9486,N_6095);
nor U10223 (N_10223,N_7858,N_8790);
nor U10224 (N_10224,N_5400,N_8083);
nor U10225 (N_10225,N_5443,N_6093);
nor U10226 (N_10226,N_8130,N_5281);
nand U10227 (N_10227,N_6953,N_6442);
nor U10228 (N_10228,N_6356,N_9729);
or U10229 (N_10229,N_8656,N_6893);
or U10230 (N_10230,N_7066,N_5931);
and U10231 (N_10231,N_9378,N_9037);
and U10232 (N_10232,N_6466,N_8826);
nor U10233 (N_10233,N_8052,N_5783);
or U10234 (N_10234,N_6342,N_9680);
nand U10235 (N_10235,N_8387,N_7073);
or U10236 (N_10236,N_7553,N_5866);
nand U10237 (N_10237,N_7595,N_6598);
nor U10238 (N_10238,N_9607,N_7571);
or U10239 (N_10239,N_8278,N_9280);
nand U10240 (N_10240,N_5474,N_6374);
nand U10241 (N_10241,N_6260,N_7227);
xor U10242 (N_10242,N_7809,N_5538);
and U10243 (N_10243,N_7472,N_7525);
nand U10244 (N_10244,N_6459,N_5814);
and U10245 (N_10245,N_7142,N_9827);
or U10246 (N_10246,N_5408,N_7917);
and U10247 (N_10247,N_5612,N_9468);
and U10248 (N_10248,N_8055,N_8727);
nand U10249 (N_10249,N_7484,N_6184);
nor U10250 (N_10250,N_6157,N_5401);
and U10251 (N_10251,N_9678,N_8148);
and U10252 (N_10252,N_9599,N_7882);
nor U10253 (N_10253,N_5886,N_7950);
nand U10254 (N_10254,N_7228,N_9018);
nor U10255 (N_10255,N_6723,N_8066);
nand U10256 (N_10256,N_6012,N_7625);
or U10257 (N_10257,N_9304,N_9564);
and U10258 (N_10258,N_7627,N_7181);
and U10259 (N_10259,N_8166,N_8970);
nand U10260 (N_10260,N_6909,N_7323);
nand U10261 (N_10261,N_7787,N_6889);
nor U10262 (N_10262,N_8861,N_8953);
nand U10263 (N_10263,N_9101,N_8881);
nor U10264 (N_10264,N_7117,N_5846);
nor U10265 (N_10265,N_5736,N_8273);
nand U10266 (N_10266,N_9248,N_8054);
nand U10267 (N_10267,N_8696,N_6694);
or U10268 (N_10268,N_7482,N_5222);
nor U10269 (N_10269,N_8087,N_5933);
nor U10270 (N_10270,N_5992,N_6480);
or U10271 (N_10271,N_6207,N_8537);
and U10272 (N_10272,N_7794,N_7517);
nand U10273 (N_10273,N_6641,N_5699);
nor U10274 (N_10274,N_8866,N_9241);
and U10275 (N_10275,N_7468,N_8605);
or U10276 (N_10276,N_7250,N_9091);
nand U10277 (N_10277,N_5496,N_8971);
or U10278 (N_10278,N_7573,N_6671);
or U10279 (N_10279,N_5982,N_5669);
and U10280 (N_10280,N_6627,N_9854);
nand U10281 (N_10281,N_6308,N_9408);
and U10282 (N_10282,N_9809,N_7382);
nor U10283 (N_10283,N_9398,N_5595);
nand U10284 (N_10284,N_5665,N_8632);
or U10285 (N_10285,N_8856,N_5565);
or U10286 (N_10286,N_6566,N_9562);
and U10287 (N_10287,N_8042,N_7254);
nor U10288 (N_10288,N_5748,N_5890);
nor U10289 (N_10289,N_9543,N_6229);
nor U10290 (N_10290,N_6133,N_7164);
and U10291 (N_10291,N_6919,N_8242);
nand U10292 (N_10292,N_8781,N_8613);
nor U10293 (N_10293,N_9229,N_6300);
nor U10294 (N_10294,N_6920,N_9999);
nand U10295 (N_10295,N_9612,N_5551);
and U10296 (N_10296,N_7895,N_6181);
nand U10297 (N_10297,N_9131,N_5899);
and U10298 (N_10298,N_7353,N_9448);
or U10299 (N_10299,N_6993,N_5076);
nor U10300 (N_10300,N_5362,N_6437);
and U10301 (N_10301,N_5872,N_5116);
nor U10302 (N_10302,N_9875,N_7590);
or U10303 (N_10303,N_8416,N_7078);
and U10304 (N_10304,N_6944,N_6326);
or U10305 (N_10305,N_9638,N_8570);
nand U10306 (N_10306,N_7973,N_8014);
nor U10307 (N_10307,N_5490,N_5207);
nand U10308 (N_10308,N_8236,N_9624);
or U10309 (N_10309,N_8425,N_9007);
and U10310 (N_10310,N_6191,N_7077);
or U10311 (N_10311,N_5578,N_6180);
and U10312 (N_10312,N_7686,N_7104);
and U10313 (N_10313,N_6623,N_9630);
nor U10314 (N_10314,N_5454,N_5521);
and U10315 (N_10315,N_5467,N_8721);
nor U10316 (N_10316,N_6502,N_6631);
and U10317 (N_10317,N_7567,N_8045);
nand U10318 (N_10318,N_9820,N_7225);
or U10319 (N_10319,N_6726,N_8901);
and U10320 (N_10320,N_9842,N_6802);
nand U10321 (N_10321,N_8767,N_5308);
and U10322 (N_10322,N_7197,N_7354);
or U10323 (N_10323,N_6083,N_8071);
nor U10324 (N_10324,N_9645,N_8474);
xor U10325 (N_10325,N_6412,N_9663);
and U10326 (N_10326,N_9272,N_8514);
nand U10327 (N_10327,N_7990,N_7939);
nor U10328 (N_10328,N_7876,N_5398);
nand U10329 (N_10329,N_9681,N_5372);
nor U10330 (N_10330,N_6949,N_5387);
nand U10331 (N_10331,N_6441,N_5173);
and U10332 (N_10332,N_7916,N_6957);
nand U10333 (N_10333,N_7725,N_9413);
nor U10334 (N_10334,N_7727,N_9296);
and U10335 (N_10335,N_6861,N_6350);
and U10336 (N_10336,N_7692,N_8817);
nand U10337 (N_10337,N_6800,N_6013);
or U10338 (N_10338,N_6842,N_5997);
and U10339 (N_10339,N_8547,N_5623);
or U10340 (N_10340,N_9888,N_6529);
or U10341 (N_10341,N_5782,N_7423);
or U10342 (N_10342,N_6901,N_6553);
or U10343 (N_10343,N_8915,N_7434);
and U10344 (N_10344,N_5192,N_9741);
nor U10345 (N_10345,N_8070,N_7498);
and U10346 (N_10346,N_7160,N_6038);
and U10347 (N_10347,N_6742,N_9473);
and U10348 (N_10348,N_5912,N_9066);
or U10349 (N_10349,N_8883,N_6626);
nor U10350 (N_10350,N_6319,N_8344);
or U10351 (N_10351,N_6640,N_8483);
nor U10352 (N_10352,N_6869,N_8485);
nand U10353 (N_10353,N_8840,N_9618);
nor U10354 (N_10354,N_6269,N_5332);
and U10355 (N_10355,N_9355,N_7552);
or U10356 (N_10356,N_9839,N_8046);
nand U10357 (N_10357,N_8490,N_9051);
nand U10358 (N_10358,N_9356,N_7827);
nor U10359 (N_10359,N_9346,N_6206);
nand U10360 (N_10360,N_7024,N_6155);
nor U10361 (N_10361,N_9959,N_6174);
and U10362 (N_10362,N_8049,N_9511);
nor U10363 (N_10363,N_8082,N_6111);
or U10364 (N_10364,N_9259,N_6575);
or U10365 (N_10365,N_5419,N_9950);
xnor U10366 (N_10366,N_9135,N_8157);
nor U10367 (N_10367,N_7068,N_5127);
or U10368 (N_10368,N_5913,N_5284);
nor U10369 (N_10369,N_5803,N_9514);
nor U10370 (N_10370,N_5489,N_7019);
nand U10371 (N_10371,N_7129,N_9001);
nand U10372 (N_10372,N_8454,N_7989);
or U10373 (N_10373,N_6516,N_5943);
nand U10374 (N_10374,N_8489,N_7237);
nand U10375 (N_10375,N_7633,N_9194);
nor U10376 (N_10376,N_8618,N_6098);
nor U10377 (N_10377,N_7923,N_6801);
or U10378 (N_10378,N_9985,N_6458);
nor U10379 (N_10379,N_9893,N_9421);
nor U10380 (N_10380,N_9620,N_5003);
nand U10381 (N_10381,N_9790,N_9434);
and U10382 (N_10382,N_9360,N_7802);
and U10383 (N_10383,N_6072,N_5666);
nand U10384 (N_10384,N_9954,N_6772);
or U10385 (N_10385,N_8854,N_6141);
and U10386 (N_10386,N_7792,N_5154);
and U10387 (N_10387,N_9347,N_8180);
nand U10388 (N_10388,N_7178,N_9619);
nor U10389 (N_10389,N_9351,N_9158);
nor U10390 (N_10390,N_8162,N_6940);
and U10391 (N_10391,N_7097,N_5841);
nor U10392 (N_10392,N_8394,N_6628);
nor U10393 (N_10393,N_8424,N_8563);
nand U10394 (N_10394,N_8879,N_8754);
or U10395 (N_10395,N_6129,N_8633);
nand U10396 (N_10396,N_8735,N_6789);
nand U10397 (N_10397,N_7072,N_6797);
nor U10398 (N_10398,N_5064,N_8779);
nand U10399 (N_10399,N_9742,N_5624);
or U10400 (N_10400,N_8386,N_8984);
nor U10401 (N_10401,N_5497,N_5334);
nor U10402 (N_10402,N_8692,N_6596);
nand U10403 (N_10403,N_8374,N_9325);
nor U10404 (N_10404,N_5194,N_8527);
nand U10405 (N_10405,N_5654,N_5646);
and U10406 (N_10406,N_7777,N_8851);
nor U10407 (N_10407,N_7308,N_7871);
nor U10408 (N_10408,N_9212,N_7036);
nand U10409 (N_10409,N_9075,N_6798);
and U10410 (N_10410,N_8952,N_9916);
xor U10411 (N_10411,N_7413,N_9435);
and U10412 (N_10412,N_9237,N_6339);
and U10413 (N_10413,N_6952,N_6716);
nand U10414 (N_10414,N_7338,N_7589);
nand U10415 (N_10415,N_9148,N_9712);
and U10416 (N_10416,N_6731,N_7400);
or U10417 (N_10417,N_9713,N_6422);
or U10418 (N_10418,N_9804,N_8597);
and U10419 (N_10419,N_7123,N_5576);
and U10420 (N_10420,N_5391,N_6110);
nor U10421 (N_10421,N_5533,N_8511);
or U10422 (N_10422,N_6750,N_7872);
nand U10423 (N_10423,N_6512,N_5326);
nand U10424 (N_10424,N_5162,N_5071);
and U10425 (N_10425,N_5949,N_8100);
nand U10426 (N_10426,N_6041,N_9121);
nor U10427 (N_10427,N_7037,N_5716);
xnor U10428 (N_10428,N_7435,N_6721);
and U10429 (N_10429,N_8176,N_5965);
nand U10430 (N_10430,N_8402,N_9682);
and U10431 (N_10431,N_6922,N_5101);
nor U10432 (N_10432,N_6539,N_8616);
or U10433 (N_10433,N_7372,N_9973);
nand U10434 (N_10434,N_6476,N_6138);
nand U10435 (N_10435,N_9952,N_8430);
nor U10436 (N_10436,N_7894,N_9086);
or U10437 (N_10437,N_8859,N_9609);
nand U10438 (N_10438,N_6929,N_5640);
nor U10439 (N_10439,N_5794,N_9927);
nand U10440 (N_10440,N_9847,N_9208);
nor U10441 (N_10441,N_8713,N_8447);
nand U10442 (N_10442,N_5375,N_8448);
nor U10443 (N_10443,N_8235,N_9891);
and U10444 (N_10444,N_9862,N_9857);
or U10445 (N_10445,N_7879,N_9275);
or U10446 (N_10446,N_5018,N_6906);
nand U10447 (N_10447,N_9019,N_6074);
nand U10448 (N_10448,N_6006,N_6246);
nand U10449 (N_10449,N_9532,N_7706);
or U10450 (N_10450,N_5682,N_6734);
or U10451 (N_10451,N_9418,N_7328);
nor U10452 (N_10452,N_9402,N_5815);
and U10453 (N_10453,N_5053,N_6975);
xor U10454 (N_10454,N_9605,N_5539);
nand U10455 (N_10455,N_8449,N_8232);
nor U10456 (N_10456,N_8928,N_6880);
or U10457 (N_10457,N_6424,N_6431);
and U10458 (N_10458,N_6885,N_9851);
nand U10459 (N_10459,N_6468,N_6574);
or U10460 (N_10460,N_9535,N_6421);
nor U10461 (N_10461,N_8361,N_7494);
or U10462 (N_10462,N_9689,N_9155);
nor U10463 (N_10463,N_6786,N_7249);
and U10464 (N_10464,N_5753,N_7937);
or U10465 (N_10465,N_7152,N_7906);
nor U10466 (N_10466,N_6810,N_5163);
nor U10467 (N_10467,N_6283,N_5962);
or U10468 (N_10468,N_6112,N_6898);
nor U10469 (N_10469,N_8155,N_5377);
or U10470 (N_10470,N_9117,N_6197);
or U10471 (N_10471,N_5312,N_8069);
nor U10472 (N_10472,N_5580,N_9127);
or U10473 (N_10473,N_9880,N_6278);
nor U10474 (N_10474,N_9256,N_9582);
or U10475 (N_10475,N_7067,N_9330);
nand U10476 (N_10476,N_8184,N_9974);
nor U10477 (N_10477,N_7693,N_8478);
nor U10478 (N_10478,N_9525,N_6086);
and U10479 (N_10479,N_7262,N_5644);
nor U10480 (N_10480,N_8279,N_7756);
or U10481 (N_10481,N_9397,N_6209);
and U10482 (N_10482,N_7185,N_6062);
xnor U10483 (N_10483,N_6523,N_5887);
or U10484 (N_10484,N_8941,N_7600);
and U10485 (N_10485,N_8577,N_6301);
nor U10486 (N_10486,N_6616,N_5613);
nand U10487 (N_10487,N_8758,N_7677);
nor U10488 (N_10488,N_5609,N_5170);
nand U10489 (N_10489,N_9379,N_5863);
or U10490 (N_10490,N_6652,N_9843);
nand U10491 (N_10491,N_9928,N_9472);
and U10492 (N_10492,N_8875,N_8290);
and U10493 (N_10493,N_6070,N_5146);
or U10494 (N_10494,N_9271,N_7399);
nand U10495 (N_10495,N_7582,N_8649);
and U10496 (N_10496,N_8466,N_5599);
and U10497 (N_10497,N_9046,N_5444);
nand U10498 (N_10498,N_5494,N_9245);
or U10499 (N_10499,N_5729,N_6131);
and U10500 (N_10500,N_9895,N_8339);
nand U10501 (N_10501,N_7510,N_5031);
or U10502 (N_10502,N_8660,N_6720);
nand U10503 (N_10503,N_9538,N_6839);
or U10504 (N_10504,N_6552,N_9865);
nand U10505 (N_10505,N_5221,N_7173);
and U10506 (N_10506,N_8575,N_9137);
nor U10507 (N_10507,N_6573,N_5940);
and U10508 (N_10508,N_7862,N_8668);
nand U10509 (N_10509,N_8233,N_8007);
nor U10510 (N_10510,N_8224,N_9937);
nand U10511 (N_10511,N_8765,N_9964);
and U10512 (N_10512,N_6891,N_9855);
and U10513 (N_10513,N_7301,N_6335);
or U10514 (N_10514,N_5761,N_9489);
nand U10515 (N_10515,N_8324,N_6495);
or U10516 (N_10516,N_9517,N_9032);
and U10517 (N_10517,N_7551,N_8428);
nor U10518 (N_10518,N_9542,N_8927);
and U10519 (N_10519,N_7830,N_7465);
nand U10520 (N_10520,N_9755,N_5944);
nor U10521 (N_10521,N_9396,N_7757);
nor U10522 (N_10522,N_8751,N_6833);
and U10523 (N_10523,N_6817,N_7218);
and U10524 (N_10524,N_5016,N_7395);
and U10525 (N_10525,N_8657,N_9459);
and U10526 (N_10526,N_9698,N_5225);
nand U10527 (N_10527,N_9062,N_5571);
or U10528 (N_10528,N_8064,N_9332);
nor U10529 (N_10529,N_7532,N_9324);
or U10530 (N_10530,N_8337,N_7139);
nor U10531 (N_10531,N_6915,N_7277);
nand U10532 (N_10532,N_7256,N_7379);
and U10533 (N_10533,N_7404,N_6467);
nand U10534 (N_10534,N_9710,N_7076);
and U10535 (N_10535,N_7883,N_8715);
nor U10536 (N_10536,N_8538,N_9876);
nor U10537 (N_10537,N_6851,N_7107);
or U10538 (N_10538,N_8918,N_5577);
nand U10539 (N_10539,N_5530,N_8379);
and U10540 (N_10540,N_5504,N_5370);
or U10541 (N_10541,N_8043,N_6960);
or U10542 (N_10542,N_8020,N_6608);
and U10543 (N_10543,N_9601,N_9600);
nor U10544 (N_10544,N_6638,N_5862);
nand U10545 (N_10545,N_8296,N_7890);
nand U10546 (N_10546,N_8682,N_9737);
or U10547 (N_10547,N_5597,N_5136);
nor U10548 (N_10548,N_8028,N_9393);
or U10549 (N_10549,N_5365,N_7169);
and U10550 (N_10550,N_8691,N_7159);
nor U10551 (N_10551,N_7536,N_6781);
nor U10552 (N_10552,N_5302,N_7703);
nand U10553 (N_10553,N_7678,N_7966);
and U10554 (N_10554,N_6149,N_9926);
nand U10555 (N_10555,N_9613,N_8096);
and U10556 (N_10556,N_6395,N_5779);
or U10557 (N_10557,N_7905,N_5718);
and U10558 (N_10558,N_5210,N_6985);
or U10559 (N_10559,N_6739,N_6820);
nor U10560 (N_10560,N_8287,N_7003);
or U10561 (N_10561,N_6315,N_8892);
nand U10562 (N_10562,N_6597,N_5730);
and U10563 (N_10563,N_9759,N_9853);
and U10564 (N_10564,N_5432,N_5291);
nor U10565 (N_10565,N_6963,N_9817);
or U10566 (N_10566,N_9626,N_8516);
nand U10567 (N_10567,N_6094,N_5328);
nand U10568 (N_10568,N_5514,N_8791);
or U10569 (N_10569,N_7206,N_7810);
nand U10570 (N_10570,N_6875,N_5252);
or U10571 (N_10571,N_7322,N_6355);
nor U10572 (N_10572,N_9986,N_5128);
nor U10573 (N_10573,N_5859,N_5750);
and U10574 (N_10574,N_5706,N_6942);
nor U10575 (N_10575,N_9111,N_8358);
nor U10576 (N_10576,N_9218,N_6371);
nor U10577 (N_10577,N_5621,N_7695);
nand U10578 (N_10578,N_8823,N_5023);
nand U10579 (N_10579,N_6545,N_6989);
nor U10580 (N_10580,N_6967,N_9794);
or U10581 (N_10581,N_9210,N_6262);
nand U10582 (N_10582,N_5201,N_8903);
nand U10583 (N_10583,N_7199,N_9572);
and U10584 (N_10584,N_7203,N_5149);
and U10585 (N_10585,N_9652,N_5854);
nor U10586 (N_10586,N_5765,N_6456);
nand U10587 (N_10587,N_9979,N_5452);
and U10588 (N_10588,N_5787,N_5891);
or U10589 (N_10589,N_8486,N_7755);
and U10590 (N_10590,N_5795,N_5893);
nand U10591 (N_10591,N_6864,N_7086);
nor U10592 (N_10592,N_8771,N_6803);
or U10593 (N_10593,N_8852,N_9220);
or U10594 (N_10594,N_5555,N_9478);
or U10595 (N_10595,N_5684,N_6432);
and U10596 (N_10596,N_9848,N_6886);
or U10597 (N_10597,N_6763,N_7402);
nor U10598 (N_10598,N_9428,N_9584);
nand U10599 (N_10599,N_6712,N_5202);
nor U10600 (N_10600,N_6295,N_8263);
and U10601 (N_10601,N_6270,N_7483);
nor U10602 (N_10602,N_5126,N_5703);
nand U10603 (N_10603,N_9384,N_8377);
or U10604 (N_10604,N_5242,N_5143);
nor U10605 (N_10605,N_7653,N_6085);
or U10606 (N_10606,N_8281,N_8961);
or U10607 (N_10607,N_8481,N_8576);
nor U10608 (N_10608,N_6214,N_5289);
nor U10609 (N_10609,N_8409,N_7014);
or U10610 (N_10610,N_7770,N_7020);
nand U10611 (N_10611,N_7932,N_9409);
nor U10612 (N_10612,N_8149,N_6780);
or U10613 (N_10613,N_9530,N_7784);
nand U10614 (N_10614,N_7084,N_9684);
or U10615 (N_10615,N_6097,N_8981);
and U10616 (N_10616,N_5987,N_5449);
and U10617 (N_10617,N_7504,N_5711);
nor U10618 (N_10618,N_9112,N_7319);
and U10619 (N_10619,N_9971,N_9228);
nand U10620 (N_10620,N_8179,N_6693);
or U10621 (N_10621,N_7847,N_8151);
and U10622 (N_10622,N_8376,N_9628);
nand U10623 (N_10623,N_5822,N_8873);
nand U10624 (N_10624,N_6717,N_8496);
or U10625 (N_10625,N_6522,N_6657);
nor U10626 (N_10626,N_7969,N_6806);
nand U10627 (N_10627,N_9181,N_8679);
and U10628 (N_10628,N_8589,N_7128);
and U10629 (N_10629,N_7859,N_6888);
nand U10630 (N_10630,N_8009,N_5459);
nor U10631 (N_10631,N_8060,N_5853);
nand U10632 (N_10632,N_9836,N_7245);
nand U10633 (N_10633,N_7647,N_5820);
nor U10634 (N_10634,N_9749,N_8667);
or U10635 (N_10635,N_6256,N_5659);
nand U10636 (N_10636,N_6073,N_9427);
nor U10637 (N_10637,N_9060,N_6856);
nand U10638 (N_10638,N_5095,N_7835);
or U10639 (N_10639,N_5875,N_5050);
nand U10640 (N_10640,N_7065,N_7900);
nand U10641 (N_10641,N_8648,N_5137);
nand U10642 (N_10642,N_5305,N_7749);
nor U10643 (N_10643,N_8569,N_7315);
nand U10644 (N_10644,N_7424,N_7304);
nand U10645 (N_10645,N_7715,N_8476);
nor U10646 (N_10646,N_9200,N_7205);
and U10647 (N_10647,N_9057,N_7539);
nand U10648 (N_10648,N_8450,N_5028);
or U10649 (N_10649,N_6190,N_5077);
nor U10650 (N_10650,N_6835,N_6302);
or U10651 (N_10651,N_9183,N_5480);
and U10652 (N_10652,N_7191,N_8581);
nor U10653 (N_10653,N_9022,N_9216);
nor U10654 (N_10654,N_6449,N_5367);
nand U10655 (N_10655,N_9923,N_5907);
nor U10656 (N_10656,N_7153,N_7850);
and U10657 (N_10657,N_8702,N_6881);
or U10658 (N_10658,N_9161,N_9072);
nand U10659 (N_10659,N_5507,N_7018);
and U10660 (N_10660,N_8111,N_6303);
nand U10661 (N_10661,N_9637,N_9188);
and U10662 (N_10662,N_5870,N_5272);
nand U10663 (N_10663,N_7839,N_8322);
and U10664 (N_10664,N_5811,N_9247);
nand U10665 (N_10665,N_6790,N_9206);
or U10666 (N_10666,N_8784,N_6340);
or U10667 (N_10667,N_5215,N_7030);
nand U10668 (N_10668,N_8796,N_5336);
and U10669 (N_10669,N_7867,N_7233);
and U10670 (N_10670,N_8534,N_7230);
and U10671 (N_10671,N_9982,N_8471);
or U10672 (N_10672,N_7661,N_7061);
and U10673 (N_10673,N_5132,N_6821);
nor U10674 (N_10674,N_7592,N_9949);
nand U10675 (N_10675,N_6369,N_5671);
nand U10676 (N_10676,N_7586,N_8182);
nand U10677 (N_10677,N_7981,N_7509);
and U10678 (N_10678,N_5777,N_6177);
nor U10679 (N_10679,N_9816,N_6841);
or U10680 (N_10680,N_5418,N_9765);
or U10681 (N_10681,N_6677,N_7035);
and U10682 (N_10682,N_5957,N_7806);
or U10683 (N_10683,N_8652,N_9874);
and U10684 (N_10684,N_5112,N_6550);
nand U10685 (N_10685,N_5180,N_7909);
or U10686 (N_10686,N_8128,N_7610);
and U10687 (N_10687,N_7217,N_9548);
or U10688 (N_10688,N_9357,N_8564);
or U10689 (N_10689,N_8920,N_6676);
or U10690 (N_10690,N_8025,N_5829);
and U10691 (N_10691,N_8559,N_8908);
nand U10692 (N_10692,N_8493,N_7156);
nand U10693 (N_10693,N_8211,N_5986);
and U10694 (N_10694,N_9463,N_6725);
nand U10695 (N_10695,N_5948,N_7219);
nor U10696 (N_10696,N_8498,N_5697);
or U10697 (N_10697,N_8065,N_6792);
and U10698 (N_10698,N_6189,N_6615);
or U10699 (N_10699,N_5083,N_7721);
nor U10700 (N_10700,N_5234,N_9995);
and U10701 (N_10701,N_7711,N_7158);
nand U10702 (N_10702,N_7431,N_6629);
or U10703 (N_10703,N_8845,N_5752);
and U10704 (N_10704,N_6609,N_5745);
or U10705 (N_10705,N_7309,N_8408);
or U10706 (N_10706,N_8203,N_7464);
and U10707 (N_10707,N_8282,N_7095);
or U10708 (N_10708,N_9105,N_9368);
nand U10709 (N_10709,N_9283,N_9897);
nor U10710 (N_10710,N_9587,N_7489);
nor U10711 (N_10711,N_7682,N_7594);
nor U10712 (N_10712,N_7507,N_6765);
nand U10713 (N_10713,N_5518,N_5939);
nor U10714 (N_10714,N_8824,N_7347);
and U10715 (N_10715,N_8531,N_9294);
and U10716 (N_10716,N_8850,N_8896);
nand U10717 (N_10717,N_9039,N_7618);
or U10718 (N_10718,N_6863,N_7884);
nand U10719 (N_10719,N_9883,N_8120);
nor U10720 (N_10720,N_5936,N_5488);
and U10721 (N_10721,N_7064,N_9056);
or U10722 (N_10722,N_7240,N_5402);
nand U10723 (N_10723,N_9735,N_6101);
nand U10724 (N_10724,N_8705,N_6498);
or U10725 (N_10725,N_7813,N_9863);
nor U10726 (N_10726,N_5486,N_8990);
nand U10727 (N_10727,N_6986,N_5984);
or U10728 (N_10728,N_9458,N_6425);
and U10729 (N_10729,N_8340,N_9038);
nor U10730 (N_10730,N_7135,N_8246);
nor U10731 (N_10731,N_5568,N_7348);
or U10732 (N_10732,N_8002,N_8541);
nor U10733 (N_10733,N_5042,N_9746);
nor U10734 (N_10734,N_8144,N_6847);
nand U10735 (N_10735,N_5134,N_8601);
and U10736 (N_10736,N_9388,N_8031);
or U10737 (N_10737,N_5069,N_6299);
nand U10738 (N_10738,N_9824,N_9996);
and U10739 (N_10739,N_9945,N_9590);
or U10740 (N_10740,N_5789,N_5950);
nand U10741 (N_10741,N_7396,N_7383);
and U10742 (N_10742,N_6645,N_6937);
and U10743 (N_10743,N_8923,N_8080);
nor U10744 (N_10744,N_6289,N_7487);
nor U10745 (N_10745,N_8205,N_9719);
or U10746 (N_10746,N_5563,N_6415);
xor U10747 (N_10747,N_6313,N_8925);
and U10748 (N_10748,N_8533,N_7956);
or U10749 (N_10749,N_5685,N_9009);
and U10750 (N_10750,N_5661,N_5323);
or U10751 (N_10751,N_6508,N_9264);
nor U10752 (N_10752,N_5065,N_6664);
nor U10753 (N_10753,N_6125,N_5587);
nor U10754 (N_10754,N_7566,N_6887);
or U10755 (N_10755,N_8145,N_7490);
nand U10756 (N_10756,N_6018,N_9481);
or U10757 (N_10757,N_5901,N_8899);
and U10758 (N_10758,N_5819,N_8115);
nor U10759 (N_10759,N_5605,N_9551);
or U10760 (N_10760,N_5306,N_6426);
or U10761 (N_10761,N_9257,N_6030);
nand U10762 (N_10762,N_5584,N_8773);
nor U10763 (N_10763,N_5797,N_6680);
or U10764 (N_10764,N_6124,N_8535);
nor U10765 (N_10765,N_7485,N_9083);
and U10766 (N_10766,N_8733,N_6193);
and U10767 (N_10767,N_9479,N_7783);
or U10768 (N_10768,N_9106,N_6710);
or U10769 (N_10769,N_5517,N_6948);
or U10770 (N_10770,N_7634,N_7229);
or U10771 (N_10771,N_9981,N_6927);
nand U10772 (N_10772,N_7843,N_7972);
nor U10773 (N_10773,N_6082,N_6932);
and U10774 (N_10774,N_8105,N_8383);
or U10775 (N_10775,N_6047,N_9316);
or U10776 (N_10776,N_9361,N_8957);
nor U10777 (N_10777,N_7557,N_6683);
and U10778 (N_10778,N_8094,N_8467);
nand U10779 (N_10779,N_7141,N_7767);
and U10780 (N_10780,N_9339,N_7888);
or U10781 (N_10781,N_8740,N_6752);
or U10782 (N_10782,N_7978,N_5498);
nor U10783 (N_10783,N_5288,N_9596);
nand U10784 (N_10784,N_6264,N_7474);
nor U10785 (N_10785,N_9724,N_8106);
nor U10786 (N_10786,N_8124,N_6106);
nand U10787 (N_10787,N_7165,N_7886);
nor U10788 (N_10788,N_7432,N_8676);
and U10789 (N_10789,N_6410,N_5865);
and U10790 (N_10790,N_7025,N_6148);
and U10791 (N_10791,N_5849,N_8770);
nor U10792 (N_10792,N_9606,N_8878);
or U10793 (N_10793,N_9340,N_7699);
nor U10794 (N_10794,N_6509,N_5049);
nand U10795 (N_10795,N_5254,N_6775);
or U10796 (N_10796,N_8451,N_7901);
and U10797 (N_10797,N_7933,N_7665);
and U10798 (N_10798,N_7521,N_9990);
or U10799 (N_10799,N_5232,N_5297);
or U10800 (N_10800,N_6393,N_6228);
and U10801 (N_10801,N_6736,N_6559);
and U10802 (N_10802,N_7747,N_6194);
or U10803 (N_10803,N_8710,N_9159);
nand U10804 (N_10804,N_6427,N_7453);
nor U10805 (N_10805,N_6610,N_8143);
or U10806 (N_10806,N_9254,N_7938);
and U10807 (N_10807,N_8664,N_7397);
and U10808 (N_10808,N_8627,N_7672);
nor U10809 (N_10809,N_7033,N_6630);
and U10810 (N_10810,N_8391,N_9726);
nand U10811 (N_10811,N_7955,N_6530);
nor U10812 (N_10812,N_7144,N_6016);
or U10813 (N_10813,N_7753,N_9013);
or U10814 (N_10814,N_7898,N_6104);
and U10815 (N_10815,N_7327,N_8980);
and U10816 (N_10816,N_6777,N_8686);
nor U10817 (N_10817,N_5970,N_5102);
nor U10818 (N_10818,N_9447,N_9392);
nor U10819 (N_10819,N_6183,N_5604);
nor U10820 (N_10820,N_6014,N_8218);
nor U10821 (N_10821,N_8004,N_5309);
nor U10822 (N_10822,N_6998,N_9329);
nor U10823 (N_10823,N_5015,N_5619);
or U10824 (N_10824,N_9287,N_6389);
nand U10825 (N_10825,N_9805,N_8507);
and U10826 (N_10826,N_8936,N_6473);
nand U10827 (N_10827,N_6089,N_5544);
and U10828 (N_10828,N_9913,N_7093);
nand U10829 (N_10829,N_5909,N_9002);
or U10830 (N_10830,N_8704,N_6791);
nand U10831 (N_10831,N_7223,N_9925);
and U10832 (N_10832,N_7982,N_9136);
nand U10833 (N_10833,N_7577,N_7411);
and U10834 (N_10834,N_9829,N_7190);
or U10835 (N_10835,N_6446,N_5734);
nand U10836 (N_10836,N_7949,N_9502);
and U10837 (N_10837,N_5998,N_9268);
nor U10838 (N_10838,N_9429,N_5399);
nand U10839 (N_10839,N_8138,N_5156);
nor U10840 (N_10840,N_8468,N_7365);
or U10841 (N_10841,N_7881,N_9911);
nand U10842 (N_10842,N_8587,N_8436);
and U10843 (N_10843,N_9491,N_5200);
or U10844 (N_10844,N_7143,N_5085);
or U10845 (N_10845,N_9695,N_6385);
and U10846 (N_10846,N_5409,N_7335);
nor U10847 (N_10847,N_6687,N_7188);
nand U10848 (N_10848,N_8472,N_8744);
nor U10849 (N_10849,N_6026,N_6558);
nand U10850 (N_10850,N_8258,N_9114);
or U10851 (N_10851,N_8153,N_8283);
or U10852 (N_10852,N_9410,N_7392);
xnor U10853 (N_10853,N_9603,N_9004);
and U10854 (N_10854,N_7915,N_6377);
and U10855 (N_10855,N_5562,N_7518);
and U10856 (N_10856,N_6587,N_9942);
nand U10857 (N_10857,N_5066,N_9627);
nand U10858 (N_10858,N_8762,N_5993);
nor U10859 (N_10859,N_8316,N_8013);
and U10860 (N_10860,N_5072,N_8567);
nor U10861 (N_10861,N_7739,N_9909);
or U10862 (N_10862,N_6535,N_7788);
and U10863 (N_10863,N_5322,N_9519);
or U10864 (N_10864,N_5760,N_6688);
nor U10865 (N_10865,N_8311,N_6572);
or U10866 (N_10866,N_9617,N_7426);
and U10867 (N_10867,N_7032,N_6220);
nand U10868 (N_10868,N_7892,N_9581);
nor U10869 (N_10869,N_9866,N_7202);
or U10870 (N_10870,N_9664,N_5702);
nand U10871 (N_10871,N_7090,N_8241);
and U10872 (N_10872,N_5626,N_5648);
and U10873 (N_10873,N_8973,N_7583);
nor U10874 (N_10874,N_6347,N_8701);
and U10875 (N_10875,N_8837,N_9010);
nor U10876 (N_10876,N_6621,N_5838);
and U10877 (N_10877,N_6154,N_5611);
and U10878 (N_10878,N_8598,N_8792);
nor U10879 (N_10879,N_9559,N_8730);
and U10880 (N_10880,N_8921,N_6053);
nand U10881 (N_10881,N_8006,N_6707);
nor U10882 (N_10882,N_9640,N_9232);
or U10883 (N_10883,N_9785,N_7776);
nand U10884 (N_10884,N_7869,N_9116);
or U10885 (N_10885,N_5421,N_9467);
and U10886 (N_10886,N_9430,N_8050);
or U10887 (N_10887,N_5959,N_5830);
nand U10888 (N_10888,N_7605,N_7151);
or U10889 (N_10889,N_5868,N_8939);
nand U10890 (N_10890,N_9772,N_5740);
or U10891 (N_10891,N_9286,N_6577);
nand U10892 (N_10892,N_9747,N_9014);
nor U10893 (N_10893,N_9797,N_6980);
nand U10894 (N_10894,N_8810,N_6481);
or U10895 (N_10895,N_6589,N_9823);
nor U10896 (N_10896,N_5278,N_7515);
and U10897 (N_10897,N_9322,N_8256);
nand U10898 (N_10898,N_6533,N_6100);
or U10899 (N_10899,N_6028,N_9674);
nand U10900 (N_10900,N_7519,N_9302);
nand U10901 (N_10901,N_8439,N_9441);
or U10902 (N_10902,N_9359,N_8766);
or U10903 (N_10903,N_7132,N_7707);
nor U10904 (N_10904,N_5223,N_7537);
or U10905 (N_10905,N_8723,N_8348);
nand U10906 (N_10906,N_7224,N_5196);
or U10907 (N_10907,N_9718,N_5352);
or U10908 (N_10908,N_5141,N_7578);
and U10909 (N_10909,N_7638,N_8058);
nand U10910 (N_10910,N_6754,N_9269);
nand U10911 (N_10911,N_6691,N_8227);
or U10912 (N_10912,N_5564,N_7119);
and U10913 (N_10913,N_6474,N_7422);
and U10914 (N_10914,N_8994,N_9503);
nor U10915 (N_10915,N_5248,N_5792);
nor U10916 (N_10916,N_8836,N_6984);
nor U10917 (N_10917,N_7381,N_7221);
and U10918 (N_10918,N_7622,N_8663);
nor U10919 (N_10919,N_5415,N_6365);
nor U10920 (N_10920,N_7918,N_5653);
and U10921 (N_10921,N_7133,N_9717);
and U10922 (N_10922,N_5989,N_7951);
nor U10923 (N_10923,N_5005,N_6245);
nand U10924 (N_10924,N_9577,N_5692);
nand U10925 (N_10925,N_7758,N_6065);
or U10926 (N_10926,N_8885,N_9145);
nand U10927 (N_10927,N_7987,N_8255);
nand U10928 (N_10928,N_5178,N_7632);
nor U10929 (N_10929,N_9554,N_8788);
and U10930 (N_10930,N_6312,N_6746);
or U10931 (N_10931,N_5812,N_5608);
nand U10932 (N_10932,N_8292,N_8196);
and U10933 (N_10933,N_6729,N_8835);
or U10934 (N_10934,N_6430,N_7591);
nand U10935 (N_10935,N_9841,N_5093);
nand U10936 (N_10936,N_7988,N_9431);
nor U10937 (N_10937,N_7697,N_6171);
or U10938 (N_10938,N_5964,N_8989);
nor U10939 (N_10939,N_7929,N_7421);
and U10940 (N_10940,N_8384,N_6293);
and U10941 (N_10941,N_6044,N_7473);
nand U10942 (N_10942,N_7079,N_8992);
nor U10943 (N_10943,N_7606,N_7946);
and U10944 (N_10944,N_6451,N_8382);
nand U10945 (N_10945,N_7470,N_9102);
nand U10946 (N_10946,N_6632,N_5188);
nor U10947 (N_10947,N_6107,N_8528);
nand U10948 (N_10948,N_9282,N_8230);
and U10949 (N_10949,N_5652,N_5439);
or U10950 (N_10950,N_5492,N_5889);
and U10951 (N_10951,N_8041,N_7659);
and U10952 (N_10952,N_5762,N_9124);
and U10953 (N_10953,N_5861,N_8097);
nand U10954 (N_10954,N_6084,N_7958);
or U10955 (N_10955,N_8458,N_6921);
nor U10956 (N_10956,N_6033,N_7623);
and U10957 (N_10957,N_8934,N_9387);
and U10958 (N_10958,N_7691,N_9395);
or U10959 (N_10959,N_6561,N_7598);
or U10960 (N_10960,N_7098,N_8799);
and U10961 (N_10961,N_6069,N_5996);
and U10962 (N_10962,N_7447,N_9570);
nor U10963 (N_10963,N_5059,N_8150);
nor U10964 (N_10964,N_7891,N_7930);
nor U10965 (N_10965,N_5081,N_5012);
or U10966 (N_10966,N_8978,N_5804);
nand U10967 (N_10967,N_6569,N_5271);
and U10968 (N_10968,N_8375,N_9089);
or U10969 (N_10969,N_9615,N_6905);
and U10970 (N_10970,N_5510,N_6348);
and U10971 (N_10971,N_7925,N_5422);
nand U10972 (N_10972,N_7732,N_9754);
nor U10973 (N_10973,N_8670,N_9270);
or U10974 (N_10974,N_6156,N_5929);
nor U10975 (N_10975,N_9094,N_9566);
or U10976 (N_10976,N_6443,N_9944);
nand U10977 (N_10977,N_8029,N_6744);
nand U10978 (N_10978,N_9425,N_5381);
nor U10979 (N_10979,N_6490,N_9110);
nor U10980 (N_10980,N_6272,N_8003);
or U10981 (N_10981,N_9052,N_7619);
nor U10982 (N_10982,N_9250,N_6506);
nor U10983 (N_10983,N_5726,N_6992);
or U10984 (N_10984,N_9677,N_5282);
and U10985 (N_10985,N_9861,N_6546);
nand U10986 (N_10986,N_5937,N_5094);
and U10987 (N_10987,N_8059,N_7511);
or U10988 (N_10988,N_5217,N_6267);
or U10989 (N_10989,N_8038,N_9622);
nor U10990 (N_10990,N_9119,N_8342);
or U10991 (N_10991,N_7831,N_6056);
nor U10992 (N_10992,N_6947,N_5955);
and U10993 (N_10993,N_8345,N_6770);
nor U10994 (N_10994,N_5837,N_9731);
or U10995 (N_10995,N_7046,N_5243);
nand U10996 (N_10996,N_9602,N_6541);
and U10997 (N_10997,N_8884,N_8216);
or U10998 (N_10998,N_6461,N_9424);
nor U10999 (N_10999,N_7127,N_9575);
or U11000 (N_11000,N_7311,N_7293);
nor U11001 (N_11001,N_8764,N_9550);
nor U11002 (N_11002,N_6849,N_8999);
nor U11003 (N_11003,N_9485,N_5914);
or U11004 (N_11004,N_8780,N_8363);
and U11005 (N_11005,N_5187,N_7576);
nor U11006 (N_11006,N_6022,N_6392);
nand U11007 (N_11007,N_7266,N_9098);
nor U11008 (N_11008,N_8102,N_5250);
and U11009 (N_11009,N_6405,N_5404);
nand U11010 (N_11010,N_5084,N_6549);
nand U11011 (N_11011,N_6962,N_8935);
and U11012 (N_11012,N_5516,N_9293);
nand U11013 (N_11013,N_7427,N_6912);
or U11014 (N_11014,N_9323,N_6266);
and U11015 (N_11015,N_8654,N_6698);
nand U11016 (N_11016,N_9242,N_8579);
nor U11017 (N_11017,N_5553,N_9625);
or U11018 (N_11018,N_8302,N_7116);
nand U11019 (N_11019,N_5633,N_6809);
and U11020 (N_11020,N_9960,N_8250);
and U11021 (N_11021,N_8741,N_6787);
nor U11022 (N_11022,N_5519,N_5502);
nand U11023 (N_11023,N_6635,N_9230);
nor U11024 (N_11024,N_8898,N_8926);
or U11025 (N_11025,N_9887,N_7506);
nor U11026 (N_11026,N_9382,N_5007);
nor U11027 (N_11027,N_8062,N_6417);
and U11028 (N_11028,N_8181,N_7842);
or U11029 (N_11029,N_8512,N_9563);
nor U11030 (N_11030,N_7928,N_6035);
and U11031 (N_11031,N_5852,N_9672);
and U11032 (N_11032,N_7817,N_8550);
nor U11033 (N_11033,N_5622,N_9171);
or U11034 (N_11034,N_6019,N_5591);
nor U11035 (N_11035,N_9654,N_5663);
or U11036 (N_11036,N_5848,N_9023);
and U11037 (N_11037,N_8016,N_5928);
nor U11038 (N_11038,N_7546,N_8807);
or U11039 (N_11039,N_7246,N_8865);
or U11040 (N_11040,N_9475,N_7082);
and U11041 (N_11041,N_9345,N_8479);
or U11042 (N_11042,N_5036,N_5902);
and U11043 (N_11043,N_6482,N_9886);
nand U11044 (N_11044,N_6793,N_7349);
or U11045 (N_11045,N_8139,N_9777);
and U11046 (N_11046,N_6286,N_5406);
nor U11047 (N_11047,N_9789,N_9498);
nand U11048 (N_11048,N_5981,N_5739);
nor U11049 (N_11049,N_7811,N_9160);
or U11050 (N_11050,N_5299,N_8666);
nor U11051 (N_11051,N_5978,N_9711);
nand U11052 (N_11052,N_9633,N_9412);
nand U11053 (N_11053,N_8213,N_5759);
or U11054 (N_11054,N_6704,N_8267);
or U11055 (N_11055,N_6460,N_6187);
and U11056 (N_11056,N_8674,N_6860);
nor U11057 (N_11057,N_8809,N_6032);
nand U11058 (N_11058,N_6238,N_8401);
nand U11059 (N_11059,N_9776,N_6946);
and U11060 (N_11060,N_9709,N_7544);
or U11061 (N_11061,N_8266,N_9417);
and U11062 (N_11062,N_8165,N_8406);
or U11063 (N_11063,N_9815,N_5376);
or U11064 (N_11064,N_8610,N_5499);
nand U11065 (N_11065,N_5802,N_8091);
nor U11066 (N_11066,N_8619,N_5704);
and U11067 (N_11067,N_9968,N_7210);
nand U11068 (N_11068,N_8309,N_6961);
nor U11069 (N_11069,N_5253,N_5546);
and U11070 (N_11070,N_6966,N_5764);
and U11071 (N_11071,N_8585,N_8986);
nor U11072 (N_11072,N_6316,N_9443);
nand U11073 (N_11073,N_6674,N_6448);
and U11074 (N_11074,N_9822,N_7337);
nand U11075 (N_11075,N_7851,N_6911);
or U11076 (N_11076,N_5043,N_6711);
nor U11077 (N_11077,N_7179,N_8335);
and U11078 (N_11078,N_5733,N_9515);
or U11079 (N_11079,N_9221,N_8398);
or U11080 (N_11080,N_7705,N_6061);
and U11081 (N_11081,N_7377,N_6896);
nand U11082 (N_11082,N_5258,N_5771);
and U11083 (N_11083,N_9107,N_8356);
nor U11084 (N_11084,N_7702,N_8739);
nor U11085 (N_11085,N_7713,N_6137);
and U11086 (N_11086,N_6227,N_9671);
nor U11087 (N_11087,N_8061,N_9631);
or U11088 (N_11088,N_5104,N_7407);
or U11089 (N_11089,N_9803,N_9598);
or U11090 (N_11090,N_9992,N_5142);
or U11091 (N_11091,N_7650,N_7055);
nand U11092 (N_11092,N_5092,N_7609);
or U11093 (N_11093,N_6351,N_7467);
nor U11094 (N_11094,N_8966,N_6637);
and U11095 (N_11095,N_7192,N_7952);
nor U11096 (N_11096,N_6759,N_6273);
nor U11097 (N_11097,N_7070,N_9757);
nand U11098 (N_11098,N_8673,N_6103);
nor U11099 (N_11099,N_7213,N_7481);
and U11100 (N_11100,N_8752,N_8640);
nand U11101 (N_11101,N_6818,N_6455);
nand U11102 (N_11102,N_6113,N_9750);
nor U11103 (N_11103,N_8417,N_5110);
nand U11104 (N_11104,N_6843,N_9426);
nand U11105 (N_11105,N_9334,N_7629);
or U11106 (N_11106,N_9400,N_9311);
nor U11107 (N_11107,N_7398,N_9333);
nor U11108 (N_11108,N_9504,N_7448);
or U11109 (N_11109,N_8254,N_6679);
nor U11110 (N_11110,N_9740,N_8306);
and U11111 (N_11111,N_6690,N_9934);
or U11112 (N_11112,N_7386,N_7318);
nor U11113 (N_11113,N_6132,N_7613);
nor U11114 (N_11114,N_6878,N_8325);
nand U11115 (N_11115,N_9082,N_8759);
nand U11116 (N_11116,N_7131,N_7344);
or U11117 (N_11117,N_8546,N_6544);
nand U11118 (N_11118,N_8280,N_9801);
or U11119 (N_11119,N_9011,N_8789);
nand U11120 (N_11120,N_8556,N_9943);
or U11121 (N_11121,N_6057,N_9015);
or U11122 (N_11122,N_6391,N_8975);
nor U11123 (N_11123,N_6639,N_5657);
or U11124 (N_11124,N_5592,N_6244);
nor U11125 (N_11125,N_8473,N_7443);
nand U11126 (N_11126,N_5884,N_7163);
or U11127 (N_11127,N_7849,N_9561);
nand U11128 (N_11128,N_8974,N_9389);
nand U11129 (N_11129,N_6913,N_6367);
xnor U11130 (N_11130,N_8198,N_9128);
nor U11131 (N_11131,N_7836,N_9683);
and U11132 (N_11132,N_9249,N_8844);
or U11133 (N_11133,N_8863,N_6622);
or U11134 (N_11134,N_6235,N_7953);
nor U11135 (N_11135,N_5021,N_7735);
or U11136 (N_11136,N_5995,N_8465);
or U11137 (N_11137,N_8215,N_5938);
or U11138 (N_11138,N_5670,N_7745);
nor U11139 (N_11139,N_9808,N_7996);
or U11140 (N_11140,N_8237,N_8419);
nand U11141 (N_11141,N_5506,N_8838);
or U11142 (N_11142,N_7231,N_6015);
and U11143 (N_11143,N_9668,N_9474);
nor U11144 (N_11144,N_8470,N_6648);
nor U11145 (N_11145,N_8578,N_6994);
nand U11146 (N_11146,N_7497,N_6296);
nand U11147 (N_11147,N_7195,N_6624);
nand U11148 (N_11148,N_5834,N_8750);
nand U11149 (N_11149,N_9882,N_9012);
and U11150 (N_11150,N_6403,N_9984);
and U11151 (N_11151,N_9941,N_6996);
or U11152 (N_11152,N_8488,N_8057);
or U11153 (N_11153,N_7171,N_8549);
and U11154 (N_11154,N_7667,N_7006);
nor U11155 (N_11155,N_7002,N_7170);
or U11156 (N_11156,N_9034,N_7122);
and U11157 (N_11157,N_9350,N_6285);
or U11158 (N_11158,N_9780,N_8170);
nand U11159 (N_11159,N_8110,N_8820);
and U11160 (N_11160,N_5145,N_7096);
nor U11161 (N_11161,N_7856,N_7527);
and U11162 (N_11162,N_9788,N_6128);
and U11163 (N_11163,N_9405,N_8270);
or U11164 (N_11164,N_5645,N_5351);
and U11165 (N_11165,N_6784,N_7350);
or U11166 (N_11166,N_7043,N_5999);
nor U11167 (N_11167,N_8834,N_9367);
nand U11168 (N_11168,N_5125,N_5335);
nand U11169 (N_11169,N_9924,N_9552);
nor U11170 (N_11170,N_9341,N_7991);
nand U11171 (N_11171,N_8127,N_5218);
and U11172 (N_11172,N_6117,N_7211);
nand U11173 (N_11173,N_9202,N_9035);
nor U11174 (N_11174,N_7698,N_5991);
nor U11175 (N_11175,N_9556,N_5714);
nand U11176 (N_11176,N_6092,N_9207);
nand U11177 (N_11177,N_8543,N_7773);
or U11178 (N_11178,N_7630,N_8314);
or U11179 (N_11179,N_8813,N_7054);
nor U11180 (N_11180,N_7708,N_7636);
or U11181 (N_11181,N_8405,N_7270);
nand U11182 (N_11182,N_7528,N_7615);
and U11183 (N_11183,N_9783,N_7674);
xor U11184 (N_11184,N_8905,N_9100);
nand U11185 (N_11185,N_9328,N_5921);
and U11186 (N_11186,N_8015,N_5185);
and U11187 (N_11187,N_7157,N_8067);
nor U11188 (N_11188,N_5450,N_8818);
and U11189 (N_11189,N_9090,N_8438);
or U11190 (N_11190,N_5827,N_5445);
nor U11191 (N_11191,N_8307,N_5255);
nand U11192 (N_11192,N_5831,N_6796);
or U11193 (N_11193,N_7275,N_6563);
nand U11194 (N_11194,N_6486,N_8249);
and U11195 (N_11195,N_7081,N_5303);
nand U11196 (N_11196,N_6352,N_9385);
nor U11197 (N_11197,N_7314,N_6670);
or U11198 (N_11198,N_5011,N_5513);
nand U11199 (N_11199,N_6122,N_7814);
and U11200 (N_11200,N_7568,N_7816);
or U11201 (N_11201,N_5058,N_9366);
nor U11202 (N_11202,N_6088,N_8204);
and U11203 (N_11203,N_8017,N_6612);
and U11204 (N_11204,N_9093,N_7196);
nand U11205 (N_11205,N_7760,N_5086);
nand U11206 (N_11206,N_6484,N_5952);
or U11207 (N_11207,N_5075,N_6567);
nor U11208 (N_11208,N_8137,N_6964);
or U11209 (N_11209,N_7263,N_5167);
nand U11210 (N_11210,N_6685,N_6865);
nor U11211 (N_11211,N_7248,N_6164);
or U11212 (N_11212,N_5017,N_7824);
or U11213 (N_11213,N_5744,N_6337);
nor U11214 (N_11214,N_5211,N_6958);
or U11215 (N_11215,N_6611,N_9224);
or U11216 (N_11216,N_7781,N_5460);
or U11217 (N_11217,N_9835,N_5157);
and U11218 (N_11218,N_7184,N_5676);
or U11219 (N_11219,N_7058,N_8275);
nand U11220 (N_11220,N_6407,N_9476);
or U11221 (N_11221,N_6811,N_9077);
and U11222 (N_11222,N_9185,N_7371);
or U11223 (N_11223,N_7829,N_5413);
nand U11224 (N_11224,N_6908,N_7330);
nor U11225 (N_11225,N_7316,N_5723);
nor U11226 (N_11226,N_7704,N_6453);
nand U11227 (N_11227,N_9660,N_8443);
and U11228 (N_11228,N_8625,N_9830);
and U11229 (N_11229,N_8338,N_7296);
or U11230 (N_11230,N_8011,N_7685);
or U11231 (N_11231,N_6776,N_7771);
nor U11232 (N_11232,N_8630,N_9850);
nor U11233 (N_11233,N_9222,N_7235);
or U11234 (N_11234,N_7641,N_6457);
nand U11235 (N_11235,N_8700,N_5378);
nand U11236 (N_11236,N_9267,N_5317);
or U11237 (N_11237,N_8603,N_9372);
and U11238 (N_11238,N_8354,N_7728);
or U11239 (N_11239,N_8048,N_5641);
or U11240 (N_11240,N_8226,N_5437);
and U11241 (N_11241,N_7841,N_8032);
or U11242 (N_11242,N_6853,N_8515);
nor U11243 (N_11243,N_5769,N_9951);
nor U11244 (N_11244,N_5625,N_7907);
or U11245 (N_11245,N_8801,N_5245);
and U11246 (N_11246,N_7575,N_5575);
or U11247 (N_11247,N_6686,N_5111);
nor U11248 (N_11248,N_7370,N_6673);
or U11249 (N_11249,N_7723,N_8725);
nor U11250 (N_11250,N_6071,N_5471);
nand U11251 (N_11251,N_9406,N_6418);
nor U11252 (N_11252,N_5158,N_6974);
or U11253 (N_11253,N_8972,N_8595);
or U11254 (N_11254,N_8592,N_5808);
nor U11255 (N_11255,N_8724,N_5715);
and U11256 (N_11256,N_7681,N_8288);
xnor U11257 (N_11257,N_9099,N_8949);
nor U11258 (N_11258,N_6003,N_5651);
and U11259 (N_11259,N_9306,N_7147);
and U11260 (N_11260,N_7737,N_7091);
and U11261 (N_11261,N_9821,N_6603);
nor U11262 (N_11262,N_6756,N_7700);
nor U11263 (N_11263,N_5390,N_6358);
or U11264 (N_11264,N_8756,N_5479);
and U11265 (N_11265,N_6039,N_5144);
or U11266 (N_11266,N_9948,N_6604);
and U11267 (N_11267,N_5535,N_7044);
and U11268 (N_11268,N_9910,N_5318);
nand U11269 (N_11269,N_9225,N_6834);
or U11270 (N_11270,N_8414,N_7789);
and U11271 (N_11271,N_5768,N_5423);
nor U11272 (N_11272,N_5574,N_7866);
or U11273 (N_11273,N_7710,N_5392);
nor U11274 (N_11274,N_7441,N_7676);
nand U11275 (N_11275,N_5639,N_9005);
or U11276 (N_11276,N_8373,N_8201);
and U11277 (N_11277,N_8622,N_7977);
or U11278 (N_11278,N_9555,N_5280);
or U11279 (N_11279,N_9922,N_7146);
nor U11280 (N_11280,N_7405,N_6519);
and U11281 (N_11281,N_6518,N_9690);
nand U11282 (N_11282,N_6995,N_5755);
nor U11283 (N_11283,N_5320,N_7101);
nor U11284 (N_11284,N_6250,N_8163);
nand U11285 (N_11285,N_5176,N_5810);
and U11286 (N_11286,N_8876,N_9623);
and U11287 (N_11287,N_8104,N_5448);
or U11288 (N_11288,N_8323,N_6234);
or U11289 (N_11289,N_7775,N_6737);
and U11290 (N_11290,N_7149,N_5359);
nand U11291 (N_11291,N_7130,N_6581);
nor U11292 (N_11292,N_6783,N_9975);
or U11293 (N_11293,N_5161,N_6163);
or U11294 (N_11294,N_6513,N_7652);
nand U11295 (N_11295,N_6663,N_5286);
xnor U11296 (N_11296,N_6202,N_8833);
and U11297 (N_11297,N_7807,N_9703);
or U11298 (N_11298,N_9047,N_5440);
nand U11299 (N_11299,N_9512,N_5032);
nand U11300 (N_11300,N_6538,N_5705);
and U11301 (N_11301,N_5350,N_5389);
or U11302 (N_11302,N_7736,N_8378);
nor U11303 (N_11303,N_5379,N_8040);
nand U11304 (N_11304,N_6733,N_9313);
nand U11305 (N_11305,N_5677,N_6496);
or U11306 (N_11306,N_6917,N_8191);
or U11307 (N_11307,N_5799,N_9115);
nand U11308 (N_11308,N_8188,N_7880);
nor U11309 (N_11309,N_5864,N_9496);
or U11310 (N_11310,N_7921,N_5472);
and U11311 (N_11311,N_6959,N_6514);
nor U11312 (N_11312,N_8867,N_7812);
or U11313 (N_11313,N_9087,N_7690);
xnor U11314 (N_11314,N_6862,N_6548);
or U11315 (N_11315,N_5785,N_8562);
nand U11316 (N_11316,N_7492,N_5655);
nand U11317 (N_11317,N_9059,N_9859);
nand U11318 (N_11318,N_8503,N_7222);
or U11319 (N_11319,N_8276,N_5429);
nand U11320 (N_11320,N_5897,N_8012);
or U11321 (N_11321,N_8551,N_5120);
or U11322 (N_11322,N_5300,N_9522);
and U11323 (N_11323,N_9231,N_9439);
or U11324 (N_11324,N_5139,N_8221);
nor U11325 (N_11325,N_7125,N_7080);
nand U11326 (N_11326,N_9113,N_8272);
nand U11327 (N_11327,N_6785,N_9068);
nand U11328 (N_11328,N_5881,N_9462);
and U11329 (N_11329,N_5034,N_7748);
nand U11330 (N_11330,N_5638,N_9967);
or U11331 (N_11331,N_5717,N_8239);
nor U11332 (N_11332,N_9929,N_9455);
and U11333 (N_11333,N_9956,N_7919);
and U11334 (N_11334,N_5174,N_8116);
nand U11335 (N_11335,N_6002,N_6034);
or U11336 (N_11336,N_7475,N_7712);
nor U11337 (N_11337,N_9571,N_7854);
and U11338 (N_11338,N_9461,N_9529);
or U11339 (N_11339,N_7440,N_6762);
nor U11340 (N_11340,N_8284,N_9440);
nor U11341 (N_11341,N_5721,N_8558);
nand U11342 (N_11342,N_6143,N_8646);
or U11343 (N_11343,N_5586,N_8073);
nor U11344 (N_11344,N_5153,N_8708);
nor U11345 (N_11345,N_7545,N_9921);
and U11346 (N_11346,N_5453,N_5388);
nand U11347 (N_11347,N_6116,N_7523);
nand U11348 (N_11348,N_7451,N_5209);
nor U11349 (N_11349,N_5239,N_5098);
or U11350 (N_11350,N_6532,N_7542);
or U11351 (N_11351,N_7267,N_7911);
or U11352 (N_11352,N_5588,N_6254);
or U11353 (N_11353,N_9751,N_6435);
and U11354 (N_11354,N_8364,N_9008);
or U11355 (N_11355,N_8757,N_8945);
or U11356 (N_11356,N_7868,N_9120);
or U11357 (N_11357,N_5600,N_7818);
nor U11358 (N_11358,N_8459,N_6447);
nand U11359 (N_11359,N_5044,N_8929);
or U11360 (N_11360,N_8698,N_9364);
nor U11361 (N_11361,N_9767,N_6108);
or U11362 (N_11362,N_6445,N_9686);
nand U11363 (N_11363,N_5405,N_6568);
nand U11364 (N_11364,N_5660,N_6584);
and U11365 (N_11365,N_9186,N_7635);
and U11366 (N_11366,N_9965,N_5477);
nand U11367 (N_11367,N_5159,N_8651);
or U11368 (N_11368,N_6576,N_8171);
nand U11369 (N_11369,N_8118,N_5650);
nand U11370 (N_11370,N_7769,N_8858);
and U11371 (N_11371,N_7599,N_6237);
nand U11372 (N_11372,N_8173,N_9024);
and U11373 (N_11373,N_9394,N_6162);
or U11374 (N_11374,N_9365,N_6230);
nand U11375 (N_11375,N_8775,N_7717);
xor U11376 (N_11376,N_5304,N_6408);
and U11377 (N_11377,N_8019,N_9201);
or U11378 (N_11378,N_8103,N_8753);
nand U11379 (N_11379,N_8160,N_6492);
nor U11380 (N_11380,N_8141,N_8129);
nand U11381 (N_11381,N_5292,N_8308);
or U11382 (N_11382,N_9953,N_5594);
nand U11383 (N_11383,N_9209,N_7791);
or U11384 (N_11384,N_8814,N_6507);
nand U11385 (N_11385,N_9763,N_7333);
nand U11386 (N_11386,N_9567,N_8370);
or U11387 (N_11387,N_7215,N_5337);
or U11388 (N_11388,N_6179,N_9336);
and U11389 (N_11389,N_5871,N_5979);
nand U11390 (N_11390,N_5643,N_5616);
nor U11391 (N_11391,N_6168,N_8916);
xnor U11392 (N_11392,N_6588,N_5695);
nand U11393 (N_11393,N_9196,N_5501);
or U11394 (N_11394,N_8366,N_7140);
nand U11395 (N_11395,N_6928,N_5737);
or U11396 (N_11396,N_5947,N_7345);
or U11397 (N_11397,N_8829,N_7057);
nor U11398 (N_11398,N_6982,N_5354);
or U11399 (N_11399,N_5935,N_5324);
and U11400 (N_11400,N_9246,N_8502);
or U11401 (N_11401,N_8518,N_5631);
or U11402 (N_11402,N_7541,N_8760);
nor U11403 (N_11403,N_7074,N_7260);
nand U11404 (N_11404,N_8831,N_6243);
and U11405 (N_11405,N_7759,N_6916);
nand U11406 (N_11406,N_6642,N_8719);
nand U11407 (N_11407,N_7359,N_7795);
nand U11408 (N_11408,N_6620,N_7094);
nand U11409 (N_11409,N_9508,N_5888);
nor U11410 (N_11410,N_8887,N_7389);
and U11411 (N_11411,N_7457,N_7269);
or U11412 (N_11412,N_5845,N_9088);
nand U11413 (N_11413,N_8608,N_8607);
nor U11414 (N_11414,N_7714,N_5585);
and U11415 (N_11415,N_7520,N_5738);
nand U11416 (N_11416,N_7329,N_7768);
or U11417 (N_11417,N_8832,N_5189);
or U11418 (N_11418,N_6515,N_6066);
and U11419 (N_11419,N_9450,N_6388);
xor U11420 (N_11420,N_5382,N_5396);
and U11421 (N_11421,N_7621,N_6279);
nor U11422 (N_11422,N_9521,N_9580);
nand U11423 (N_11423,N_6831,N_7893);
nand U11424 (N_11424,N_9132,N_5675);
nand U11425 (N_11425,N_5462,N_5019);
or U11426 (N_11426,N_7302,N_8131);
nor U11427 (N_11427,N_7027,N_8047);
nor U11428 (N_11428,N_9534,N_7980);
nor U11429 (N_11429,N_9126,N_5876);
nand U11430 (N_11430,N_8441,N_7134);
nor U11431 (N_11431,N_6852,N_9576);
nand U11432 (N_11432,N_5728,N_9541);
and U11433 (N_11433,N_8389,N_5426);
xnor U11434 (N_11434,N_5205,N_6551);
nand U11435 (N_11435,N_9146,N_7013);
xnor U11436 (N_11436,N_6951,N_6653);
or U11437 (N_11437,N_7522,N_7584);
nand U11438 (N_11438,N_5572,N_9976);
nand U11439 (N_11439,N_9500,N_6773);
nand U11440 (N_11440,N_5874,N_8352);
and U11441 (N_11441,N_9994,N_9217);
nand U11442 (N_11442,N_9030,N_5476);
nand U11443 (N_11443,N_8260,N_6438);
nor U11444 (N_11444,N_7390,N_5247);
or U11445 (N_11445,N_6170,N_9203);
or U11446 (N_11446,N_5373,N_9383);
or U11447 (N_11447,N_8522,N_5457);
nand U11448 (N_11448,N_6971,N_8690);
nor U11449 (N_11449,N_8857,N_8222);
nand U11450 (N_11450,N_6147,N_8159);
and U11451 (N_11451,N_7075,N_9103);
or U11452 (N_11452,N_5341,N_5687);
or U11453 (N_11453,N_8924,N_7038);
and U11454 (N_11454,N_5257,N_7118);
and U11455 (N_11455,N_6494,N_9466);
nand U11456 (N_11456,N_6321,N_7885);
nand U11457 (N_11457,N_7059,N_9845);
or U11458 (N_11458,N_9471,N_5010);
and U11459 (N_11459,N_6274,N_8193);
nand U11460 (N_11460,N_5746,N_6290);
nand U11461 (N_11461,N_8922,N_9787);
nand U11462 (N_11462,N_5526,N_6102);
or U11463 (N_11463,N_7805,N_7718);
nand U11464 (N_11464,N_5030,N_6939);
nand U11465 (N_11465,N_9092,N_8289);
and U11466 (N_11466,N_5710,N_6464);
or U11467 (N_11467,N_5541,N_8505);
nand U11468 (N_11468,N_5296,N_6320);
and U11469 (N_11469,N_6832,N_6462);
nand U11470 (N_11470,N_6087,N_6341);
or U11471 (N_11471,N_7954,N_5135);
or U11472 (N_11472,N_9167,N_7550);
nand U11473 (N_11473,N_9044,N_6979);
and U11474 (N_11474,N_9536,N_7968);
nor U11475 (N_11475,N_8510,N_5238);
and U11476 (N_11476,N_7480,N_9867);
and U11477 (N_11477,N_9670,N_5190);
nor U11478 (N_11478,N_6134,N_5598);
and U11479 (N_11479,N_9036,N_5615);
or U11480 (N_11480,N_9320,N_8772);
nand U11481 (N_11481,N_8943,N_8271);
and U11482 (N_11482,N_7556,N_8135);
and U11483 (N_11483,N_8351,N_6051);
or U11484 (N_11484,N_7657,N_5356);
and U11485 (N_11485,N_5353,N_8848);
or U11486 (N_11486,N_6730,N_9149);
or U11487 (N_11487,N_6307,N_6263);
nor U11488 (N_11488,N_5850,N_8295);
xnor U11489 (N_11489,N_8186,N_8484);
or U11490 (N_11490,N_8968,N_5228);
or U11491 (N_11491,N_7782,N_7029);
or U11492 (N_11492,N_8882,N_9885);
or U11493 (N_11493,N_6585,N_9810);
or U11494 (N_11494,N_8229,N_9773);
nor U11495 (N_11495,N_8983,N_6537);
nor U11496 (N_11496,N_8774,N_7292);
nor U11497 (N_11497,N_8768,N_8411);
nor U11498 (N_11498,N_5751,N_9025);
nand U11499 (N_11499,N_7660,N_7587);
and U11500 (N_11500,N_5152,N_6617);
nor U11501 (N_11501,N_5117,N_9151);
or U11502 (N_11502,N_7804,N_6678);
and U11503 (N_11503,N_5340,N_9872);
or U11504 (N_11504,N_8400,N_7312);
or U11505 (N_11505,N_8326,N_5696);
and U11506 (N_11506,N_7815,N_9651);
nor U11507 (N_11507,N_7439,N_9936);
or U11508 (N_11508,N_6651,N_5790);
or U11509 (N_11509,N_5485,N_7288);
nor U11510 (N_11510,N_8444,N_5840);
nand U11511 (N_11511,N_7762,N_7834);
nand U11512 (N_11512,N_9665,N_7247);
nand U11513 (N_11513,N_7935,N_9140);
nor U11514 (N_11514,N_5731,N_7285);
and U11515 (N_11515,N_9745,N_9363);
and U11516 (N_11516,N_8609,N_8588);
nor U11517 (N_11517,N_5045,N_7833);
or U11518 (N_11518,N_5226,N_7488);
nor U11519 (N_11519,N_8187,N_8415);
nor U11520 (N_11520,N_7764,N_8629);
or U11521 (N_11521,N_5860,N_7401);
and U11522 (N_11522,N_7021,N_9244);
nand U11523 (N_11523,N_9006,N_6196);
and U11524 (N_11524,N_7456,N_9080);
and U11525 (N_11525,N_6450,N_9901);
nand U11526 (N_11526,N_7870,N_9513);
and U11527 (N_11527,N_8946,N_9097);
or U11528 (N_11528,N_6345,N_9420);
nand U11529 (N_11529,N_7547,N_8418);
nand U11530 (N_11530,N_6200,N_6719);
and U11531 (N_11531,N_5693,N_8862);
and U11532 (N_11532,N_5880,N_7624);
or U11533 (N_11533,N_7549,N_8996);
and U11534 (N_11534,N_8136,N_9700);
or U11535 (N_11535,N_9407,N_9452);
and U11536 (N_11536,N_9211,N_7168);
nor U11537 (N_11537,N_5961,N_7853);
nand U11538 (N_11538,N_5798,N_6606);
or U11539 (N_11539,N_8797,N_5628);
xnor U11540 (N_11540,N_8075,N_8914);
or U11541 (N_11541,N_6219,N_7351);
nand U11542 (N_11542,N_9172,N_9878);
or U11543 (N_11543,N_9752,N_8294);
or U11544 (N_11544,N_7945,N_9621);
xor U11545 (N_11545,N_8795,N_8433);
or U11546 (N_11546,N_5898,N_7462);
or U11547 (N_11547,N_9989,N_6025);
nand U11548 (N_11548,N_9819,N_6370);
or U11549 (N_11549,N_8526,N_9219);
or U11550 (N_11550,N_9227,N_7045);
nor U11551 (N_11551,N_9579,N_7209);
and U11552 (N_11552,N_5344,N_9704);
or U11553 (N_11553,N_9778,N_8868);
nand U11554 (N_11554,N_8231,N_5844);
or U11555 (N_11555,N_5873,N_5773);
nand U11556 (N_11556,N_9509,N_5287);
and U11557 (N_11557,N_5172,N_5892);
nor U11558 (N_11558,N_7733,N_6547);
nand U11559 (N_11559,N_6634,N_5683);
nor U11560 (N_11560,N_8947,N_7326);
and U11561 (N_11561,N_8492,N_6055);
or U11562 (N_11562,N_7216,N_9505);
and U11563 (N_11563,N_9565,N_8259);
xnor U11564 (N_11564,N_9318,N_7658);
and U11565 (N_11565,N_7975,N_7731);
nor U11566 (N_11566,N_7403,N_9308);
nor U11567 (N_11567,N_5975,N_6471);
nor U11568 (N_11568,N_8053,N_8860);
nor U11569 (N_11569,N_5735,N_9432);
or U11570 (N_11570,N_5198,N_5532);
and U11571 (N_11571,N_7273,N_5926);
nor U11572 (N_11572,N_8736,N_5395);
or U11573 (N_11573,N_5090,N_8783);
or U11574 (N_11574,N_9868,N_5515);
and U11575 (N_11575,N_6805,N_9970);
nor U11576 (N_11576,N_9593,N_8658);
or U11577 (N_11577,N_8819,N_6161);
and U11578 (N_11578,N_9058,N_5573);
and U11579 (N_11579,N_6669,N_6252);
and U11580 (N_11580,N_5922,N_7766);
and U11581 (N_11581,N_6076,N_7167);
nor U11582 (N_11582,N_6619,N_5977);
or U11583 (N_11583,N_9262,N_6357);
and U11584 (N_11584,N_8747,N_9162);
or U11585 (N_11585,N_6528,N_9187);
and U11586 (N_11586,N_7201,N_7362);
nor U11587 (N_11587,N_5469,N_5433);
nor U11588 (N_11588,N_6857,N_7278);
nand U11589 (N_11589,N_5331,N_9939);
nand U11590 (N_11590,N_7992,N_8532);
nor U11591 (N_11591,N_9837,N_5233);
or U11592 (N_11592,N_6819,N_6253);
xor U11593 (N_11593,N_8248,N_6479);
nor U11594 (N_11594,N_8334,N_8816);
or U11595 (N_11595,N_8208,N_7145);
and U11596 (N_11596,N_7720,N_7388);
nor U11597 (N_11597,N_9825,N_7765);
nor U11598 (N_11598,N_5386,N_7750);
or U11599 (N_11599,N_5184,N_8964);
or U11600 (N_11600,N_8134,N_5313);
nand U11601 (N_11601,N_7088,N_6900);
nor U11602 (N_11602,N_8300,N_6401);
nor U11603 (N_11603,N_6119,N_8536);
and U11604 (N_11604,N_8332,N_6914);
and U11605 (N_11605,N_7501,N_7730);
nand U11606 (N_11606,N_8617,N_8084);
nor U11607 (N_11607,N_7608,N_6910);
nor U11608 (N_11608,N_9890,N_7979);
or U11609 (N_11609,N_9915,N_7310);
nand U11610 (N_11610,N_8675,N_6199);
nor U11611 (N_11611,N_5596,N_8830);
nand U11612 (N_11612,N_8174,N_8909);
nor U11613 (N_11613,N_6259,N_8305);
or U11614 (N_11614,N_5412,N_5130);
and U11615 (N_11615,N_6166,N_5212);
nand U11616 (N_11616,N_8085,N_8392);
nor U11617 (N_11617,N_8987,N_9195);
nand U11618 (N_11618,N_7007,N_5882);
nand U11619 (N_11619,N_7962,N_8985);
or U11620 (N_11620,N_8650,N_9199);
or U11621 (N_11621,N_7298,N_9238);
nor U11622 (N_11622,N_9331,N_8555);
nor U11623 (N_11623,N_5727,N_8089);
and U11624 (N_11624,N_9610,N_9017);
or U11625 (N_11625,N_6029,N_6897);
or U11626 (N_11626,N_9844,N_5885);
or U11627 (N_11627,N_7418,N_5277);
or U11628 (N_11628,N_8200,N_5869);
nand U11629 (N_11629,N_7861,N_8368);
or U11630 (N_11630,N_9236,N_5041);
and U11631 (N_11631,N_5355,N_6643);
or U11632 (N_11632,N_5842,N_9795);
nand U11633 (N_11633,N_9983,N_9129);
or U11634 (N_11634,N_5910,N_7683);
or U11635 (N_11635,N_8371,N_7455);
nand U11636 (N_11636,N_5847,N_6735);
or U11637 (N_11637,N_8431,N_6360);
or U11638 (N_11638,N_9540,N_7010);
and U11639 (N_11639,N_9658,N_8277);
and U11640 (N_11640,N_8963,N_9422);
and U11641 (N_11641,N_8932,N_7671);
nor U11642 (N_11642,N_5414,N_6542);
nor U11643 (N_11643,N_5567,N_7798);
nor U11644 (N_11644,N_6872,N_5403);
nand U11645 (N_11645,N_5582,N_5832);
or U11646 (N_11646,N_8530,N_9608);
or U11647 (N_11647,N_6224,N_8262);
nand U11648 (N_11648,N_9050,N_5006);
and U11649 (N_11649,N_6779,N_7114);
nand U11650 (N_11650,N_5263,N_7903);
nand U11651 (N_11651,N_9239,N_8871);
or U11652 (N_11652,N_8388,N_9438);
and U11653 (N_11653,N_7558,N_6760);
or U11654 (N_11654,N_8615,N_6277);
and U11655 (N_11655,N_6297,N_9597);
nand U11656 (N_11656,N_8194,N_8805);
xnor U11657 (N_11657,N_7533,N_7662);
or U11658 (N_11658,N_5063,N_5634);
or U11659 (N_11659,N_8612,N_8841);
nor U11660 (N_11660,N_9176,N_5147);
and U11661 (N_11661,N_7602,N_6242);
or U11662 (N_11662,N_6557,N_6292);
nor U11663 (N_11663,N_5121,N_5821);
and U11664 (N_11664,N_9163,N_6877);
nand U11665 (N_11665,N_7182,N_7255);
and U11666 (N_11666,N_7051,N_9223);
and U11667 (N_11667,N_7601,N_8008);
nor U11668 (N_11668,N_8699,N_9646);
nor U11669 (N_11669,N_5427,N_6732);
and U11670 (N_11670,N_6144,N_5967);
nand U11671 (N_11671,N_8044,N_5343);
and U11672 (N_11672,N_6935,N_9494);
nor U11673 (N_11673,N_5525,N_7042);
and U11674 (N_11674,N_5566,N_5251);
and U11675 (N_11675,N_9748,N_7137);
nand U11676 (N_11676,N_7626,N_9177);
nor U11677 (N_11677,N_5786,N_9263);
or U11678 (N_11678,N_7126,N_7845);
or U11679 (N_11679,N_5857,N_6380);
nand U11680 (N_11680,N_5971,N_7924);
nand U11681 (N_11681,N_6850,N_9549);
nand U11682 (N_11682,N_6436,N_7017);
and U11683 (N_11683,N_8212,N_7108);
or U11684 (N_11684,N_6152,N_7004);
xor U11685 (N_11685,N_8318,N_8313);
and U11686 (N_11686,N_6564,N_5193);
nand U11687 (N_11687,N_7687,N_5559);
and U11688 (N_11688,N_8712,N_8092);
nand U11689 (N_11689,N_8140,N_8257);
nand U11690 (N_11690,N_6211,N_7564);
or U11691 (N_11691,N_9611,N_5983);
or U11692 (N_11692,N_8804,N_6823);
nor U11693 (N_11693,N_5256,N_6924);
nor U11694 (N_11694,N_8993,N_6918);
nor U11695 (N_11695,N_9477,N_8886);
nand U11696 (N_11696,N_7416,N_8397);
or U11697 (N_11697,N_8210,N_6804);
nand U11698 (N_11698,N_9348,N_9828);
and U11699 (N_11699,N_9659,N_9260);
nand U11700 (N_11700,N_7450,N_7280);
or U11701 (N_11701,N_9031,N_5241);
or U11702 (N_11702,N_8959,N_7822);
nor U11703 (N_11703,N_6866,N_6251);
nand U11704 (N_11704,N_7668,N_7406);
nand U11705 (N_11705,N_8716,N_6970);
and U11706 (N_11706,N_7820,N_7306);
nor U11707 (N_11707,N_5325,N_6325);
nand U11708 (N_11708,N_8330,N_6649);
nand U11709 (N_11709,N_8506,N_9411);
and U11710 (N_11710,N_6130,N_9762);
nand U11711 (N_11711,N_7352,N_9480);
and U11712 (N_11712,N_6936,N_9154);
nor U11713 (N_11713,N_7056,N_5851);
or U11714 (N_11714,N_7023,N_9812);
nand U11715 (N_11715,N_9641,N_9938);
nor U11716 (N_11716,N_5138,N_9456);
or U11717 (N_11717,N_5231,N_5698);
or U11718 (N_11718,N_5080,N_6708);
or U11719 (N_11719,N_5481,N_8452);
nor U11720 (N_11720,N_6332,N_7226);
nor U11721 (N_11721,N_9310,N_8393);
nand U11722 (N_11722,N_5478,N_5383);
or U11723 (N_11723,N_5520,N_6323);
and U11724 (N_11724,N_5038,N_5509);
or U11725 (N_11725,N_5934,N_6248);
nand U11726 (N_11726,N_7321,N_5954);
nor U11727 (N_11727,N_9375,N_7284);
nand U11728 (N_11728,N_7336,N_8482);
nor U11729 (N_11729,N_5583,N_7373);
nand U11730 (N_11730,N_6607,N_9537);
nand U11731 (N_11731,N_8842,N_5430);
nor U11732 (N_11732,N_8910,N_6997);
nand U11733 (N_11733,N_5047,N_9354);
or U11734 (N_11734,N_7534,N_9649);
nand U11735 (N_11735,N_9309,N_9586);
or U11736 (N_11736,N_7369,N_7419);
or U11737 (N_11737,N_8815,N_5579);
and U11738 (N_11738,N_5039,N_8079);
nor U11739 (N_11739,N_6825,N_7585);
or U11740 (N_11740,N_6322,N_5915);
or U11741 (N_11741,N_6824,N_5635);
nand U11742 (N_11742,N_9933,N_7967);
or U11743 (N_11743,N_6873,N_5346);
or U11744 (N_11744,N_9204,N_5169);
nor U11745 (N_11745,N_6536,N_7524);
and U11746 (N_11746,N_7934,N_9932);
nand U11747 (N_11747,N_7295,N_7272);
nor U11748 (N_11748,N_8068,N_9814);
nand U11749 (N_11749,N_6904,N_7666);
nand U11750 (N_11750,N_6381,N_8074);
or U11751 (N_11751,N_7680,N_9634);
or U11752 (N_11752,N_9003,N_7786);
nor U11753 (N_11753,N_7603,N_7154);
nor U11754 (N_11754,N_6595,N_7819);
nand U11755 (N_11755,N_6439,N_8244);
nor U11756 (N_11756,N_7324,N_8524);
nand U11757 (N_11757,N_9644,N_7612);
and U11758 (N_11758,N_9779,N_8811);
nor U11759 (N_11759,N_7452,N_8169);
and U11760 (N_11760,N_9233,N_9192);
nor U11761 (N_11761,N_5968,N_8301);
nor U11762 (N_11762,N_9635,N_9906);
or U11763 (N_11763,N_6890,N_7052);
nor U11764 (N_11764,N_7796,N_9469);
or U11765 (N_11765,N_7679,N_7772);
nor U11766 (N_11766,N_6956,N_6067);
nor U11767 (N_11767,N_6394,N_5770);
or U11768 (N_11768,N_8611,N_9358);
nor U11769 (N_11769,N_8077,N_5793);
xnor U11770 (N_11770,N_9349,N_5004);
or U11771 (N_11771,N_7508,N_6406);
and U11772 (N_11772,N_8353,N_8228);
nor U11773 (N_11773,N_7279,N_9289);
nand U11774 (N_11774,N_8685,N_7412);
nor U11775 (N_11775,N_8634,N_6692);
nand U11776 (N_11776,N_6173,N_8072);
nand U11777 (N_11777,N_5160,N_7947);
nand U11778 (N_11778,N_5956,N_9873);
nor U11779 (N_11779,N_7150,N_6665);
nand U11780 (N_11780,N_8341,N_6305);
and U11781 (N_11781,N_7120,N_7331);
nor U11782 (N_11782,N_5366,N_9775);
and U11783 (N_11783,N_7505,N_7863);
or U11784 (N_11784,N_5347,N_6753);
or U11785 (N_11785,N_7514,N_9133);
nor U11786 (N_11786,N_6540,N_8158);
and U11787 (N_11787,N_6718,N_8737);
nor U11788 (N_11788,N_5182,N_9288);
xor U11789 (N_11789,N_6058,N_9020);
or U11790 (N_11790,N_5618,N_7112);
or U11791 (N_11791,N_5279,N_8742);
and U11792 (N_11792,N_6387,N_5269);
and U11793 (N_11793,N_9490,N_9381);
nand U11794 (N_11794,N_6505,N_9578);
or U11795 (N_11795,N_7855,N_9391);
nor U11796 (N_11796,N_6282,N_9193);
nor U11797 (N_11797,N_9583,N_5732);
and U11798 (N_11798,N_7823,N_6854);
nand U11799 (N_11799,N_5630,N_8782);
or U11800 (N_11800,N_5301,N_7985);
and U11801 (N_11801,N_9811,N_8252);
and U11802 (N_11802,N_9026,N_5896);
nand U11803 (N_11803,N_9736,N_6000);
or U11804 (N_11804,N_7675,N_8911);
and U11805 (N_11805,N_9401,N_7995);
nor U11806 (N_11806,N_8183,N_5547);
or U11807 (N_11807,N_8956,N_8645);
or U11808 (N_11808,N_8544,N_6127);
and U11809 (N_11809,N_9722,N_9174);
nor U11810 (N_11810,N_8894,N_7752);
and U11811 (N_11811,N_6695,N_6938);
or U11812 (N_11812,N_8303,N_9464);
nor U11813 (N_11813,N_6343,N_9096);
nand U11814 (N_11814,N_7531,N_6192);
or U11815 (N_11815,N_6968,N_6231);
and U11816 (N_11816,N_5742,N_9123);
nor U11817 (N_11817,N_7722,N_8426);
nand U11818 (N_11818,N_6614,N_8081);
or U11819 (N_11819,N_7913,N_9314);
or U11820 (N_11820,N_8463,N_9449);
nand U11821 (N_11821,N_8495,N_5224);
or U11822 (N_11822,N_6349,N_8695);
or U11823 (N_11823,N_9416,N_8694);
and U11824 (N_11824,N_8298,N_5932);
nand U11825 (N_11825,N_5906,N_9142);
and U11826 (N_11826,N_6398,N_7433);
and U11827 (N_11827,N_9454,N_5339);
or U11828 (N_11828,N_8960,N_6830);
or U11829 (N_11829,N_7744,N_7180);
and U11830 (N_11830,N_7997,N_7317);
and U11831 (N_11831,N_8207,N_5214);
and U11832 (N_11832,N_7826,N_6583);
nor U11833 (N_11833,N_6525,N_5290);
and U11834 (N_11834,N_7060,N_7385);
or U11835 (N_11835,N_7265,N_7048);
and U11836 (N_11836,N_9444,N_6379);
nand U11837 (N_11837,N_5843,N_6115);
nor U11838 (N_11838,N_5554,N_5558);
or U11839 (N_11839,N_5524,N_8437);
and U11840 (N_11840,N_6024,N_8869);
nor U11841 (N_11841,N_5772,N_8346);
nand U11842 (N_11842,N_9104,N_9033);
or U11843 (N_11843,N_9130,N_8167);
nand U11844 (N_11844,N_6855,N_9966);
and U11845 (N_11845,N_5818,N_8778);
nand U11846 (N_11846,N_5976,N_8888);
or U11847 (N_11847,N_8035,N_9898);
and U11848 (N_11848,N_9935,N_7579);
nand U11849 (N_11849,N_8265,N_5206);
nand U11850 (N_11850,N_8707,N_8919);
nor U11851 (N_11851,N_5394,N_5988);
nor U11852 (N_11852,N_7502,N_9213);
nor U11853 (N_11853,N_7963,N_5606);
nor U11854 (N_11854,N_8245,N_6210);
nand U11855 (N_11855,N_8624,N_9715);
or U11856 (N_11856,N_7825,N_5766);
or U11857 (N_11857,N_9470,N_6794);
nand U11858 (N_11858,N_5195,N_5082);
nor U11859 (N_11859,N_6091,N_7910);
or U11860 (N_11860,N_9048,N_7530);
or U11861 (N_11861,N_5148,N_6976);
or U11862 (N_11862,N_8304,N_7944);
and U11863 (N_11863,N_8423,N_5903);
nor U11864 (N_11864,N_7415,N_6722);
nor U11865 (N_11865,N_5709,N_8586);
and U11866 (N_11866,N_5817,N_7410);
nor U11867 (N_11867,N_9676,N_7271);
or U11868 (N_11868,N_8897,N_5026);
nor U11869 (N_11869,N_9727,N_5447);
nand U11870 (N_11870,N_7957,N_5106);
and U11871 (N_11871,N_8422,N_8889);
and U11872 (N_11872,N_8420,N_5431);
or U11873 (N_11873,N_7238,N_7259);
and U11874 (N_11874,N_7999,N_6400);
or U11875 (N_11875,N_5522,N_5686);
and U11876 (N_11876,N_5294,N_8477);
nor U11877 (N_11877,N_9771,N_9415);
nand U11878 (N_11878,N_9169,N_5073);
and U11879 (N_11879,N_7899,N_7993);
nor U11880 (N_11880,N_5823,N_6121);
nor U11881 (N_11881,N_6662,N_8846);
nand U11882 (N_11882,N_8453,N_5109);
nand U11883 (N_11883,N_9902,N_8310);
nand U11884 (N_11884,N_7387,N_5262);
and U11885 (N_11885,N_9701,N_9273);
or U11886 (N_11886,N_9675,N_8018);
nand U11887 (N_11887,N_9027,N_9730);
nand U11888 (N_11888,N_5463,N_8413);
or U11889 (N_11889,N_5275,N_6907);
nor U11890 (N_11890,N_6195,N_6838);
nor U11891 (N_11891,N_7039,N_5374);
or U11892 (N_11892,N_8548,N_9643);
or U11893 (N_11893,N_5436,N_9931);
and U11894 (N_11894,N_9679,N_5220);
and U11895 (N_11895,N_9404,N_9723);
nand U11896 (N_11896,N_7646,N_7053);
nor U11897 (N_11897,N_5151,N_6543);
nand U11898 (N_11898,N_9818,N_6728);
nor U11899 (N_11899,N_5244,N_9457);
or U11900 (N_11900,N_5990,N_5966);
and U11901 (N_11901,N_5333,N_8381);
nor U11902 (N_11902,N_6077,N_8261);
and U11903 (N_11903,N_8891,N_9403);
nand U11904 (N_11904,N_8662,N_8435);
and U11905 (N_11905,N_5614,N_9487);
or U11906 (N_11906,N_8369,N_9076);
nand U11907 (N_11907,N_5877,N_7670);
nor U11908 (N_11908,N_6353,N_9164);
nand U11909 (N_11909,N_7291,N_9545);
nand U11910 (N_11910,N_7808,N_5273);
and U11911 (N_11911,N_5168,N_5972);
nor U11912 (N_11912,N_7669,N_9988);
nor U11913 (N_11913,N_5113,N_9912);
nor U11914 (N_11914,N_6280,N_9706);
nor U11915 (N_11915,N_6363,N_9078);
nor U11916 (N_11916,N_8906,N_7454);
nor U11917 (N_11917,N_7793,N_5295);
or U11918 (N_11918,N_6605,N_6879);
or U11919 (N_11919,N_6188,N_5055);
and U11920 (N_11920,N_6396,N_8264);
or U11921 (N_11921,N_5545,N_9892);
and U11922 (N_11922,N_9095,N_7580);
nor U11923 (N_11923,N_7837,N_8800);
nor U11924 (N_11924,N_7628,N_9705);
nand U11925 (N_11925,N_7961,N_7183);
or U11926 (N_11926,N_9963,N_7832);
nand U11927 (N_11927,N_7645,N_5673);
nor U11928 (N_11928,N_9070,N_5393);
or U11929 (N_11929,N_8849,N_9799);
nor U11930 (N_11930,N_5027,N_8033);
or U11931 (N_11931,N_5096,N_5103);
and U11932 (N_11932,N_6761,N_8998);
nor U11933 (N_11933,N_8238,N_5025);
nor U11934 (N_11934,N_6226,N_6493);
or U11935 (N_11935,N_7109,N_7189);
and U11936 (N_11936,N_7286,N_9134);
nor U11937 (N_11937,N_9852,N_9792);
nand U11938 (N_11938,N_5465,N_7922);
nor U11939 (N_11939,N_8051,N_5688);
nor U11940 (N_11940,N_9958,N_5552);
and U11941 (N_11941,N_5700,N_5179);
nor U11942 (N_11942,N_8521,N_8902);
or U11943 (N_11943,N_6925,N_7005);
nand U11944 (N_11944,N_7644,N_6378);
or U11945 (N_11945,N_8519,N_8542);
nand U11946 (N_11946,N_5369,N_7912);
or U11947 (N_11947,N_6868,N_8839);
or U11948 (N_11948,N_7500,N_5140);
and U11949 (N_11949,N_6923,N_7001);
or U11950 (N_11950,N_7513,N_6488);
nor U11951 (N_11951,N_8606,N_5557);
nand U11952 (N_11952,N_5181,N_8877);
nor U11953 (N_11953,N_7268,N_5013);
or U11954 (N_11954,N_7729,N_5629);
xor U11955 (N_11955,N_6829,N_9516);
nand U11956 (N_11956,N_5963,N_8853);
nand U11957 (N_11957,N_9791,N_8969);
and U11958 (N_11958,N_9661,N_5589);
nor U11959 (N_11959,N_8098,N_6701);
or U11960 (N_11960,N_9732,N_8938);
and U11961 (N_11961,N_9544,N_9261);
or U11962 (N_11962,N_8626,N_5701);
and U11963 (N_11963,N_7471,N_9205);
or U11964 (N_11964,N_6001,N_6599);
and U11965 (N_11965,N_9141,N_9846);
xor U11966 (N_11966,N_5942,N_8125);
nor U11967 (N_11967,N_9168,N_6758);
and U11968 (N_11968,N_9616,N_5813);
or U11969 (N_11969,N_6205,N_8234);
nor U11970 (N_11970,N_9055,N_9442);
or U11971 (N_11971,N_9042,N_6213);
nand U11972 (N_11972,N_7479,N_7800);
and U11973 (N_11973,N_6042,N_5183);
or U11974 (N_11974,N_5581,N_5000);
or U11975 (N_11975,N_9520,N_6845);
nand U11976 (N_11976,N_6045,N_9198);
nor U11977 (N_11977,N_8464,N_6815);
nand U11978 (N_11978,N_9807,N_7828);
nand U11979 (N_11979,N_7294,N_8954);
nand U11980 (N_11980,N_5114,N_8872);
nand U11981 (N_11981,N_6526,N_7596);
nor U11982 (N_11982,N_8172,N_6894);
xor U11983 (N_11983,N_7887,N_9877);
or U11984 (N_11984,N_5756,N_9369);
nor U11985 (N_11985,N_9147,N_6146);
xor U11986 (N_11986,N_5758,N_9507);
and U11987 (N_11987,N_5560,N_6655);
nor U11988 (N_11988,N_8291,N_6520);
nor U11989 (N_11989,N_7927,N_6524);
nor U11990 (N_11990,N_6276,N_7026);
and U11991 (N_11991,N_8497,N_5642);
nand U11992 (N_11992,N_8785,N_5060);
and U11993 (N_11993,N_9049,N_6368);
nand U11994 (N_11994,N_6096,N_7378);
or U11995 (N_11995,N_5131,N_6848);
nor U11996 (N_11996,N_5712,N_8126);
and U11997 (N_11997,N_8217,N_9721);
nor U11998 (N_11998,N_9045,N_8349);
and U11999 (N_11999,N_7694,N_9553);
and U12000 (N_12000,N_6046,N_8336);
nor U12001 (N_12001,N_9274,N_5420);
nand U12002 (N_12002,N_6304,N_7607);
nor U12003 (N_12003,N_8942,N_9756);
and U12004 (N_12004,N_5534,N_7478);
nand U12005 (N_12005,N_5371,N_8501);
or U12006 (N_12006,N_8979,N_6031);
and U12007 (N_12007,N_8010,N_5620);
nand U12008 (N_12008,N_6416,N_9539);
nor U12009 (N_12009,N_8574,N_5487);
nor U12010 (N_12010,N_7516,N_6167);
nor U12011 (N_12011,N_7548,N_8240);
and U12012 (N_12012,N_9798,N_8930);
xnor U12013 (N_12013,N_6988,N_7604);
nand U12014 (N_12014,N_7696,N_6991);
nor U12015 (N_12015,N_5895,N_9738);
nand U12016 (N_12016,N_7161,N_6054);
nor U12017 (N_12017,N_8192,N_8223);
or U12018 (N_12018,N_9255,N_5358);
and U12019 (N_12019,N_9170,N_8268);
or U12020 (N_12020,N_5213,N_6176);
nor U12021 (N_12021,N_5548,N_8457);
nor U12022 (N_12022,N_5883,N_6271);
nand U12023 (N_12023,N_5523,N_6965);
or U12024 (N_12024,N_6288,N_7258);
nand U12025 (N_12025,N_7138,N_8944);
and U12026 (N_12026,N_6469,N_6601);
and U12027 (N_12027,N_5757,N_6384);
and U12028 (N_12028,N_6755,N_5155);
nand U12029 (N_12029,N_7384,N_9692);
or U12030 (N_12030,N_8247,N_8168);
nor U12031 (N_12031,N_7649,N_5691);
or U12032 (N_12032,N_8827,N_9414);
and U12033 (N_12033,N_7799,N_5166);
or U12034 (N_12034,N_7274,N_6005);
nand U12035 (N_12035,N_9122,N_5791);
or U12036 (N_12036,N_7535,N_6895);
nor U12037 (N_12037,N_8487,N_5946);
or U12038 (N_12038,N_5919,N_9125);
and U12039 (N_12039,N_9531,N_5537);
nor U12040 (N_12040,N_9527,N_8090);
or U12041 (N_12041,N_9235,N_6884);
and U12042 (N_12042,N_6769,N_5349);
or U12043 (N_12043,N_5925,N_6778);
nand U12044 (N_12044,N_7574,N_5100);
or U12045 (N_12045,N_8639,N_9499);
or U12046 (N_12046,N_5681,N_6440);
or U12047 (N_12047,N_6822,N_8001);
nand U12048 (N_12048,N_6684,N_7186);
nand U12049 (N_12049,N_6382,N_8225);
and U12050 (N_12050,N_5828,N_7009);
or U12051 (N_12051,N_7103,N_9041);
nand U12052 (N_12052,N_8114,N_9588);
nand U12053 (N_12053,N_8643,N_6043);
nand U12054 (N_12054,N_9707,N_5165);
xnor U12055 (N_12055,N_6376,N_8475);
nand U12056 (N_12056,N_7241,N_5754);
and U12057 (N_12057,N_9297,N_9301);
and U12058 (N_12058,N_8678,N_8446);
or U12059 (N_12059,N_7908,N_5074);
nor U12060 (N_12060,N_5973,N_5985);
or U12061 (N_12061,N_6517,N_7790);
nor U12062 (N_12062,N_7844,N_5068);
nor U12063 (N_12063,N_9955,N_9064);
or U12064 (N_12064,N_5601,N_5809);
nand U12065 (N_12065,N_8803,N_7562);
nor U12066 (N_12066,N_7115,N_9946);
and U12067 (N_12067,N_8286,N_8156);
nand U12068 (N_12068,N_8491,N_7307);
nor U12069 (N_12069,N_9305,N_9191);
nand U12070 (N_12070,N_8895,N_8460);
and U12071 (N_12071,N_7974,N_9685);
nand U12072 (N_12072,N_9760,N_8655);
and U12073 (N_12073,N_6334,N_7363);
or U12074 (N_12074,N_7466,N_6142);
or U12075 (N_12075,N_7738,N_6007);
and U12076 (N_12076,N_8554,N_5719);
or U12077 (N_12077,N_6354,N_9451);
nor U12078 (N_12078,N_8206,N_8078);
nand U12079 (N_12079,N_8500,N_7193);
nand U12080 (N_12080,N_7503,N_9118);
nand U12081 (N_12081,N_9669,N_8706);
and U12082 (N_12082,N_9178,N_5342);
nor U12083 (N_12083,N_9774,N_8900);
and U12084 (N_12084,N_7257,N_7463);
or U12085 (N_12085,N_6813,N_9157);
and U12086 (N_12086,N_7049,N_6840);
and U12087 (N_12087,N_9744,N_6771);
nand U12088 (N_12088,N_5338,N_7572);
nor U12089 (N_12089,N_6215,N_7391);
nor U12090 (N_12090,N_7099,N_8175);
or U12091 (N_12091,N_8407,N_9386);
nand U12092 (N_12092,N_6059,N_5917);
nand U12093 (N_12093,N_9493,N_9189);
and U12094 (N_12094,N_5321,N_6483);
nand U12095 (N_12095,N_8440,N_7358);
nand U12096 (N_12096,N_6945,N_9833);
and U12097 (N_12097,N_8672,N_5747);
and U12098 (N_12098,N_7303,N_9376);
or U12099 (N_12099,N_8631,N_6078);
nand U12100 (N_12100,N_9734,N_5384);
or U12101 (N_12101,N_9492,N_9300);
and U12102 (N_12102,N_5177,N_6079);
and U12103 (N_12103,N_8659,N_7232);
nor U12104 (N_12104,N_8037,N_6009);
or U12105 (N_12105,N_5107,N_6399);
nor U12106 (N_12106,N_7476,N_7214);
nand U12107 (N_12107,N_8132,N_7631);
nand U12108 (N_12108,N_7865,N_9889);
and U12109 (N_12109,N_7561,N_9342);
xor U12110 (N_12110,N_5656,N_9258);
and U12111 (N_12111,N_6591,N_6362);
nand U12112 (N_12112,N_7942,N_7512);
nand U12113 (N_12113,N_5311,N_6160);
nor U12114 (N_12114,N_6411,N_5667);
or U12115 (N_12115,N_6867,N_8445);
or U12116 (N_12116,N_8812,N_5380);
nor U12117 (N_12117,N_7442,N_7651);
nand U12118 (N_12118,N_9278,N_9021);
nand U12119 (N_12119,N_9085,N_6232);
nand U12120 (N_12120,N_6625,N_9595);
or U12121 (N_12121,N_7904,N_6201);
or U12122 (N_12122,N_7071,N_9069);
nand U12123 (N_12123,N_7588,N_6556);
and U12124 (N_12124,N_7187,N_6298);
and U12125 (N_12125,N_5531,N_6727);
nor U12126 (N_12126,N_6261,N_7611);
nor U12127 (N_12127,N_6255,N_6646);
or U12128 (N_12128,N_8529,N_5482);
or U12129 (N_12129,N_9796,N_8385);
and U12130 (N_12130,N_5668,N_6682);
nor U12131 (N_12131,N_6310,N_8843);
or U12132 (N_12132,N_7734,N_8732);
and U12133 (N_12133,N_5511,N_6501);
nor U12134 (N_12134,N_5008,N_8880);
or U12135 (N_12135,N_5097,N_5014);
nor U12136 (N_12136,N_5927,N_8372);
nor U12137 (N_12137,N_5500,N_8962);
nand U12138 (N_12138,N_5905,N_9962);
nor U12139 (N_12139,N_9957,N_9940);
nand U12140 (N_12140,N_8798,N_6423);
nor U12141 (N_12141,N_5980,N_5994);
nand U12142 (N_12142,N_7941,N_7654);
and U12143 (N_12143,N_6745,N_5466);
and U12144 (N_12144,N_5930,N_9733);
or U12145 (N_12145,N_5529,N_5569);
nand U12146 (N_12146,N_8101,N_7355);
or U12147 (N_12147,N_5694,N_8893);
or U12148 (N_12148,N_8121,N_5464);
nand U12149 (N_12149,N_9896,N_8637);
or U12150 (N_12150,N_5425,N_7673);
and U12151 (N_12151,N_5091,N_8161);
nand U12152 (N_12152,N_8462,N_6902);
nand U12153 (N_12153,N_7688,N_6186);
and U12154 (N_12154,N_8647,N_5780);
nor U12155 (N_12155,N_8509,N_9419);
or U12156 (N_12156,N_6892,N_6983);
nand U12157 (N_12157,N_8513,N_8113);
nand U12158 (N_12158,N_6419,N_8195);
nand U12159 (N_12159,N_9930,N_6221);
or U12160 (N_12160,N_6656,N_5040);
and U12161 (N_12161,N_5259,N_9144);
nand U12162 (N_12162,N_7261,N_5763);
and U12163 (N_12163,N_6527,N_7414);
nor U12164 (N_12164,N_9484,N_5816);
nand U12165 (N_12165,N_9716,N_7526);
and U12166 (N_12166,N_9182,N_8937);
and U12167 (N_12167,N_5363,N_8718);
nand U12168 (N_12168,N_5664,N_9446);
nand U12169 (N_12169,N_5836,N_5805);
nor U12170 (N_12170,N_9528,N_9650);
or U12171 (N_12171,N_9281,N_8628);
nand U12172 (N_12172,N_8553,N_5236);
and U12173 (N_12173,N_7340,N_8154);
or U12174 (N_12174,N_5774,N_7491);
or U12175 (N_12175,N_6660,N_5052);
nand U12176 (N_12176,N_8523,N_5484);
nand U12177 (N_12177,N_9648,N_5348);
or U12178 (N_12178,N_6265,N_8243);
and U12179 (N_12179,N_7499,N_5662);
nor U12180 (N_12180,N_7361,N_9708);
nand U12181 (N_12181,N_7458,N_6594);
nor U12182 (N_12182,N_5649,N_5035);
or U12183 (N_12183,N_9969,N_6578);
nor U12184 (N_12184,N_9632,N_7559);
nor U12185 (N_12185,N_7300,N_9769);
nand U12186 (N_12186,N_5203,N_6159);
nand U12187 (N_12187,N_5749,N_6858);
or U12188 (N_12188,N_6702,N_8636);
nand U12189 (N_12189,N_8220,N_8107);
nor U12190 (N_12190,N_8572,N_7529);
and U12191 (N_12191,N_7716,N_6602);
nor U12192 (N_12192,N_6592,N_5411);
or U12193 (N_12193,N_5725,N_8199);
nor U12194 (N_12194,N_5679,N_7664);
or U12195 (N_12195,N_6212,N_9214);
nand U12196 (N_12196,N_5945,N_8681);
or U12197 (N_12197,N_7239,N_9919);
nand U12198 (N_12198,N_9081,N_9591);
nand U12199 (N_12199,N_6859,N_8738);
nand U12200 (N_12200,N_8455,N_6570);
nor U12201 (N_12201,N_6714,N_9558);
and U12202 (N_12202,N_8761,N_6185);
and U12203 (N_12203,N_5033,N_8988);
nor U12204 (N_12204,N_8026,N_9725);
nor U12205 (N_12205,N_7742,N_8380);
or U12206 (N_12206,N_7543,N_8214);
nand U12207 (N_12207,N_8456,N_8039);
nand U12208 (N_12208,N_7643,N_6140);
and U12209 (N_12209,N_7236,N_5197);
or U12210 (N_12210,N_7964,N_9978);
nand U12211 (N_12211,N_9266,N_9879);
nand U12212 (N_12212,N_9291,N_9666);
or U12213 (N_12213,N_8285,N_6268);
nor U12214 (N_12214,N_6504,N_8602);
or U12215 (N_12215,N_5904,N_5267);
or U12216 (N_12216,N_5407,N_7062);
and U12217 (N_12217,N_7994,N_5123);
and U12218 (N_12218,N_6774,N_8269);
nand U12219 (N_12219,N_7367,N_7846);
nand U12220 (N_12220,N_8931,N_5216);
or U12221 (N_12221,N_9662,N_6987);
and U12222 (N_12222,N_6153,N_8855);
nor U12223 (N_12223,N_8688,N_8822);
nand U12224 (N_12224,N_9152,N_6562);
or U12225 (N_12225,N_8109,N_5570);
nor U12226 (N_12226,N_8333,N_8951);
nand U12227 (N_12227,N_5089,N_6344);
or U12228 (N_12228,N_5360,N_9043);
nand U12229 (N_12229,N_5298,N_6135);
nand U12230 (N_12230,N_8093,N_7124);
nor U12231 (N_12231,N_5385,N_6586);
nand U12232 (N_12232,N_9108,N_5099);
and U12233 (N_12233,N_7276,N_7840);
or U12234 (N_12234,N_6560,N_8202);
nand U12235 (N_12235,N_8560,N_6465);
and U12236 (N_12236,N_7376,N_5542);
nor U12237 (N_12237,N_9574,N_8571);
or U12238 (N_12238,N_9784,N_5781);
nor U12239 (N_12239,N_7100,N_9802);
or U12240 (N_12240,N_8693,N_8745);
nor U12241 (N_12241,N_7425,N_7177);
xor U12242 (N_12242,N_5824,N_7642);
and U12243 (N_12243,N_9143,N_5833);
nand U12244 (N_12244,N_9904,N_8584);
nand U12245 (N_12245,N_8315,N_8621);
or U12246 (N_12246,N_5274,N_9869);
nand U12247 (N_12247,N_9226,N_5900);
or U12248 (N_12248,N_6375,N_7430);
nor U12249 (N_12249,N_5835,N_5974);
nand U12250 (N_12250,N_8958,N_8525);
or U12251 (N_12251,N_6903,N_6008);
or U12252 (N_12252,N_9614,N_7902);
nor U12253 (N_12253,N_6249,N_7040);
nor U12254 (N_12254,N_5920,N_9849);
nor U12255 (N_12255,N_6699,N_6844);
nand U12256 (N_12256,N_5029,N_8620);
nor U12257 (N_12257,N_7393,N_6600);
or U12258 (N_12258,N_6208,N_7102);
or U12259 (N_12259,N_5293,N_5062);
or U12260 (N_12260,N_6666,N_6933);
and U12261 (N_12261,N_9977,N_5315);
nand U12262 (N_12262,N_8982,N_8787);
or U12263 (N_12263,N_8099,N_9980);
or U12264 (N_12264,N_8802,N_9826);
nand U12265 (N_12265,N_8711,N_8977);
or U12266 (N_12266,N_5230,N_6222);
or U12267 (N_12267,N_7709,N_6311);
nor U12268 (N_12268,N_6990,N_6724);
nor U12269 (N_12269,N_5767,N_9153);
and U12270 (N_12270,N_7554,N_6870);
nor U12271 (N_12271,N_8948,N_6004);
nor U12272 (N_12272,N_8623,N_7936);
nor U12273 (N_12273,N_6931,N_5543);
or U12274 (N_12274,N_7565,N_7617);
and U12275 (N_12275,N_9914,N_8593);
and U12276 (N_12276,N_9908,N_5001);
or U12277 (N_12277,N_5171,N_8680);
or U12278 (N_12278,N_7380,N_9173);
nand U12279 (N_12279,N_6203,N_6703);
or U12280 (N_12280,N_5020,N_7877);
and U12281 (N_12281,N_5617,N_6060);
nor U12282 (N_12282,N_7022,N_9338);
and U12283 (N_12283,N_7914,N_7417);
nand U12284 (N_12284,N_9362,N_6650);
nor U12285 (N_12285,N_7446,N_6118);
or U12286 (N_12286,N_9813,N_8566);
or U12287 (N_12287,N_8786,N_5088);
nand U12288 (N_12288,N_8122,N_7920);
and U12289 (N_12289,N_5057,N_6969);
nand U12290 (N_12290,N_7220,N_9728);
and U12291 (N_12291,N_7563,N_5647);
and U12292 (N_12292,N_6644,N_8190);
nand U12293 (N_12293,N_7838,N_9053);
and U12294 (N_12294,N_8005,N_5129);
or U12295 (N_12295,N_6883,N_7848);
nand U12296 (N_12296,N_6331,N_7234);
and U12297 (N_12297,N_6145,N_7746);
nor U12298 (N_12298,N_6654,N_8360);
nor U12299 (N_12299,N_6999,N_5219);
and U12300 (N_12300,N_9781,N_7339);
nand U12301 (N_12301,N_8755,N_6808);
and U12302 (N_12302,N_8520,N_9997);
and U12303 (N_12303,N_5002,N_8763);
nand U12304 (N_12304,N_9761,N_5435);
nand U12305 (N_12305,N_6934,N_5105);
nand U12306 (N_12306,N_7366,N_6109);
nand U12307 (N_12307,N_9687,N_8480);
nor U12308 (N_12308,N_5707,N_8728);
nor U12309 (N_12309,N_7089,N_6010);
or U12310 (N_12310,N_5825,N_6972);
nor U12311 (N_12311,N_9433,N_8604);
nand U12312 (N_12312,N_9292,N_5483);
and U12313 (N_12313,N_6782,N_9084);
nand U12314 (N_12314,N_9295,N_8726);
nand U12315 (N_12315,N_6876,N_7986);
nand U12316 (N_12316,N_9546,N_9190);
or U12317 (N_12317,N_6258,N_7289);
or U12318 (N_12318,N_8912,N_9557);
and U12319 (N_12319,N_7420,N_8714);
and U12320 (N_12320,N_9390,N_8967);
or U12321 (N_12321,N_8599,N_7741);
nor U12322 (N_12322,N_7754,N_5037);
and U12323 (N_12323,N_8709,N_7743);
and U12324 (N_12324,N_5610,N_6582);
nor U12325 (N_12325,N_8297,N_6366);
nand U12326 (N_12326,N_8870,N_7290);
nor U12327 (N_12327,N_7984,N_9987);
or U12328 (N_12328,N_7341,N_6740);
and U12329 (N_12329,N_6826,N_6633);
and U12330 (N_12330,N_5924,N_8359);
nand U12331 (N_12331,N_5424,N_6661);
nand U12332 (N_12332,N_6324,N_8874);
or U12333 (N_12333,N_7637,N_9497);
nand U12334 (N_12334,N_7889,N_8776);
or U12335 (N_12335,N_5528,N_8274);
nand U12336 (N_12336,N_5438,N_7797);
or U12337 (N_12337,N_9524,N_9753);
nor U12338 (N_12338,N_6123,N_7774);
or U12339 (N_12339,N_9353,N_9307);
or U12340 (N_12340,N_9871,N_6328);
nor U12341 (N_12341,N_5916,N_6020);
or U12342 (N_12342,N_6697,N_9657);
nand U12343 (N_12343,N_9693,N_6309);
nand U12344 (N_12344,N_6747,N_7436);
nand U12345 (N_12345,N_7896,N_8088);
or U12346 (N_12346,N_5108,N_7204);
or U12347 (N_12347,N_8421,N_7570);
and U12348 (N_12348,N_6218,N_8499);
and U12349 (N_12349,N_6233,N_7852);
nor U12350 (N_12350,N_5788,N_5175);
or U12351 (N_12351,N_6764,N_8367);
or U12352 (N_12352,N_8412,N_7092);
and U12353 (N_12353,N_7320,N_6040);
xor U12354 (N_12354,N_8299,N_8793);
nand U12355 (N_12355,N_9029,N_9465);
nor U12356 (N_12356,N_7460,N_5368);
or U12357 (N_12357,N_5307,N_8669);
nor U12358 (N_12358,N_8362,N_7926);
nor U12359 (N_12359,N_9642,N_9437);
and U12360 (N_12360,N_6749,N_9903);
nand U12361 (N_12361,N_9714,N_6510);
or U12362 (N_12362,N_9793,N_5878);
or U12363 (N_12363,N_7113,N_9569);
nand U12364 (N_12364,N_6954,N_6706);
nor U12365 (N_12365,N_6223,N_9770);
nand U12366 (N_12366,N_7282,N_8365);
nand U12367 (N_12367,N_8146,N_8907);
xor U12368 (N_12368,N_8133,N_5240);
or U12369 (N_12369,N_7243,N_6715);
and U12370 (N_12370,N_8024,N_6182);
and U12371 (N_12371,N_6120,N_9251);
and U12372 (N_12372,N_8404,N_9279);
and U12373 (N_12373,N_9860,N_9696);
nor U12374 (N_12374,N_7569,N_6926);
and U12375 (N_12375,N_5070,N_7087);
nand U12376 (N_12376,N_5801,N_8119);
nand U12377 (N_12377,N_8638,N_5807);
nor U12378 (N_12378,N_7111,N_5911);
and U12379 (N_12379,N_9918,N_7342);
nand U12380 (N_12380,N_8731,N_5839);
and U12381 (N_12381,N_6318,N_5867);
or U12382 (N_12382,N_5593,N_5858);
or U12383 (N_12383,N_7614,N_8108);
nor U12384 (N_12384,N_8350,N_7375);
and U12385 (N_12385,N_8197,N_9285);
nor U12386 (N_12386,N_5285,N_8890);
nand U12387 (N_12387,N_5458,N_6491);
nand U12388 (N_12388,N_7965,N_9533);
or U12389 (N_12389,N_5461,N_5713);
and U12390 (N_12390,N_5495,N_9184);
nor U12391 (N_12391,N_5199,N_6386);
and U12392 (N_12392,N_9374,N_6236);
nor U12393 (N_12393,N_6329,N_6247);
or U12394 (N_12394,N_7207,N_6837);
and U12395 (N_12395,N_6470,N_9399);
and U12396 (N_12396,N_5124,N_6433);
and U12397 (N_12397,N_8317,N_7429);
nor U12398 (N_12398,N_7469,N_7495);
and U12399 (N_12399,N_9639,N_8429);
and U12400 (N_12400,N_5150,N_5264);
and U12401 (N_12401,N_8689,N_8403);
nor U12402 (N_12402,N_9352,N_5680);
or U12403 (N_12403,N_5246,N_7409);
or U12404 (N_12404,N_7121,N_7408);
or U12405 (N_12405,N_6361,N_8729);
xor U12406 (N_12406,N_7931,N_5235);
or U12407 (N_12407,N_7486,N_6814);
nor U12408 (N_12408,N_5009,N_7875);
and U12409 (N_12409,N_8022,N_9647);
or U12410 (N_12410,N_7689,N_6434);
or U12411 (N_12411,N_5550,N_6306);
nor U12412 (N_12412,N_6579,N_9560);
or U12413 (N_12413,N_5265,N_6364);
or U12414 (N_12414,N_9197,N_9568);
and U12415 (N_12415,N_7299,N_6383);
nand U12416 (N_12416,N_7242,N_9653);
nand U12417 (N_12417,N_9315,N_7357);
and U12418 (N_12418,N_7428,N_6941);
or U12419 (N_12419,N_7540,N_5208);
nand U12420 (N_12420,N_5118,N_9488);
and U12421 (N_12421,N_5894,N_5314);
nand U12422 (N_12422,N_8469,N_9758);
or U12423 (N_12423,N_5283,N_7663);
nand U12424 (N_12424,N_6743,N_5191);
and U12425 (N_12425,N_7063,N_8399);
or U12426 (N_12426,N_7751,N_9655);
or U12427 (N_12427,N_9165,N_9766);
or U12428 (N_12428,N_5775,N_6257);
nand U12429 (N_12429,N_5627,N_6052);
nor U12430 (N_12430,N_5918,N_6705);
nand U12431 (N_12431,N_6485,N_7597);
nand U12432 (N_12432,N_8517,N_7047);
or U12433 (N_12433,N_5561,N_5602);
or U12434 (N_12434,N_9460,N_5022);
or U12435 (N_12435,N_6139,N_5361);
nand U12436 (N_12436,N_6767,N_8940);
or U12437 (N_12437,N_6454,N_6871);
nand U12438 (N_12438,N_9277,N_6150);
or U12439 (N_12439,N_6169,N_6330);
nand U12440 (N_12440,N_6477,N_7015);
and U12441 (N_12441,N_8677,N_8635);
xnor U12442 (N_12442,N_9303,N_7857);
or U12443 (N_12443,N_8442,N_8461);
or U12444 (N_12444,N_8653,N_6397);
and U12445 (N_12445,N_6788,N_5951);
nor U12446 (N_12446,N_5720,N_8432);
nand U12447 (N_12447,N_5855,N_8913);
and U12448 (N_12448,N_6225,N_7639);
nor U12449 (N_12449,N_8904,N_5316);
and U12450 (N_12450,N_8112,N_5708);
or U12451 (N_12451,N_9109,N_6636);
nor U12452 (N_12452,N_8683,N_5536);
and U12453 (N_12453,N_5327,N_6950);
nor U12454 (N_12454,N_7874,N_5330);
and U12455 (N_12455,N_7620,N_6955);
nor U12456 (N_12456,N_6068,N_5310);
nand U12457 (N_12457,N_6521,N_6294);
and U12458 (N_12458,N_5260,N_8997);
nor U12459 (N_12459,N_7031,N_9483);
nor U12460 (N_12460,N_7297,N_8950);
nand U12461 (N_12461,N_8748,N_9782);
nand U12462 (N_12462,N_6240,N_7166);
nor U12463 (N_12463,N_9972,N_8665);
or U12464 (N_12464,N_8178,N_7960);
and U12465 (N_12465,N_9252,N_9688);
and U12466 (N_12466,N_6075,N_6659);
and U12467 (N_12467,N_6239,N_9371);
nor U12468 (N_12468,N_6836,N_6372);
and U12469 (N_12469,N_6275,N_6511);
nor U12470 (N_12470,N_6738,N_7136);
and U12471 (N_12471,N_8117,N_7041);
and U12472 (N_12472,N_8828,N_8720);
xnor U12473 (N_12473,N_9667,N_9240);
and U12474 (N_12474,N_5087,N_6081);
nor U12475 (N_12475,N_5776,N_6768);
or U12476 (N_12476,N_8743,N_8864);
nand U12477 (N_12477,N_7538,N_5470);
or U12478 (N_12478,N_9138,N_5024);
nand U12479 (N_12479,N_6390,N_8319);
nand U12480 (N_12480,N_5806,N_7581);
nor U12481 (N_12481,N_5451,N_6017);
or U12482 (N_12482,N_6681,N_9961);
nand U12483 (N_12483,N_8123,N_7873);
nor U12484 (N_12484,N_8494,N_9312);
and U12485 (N_12485,N_6452,N_6943);
nand U12486 (N_12486,N_9028,N_7069);
nand U12487 (N_12487,N_8540,N_7174);
and U12488 (N_12488,N_6475,N_8614);
nand U12489 (N_12489,N_6023,N_6757);
or U12490 (N_12490,N_6930,N_7360);
nand U12491 (N_12491,N_7244,N_5186);
nor U12492 (N_12492,N_7251,N_6554);
nor U12493 (N_12493,N_9175,N_8568);
or U12494 (N_12494,N_9510,N_7821);
nor U12495 (N_12495,N_8355,N_9156);
nand U12496 (N_12496,N_9370,N_6816);
and U12497 (N_12497,N_5051,N_5319);
nand U12498 (N_12498,N_6064,N_9000);
nand U12499 (N_12499,N_9884,N_5493);
or U12500 (N_12500,N_6872,N_7638);
nand U12501 (N_12501,N_8593,N_6400);
nand U12502 (N_12502,N_7834,N_7324);
nor U12503 (N_12503,N_9892,N_8319);
or U12504 (N_12504,N_5218,N_7791);
nor U12505 (N_12505,N_5817,N_8162);
xnor U12506 (N_12506,N_9885,N_8546);
nor U12507 (N_12507,N_8496,N_6434);
and U12508 (N_12508,N_5216,N_6151);
or U12509 (N_12509,N_9414,N_5958);
nand U12510 (N_12510,N_5404,N_5646);
nand U12511 (N_12511,N_9739,N_8913);
and U12512 (N_12512,N_7839,N_6729);
nand U12513 (N_12513,N_9938,N_9189);
nand U12514 (N_12514,N_6798,N_7789);
and U12515 (N_12515,N_9194,N_7892);
and U12516 (N_12516,N_9047,N_9454);
or U12517 (N_12517,N_8193,N_9611);
nor U12518 (N_12518,N_6532,N_7170);
or U12519 (N_12519,N_7169,N_7807);
nand U12520 (N_12520,N_7484,N_5016);
and U12521 (N_12521,N_8835,N_8845);
and U12522 (N_12522,N_5629,N_5170);
xnor U12523 (N_12523,N_9812,N_7575);
and U12524 (N_12524,N_8398,N_5084);
and U12525 (N_12525,N_8824,N_7398);
nor U12526 (N_12526,N_9941,N_8802);
nor U12527 (N_12527,N_8037,N_7560);
and U12528 (N_12528,N_9842,N_5557);
nand U12529 (N_12529,N_5975,N_7631);
nor U12530 (N_12530,N_5248,N_6350);
nand U12531 (N_12531,N_8970,N_8362);
nor U12532 (N_12532,N_7963,N_9259);
and U12533 (N_12533,N_7673,N_9166);
and U12534 (N_12534,N_6235,N_6354);
and U12535 (N_12535,N_5252,N_6327);
nor U12536 (N_12536,N_8159,N_6338);
nand U12537 (N_12537,N_6930,N_7135);
nand U12538 (N_12538,N_6545,N_5042);
or U12539 (N_12539,N_8857,N_7858);
nor U12540 (N_12540,N_8959,N_6966);
nor U12541 (N_12541,N_9263,N_6708);
nor U12542 (N_12542,N_5266,N_7587);
nor U12543 (N_12543,N_9584,N_7167);
nand U12544 (N_12544,N_7302,N_7291);
nand U12545 (N_12545,N_9651,N_8067);
or U12546 (N_12546,N_9222,N_7596);
or U12547 (N_12547,N_6999,N_6751);
nand U12548 (N_12548,N_6230,N_6525);
xor U12549 (N_12549,N_8915,N_7057);
or U12550 (N_12550,N_8709,N_7739);
nor U12551 (N_12551,N_9798,N_9600);
and U12552 (N_12552,N_9352,N_8912);
nor U12553 (N_12553,N_5861,N_6160);
nand U12554 (N_12554,N_5351,N_5808);
and U12555 (N_12555,N_9618,N_9965);
or U12556 (N_12556,N_9931,N_9371);
nand U12557 (N_12557,N_5555,N_6510);
and U12558 (N_12558,N_6160,N_7214);
nand U12559 (N_12559,N_6739,N_9245);
nor U12560 (N_12560,N_6722,N_7899);
nor U12561 (N_12561,N_5505,N_9872);
or U12562 (N_12562,N_9798,N_7451);
and U12563 (N_12563,N_5524,N_9023);
and U12564 (N_12564,N_7673,N_9705);
xor U12565 (N_12565,N_9389,N_6662);
or U12566 (N_12566,N_9311,N_7823);
and U12567 (N_12567,N_6346,N_5133);
nand U12568 (N_12568,N_7306,N_9850);
or U12569 (N_12569,N_8651,N_5451);
or U12570 (N_12570,N_7170,N_9794);
nand U12571 (N_12571,N_9528,N_5673);
nand U12572 (N_12572,N_6737,N_5346);
or U12573 (N_12573,N_6538,N_9682);
or U12574 (N_12574,N_8899,N_5163);
and U12575 (N_12575,N_5859,N_6045);
and U12576 (N_12576,N_8200,N_6537);
nand U12577 (N_12577,N_5021,N_7304);
nor U12578 (N_12578,N_5192,N_7165);
and U12579 (N_12579,N_9552,N_6333);
nor U12580 (N_12580,N_8365,N_9964);
nand U12581 (N_12581,N_9394,N_8285);
nand U12582 (N_12582,N_5853,N_8882);
nand U12583 (N_12583,N_6335,N_9680);
nand U12584 (N_12584,N_5666,N_7802);
and U12585 (N_12585,N_6404,N_6500);
and U12586 (N_12586,N_7999,N_9368);
or U12587 (N_12587,N_8755,N_8456);
or U12588 (N_12588,N_9584,N_9572);
nor U12589 (N_12589,N_7229,N_8619);
nand U12590 (N_12590,N_5902,N_5813);
nand U12591 (N_12591,N_8905,N_7280);
nand U12592 (N_12592,N_5864,N_5721);
nand U12593 (N_12593,N_9550,N_7583);
or U12594 (N_12594,N_6990,N_8577);
xor U12595 (N_12595,N_9533,N_8179);
nand U12596 (N_12596,N_5909,N_8039);
and U12597 (N_12597,N_8730,N_6608);
or U12598 (N_12598,N_8740,N_6074);
and U12599 (N_12599,N_9004,N_9645);
and U12600 (N_12600,N_8851,N_6151);
nand U12601 (N_12601,N_6492,N_9102);
nand U12602 (N_12602,N_6911,N_9472);
nand U12603 (N_12603,N_7593,N_5540);
and U12604 (N_12604,N_9277,N_9556);
or U12605 (N_12605,N_9502,N_8450);
nand U12606 (N_12606,N_9674,N_7405);
and U12607 (N_12607,N_5142,N_9868);
or U12608 (N_12608,N_9909,N_7193);
and U12609 (N_12609,N_6988,N_7704);
nand U12610 (N_12610,N_6258,N_5316);
or U12611 (N_12611,N_9701,N_6951);
or U12612 (N_12612,N_7357,N_7406);
or U12613 (N_12613,N_6172,N_8249);
nand U12614 (N_12614,N_5139,N_8943);
nor U12615 (N_12615,N_7340,N_5235);
nand U12616 (N_12616,N_7350,N_8050);
nand U12617 (N_12617,N_6998,N_9811);
or U12618 (N_12618,N_5593,N_9355);
and U12619 (N_12619,N_6824,N_5604);
or U12620 (N_12620,N_7267,N_7215);
nor U12621 (N_12621,N_6764,N_6359);
nor U12622 (N_12622,N_7599,N_7247);
or U12623 (N_12623,N_7788,N_6069);
nor U12624 (N_12624,N_5821,N_7331);
and U12625 (N_12625,N_5367,N_5402);
nor U12626 (N_12626,N_5437,N_6492);
or U12627 (N_12627,N_7630,N_9218);
nand U12628 (N_12628,N_6400,N_6938);
nand U12629 (N_12629,N_5309,N_6436);
nand U12630 (N_12630,N_6609,N_6222);
nor U12631 (N_12631,N_5691,N_6861);
nand U12632 (N_12632,N_8146,N_7636);
nand U12633 (N_12633,N_8527,N_8938);
nand U12634 (N_12634,N_5214,N_7672);
nor U12635 (N_12635,N_6512,N_9695);
and U12636 (N_12636,N_9100,N_6918);
nor U12637 (N_12637,N_7844,N_7398);
or U12638 (N_12638,N_5218,N_9012);
and U12639 (N_12639,N_6608,N_5856);
or U12640 (N_12640,N_9981,N_8304);
nand U12641 (N_12641,N_7431,N_8175);
nand U12642 (N_12642,N_6665,N_7387);
nand U12643 (N_12643,N_6575,N_6004);
or U12644 (N_12644,N_7688,N_9055);
or U12645 (N_12645,N_6776,N_5555);
or U12646 (N_12646,N_8631,N_7996);
nor U12647 (N_12647,N_7205,N_7498);
nor U12648 (N_12648,N_9044,N_5971);
nand U12649 (N_12649,N_7054,N_7910);
and U12650 (N_12650,N_7790,N_6558);
nand U12651 (N_12651,N_6858,N_8237);
nor U12652 (N_12652,N_5678,N_7341);
nor U12653 (N_12653,N_8339,N_7922);
xnor U12654 (N_12654,N_5673,N_7174);
nor U12655 (N_12655,N_5488,N_9281);
and U12656 (N_12656,N_6632,N_9782);
nor U12657 (N_12657,N_5540,N_6578);
and U12658 (N_12658,N_7688,N_6733);
nor U12659 (N_12659,N_7026,N_5307);
and U12660 (N_12660,N_9074,N_9535);
or U12661 (N_12661,N_6590,N_9218);
nor U12662 (N_12662,N_5571,N_5121);
nor U12663 (N_12663,N_9354,N_9102);
and U12664 (N_12664,N_6873,N_9512);
or U12665 (N_12665,N_7357,N_8142);
or U12666 (N_12666,N_9170,N_5388);
nand U12667 (N_12667,N_5409,N_6425);
nor U12668 (N_12668,N_9881,N_7823);
nor U12669 (N_12669,N_8291,N_6817);
or U12670 (N_12670,N_5151,N_8824);
nand U12671 (N_12671,N_5209,N_6965);
or U12672 (N_12672,N_9997,N_5599);
nand U12673 (N_12673,N_9142,N_8785);
or U12674 (N_12674,N_5010,N_6897);
or U12675 (N_12675,N_6074,N_5953);
nor U12676 (N_12676,N_8942,N_5748);
nor U12677 (N_12677,N_9752,N_7864);
and U12678 (N_12678,N_7184,N_6646);
nor U12679 (N_12679,N_8070,N_9629);
nor U12680 (N_12680,N_8967,N_6357);
or U12681 (N_12681,N_8560,N_7390);
and U12682 (N_12682,N_8148,N_9043);
nand U12683 (N_12683,N_5852,N_9126);
and U12684 (N_12684,N_9162,N_7184);
or U12685 (N_12685,N_8417,N_8384);
nor U12686 (N_12686,N_8593,N_8772);
nor U12687 (N_12687,N_9242,N_5070);
and U12688 (N_12688,N_5810,N_7623);
or U12689 (N_12689,N_5583,N_9999);
and U12690 (N_12690,N_6666,N_6738);
nor U12691 (N_12691,N_8815,N_6532);
or U12692 (N_12692,N_5664,N_5585);
nor U12693 (N_12693,N_7399,N_6512);
nand U12694 (N_12694,N_6912,N_7901);
nor U12695 (N_12695,N_6249,N_8353);
or U12696 (N_12696,N_6354,N_7394);
and U12697 (N_12697,N_5082,N_7846);
nand U12698 (N_12698,N_7818,N_7883);
nand U12699 (N_12699,N_5631,N_5847);
or U12700 (N_12700,N_5147,N_7680);
nand U12701 (N_12701,N_8945,N_7678);
or U12702 (N_12702,N_6225,N_6875);
and U12703 (N_12703,N_7926,N_6742);
and U12704 (N_12704,N_6453,N_6185);
and U12705 (N_12705,N_9362,N_8374);
and U12706 (N_12706,N_9277,N_9219);
or U12707 (N_12707,N_7941,N_9713);
nand U12708 (N_12708,N_7519,N_6539);
nor U12709 (N_12709,N_5556,N_8322);
nor U12710 (N_12710,N_8963,N_8142);
nor U12711 (N_12711,N_8205,N_7370);
nand U12712 (N_12712,N_8226,N_9613);
or U12713 (N_12713,N_5841,N_9460);
or U12714 (N_12714,N_7583,N_6782);
nor U12715 (N_12715,N_8809,N_7813);
nor U12716 (N_12716,N_8574,N_5561);
nand U12717 (N_12717,N_5818,N_9729);
nand U12718 (N_12718,N_6939,N_5244);
and U12719 (N_12719,N_5934,N_8688);
nor U12720 (N_12720,N_8030,N_9866);
or U12721 (N_12721,N_5422,N_9430);
and U12722 (N_12722,N_9938,N_6090);
nor U12723 (N_12723,N_7170,N_7560);
nor U12724 (N_12724,N_7000,N_9978);
and U12725 (N_12725,N_8732,N_5109);
and U12726 (N_12726,N_6682,N_6090);
nand U12727 (N_12727,N_6595,N_9765);
nor U12728 (N_12728,N_7252,N_8833);
nor U12729 (N_12729,N_7568,N_7233);
nor U12730 (N_12730,N_7239,N_5311);
or U12731 (N_12731,N_5625,N_8178);
nand U12732 (N_12732,N_8464,N_6860);
nor U12733 (N_12733,N_8650,N_8842);
nand U12734 (N_12734,N_9871,N_6315);
and U12735 (N_12735,N_5772,N_8660);
nand U12736 (N_12736,N_9851,N_7262);
and U12737 (N_12737,N_6821,N_5435);
nor U12738 (N_12738,N_6460,N_9598);
nor U12739 (N_12739,N_7387,N_8334);
nor U12740 (N_12740,N_8101,N_9149);
nor U12741 (N_12741,N_5561,N_9366);
or U12742 (N_12742,N_7870,N_8364);
or U12743 (N_12743,N_6952,N_6196);
or U12744 (N_12744,N_7542,N_9940);
nor U12745 (N_12745,N_5144,N_6068);
nand U12746 (N_12746,N_9866,N_7012);
nor U12747 (N_12747,N_5887,N_8449);
nor U12748 (N_12748,N_9736,N_6161);
and U12749 (N_12749,N_6038,N_6640);
or U12750 (N_12750,N_5154,N_9086);
and U12751 (N_12751,N_8276,N_7754);
or U12752 (N_12752,N_9954,N_6876);
and U12753 (N_12753,N_7427,N_8333);
or U12754 (N_12754,N_6512,N_5697);
and U12755 (N_12755,N_7974,N_6789);
and U12756 (N_12756,N_6735,N_8548);
or U12757 (N_12757,N_9254,N_6724);
or U12758 (N_12758,N_6058,N_9752);
and U12759 (N_12759,N_8414,N_6980);
or U12760 (N_12760,N_6516,N_9728);
and U12761 (N_12761,N_5480,N_5810);
or U12762 (N_12762,N_5676,N_8893);
or U12763 (N_12763,N_6483,N_7041);
or U12764 (N_12764,N_7764,N_9283);
xor U12765 (N_12765,N_6592,N_8249);
nor U12766 (N_12766,N_7140,N_7234);
and U12767 (N_12767,N_7538,N_8148);
nor U12768 (N_12768,N_6055,N_9473);
nand U12769 (N_12769,N_9528,N_9095);
nand U12770 (N_12770,N_9802,N_9237);
or U12771 (N_12771,N_5565,N_9122);
or U12772 (N_12772,N_5793,N_9578);
nor U12773 (N_12773,N_9380,N_5170);
nand U12774 (N_12774,N_8883,N_9685);
nor U12775 (N_12775,N_5821,N_5317);
nand U12776 (N_12776,N_9513,N_8786);
or U12777 (N_12777,N_7925,N_7440);
or U12778 (N_12778,N_5338,N_9497);
nor U12779 (N_12779,N_9112,N_7165);
and U12780 (N_12780,N_8099,N_6278);
nand U12781 (N_12781,N_6482,N_8987);
nor U12782 (N_12782,N_9624,N_6850);
or U12783 (N_12783,N_5637,N_7392);
and U12784 (N_12784,N_5826,N_5126);
xnor U12785 (N_12785,N_7245,N_5471);
or U12786 (N_12786,N_6447,N_6831);
and U12787 (N_12787,N_9771,N_9548);
or U12788 (N_12788,N_7699,N_7100);
nand U12789 (N_12789,N_7997,N_5373);
nor U12790 (N_12790,N_7111,N_9368);
or U12791 (N_12791,N_9005,N_6179);
xnor U12792 (N_12792,N_7211,N_6577);
and U12793 (N_12793,N_9575,N_7099);
or U12794 (N_12794,N_9806,N_5796);
and U12795 (N_12795,N_9503,N_6569);
and U12796 (N_12796,N_9008,N_9928);
or U12797 (N_12797,N_8806,N_5891);
nand U12798 (N_12798,N_7775,N_8552);
and U12799 (N_12799,N_5260,N_8358);
and U12800 (N_12800,N_9638,N_8325);
nor U12801 (N_12801,N_6003,N_6368);
or U12802 (N_12802,N_5108,N_8745);
or U12803 (N_12803,N_7309,N_8158);
and U12804 (N_12804,N_7900,N_7746);
and U12805 (N_12805,N_6468,N_8066);
nand U12806 (N_12806,N_9052,N_6656);
nor U12807 (N_12807,N_8378,N_6941);
and U12808 (N_12808,N_8436,N_8828);
or U12809 (N_12809,N_9529,N_5632);
nor U12810 (N_12810,N_5624,N_7013);
nand U12811 (N_12811,N_8005,N_9406);
or U12812 (N_12812,N_6532,N_5178);
nor U12813 (N_12813,N_8275,N_6021);
nor U12814 (N_12814,N_5363,N_9063);
or U12815 (N_12815,N_6872,N_9054);
or U12816 (N_12816,N_8331,N_8240);
and U12817 (N_12817,N_6829,N_8188);
and U12818 (N_12818,N_9670,N_6865);
or U12819 (N_12819,N_8618,N_7613);
or U12820 (N_12820,N_6765,N_5786);
or U12821 (N_12821,N_9490,N_8316);
and U12822 (N_12822,N_9019,N_8399);
and U12823 (N_12823,N_9748,N_6334);
and U12824 (N_12824,N_9054,N_8730);
nand U12825 (N_12825,N_6121,N_8637);
nand U12826 (N_12826,N_5924,N_7353);
or U12827 (N_12827,N_5809,N_8307);
nand U12828 (N_12828,N_5621,N_9137);
xor U12829 (N_12829,N_5669,N_5598);
or U12830 (N_12830,N_9633,N_9417);
and U12831 (N_12831,N_8232,N_6413);
xor U12832 (N_12832,N_7387,N_8897);
or U12833 (N_12833,N_8671,N_8781);
nand U12834 (N_12834,N_7097,N_5557);
or U12835 (N_12835,N_5031,N_9869);
nand U12836 (N_12836,N_8335,N_7320);
xnor U12837 (N_12837,N_8779,N_7495);
or U12838 (N_12838,N_5101,N_8346);
or U12839 (N_12839,N_6236,N_8306);
nand U12840 (N_12840,N_9474,N_8732);
and U12841 (N_12841,N_7686,N_6903);
or U12842 (N_12842,N_5500,N_7077);
or U12843 (N_12843,N_9766,N_6144);
or U12844 (N_12844,N_5058,N_8394);
nand U12845 (N_12845,N_8505,N_5197);
nand U12846 (N_12846,N_7446,N_9959);
and U12847 (N_12847,N_8571,N_6725);
or U12848 (N_12848,N_7531,N_6806);
and U12849 (N_12849,N_9822,N_6674);
and U12850 (N_12850,N_5571,N_6226);
nor U12851 (N_12851,N_7820,N_7156);
and U12852 (N_12852,N_7305,N_6764);
nand U12853 (N_12853,N_9664,N_7092);
nor U12854 (N_12854,N_9844,N_8410);
nand U12855 (N_12855,N_5193,N_9394);
nand U12856 (N_12856,N_7992,N_8186);
nand U12857 (N_12857,N_5799,N_6574);
nand U12858 (N_12858,N_8107,N_5131);
nor U12859 (N_12859,N_6705,N_5799);
or U12860 (N_12860,N_8326,N_8539);
and U12861 (N_12861,N_5930,N_5821);
and U12862 (N_12862,N_9799,N_6002);
nor U12863 (N_12863,N_6251,N_6105);
nand U12864 (N_12864,N_6073,N_6696);
nor U12865 (N_12865,N_7099,N_8982);
or U12866 (N_12866,N_7123,N_5044);
and U12867 (N_12867,N_7469,N_6155);
and U12868 (N_12868,N_9641,N_8044);
or U12869 (N_12869,N_9056,N_5333);
nor U12870 (N_12870,N_8101,N_5912);
nor U12871 (N_12871,N_5361,N_8116);
nand U12872 (N_12872,N_5949,N_7796);
or U12873 (N_12873,N_8576,N_8661);
nor U12874 (N_12874,N_6026,N_5106);
or U12875 (N_12875,N_5383,N_9134);
and U12876 (N_12876,N_7564,N_7390);
nand U12877 (N_12877,N_5278,N_5221);
or U12878 (N_12878,N_7779,N_6241);
and U12879 (N_12879,N_7054,N_6683);
nand U12880 (N_12880,N_9299,N_8477);
nand U12881 (N_12881,N_8117,N_5753);
nand U12882 (N_12882,N_8404,N_5844);
or U12883 (N_12883,N_9958,N_6060);
or U12884 (N_12884,N_5526,N_9303);
nor U12885 (N_12885,N_9103,N_7079);
and U12886 (N_12886,N_7509,N_8136);
or U12887 (N_12887,N_6911,N_6419);
nor U12888 (N_12888,N_7978,N_5431);
nand U12889 (N_12889,N_6881,N_7233);
nand U12890 (N_12890,N_5484,N_6426);
or U12891 (N_12891,N_9630,N_9416);
and U12892 (N_12892,N_7280,N_7631);
or U12893 (N_12893,N_8139,N_6715);
or U12894 (N_12894,N_5367,N_5106);
and U12895 (N_12895,N_5917,N_9904);
or U12896 (N_12896,N_6642,N_6133);
nand U12897 (N_12897,N_5433,N_6147);
nor U12898 (N_12898,N_9907,N_5571);
and U12899 (N_12899,N_7022,N_9041);
or U12900 (N_12900,N_9308,N_7337);
or U12901 (N_12901,N_5759,N_6153);
nand U12902 (N_12902,N_9042,N_5782);
or U12903 (N_12903,N_8340,N_8209);
or U12904 (N_12904,N_9030,N_9731);
and U12905 (N_12905,N_8862,N_5800);
or U12906 (N_12906,N_9140,N_7401);
nand U12907 (N_12907,N_6329,N_6157);
and U12908 (N_12908,N_8696,N_5091);
nor U12909 (N_12909,N_5525,N_8955);
nand U12910 (N_12910,N_8715,N_7644);
or U12911 (N_12911,N_7655,N_6410);
and U12912 (N_12912,N_9844,N_9986);
or U12913 (N_12913,N_8252,N_8130);
or U12914 (N_12914,N_8687,N_5183);
and U12915 (N_12915,N_6882,N_7871);
or U12916 (N_12916,N_6986,N_6108);
nor U12917 (N_12917,N_8991,N_6424);
nand U12918 (N_12918,N_9371,N_6933);
and U12919 (N_12919,N_9151,N_5284);
or U12920 (N_12920,N_6621,N_8999);
nand U12921 (N_12921,N_9052,N_6761);
or U12922 (N_12922,N_6605,N_8315);
and U12923 (N_12923,N_8342,N_9725);
and U12924 (N_12924,N_7522,N_6513);
and U12925 (N_12925,N_6214,N_9011);
nor U12926 (N_12926,N_9581,N_8790);
and U12927 (N_12927,N_5944,N_7096);
nor U12928 (N_12928,N_6781,N_6005);
nor U12929 (N_12929,N_7218,N_6525);
nor U12930 (N_12930,N_9104,N_9651);
or U12931 (N_12931,N_6032,N_7283);
nor U12932 (N_12932,N_7634,N_9804);
nand U12933 (N_12933,N_8984,N_5248);
or U12934 (N_12934,N_7008,N_5699);
and U12935 (N_12935,N_8499,N_7912);
nand U12936 (N_12936,N_8273,N_8443);
nand U12937 (N_12937,N_9285,N_7714);
nor U12938 (N_12938,N_5411,N_7498);
nand U12939 (N_12939,N_8813,N_8523);
nor U12940 (N_12940,N_9206,N_5967);
or U12941 (N_12941,N_5015,N_5568);
or U12942 (N_12942,N_9714,N_5676);
and U12943 (N_12943,N_5328,N_9692);
nand U12944 (N_12944,N_5117,N_8197);
nor U12945 (N_12945,N_7647,N_9389);
nor U12946 (N_12946,N_8206,N_6379);
and U12947 (N_12947,N_7376,N_5106);
nor U12948 (N_12948,N_7128,N_9428);
and U12949 (N_12949,N_8693,N_6223);
nand U12950 (N_12950,N_6960,N_5452);
and U12951 (N_12951,N_5277,N_5524);
nand U12952 (N_12952,N_5766,N_7597);
and U12953 (N_12953,N_9971,N_6519);
nor U12954 (N_12954,N_6515,N_9348);
nor U12955 (N_12955,N_5356,N_5308);
nand U12956 (N_12956,N_9513,N_9207);
and U12957 (N_12957,N_7600,N_7277);
or U12958 (N_12958,N_7818,N_5725);
nand U12959 (N_12959,N_7101,N_5830);
or U12960 (N_12960,N_7624,N_8390);
nor U12961 (N_12961,N_7327,N_9534);
nor U12962 (N_12962,N_8261,N_6204);
nor U12963 (N_12963,N_6577,N_7854);
and U12964 (N_12964,N_5475,N_5173);
nor U12965 (N_12965,N_9680,N_8483);
or U12966 (N_12966,N_7647,N_5834);
nor U12967 (N_12967,N_8034,N_6820);
or U12968 (N_12968,N_8805,N_9781);
nor U12969 (N_12969,N_8381,N_5993);
nor U12970 (N_12970,N_8521,N_8438);
and U12971 (N_12971,N_6368,N_6269);
nor U12972 (N_12972,N_6077,N_7323);
and U12973 (N_12973,N_5950,N_9593);
or U12974 (N_12974,N_7137,N_8045);
nand U12975 (N_12975,N_6248,N_6313);
nor U12976 (N_12976,N_6001,N_8976);
and U12977 (N_12977,N_8461,N_7683);
and U12978 (N_12978,N_8432,N_8493);
or U12979 (N_12979,N_6560,N_6728);
nor U12980 (N_12980,N_5706,N_8868);
nand U12981 (N_12981,N_5458,N_8500);
or U12982 (N_12982,N_5836,N_5815);
or U12983 (N_12983,N_9889,N_6881);
and U12984 (N_12984,N_7167,N_6153);
and U12985 (N_12985,N_9882,N_9261);
and U12986 (N_12986,N_8360,N_6749);
and U12987 (N_12987,N_6162,N_8584);
and U12988 (N_12988,N_8426,N_7714);
and U12989 (N_12989,N_6002,N_8637);
and U12990 (N_12990,N_7461,N_9842);
nand U12991 (N_12991,N_6925,N_9686);
or U12992 (N_12992,N_5100,N_8870);
or U12993 (N_12993,N_6911,N_8814);
nand U12994 (N_12994,N_7620,N_8126);
nor U12995 (N_12995,N_5968,N_8463);
nand U12996 (N_12996,N_9295,N_5755);
nor U12997 (N_12997,N_8278,N_5836);
and U12998 (N_12998,N_6471,N_5340);
nor U12999 (N_12999,N_6842,N_7419);
nor U13000 (N_13000,N_5724,N_8055);
or U13001 (N_13001,N_9438,N_8735);
or U13002 (N_13002,N_9588,N_8098);
and U13003 (N_13003,N_7604,N_5385);
nor U13004 (N_13004,N_5872,N_9726);
nor U13005 (N_13005,N_9128,N_6369);
nor U13006 (N_13006,N_8088,N_8705);
or U13007 (N_13007,N_6798,N_8582);
nor U13008 (N_13008,N_5548,N_5698);
and U13009 (N_13009,N_6549,N_8706);
nor U13010 (N_13010,N_6371,N_5186);
or U13011 (N_13011,N_5421,N_8491);
nor U13012 (N_13012,N_8778,N_7171);
nor U13013 (N_13013,N_9888,N_6865);
or U13014 (N_13014,N_9274,N_5560);
and U13015 (N_13015,N_8493,N_8024);
nand U13016 (N_13016,N_6425,N_6181);
nor U13017 (N_13017,N_7093,N_7499);
nor U13018 (N_13018,N_9660,N_8781);
and U13019 (N_13019,N_5164,N_6743);
nor U13020 (N_13020,N_5442,N_5750);
and U13021 (N_13021,N_6564,N_6691);
nor U13022 (N_13022,N_7311,N_7869);
or U13023 (N_13023,N_8164,N_6742);
nand U13024 (N_13024,N_5058,N_9478);
and U13025 (N_13025,N_6448,N_7907);
xor U13026 (N_13026,N_8220,N_9298);
or U13027 (N_13027,N_6512,N_5343);
or U13028 (N_13028,N_7380,N_6395);
and U13029 (N_13029,N_6007,N_5698);
nor U13030 (N_13030,N_9784,N_9474);
or U13031 (N_13031,N_5265,N_7559);
or U13032 (N_13032,N_5872,N_8414);
nand U13033 (N_13033,N_5569,N_9784);
and U13034 (N_13034,N_7353,N_6901);
nor U13035 (N_13035,N_9322,N_5145);
and U13036 (N_13036,N_9638,N_5541);
and U13037 (N_13037,N_6634,N_8986);
and U13038 (N_13038,N_5827,N_7018);
and U13039 (N_13039,N_5658,N_9624);
or U13040 (N_13040,N_5661,N_8156);
and U13041 (N_13041,N_7258,N_8808);
nor U13042 (N_13042,N_9328,N_8026);
nor U13043 (N_13043,N_8352,N_5062);
or U13044 (N_13044,N_5060,N_5665);
or U13045 (N_13045,N_5516,N_5749);
nor U13046 (N_13046,N_6083,N_7340);
nor U13047 (N_13047,N_7046,N_7610);
nand U13048 (N_13048,N_9849,N_5219);
nor U13049 (N_13049,N_8449,N_8588);
nand U13050 (N_13050,N_7920,N_8841);
and U13051 (N_13051,N_7385,N_8325);
nand U13052 (N_13052,N_9806,N_8258);
nor U13053 (N_13053,N_6915,N_5225);
or U13054 (N_13054,N_6530,N_8455);
and U13055 (N_13055,N_7238,N_7499);
nand U13056 (N_13056,N_5718,N_6869);
and U13057 (N_13057,N_7786,N_9283);
and U13058 (N_13058,N_6461,N_9403);
nor U13059 (N_13059,N_8094,N_5035);
nand U13060 (N_13060,N_8718,N_8459);
or U13061 (N_13061,N_6180,N_8969);
nand U13062 (N_13062,N_9912,N_8333);
and U13063 (N_13063,N_9622,N_9026);
and U13064 (N_13064,N_9217,N_8017);
and U13065 (N_13065,N_8745,N_7199);
nand U13066 (N_13066,N_5106,N_7339);
nor U13067 (N_13067,N_6044,N_5621);
or U13068 (N_13068,N_9889,N_7038);
or U13069 (N_13069,N_9255,N_7777);
or U13070 (N_13070,N_8251,N_8478);
or U13071 (N_13071,N_7767,N_7513);
and U13072 (N_13072,N_8253,N_7088);
or U13073 (N_13073,N_8090,N_7161);
nand U13074 (N_13074,N_9570,N_5401);
or U13075 (N_13075,N_5149,N_8896);
nand U13076 (N_13076,N_6801,N_8509);
nand U13077 (N_13077,N_6654,N_8609);
and U13078 (N_13078,N_8223,N_9171);
and U13079 (N_13079,N_6390,N_6769);
nand U13080 (N_13080,N_6245,N_6360);
nand U13081 (N_13081,N_6356,N_7694);
and U13082 (N_13082,N_5138,N_9655);
nor U13083 (N_13083,N_5936,N_7712);
or U13084 (N_13084,N_9853,N_5691);
or U13085 (N_13085,N_8527,N_5718);
nand U13086 (N_13086,N_8467,N_7461);
nor U13087 (N_13087,N_5088,N_6082);
and U13088 (N_13088,N_7586,N_7934);
or U13089 (N_13089,N_6618,N_7327);
nand U13090 (N_13090,N_8747,N_6602);
nand U13091 (N_13091,N_8319,N_5094);
nor U13092 (N_13092,N_9023,N_8955);
or U13093 (N_13093,N_7149,N_7594);
and U13094 (N_13094,N_7840,N_8890);
or U13095 (N_13095,N_7091,N_5058);
nand U13096 (N_13096,N_5883,N_6395);
or U13097 (N_13097,N_8768,N_9722);
and U13098 (N_13098,N_8665,N_5288);
nand U13099 (N_13099,N_8542,N_8352);
nand U13100 (N_13100,N_8059,N_9912);
nand U13101 (N_13101,N_8304,N_7762);
and U13102 (N_13102,N_8880,N_9379);
nor U13103 (N_13103,N_9240,N_9279);
nor U13104 (N_13104,N_7735,N_7650);
and U13105 (N_13105,N_7753,N_6424);
nor U13106 (N_13106,N_9631,N_5978);
and U13107 (N_13107,N_7690,N_9211);
and U13108 (N_13108,N_5594,N_8398);
and U13109 (N_13109,N_8154,N_7691);
and U13110 (N_13110,N_9311,N_9880);
nor U13111 (N_13111,N_9695,N_6135);
nand U13112 (N_13112,N_9463,N_8723);
nor U13113 (N_13113,N_5945,N_5692);
and U13114 (N_13114,N_5677,N_9114);
xor U13115 (N_13115,N_8690,N_6140);
and U13116 (N_13116,N_6201,N_5987);
nor U13117 (N_13117,N_5610,N_5421);
and U13118 (N_13118,N_6578,N_5909);
nand U13119 (N_13119,N_7591,N_9768);
nor U13120 (N_13120,N_8323,N_5208);
nor U13121 (N_13121,N_9847,N_6001);
and U13122 (N_13122,N_7922,N_5263);
or U13123 (N_13123,N_7096,N_9624);
or U13124 (N_13124,N_9108,N_6654);
and U13125 (N_13125,N_9562,N_7538);
nor U13126 (N_13126,N_5510,N_6429);
or U13127 (N_13127,N_6172,N_9816);
or U13128 (N_13128,N_8793,N_5264);
or U13129 (N_13129,N_9826,N_8483);
nor U13130 (N_13130,N_5237,N_9386);
or U13131 (N_13131,N_5717,N_8276);
or U13132 (N_13132,N_7867,N_9497);
and U13133 (N_13133,N_6754,N_9289);
nand U13134 (N_13134,N_6317,N_5087);
nand U13135 (N_13135,N_8909,N_7663);
nor U13136 (N_13136,N_6128,N_5859);
and U13137 (N_13137,N_8451,N_9855);
nand U13138 (N_13138,N_5995,N_6008);
nand U13139 (N_13139,N_8758,N_9476);
nand U13140 (N_13140,N_8305,N_6458);
and U13141 (N_13141,N_9501,N_7884);
and U13142 (N_13142,N_5175,N_9662);
nand U13143 (N_13143,N_7544,N_7706);
nor U13144 (N_13144,N_5869,N_5264);
nand U13145 (N_13145,N_7799,N_8400);
nand U13146 (N_13146,N_6737,N_6877);
nand U13147 (N_13147,N_6428,N_6666);
or U13148 (N_13148,N_6539,N_9779);
or U13149 (N_13149,N_5957,N_6291);
nand U13150 (N_13150,N_5082,N_9577);
xnor U13151 (N_13151,N_8416,N_5734);
nand U13152 (N_13152,N_7792,N_6346);
and U13153 (N_13153,N_5327,N_6699);
nand U13154 (N_13154,N_6127,N_9377);
nand U13155 (N_13155,N_9073,N_7053);
nor U13156 (N_13156,N_5596,N_5974);
and U13157 (N_13157,N_5639,N_6447);
or U13158 (N_13158,N_9062,N_8473);
nand U13159 (N_13159,N_9312,N_8736);
nor U13160 (N_13160,N_7772,N_9957);
nand U13161 (N_13161,N_9018,N_5374);
or U13162 (N_13162,N_8308,N_5425);
nand U13163 (N_13163,N_5105,N_8268);
and U13164 (N_13164,N_7336,N_6916);
nand U13165 (N_13165,N_9775,N_7753);
nor U13166 (N_13166,N_7804,N_5635);
nand U13167 (N_13167,N_5068,N_8054);
nand U13168 (N_13168,N_9896,N_6893);
nor U13169 (N_13169,N_5473,N_7131);
and U13170 (N_13170,N_6417,N_6739);
and U13171 (N_13171,N_9771,N_5409);
nor U13172 (N_13172,N_8757,N_8637);
and U13173 (N_13173,N_6805,N_5484);
nor U13174 (N_13174,N_5370,N_7904);
nor U13175 (N_13175,N_7880,N_7559);
and U13176 (N_13176,N_6034,N_6001);
and U13177 (N_13177,N_7446,N_7320);
and U13178 (N_13178,N_8465,N_9719);
nor U13179 (N_13179,N_8021,N_7019);
nand U13180 (N_13180,N_5560,N_8190);
nor U13181 (N_13181,N_5870,N_6456);
nor U13182 (N_13182,N_9866,N_6968);
and U13183 (N_13183,N_7751,N_5088);
or U13184 (N_13184,N_7771,N_5016);
nor U13185 (N_13185,N_6569,N_9923);
nor U13186 (N_13186,N_9371,N_5207);
and U13187 (N_13187,N_7351,N_9352);
nor U13188 (N_13188,N_9312,N_9047);
nand U13189 (N_13189,N_5368,N_8455);
nand U13190 (N_13190,N_5112,N_8850);
and U13191 (N_13191,N_5367,N_6776);
nor U13192 (N_13192,N_5272,N_9211);
nand U13193 (N_13193,N_6574,N_8856);
and U13194 (N_13194,N_6627,N_5517);
and U13195 (N_13195,N_5969,N_5618);
nor U13196 (N_13196,N_7396,N_5231);
or U13197 (N_13197,N_8075,N_9137);
or U13198 (N_13198,N_6633,N_7042);
or U13199 (N_13199,N_5132,N_6435);
and U13200 (N_13200,N_5741,N_8129);
and U13201 (N_13201,N_5463,N_9151);
and U13202 (N_13202,N_8690,N_9687);
nor U13203 (N_13203,N_5941,N_5873);
and U13204 (N_13204,N_5748,N_7161);
nand U13205 (N_13205,N_5949,N_7653);
nand U13206 (N_13206,N_9769,N_5403);
nand U13207 (N_13207,N_9332,N_6411);
and U13208 (N_13208,N_6140,N_6687);
and U13209 (N_13209,N_6553,N_6496);
or U13210 (N_13210,N_5782,N_7824);
nor U13211 (N_13211,N_9691,N_7678);
or U13212 (N_13212,N_7811,N_8491);
nand U13213 (N_13213,N_5015,N_5760);
nor U13214 (N_13214,N_9664,N_6749);
nor U13215 (N_13215,N_9270,N_7119);
and U13216 (N_13216,N_6566,N_8730);
nand U13217 (N_13217,N_8376,N_7092);
nor U13218 (N_13218,N_9353,N_7535);
nor U13219 (N_13219,N_8115,N_9126);
or U13220 (N_13220,N_8890,N_9984);
nand U13221 (N_13221,N_8151,N_6528);
nor U13222 (N_13222,N_6593,N_9344);
nand U13223 (N_13223,N_8209,N_5386);
nor U13224 (N_13224,N_6747,N_5908);
and U13225 (N_13225,N_5765,N_6855);
nand U13226 (N_13226,N_6384,N_7664);
and U13227 (N_13227,N_8394,N_6994);
nor U13228 (N_13228,N_9487,N_7337);
and U13229 (N_13229,N_7076,N_5852);
or U13230 (N_13230,N_6351,N_6896);
nor U13231 (N_13231,N_6303,N_5838);
nand U13232 (N_13232,N_9328,N_7268);
or U13233 (N_13233,N_8231,N_5698);
nor U13234 (N_13234,N_7113,N_8609);
nor U13235 (N_13235,N_9486,N_7565);
nand U13236 (N_13236,N_6408,N_6138);
and U13237 (N_13237,N_5279,N_9192);
nand U13238 (N_13238,N_9338,N_5724);
nand U13239 (N_13239,N_8431,N_6895);
nor U13240 (N_13240,N_8381,N_5100);
or U13241 (N_13241,N_8714,N_8581);
nor U13242 (N_13242,N_9437,N_9527);
nor U13243 (N_13243,N_5605,N_8648);
or U13244 (N_13244,N_6036,N_7778);
and U13245 (N_13245,N_9560,N_7339);
nand U13246 (N_13246,N_5318,N_5692);
nand U13247 (N_13247,N_7513,N_7837);
and U13248 (N_13248,N_5576,N_5794);
nand U13249 (N_13249,N_9808,N_8652);
or U13250 (N_13250,N_6999,N_9846);
or U13251 (N_13251,N_7485,N_8321);
nand U13252 (N_13252,N_6342,N_6909);
and U13253 (N_13253,N_7256,N_7464);
nor U13254 (N_13254,N_5216,N_7921);
nor U13255 (N_13255,N_5325,N_5720);
or U13256 (N_13256,N_8667,N_5000);
nor U13257 (N_13257,N_5751,N_7862);
nand U13258 (N_13258,N_9304,N_9036);
and U13259 (N_13259,N_6139,N_6429);
or U13260 (N_13260,N_8395,N_8360);
nor U13261 (N_13261,N_9902,N_9363);
nor U13262 (N_13262,N_9164,N_5506);
xor U13263 (N_13263,N_5113,N_6077);
or U13264 (N_13264,N_5015,N_8018);
or U13265 (N_13265,N_8392,N_7506);
nor U13266 (N_13266,N_5254,N_5562);
nand U13267 (N_13267,N_9845,N_5460);
or U13268 (N_13268,N_7303,N_6255);
nor U13269 (N_13269,N_8072,N_7223);
or U13270 (N_13270,N_6187,N_7529);
or U13271 (N_13271,N_8205,N_8802);
nand U13272 (N_13272,N_7416,N_8479);
and U13273 (N_13273,N_5233,N_8543);
nor U13274 (N_13274,N_9440,N_9645);
xnor U13275 (N_13275,N_6271,N_8753);
nor U13276 (N_13276,N_9989,N_5804);
and U13277 (N_13277,N_5521,N_6923);
and U13278 (N_13278,N_6061,N_6423);
or U13279 (N_13279,N_8680,N_8011);
and U13280 (N_13280,N_9784,N_9302);
and U13281 (N_13281,N_7481,N_5028);
nor U13282 (N_13282,N_8108,N_7288);
or U13283 (N_13283,N_6867,N_9496);
nor U13284 (N_13284,N_9579,N_5593);
and U13285 (N_13285,N_6721,N_9993);
nor U13286 (N_13286,N_7500,N_5788);
or U13287 (N_13287,N_6784,N_8176);
and U13288 (N_13288,N_6940,N_9211);
nand U13289 (N_13289,N_6513,N_6612);
nand U13290 (N_13290,N_8430,N_5493);
nor U13291 (N_13291,N_5970,N_7389);
nor U13292 (N_13292,N_8911,N_9989);
nand U13293 (N_13293,N_9813,N_7758);
nor U13294 (N_13294,N_7295,N_5133);
or U13295 (N_13295,N_8160,N_5760);
nand U13296 (N_13296,N_9154,N_8923);
xnor U13297 (N_13297,N_8054,N_5550);
or U13298 (N_13298,N_6361,N_8084);
or U13299 (N_13299,N_7284,N_8559);
and U13300 (N_13300,N_6801,N_8725);
nand U13301 (N_13301,N_7415,N_9834);
or U13302 (N_13302,N_9410,N_7184);
or U13303 (N_13303,N_9519,N_7779);
nor U13304 (N_13304,N_5863,N_9332);
nand U13305 (N_13305,N_8589,N_5022);
and U13306 (N_13306,N_9201,N_5592);
nor U13307 (N_13307,N_9663,N_6393);
nand U13308 (N_13308,N_6863,N_7172);
nor U13309 (N_13309,N_6330,N_9461);
or U13310 (N_13310,N_9352,N_8082);
nand U13311 (N_13311,N_8397,N_7246);
and U13312 (N_13312,N_6681,N_7558);
nor U13313 (N_13313,N_9819,N_9221);
nor U13314 (N_13314,N_6138,N_5760);
nand U13315 (N_13315,N_5049,N_6251);
nand U13316 (N_13316,N_5070,N_5513);
nand U13317 (N_13317,N_9746,N_5126);
and U13318 (N_13318,N_9335,N_8023);
nor U13319 (N_13319,N_9823,N_9117);
and U13320 (N_13320,N_5971,N_5103);
and U13321 (N_13321,N_6724,N_6569);
and U13322 (N_13322,N_9062,N_9114);
nor U13323 (N_13323,N_7086,N_6400);
nor U13324 (N_13324,N_5503,N_9408);
or U13325 (N_13325,N_8955,N_6095);
and U13326 (N_13326,N_9282,N_5629);
or U13327 (N_13327,N_8596,N_5989);
nand U13328 (N_13328,N_8467,N_5766);
and U13329 (N_13329,N_6544,N_9794);
nor U13330 (N_13330,N_6430,N_9339);
or U13331 (N_13331,N_8783,N_8694);
or U13332 (N_13332,N_7791,N_9302);
and U13333 (N_13333,N_9790,N_7547);
nand U13334 (N_13334,N_6715,N_6422);
and U13335 (N_13335,N_7023,N_8017);
nor U13336 (N_13336,N_7501,N_9388);
and U13337 (N_13337,N_6449,N_9331);
nor U13338 (N_13338,N_6503,N_5151);
nor U13339 (N_13339,N_5427,N_5367);
and U13340 (N_13340,N_6674,N_8282);
nand U13341 (N_13341,N_5289,N_7849);
nand U13342 (N_13342,N_9336,N_6940);
nor U13343 (N_13343,N_6567,N_8144);
nand U13344 (N_13344,N_9909,N_5690);
nor U13345 (N_13345,N_7595,N_5356);
nor U13346 (N_13346,N_7778,N_6396);
nand U13347 (N_13347,N_5034,N_7710);
nand U13348 (N_13348,N_7718,N_6278);
and U13349 (N_13349,N_7590,N_8074);
or U13350 (N_13350,N_7639,N_8317);
nand U13351 (N_13351,N_7031,N_9305);
nor U13352 (N_13352,N_6335,N_9830);
nor U13353 (N_13353,N_7181,N_9387);
or U13354 (N_13354,N_6565,N_9977);
xnor U13355 (N_13355,N_7206,N_6287);
and U13356 (N_13356,N_9678,N_8731);
xor U13357 (N_13357,N_9389,N_6475);
xnor U13358 (N_13358,N_5471,N_6239);
nand U13359 (N_13359,N_5616,N_9117);
and U13360 (N_13360,N_7969,N_8158);
nand U13361 (N_13361,N_7597,N_8273);
nor U13362 (N_13362,N_7909,N_6502);
and U13363 (N_13363,N_9842,N_7900);
nor U13364 (N_13364,N_7947,N_5441);
nor U13365 (N_13365,N_5791,N_5793);
nor U13366 (N_13366,N_6015,N_7715);
and U13367 (N_13367,N_5449,N_8803);
nor U13368 (N_13368,N_5341,N_8437);
or U13369 (N_13369,N_9138,N_6828);
nor U13370 (N_13370,N_7963,N_7705);
and U13371 (N_13371,N_9652,N_8838);
nand U13372 (N_13372,N_6355,N_7779);
and U13373 (N_13373,N_6555,N_9333);
and U13374 (N_13374,N_7886,N_9990);
or U13375 (N_13375,N_7178,N_9237);
xnor U13376 (N_13376,N_9170,N_7041);
and U13377 (N_13377,N_7490,N_5285);
or U13378 (N_13378,N_5951,N_7569);
nor U13379 (N_13379,N_5172,N_8056);
or U13380 (N_13380,N_6049,N_6437);
and U13381 (N_13381,N_8069,N_9442);
and U13382 (N_13382,N_8183,N_7612);
nand U13383 (N_13383,N_8245,N_9542);
nand U13384 (N_13384,N_9631,N_7664);
or U13385 (N_13385,N_7512,N_7552);
or U13386 (N_13386,N_8237,N_9387);
and U13387 (N_13387,N_9435,N_7506);
nand U13388 (N_13388,N_8618,N_5859);
nand U13389 (N_13389,N_8845,N_6925);
and U13390 (N_13390,N_9704,N_9630);
and U13391 (N_13391,N_6154,N_9604);
nor U13392 (N_13392,N_7533,N_6392);
or U13393 (N_13393,N_5216,N_6280);
nand U13394 (N_13394,N_7440,N_7088);
or U13395 (N_13395,N_5908,N_5012);
or U13396 (N_13396,N_5944,N_7845);
or U13397 (N_13397,N_5892,N_8064);
nand U13398 (N_13398,N_7105,N_7359);
nor U13399 (N_13399,N_6880,N_8132);
nor U13400 (N_13400,N_5613,N_9727);
nand U13401 (N_13401,N_8618,N_9488);
and U13402 (N_13402,N_8659,N_7214);
nor U13403 (N_13403,N_6075,N_9701);
or U13404 (N_13404,N_9118,N_9159);
or U13405 (N_13405,N_9967,N_5762);
or U13406 (N_13406,N_9540,N_5743);
or U13407 (N_13407,N_8597,N_6851);
and U13408 (N_13408,N_7087,N_7878);
nor U13409 (N_13409,N_5033,N_8452);
and U13410 (N_13410,N_9504,N_6470);
nor U13411 (N_13411,N_7351,N_5801);
nor U13412 (N_13412,N_5828,N_5766);
or U13413 (N_13413,N_6564,N_7820);
or U13414 (N_13414,N_5670,N_5278);
or U13415 (N_13415,N_5851,N_6472);
or U13416 (N_13416,N_6532,N_7204);
nand U13417 (N_13417,N_7100,N_8694);
and U13418 (N_13418,N_7119,N_7294);
nor U13419 (N_13419,N_5309,N_7174);
xnor U13420 (N_13420,N_8555,N_9625);
or U13421 (N_13421,N_6037,N_8999);
and U13422 (N_13422,N_9021,N_7570);
nor U13423 (N_13423,N_8304,N_5901);
or U13424 (N_13424,N_6114,N_6543);
nor U13425 (N_13425,N_7838,N_6539);
nand U13426 (N_13426,N_9831,N_7219);
or U13427 (N_13427,N_9320,N_8785);
or U13428 (N_13428,N_8656,N_8662);
or U13429 (N_13429,N_7484,N_8788);
or U13430 (N_13430,N_5679,N_6004);
and U13431 (N_13431,N_6353,N_8842);
and U13432 (N_13432,N_9700,N_8152);
or U13433 (N_13433,N_5267,N_6425);
or U13434 (N_13434,N_8952,N_7242);
or U13435 (N_13435,N_6311,N_9859);
and U13436 (N_13436,N_5737,N_9814);
or U13437 (N_13437,N_8052,N_7597);
or U13438 (N_13438,N_7425,N_7350);
nor U13439 (N_13439,N_7986,N_8118);
nand U13440 (N_13440,N_7940,N_9330);
or U13441 (N_13441,N_9080,N_8730);
nor U13442 (N_13442,N_5086,N_8844);
or U13443 (N_13443,N_8942,N_8317);
nand U13444 (N_13444,N_8078,N_7669);
or U13445 (N_13445,N_5501,N_7189);
and U13446 (N_13446,N_7490,N_8673);
nor U13447 (N_13447,N_9116,N_8921);
nor U13448 (N_13448,N_6496,N_7977);
or U13449 (N_13449,N_5584,N_9170);
nor U13450 (N_13450,N_6835,N_9618);
nand U13451 (N_13451,N_7610,N_6702);
and U13452 (N_13452,N_8043,N_6171);
or U13453 (N_13453,N_5932,N_8556);
and U13454 (N_13454,N_9772,N_6585);
or U13455 (N_13455,N_7242,N_7066);
or U13456 (N_13456,N_5014,N_8108);
and U13457 (N_13457,N_8777,N_5561);
or U13458 (N_13458,N_8772,N_6448);
or U13459 (N_13459,N_5090,N_6466);
and U13460 (N_13460,N_8973,N_7124);
and U13461 (N_13461,N_5196,N_5528);
nand U13462 (N_13462,N_6001,N_9569);
nand U13463 (N_13463,N_8620,N_7622);
nor U13464 (N_13464,N_6701,N_8517);
or U13465 (N_13465,N_9156,N_9383);
and U13466 (N_13466,N_9177,N_7021);
nand U13467 (N_13467,N_8217,N_6502);
nor U13468 (N_13468,N_7407,N_9603);
nand U13469 (N_13469,N_5809,N_8733);
nand U13470 (N_13470,N_5470,N_7212);
nor U13471 (N_13471,N_6141,N_9098);
and U13472 (N_13472,N_6991,N_8973);
or U13473 (N_13473,N_5206,N_6653);
nor U13474 (N_13474,N_6376,N_6615);
nand U13475 (N_13475,N_5779,N_9388);
or U13476 (N_13476,N_8131,N_6411);
or U13477 (N_13477,N_5283,N_5430);
and U13478 (N_13478,N_6295,N_9772);
or U13479 (N_13479,N_7533,N_9862);
or U13480 (N_13480,N_5747,N_9758);
and U13481 (N_13481,N_7067,N_8084);
nand U13482 (N_13482,N_7205,N_5293);
or U13483 (N_13483,N_8879,N_5104);
and U13484 (N_13484,N_9687,N_5014);
nor U13485 (N_13485,N_9640,N_9439);
nand U13486 (N_13486,N_9764,N_7027);
nand U13487 (N_13487,N_5285,N_8869);
nand U13488 (N_13488,N_7871,N_8351);
or U13489 (N_13489,N_8959,N_8766);
nor U13490 (N_13490,N_9454,N_9199);
or U13491 (N_13491,N_5041,N_7307);
and U13492 (N_13492,N_7126,N_7524);
or U13493 (N_13493,N_6546,N_9581);
nand U13494 (N_13494,N_5401,N_5532);
nor U13495 (N_13495,N_8906,N_5206);
and U13496 (N_13496,N_7468,N_7843);
or U13497 (N_13497,N_8692,N_8542);
nand U13498 (N_13498,N_5687,N_9375);
and U13499 (N_13499,N_6644,N_7606);
or U13500 (N_13500,N_6447,N_6472);
xor U13501 (N_13501,N_8710,N_9474);
nand U13502 (N_13502,N_8820,N_6183);
and U13503 (N_13503,N_7943,N_8499);
nor U13504 (N_13504,N_5268,N_8563);
nand U13505 (N_13505,N_5088,N_6662);
or U13506 (N_13506,N_5457,N_6481);
nand U13507 (N_13507,N_9513,N_8088);
or U13508 (N_13508,N_9798,N_9445);
or U13509 (N_13509,N_8503,N_5535);
nand U13510 (N_13510,N_7951,N_5943);
nand U13511 (N_13511,N_8530,N_7343);
nand U13512 (N_13512,N_8871,N_9104);
or U13513 (N_13513,N_5218,N_9104);
or U13514 (N_13514,N_8732,N_6387);
and U13515 (N_13515,N_7909,N_7466);
or U13516 (N_13516,N_9212,N_6182);
and U13517 (N_13517,N_9816,N_9688);
nand U13518 (N_13518,N_7538,N_7220);
nand U13519 (N_13519,N_6316,N_6485);
nand U13520 (N_13520,N_6002,N_5057);
nand U13521 (N_13521,N_6309,N_9271);
nand U13522 (N_13522,N_9255,N_7219);
and U13523 (N_13523,N_8157,N_7415);
or U13524 (N_13524,N_8351,N_9470);
xnor U13525 (N_13525,N_6218,N_7915);
nand U13526 (N_13526,N_6104,N_7068);
nand U13527 (N_13527,N_9818,N_5043);
nor U13528 (N_13528,N_6638,N_6954);
nor U13529 (N_13529,N_5452,N_7669);
nor U13530 (N_13530,N_5220,N_8982);
nor U13531 (N_13531,N_8859,N_7631);
or U13532 (N_13532,N_5999,N_6901);
nand U13533 (N_13533,N_5018,N_9546);
nor U13534 (N_13534,N_8046,N_9129);
or U13535 (N_13535,N_9835,N_6809);
and U13536 (N_13536,N_9140,N_7476);
and U13537 (N_13537,N_5717,N_8522);
or U13538 (N_13538,N_6994,N_6424);
nor U13539 (N_13539,N_8178,N_5423);
nand U13540 (N_13540,N_8178,N_7197);
nor U13541 (N_13541,N_7376,N_8584);
or U13542 (N_13542,N_7948,N_8710);
nand U13543 (N_13543,N_6131,N_6047);
nand U13544 (N_13544,N_6642,N_9675);
nor U13545 (N_13545,N_9933,N_6299);
nand U13546 (N_13546,N_8123,N_8294);
nor U13547 (N_13547,N_8241,N_5437);
and U13548 (N_13548,N_9498,N_5396);
and U13549 (N_13549,N_6772,N_9090);
nand U13550 (N_13550,N_5989,N_8261);
or U13551 (N_13551,N_7869,N_7712);
nor U13552 (N_13552,N_9109,N_9338);
and U13553 (N_13553,N_8237,N_5098);
and U13554 (N_13554,N_5006,N_7887);
nand U13555 (N_13555,N_8216,N_5427);
nor U13556 (N_13556,N_5842,N_8902);
and U13557 (N_13557,N_8505,N_6601);
nand U13558 (N_13558,N_7607,N_8411);
nor U13559 (N_13559,N_7560,N_8695);
or U13560 (N_13560,N_7883,N_6381);
and U13561 (N_13561,N_8060,N_7916);
or U13562 (N_13562,N_9046,N_6351);
nand U13563 (N_13563,N_6446,N_5710);
or U13564 (N_13564,N_5486,N_8459);
nand U13565 (N_13565,N_9358,N_7202);
or U13566 (N_13566,N_5633,N_6454);
or U13567 (N_13567,N_6506,N_9579);
or U13568 (N_13568,N_9080,N_9696);
and U13569 (N_13569,N_6667,N_6039);
or U13570 (N_13570,N_5525,N_5589);
and U13571 (N_13571,N_9294,N_6203);
and U13572 (N_13572,N_6074,N_6858);
or U13573 (N_13573,N_5858,N_5355);
nor U13574 (N_13574,N_9680,N_8902);
nand U13575 (N_13575,N_8336,N_8159);
xor U13576 (N_13576,N_7520,N_7868);
nor U13577 (N_13577,N_9524,N_8125);
nor U13578 (N_13578,N_8453,N_6569);
nand U13579 (N_13579,N_6057,N_8476);
nand U13580 (N_13580,N_5654,N_5748);
nand U13581 (N_13581,N_9705,N_6276);
nand U13582 (N_13582,N_9192,N_7265);
nor U13583 (N_13583,N_8143,N_7955);
nor U13584 (N_13584,N_8672,N_7822);
nand U13585 (N_13585,N_7920,N_8969);
nor U13586 (N_13586,N_5552,N_6052);
nor U13587 (N_13587,N_5682,N_8038);
or U13588 (N_13588,N_7574,N_9424);
or U13589 (N_13589,N_8853,N_9372);
nor U13590 (N_13590,N_6777,N_6286);
and U13591 (N_13591,N_8742,N_8162);
nand U13592 (N_13592,N_5286,N_6240);
nand U13593 (N_13593,N_7172,N_9321);
or U13594 (N_13594,N_5333,N_7879);
nor U13595 (N_13595,N_7542,N_9260);
nor U13596 (N_13596,N_6787,N_7272);
or U13597 (N_13597,N_7644,N_6617);
and U13598 (N_13598,N_5224,N_8159);
and U13599 (N_13599,N_6460,N_5262);
or U13600 (N_13600,N_5505,N_7228);
or U13601 (N_13601,N_7338,N_5085);
nand U13602 (N_13602,N_6263,N_7125);
nor U13603 (N_13603,N_8343,N_7406);
or U13604 (N_13604,N_9758,N_6229);
or U13605 (N_13605,N_8051,N_7054);
nand U13606 (N_13606,N_9074,N_6957);
nand U13607 (N_13607,N_5043,N_8155);
and U13608 (N_13608,N_5911,N_7336);
nor U13609 (N_13609,N_9530,N_8068);
nor U13610 (N_13610,N_5377,N_7869);
nor U13611 (N_13611,N_8348,N_9356);
nand U13612 (N_13612,N_8000,N_6001);
or U13613 (N_13613,N_6389,N_8040);
and U13614 (N_13614,N_8831,N_7124);
nand U13615 (N_13615,N_9693,N_9535);
nand U13616 (N_13616,N_5231,N_5332);
or U13617 (N_13617,N_9821,N_9928);
nand U13618 (N_13618,N_9091,N_9986);
nand U13619 (N_13619,N_8699,N_8240);
nor U13620 (N_13620,N_6975,N_8335);
nor U13621 (N_13621,N_8917,N_8338);
or U13622 (N_13622,N_8800,N_9427);
nor U13623 (N_13623,N_7101,N_6084);
nand U13624 (N_13624,N_9722,N_8427);
nor U13625 (N_13625,N_8942,N_7927);
nor U13626 (N_13626,N_9235,N_6971);
and U13627 (N_13627,N_7605,N_6383);
and U13628 (N_13628,N_6077,N_5369);
or U13629 (N_13629,N_5269,N_6990);
nor U13630 (N_13630,N_9676,N_6444);
nand U13631 (N_13631,N_5538,N_7198);
and U13632 (N_13632,N_5168,N_8932);
nor U13633 (N_13633,N_7139,N_5797);
nor U13634 (N_13634,N_7948,N_6589);
or U13635 (N_13635,N_8002,N_9737);
nand U13636 (N_13636,N_8987,N_8111);
and U13637 (N_13637,N_6231,N_5996);
nor U13638 (N_13638,N_8346,N_9939);
and U13639 (N_13639,N_8839,N_6691);
and U13640 (N_13640,N_7517,N_5407);
or U13641 (N_13641,N_5393,N_8787);
nor U13642 (N_13642,N_7548,N_7726);
nand U13643 (N_13643,N_8950,N_7776);
nor U13644 (N_13644,N_6179,N_7215);
or U13645 (N_13645,N_8192,N_7666);
and U13646 (N_13646,N_5086,N_5473);
xor U13647 (N_13647,N_5821,N_6350);
nor U13648 (N_13648,N_9162,N_7708);
or U13649 (N_13649,N_8630,N_9406);
or U13650 (N_13650,N_5935,N_8126);
xor U13651 (N_13651,N_7271,N_8783);
or U13652 (N_13652,N_9107,N_8773);
and U13653 (N_13653,N_8151,N_9455);
or U13654 (N_13654,N_6130,N_5878);
nand U13655 (N_13655,N_9576,N_9256);
and U13656 (N_13656,N_5263,N_5709);
and U13657 (N_13657,N_6792,N_6263);
nand U13658 (N_13658,N_6463,N_5463);
and U13659 (N_13659,N_6216,N_5746);
nand U13660 (N_13660,N_9781,N_9416);
nor U13661 (N_13661,N_8780,N_9747);
nor U13662 (N_13662,N_5056,N_8474);
nand U13663 (N_13663,N_8776,N_8886);
or U13664 (N_13664,N_5215,N_9655);
and U13665 (N_13665,N_9069,N_6876);
nor U13666 (N_13666,N_7297,N_8501);
nand U13667 (N_13667,N_7453,N_5497);
nand U13668 (N_13668,N_8748,N_5640);
nand U13669 (N_13669,N_6527,N_6403);
and U13670 (N_13670,N_9027,N_8792);
nor U13671 (N_13671,N_9214,N_6118);
nor U13672 (N_13672,N_6656,N_5911);
and U13673 (N_13673,N_8690,N_7206);
or U13674 (N_13674,N_5943,N_6383);
nor U13675 (N_13675,N_9643,N_7596);
nand U13676 (N_13676,N_9563,N_7746);
nand U13677 (N_13677,N_6335,N_5928);
nand U13678 (N_13678,N_6244,N_5837);
nor U13679 (N_13679,N_6487,N_5311);
or U13680 (N_13680,N_6510,N_7784);
nand U13681 (N_13681,N_5018,N_5987);
nand U13682 (N_13682,N_6246,N_6031);
nand U13683 (N_13683,N_7751,N_6030);
nand U13684 (N_13684,N_8420,N_9808);
nor U13685 (N_13685,N_5536,N_8159);
and U13686 (N_13686,N_8869,N_8537);
or U13687 (N_13687,N_8200,N_9186);
and U13688 (N_13688,N_7888,N_5286);
nor U13689 (N_13689,N_8276,N_9445);
or U13690 (N_13690,N_9774,N_6124);
nor U13691 (N_13691,N_9833,N_8824);
nand U13692 (N_13692,N_6848,N_5097);
nor U13693 (N_13693,N_8143,N_9859);
nand U13694 (N_13694,N_8266,N_7529);
or U13695 (N_13695,N_9035,N_6928);
and U13696 (N_13696,N_9505,N_6532);
or U13697 (N_13697,N_5094,N_6703);
nor U13698 (N_13698,N_5804,N_7775);
or U13699 (N_13699,N_9586,N_7084);
nor U13700 (N_13700,N_8331,N_5930);
nand U13701 (N_13701,N_8862,N_5049);
nand U13702 (N_13702,N_7013,N_5997);
and U13703 (N_13703,N_7762,N_7835);
and U13704 (N_13704,N_9938,N_7182);
or U13705 (N_13705,N_7473,N_8601);
nand U13706 (N_13706,N_8586,N_9666);
nor U13707 (N_13707,N_6001,N_8939);
nor U13708 (N_13708,N_5133,N_7435);
or U13709 (N_13709,N_9190,N_9140);
nand U13710 (N_13710,N_5230,N_7543);
nor U13711 (N_13711,N_6456,N_9717);
xnor U13712 (N_13712,N_8548,N_6520);
nor U13713 (N_13713,N_6275,N_7010);
nand U13714 (N_13714,N_7697,N_6594);
and U13715 (N_13715,N_9907,N_8023);
nand U13716 (N_13716,N_6397,N_5872);
nand U13717 (N_13717,N_5781,N_5921);
nor U13718 (N_13718,N_5725,N_6862);
nand U13719 (N_13719,N_8967,N_7306);
nor U13720 (N_13720,N_5790,N_8469);
and U13721 (N_13721,N_5483,N_6904);
nand U13722 (N_13722,N_9435,N_6727);
and U13723 (N_13723,N_9636,N_5526);
and U13724 (N_13724,N_8303,N_7416);
nor U13725 (N_13725,N_5500,N_9798);
nor U13726 (N_13726,N_8687,N_5817);
nor U13727 (N_13727,N_5691,N_6960);
or U13728 (N_13728,N_8987,N_8077);
nand U13729 (N_13729,N_8654,N_9329);
or U13730 (N_13730,N_7183,N_6423);
nor U13731 (N_13731,N_6784,N_9720);
nor U13732 (N_13732,N_6212,N_9726);
nor U13733 (N_13733,N_6141,N_5021);
nor U13734 (N_13734,N_8351,N_9252);
or U13735 (N_13735,N_6352,N_8925);
nor U13736 (N_13736,N_7186,N_5722);
nand U13737 (N_13737,N_9840,N_9704);
nand U13738 (N_13738,N_7508,N_8285);
nand U13739 (N_13739,N_7928,N_6756);
nand U13740 (N_13740,N_7875,N_8715);
or U13741 (N_13741,N_8219,N_6269);
nand U13742 (N_13742,N_5885,N_7027);
and U13743 (N_13743,N_5704,N_7570);
or U13744 (N_13744,N_5535,N_8913);
nor U13745 (N_13745,N_6379,N_8593);
nand U13746 (N_13746,N_6994,N_5118);
nand U13747 (N_13747,N_7230,N_7527);
or U13748 (N_13748,N_5057,N_9151);
or U13749 (N_13749,N_8853,N_5570);
nor U13750 (N_13750,N_6439,N_6362);
nor U13751 (N_13751,N_9748,N_9828);
nor U13752 (N_13752,N_7701,N_7222);
nand U13753 (N_13753,N_9868,N_5555);
nor U13754 (N_13754,N_5645,N_5421);
nand U13755 (N_13755,N_5199,N_8038);
nand U13756 (N_13756,N_5885,N_9146);
or U13757 (N_13757,N_6506,N_5014);
and U13758 (N_13758,N_6120,N_9173);
nor U13759 (N_13759,N_8285,N_6228);
nand U13760 (N_13760,N_9080,N_5958);
nand U13761 (N_13761,N_9056,N_8377);
and U13762 (N_13762,N_7002,N_9897);
or U13763 (N_13763,N_7579,N_8034);
or U13764 (N_13764,N_7873,N_6803);
nand U13765 (N_13765,N_9193,N_7151);
or U13766 (N_13766,N_8102,N_7892);
nor U13767 (N_13767,N_6424,N_5078);
or U13768 (N_13768,N_9375,N_6445);
nand U13769 (N_13769,N_5395,N_6292);
nor U13770 (N_13770,N_5676,N_5571);
nor U13771 (N_13771,N_9796,N_7657);
nor U13772 (N_13772,N_9692,N_8445);
nor U13773 (N_13773,N_8208,N_8790);
nand U13774 (N_13774,N_9906,N_6127);
nor U13775 (N_13775,N_7938,N_7113);
or U13776 (N_13776,N_6305,N_7373);
nand U13777 (N_13777,N_6556,N_7386);
nor U13778 (N_13778,N_9522,N_7443);
nor U13779 (N_13779,N_9960,N_7235);
nand U13780 (N_13780,N_8126,N_6369);
or U13781 (N_13781,N_9226,N_5973);
or U13782 (N_13782,N_6398,N_9058);
or U13783 (N_13783,N_5668,N_9748);
nor U13784 (N_13784,N_8882,N_5670);
and U13785 (N_13785,N_6073,N_5824);
nor U13786 (N_13786,N_7591,N_8130);
or U13787 (N_13787,N_8601,N_7725);
or U13788 (N_13788,N_9287,N_8441);
or U13789 (N_13789,N_8587,N_7924);
nand U13790 (N_13790,N_6092,N_8371);
nand U13791 (N_13791,N_8661,N_7863);
or U13792 (N_13792,N_7578,N_6994);
nand U13793 (N_13793,N_9802,N_7672);
and U13794 (N_13794,N_6716,N_8031);
or U13795 (N_13795,N_5910,N_5974);
nand U13796 (N_13796,N_6355,N_6570);
or U13797 (N_13797,N_9597,N_7805);
nand U13798 (N_13798,N_5935,N_5425);
nor U13799 (N_13799,N_6582,N_9934);
and U13800 (N_13800,N_5145,N_8034);
nand U13801 (N_13801,N_8330,N_6801);
and U13802 (N_13802,N_6899,N_6567);
nor U13803 (N_13803,N_8385,N_9071);
nor U13804 (N_13804,N_6340,N_9840);
and U13805 (N_13805,N_7741,N_6301);
nand U13806 (N_13806,N_5483,N_7809);
nand U13807 (N_13807,N_9773,N_5356);
nor U13808 (N_13808,N_6316,N_7675);
nor U13809 (N_13809,N_8099,N_6686);
nand U13810 (N_13810,N_8897,N_5067);
nand U13811 (N_13811,N_7880,N_5716);
nand U13812 (N_13812,N_5181,N_8198);
and U13813 (N_13813,N_6322,N_9029);
nand U13814 (N_13814,N_5236,N_5571);
nor U13815 (N_13815,N_8578,N_8866);
nand U13816 (N_13816,N_5205,N_6002);
nand U13817 (N_13817,N_8475,N_7552);
and U13818 (N_13818,N_9976,N_8516);
nor U13819 (N_13819,N_8218,N_8889);
nand U13820 (N_13820,N_6264,N_6869);
nor U13821 (N_13821,N_7988,N_9650);
nor U13822 (N_13822,N_6628,N_8621);
nand U13823 (N_13823,N_8588,N_9110);
nor U13824 (N_13824,N_7846,N_6778);
and U13825 (N_13825,N_7331,N_9612);
nor U13826 (N_13826,N_5697,N_8636);
or U13827 (N_13827,N_5813,N_7969);
and U13828 (N_13828,N_8020,N_9487);
and U13829 (N_13829,N_5194,N_7579);
xnor U13830 (N_13830,N_5089,N_9761);
and U13831 (N_13831,N_7678,N_5177);
nor U13832 (N_13832,N_6466,N_5883);
nand U13833 (N_13833,N_8243,N_5387);
or U13834 (N_13834,N_7810,N_7772);
or U13835 (N_13835,N_8957,N_8159);
xor U13836 (N_13836,N_6163,N_5182);
and U13837 (N_13837,N_5451,N_5688);
nor U13838 (N_13838,N_5415,N_9640);
nor U13839 (N_13839,N_7697,N_7756);
and U13840 (N_13840,N_8513,N_9428);
nand U13841 (N_13841,N_6725,N_7819);
or U13842 (N_13842,N_8630,N_7283);
or U13843 (N_13843,N_8294,N_6196);
and U13844 (N_13844,N_6328,N_9623);
or U13845 (N_13845,N_5917,N_7427);
and U13846 (N_13846,N_9141,N_8935);
and U13847 (N_13847,N_9928,N_8372);
or U13848 (N_13848,N_8367,N_9771);
or U13849 (N_13849,N_8322,N_5185);
nand U13850 (N_13850,N_5303,N_6250);
and U13851 (N_13851,N_7372,N_6024);
or U13852 (N_13852,N_7516,N_9316);
nand U13853 (N_13853,N_6793,N_9490);
nor U13854 (N_13854,N_6857,N_5763);
nand U13855 (N_13855,N_8388,N_6564);
nor U13856 (N_13856,N_9416,N_8926);
and U13857 (N_13857,N_5849,N_7250);
or U13858 (N_13858,N_8826,N_8093);
nand U13859 (N_13859,N_8972,N_5881);
nor U13860 (N_13860,N_5131,N_6249);
xor U13861 (N_13861,N_9113,N_6688);
or U13862 (N_13862,N_9769,N_6809);
and U13863 (N_13863,N_8462,N_8357);
nand U13864 (N_13864,N_6105,N_8011);
and U13865 (N_13865,N_5143,N_7100);
and U13866 (N_13866,N_8951,N_6067);
nor U13867 (N_13867,N_8769,N_5957);
nor U13868 (N_13868,N_9870,N_9865);
nor U13869 (N_13869,N_8083,N_5262);
and U13870 (N_13870,N_7321,N_5156);
nor U13871 (N_13871,N_9496,N_9324);
nand U13872 (N_13872,N_8664,N_9259);
xor U13873 (N_13873,N_5613,N_5502);
and U13874 (N_13874,N_9162,N_6502);
nor U13875 (N_13875,N_6257,N_7903);
nand U13876 (N_13876,N_6809,N_6233);
nand U13877 (N_13877,N_6036,N_5487);
nor U13878 (N_13878,N_7641,N_7575);
or U13879 (N_13879,N_5964,N_6112);
or U13880 (N_13880,N_5858,N_6154);
nand U13881 (N_13881,N_8793,N_7179);
and U13882 (N_13882,N_6818,N_7091);
and U13883 (N_13883,N_7840,N_8288);
nor U13884 (N_13884,N_7276,N_7908);
or U13885 (N_13885,N_7992,N_8814);
nor U13886 (N_13886,N_7366,N_6028);
and U13887 (N_13887,N_7208,N_7631);
nand U13888 (N_13888,N_6934,N_9843);
or U13889 (N_13889,N_8198,N_7885);
nand U13890 (N_13890,N_7947,N_9036);
and U13891 (N_13891,N_8841,N_7546);
nor U13892 (N_13892,N_9847,N_9446);
or U13893 (N_13893,N_5936,N_7677);
nor U13894 (N_13894,N_6508,N_5179);
and U13895 (N_13895,N_5695,N_9927);
nor U13896 (N_13896,N_8618,N_6441);
or U13897 (N_13897,N_8953,N_5838);
nand U13898 (N_13898,N_8174,N_5319);
nor U13899 (N_13899,N_8204,N_5003);
nand U13900 (N_13900,N_5667,N_7269);
nand U13901 (N_13901,N_5879,N_7603);
nor U13902 (N_13902,N_8640,N_9508);
nor U13903 (N_13903,N_6208,N_5945);
or U13904 (N_13904,N_9437,N_9930);
or U13905 (N_13905,N_7166,N_6176);
nand U13906 (N_13906,N_7711,N_9293);
nand U13907 (N_13907,N_6150,N_6549);
nand U13908 (N_13908,N_6022,N_7590);
or U13909 (N_13909,N_8938,N_7032);
nand U13910 (N_13910,N_7293,N_6855);
nand U13911 (N_13911,N_6992,N_8092);
nor U13912 (N_13912,N_6672,N_9855);
nand U13913 (N_13913,N_5061,N_5819);
and U13914 (N_13914,N_9721,N_5066);
and U13915 (N_13915,N_9469,N_8440);
nor U13916 (N_13916,N_8214,N_6239);
and U13917 (N_13917,N_6335,N_7941);
nand U13918 (N_13918,N_9084,N_8155);
and U13919 (N_13919,N_5486,N_9308);
nor U13920 (N_13920,N_8886,N_7368);
or U13921 (N_13921,N_5231,N_8396);
nor U13922 (N_13922,N_6545,N_7553);
or U13923 (N_13923,N_5047,N_6374);
or U13924 (N_13924,N_5067,N_8613);
nor U13925 (N_13925,N_7829,N_5821);
or U13926 (N_13926,N_5637,N_5455);
and U13927 (N_13927,N_8442,N_5958);
and U13928 (N_13928,N_6629,N_7276);
nand U13929 (N_13929,N_9006,N_9494);
nand U13930 (N_13930,N_9500,N_6944);
and U13931 (N_13931,N_6112,N_6237);
and U13932 (N_13932,N_6833,N_6420);
nand U13933 (N_13933,N_9011,N_9691);
or U13934 (N_13934,N_6123,N_8935);
and U13935 (N_13935,N_7156,N_8263);
or U13936 (N_13936,N_8184,N_7693);
and U13937 (N_13937,N_6556,N_6233);
nor U13938 (N_13938,N_5902,N_9268);
nor U13939 (N_13939,N_5399,N_6104);
and U13940 (N_13940,N_9508,N_5061);
or U13941 (N_13941,N_7094,N_6944);
and U13942 (N_13942,N_5766,N_8183);
and U13943 (N_13943,N_8759,N_7519);
nor U13944 (N_13944,N_9401,N_5039);
nor U13945 (N_13945,N_5566,N_9633);
or U13946 (N_13946,N_7251,N_9555);
or U13947 (N_13947,N_7397,N_8182);
or U13948 (N_13948,N_9159,N_8790);
nor U13949 (N_13949,N_6666,N_8450);
and U13950 (N_13950,N_5885,N_8332);
and U13951 (N_13951,N_7646,N_6082);
and U13952 (N_13952,N_8969,N_6904);
nand U13953 (N_13953,N_6259,N_8124);
and U13954 (N_13954,N_9984,N_6928);
nor U13955 (N_13955,N_7908,N_8221);
or U13956 (N_13956,N_9901,N_6889);
nand U13957 (N_13957,N_7480,N_5666);
and U13958 (N_13958,N_8077,N_6878);
nand U13959 (N_13959,N_7659,N_7573);
nor U13960 (N_13960,N_9566,N_5048);
or U13961 (N_13961,N_7448,N_7304);
or U13962 (N_13962,N_8333,N_9207);
and U13963 (N_13963,N_9801,N_7900);
and U13964 (N_13964,N_9281,N_7998);
nand U13965 (N_13965,N_7559,N_5275);
or U13966 (N_13966,N_6825,N_6191);
nand U13967 (N_13967,N_8120,N_7251);
nand U13968 (N_13968,N_8482,N_6192);
nor U13969 (N_13969,N_5181,N_6704);
nand U13970 (N_13970,N_9401,N_9480);
nor U13971 (N_13971,N_9393,N_5313);
nor U13972 (N_13972,N_5142,N_5433);
and U13973 (N_13973,N_9507,N_6788);
nand U13974 (N_13974,N_5161,N_9634);
or U13975 (N_13975,N_8443,N_5897);
or U13976 (N_13976,N_5737,N_7862);
nand U13977 (N_13977,N_8676,N_5440);
nand U13978 (N_13978,N_8592,N_7341);
nand U13979 (N_13979,N_9096,N_8249);
and U13980 (N_13980,N_5380,N_8302);
nand U13981 (N_13981,N_5683,N_6894);
and U13982 (N_13982,N_6929,N_6063);
or U13983 (N_13983,N_9401,N_9728);
nor U13984 (N_13984,N_7799,N_6616);
and U13985 (N_13985,N_6786,N_7147);
nor U13986 (N_13986,N_8462,N_9620);
nor U13987 (N_13987,N_7230,N_5407);
or U13988 (N_13988,N_5230,N_5373);
xor U13989 (N_13989,N_6898,N_7925);
nor U13990 (N_13990,N_7081,N_7835);
nand U13991 (N_13991,N_7195,N_7356);
nor U13992 (N_13992,N_6937,N_6848);
nor U13993 (N_13993,N_7653,N_9149);
nand U13994 (N_13994,N_6929,N_5505);
or U13995 (N_13995,N_9570,N_9701);
nand U13996 (N_13996,N_7911,N_5315);
and U13997 (N_13997,N_6148,N_8350);
and U13998 (N_13998,N_9634,N_7461);
or U13999 (N_13999,N_9172,N_8596);
nor U14000 (N_14000,N_9780,N_5882);
nor U14001 (N_14001,N_7515,N_6889);
nor U14002 (N_14002,N_7706,N_9954);
and U14003 (N_14003,N_6097,N_6880);
or U14004 (N_14004,N_6443,N_6738);
or U14005 (N_14005,N_9023,N_5353);
nor U14006 (N_14006,N_9471,N_7864);
or U14007 (N_14007,N_6312,N_9951);
nor U14008 (N_14008,N_7573,N_8172);
nand U14009 (N_14009,N_5352,N_8329);
or U14010 (N_14010,N_9208,N_7492);
nand U14011 (N_14011,N_7369,N_8396);
nand U14012 (N_14012,N_5477,N_8736);
and U14013 (N_14013,N_7253,N_6383);
nand U14014 (N_14014,N_8907,N_5823);
nor U14015 (N_14015,N_6963,N_6734);
or U14016 (N_14016,N_5538,N_7461);
nand U14017 (N_14017,N_7467,N_7008);
nand U14018 (N_14018,N_7478,N_8277);
or U14019 (N_14019,N_6665,N_9834);
nor U14020 (N_14020,N_6772,N_8044);
and U14021 (N_14021,N_9416,N_5673);
nor U14022 (N_14022,N_7594,N_7382);
or U14023 (N_14023,N_5710,N_9442);
and U14024 (N_14024,N_7226,N_8823);
nand U14025 (N_14025,N_6657,N_6614);
or U14026 (N_14026,N_9969,N_6295);
or U14027 (N_14027,N_5720,N_5364);
and U14028 (N_14028,N_6666,N_8002);
nor U14029 (N_14029,N_9491,N_6304);
or U14030 (N_14030,N_9244,N_5830);
or U14031 (N_14031,N_8516,N_7199);
nand U14032 (N_14032,N_6647,N_8638);
nor U14033 (N_14033,N_9217,N_5850);
and U14034 (N_14034,N_6357,N_9797);
nor U14035 (N_14035,N_7112,N_8234);
and U14036 (N_14036,N_9664,N_5018);
or U14037 (N_14037,N_9297,N_7932);
or U14038 (N_14038,N_9135,N_6994);
nand U14039 (N_14039,N_7766,N_5558);
nand U14040 (N_14040,N_6650,N_5788);
nand U14041 (N_14041,N_9405,N_6448);
and U14042 (N_14042,N_9210,N_8034);
and U14043 (N_14043,N_5448,N_6658);
nand U14044 (N_14044,N_5142,N_6169);
nor U14045 (N_14045,N_5258,N_5103);
nor U14046 (N_14046,N_9793,N_9915);
nor U14047 (N_14047,N_6858,N_7578);
nand U14048 (N_14048,N_8467,N_7428);
and U14049 (N_14049,N_6025,N_8944);
or U14050 (N_14050,N_5953,N_9437);
nor U14051 (N_14051,N_9730,N_7399);
nand U14052 (N_14052,N_8870,N_7542);
nand U14053 (N_14053,N_7621,N_9364);
or U14054 (N_14054,N_6809,N_7242);
or U14055 (N_14055,N_9058,N_5912);
nand U14056 (N_14056,N_8021,N_7141);
nor U14057 (N_14057,N_5918,N_5289);
nand U14058 (N_14058,N_8055,N_8387);
or U14059 (N_14059,N_5925,N_6740);
nor U14060 (N_14060,N_7588,N_7871);
nand U14061 (N_14061,N_8686,N_7751);
nand U14062 (N_14062,N_9013,N_6089);
or U14063 (N_14063,N_6187,N_9921);
or U14064 (N_14064,N_6158,N_6886);
and U14065 (N_14065,N_8840,N_6894);
and U14066 (N_14066,N_5140,N_9246);
and U14067 (N_14067,N_9857,N_8089);
and U14068 (N_14068,N_7631,N_7867);
and U14069 (N_14069,N_5400,N_9317);
nand U14070 (N_14070,N_7505,N_5833);
nor U14071 (N_14071,N_8255,N_5597);
or U14072 (N_14072,N_6276,N_9520);
nor U14073 (N_14073,N_8876,N_8711);
nor U14074 (N_14074,N_5816,N_7718);
nand U14075 (N_14075,N_9594,N_5511);
or U14076 (N_14076,N_5402,N_5847);
and U14077 (N_14077,N_6265,N_6392);
or U14078 (N_14078,N_6352,N_7745);
nand U14079 (N_14079,N_5045,N_7981);
nor U14080 (N_14080,N_7844,N_7982);
and U14081 (N_14081,N_9318,N_5074);
and U14082 (N_14082,N_9550,N_5647);
nand U14083 (N_14083,N_8806,N_6950);
or U14084 (N_14084,N_8455,N_7508);
and U14085 (N_14085,N_8296,N_6835);
nor U14086 (N_14086,N_7975,N_5187);
nand U14087 (N_14087,N_9038,N_6736);
or U14088 (N_14088,N_8206,N_9050);
nor U14089 (N_14089,N_5891,N_8586);
or U14090 (N_14090,N_8858,N_9060);
or U14091 (N_14091,N_5938,N_8122);
nor U14092 (N_14092,N_8083,N_8714);
or U14093 (N_14093,N_6119,N_7016);
and U14094 (N_14094,N_6715,N_5803);
and U14095 (N_14095,N_9407,N_6326);
or U14096 (N_14096,N_9426,N_9986);
and U14097 (N_14097,N_6728,N_9754);
and U14098 (N_14098,N_7811,N_5206);
and U14099 (N_14099,N_7809,N_7733);
nor U14100 (N_14100,N_9157,N_6647);
or U14101 (N_14101,N_5615,N_6775);
nand U14102 (N_14102,N_5631,N_8259);
nand U14103 (N_14103,N_6377,N_5858);
nor U14104 (N_14104,N_5212,N_5931);
nand U14105 (N_14105,N_6448,N_5872);
and U14106 (N_14106,N_5972,N_7074);
or U14107 (N_14107,N_8198,N_6188);
nand U14108 (N_14108,N_5867,N_9889);
nand U14109 (N_14109,N_9151,N_5678);
nor U14110 (N_14110,N_8373,N_9229);
nor U14111 (N_14111,N_6951,N_5539);
or U14112 (N_14112,N_7540,N_8055);
or U14113 (N_14113,N_8296,N_7301);
nor U14114 (N_14114,N_6742,N_8294);
and U14115 (N_14115,N_5574,N_9073);
nor U14116 (N_14116,N_5804,N_5263);
nor U14117 (N_14117,N_7857,N_6676);
nand U14118 (N_14118,N_6524,N_7843);
and U14119 (N_14119,N_7931,N_8472);
and U14120 (N_14120,N_5793,N_7850);
nand U14121 (N_14121,N_9328,N_6882);
or U14122 (N_14122,N_8933,N_8628);
or U14123 (N_14123,N_7808,N_9909);
nand U14124 (N_14124,N_6846,N_9112);
nor U14125 (N_14125,N_8945,N_7398);
or U14126 (N_14126,N_7109,N_5094);
and U14127 (N_14127,N_8234,N_7510);
xor U14128 (N_14128,N_5455,N_6361);
or U14129 (N_14129,N_5702,N_6925);
and U14130 (N_14130,N_8575,N_8972);
or U14131 (N_14131,N_8471,N_6044);
nor U14132 (N_14132,N_5649,N_9602);
or U14133 (N_14133,N_5471,N_9988);
nand U14134 (N_14134,N_6001,N_7759);
nand U14135 (N_14135,N_7295,N_8783);
and U14136 (N_14136,N_9091,N_5984);
nor U14137 (N_14137,N_7433,N_9209);
nand U14138 (N_14138,N_5458,N_7162);
nand U14139 (N_14139,N_5696,N_8734);
nand U14140 (N_14140,N_6762,N_6690);
and U14141 (N_14141,N_6205,N_9164);
nand U14142 (N_14142,N_5274,N_7368);
nand U14143 (N_14143,N_6961,N_7789);
nand U14144 (N_14144,N_7457,N_8383);
and U14145 (N_14145,N_9531,N_7208);
nand U14146 (N_14146,N_5794,N_9489);
or U14147 (N_14147,N_9015,N_5121);
and U14148 (N_14148,N_6317,N_5302);
and U14149 (N_14149,N_5915,N_7897);
nand U14150 (N_14150,N_8814,N_6856);
nor U14151 (N_14151,N_8585,N_9422);
nand U14152 (N_14152,N_6757,N_6817);
nor U14153 (N_14153,N_5495,N_7855);
nor U14154 (N_14154,N_5118,N_5149);
or U14155 (N_14155,N_5625,N_9353);
nor U14156 (N_14156,N_9624,N_7256);
nand U14157 (N_14157,N_7351,N_7512);
and U14158 (N_14158,N_8485,N_7267);
nor U14159 (N_14159,N_5798,N_7666);
nand U14160 (N_14160,N_9920,N_6089);
nor U14161 (N_14161,N_5957,N_9471);
nor U14162 (N_14162,N_6732,N_5363);
nand U14163 (N_14163,N_5569,N_9488);
or U14164 (N_14164,N_8024,N_5849);
nand U14165 (N_14165,N_7945,N_6941);
or U14166 (N_14166,N_5057,N_6401);
nand U14167 (N_14167,N_8097,N_7606);
and U14168 (N_14168,N_6304,N_5943);
nor U14169 (N_14169,N_7385,N_9598);
nand U14170 (N_14170,N_6349,N_6137);
nand U14171 (N_14171,N_7100,N_8837);
nand U14172 (N_14172,N_7573,N_6759);
nor U14173 (N_14173,N_6624,N_9530);
nand U14174 (N_14174,N_8919,N_7405);
and U14175 (N_14175,N_6329,N_5029);
or U14176 (N_14176,N_9264,N_9861);
nand U14177 (N_14177,N_9671,N_8307);
nand U14178 (N_14178,N_8245,N_5442);
and U14179 (N_14179,N_6144,N_6067);
and U14180 (N_14180,N_7964,N_7487);
nand U14181 (N_14181,N_5978,N_9761);
nand U14182 (N_14182,N_8902,N_5634);
nor U14183 (N_14183,N_5469,N_5326);
or U14184 (N_14184,N_9092,N_9300);
and U14185 (N_14185,N_9686,N_7752);
nand U14186 (N_14186,N_9344,N_8349);
nand U14187 (N_14187,N_9221,N_8208);
nor U14188 (N_14188,N_5722,N_8781);
nand U14189 (N_14189,N_5201,N_9019);
nor U14190 (N_14190,N_5835,N_8413);
and U14191 (N_14191,N_5404,N_7506);
and U14192 (N_14192,N_7010,N_7507);
nor U14193 (N_14193,N_5676,N_5178);
nor U14194 (N_14194,N_8761,N_6848);
and U14195 (N_14195,N_5612,N_9875);
nor U14196 (N_14196,N_6948,N_7605);
nor U14197 (N_14197,N_8063,N_8334);
nor U14198 (N_14198,N_6246,N_5723);
nand U14199 (N_14199,N_7634,N_7414);
nor U14200 (N_14200,N_9031,N_7257);
nor U14201 (N_14201,N_6312,N_7307);
nor U14202 (N_14202,N_7768,N_9150);
nor U14203 (N_14203,N_7093,N_9947);
or U14204 (N_14204,N_7416,N_9227);
nand U14205 (N_14205,N_5836,N_5275);
nor U14206 (N_14206,N_5329,N_8057);
nand U14207 (N_14207,N_8114,N_9282);
nor U14208 (N_14208,N_6142,N_7806);
nor U14209 (N_14209,N_7779,N_5429);
and U14210 (N_14210,N_8577,N_5970);
nor U14211 (N_14211,N_7084,N_5743);
or U14212 (N_14212,N_8407,N_9147);
and U14213 (N_14213,N_6239,N_5487);
and U14214 (N_14214,N_7280,N_6308);
xnor U14215 (N_14215,N_9700,N_6146);
and U14216 (N_14216,N_7399,N_9423);
nand U14217 (N_14217,N_8793,N_9283);
and U14218 (N_14218,N_5896,N_9013);
or U14219 (N_14219,N_6602,N_5576);
and U14220 (N_14220,N_8276,N_5986);
or U14221 (N_14221,N_5461,N_7647);
and U14222 (N_14222,N_5206,N_7166);
nor U14223 (N_14223,N_8448,N_8122);
nor U14224 (N_14224,N_5199,N_5519);
and U14225 (N_14225,N_6755,N_9609);
or U14226 (N_14226,N_8000,N_9724);
and U14227 (N_14227,N_6547,N_6881);
nand U14228 (N_14228,N_5144,N_9806);
nand U14229 (N_14229,N_9699,N_5312);
and U14230 (N_14230,N_6017,N_5049);
nand U14231 (N_14231,N_6676,N_9242);
and U14232 (N_14232,N_6727,N_9217);
nor U14233 (N_14233,N_6457,N_6292);
and U14234 (N_14234,N_8696,N_5939);
and U14235 (N_14235,N_5417,N_7968);
and U14236 (N_14236,N_7932,N_7158);
and U14237 (N_14237,N_8846,N_6934);
nor U14238 (N_14238,N_5007,N_7222);
or U14239 (N_14239,N_6970,N_6979);
and U14240 (N_14240,N_6241,N_5576);
and U14241 (N_14241,N_6186,N_9030);
or U14242 (N_14242,N_9106,N_6761);
nor U14243 (N_14243,N_8691,N_9482);
and U14244 (N_14244,N_7263,N_8089);
nand U14245 (N_14245,N_7237,N_7340);
nand U14246 (N_14246,N_9815,N_7050);
and U14247 (N_14247,N_9410,N_7267);
and U14248 (N_14248,N_9546,N_5927);
and U14249 (N_14249,N_9448,N_7457);
and U14250 (N_14250,N_9862,N_8128);
nor U14251 (N_14251,N_7552,N_7307);
and U14252 (N_14252,N_8547,N_5164);
nor U14253 (N_14253,N_8861,N_8408);
and U14254 (N_14254,N_7503,N_7829);
nand U14255 (N_14255,N_7513,N_9662);
nand U14256 (N_14256,N_5215,N_6219);
and U14257 (N_14257,N_5821,N_6566);
nor U14258 (N_14258,N_5582,N_8482);
or U14259 (N_14259,N_6197,N_8063);
or U14260 (N_14260,N_8992,N_9459);
nor U14261 (N_14261,N_6813,N_9113);
and U14262 (N_14262,N_9039,N_7307);
and U14263 (N_14263,N_6789,N_5724);
nand U14264 (N_14264,N_8723,N_5435);
nor U14265 (N_14265,N_9073,N_5189);
and U14266 (N_14266,N_5312,N_7259);
nand U14267 (N_14267,N_9253,N_7630);
nand U14268 (N_14268,N_7720,N_8421);
nor U14269 (N_14269,N_7644,N_7525);
nand U14270 (N_14270,N_8185,N_9280);
and U14271 (N_14271,N_8445,N_7092);
or U14272 (N_14272,N_5520,N_8892);
or U14273 (N_14273,N_6763,N_6671);
nand U14274 (N_14274,N_5640,N_8810);
nand U14275 (N_14275,N_7690,N_8894);
nor U14276 (N_14276,N_7990,N_7548);
nor U14277 (N_14277,N_7680,N_8167);
and U14278 (N_14278,N_9749,N_7257);
nand U14279 (N_14279,N_5663,N_8547);
nand U14280 (N_14280,N_9146,N_7067);
nand U14281 (N_14281,N_9986,N_6755);
or U14282 (N_14282,N_9186,N_7147);
nand U14283 (N_14283,N_5299,N_6477);
nand U14284 (N_14284,N_6046,N_8145);
or U14285 (N_14285,N_8080,N_8925);
and U14286 (N_14286,N_8975,N_9503);
and U14287 (N_14287,N_7782,N_7285);
and U14288 (N_14288,N_6993,N_9083);
or U14289 (N_14289,N_7882,N_6074);
nand U14290 (N_14290,N_8697,N_6284);
or U14291 (N_14291,N_5118,N_9409);
nor U14292 (N_14292,N_5918,N_9568);
nor U14293 (N_14293,N_6600,N_5626);
nor U14294 (N_14294,N_6162,N_7212);
and U14295 (N_14295,N_8837,N_7617);
and U14296 (N_14296,N_8371,N_6553);
and U14297 (N_14297,N_5015,N_5073);
nand U14298 (N_14298,N_9913,N_8148);
nand U14299 (N_14299,N_7646,N_9215);
or U14300 (N_14300,N_5211,N_7133);
or U14301 (N_14301,N_8831,N_5418);
and U14302 (N_14302,N_5431,N_6110);
nor U14303 (N_14303,N_9227,N_6299);
nor U14304 (N_14304,N_8563,N_7383);
xnor U14305 (N_14305,N_7053,N_6606);
nor U14306 (N_14306,N_8842,N_5072);
nand U14307 (N_14307,N_9739,N_7153);
or U14308 (N_14308,N_7296,N_8205);
nor U14309 (N_14309,N_5312,N_9828);
and U14310 (N_14310,N_7124,N_8511);
nor U14311 (N_14311,N_6366,N_9546);
or U14312 (N_14312,N_6595,N_7374);
nand U14313 (N_14313,N_7791,N_9213);
or U14314 (N_14314,N_6947,N_5585);
nor U14315 (N_14315,N_5958,N_9326);
nor U14316 (N_14316,N_7788,N_9021);
and U14317 (N_14317,N_5354,N_6169);
and U14318 (N_14318,N_7777,N_7364);
or U14319 (N_14319,N_9942,N_6642);
and U14320 (N_14320,N_5929,N_9492);
or U14321 (N_14321,N_9514,N_5280);
and U14322 (N_14322,N_8091,N_6613);
and U14323 (N_14323,N_6700,N_9160);
nand U14324 (N_14324,N_7721,N_7789);
and U14325 (N_14325,N_6018,N_7103);
and U14326 (N_14326,N_7586,N_8284);
nand U14327 (N_14327,N_7336,N_8978);
and U14328 (N_14328,N_9040,N_9144);
or U14329 (N_14329,N_8415,N_8584);
and U14330 (N_14330,N_8128,N_8846);
nand U14331 (N_14331,N_8548,N_6553);
nand U14332 (N_14332,N_5422,N_6384);
nand U14333 (N_14333,N_7278,N_8271);
or U14334 (N_14334,N_5756,N_9926);
and U14335 (N_14335,N_8449,N_8399);
or U14336 (N_14336,N_8351,N_5892);
or U14337 (N_14337,N_8272,N_7378);
nand U14338 (N_14338,N_6048,N_6403);
and U14339 (N_14339,N_6095,N_9427);
nor U14340 (N_14340,N_7539,N_7301);
and U14341 (N_14341,N_6504,N_5920);
or U14342 (N_14342,N_7515,N_6211);
nor U14343 (N_14343,N_7171,N_6940);
nand U14344 (N_14344,N_5097,N_5126);
xnor U14345 (N_14345,N_5594,N_8462);
nor U14346 (N_14346,N_7672,N_7062);
nor U14347 (N_14347,N_7272,N_8110);
or U14348 (N_14348,N_9829,N_8705);
xor U14349 (N_14349,N_9541,N_5451);
nor U14350 (N_14350,N_9362,N_5510);
nand U14351 (N_14351,N_6946,N_8966);
nor U14352 (N_14352,N_8236,N_6928);
nor U14353 (N_14353,N_5215,N_7932);
and U14354 (N_14354,N_9127,N_7250);
and U14355 (N_14355,N_7722,N_6166);
nand U14356 (N_14356,N_7461,N_9997);
or U14357 (N_14357,N_6270,N_9184);
and U14358 (N_14358,N_6786,N_9419);
nor U14359 (N_14359,N_7648,N_7230);
nand U14360 (N_14360,N_6236,N_7319);
and U14361 (N_14361,N_6839,N_8127);
nand U14362 (N_14362,N_6698,N_5513);
xor U14363 (N_14363,N_6420,N_7760);
nand U14364 (N_14364,N_6953,N_6661);
nand U14365 (N_14365,N_9190,N_6512);
nand U14366 (N_14366,N_8952,N_6037);
or U14367 (N_14367,N_5617,N_9571);
nand U14368 (N_14368,N_7718,N_9545);
or U14369 (N_14369,N_9155,N_6623);
or U14370 (N_14370,N_7779,N_5010);
xor U14371 (N_14371,N_5522,N_8656);
and U14372 (N_14372,N_7578,N_8943);
nor U14373 (N_14373,N_9560,N_6196);
or U14374 (N_14374,N_6193,N_6436);
or U14375 (N_14375,N_5859,N_6531);
or U14376 (N_14376,N_6158,N_9764);
or U14377 (N_14377,N_8419,N_6493);
nand U14378 (N_14378,N_9390,N_9758);
nand U14379 (N_14379,N_5033,N_6943);
nand U14380 (N_14380,N_7337,N_8439);
and U14381 (N_14381,N_5425,N_9276);
or U14382 (N_14382,N_8476,N_9312);
nand U14383 (N_14383,N_8901,N_9774);
nand U14384 (N_14384,N_5824,N_6451);
or U14385 (N_14385,N_5726,N_5292);
nand U14386 (N_14386,N_9702,N_6211);
or U14387 (N_14387,N_5691,N_6151);
nor U14388 (N_14388,N_7491,N_7517);
and U14389 (N_14389,N_5137,N_7252);
or U14390 (N_14390,N_9014,N_6900);
or U14391 (N_14391,N_6660,N_6965);
and U14392 (N_14392,N_7250,N_7485);
nor U14393 (N_14393,N_7386,N_8901);
nor U14394 (N_14394,N_8893,N_8681);
and U14395 (N_14395,N_5932,N_8090);
nor U14396 (N_14396,N_5059,N_9079);
or U14397 (N_14397,N_5540,N_5535);
or U14398 (N_14398,N_7438,N_7774);
nor U14399 (N_14399,N_9870,N_8494);
nor U14400 (N_14400,N_7005,N_9929);
nor U14401 (N_14401,N_5562,N_7814);
nor U14402 (N_14402,N_8810,N_8514);
nand U14403 (N_14403,N_7994,N_9380);
and U14404 (N_14404,N_6727,N_6754);
and U14405 (N_14405,N_7095,N_5208);
and U14406 (N_14406,N_5139,N_6989);
nor U14407 (N_14407,N_7875,N_6604);
nor U14408 (N_14408,N_9014,N_5763);
nor U14409 (N_14409,N_8286,N_8391);
and U14410 (N_14410,N_9709,N_5135);
or U14411 (N_14411,N_8280,N_5434);
and U14412 (N_14412,N_7834,N_6165);
nor U14413 (N_14413,N_8590,N_6791);
nor U14414 (N_14414,N_9518,N_9204);
and U14415 (N_14415,N_5578,N_9963);
nand U14416 (N_14416,N_9903,N_7954);
nor U14417 (N_14417,N_9373,N_9333);
and U14418 (N_14418,N_5301,N_5646);
nor U14419 (N_14419,N_8849,N_9986);
nor U14420 (N_14420,N_8875,N_9602);
nor U14421 (N_14421,N_5389,N_8616);
and U14422 (N_14422,N_5156,N_9120);
and U14423 (N_14423,N_7759,N_5726);
or U14424 (N_14424,N_7198,N_5752);
nand U14425 (N_14425,N_6016,N_6775);
or U14426 (N_14426,N_5648,N_6435);
nand U14427 (N_14427,N_8606,N_6963);
nand U14428 (N_14428,N_6832,N_8950);
or U14429 (N_14429,N_7068,N_6574);
nand U14430 (N_14430,N_8873,N_7212);
or U14431 (N_14431,N_6186,N_8924);
and U14432 (N_14432,N_9738,N_5133);
or U14433 (N_14433,N_7515,N_8231);
nand U14434 (N_14434,N_7657,N_7479);
nand U14435 (N_14435,N_6026,N_9474);
nand U14436 (N_14436,N_6725,N_9294);
xnor U14437 (N_14437,N_6718,N_5523);
nor U14438 (N_14438,N_8856,N_5443);
nand U14439 (N_14439,N_7864,N_9633);
or U14440 (N_14440,N_8697,N_7087);
and U14441 (N_14441,N_8883,N_7334);
nand U14442 (N_14442,N_8536,N_5736);
nand U14443 (N_14443,N_7536,N_9093);
and U14444 (N_14444,N_7990,N_6874);
nor U14445 (N_14445,N_5091,N_5855);
nor U14446 (N_14446,N_9889,N_5675);
nor U14447 (N_14447,N_5253,N_8668);
or U14448 (N_14448,N_8895,N_8429);
or U14449 (N_14449,N_7216,N_9152);
and U14450 (N_14450,N_7820,N_9074);
nor U14451 (N_14451,N_5590,N_8908);
nand U14452 (N_14452,N_9396,N_8626);
or U14453 (N_14453,N_7953,N_6538);
and U14454 (N_14454,N_6171,N_5097);
nand U14455 (N_14455,N_5466,N_8774);
nor U14456 (N_14456,N_7530,N_8851);
nor U14457 (N_14457,N_7741,N_9013);
nand U14458 (N_14458,N_7880,N_9371);
nor U14459 (N_14459,N_5664,N_9555);
nor U14460 (N_14460,N_8654,N_6031);
or U14461 (N_14461,N_9952,N_9694);
nand U14462 (N_14462,N_9012,N_6992);
and U14463 (N_14463,N_7501,N_9761);
nor U14464 (N_14464,N_7467,N_7891);
or U14465 (N_14465,N_7559,N_9531);
and U14466 (N_14466,N_8427,N_8779);
or U14467 (N_14467,N_6747,N_6892);
or U14468 (N_14468,N_8029,N_7767);
nor U14469 (N_14469,N_5587,N_9451);
and U14470 (N_14470,N_5498,N_8890);
or U14471 (N_14471,N_6133,N_9629);
nand U14472 (N_14472,N_8416,N_9984);
or U14473 (N_14473,N_6040,N_7717);
or U14474 (N_14474,N_6767,N_6507);
xnor U14475 (N_14475,N_8197,N_6989);
nand U14476 (N_14476,N_5258,N_8391);
nand U14477 (N_14477,N_5930,N_5625);
or U14478 (N_14478,N_9632,N_6505);
nand U14479 (N_14479,N_8668,N_6641);
and U14480 (N_14480,N_7229,N_7225);
or U14481 (N_14481,N_7792,N_6165);
or U14482 (N_14482,N_7188,N_8025);
nor U14483 (N_14483,N_8183,N_8798);
or U14484 (N_14484,N_7886,N_8527);
or U14485 (N_14485,N_6957,N_9958);
or U14486 (N_14486,N_8816,N_5220);
nand U14487 (N_14487,N_5082,N_5003);
or U14488 (N_14488,N_5841,N_5664);
nand U14489 (N_14489,N_6397,N_8269);
or U14490 (N_14490,N_8421,N_6206);
nor U14491 (N_14491,N_8108,N_7339);
and U14492 (N_14492,N_7220,N_8535);
and U14493 (N_14493,N_9157,N_5627);
and U14494 (N_14494,N_9943,N_9493);
and U14495 (N_14495,N_5382,N_8073);
nand U14496 (N_14496,N_8485,N_5806);
nor U14497 (N_14497,N_9423,N_7724);
and U14498 (N_14498,N_7673,N_8280);
nor U14499 (N_14499,N_6564,N_9478);
and U14500 (N_14500,N_8015,N_8560);
nand U14501 (N_14501,N_9987,N_7624);
nor U14502 (N_14502,N_6545,N_7605);
or U14503 (N_14503,N_8284,N_6774);
or U14504 (N_14504,N_9305,N_9949);
nand U14505 (N_14505,N_7930,N_9691);
and U14506 (N_14506,N_9551,N_6961);
nand U14507 (N_14507,N_8306,N_7394);
nand U14508 (N_14508,N_8257,N_5066);
nor U14509 (N_14509,N_9726,N_5301);
or U14510 (N_14510,N_7131,N_7590);
and U14511 (N_14511,N_8176,N_6559);
and U14512 (N_14512,N_5641,N_5817);
nand U14513 (N_14513,N_7301,N_9735);
or U14514 (N_14514,N_9667,N_8752);
nor U14515 (N_14515,N_9781,N_5194);
and U14516 (N_14516,N_9136,N_7482);
nand U14517 (N_14517,N_5475,N_6153);
xnor U14518 (N_14518,N_7082,N_7718);
and U14519 (N_14519,N_5921,N_6984);
nor U14520 (N_14520,N_7470,N_9703);
or U14521 (N_14521,N_5084,N_5715);
nor U14522 (N_14522,N_6422,N_6328);
and U14523 (N_14523,N_7768,N_5602);
and U14524 (N_14524,N_8203,N_9143);
nand U14525 (N_14525,N_8911,N_9532);
nor U14526 (N_14526,N_9888,N_6689);
and U14527 (N_14527,N_8864,N_8242);
and U14528 (N_14528,N_6182,N_8774);
nor U14529 (N_14529,N_9920,N_7763);
nand U14530 (N_14530,N_7525,N_8416);
or U14531 (N_14531,N_7558,N_9683);
nand U14532 (N_14532,N_6042,N_6455);
or U14533 (N_14533,N_9386,N_9107);
xor U14534 (N_14534,N_8593,N_7337);
and U14535 (N_14535,N_6787,N_7068);
nand U14536 (N_14536,N_8005,N_5743);
xor U14537 (N_14537,N_9199,N_5868);
or U14538 (N_14538,N_5031,N_7229);
and U14539 (N_14539,N_7617,N_9035);
and U14540 (N_14540,N_9936,N_5976);
nand U14541 (N_14541,N_8198,N_7836);
or U14542 (N_14542,N_8633,N_5508);
and U14543 (N_14543,N_9437,N_8148);
and U14544 (N_14544,N_9369,N_9003);
or U14545 (N_14545,N_8104,N_5630);
nand U14546 (N_14546,N_9967,N_8398);
nand U14547 (N_14547,N_7549,N_7678);
nor U14548 (N_14548,N_7904,N_9606);
nor U14549 (N_14549,N_5590,N_9131);
nor U14550 (N_14550,N_5965,N_8533);
or U14551 (N_14551,N_5299,N_8375);
nor U14552 (N_14552,N_7422,N_9127);
nand U14553 (N_14553,N_6545,N_7196);
nor U14554 (N_14554,N_9548,N_9974);
nor U14555 (N_14555,N_9016,N_7157);
and U14556 (N_14556,N_6241,N_8591);
nand U14557 (N_14557,N_7352,N_5237);
or U14558 (N_14558,N_6543,N_7425);
or U14559 (N_14559,N_9553,N_9218);
nor U14560 (N_14560,N_6035,N_8364);
nand U14561 (N_14561,N_9815,N_6260);
nand U14562 (N_14562,N_5572,N_9191);
and U14563 (N_14563,N_9321,N_7875);
nor U14564 (N_14564,N_6598,N_6316);
nor U14565 (N_14565,N_8311,N_9878);
and U14566 (N_14566,N_5250,N_5188);
nor U14567 (N_14567,N_9518,N_7937);
nor U14568 (N_14568,N_6317,N_9959);
or U14569 (N_14569,N_7250,N_9555);
or U14570 (N_14570,N_9039,N_6320);
and U14571 (N_14571,N_6031,N_8128);
nor U14572 (N_14572,N_6341,N_8743);
or U14573 (N_14573,N_5527,N_9199);
nand U14574 (N_14574,N_9661,N_9606);
or U14575 (N_14575,N_5287,N_9895);
or U14576 (N_14576,N_7765,N_5719);
nor U14577 (N_14577,N_5645,N_6552);
nand U14578 (N_14578,N_9498,N_6613);
nand U14579 (N_14579,N_5991,N_8329);
nor U14580 (N_14580,N_8512,N_8233);
nand U14581 (N_14581,N_8171,N_7294);
nand U14582 (N_14582,N_5897,N_7392);
and U14583 (N_14583,N_9578,N_9720);
or U14584 (N_14584,N_5004,N_6099);
nand U14585 (N_14585,N_9174,N_9916);
nand U14586 (N_14586,N_9786,N_5260);
or U14587 (N_14587,N_9530,N_6172);
and U14588 (N_14588,N_7899,N_8979);
nor U14589 (N_14589,N_6412,N_9130);
nand U14590 (N_14590,N_6347,N_6505);
xor U14591 (N_14591,N_5063,N_8439);
or U14592 (N_14592,N_7750,N_5476);
nand U14593 (N_14593,N_7514,N_5120);
xnor U14594 (N_14594,N_8010,N_5356);
and U14595 (N_14595,N_5703,N_6108);
nor U14596 (N_14596,N_9845,N_5353);
and U14597 (N_14597,N_7313,N_6193);
or U14598 (N_14598,N_5036,N_7127);
and U14599 (N_14599,N_9986,N_7625);
nand U14600 (N_14600,N_5673,N_5341);
and U14601 (N_14601,N_9022,N_9098);
or U14602 (N_14602,N_7672,N_7210);
nand U14603 (N_14603,N_9523,N_6566);
or U14604 (N_14604,N_9662,N_6229);
or U14605 (N_14605,N_5065,N_8395);
nand U14606 (N_14606,N_5298,N_7552);
or U14607 (N_14607,N_7403,N_6667);
nand U14608 (N_14608,N_5490,N_7235);
and U14609 (N_14609,N_8811,N_9182);
or U14610 (N_14610,N_5921,N_6866);
nor U14611 (N_14611,N_8985,N_9125);
nor U14612 (N_14612,N_8487,N_6701);
or U14613 (N_14613,N_8812,N_6719);
or U14614 (N_14614,N_5621,N_9535);
or U14615 (N_14615,N_8515,N_7637);
and U14616 (N_14616,N_6352,N_9197);
nand U14617 (N_14617,N_8351,N_9609);
and U14618 (N_14618,N_7051,N_6905);
nand U14619 (N_14619,N_9853,N_9667);
nand U14620 (N_14620,N_9437,N_8815);
nand U14621 (N_14621,N_8362,N_9912);
and U14622 (N_14622,N_6762,N_8863);
nand U14623 (N_14623,N_6897,N_5624);
nor U14624 (N_14624,N_7840,N_7474);
nor U14625 (N_14625,N_9831,N_6951);
nor U14626 (N_14626,N_8031,N_9589);
nand U14627 (N_14627,N_5710,N_6452);
and U14628 (N_14628,N_7091,N_8276);
nor U14629 (N_14629,N_7606,N_6757);
nand U14630 (N_14630,N_9863,N_8768);
and U14631 (N_14631,N_5984,N_5306);
or U14632 (N_14632,N_8510,N_6926);
nand U14633 (N_14633,N_5075,N_6380);
or U14634 (N_14634,N_8118,N_9795);
or U14635 (N_14635,N_6395,N_9919);
nor U14636 (N_14636,N_8915,N_7013);
and U14637 (N_14637,N_9203,N_9666);
nor U14638 (N_14638,N_5404,N_7492);
nand U14639 (N_14639,N_6203,N_9843);
and U14640 (N_14640,N_9487,N_8129);
or U14641 (N_14641,N_8701,N_9249);
nor U14642 (N_14642,N_9161,N_9217);
and U14643 (N_14643,N_5627,N_6585);
or U14644 (N_14644,N_7143,N_5498);
or U14645 (N_14645,N_6176,N_9678);
or U14646 (N_14646,N_6273,N_7607);
and U14647 (N_14647,N_6895,N_6745);
nand U14648 (N_14648,N_9682,N_9030);
nor U14649 (N_14649,N_6262,N_8097);
or U14650 (N_14650,N_9634,N_5424);
nand U14651 (N_14651,N_9653,N_6691);
nor U14652 (N_14652,N_5831,N_9160);
nand U14653 (N_14653,N_8375,N_9501);
nor U14654 (N_14654,N_5176,N_7066);
and U14655 (N_14655,N_7910,N_7887);
nor U14656 (N_14656,N_9866,N_7051);
nor U14657 (N_14657,N_8450,N_8819);
and U14658 (N_14658,N_7228,N_9542);
nor U14659 (N_14659,N_5371,N_8754);
nor U14660 (N_14660,N_6421,N_8468);
nand U14661 (N_14661,N_6436,N_6637);
nand U14662 (N_14662,N_7711,N_9799);
or U14663 (N_14663,N_7775,N_9314);
nor U14664 (N_14664,N_9243,N_5395);
and U14665 (N_14665,N_6079,N_8652);
or U14666 (N_14666,N_5356,N_7944);
or U14667 (N_14667,N_7792,N_5190);
nor U14668 (N_14668,N_5949,N_9883);
nand U14669 (N_14669,N_5302,N_7411);
nor U14670 (N_14670,N_7829,N_9330);
or U14671 (N_14671,N_6119,N_7677);
and U14672 (N_14672,N_8934,N_6297);
nor U14673 (N_14673,N_7128,N_9298);
nand U14674 (N_14674,N_7591,N_5430);
nand U14675 (N_14675,N_9303,N_8373);
nor U14676 (N_14676,N_9646,N_8354);
nand U14677 (N_14677,N_7784,N_6608);
nor U14678 (N_14678,N_5402,N_9396);
nand U14679 (N_14679,N_8884,N_6650);
nor U14680 (N_14680,N_8317,N_8384);
or U14681 (N_14681,N_5694,N_8148);
nor U14682 (N_14682,N_9048,N_7073);
and U14683 (N_14683,N_9530,N_9277);
or U14684 (N_14684,N_9757,N_9354);
nand U14685 (N_14685,N_6556,N_5232);
nand U14686 (N_14686,N_8018,N_7710);
nand U14687 (N_14687,N_6339,N_9390);
nand U14688 (N_14688,N_6318,N_8482);
nor U14689 (N_14689,N_8505,N_8756);
and U14690 (N_14690,N_8956,N_7487);
nor U14691 (N_14691,N_6158,N_7657);
and U14692 (N_14692,N_5301,N_5583);
and U14693 (N_14693,N_6915,N_8060);
nand U14694 (N_14694,N_6385,N_7786);
nand U14695 (N_14695,N_9785,N_8168);
or U14696 (N_14696,N_5045,N_8053);
and U14697 (N_14697,N_7490,N_7353);
and U14698 (N_14698,N_6500,N_8553);
and U14699 (N_14699,N_7287,N_8160);
nand U14700 (N_14700,N_6868,N_9263);
nor U14701 (N_14701,N_9975,N_9692);
nor U14702 (N_14702,N_8098,N_5269);
or U14703 (N_14703,N_5854,N_5164);
nand U14704 (N_14704,N_8982,N_9952);
nor U14705 (N_14705,N_9499,N_8866);
nand U14706 (N_14706,N_8882,N_6164);
nor U14707 (N_14707,N_7672,N_9887);
or U14708 (N_14708,N_8951,N_7408);
nor U14709 (N_14709,N_5118,N_6787);
nand U14710 (N_14710,N_8978,N_7930);
or U14711 (N_14711,N_9501,N_9792);
or U14712 (N_14712,N_8787,N_7792);
or U14713 (N_14713,N_7931,N_7330);
and U14714 (N_14714,N_8232,N_9586);
and U14715 (N_14715,N_9146,N_7305);
nor U14716 (N_14716,N_7275,N_8339);
nor U14717 (N_14717,N_8325,N_7607);
nor U14718 (N_14718,N_5730,N_8900);
nand U14719 (N_14719,N_9254,N_7304);
nor U14720 (N_14720,N_9819,N_8330);
and U14721 (N_14721,N_8850,N_7292);
nor U14722 (N_14722,N_8020,N_9076);
or U14723 (N_14723,N_7510,N_9747);
and U14724 (N_14724,N_7396,N_5308);
or U14725 (N_14725,N_8316,N_7740);
or U14726 (N_14726,N_9017,N_8328);
nor U14727 (N_14727,N_8445,N_6481);
nor U14728 (N_14728,N_6404,N_9857);
nor U14729 (N_14729,N_9727,N_7031);
or U14730 (N_14730,N_9668,N_8513);
nor U14731 (N_14731,N_8246,N_6511);
or U14732 (N_14732,N_8041,N_9874);
or U14733 (N_14733,N_9491,N_5749);
or U14734 (N_14734,N_7736,N_7124);
and U14735 (N_14735,N_6440,N_5655);
or U14736 (N_14736,N_7876,N_8783);
or U14737 (N_14737,N_7076,N_5377);
or U14738 (N_14738,N_8382,N_7316);
or U14739 (N_14739,N_9273,N_9837);
nor U14740 (N_14740,N_5834,N_5294);
or U14741 (N_14741,N_9515,N_7595);
nor U14742 (N_14742,N_5975,N_8595);
nand U14743 (N_14743,N_8693,N_6936);
or U14744 (N_14744,N_7769,N_8524);
or U14745 (N_14745,N_8465,N_9417);
or U14746 (N_14746,N_8282,N_9298);
nor U14747 (N_14747,N_5176,N_9394);
nor U14748 (N_14748,N_5590,N_7642);
or U14749 (N_14749,N_7861,N_7246);
and U14750 (N_14750,N_9287,N_7805);
nor U14751 (N_14751,N_5106,N_8533);
and U14752 (N_14752,N_6009,N_5182);
and U14753 (N_14753,N_8533,N_6993);
nand U14754 (N_14754,N_7861,N_7046);
and U14755 (N_14755,N_5339,N_5449);
nand U14756 (N_14756,N_9633,N_5020);
nor U14757 (N_14757,N_7579,N_8426);
or U14758 (N_14758,N_8884,N_6156);
and U14759 (N_14759,N_8193,N_9262);
or U14760 (N_14760,N_5324,N_8480);
nor U14761 (N_14761,N_7811,N_8821);
or U14762 (N_14762,N_9483,N_8826);
nor U14763 (N_14763,N_8830,N_9005);
nor U14764 (N_14764,N_9131,N_7520);
and U14765 (N_14765,N_6099,N_6377);
or U14766 (N_14766,N_9815,N_5034);
and U14767 (N_14767,N_9828,N_8549);
nand U14768 (N_14768,N_5237,N_9693);
and U14769 (N_14769,N_9541,N_8938);
or U14770 (N_14770,N_9241,N_9234);
nor U14771 (N_14771,N_9966,N_8126);
or U14772 (N_14772,N_5175,N_5455);
nand U14773 (N_14773,N_9981,N_8583);
and U14774 (N_14774,N_8851,N_8060);
nand U14775 (N_14775,N_6147,N_9041);
or U14776 (N_14776,N_9966,N_5922);
nor U14777 (N_14777,N_8797,N_9690);
nor U14778 (N_14778,N_7832,N_5728);
and U14779 (N_14779,N_7884,N_7775);
nor U14780 (N_14780,N_6527,N_7307);
or U14781 (N_14781,N_6494,N_8829);
nand U14782 (N_14782,N_9826,N_8895);
or U14783 (N_14783,N_6366,N_6653);
nor U14784 (N_14784,N_7516,N_6618);
and U14785 (N_14785,N_7682,N_7557);
and U14786 (N_14786,N_6267,N_8766);
nor U14787 (N_14787,N_6453,N_8643);
nand U14788 (N_14788,N_9607,N_5109);
nand U14789 (N_14789,N_6029,N_8439);
nor U14790 (N_14790,N_5249,N_5202);
or U14791 (N_14791,N_8953,N_6612);
and U14792 (N_14792,N_9702,N_7980);
nor U14793 (N_14793,N_7844,N_6627);
nand U14794 (N_14794,N_7538,N_6283);
and U14795 (N_14795,N_6061,N_9080);
nand U14796 (N_14796,N_8732,N_9609);
and U14797 (N_14797,N_5615,N_5734);
nand U14798 (N_14798,N_9864,N_9108);
or U14799 (N_14799,N_8867,N_8556);
or U14800 (N_14800,N_6630,N_7852);
or U14801 (N_14801,N_6438,N_7607);
xor U14802 (N_14802,N_6412,N_5639);
nor U14803 (N_14803,N_6423,N_8243);
nand U14804 (N_14804,N_7260,N_7831);
nor U14805 (N_14805,N_5554,N_6990);
or U14806 (N_14806,N_7026,N_7792);
nand U14807 (N_14807,N_5931,N_5219);
or U14808 (N_14808,N_8738,N_8505);
or U14809 (N_14809,N_7398,N_6686);
and U14810 (N_14810,N_5542,N_9081);
nand U14811 (N_14811,N_9697,N_7706);
or U14812 (N_14812,N_6504,N_8813);
xnor U14813 (N_14813,N_6693,N_6265);
nor U14814 (N_14814,N_7405,N_8350);
nor U14815 (N_14815,N_9942,N_9013);
nand U14816 (N_14816,N_7793,N_9271);
nand U14817 (N_14817,N_7487,N_6813);
and U14818 (N_14818,N_5186,N_7637);
xor U14819 (N_14819,N_6385,N_7366);
or U14820 (N_14820,N_9881,N_7492);
and U14821 (N_14821,N_5987,N_7750);
nor U14822 (N_14822,N_5153,N_5882);
or U14823 (N_14823,N_5486,N_5541);
nor U14824 (N_14824,N_9234,N_7280);
and U14825 (N_14825,N_8973,N_9506);
nand U14826 (N_14826,N_9431,N_9444);
and U14827 (N_14827,N_9430,N_8511);
and U14828 (N_14828,N_7671,N_8402);
nor U14829 (N_14829,N_5598,N_6828);
nor U14830 (N_14830,N_8993,N_6705);
and U14831 (N_14831,N_9365,N_9081);
nor U14832 (N_14832,N_7268,N_9433);
nor U14833 (N_14833,N_9778,N_5710);
nand U14834 (N_14834,N_7643,N_5078);
and U14835 (N_14835,N_7924,N_9165);
or U14836 (N_14836,N_5808,N_9470);
and U14837 (N_14837,N_6004,N_8872);
nor U14838 (N_14838,N_5751,N_6201);
or U14839 (N_14839,N_5725,N_7800);
or U14840 (N_14840,N_5776,N_5382);
and U14841 (N_14841,N_8846,N_6660);
and U14842 (N_14842,N_8292,N_6037);
nor U14843 (N_14843,N_6542,N_8143);
nor U14844 (N_14844,N_6432,N_7064);
nand U14845 (N_14845,N_8403,N_7724);
or U14846 (N_14846,N_5038,N_5804);
and U14847 (N_14847,N_6079,N_8355);
or U14848 (N_14848,N_9018,N_5424);
nand U14849 (N_14849,N_6841,N_6011);
nand U14850 (N_14850,N_8920,N_5041);
nor U14851 (N_14851,N_7309,N_9386);
and U14852 (N_14852,N_9140,N_6544);
or U14853 (N_14853,N_9167,N_9523);
nand U14854 (N_14854,N_7512,N_7694);
and U14855 (N_14855,N_8603,N_9324);
nor U14856 (N_14856,N_5839,N_6710);
nand U14857 (N_14857,N_7358,N_5915);
and U14858 (N_14858,N_5643,N_8077);
nor U14859 (N_14859,N_9675,N_9324);
and U14860 (N_14860,N_7579,N_8131);
or U14861 (N_14861,N_9140,N_8982);
and U14862 (N_14862,N_6285,N_5399);
nor U14863 (N_14863,N_9515,N_6132);
and U14864 (N_14864,N_5296,N_7563);
or U14865 (N_14865,N_5345,N_5149);
nand U14866 (N_14866,N_9034,N_7217);
nor U14867 (N_14867,N_5875,N_5487);
nand U14868 (N_14868,N_9111,N_9772);
nand U14869 (N_14869,N_7020,N_5999);
and U14870 (N_14870,N_8721,N_6076);
nor U14871 (N_14871,N_5420,N_9060);
nor U14872 (N_14872,N_8733,N_8408);
and U14873 (N_14873,N_5676,N_8073);
nor U14874 (N_14874,N_6884,N_7600);
or U14875 (N_14875,N_9588,N_5073);
or U14876 (N_14876,N_5826,N_8251);
or U14877 (N_14877,N_9460,N_7499);
nor U14878 (N_14878,N_6606,N_7770);
or U14879 (N_14879,N_5718,N_8395);
nand U14880 (N_14880,N_6600,N_9662);
nand U14881 (N_14881,N_7076,N_5610);
and U14882 (N_14882,N_6700,N_9032);
nand U14883 (N_14883,N_8104,N_9531);
nor U14884 (N_14884,N_6370,N_5171);
nand U14885 (N_14885,N_8946,N_9196);
nand U14886 (N_14886,N_9771,N_9894);
and U14887 (N_14887,N_9593,N_7662);
and U14888 (N_14888,N_6408,N_8563);
nand U14889 (N_14889,N_8144,N_7186);
nand U14890 (N_14890,N_6490,N_7715);
or U14891 (N_14891,N_8083,N_9068);
nor U14892 (N_14892,N_5818,N_9691);
or U14893 (N_14893,N_7652,N_6615);
nor U14894 (N_14894,N_7773,N_8172);
nand U14895 (N_14895,N_7532,N_8027);
and U14896 (N_14896,N_7204,N_8034);
and U14897 (N_14897,N_7798,N_6131);
nor U14898 (N_14898,N_7056,N_5305);
nor U14899 (N_14899,N_6891,N_9992);
and U14900 (N_14900,N_7614,N_7569);
and U14901 (N_14901,N_6132,N_8488);
and U14902 (N_14902,N_9354,N_7723);
nor U14903 (N_14903,N_7936,N_6831);
nand U14904 (N_14904,N_6757,N_5806);
or U14905 (N_14905,N_9027,N_7133);
nor U14906 (N_14906,N_5076,N_6317);
and U14907 (N_14907,N_9886,N_5075);
and U14908 (N_14908,N_9157,N_5743);
nor U14909 (N_14909,N_8796,N_5756);
or U14910 (N_14910,N_9912,N_7395);
or U14911 (N_14911,N_7270,N_7403);
or U14912 (N_14912,N_6934,N_6940);
or U14913 (N_14913,N_5458,N_8460);
or U14914 (N_14914,N_7208,N_6480);
nand U14915 (N_14915,N_8648,N_9349);
nor U14916 (N_14916,N_6134,N_6348);
nand U14917 (N_14917,N_7161,N_6051);
and U14918 (N_14918,N_8890,N_7258);
or U14919 (N_14919,N_9390,N_9886);
nor U14920 (N_14920,N_8931,N_6122);
and U14921 (N_14921,N_9888,N_8477);
or U14922 (N_14922,N_8118,N_9331);
or U14923 (N_14923,N_8753,N_6803);
and U14924 (N_14924,N_9627,N_5783);
nand U14925 (N_14925,N_8698,N_8433);
nand U14926 (N_14926,N_5827,N_8210);
nor U14927 (N_14927,N_5287,N_9461);
or U14928 (N_14928,N_6773,N_6694);
nand U14929 (N_14929,N_6792,N_9810);
or U14930 (N_14930,N_9641,N_5968);
nor U14931 (N_14931,N_7015,N_8642);
or U14932 (N_14932,N_9441,N_7968);
and U14933 (N_14933,N_5588,N_6066);
nor U14934 (N_14934,N_5477,N_7015);
nor U14935 (N_14935,N_5835,N_5283);
and U14936 (N_14936,N_5560,N_6855);
nor U14937 (N_14937,N_6096,N_8231);
nor U14938 (N_14938,N_6758,N_7191);
and U14939 (N_14939,N_7323,N_9074);
or U14940 (N_14940,N_6634,N_9222);
nor U14941 (N_14941,N_9134,N_5720);
nand U14942 (N_14942,N_9697,N_9180);
nor U14943 (N_14943,N_6315,N_6805);
nand U14944 (N_14944,N_7242,N_9283);
or U14945 (N_14945,N_7868,N_9710);
or U14946 (N_14946,N_5217,N_8678);
xor U14947 (N_14947,N_5323,N_9721);
nand U14948 (N_14948,N_5729,N_8621);
nand U14949 (N_14949,N_8187,N_6686);
nand U14950 (N_14950,N_7437,N_7066);
nand U14951 (N_14951,N_7135,N_6995);
nand U14952 (N_14952,N_6864,N_9140);
or U14953 (N_14953,N_5304,N_5831);
and U14954 (N_14954,N_6124,N_8972);
and U14955 (N_14955,N_9282,N_8258);
or U14956 (N_14956,N_5932,N_7400);
and U14957 (N_14957,N_8588,N_7627);
nor U14958 (N_14958,N_8509,N_7849);
and U14959 (N_14959,N_5290,N_9411);
and U14960 (N_14960,N_7051,N_9371);
or U14961 (N_14961,N_6257,N_8391);
and U14962 (N_14962,N_5524,N_9781);
or U14963 (N_14963,N_7629,N_7998);
nand U14964 (N_14964,N_5480,N_9333);
or U14965 (N_14965,N_8560,N_8718);
and U14966 (N_14966,N_6814,N_7670);
nor U14967 (N_14967,N_6787,N_5421);
nor U14968 (N_14968,N_5414,N_5652);
or U14969 (N_14969,N_6463,N_9363);
and U14970 (N_14970,N_6760,N_6236);
nor U14971 (N_14971,N_6762,N_6198);
and U14972 (N_14972,N_6838,N_8702);
nand U14973 (N_14973,N_6876,N_7219);
nand U14974 (N_14974,N_7196,N_9289);
or U14975 (N_14975,N_8672,N_8640);
and U14976 (N_14976,N_5485,N_7917);
or U14977 (N_14977,N_6711,N_7272);
nand U14978 (N_14978,N_9718,N_7459);
xnor U14979 (N_14979,N_6635,N_9332);
or U14980 (N_14980,N_6836,N_6390);
or U14981 (N_14981,N_6817,N_7849);
or U14982 (N_14982,N_5316,N_6050);
and U14983 (N_14983,N_9104,N_6327);
and U14984 (N_14984,N_6324,N_9137);
and U14985 (N_14985,N_8796,N_8638);
xor U14986 (N_14986,N_9890,N_8166);
nor U14987 (N_14987,N_6966,N_5351);
nand U14988 (N_14988,N_5252,N_9872);
or U14989 (N_14989,N_8097,N_7947);
nor U14990 (N_14990,N_7990,N_8010);
nand U14991 (N_14991,N_6609,N_6530);
or U14992 (N_14992,N_7740,N_6751);
nand U14993 (N_14993,N_8139,N_6094);
nand U14994 (N_14994,N_7951,N_6877);
nor U14995 (N_14995,N_8485,N_8205);
nand U14996 (N_14996,N_6047,N_8321);
nor U14997 (N_14997,N_7800,N_9690);
nand U14998 (N_14998,N_6053,N_5475);
nor U14999 (N_14999,N_5997,N_6183);
nor UO_0 (O_0,N_10435,N_12880);
or UO_1 (O_1,N_13568,N_12339);
nand UO_2 (O_2,N_12508,N_10779);
nand UO_3 (O_3,N_14176,N_10524);
or UO_4 (O_4,N_10816,N_11690);
nand UO_5 (O_5,N_10665,N_10152);
nand UO_6 (O_6,N_12686,N_11276);
or UO_7 (O_7,N_11491,N_13930);
or UO_8 (O_8,N_12451,N_10089);
nor UO_9 (O_9,N_14611,N_10990);
and UO_10 (O_10,N_10142,N_11445);
or UO_11 (O_11,N_12008,N_11708);
nor UO_12 (O_12,N_12479,N_10730);
or UO_13 (O_13,N_13501,N_14454);
nand UO_14 (O_14,N_12531,N_12990);
nor UO_15 (O_15,N_11751,N_13510);
or UO_16 (O_16,N_12722,N_11755);
nor UO_17 (O_17,N_11669,N_13609);
nand UO_18 (O_18,N_12375,N_14023);
nand UO_19 (O_19,N_12678,N_13406);
nor UO_20 (O_20,N_12675,N_13239);
and UO_21 (O_21,N_14047,N_14579);
nand UO_22 (O_22,N_14029,N_14581);
nand UO_23 (O_23,N_10335,N_11726);
nand UO_24 (O_24,N_13646,N_14988);
or UO_25 (O_25,N_12510,N_12632);
or UO_26 (O_26,N_10925,N_12007);
or UO_27 (O_27,N_11457,N_14106);
nand UO_28 (O_28,N_12391,N_11737);
nor UO_29 (O_29,N_14757,N_12061);
nand UO_30 (O_30,N_12355,N_13002);
or UO_31 (O_31,N_10347,N_10204);
nor UO_32 (O_32,N_10353,N_14823);
and UO_33 (O_33,N_14278,N_10500);
and UO_34 (O_34,N_12025,N_11480);
or UO_35 (O_35,N_13608,N_14496);
or UO_36 (O_36,N_11487,N_14478);
and UO_37 (O_37,N_13348,N_14596);
or UO_38 (O_38,N_11113,N_11109);
nand UO_39 (O_39,N_14699,N_10520);
and UO_40 (O_40,N_10140,N_10410);
and UO_41 (O_41,N_14881,N_10162);
and UO_42 (O_42,N_14162,N_11412);
and UO_43 (O_43,N_14840,N_10409);
nor UO_44 (O_44,N_10422,N_11250);
nand UO_45 (O_45,N_14769,N_14531);
nand UO_46 (O_46,N_12096,N_14755);
nor UO_47 (O_47,N_12644,N_10749);
and UO_48 (O_48,N_12705,N_13289);
or UO_49 (O_49,N_14366,N_14097);
nand UO_50 (O_50,N_13952,N_12081);
and UO_51 (O_51,N_13386,N_13889);
and UO_52 (O_52,N_10436,N_14316);
or UO_53 (O_53,N_11279,N_12165);
nor UO_54 (O_54,N_11333,N_11204);
nor UO_55 (O_55,N_14244,N_11811);
nor UO_56 (O_56,N_14020,N_12435);
nand UO_57 (O_57,N_11927,N_11256);
nor UO_58 (O_58,N_14888,N_11298);
and UO_59 (O_59,N_11285,N_10263);
nor UO_60 (O_60,N_14400,N_10589);
and UO_61 (O_61,N_14975,N_10931);
nand UO_62 (O_62,N_12643,N_14025);
nor UO_63 (O_63,N_10359,N_14367);
nor UO_64 (O_64,N_11799,N_11073);
and UO_65 (O_65,N_14335,N_12489);
nand UO_66 (O_66,N_12604,N_12297);
or UO_67 (O_67,N_11240,N_13718);
nor UO_68 (O_68,N_11676,N_14433);
or UO_69 (O_69,N_14756,N_14657);
nor UO_70 (O_70,N_12173,N_13325);
and UO_71 (O_71,N_12905,N_13792);
and UO_72 (O_72,N_12517,N_12579);
and UO_73 (O_73,N_12665,N_13147);
or UO_74 (O_74,N_11000,N_11785);
or UO_75 (O_75,N_13059,N_14659);
and UO_76 (O_76,N_14820,N_11937);
or UO_77 (O_77,N_13920,N_10293);
and UO_78 (O_78,N_10241,N_12121);
nand UO_79 (O_79,N_14908,N_12129);
nor UO_80 (O_80,N_13111,N_11167);
or UO_81 (O_81,N_14224,N_10228);
nor UO_82 (O_82,N_14718,N_12284);
nand UO_83 (O_83,N_12878,N_10016);
or UO_84 (O_84,N_10010,N_13363);
nand UO_85 (O_85,N_11241,N_14972);
or UO_86 (O_86,N_11053,N_10901);
or UO_87 (O_87,N_14222,N_13192);
and UO_88 (O_88,N_11354,N_10291);
or UO_89 (O_89,N_14683,N_13915);
nor UO_90 (O_90,N_10394,N_11035);
nor UO_91 (O_91,N_11527,N_10273);
and UO_92 (O_92,N_12358,N_14515);
nand UO_93 (O_93,N_13996,N_10610);
and UO_94 (O_94,N_12866,N_10547);
nor UO_95 (O_95,N_12820,N_10604);
and UO_96 (O_96,N_10736,N_11237);
nor UO_97 (O_97,N_11482,N_11492);
and UO_98 (O_98,N_12023,N_13546);
nand UO_99 (O_99,N_10629,N_13799);
nand UO_100 (O_100,N_14185,N_12901);
nor UO_101 (O_101,N_11621,N_13193);
or UO_102 (O_102,N_10586,N_11779);
nor UO_103 (O_103,N_12246,N_13019);
nand UO_104 (O_104,N_13940,N_12271);
or UO_105 (O_105,N_11086,N_12563);
nor UO_106 (O_106,N_10402,N_13218);
nor UO_107 (O_107,N_10747,N_11414);
and UO_108 (O_108,N_11627,N_13808);
nor UO_109 (O_109,N_14261,N_11586);
nand UO_110 (O_110,N_10956,N_10888);
nor UO_111 (O_111,N_14548,N_13993);
nor UO_112 (O_112,N_11367,N_10783);
and UO_113 (O_113,N_14050,N_12884);
nand UO_114 (O_114,N_13999,N_13012);
nand UO_115 (O_115,N_10835,N_14605);
nand UO_116 (O_116,N_11997,N_11008);
or UO_117 (O_117,N_10302,N_10416);
or UO_118 (O_118,N_11743,N_13252);
or UO_119 (O_119,N_12960,N_12306);
and UO_120 (O_120,N_13593,N_11775);
or UO_121 (O_121,N_11433,N_11582);
and UO_122 (O_122,N_13702,N_10337);
or UO_123 (O_123,N_14110,N_10451);
xnor UO_124 (O_124,N_14502,N_13944);
and UO_125 (O_125,N_14633,N_13281);
nand UO_126 (O_126,N_11715,N_12337);
nor UO_127 (O_127,N_10289,N_10066);
nand UO_128 (O_128,N_14951,N_14242);
and UO_129 (O_129,N_12349,N_11254);
and UO_130 (O_130,N_12608,N_13500);
and UO_131 (O_131,N_10120,N_11233);
nand UO_132 (O_132,N_11520,N_10671);
nand UO_133 (O_133,N_10499,N_10275);
nor UO_134 (O_134,N_14814,N_11837);
nand UO_135 (O_135,N_12663,N_13732);
or UO_136 (O_136,N_13404,N_13277);
or UO_137 (O_137,N_12591,N_11385);
or UO_138 (O_138,N_14929,N_10576);
and UO_139 (O_139,N_11474,N_13734);
or UO_140 (O_140,N_14594,N_11776);
nand UO_141 (O_141,N_11853,N_12917);
and UO_142 (O_142,N_10578,N_11805);
and UO_143 (O_143,N_12017,N_13956);
and UO_144 (O_144,N_10869,N_13575);
or UO_145 (O_145,N_12352,N_12595);
or UO_146 (O_146,N_13443,N_11056);
or UO_147 (O_147,N_12660,N_13382);
nor UO_148 (O_148,N_14737,N_10488);
and UO_149 (O_149,N_13463,N_13138);
or UO_150 (O_150,N_13290,N_13372);
nand UO_151 (O_151,N_12412,N_13830);
nand UO_152 (O_152,N_14290,N_12523);
and UO_153 (O_153,N_11691,N_13592);
nor UO_154 (O_154,N_13384,N_14696);
nand UO_155 (O_155,N_11484,N_14318);
and UO_156 (O_156,N_13742,N_14093);
and UO_157 (O_157,N_12806,N_13376);
or UO_158 (O_158,N_12389,N_11351);
nor UO_159 (O_159,N_14917,N_14187);
or UO_160 (O_160,N_12743,N_11835);
nor UO_161 (O_161,N_13194,N_11659);
nor UO_162 (O_162,N_13211,N_14810);
nand UO_163 (O_163,N_13369,N_14918);
nor UO_164 (O_164,N_11666,N_14295);
nand UO_165 (O_165,N_11136,N_13445);
or UO_166 (O_166,N_14781,N_10360);
nand UO_167 (O_167,N_12317,N_13246);
nor UO_168 (O_168,N_10075,N_11894);
or UO_169 (O_169,N_14248,N_10766);
nor UO_170 (O_170,N_12461,N_10542);
nor UO_171 (O_171,N_13144,N_12252);
or UO_172 (O_172,N_13954,N_12243);
nor UO_173 (O_173,N_11982,N_11009);
and UO_174 (O_174,N_11832,N_11983);
and UO_175 (O_175,N_10452,N_11312);
or UO_176 (O_176,N_11704,N_10770);
nand UO_177 (O_177,N_12761,N_12739);
nor UO_178 (O_178,N_10174,N_12970);
nor UO_179 (O_179,N_11922,N_14450);
and UO_180 (O_180,N_10019,N_11038);
nor UO_181 (O_181,N_10871,N_14872);
nand UO_182 (O_182,N_10808,N_14526);
nand UO_183 (O_183,N_12215,N_13370);
and UO_184 (O_184,N_12609,N_12456);
nor UO_185 (O_185,N_13397,N_14382);
nand UO_186 (O_186,N_12377,N_10294);
and UO_187 (O_187,N_13971,N_14505);
nand UO_188 (O_188,N_10419,N_11738);
nor UO_189 (O_189,N_11398,N_13907);
nor UO_190 (O_190,N_13823,N_14252);
or UO_191 (O_191,N_12431,N_11514);
nand UO_192 (O_192,N_12589,N_11238);
or UO_193 (O_193,N_11848,N_10205);
nand UO_194 (O_194,N_10717,N_10048);
and UO_195 (O_195,N_14983,N_14238);
nand UO_196 (O_196,N_11323,N_14472);
or UO_197 (O_197,N_12285,N_10509);
nor UO_198 (O_198,N_11375,N_12136);
nand UO_199 (O_199,N_10992,N_14161);
or UO_200 (O_200,N_12583,N_10765);
nand UO_201 (O_201,N_10916,N_12372);
and UO_202 (O_202,N_10407,N_10200);
nor UO_203 (O_203,N_11089,N_11419);
or UO_204 (O_204,N_10919,N_13033);
or UO_205 (O_205,N_14939,N_11470);
nor UO_206 (O_206,N_10180,N_11325);
or UO_207 (O_207,N_14671,N_10071);
nor UO_208 (O_208,N_11609,N_12718);
or UO_209 (O_209,N_13197,N_11155);
or UO_210 (O_210,N_13673,N_10687);
nor UO_211 (O_211,N_11060,N_13894);
nand UO_212 (O_212,N_10889,N_14417);
nor UO_213 (O_213,N_11243,N_11189);
nor UO_214 (O_214,N_10366,N_14650);
nor UO_215 (O_215,N_14119,N_14285);
nor UO_216 (O_216,N_13577,N_12657);
and UO_217 (O_217,N_11436,N_13648);
nor UO_218 (O_218,N_12757,N_10978);
nand UO_219 (O_219,N_13474,N_13735);
nand UO_220 (O_220,N_11761,N_10083);
nor UO_221 (O_221,N_12942,N_10232);
nor UO_222 (O_222,N_10530,N_13403);
or UO_223 (O_223,N_12336,N_14172);
nor UO_224 (O_224,N_11526,N_11045);
nand UO_225 (O_225,N_13805,N_13900);
or UO_226 (O_226,N_11230,N_13257);
and UO_227 (O_227,N_13263,N_13773);
nand UO_228 (O_228,N_14432,N_11064);
or UO_229 (O_229,N_11663,N_12505);
nor UO_230 (O_230,N_12142,N_14443);
or UO_231 (O_231,N_13366,N_10713);
nand UO_232 (O_232,N_11022,N_14114);
and UO_233 (O_233,N_14070,N_13630);
nand UO_234 (O_234,N_10601,N_10179);
or UO_235 (O_235,N_13824,N_12645);
and UO_236 (O_236,N_14049,N_13662);
nand UO_237 (O_237,N_14036,N_12842);
and UO_238 (O_238,N_11332,N_13583);
and UO_239 (O_239,N_11773,N_12498);
nand UO_240 (O_240,N_14901,N_11786);
and UO_241 (O_241,N_12185,N_13187);
or UO_242 (O_242,N_13628,N_13417);
or UO_243 (O_243,N_10572,N_10677);
nand UO_244 (O_244,N_13846,N_12350);
nor UO_245 (O_245,N_12500,N_12790);
or UO_246 (O_246,N_13330,N_11075);
nand UO_247 (O_247,N_11434,N_12259);
nand UO_248 (O_248,N_14747,N_12216);
nand UO_249 (O_249,N_11636,N_14619);
or UO_250 (O_250,N_11464,N_10235);
and UO_251 (O_251,N_12378,N_10989);
and UO_252 (O_252,N_13795,N_12035);
nor UO_253 (O_253,N_11529,N_13709);
and UO_254 (O_254,N_13763,N_11789);
and UO_255 (O_255,N_10627,N_13431);
nor UO_256 (O_256,N_12810,N_13396);
and UO_257 (O_257,N_10033,N_13292);
nor UO_258 (O_258,N_12405,N_11424);
nor UO_259 (O_259,N_10065,N_12574);
nand UO_260 (O_260,N_12542,N_12445);
nor UO_261 (O_261,N_11163,N_13635);
and UO_262 (O_262,N_11320,N_10551);
nor UO_263 (O_263,N_14039,N_11069);
or UO_264 (O_264,N_10026,N_11407);
nand UO_265 (O_265,N_14796,N_10073);
nand UO_266 (O_266,N_12824,N_10350);
nand UO_267 (O_267,N_13333,N_14380);
and UO_268 (O_268,N_13442,N_13833);
or UO_269 (O_269,N_11680,N_10467);
and UO_270 (O_270,N_11742,N_13522);
and UO_271 (O_271,N_10288,N_13477);
nor UO_272 (O_272,N_14199,N_10534);
or UO_273 (O_273,N_12898,N_11130);
or UO_274 (O_274,N_11754,N_13137);
nand UO_275 (O_275,N_14846,N_10039);
and UO_276 (O_276,N_13109,N_12545);
or UO_277 (O_277,N_14542,N_11435);
nand UO_278 (O_278,N_13615,N_12254);
or UO_279 (O_279,N_11865,N_13312);
and UO_280 (O_280,N_11287,N_13960);
or UO_281 (O_281,N_13625,N_11536);
or UO_282 (O_282,N_13199,N_13004);
nor UO_283 (O_283,N_11843,N_10119);
and UO_284 (O_284,N_11483,N_13320);
or UO_285 (O_285,N_13947,N_10744);
or UO_286 (O_286,N_13746,N_14758);
xnor UO_287 (O_287,N_11215,N_10003);
and UO_288 (O_288,N_14628,N_10845);
nor UO_289 (O_289,N_14546,N_14639);
nand UO_290 (O_290,N_14809,N_11990);
nor UO_291 (O_291,N_11423,N_14326);
nand UO_292 (O_292,N_13255,N_13184);
nor UO_293 (O_293,N_11639,N_11314);
nor UO_294 (O_294,N_14640,N_14071);
and UO_295 (O_295,N_13994,N_10833);
and UO_296 (O_296,N_11583,N_12894);
nand UO_297 (O_297,N_12039,N_10902);
or UO_298 (O_298,N_13007,N_12274);
nand UO_299 (O_299,N_14600,N_12200);
or UO_300 (O_300,N_10387,N_12487);
nor UO_301 (O_301,N_14419,N_13280);
or UO_302 (O_302,N_12698,N_11833);
or UO_303 (O_303,N_14506,N_11471);
and UO_304 (O_304,N_12114,N_13943);
nor UO_305 (O_305,N_13741,N_14572);
or UO_306 (O_306,N_10683,N_12813);
and UO_307 (O_307,N_13173,N_11784);
nor UO_308 (O_308,N_10169,N_14456);
nand UO_309 (O_309,N_14006,N_12615);
or UO_310 (O_310,N_12852,N_10151);
and UO_311 (O_311,N_12086,N_11970);
and UO_312 (O_312,N_14276,N_12839);
nand UO_313 (O_313,N_14903,N_13284);
nand UO_314 (O_314,N_14484,N_11643);
nand UO_315 (O_315,N_12991,N_13163);
and UO_316 (O_316,N_10042,N_11037);
or UO_317 (O_317,N_13306,N_11846);
or UO_318 (O_318,N_11186,N_14815);
nor UO_319 (O_319,N_12703,N_11386);
or UO_320 (O_320,N_10655,N_10389);
or UO_321 (O_321,N_13326,N_10094);
or UO_322 (O_322,N_10706,N_14632);
and UO_323 (O_323,N_12413,N_14653);
nand UO_324 (O_324,N_11615,N_12881);
or UO_325 (O_325,N_14919,N_14794);
and UO_326 (O_326,N_11548,N_14381);
or UO_327 (O_327,N_13948,N_14100);
nand UO_328 (O_328,N_13261,N_13722);
nand UO_329 (O_329,N_11402,N_14943);
nor UO_330 (O_330,N_12571,N_11898);
nand UO_331 (O_331,N_10946,N_14587);
and UO_332 (O_332,N_13549,N_13119);
or UO_333 (O_333,N_12631,N_10050);
and UO_334 (O_334,N_10987,N_13975);
nor UO_335 (O_335,N_11809,N_12930);
and UO_336 (O_336,N_11866,N_13832);
or UO_337 (O_337,N_11216,N_11498);
nor UO_338 (O_338,N_11503,N_12829);
nor UO_339 (O_339,N_10274,N_12734);
or UO_340 (O_340,N_12276,N_14524);
or UO_341 (O_341,N_12731,N_10260);
and UO_342 (O_342,N_11379,N_14841);
or UO_343 (O_343,N_14974,N_10093);
nand UO_344 (O_344,N_14338,N_12834);
nand UO_345 (O_345,N_11309,N_10914);
or UO_346 (O_346,N_13053,N_13989);
and UO_347 (O_347,N_12776,N_11284);
nand UO_348 (O_348,N_14179,N_12701);
nand UO_349 (O_349,N_12573,N_14759);
nand UO_350 (O_350,N_11569,N_12109);
and UO_351 (O_351,N_10265,N_12626);
nor UO_352 (O_352,N_13991,N_13440);
and UO_353 (O_353,N_13169,N_12194);
nand UO_354 (O_354,N_11652,N_14314);
and UO_355 (O_355,N_11018,N_10025);
or UO_356 (O_356,N_14453,N_14607);
and UO_357 (O_357,N_14751,N_14164);
and UO_358 (O_358,N_10052,N_10284);
and UO_359 (O_359,N_10156,N_14965);
and UO_360 (O_360,N_14152,N_11347);
nor UO_361 (O_361,N_11549,N_13291);
nor UO_362 (O_362,N_14763,N_13961);
or UO_363 (O_363,N_11362,N_11063);
or UO_364 (O_364,N_13769,N_13843);
nor UO_365 (O_365,N_11883,N_10958);
or UO_366 (O_366,N_14218,N_10827);
and UO_367 (O_367,N_11887,N_10596);
nand UO_368 (O_368,N_11769,N_10815);
and UO_369 (O_369,N_10543,N_12802);
and UO_370 (O_370,N_14291,N_11051);
nand UO_371 (O_371,N_13738,N_10068);
nand UO_372 (O_372,N_11978,N_13432);
nand UO_373 (O_373,N_12097,N_10176);
or UO_374 (O_374,N_12180,N_12633);
or UO_375 (O_375,N_13644,N_11561);
nand UO_376 (O_376,N_10087,N_14402);
nor UO_377 (O_377,N_14702,N_11816);
or UO_378 (O_378,N_14442,N_14824);
nand UO_379 (O_379,N_13654,N_13565);
nand UO_380 (O_380,N_14625,N_10121);
nor UO_381 (O_381,N_10972,N_10984);
nand UO_382 (O_382,N_14083,N_14061);
and UO_383 (O_383,N_11460,N_13078);
nor UO_384 (O_384,N_13216,N_14723);
nor UO_385 (O_385,N_12899,N_11689);
nor UO_386 (O_386,N_13154,N_14099);
and UO_387 (O_387,N_13409,N_10403);
nor UO_388 (O_388,N_14800,N_13032);
nor UO_389 (O_389,N_10590,N_14236);
and UO_390 (O_390,N_11858,N_12214);
and UO_391 (O_391,N_13887,N_14553);
or UO_392 (O_392,N_14925,N_13516);
or UO_393 (O_393,N_14150,N_13998);
nor UO_394 (O_394,N_11261,N_14068);
nand UO_395 (O_395,N_11272,N_13075);
or UO_396 (O_396,N_11355,N_14547);
nor UO_397 (O_397,N_13120,N_13884);
and UO_398 (O_398,N_14107,N_13498);
nor UO_399 (O_399,N_11083,N_10312);
and UO_400 (O_400,N_11534,N_13438);
or UO_401 (O_401,N_11513,N_13816);
or UO_402 (O_402,N_14220,N_13942);
and UO_403 (O_403,N_11026,N_11550);
or UO_404 (O_404,N_12493,N_12837);
nand UO_405 (O_405,N_14365,N_11229);
or UO_406 (O_406,N_11533,N_11611);
nand UO_407 (O_407,N_10096,N_11670);
and UO_408 (O_408,N_11100,N_12295);
nor UO_409 (O_409,N_14679,N_12019);
nor UO_410 (O_410,N_12580,N_14171);
or UO_411 (O_411,N_10980,N_12313);
or UO_412 (O_412,N_14158,N_12092);
and UO_413 (O_413,N_11617,N_12607);
or UO_414 (O_414,N_14778,N_14511);
nand UO_415 (O_415,N_10771,N_14554);
or UO_416 (O_416,N_13204,N_14339);
nor UO_417 (O_417,N_14518,N_14590);
or UO_418 (O_418,N_13241,N_12376);
nand UO_419 (O_419,N_10698,N_11203);
nand UO_420 (O_420,N_12885,N_14602);
nand UO_421 (O_421,N_11633,N_13115);
nand UO_422 (O_422,N_14256,N_13098);
or UO_423 (O_423,N_12241,N_13422);
and UO_424 (O_424,N_14231,N_12934);
nand UO_425 (O_425,N_12639,N_14232);
and UO_426 (O_426,N_10144,N_12753);
and UO_427 (O_427,N_11310,N_10510);
or UO_428 (O_428,N_11370,N_11886);
nand UO_429 (O_429,N_14096,N_10367);
nand UO_430 (O_430,N_10053,N_14120);
nand UO_431 (O_431,N_14520,N_12100);
and UO_432 (O_432,N_11376,N_10774);
or UO_433 (O_433,N_11213,N_11860);
or UO_434 (O_434,N_10664,N_10790);
nand UO_435 (O_435,N_11981,N_13914);
and UO_436 (O_436,N_14234,N_12959);
and UO_437 (O_437,N_12380,N_14069);
nor UO_438 (O_438,N_12588,N_10759);
nand UO_439 (O_439,N_10540,N_13214);
nand UO_440 (O_440,N_11950,N_13767);
and UO_441 (O_441,N_13454,N_13863);
and UO_442 (O_442,N_13383,N_12006);
nor UO_443 (O_443,N_13847,N_13754);
and UO_444 (O_444,N_12797,N_10876);
nand UO_445 (O_445,N_13131,N_11645);
and UO_446 (O_446,N_13928,N_13341);
and UO_447 (O_447,N_10692,N_13771);
nand UO_448 (O_448,N_14147,N_11671);
and UO_449 (O_449,N_13287,N_13626);
nor UO_450 (O_450,N_11528,N_11608);
and UO_451 (O_451,N_10161,N_12982);
nand UO_452 (O_452,N_12597,N_13411);
nor UO_453 (O_453,N_14010,N_11182);
nand UO_454 (O_454,N_12382,N_14125);
and UO_455 (O_455,N_14510,N_10734);
nand UO_456 (O_456,N_10796,N_10290);
and UO_457 (O_457,N_11818,N_11348);
and UO_458 (O_458,N_12002,N_10357);
or UO_459 (O_459,N_11951,N_12666);
and UO_460 (O_460,N_10787,N_12099);
or UO_461 (O_461,N_11600,N_13641);
nand UO_462 (O_462,N_14475,N_14821);
nor UO_463 (O_463,N_12728,N_14112);
nand UO_464 (O_464,N_14585,N_12108);
nor UO_465 (O_465,N_10806,N_10591);
nor UO_466 (O_466,N_12370,N_11205);
and UO_467 (O_467,N_12427,N_10253);
and UO_468 (O_468,N_14298,N_12258);
nand UO_469 (O_469,N_12590,N_13177);
or UO_470 (O_470,N_10202,N_10805);
nor UO_471 (O_471,N_12953,N_14237);
and UO_472 (O_472,N_12208,N_11546);
and UO_473 (O_473,N_12702,N_14151);
nand UO_474 (O_474,N_12484,N_10047);
nand UO_475 (O_475,N_14738,N_12430);
nor UO_476 (O_476,N_11074,N_14904);
or UO_477 (O_477,N_10494,N_12331);
or UO_478 (O_478,N_14159,N_10872);
nor UO_479 (O_479,N_10951,N_11172);
or UO_480 (O_480,N_14205,N_12688);
and UO_481 (O_481,N_12361,N_12357);
and UO_482 (O_482,N_12268,N_14805);
nand UO_483 (O_483,N_10371,N_13353);
nand UO_484 (O_484,N_13707,N_14952);
nand UO_485 (O_485,N_12715,N_12137);
and UO_486 (O_486,N_12244,N_12592);
and UO_487 (O_487,N_13113,N_14570);
nand UO_488 (O_488,N_12094,N_10653);
nor UO_489 (O_489,N_12809,N_12988);
and UO_490 (O_490,N_11646,N_11606);
nand UO_491 (O_491,N_12400,N_11427);
nor UO_492 (O_492,N_11387,N_10362);
and UO_493 (O_493,N_12710,N_10814);
nand UO_494 (O_494,N_12069,N_13414);
and UO_495 (O_495,N_11634,N_12814);
nor UO_496 (O_496,N_12012,N_13174);
nand UO_497 (O_497,N_13774,N_13621);
nor UO_498 (O_498,N_10667,N_12272);
nor UO_499 (O_499,N_11411,N_11359);
nand UO_500 (O_500,N_10172,N_11448);
nor UO_501 (O_501,N_10245,N_13797);
nor UO_502 (O_502,N_13129,N_12619);
or UO_503 (O_503,N_10646,N_13031);
and UO_504 (O_504,N_11834,N_14771);
or UO_505 (O_505,N_12733,N_10224);
nor UO_506 (O_506,N_11342,N_10841);
or UO_507 (O_507,N_12112,N_13433);
and UO_508 (O_508,N_13594,N_12348);
nand UO_509 (O_509,N_10738,N_12196);
and UO_510 (O_510,N_13141,N_12176);
and UO_511 (O_511,N_14928,N_14998);
nor UO_512 (O_512,N_13269,N_10115);
and UO_513 (O_513,N_13125,N_12973);
or UO_514 (O_514,N_13781,N_10983);
nor UO_515 (O_515,N_10194,N_12090);
nand UO_516 (O_516,N_11245,N_10127);
nor UO_517 (O_517,N_10557,N_11199);
nor UO_518 (O_518,N_11093,N_11267);
or UO_519 (O_519,N_10619,N_11451);
nor UO_520 (O_520,N_12038,N_12746);
or UO_521 (O_521,N_12566,N_10060);
nand UO_522 (O_522,N_10758,N_10086);
or UO_523 (O_523,N_12532,N_11331);
nor UO_524 (O_524,N_13323,N_13564);
nand UO_525 (O_525,N_14961,N_14007);
or UO_526 (O_526,N_14870,N_10642);
or UO_527 (O_527,N_14533,N_11788);
nor UO_528 (O_528,N_10100,N_11696);
nand UO_529 (O_529,N_14977,N_10781);
and UO_530 (O_530,N_13451,N_11655);
or UO_531 (O_531,N_10754,N_10213);
and UO_532 (O_532,N_14793,N_14355);
or UO_533 (O_533,N_12777,N_11949);
nor UO_534 (O_534,N_12578,N_13789);
nand UO_535 (O_535,N_13585,N_12153);
nand UO_536 (O_536,N_13649,N_10309);
or UO_537 (O_537,N_11308,N_14391);
nand UO_538 (O_538,N_14425,N_12332);
nor UO_539 (O_539,N_12692,N_10046);
and UO_540 (O_540,N_12290,N_10056);
and UO_541 (O_541,N_12527,N_10095);
nor UO_542 (O_542,N_10514,N_13202);
or UO_543 (O_543,N_11227,N_14710);
xnor UO_544 (O_544,N_11102,N_12045);
and UO_545 (O_545,N_14411,N_12762);
or UO_546 (O_546,N_11668,N_14255);
nor UO_547 (O_547,N_11185,N_11292);
or UO_548 (O_548,N_13096,N_14656);
and UO_549 (O_549,N_14788,N_13201);
and UO_550 (O_550,N_11766,N_10193);
or UO_551 (O_551,N_13095,N_14190);
and UO_552 (O_552,N_12163,N_12062);
nand UO_553 (O_553,N_12315,N_13534);
nor UO_554 (O_554,N_11588,N_13879);
and UO_555 (O_555,N_10440,N_14874);
nand UO_556 (O_556,N_13416,N_10102);
nand UO_557 (O_557,N_10750,N_11762);
nand UO_558 (O_558,N_14953,N_13161);
or UO_559 (O_559,N_14088,N_12020);
or UO_560 (O_560,N_10632,N_10148);
nor UO_561 (O_561,N_13021,N_10763);
and UO_562 (O_562,N_12966,N_10474);
and UO_563 (O_563,N_11345,N_11807);
and UO_564 (O_564,N_12551,N_11059);
or UO_565 (O_565,N_13343,N_12183);
nor UO_566 (O_566,N_12693,N_13273);
nor UO_567 (O_567,N_13664,N_13651);
and UO_568 (O_568,N_10842,N_12996);
nand UO_569 (O_569,N_14749,N_14368);
nand UO_570 (O_570,N_12998,N_10030);
and UO_571 (O_571,N_12472,N_12983);
and UO_572 (O_572,N_11810,N_10113);
or UO_573 (O_573,N_12676,N_10875);
or UO_574 (O_574,N_14745,N_11209);
or UO_575 (O_575,N_10624,N_13185);
nand UO_576 (O_576,N_11468,N_14890);
or UO_577 (O_577,N_11120,N_10573);
nand UO_578 (O_578,N_11221,N_11772);
nand UO_579 (O_579,N_10333,N_13044);
nor UO_580 (O_580,N_13380,N_10940);
and UO_581 (O_581,N_14500,N_10885);
and UO_582 (O_582,N_10463,N_10233);
nand UO_583 (O_583,N_14243,N_13640);
and UO_584 (O_584,N_11757,N_11914);
xnor UO_585 (O_585,N_11425,N_13022);
nor UO_586 (O_586,N_14307,N_10823);
and UO_587 (O_587,N_11593,N_12862);
nand UO_588 (O_588,N_11901,N_10800);
nor UO_589 (O_589,N_14930,N_13365);
and UO_590 (O_590,N_10733,N_11259);
or UO_591 (O_591,N_12047,N_12792);
and UO_592 (O_592,N_14662,N_10712);
and UO_593 (O_593,N_10346,N_12811);
nand UO_594 (O_594,N_10420,N_11735);
nor UO_595 (O_595,N_12362,N_14497);
or UO_596 (O_596,N_14153,N_10379);
or UO_597 (O_597,N_10375,N_14354);
and UO_598 (O_598,N_10430,N_12903);
nand UO_599 (O_599,N_13245,N_12307);
and UO_600 (O_600,N_13647,N_10308);
and UO_601 (O_601,N_12817,N_14384);
nand UO_602 (O_602,N_11845,N_14825);
nor UO_603 (O_603,N_11944,N_12425);
or UO_604 (O_604,N_14779,N_11191);
or UO_605 (O_605,N_14543,N_12197);
and UO_606 (O_606,N_13992,N_12858);
and UO_607 (O_607,N_12037,N_13878);
and UO_608 (O_608,N_10908,N_12544);
and UO_609 (O_609,N_11725,N_13704);
nand UO_610 (O_610,N_14155,N_14626);
nand UO_611 (O_611,N_13721,N_10154);
and UO_612 (O_612,N_11543,N_14996);
and UO_613 (O_613,N_14011,N_10131);
and UO_614 (O_614,N_14058,N_13232);
xor UO_615 (O_615,N_10457,N_10132);
or UO_616 (O_616,N_12638,N_14703);
or UO_617 (O_617,N_11306,N_10130);
or UO_618 (O_618,N_12171,N_11247);
and UO_619 (O_619,N_10225,N_10924);
and UO_620 (O_620,N_13814,N_13436);
nand UO_621 (O_621,N_13061,N_11651);
and UO_622 (O_622,N_12725,N_10314);
or UO_623 (O_623,N_11149,N_11097);
nand UO_624 (O_624,N_14102,N_11044);
nor UO_625 (O_625,N_10183,N_11393);
nor UO_626 (O_626,N_11595,N_12871);
nand UO_627 (O_627,N_10569,N_10168);
nand UO_628 (O_628,N_10501,N_10276);
nand UO_629 (O_629,N_11749,N_12177);
nand UO_630 (O_630,N_10877,N_14829);
nand UO_631 (O_631,N_14048,N_12750);
nand UO_632 (O_632,N_10941,N_13953);
or UO_633 (O_633,N_11804,N_14964);
nor UO_634 (O_634,N_11605,N_11364);
or UO_635 (O_635,N_12204,N_14235);
nor UO_636 (O_636,N_11535,N_10963);
or UO_637 (O_637,N_14487,N_14866);
or UO_638 (O_638,N_11787,N_12221);
and UO_639 (O_639,N_14461,N_14857);
and UO_640 (O_640,N_12727,N_13981);
nor UO_641 (O_641,N_11358,N_13473);
or UO_642 (O_642,N_10899,N_12293);
nor UO_643 (O_643,N_12301,N_12147);
and UO_644 (O_644,N_10069,N_10920);
or UO_645 (O_645,N_10186,N_10320);
or UO_646 (O_646,N_13260,N_10190);
or UO_647 (O_647,N_11910,N_13278);
or UO_648 (O_648,N_14892,N_12717);
and UO_649 (O_649,N_14528,N_10745);
nor UO_650 (O_650,N_12220,N_14066);
and UO_651 (O_651,N_12059,N_13906);
nand UO_652 (O_652,N_14195,N_12821);
and UO_653 (O_653,N_10803,N_13165);
nor UO_654 (O_654,N_13537,N_13127);
nor UO_655 (O_655,N_11244,N_11953);
nor UO_656 (O_656,N_10895,N_10864);
nor UO_657 (O_657,N_14945,N_10843);
nor UO_658 (O_658,N_13488,N_14651);
nor UO_659 (O_659,N_12771,N_12640);
nand UO_660 (O_660,N_12247,N_13871);
or UO_661 (O_661,N_10696,N_13076);
nand UO_662 (O_662,N_14075,N_11752);
and UO_663 (O_663,N_10866,N_12237);
or UO_664 (O_664,N_10702,N_14300);
nand UO_665 (O_665,N_10182,N_14540);
and UO_666 (O_666,N_13970,N_11441);
and UO_667 (O_667,N_13835,N_10104);
and UO_668 (O_668,N_10203,N_10399);
nor UO_669 (O_669,N_13497,N_10336);
nand UO_670 (O_670,N_12606,N_11729);
nor UO_671 (O_671,N_12584,N_14428);
or UO_672 (O_672,N_12044,N_12864);
or UO_673 (O_673,N_14351,N_12835);
and UO_674 (O_674,N_11985,N_10769);
nor UO_675 (O_675,N_11311,N_13143);
and UO_676 (O_676,N_14534,N_10997);
nor UO_677 (O_677,N_11620,N_14942);
nand UO_678 (O_678,N_13850,N_13085);
nand UO_679 (O_679,N_14359,N_13456);
and UO_680 (O_680,N_12714,N_13217);
nor UO_681 (O_681,N_10607,N_13469);
and UO_682 (O_682,N_13496,N_14732);
and UO_683 (O_683,N_11984,N_11187);
and UO_684 (O_684,N_14556,N_11313);
and UO_685 (O_685,N_12233,N_11870);
or UO_686 (O_686,N_12286,N_13317);
nor UO_687 (O_687,N_14583,N_11132);
and UO_688 (O_688,N_10443,N_11105);
nor UO_689 (O_689,N_10942,N_11974);
and UO_690 (O_690,N_14869,N_14675);
or UO_691 (O_691,N_14340,N_14439);
or UO_692 (O_692,N_11129,N_12696);
and UO_693 (O_693,N_13458,N_13688);
nand UO_694 (O_694,N_12083,N_10661);
or UO_695 (O_695,N_12457,N_14198);
nand UO_696 (O_696,N_12711,N_12796);
xor UO_697 (O_697,N_10341,N_13968);
and UO_698 (O_698,N_14347,N_13003);
nand UO_699 (O_699,N_11297,N_10076);
or UO_700 (O_700,N_14086,N_13051);
and UO_701 (O_701,N_13719,N_13679);
and UO_702 (O_702,N_12667,N_10306);
and UO_703 (O_703,N_10282,N_10789);
or UO_704 (O_704,N_14539,N_12463);
or UO_705 (O_705,N_11640,N_12065);
xnor UO_706 (O_706,N_11257,N_13100);
nand UO_707 (O_707,N_13225,N_10614);
nor UO_708 (O_708,N_13123,N_10088);
or UO_709 (O_709,N_13582,N_10810);
or UO_710 (O_710,N_11438,N_14514);
and UO_711 (O_711,N_10880,N_14207);
nand UO_712 (O_712,N_14863,N_12210);
nor UO_713 (O_713,N_11879,N_13619);
or UO_714 (O_714,N_12422,N_12119);
or UO_715 (O_715,N_14742,N_14783);
or UO_716 (O_716,N_13013,N_10945);
or UO_717 (O_717,N_11733,N_14170);
nor UO_718 (O_718,N_12536,N_11713);
xnor UO_719 (O_719,N_13248,N_12873);
nand UO_720 (O_720,N_12428,N_14568);
or UO_721 (O_721,N_11353,N_12262);
nand UO_722 (O_722,N_12933,N_10486);
nand UO_723 (O_723,N_11397,N_11730);
and UO_724 (O_724,N_13517,N_11036);
nand UO_725 (O_725,N_13931,N_10361);
nand UO_726 (O_726,N_13118,N_14713);
or UO_727 (O_727,N_12503,N_13374);
and UO_728 (O_728,N_13135,N_11632);
and UO_729 (O_729,N_12368,N_10133);
and UO_730 (O_730,N_13925,N_12863);
nand UO_731 (O_731,N_12736,N_13806);
nand UO_732 (O_732,N_12249,N_13427);
or UO_733 (O_733,N_11004,N_11081);
or UO_734 (O_734,N_12708,N_12016);
and UO_735 (O_735,N_12155,N_11966);
and UO_736 (O_736,N_11151,N_13308);
nor UO_737 (O_737,N_14833,N_14560);
and UO_738 (O_738,N_11068,N_14228);
nand UO_739 (O_739,N_12470,N_11381);
nand UO_740 (O_740,N_12504,N_10731);
and UO_741 (O_741,N_14858,N_11890);
or UO_742 (O_742,N_12270,N_13344);
nor UO_743 (O_743,N_12927,N_14377);
or UO_744 (O_744,N_11638,N_14692);
or UO_745 (O_745,N_14272,N_11774);
nand UO_746 (O_746,N_13237,N_12610);
xor UO_747 (O_747,N_14142,N_10490);
or UO_748 (O_748,N_14652,N_10574);
nor UO_749 (O_749,N_13512,N_14849);
or UO_750 (O_750,N_11933,N_13812);
nor UO_751 (O_751,N_14465,N_10735);
and UO_752 (O_752,N_11792,N_10727);
and UO_753 (O_753,N_12223,N_10977);
or UO_754 (O_754,N_11578,N_10560);
and UO_755 (O_755,N_10536,N_11281);
and UO_756 (O_756,N_14938,N_13164);
or UO_757 (O_757,N_14704,N_13430);
and UO_758 (O_758,N_13837,N_11295);
nand UO_759 (O_759,N_14962,N_13725);
nor UO_760 (O_760,N_10881,N_11706);
and UO_761 (O_761,N_13672,N_12747);
and UO_762 (O_762,N_10545,N_10492);
nor UO_763 (O_763,N_11629,N_12187);
nor UO_764 (O_764,N_11783,N_13077);
or UO_765 (O_765,N_11231,N_11905);
or UO_766 (O_766,N_13807,N_14864);
xor UO_767 (O_767,N_13408,N_11570);
nor UO_768 (O_768,N_14837,N_12507);
or UO_769 (O_769,N_10207,N_10106);
and UO_770 (O_770,N_10462,N_10999);
nand UO_771 (O_771,N_10411,N_13840);
nand UO_772 (O_772,N_13728,N_12672);
nor UO_773 (O_773,N_14293,N_12490);
nor UO_774 (O_774,N_10214,N_13311);
nor UO_775 (O_775,N_14309,N_13965);
or UO_776 (O_776,N_13471,N_13620);
or UO_777 (O_777,N_12992,N_13336);
and UO_778 (O_778,N_12758,N_14270);
and UO_779 (O_779,N_10602,N_12126);
nand UO_780 (O_780,N_12347,N_14301);
nor UO_781 (O_781,N_13759,N_13364);
and UO_782 (O_782,N_12316,N_10794);
nor UO_783 (O_783,N_10605,N_11664);
or UO_784 (O_784,N_12553,N_12184);
nand UO_785 (O_785,N_12649,N_14498);
and UO_786 (O_786,N_13819,N_12944);
or UO_787 (O_787,N_12421,N_14935);
nor UO_788 (O_788,N_12379,N_14804);
nor UO_789 (O_789,N_12289,N_13097);
and UO_790 (O_790,N_10386,N_14379);
and UO_791 (O_791,N_13882,N_12636);
nor UO_792 (O_792,N_12841,N_13782);
nor UO_793 (O_793,N_10022,N_13558);
and UO_794 (O_794,N_10838,N_13182);
nor UO_795 (O_795,N_11011,N_13650);
nand UO_796 (O_796,N_12070,N_11539);
or UO_797 (O_797,N_14322,N_10959);
and UO_798 (O_798,N_10175,N_10423);
nor UO_799 (O_799,N_12402,N_10897);
and UO_800 (O_800,N_13890,N_11431);
and UO_801 (O_801,N_13043,N_11365);
or UO_802 (O_802,N_11417,N_13883);
or UO_803 (O_803,N_11656,N_11672);
or UO_804 (O_804,N_10028,N_12518);
xor UO_805 (O_805,N_11505,N_14898);
or UO_806 (O_806,N_13618,N_11494);
nand UO_807 (O_807,N_13238,N_13757);
or UO_808 (O_808,N_11893,N_10339);
and UO_809 (O_809,N_11959,N_10844);
or UO_810 (O_810,N_10884,N_12916);
nor UO_811 (O_811,N_13778,N_12972);
nand UO_812 (O_812,N_11891,N_10645);
or UO_813 (O_813,N_12113,N_11125);
and UO_814 (O_814,N_12148,N_11192);
nor UO_815 (O_815,N_11771,N_11971);
or UO_816 (O_816,N_12042,N_11225);
or UO_817 (O_817,N_12459,N_13748);
xnor UO_818 (O_818,N_14466,N_11897);
nor UO_819 (O_819,N_13503,N_14101);
and UO_820 (O_820,N_10329,N_13793);
nor UO_821 (O_821,N_14695,N_14618);
or UO_822 (O_822,N_10321,N_10849);
and UO_823 (O_823,N_12828,N_12524);
and UO_824 (O_824,N_14040,N_13060);
nor UO_825 (O_825,N_11924,N_12742);
or UO_826 (O_826,N_11133,N_11625);
and UO_827 (O_827,N_11200,N_11707);
nand UO_828 (O_828,N_10001,N_10685);
nor UO_829 (O_829,N_10882,N_10651);
nand UO_830 (O_830,N_11803,N_11798);
or UO_831 (O_831,N_12334,N_11006);
nor UO_832 (O_832,N_13561,N_11062);
or UO_833 (O_833,N_11223,N_12125);
nor UO_834 (O_834,N_10352,N_12808);
nand UO_835 (O_835,N_11194,N_14077);
nand UO_836 (O_836,N_14707,N_10023);
and UO_837 (O_837,N_11114,N_11196);
nor UO_838 (O_838,N_10111,N_10672);
nor UO_839 (O_839,N_11252,N_10812);
or UO_840 (O_840,N_11802,N_13749);
or UO_841 (O_841,N_14850,N_13876);
and UO_842 (O_842,N_14693,N_11122);
or UO_843 (O_843,N_10472,N_11987);
nand UO_844 (O_844,N_10684,N_10377);
and UO_845 (O_845,N_14798,N_14397);
nand UO_846 (O_846,N_12468,N_13838);
and UO_847 (O_847,N_13345,N_11698);
or UO_848 (O_848,N_13071,N_14206);
or UO_849 (O_849,N_10623,N_13652);
or UO_850 (O_850,N_14350,N_14812);
xnor UO_851 (O_851,N_10571,N_12494);
nand UO_852 (O_852,N_11763,N_13319);
or UO_853 (O_853,N_14729,N_14822);
or UO_854 (O_854,N_14390,N_11589);
or UO_855 (O_855,N_12464,N_13254);
or UO_856 (O_856,N_12106,N_14200);
or UO_857 (O_857,N_12582,N_10979);
or UO_858 (O_858,N_11116,N_12570);
nor UO_859 (O_859,N_14663,N_14480);
and UO_860 (O_860,N_12967,N_12105);
or UO_861 (O_861,N_12231,N_14883);
nor UO_862 (O_862,N_11667,N_10993);
nor UO_863 (O_863,N_13064,N_12654);
nor UO_864 (O_864,N_11099,N_12876);
nor UO_865 (O_865,N_10040,N_12653);
nand UO_866 (O_866,N_13859,N_10861);
nand UO_867 (O_867,N_14045,N_13055);
or UO_868 (O_868,N_10431,N_12807);
nor UO_869 (O_869,N_12950,N_12154);
or UO_870 (O_870,N_10818,N_14254);
nand UO_871 (O_871,N_12805,N_14395);
nor UO_872 (O_872,N_14753,N_13801);
nor UO_873 (O_873,N_11685,N_13091);
and UO_874 (O_874,N_12529,N_13358);
or UO_875 (O_875,N_13962,N_10907);
nand UO_876 (O_876,N_13509,N_14766);
nand UO_877 (O_877,N_13519,N_12050);
nand UO_878 (O_878,N_12475,N_10928);
or UO_879 (O_879,N_12120,N_12832);
and UO_880 (O_880,N_10846,N_14091);
and UO_881 (O_881,N_11962,N_14446);
nand UO_882 (O_882,N_10244,N_13486);
nand UO_883 (O_883,N_11532,N_14464);
and UO_884 (O_884,N_10406,N_10757);
nand UO_885 (O_885,N_12001,N_12549);
nand UO_886 (O_886,N_13067,N_14286);
or UO_887 (O_887,N_14044,N_12401);
xor UO_888 (O_888,N_13880,N_12133);
nor UO_889 (O_889,N_11177,N_13136);
nor UO_890 (O_890,N_12043,N_12843);
or UO_891 (O_891,N_11753,N_11165);
or UO_892 (O_892,N_10926,N_10826);
or UO_893 (O_893,N_10726,N_11734);
nand UO_894 (O_894,N_10044,N_13418);
and UO_895 (O_895,N_13934,N_12838);
nor UO_896 (O_896,N_14289,N_12913);
or UO_897 (O_897,N_14186,N_12514);
nor UO_898 (O_898,N_12363,N_14327);
and UO_899 (O_899,N_14997,N_11571);
and UO_900 (O_900,N_14208,N_14912);
and UO_901 (O_901,N_14669,N_10299);
and UO_902 (O_902,N_12786,N_14468);
nor UO_903 (O_903,N_11830,N_10280);
and UO_904 (O_904,N_11080,N_14993);
and UO_905 (O_905,N_12923,N_10502);
nor UO_906 (O_906,N_14604,N_13152);
or UO_907 (O_907,N_14383,N_11264);
or UO_908 (O_908,N_11091,N_11139);
or UO_909 (O_909,N_10476,N_11599);
nor UO_910 (O_910,N_14686,N_11070);
nor UO_911 (O_911,N_10515,N_11642);
nand UO_912 (O_912,N_11224,N_14343);
and UO_913 (O_913,N_10461,N_14462);
nand UO_914 (O_914,N_10974,N_14999);
nand UO_915 (O_915,N_14388,N_14887);
nor UO_916 (O_916,N_10649,N_14574);
and UO_917 (O_917,N_13825,N_12124);
and UO_918 (O_918,N_11317,N_14595);
and UO_919 (O_919,N_11510,N_14565);
or UO_920 (O_920,N_10797,N_14958);
or UO_921 (O_921,N_10799,N_10220);
nand UO_922 (O_922,N_12203,N_14603);
nand UO_923 (O_923,N_11092,N_11301);
and UO_924 (O_924,N_12227,N_10630);
nand UO_925 (O_925,N_11654,N_11029);
and UO_926 (O_926,N_14470,N_11956);
or UO_927 (O_927,N_10482,N_12931);
nor UO_928 (O_928,N_13923,N_14791);
nand UO_929 (O_929,N_12585,N_10143);
or UO_930 (O_930,N_14079,N_11869);
nand UO_931 (O_931,N_12684,N_10824);
or UO_932 (O_932,N_12051,N_11619);
nand UO_933 (O_933,N_13978,N_13901);
or UO_934 (O_934,N_11936,N_13877);
or UO_935 (O_935,N_12088,N_12756);
nor UO_936 (O_936,N_13266,N_11744);
nand UO_937 (O_937,N_13870,N_13987);
nor UO_938 (O_938,N_10539,N_14028);
or UO_939 (O_939,N_11745,N_10222);
nand UO_940 (O_940,N_13677,N_13126);
and UO_941 (O_941,N_14676,N_14376);
nor UO_942 (O_942,N_12281,N_10834);
or UO_943 (O_943,N_10378,N_13233);
nor UO_944 (O_944,N_10851,N_13964);
nand UO_945 (O_945,N_14799,N_11682);
and UO_946 (O_946,N_14584,N_10077);
or UO_947 (O_947,N_11723,N_12823);
or UO_948 (O_948,N_14034,N_12946);
nor UO_949 (O_949,N_10592,N_11178);
nor UO_950 (O_950,N_10710,N_12248);
and UO_951 (O_951,N_10018,N_14673);
nand UO_952 (O_952,N_11319,N_12526);
and UO_953 (O_953,N_13017,N_14132);
and UO_954 (O_954,N_12027,N_10091);
or UO_955 (O_955,N_11202,N_11478);
nor UO_956 (O_956,N_10793,N_11330);
and UO_957 (O_957,N_11709,N_12738);
nand UO_958 (O_958,N_11027,N_14970);
nand UO_959 (O_959,N_10565,N_12443);
nor UO_960 (O_960,N_10210,N_14129);
nand UO_961 (O_961,N_12003,N_14288);
or UO_962 (O_962,N_14245,N_11562);
and UO_963 (O_963,N_13203,N_12222);
or UO_964 (O_964,N_11544,N_10415);
and UO_965 (O_965,N_10628,N_13681);
nand UO_966 (O_966,N_14115,N_11906);
nor UO_967 (O_967,N_14144,N_14434);
nand UO_968 (O_968,N_12668,N_14260);
and UO_969 (O_969,N_12877,N_14246);
nor UO_970 (O_970,N_13623,N_10303);
nand UO_971 (O_971,N_12415,N_13888);
and UO_972 (O_972,N_14213,N_12655);
nor UO_973 (O_973,N_14441,N_13133);
nor UO_974 (O_974,N_11085,N_11658);
or UO_975 (O_975,N_14089,N_12624);
and UO_976 (O_976,N_13352,N_14319);
nand UO_977 (O_977,N_14986,N_10654);
and UO_978 (O_978,N_14768,N_10855);
or UO_979 (O_979,N_13446,N_14067);
nor UO_980 (O_980,N_14160,N_12989);
or UO_981 (O_981,N_11171,N_14042);
nor UO_982 (O_982,N_14267,N_10149);
nor UO_983 (O_983,N_11838,N_11509);
nand UO_984 (O_984,N_13101,N_12849);
and UO_985 (O_985,N_12769,N_11568);
nand UO_986 (O_986,N_10933,N_10935);
nand UO_987 (O_987,N_13130,N_14128);
nand UO_988 (O_988,N_14950,N_13536);
or UO_989 (O_989,N_10109,N_12656);
and UO_990 (O_990,N_10549,N_12476);
or UO_991 (O_991,N_10857,N_11360);
or UO_992 (O_992,N_10448,N_14853);
nor UO_993 (O_993,N_12257,N_11674);
or UO_994 (O_994,N_13706,N_14776);
nand UO_995 (O_995,N_12775,N_11372);
or UO_996 (O_996,N_12793,N_12269);
and UO_997 (O_997,N_14296,N_12506);
nand UO_998 (O_998,N_10955,N_11422);
and UO_999 (O_999,N_10187,N_10470);
and UO_1000 (O_1000,N_12167,N_10295);
nor UO_1001 (O_1001,N_12683,N_10101);
nor UO_1002 (O_1002,N_12621,N_11401);
and UO_1003 (O_1003,N_10768,N_11523);
nor UO_1004 (O_1004,N_14770,N_11346);
and UO_1005 (O_1005,N_12941,N_10153);
and UO_1006 (O_1006,N_11842,N_14995);
nor UO_1007 (O_1007,N_13813,N_10715);
nand UO_1008 (O_1008,N_10660,N_11095);
nand UO_1009 (O_1009,N_10711,N_11307);
or UO_1010 (O_1010,N_14303,N_12238);
nor UO_1011 (O_1011,N_14645,N_14914);
and UO_1012 (O_1012,N_14357,N_11607);
or UO_1013 (O_1013,N_10585,N_14561);
nand UO_1014 (O_1014,N_12999,N_11294);
nand UO_1015 (O_1015,N_10242,N_10756);
and UO_1016 (O_1016,N_10716,N_14165);
nor UO_1017 (O_1017,N_13636,N_13969);
and UO_1018 (O_1018,N_13856,N_13304);
and UO_1019 (O_1019,N_11399,N_13936);
nor UO_1020 (O_1020,N_13524,N_14754);
and UO_1021 (O_1021,N_10118,N_10123);
or UO_1022 (O_1022,N_11884,N_14891);
and UO_1023 (O_1023,N_14963,N_12798);
and UO_1024 (O_1024,N_11943,N_12466);
nand UO_1025 (O_1025,N_10617,N_12617);
nor UO_1026 (O_1026,N_13866,N_14062);
nand UO_1027 (O_1027,N_11741,N_10985);
and UO_1028 (O_1028,N_12540,N_13466);
nand UO_1029 (O_1029,N_11989,N_12976);
and UO_1030 (O_1030,N_11557,N_14315);
and UO_1031 (O_1031,N_13584,N_11180);
nor UO_1032 (O_1032,N_13573,N_11148);
and UO_1033 (O_1033,N_13560,N_13482);
nand UO_1034 (O_1034,N_13529,N_14991);
and UO_1035 (O_1035,N_14535,N_14960);
and UO_1036 (O_1036,N_11072,N_13690);
nand UO_1037 (O_1037,N_12569,N_13656);
nor UO_1038 (O_1038,N_13794,N_13784);
and UO_1039 (O_1039,N_14342,N_12605);
or UO_1040 (O_1040,N_10873,N_10445);
and UO_1041 (O_1041,N_10725,N_12690);
nand UO_1042 (O_1042,N_12409,N_14191);
and UO_1043 (O_1043,N_11190,N_10421);
nor UO_1044 (O_1044,N_14687,N_14032);
or UO_1045 (O_1045,N_14989,N_12366);
nor UO_1046 (O_1046,N_13357,N_12670);
nand UO_1047 (O_1047,N_11497,N_12116);
and UO_1048 (O_1048,N_11705,N_11840);
and UO_1049 (O_1049,N_13590,N_11911);
or UO_1050 (O_1050,N_14493,N_12525);
xnor UO_1051 (O_1051,N_12760,N_12117);
nand UO_1052 (O_1052,N_14557,N_14517);
and UO_1053 (O_1053,N_12201,N_11912);
nand UO_1054 (O_1054,N_14835,N_12924);
and UO_1055 (O_1055,N_14277,N_13339);
and UO_1056 (O_1056,N_12478,N_10254);
or UO_1057 (O_1057,N_14356,N_12765);
nor UO_1058 (O_1058,N_14216,N_11881);
or UO_1059 (O_1059,N_14209,N_13068);
nand UO_1060 (O_1060,N_10775,N_13765);
nor UO_1061 (O_1061,N_10613,N_14813);
and UO_1062 (O_1062,N_12833,N_10533);
nor UO_1063 (O_1063,N_11821,N_11485);
and UO_1064 (O_1064,N_10839,N_10894);
and UO_1065 (O_1065,N_12681,N_14752);
or UO_1066 (O_1066,N_13924,N_12166);
nor UO_1067 (O_1067,N_13244,N_11168);
nand UO_1068 (O_1068,N_12642,N_12895);
and UO_1069 (O_1069,N_10117,N_14609);
nand UO_1070 (O_1070,N_13063,N_13788);
and UO_1071 (O_1071,N_13014,N_13697);
nor UO_1072 (O_1072,N_14413,N_13167);
and UO_1073 (O_1073,N_13518,N_10678);
and UO_1074 (O_1074,N_10318,N_10468);
nand UO_1075 (O_1075,N_13159,N_11695);
nor UO_1076 (O_1076,N_12369,N_11554);
or UO_1077 (O_1077,N_11157,N_11808);
nor UO_1078 (O_1078,N_13168,N_14660);
or UO_1079 (O_1079,N_14452,N_10304);
nand UO_1080 (O_1080,N_13511,N_12677);
and UO_1081 (O_1081,N_12907,N_13271);
nor UO_1082 (O_1082,N_12066,N_13010);
and UO_1083 (O_1083,N_11394,N_11408);
or UO_1084 (O_1084,N_11900,N_10012);
and UO_1085 (O_1085,N_11248,N_13745);
nand UO_1086 (O_1086,N_13988,N_10277);
nand UO_1087 (O_1087,N_12414,N_13139);
and UO_1088 (O_1088,N_12320,N_11161);
and UO_1089 (O_1089,N_12985,N_10900);
nand UO_1090 (O_1090,N_12191,N_10432);
nor UO_1091 (O_1091,N_14992,N_12448);
nor UO_1092 (O_1092,N_13858,N_13508);
and UO_1093 (O_1093,N_10405,N_10266);
nand UO_1094 (O_1094,N_10647,N_13557);
or UO_1095 (O_1095,N_14073,N_11023);
nor UO_1096 (O_1096,N_11717,N_14041);
and UO_1097 (O_1097,N_13426,N_11007);
nand UO_1098 (O_1098,N_13770,N_10652);
nand UO_1099 (O_1099,N_11892,N_13502);
or UO_1100 (O_1100,N_12887,N_10753);
nand UO_1101 (O_1101,N_10229,N_10746);
or UO_1102 (O_1102,N_14927,N_11631);
nor UO_1103 (O_1103,N_12311,N_11560);
nor UO_1104 (O_1104,N_11817,N_13250);
or UO_1105 (O_1105,N_12015,N_14691);
nor UO_1106 (O_1106,N_12872,N_10527);
and UO_1107 (O_1107,N_12719,N_14370);
xnor UO_1108 (O_1108,N_14302,N_13268);
nand UO_1109 (O_1109,N_14861,N_11731);
or UO_1110 (O_1110,N_13634,N_10128);
and UO_1111 (O_1111,N_11343,N_10910);
or UO_1112 (O_1112,N_13399,N_10465);
and UO_1113 (O_1113,N_14087,N_13556);
nor UO_1114 (O_1114,N_10564,N_13321);
and UO_1115 (O_1115,N_11782,N_10007);
nand UO_1116 (O_1116,N_10110,N_13958);
and UO_1117 (O_1117,N_10615,N_11283);
nor UO_1118 (O_1118,N_10434,N_10934);
or UO_1119 (O_1119,N_10124,N_11459);
nor UO_1120 (O_1120,N_14509,N_11531);
and UO_1121 (O_1121,N_12101,N_11222);
and UO_1122 (O_1122,N_13398,N_11065);
or UO_1123 (O_1123,N_14392,N_10508);
or UO_1124 (O_1124,N_12471,N_13006);
or UO_1125 (O_1125,N_11039,N_11413);
and UO_1126 (O_1126,N_12132,N_14868);
and UO_1127 (O_1127,N_14330,N_14735);
and UO_1128 (O_1128,N_14043,N_10201);
or UO_1129 (O_1129,N_14104,N_10011);
and UO_1130 (O_1130,N_13531,N_10523);
or UO_1131 (O_1131,N_11300,N_11878);
nor UO_1132 (O_1132,N_13258,N_10720);
nor UO_1133 (O_1133,N_11849,N_11806);
or UO_1134 (O_1134,N_14103,N_11268);
or UO_1135 (O_1135,N_11999,N_11575);
nand UO_1136 (O_1136,N_11082,N_12029);
nand UO_1137 (O_1137,N_10466,N_12854);
and UO_1138 (O_1138,N_10418,N_10791);
or UO_1139 (O_1139,N_12277,N_12077);
nand UO_1140 (O_1140,N_14332,N_13104);
or UO_1141 (O_1141,N_14612,N_10103);
or UO_1142 (O_1142,N_10552,N_10691);
and UO_1143 (O_1143,N_10126,N_13464);
nand UO_1144 (O_1144,N_14055,N_13029);
nor UO_1145 (O_1145,N_14832,N_11324);
nor UO_1146 (O_1146,N_10116,N_12712);
nand UO_1147 (O_1147,N_13764,N_11604);
or UO_1148 (O_1148,N_14108,N_12501);
and UO_1149 (O_1149,N_13114,N_14081);
or UO_1150 (O_1150,N_12383,N_14156);
nand UO_1151 (O_1151,N_11537,N_14967);
or UO_1152 (O_1152,N_10013,N_13470);
nor UO_1153 (O_1153,N_12048,N_12937);
nor UO_1154 (O_1154,N_13090,N_10762);
nand UO_1155 (O_1155,N_12179,N_13632);
and UO_1156 (O_1156,N_13178,N_12437);
and UO_1157 (O_1157,N_11839,N_13804);
nand UO_1158 (O_1158,N_14816,N_11442);
or UO_1159 (O_1159,N_11530,N_11872);
nand UO_1160 (O_1160,N_14947,N_10600);
and UO_1161 (O_1161,N_10927,N_11024);
and UO_1162 (O_1162,N_13079,N_10804);
and UO_1163 (O_1163,N_14064,N_14334);
nand UO_1164 (O_1164,N_14646,N_11049);
or UO_1165 (O_1165,N_12737,N_14264);
or UO_1166 (O_1166,N_13359,N_12028);
and UO_1167 (O_1167,N_14876,N_11867);
nor UO_1168 (O_1168,N_11828,N_10883);
nand UO_1169 (O_1169,N_12359,N_12994);
or UO_1170 (O_1170,N_14280,N_12418);
nor UO_1171 (O_1171,N_14467,N_13394);
nand UO_1172 (O_1172,N_10968,N_12691);
nor UO_1173 (O_1173,N_14015,N_11623);
nor UO_1174 (O_1174,N_12251,N_13229);
nor UO_1175 (O_1175,N_12707,N_11101);
nand UO_1176 (O_1176,N_12564,N_13530);
or UO_1177 (O_1177,N_14019,N_13294);
nand UO_1178 (O_1178,N_10455,N_12462);
nand UO_1179 (O_1179,N_13084,N_10313);
and UO_1180 (O_1180,N_12392,N_10246);
nand UO_1181 (O_1181,N_12123,N_11328);
and UO_1182 (O_1182,N_14674,N_14921);
xor UO_1183 (O_1183,N_13841,N_14435);
or UO_1184 (O_1184,N_10638,N_11430);
or UO_1185 (O_1185,N_13535,N_12781);
and UO_1186 (O_1186,N_12618,N_12630);
nand UO_1187 (O_1187,N_12974,N_11415);
nor UO_1188 (O_1188,N_13407,N_10739);
nand UO_1189 (O_1189,N_10723,N_11077);
and UO_1190 (O_1190,N_10778,N_13156);
or UO_1191 (O_1191,N_10286,N_11326);
nor UO_1192 (O_1192,N_10181,N_12469);
nor UO_1193 (O_1193,N_13548,N_14680);
xor UO_1194 (O_1194,N_11686,N_14878);
and UO_1195 (O_1195,N_14123,N_10577);
nand UO_1196 (O_1196,N_13633,N_14641);
nand UO_1197 (O_1197,N_13708,N_13367);
and UO_1198 (O_1198,N_10656,N_13132);
nor UO_1199 (O_1199,N_10240,N_12058);
or UO_1200 (O_1200,N_11993,N_13693);
or UO_1201 (O_1201,N_11857,N_12926);
nor UO_1202 (O_1202,N_14146,N_12393);
and UO_1203 (O_1203,N_12662,N_14772);
nor UO_1204 (O_1204,N_10446,N_11948);
and UO_1205 (O_1205,N_14700,N_10045);
nor UO_1206 (O_1206,N_10404,N_10327);
and UO_1207 (O_1207,N_11031,N_10896);
and UO_1208 (O_1208,N_11025,N_13834);
nand UO_1209 (O_1209,N_11106,N_13526);
nand UO_1210 (O_1210,N_13293,N_10772);
nor UO_1211 (O_1211,N_13945,N_12651);
nor UO_1212 (O_1212,N_13423,N_13297);
nor UO_1213 (O_1213,N_12474,N_11005);
nor UO_1214 (O_1214,N_12848,N_10709);
or UO_1215 (O_1215,N_10626,N_12889);
or UO_1216 (O_1216,N_13976,N_10424);
and UO_1217 (O_1217,N_11088,N_13272);
and UO_1218 (O_1218,N_10231,N_13896);
or UO_1219 (O_1219,N_11657,N_10995);
nand UO_1220 (O_1220,N_13616,N_11490);
nor UO_1221 (O_1221,N_10634,N_11710);
or UO_1222 (O_1222,N_14620,N_13533);
or UO_1223 (O_1223,N_14423,N_12338);
nand UO_1224 (O_1224,N_13210,N_12496);
or UO_1225 (O_1225,N_14459,N_10579);
or UO_1226 (O_1226,N_10079,N_13525);
or UO_1227 (O_1227,N_12287,N_12454);
nand UO_1228 (O_1228,N_14063,N_10483);
nor UO_1229 (O_1229,N_10487,N_10326);
nand UO_1230 (O_1230,N_14445,N_14907);
nand UO_1231 (O_1231,N_11249,N_11371);
or UO_1232 (O_1232,N_13758,N_13468);
and UO_1233 (O_1233,N_14971,N_14271);
nand UO_1234 (O_1234,N_12283,N_11174);
nor UO_1235 (O_1235,N_13731,N_12318);
or UO_1236 (O_1236,N_14094,N_10938);
nor UO_1237 (O_1237,N_11275,N_12477);
nand UO_1238 (O_1238,N_10988,N_11340);
nor UO_1239 (O_1239,N_11928,N_14865);
nor UO_1240 (O_1240,N_10459,N_13066);
and UO_1241 (O_1241,N_14635,N_13780);
and UO_1242 (O_1242,N_11066,N_14118);
or UO_1243 (O_1243,N_13231,N_14481);
or UO_1244 (O_1244,N_11662,N_11661);
nor UO_1245 (O_1245,N_11585,N_13815);
nor UO_1246 (O_1246,N_13459,N_10922);
nand UO_1247 (O_1247,N_11043,N_13772);
nor UO_1248 (O_1248,N_12874,N_11048);
and UO_1249 (O_1249,N_10913,N_14328);
nor UO_1250 (O_1250,N_12013,N_11392);
or UO_1251 (O_1251,N_13412,N_11246);
nand UO_1252 (O_1252,N_10704,N_10485);
or UO_1253 (O_1253,N_13986,N_14488);
nand UO_1254 (O_1254,N_14666,N_14844);
nor UO_1255 (O_1255,N_14569,N_12622);
nand UO_1256 (O_1256,N_12162,N_10554);
or UO_1257 (O_1257,N_10258,N_11968);
nor UO_1258 (O_1258,N_13720,N_11429);
nor UO_1259 (O_1259,N_13680,N_11103);
or UO_1260 (O_1260,N_13362,N_12102);
nor UO_1261 (O_1261,N_11699,N_13234);
nor UO_1262 (O_1262,N_12647,N_11469);
and UO_1263 (O_1263,N_14900,N_11955);
and UO_1264 (O_1264,N_12024,N_10385);
nor UO_1265 (O_1265,N_10755,N_11214);
xnor UO_1266 (O_1266,N_12784,N_13093);
and UO_1267 (O_1267,N_14035,N_12995);
nand UO_1268 (O_1268,N_14690,N_14447);
nor UO_1269 (O_1269,N_10532,N_14060);
nor UO_1270 (O_1270,N_11925,N_10528);
or UO_1271 (O_1271,N_12181,N_14644);
nor UO_1272 (O_1272,N_14827,N_13453);
or UO_1273 (O_1273,N_10918,N_10249);
and UO_1274 (O_1274,N_13039,N_13134);
and UO_1275 (O_1275,N_13140,N_12980);
nand UO_1276 (O_1276,N_10285,N_12831);
or UO_1277 (O_1277,N_12319,N_11286);
or UO_1278 (O_1278,N_11863,N_12141);
or UO_1279 (O_1279,N_10243,N_10760);
and UO_1280 (O_1280,N_11349,N_14407);
nor UO_1281 (O_1281,N_12502,N_11463);
nor UO_1282 (O_1282,N_14615,N_10975);
nand UO_1283 (O_1283,N_13760,N_14658);
nand UO_1284 (O_1284,N_12033,N_10563);
or UO_1285 (O_1285,N_11405,N_11179);
and UO_1286 (O_1286,N_10807,N_13865);
and UO_1287 (O_1287,N_11265,N_10498);
and UO_1288 (O_1288,N_10433,N_13390);
xor UO_1289 (O_1289,N_12282,N_11115);
nand UO_1290 (O_1290,N_14923,N_10904);
nor UO_1291 (O_1291,N_12288,N_12021);
nand UO_1292 (O_1292,N_13122,N_13388);
or UO_1293 (O_1293,N_13219,N_14733);
nand UO_1294 (O_1294,N_13242,N_10801);
and UO_1295 (O_1295,N_11574,N_10426);
or UO_1296 (O_1296,N_13183,N_13514);
nor UO_1297 (O_1297,N_13683,N_12612);
xnor UO_1298 (O_1298,N_11142,N_13467);
or UO_1299 (O_1299,N_10027,N_11555);
and UO_1300 (O_1300,N_12925,N_12305);
or UO_1301 (O_1301,N_10270,N_14477);
nand UO_1302 (O_1302,N_11421,N_11681);
xor UO_1303 (O_1303,N_12981,N_11472);
and UO_1304 (O_1304,N_11903,N_14361);
and UO_1305 (O_1305,N_14847,N_14716);
nand UO_1306 (O_1306,N_14166,N_14944);
nor UO_1307 (O_1307,N_10085,N_14084);
and UO_1308 (O_1308,N_12689,N_14728);
nor UO_1309 (O_1309,N_12780,N_13572);
nand UO_1310 (O_1310,N_13175,N_10332);
and UO_1311 (O_1311,N_14643,N_12022);
or UO_1312 (O_1312,N_10535,N_10892);
or UO_1313 (O_1313,N_12957,N_12699);
or UO_1314 (O_1314,N_11495,N_11255);
or UO_1315 (O_1315,N_11644,N_13596);
nand UO_1316 (O_1316,N_14984,N_11992);
and UO_1317 (O_1317,N_13762,N_10905);
nand UO_1318 (O_1318,N_10567,N_14521);
and UO_1319 (O_1319,N_13504,N_10639);
and UO_1320 (O_1320,N_10917,N_11524);
or UO_1321 (O_1321,N_13267,N_10428);
nor UO_1322 (O_1322,N_14834,N_13779);
nand UO_1323 (O_1323,N_13713,N_13444);
nor UO_1324 (O_1324,N_13157,N_11395);
nand UO_1325 (O_1325,N_12384,N_13327);
nand UO_1326 (O_1326,N_12230,N_14398);
nand UO_1327 (O_1327,N_14648,N_10105);
nand UO_1328 (O_1328,N_12441,N_11449);
nor UO_1329 (O_1329,N_14053,N_10856);
or UO_1330 (O_1330,N_13990,N_13196);
and UO_1331 (O_1331,N_12575,N_14148);
and UO_1332 (O_1332,N_14987,N_11703);
or UO_1333 (O_1333,N_10114,N_13667);
and UO_1334 (O_1334,N_13684,N_12381);
and UO_1335 (O_1335,N_12825,N_10659);
or UO_1336 (O_1336,N_13848,N_11624);
and UO_1337 (O_1337,N_10622,N_13598);
nor UO_1338 (O_1338,N_13413,N_14830);
nor UO_1339 (O_1339,N_11321,N_14576);
or UO_1340 (O_1340,N_11909,N_13166);
and UO_1341 (O_1341,N_10982,N_12886);
or UO_1342 (O_1342,N_14121,N_10479);
or UO_1343 (O_1343,N_11630,N_12979);
nor UO_1344 (O_1344,N_14369,N_12365);
nand UO_1345 (O_1345,N_14429,N_10383);
or UO_1346 (O_1346,N_14323,N_12900);
or UO_1347 (O_1347,N_13957,N_12652);
nand UO_1348 (O_1348,N_13729,N_10195);
nand UO_1349 (O_1349,N_14711,N_10598);
nor UO_1350 (O_1350,N_12308,N_12280);
nand UO_1351 (O_1351,N_12741,N_10994);
nor UO_1352 (O_1352,N_13226,N_12264);
and UO_1353 (O_1353,N_14052,N_10819);
and UO_1354 (O_1354,N_12548,N_12565);
and UO_1355 (O_1355,N_13927,N_14333);
nor UO_1356 (O_1356,N_10830,N_10268);
and UO_1357 (O_1357,N_14818,N_14599);
or UO_1358 (O_1358,N_14137,N_13198);
and UO_1359 (O_1359,N_14479,N_10138);
nor UO_1360 (O_1360,N_10188,N_10777);
nand UO_1361 (O_1361,N_12534,N_12774);
nand UO_1362 (O_1362,N_10674,N_13790);
nor UO_1363 (O_1363,N_13591,N_13997);
nor UO_1364 (O_1364,N_12770,N_14845);
or UO_1365 (O_1365,N_12918,N_14536);
nor UO_1366 (O_1366,N_14211,N_12110);
nand UO_1367 (O_1367,N_11746,N_12892);
nand UO_1368 (O_1368,N_10473,N_14414);
nor UO_1369 (O_1369,N_11479,N_11280);
nand UO_1370 (O_1370,N_11902,N_10960);
nor UO_1371 (O_1371,N_12174,N_10891);
nor UO_1372 (O_1372,N_12671,N_12198);
or UO_1373 (O_1373,N_14529,N_13190);
and UO_1374 (O_1374,N_10064,N_12060);
nand UO_1375 (O_1375,N_11003,N_11967);
nand UO_1376 (O_1376,N_11420,N_10516);
nor UO_1377 (O_1377,N_14926,N_14668);
nand UO_1378 (O_1378,N_10215,N_10570);
or UO_1379 (O_1379,N_14018,N_14851);
and UO_1380 (O_1380,N_10644,N_14024);
or UO_1381 (O_1381,N_12556,N_11477);
or UO_1382 (O_1382,N_10331,N_12751);
nand UO_1383 (O_1383,N_11824,N_14897);
and UO_1384 (O_1384,N_14448,N_12140);
nand UO_1385 (O_1385,N_14492,N_12897);
nor UO_1386 (O_1386,N_13658,N_12559);
and UO_1387 (O_1387,N_10322,N_11795);
or UO_1388 (O_1388,N_10037,N_14169);
nor UO_1389 (O_1389,N_10189,N_10269);
nor UO_1390 (O_1390,N_10191,N_10505);
nand UO_1391 (O_1391,N_12072,N_12232);
and UO_1392 (O_1392,N_13264,N_13542);
and UO_1393 (O_1393,N_14740,N_14573);
or UO_1394 (O_1394,N_12987,N_12442);
nand UO_1395 (O_1395,N_10682,N_11131);
nand UO_1396 (O_1396,N_11764,N_11952);
or UO_1397 (O_1397,N_14636,N_13315);
nor UO_1398 (O_1398,N_13853,N_14920);
or UO_1399 (O_1399,N_10417,N_11700);
or UO_1400 (O_1400,N_12239,N_14685);
nand UO_1401 (O_1401,N_13755,N_14105);
nand UO_1402 (O_1402,N_11947,N_11941);
or UO_1403 (O_1403,N_11873,N_11143);
nor UO_1404 (O_1404,N_10196,N_12641);
and UO_1405 (O_1405,N_14017,N_12772);
and UO_1406 (O_1406,N_12791,N_11170);
nand UO_1407 (O_1407,N_11584,N_13821);
nor UO_1408 (O_1408,N_10376,N_11958);
xnor UO_1409 (O_1409,N_14586,N_14223);
nand UO_1410 (O_1410,N_11119,N_14471);
nor UO_1411 (O_1411,N_11822,N_12759);
or UO_1412 (O_1412,N_10281,N_13016);
nor UO_1413 (O_1413,N_13740,N_11961);
or UO_1414 (O_1414,N_14623,N_10853);
or UO_1415 (O_1415,N_11338,N_10658);
nor UO_1416 (O_1416,N_11207,N_12009);
nand UO_1417 (O_1417,N_10761,N_10550);
or UO_1418 (O_1418,N_13030,N_11500);
xor UO_1419 (O_1419,N_10158,N_11046);
nand UO_1420 (O_1420,N_13235,N_12449);
or UO_1421 (O_1421,N_10226,N_12193);
nor UO_1422 (O_1422,N_10635,N_12794);
and UO_1423 (O_1423,N_10355,N_14082);
or UO_1424 (O_1424,N_10699,N_14744);
or UO_1425 (O_1425,N_10292,N_12397);
nand UO_1426 (O_1426,N_10829,N_11739);
nor UO_1427 (O_1427,N_12730,N_13279);
nand UO_1428 (O_1428,N_10469,N_11721);
and UO_1429 (O_1429,N_13922,N_14588);
or UO_1430 (O_1430,N_11052,N_14194);
xnor UO_1431 (O_1431,N_12962,N_13286);
nor UO_1432 (O_1432,N_12726,N_10867);
nand UO_1433 (O_1433,N_10374,N_11041);
xor UO_1434 (O_1434,N_11540,N_10970);
nor UO_1435 (O_1435,N_10566,N_10513);
or UO_1436 (O_1436,N_11050,N_10732);
and UO_1437 (O_1437,N_13768,N_13256);
or UO_1438 (O_1438,N_13191,N_10798);
nor UO_1439 (O_1439,N_10150,N_12783);
and UO_1440 (O_1440,N_14373,N_11242);
xor UO_1441 (O_1441,N_12087,N_10319);
and UO_1442 (O_1442,N_11940,N_12661);
nor UO_1443 (O_1443,N_14879,N_13450);
or UO_1444 (O_1444,N_13726,N_11794);
nand UO_1445 (O_1445,N_10832,N_13047);
nor UO_1446 (O_1446,N_10886,N_13082);
or UO_1447 (O_1447,N_14743,N_11154);
and UO_1448 (O_1448,N_11826,N_13950);
nor UO_1449 (O_1449,N_11815,N_14426);
nand UO_1450 (O_1450,N_11768,N_12627);
nor UO_1451 (O_1451,N_13089,N_13251);
nand UO_1452 (O_1452,N_14230,N_10334);
nand UO_1453 (O_1453,N_11030,N_14859);
and UO_1454 (O_1454,N_12236,N_13062);
nor UO_1455 (O_1455,N_11665,N_14292);
and UO_1456 (O_1456,N_10000,N_10782);
nand UO_1457 (O_1457,N_10854,N_14188);
or UO_1458 (O_1458,N_13322,N_10595);
and UO_1459 (O_1459,N_14268,N_11305);
and UO_1460 (O_1460,N_14026,N_14708);
and UO_1461 (O_1461,N_13570,N_11181);
and UO_1462 (O_1462,N_11564,N_10714);
nand UO_1463 (O_1463,N_11446,N_11899);
nand UO_1464 (O_1464,N_13354,N_13867);
nor UO_1465 (O_1465,N_10821,N_10879);
nor UO_1466 (O_1466,N_14180,N_13689);
xor UO_1467 (O_1467,N_10643,N_14549);
and UO_1468 (O_1468,N_12948,N_12929);
or UO_1469 (O_1469,N_13377,N_13972);
nand UO_1470 (O_1470,N_13351,N_12426);
and UO_1471 (O_1471,N_11488,N_13310);
and UO_1472 (O_1472,N_14460,N_12906);
and UO_1473 (O_1473,N_14389,N_11057);
nand UO_1474 (O_1474,N_14562,N_10342);
nor UO_1475 (O_1475,N_14494,N_11162);
and UO_1476 (O_1476,N_14715,N_12674);
nor UO_1477 (O_1477,N_10074,N_11373);
nand UO_1478 (O_1478,N_11673,N_14969);
nand UO_1479 (O_1479,N_12175,N_14843);
nor UO_1480 (O_1480,N_12491,N_12323);
nand UO_1481 (O_1481,N_12968,N_13828);
nand UO_1482 (O_1482,N_11453,N_14192);
nand UO_1483 (O_1483,N_10583,N_13682);
and UO_1484 (O_1484,N_10751,N_14014);
nand UO_1485 (O_1485,N_12309,N_10944);
or UO_1486 (O_1486,N_14240,N_13600);
and UO_1487 (O_1487,N_11930,N_10784);
and UO_1488 (O_1488,N_12160,N_13381);
and UO_1489 (O_1489,N_13610,N_12164);
nand UO_1490 (O_1490,N_13983,N_14403);
nand UO_1491 (O_1491,N_10612,N_14931);
nor UO_1492 (O_1492,N_13982,N_10518);
nand UO_1493 (O_1493,N_12398,N_11923);
nor UO_1494 (O_1494,N_11641,N_11637);
or UO_1495 (O_1495,N_13487,N_12145);
or UO_1496 (O_1496,N_14134,N_14420);
nor UO_1497 (O_1497,N_11262,N_12745);
nand UO_1498 (O_1498,N_11071,N_11164);
nor UO_1499 (O_1499,N_14344,N_10078);
and UO_1500 (O_1500,N_10802,N_10311);
nand UO_1501 (O_1501,N_11206,N_11977);
or UO_1502 (O_1502,N_13544,N_13368);
nand UO_1503 (O_1503,N_10369,N_14968);
nor UO_1504 (O_1504,N_10401,N_12541);
nor UO_1505 (O_1505,N_13428,N_11304);
xor UO_1506 (O_1506,N_13307,N_13105);
nand UO_1507 (O_1507,N_11885,N_13223);
nand UO_1508 (O_1508,N_11904,N_14855);
or UO_1509 (O_1509,N_10155,N_11814);
nor UO_1510 (O_1510,N_14476,N_12211);
nor UO_1511 (O_1511,N_13851,N_10454);
or UO_1512 (O_1512,N_13655,N_12291);
nand UO_1513 (O_1513,N_14889,N_13224);
and UO_1514 (O_1514,N_13011,N_12328);
and UO_1515 (O_1515,N_14712,N_11577);
nor UO_1516 (O_1516,N_13775,N_14037);
or UO_1517 (O_1517,N_13041,N_14183);
nand UO_1518 (O_1518,N_11013,N_12596);
nor UO_1519 (O_1519,N_13966,N_12385);
and UO_1520 (O_1520,N_13274,N_10122);
and UO_1521 (O_1521,N_12467,N_14385);
and UO_1522 (O_1522,N_11647,N_14667);
nor UO_1523 (O_1523,N_13484,N_13332);
and UO_1524 (O_1524,N_11374,N_12404);
and UO_1525 (O_1525,N_10688,N_13710);
nand UO_1526 (O_1526,N_14000,N_14877);
or UO_1527 (O_1527,N_14274,N_14308);
or UO_1528 (O_1528,N_10255,N_13826);
and UO_1529 (O_1529,N_13811,N_10082);
nand UO_1530 (O_1530,N_13455,N_13885);
and UO_1531 (O_1531,N_12245,N_11718);
nand UO_1532 (O_1532,N_13385,N_10966);
nand UO_1533 (O_1533,N_13441,N_13724);
or UO_1534 (O_1534,N_11841,N_14811);
or UO_1535 (O_1535,N_14785,N_10582);
nand UO_1536 (O_1536,N_11117,N_13663);
nand UO_1537 (O_1537,N_12356,N_11318);
or UO_1538 (O_1538,N_10237,N_13761);
and UO_1539 (O_1539,N_12978,N_14954);
nor UO_1540 (O_1540,N_10199,N_11378);
and UO_1541 (O_1541,N_11747,N_14937);
or UO_1542 (O_1542,N_11390,N_12314);
nand UO_1543 (O_1543,N_13836,N_11014);
nor UO_1544 (O_1544,N_11361,N_13479);
nor UO_1545 (O_1545,N_12782,N_11409);
or UO_1546 (O_1546,N_11683,N_12513);
and UO_1547 (O_1547,N_12669,N_11094);
nand UO_1548 (O_1548,N_10408,N_11697);
nor UO_1549 (O_1549,N_14281,N_12859);
nor UO_1550 (O_1550,N_13559,N_14709);
xnor UO_1551 (O_1551,N_14149,N_10887);
nor UO_1552 (O_1552,N_11270,N_10256);
nand UO_1553 (O_1553,N_11266,N_14287);
nand UO_1554 (O_1554,N_11079,N_13439);
and UO_1555 (O_1555,N_13313,N_10584);
or UO_1556 (O_1556,N_12458,N_10561);
or UO_1557 (O_1557,N_11973,N_13034);
or UO_1558 (O_1558,N_14885,N_14251);
nand UO_1559 (O_1559,N_14717,N_13049);
nor UO_1560 (O_1560,N_12778,N_12971);
nand UO_1561 (O_1561,N_14795,N_11855);
or UO_1562 (O_1562,N_11819,N_13917);
and UO_1563 (O_1563,N_12752,N_14421);
and UO_1564 (O_1564,N_13000,N_14051);
nand UO_1565 (O_1565,N_11447,N_11888);
nor UO_1566 (O_1566,N_12074,N_10252);
or UO_1567 (O_1567,N_10323,N_10506);
or UO_1568 (O_1568,N_11660,N_10517);
or UO_1569 (O_1569,N_14558,N_10512);
nor UO_1570 (O_1570,N_11934,N_14630);
and UO_1571 (O_1571,N_11337,N_13685);
or UO_1572 (O_1572,N_14154,N_10525);
nor UO_1573 (O_1573,N_12046,N_10764);
nor UO_1574 (O_1574,N_14349,N_14724);
and UO_1575 (O_1575,N_10368,N_12928);
nand UO_1576 (O_1576,N_11327,N_10496);
and UO_1577 (O_1577,N_10893,N_13073);
nand UO_1578 (O_1578,N_13373,N_11028);
nand UO_1579 (O_1579,N_12005,N_10825);
nor UO_1580 (O_1580,N_14474,N_13547);
or UO_1581 (O_1581,N_11991,N_12407);
and UO_1582 (O_1582,N_10676,N_12911);
nand UO_1583 (O_1583,N_12961,N_13065);
or UO_1584 (O_1584,N_13860,N_14364);
and UO_1585 (O_1585,N_10868,N_14140);
nand UO_1586 (O_1586,N_13018,N_11352);
nand UO_1587 (O_1587,N_12010,N_13576);
xnor UO_1588 (O_1588,N_12075,N_11258);
nor UO_1589 (O_1589,N_14210,N_14670);
or UO_1590 (O_1590,N_12724,N_14895);
nand UO_1591 (O_1591,N_14617,N_10099);
nand UO_1592 (O_1592,N_14265,N_12958);
and UO_1593 (O_1593,N_14916,N_10072);
nand UO_1594 (O_1594,N_12395,N_13750);
nor UO_1595 (O_1595,N_10330,N_11512);
or UO_1596 (O_1596,N_10177,N_12224);
and UO_1597 (O_1597,N_10964,N_13617);
nand UO_1598 (O_1598,N_13973,N_14219);
nor UO_1599 (O_1599,N_12576,N_10008);
and UO_1600 (O_1600,N_12340,N_10773);
or UO_1601 (O_1601,N_10477,N_13756);
nor UO_1602 (O_1602,N_10135,N_14030);
or UO_1603 (O_1603,N_11596,N_11622);
and UO_1604 (O_1604,N_13181,N_13727);
or UO_1605 (O_1605,N_14113,N_12614);
nor UO_1606 (O_1606,N_10780,N_12685);
and UO_1607 (O_1607,N_14684,N_10004);
or UO_1608 (O_1608,N_12302,N_13401);
nor UO_1609 (O_1609,N_14279,N_13622);
nand UO_1610 (O_1610,N_13995,N_14008);
nand UO_1611 (O_1611,N_12818,N_14002);
or UO_1612 (O_1612,N_11277,N_14056);
nor UO_1613 (O_1613,N_13275,N_14802);
or UO_1614 (O_1614,N_10952,N_14750);
or UO_1615 (O_1615,N_12890,N_12735);
nor UO_1616 (O_1616,N_12952,N_14551);
nor UO_1617 (O_1617,N_10279,N_12275);
nand UO_1618 (O_1618,N_13028,N_10381);
and UO_1619 (O_1619,N_11552,N_11694);
and UO_1620 (O_1620,N_14760,N_13495);
nor UO_1621 (O_1621,N_11594,N_11336);
nand UO_1622 (O_1622,N_12240,N_14697);
nor UO_1623 (O_1623,N_11553,N_10675);
and UO_1624 (O_1624,N_10767,N_13179);
nand UO_1625 (O_1625,N_14092,N_13527);
nand UO_1626 (O_1626,N_11388,N_13371);
nand UO_1627 (O_1627,N_10147,N_14714);
and UO_1628 (O_1628,N_10005,N_11844);
nand UO_1629 (O_1629,N_12157,N_14748);
nor UO_1630 (O_1630,N_11271,N_12170);
and UO_1631 (O_1631,N_12768,N_10373);
nand UO_1632 (O_1632,N_10447,N_13796);
nand UO_1633 (O_1633,N_12914,N_13379);
nor UO_1634 (O_1634,N_10906,N_12519);
nand UO_1635 (O_1635,N_10947,N_11439);
or UO_1636 (O_1636,N_14320,N_13909);
or UO_1637 (O_1637,N_13162,N_13614);
and UO_1638 (O_1638,N_14722,N_12073);
or UO_1639 (O_1639,N_14842,N_14491);
nor UO_1640 (O_1640,N_13476,N_10903);
or UO_1641 (O_1641,N_12803,N_10728);
or UO_1642 (O_1642,N_13550,N_12749);
and UO_1643 (O_1643,N_13977,N_11675);
nand UO_1644 (O_1644,N_11368,N_12168);
nand UO_1645 (O_1645,N_12593,N_14513);
or UO_1646 (O_1646,N_10998,N_13552);
and UO_1647 (O_1647,N_11456,N_10460);
nand UO_1648 (O_1648,N_14698,N_14317);
or UO_1649 (O_1649,N_13777,N_14221);
nor UO_1650 (O_1650,N_14852,N_14787);
nand UO_1651 (O_1651,N_13490,N_14297);
or UO_1652 (O_1652,N_10217,N_13919);
nand UO_1653 (O_1653,N_14933,N_12344);
and UO_1654 (O_1654,N_12697,N_14451);
or UO_1655 (O_1655,N_14444,N_12748);
xor UO_1656 (O_1656,N_10015,N_13691);
and UO_1657 (O_1657,N_11357,N_12827);
nand UO_1658 (O_1658,N_13103,N_12218);
or UO_1659 (O_1659,N_11341,N_12740);
nor UO_1660 (O_1660,N_14249,N_12261);
nand UO_1661 (O_1661,N_10328,N_13822);
or UO_1662 (O_1662,N_13694,N_13160);
nand UO_1663 (O_1663,N_13714,N_11462);
nand UO_1664 (O_1664,N_12263,N_14530);
nor UO_1665 (O_1665,N_10705,N_12700);
nor UO_1666 (O_1666,N_12955,N_12754);
or UO_1667 (O_1667,N_14404,N_13424);
nor UO_1668 (O_1668,N_12199,N_11551);
nand UO_1669 (O_1669,N_12255,N_12433);
and UO_1670 (O_1670,N_11796,N_13579);
and UO_1671 (O_1671,N_13959,N_11684);
and UO_1672 (O_1672,N_11032,N_13262);
or UO_1673 (O_1673,N_12436,N_14782);
or UO_1674 (O_1674,N_10686,N_13395);
or UO_1675 (O_1675,N_12659,N_12853);
nor UO_1676 (O_1676,N_10272,N_11592);
or UO_1677 (O_1677,N_10703,N_13523);
and UO_1678 (O_1678,N_12144,N_10673);
nand UO_1679 (O_1679,N_13142,N_12909);
nand UO_1680 (O_1680,N_12521,N_10450);
nor UO_1681 (O_1681,N_12482,N_11108);
or UO_1682 (O_1682,N_10701,N_14184);
nand UO_1683 (O_1683,N_10108,N_12779);
or UO_1684 (O_1684,N_11296,N_11135);
or UO_1685 (O_1685,N_11084,N_14762);
and UO_1686 (O_1686,N_10531,N_14882);
and UO_1687 (O_1687,N_11515,N_12345);
or UO_1688 (O_1688,N_14012,N_10981);
nor UO_1689 (O_1689,N_10859,N_13117);
nor UO_1690 (O_1690,N_14622,N_11648);
nand UO_1691 (O_1691,N_13420,N_10953);
nor UO_1692 (O_1692,N_12335,N_14790);
nor UO_1693 (O_1693,N_10388,N_13872);
nor UO_1694 (O_1694,N_11711,N_13566);
nor UO_1695 (O_1695,N_12452,N_13532);
nor UO_1696 (O_1696,N_14306,N_12371);
and UO_1697 (O_1697,N_10358,N_12188);
or UO_1698 (O_1698,N_13562,N_11138);
or UO_1699 (O_1699,N_10611,N_13660);
or UO_1700 (O_1700,N_13810,N_11587);
and UO_1701 (O_1701,N_11847,N_10471);
nand UO_1702 (O_1702,N_14746,N_12146);
or UO_1703 (O_1703,N_13607,N_14980);
nor UO_1704 (O_1704,N_12158,N_10372);
nand UO_1705 (O_1705,N_12410,N_14458);
nand UO_1706 (O_1706,N_10544,N_11263);
nor UO_1707 (O_1707,N_13305,N_10157);
nor UO_1708 (O_1708,N_10363,N_12856);
and UO_1709 (O_1709,N_14485,N_14438);
nor UO_1710 (O_1710,N_13666,N_11938);
and UO_1711 (O_1711,N_11994,N_11590);
and UO_1712 (O_1712,N_13733,N_11126);
and UO_1713 (O_1713,N_11334,N_10209);
and UO_1714 (O_1714,N_13475,N_14880);
and UO_1715 (O_1715,N_12234,N_14591);
nand UO_1716 (O_1716,N_14358,N_10538);
and UO_1717 (O_1717,N_12695,N_10031);
or UO_1718 (O_1718,N_14001,N_13400);
nor UO_1719 (O_1719,N_12919,N_10380);
nand UO_1720 (O_1720,N_14098,N_14862);
nor UO_1721 (O_1721,N_14266,N_11455);
or UO_1722 (O_1722,N_11781,N_11864);
and UO_1723 (O_1723,N_11010,N_10356);
nand UO_1724 (O_1724,N_14173,N_10657);
and UO_1725 (O_1725,N_12664,N_13116);
nand UO_1726 (O_1726,N_14501,N_11559);
xnor UO_1727 (O_1727,N_14233,N_12330);
nor UO_1728 (O_1728,N_13259,N_14122);
and UO_1729 (O_1729,N_14353,N_13329);
or UO_1730 (O_1730,N_10020,N_10305);
nor UO_1731 (O_1731,N_14682,N_11228);
nor UO_1732 (O_1732,N_11158,N_11232);
or UO_1733 (O_1733,N_14934,N_13447);
or UO_1734 (O_1734,N_12846,N_12785);
nand UO_1735 (O_1735,N_13285,N_13730);
and UO_1736 (O_1736,N_13903,N_11996);
or UO_1737 (O_1737,N_13875,N_13791);
nand UO_1738 (O_1738,N_13638,N_14372);
and UO_1739 (O_1739,N_11377,N_12343);
or UO_1740 (O_1740,N_10581,N_11932);
and UO_1741 (O_1741,N_11616,N_10262);
or UO_1742 (O_1742,N_12434,N_11201);
or UO_1743 (O_1743,N_11547,N_11197);
nand UO_1744 (O_1744,N_11728,N_13868);
or UO_1745 (O_1745,N_11440,N_14201);
and UO_1746 (O_1746,N_13554,N_14508);
or UO_1747 (O_1747,N_14135,N_11380);
or UO_1748 (O_1748,N_10480,N_11293);
nor UO_1749 (O_1749,N_12598,N_13657);
or UO_1750 (O_1750,N_14973,N_12977);
nand UO_1751 (O_1751,N_13545,N_14911);
nand UO_1752 (O_1752,N_11489,N_10603);
nand UO_1753 (O_1753,N_14193,N_13911);
nand UO_1754 (O_1754,N_11504,N_11791);
and UO_1755 (O_1755,N_12509,N_14196);
nand UO_1756 (O_1756,N_14157,N_13228);
or UO_1757 (O_1757,N_14624,N_11465);
nand UO_1758 (O_1758,N_11152,N_13207);
and UO_1759 (O_1759,N_14163,N_13507);
nor UO_1760 (O_1760,N_10788,N_14005);
and UO_1761 (O_1761,N_13350,N_10668);
nor UO_1762 (O_1762,N_12408,N_13375);
nor UO_1763 (O_1763,N_10923,N_12861);
and UO_1764 (O_1764,N_10813,N_13974);
nor UO_1765 (O_1765,N_13057,N_13671);
or UO_1766 (O_1766,N_11067,N_14436);
and UO_1767 (O_1767,N_12394,N_13845);
nor UO_1768 (O_1768,N_10444,N_14976);
nor UO_1769 (O_1769,N_10185,N_10809);
nand UO_1770 (O_1770,N_13521,N_13227);
and UO_1771 (O_1771,N_10507,N_11339);
or UO_1772 (O_1772,N_10909,N_11476);
or UO_1773 (O_1773,N_12836,N_11012);
or UO_1774 (O_1774,N_13378,N_10828);
nor UO_1775 (O_1775,N_12014,N_10067);
or UO_1776 (O_1776,N_13595,N_10742);
nand UO_1777 (O_1777,N_12054,N_14678);
nand UO_1778 (O_1778,N_11521,N_11556);
nor UO_1779 (O_1779,N_11793,N_13723);
or UO_1780 (O_1780,N_14440,N_10621);
and UO_1781 (O_1781,N_12755,N_10456);
and UO_1782 (O_1782,N_11542,N_10522);
or UO_1783 (O_1783,N_10707,N_12353);
nand UO_1784 (O_1784,N_11538,N_14250);
nor UO_1785 (O_1785,N_13669,N_14819);
nor UO_1786 (O_1786,N_13895,N_11034);
or UO_1787 (O_1787,N_10139,N_12321);
or UO_1788 (O_1788,N_13172,N_14095);
nor UO_1789 (O_1789,N_10743,N_10860);
nand UO_1790 (O_1790,N_13301,N_14803);
nand UO_1791 (O_1791,N_13492,N_13692);
or UO_1792 (O_1792,N_12855,N_10137);
nand UO_1793 (O_1793,N_14922,N_12026);
nor UO_1794 (O_1794,N_11322,N_13699);
and UO_1795 (O_1795,N_10129,N_10070);
or UO_1796 (O_1796,N_12351,N_14910);
nor UO_1797 (O_1797,N_11954,N_10484);
or UO_1798 (O_1798,N_13933,N_12904);
or UO_1799 (O_1799,N_14831,N_14902);
and UO_1800 (O_1800,N_10035,N_14532);
or UO_1801 (O_1801,N_13861,N_13128);
nand UO_1802 (O_1802,N_14072,N_12682);
nand UO_1803 (O_1803,N_11384,N_13037);
nor UO_1804 (O_1804,N_12432,N_14701);
or UO_1805 (O_1805,N_10847,N_13899);
or UO_1806 (O_1806,N_13676,N_14777);
or UO_1807 (O_1807,N_13180,N_11918);
nor UO_1808 (O_1808,N_10338,N_14689);
nor UO_1809 (O_1809,N_10521,N_11260);
nand UO_1810 (O_1810,N_13195,N_13873);
and UO_1811 (O_1811,N_12195,N_14003);
nand UO_1812 (O_1812,N_14775,N_13460);
and UO_1813 (O_1813,N_14057,N_13553);
nand UO_1814 (O_1814,N_10354,N_10043);
nand UO_1815 (O_1815,N_11055,N_10398);
nor UO_1816 (O_1816,N_13580,N_11302);
nand UO_1817 (O_1817,N_14525,N_14629);
or UO_1818 (O_1818,N_11400,N_11021);
nor UO_1819 (O_1819,N_13425,N_11150);
nor UO_1820 (O_1820,N_12815,N_13817);
and UO_1821 (O_1821,N_10219,N_12213);
nand UO_1822 (O_1822,N_12390,N_10392);
or UO_1823 (O_1823,N_11862,N_11895);
or UO_1824 (O_1824,N_14886,N_13389);
or UO_1825 (O_1825,N_14174,N_11581);
nor UO_1826 (O_1826,N_10300,N_12068);
or UO_1827 (O_1827,N_11160,N_13955);
or UO_1828 (O_1828,N_10024,N_10192);
or UO_1829 (O_1829,N_10364,N_11253);
or UO_1830 (O_1830,N_11087,N_12093);
nand UO_1831 (O_1831,N_11913,N_13015);
or UO_1832 (O_1832,N_14258,N_12687);
nand UO_1833 (O_1833,N_11183,N_13820);
or UO_1834 (O_1834,N_14541,N_12324);
nor UO_1835 (O_1835,N_13240,N_14948);
nand UO_1836 (O_1836,N_10594,N_14725);
nor UO_1837 (O_1837,N_10636,N_14567);
and UO_1838 (O_1838,N_12192,N_11096);
nor UO_1839 (O_1839,N_13588,N_14412);
nand UO_1840 (O_1840,N_11756,N_13891);
nor UO_1841 (O_1841,N_10697,N_13361);
nand UO_1842 (O_1842,N_14117,N_13643);
nor UO_1843 (O_1843,N_10529,N_13209);
xor UO_1844 (O_1844,N_10669,N_12954);
nand UO_1845 (O_1845,N_14282,N_13083);
or UO_1846 (O_1846,N_12226,N_14978);
or UO_1847 (O_1847,N_10391,N_12267);
nor UO_1848 (O_1848,N_12018,N_14362);
or UO_1849 (O_1849,N_10216,N_12080);
or UO_1850 (O_1850,N_14789,N_12182);
and UO_1851 (O_1851,N_13025,N_14378);
nor UO_1852 (O_1852,N_10588,N_10503);
and UO_1853 (O_1853,N_13247,N_12209);
or UO_1854 (O_1854,N_10748,N_11437);
and UO_1855 (O_1855,N_11107,N_14780);
nand UO_1856 (O_1856,N_12429,N_13001);
nand UO_1857 (O_1857,N_13506,N_12723);
or UO_1858 (O_1858,N_11299,N_10163);
and UO_1859 (O_1859,N_10234,N_12616);
and UO_1860 (O_1860,N_12346,N_13435);
nor UO_1861 (O_1861,N_12450,N_11572);
nand UO_1862 (O_1862,N_12850,N_13314);
or UO_1863 (O_1863,N_11173,N_11061);
and UO_1864 (O_1864,N_12512,N_12473);
nor UO_1865 (O_1865,N_11269,N_14336);
and UO_1866 (O_1866,N_13036,N_10562);
nand UO_1867 (O_1867,N_12875,N_10400);
and UO_1868 (O_1868,N_13265,N_12488);
nand UO_1869 (O_1869,N_13908,N_12217);
nor UO_1870 (O_1870,N_13984,N_12151);
or UO_1871 (O_1871,N_13215,N_12561);
nor UO_1872 (O_1872,N_10967,N_12602);
nand UO_1873 (O_1873,N_12646,N_12278);
or UO_1874 (O_1874,N_12629,N_11111);
nand UO_1875 (O_1875,N_13798,N_13921);
nor UO_1876 (O_1876,N_14143,N_14405);
nor UO_1877 (O_1877,N_12800,N_14736);
and UO_1878 (O_1878,N_12869,N_10954);
nor UO_1879 (O_1879,N_10568,N_11090);
and UO_1880 (O_1880,N_14182,N_12292);
nand UO_1881 (O_1881,N_13392,N_10831);
nand UO_1882 (O_1882,N_13967,N_11175);
and UO_1883 (O_1883,N_10395,N_13674);
or UO_1884 (O_1884,N_13893,N_14741);
or UO_1885 (O_1885,N_12943,N_14215);
nand UO_1886 (O_1886,N_10663,N_12572);
and UO_1887 (O_1887,N_10134,N_10259);
or UO_1888 (O_1888,N_11859,N_10837);
nand UO_1889 (O_1889,N_14124,N_13602);
nand UO_1890 (O_1890,N_12235,N_11567);
or UO_1891 (O_1891,N_11140,N_12920);
nor UO_1892 (O_1892,N_14046,N_12161);
and UO_1893 (O_1893,N_12984,N_11926);
and UO_1894 (O_1894,N_14706,N_12388);
or UO_1895 (O_1895,N_12567,N_11732);
or UO_1896 (O_1896,N_10786,N_13052);
and UO_1897 (O_1897,N_14463,N_10915);
and UO_1898 (O_1898,N_14512,N_13739);
nand UO_1899 (O_1899,N_12253,N_10316);
nand UO_1900 (O_1900,N_10962,N_11288);
and UO_1901 (O_1901,N_12888,N_11078);
nor UO_1902 (O_1902,N_13045,N_12789);
and UO_1903 (O_1903,N_10429,N_12373);
nor UO_1904 (O_1904,N_11452,N_10390);
nor UO_1905 (O_1905,N_12879,N_10519);
and UO_1906 (O_1906,N_14262,N_14990);
or UO_1907 (O_1907,N_13862,N_11692);
or UO_1908 (O_1908,N_12260,N_10556);
nand UO_1909 (O_1909,N_13220,N_11239);
and UO_1910 (O_1910,N_13586,N_14655);
nor UO_1911 (O_1911,N_10212,N_13485);
and UO_1912 (O_1912,N_14074,N_13056);
or UO_1913 (O_1913,N_13040,N_14241);
nand UO_1914 (O_1914,N_12552,N_11907);
xor UO_1915 (O_1915,N_10438,N_12416);
and UO_1916 (O_1916,N_13480,N_11980);
or UO_1917 (O_1917,N_10497,N_13624);
or UO_1918 (O_1918,N_14598,N_13854);
or UO_1919 (O_1919,N_14214,N_13493);
nor UO_1920 (O_1920,N_11678,N_10208);
nor UO_1921 (O_1921,N_10307,N_14884);
or UO_1922 (O_1922,N_12637,N_14204);
and UO_1923 (O_1923,N_10537,N_14054);
nor UO_1924 (O_1924,N_13864,N_11220);
and UO_1925 (O_1925,N_12327,N_14784);
nand UO_1926 (O_1926,N_10548,N_11454);
nor UO_1927 (O_1927,N_11350,N_13081);
or UO_1928 (O_1928,N_13803,N_11829);
nand UO_1929 (O_1929,N_10932,N_12528);
nor UO_1930 (O_1930,N_14856,N_14424);
nor UO_1931 (O_1931,N_13904,N_11076);
nand UO_1932 (O_1932,N_10817,N_13601);
or UO_1933 (O_1933,N_10606,N_13589);
nor UO_1934 (O_1934,N_11836,N_10820);
nor UO_1935 (O_1935,N_13360,N_14894);
and UO_1936 (O_1936,N_10365,N_10055);
or UO_1937 (O_1937,N_13941,N_12481);
or UO_1938 (O_1938,N_13604,N_11291);
nor UO_1939 (O_1939,N_10453,N_12424);
and UO_1940 (O_1940,N_12417,N_10741);
nand UO_1941 (O_1941,N_13437,N_12706);
nor UO_1942 (O_1942,N_12055,N_12095);
and UO_1943 (O_1943,N_11827,N_13665);
or UO_1944 (O_1944,N_13703,N_13574);
and UO_1945 (O_1945,N_11134,N_11736);
nand UO_1946 (O_1946,N_10991,N_13462);
and UO_1947 (O_1947,N_11969,N_11525);
nand UO_1948 (O_1948,N_13023,N_12625);
or UO_1949 (O_1949,N_12034,N_14681);
or UO_1950 (O_1950,N_12440,N_14430);
and UO_1951 (O_1951,N_12965,N_11976);
or UO_1952 (O_1952,N_14909,N_12932);
nand UO_1953 (O_1953,N_10349,N_12568);
and UO_1954 (O_1954,N_14773,N_11212);
nand UO_1955 (O_1955,N_13831,N_12558);
nor UO_1956 (O_1956,N_12396,N_13939);
nand UO_1957 (O_1957,N_14299,N_14734);
and UO_1958 (O_1958,N_10852,N_10948);
and UO_1959 (O_1959,N_10080,N_10097);
or UO_1960 (O_1960,N_11198,N_11942);
and UO_1961 (O_1961,N_12516,N_13070);
and UO_1962 (O_1962,N_10863,N_11573);
or UO_1963 (O_1963,N_12056,N_12219);
and UO_1964 (O_1964,N_13898,N_12804);
nand UO_1965 (O_1965,N_13499,N_14721);
nor UO_1966 (O_1966,N_10197,N_12207);
and UO_1967 (O_1967,N_10171,N_13985);
nand UO_1968 (O_1968,N_13124,N_14387);
nor UO_1969 (O_1969,N_14627,N_10478);
or UO_1970 (O_1970,N_13074,N_11144);
or UO_1971 (O_1971,N_13949,N_11919);
and UO_1972 (O_1972,N_13421,N_14080);
and UO_1973 (O_1973,N_12812,N_11329);
nand UO_1974 (O_1974,N_10425,N_10587);
nand UO_1975 (O_1975,N_13551,N_13645);
or UO_1976 (O_1976,N_12374,N_11002);
nand UO_1977 (O_1977,N_13087,N_12763);
nand UO_1978 (O_1978,N_11001,N_11868);
nor UO_1979 (O_1979,N_10541,N_10599);
and UO_1980 (O_1980,N_11112,N_12004);
and UO_1981 (O_1981,N_13929,N_13659);
or UO_1982 (O_1982,N_10921,N_11493);
nor UO_1983 (O_1983,N_11290,N_13916);
nor UO_1984 (O_1984,N_12673,N_12143);
nor UO_1985 (O_1985,N_12178,N_14312);
and UO_1986 (O_1986,N_12922,N_12138);
or UO_1987 (O_1987,N_13705,N_10059);
and UO_1988 (O_1988,N_14637,N_12599);
and UO_1989 (O_1989,N_14985,N_14016);
nand UO_1990 (O_1990,N_10296,N_14227);
nand UO_1991 (O_1991,N_11118,N_11486);
or UO_1992 (O_1992,N_10949,N_13008);
xnor UO_1993 (O_1993,N_13661,N_10014);
and UO_1994 (O_1994,N_14764,N_11812);
and UO_1995 (O_1995,N_10414,N_11016);
or UO_1996 (O_1996,N_10198,N_12801);
or UO_1997 (O_1997,N_11428,N_11929);
and UO_1998 (O_1998,N_14580,N_14899);
and UO_1999 (O_1999,N_12273,N_12956);
endmodule