module basic_2500_25000_3000_4_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18883,N_18884,N_18885,N_18886,N_18887,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19032,N_19033,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19103,N_19105,N_19106,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19241,N_19242,N_19243,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19472,N_19473,N_19474,N_19475,N_19476,N_19478,N_19479,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19493,N_19494,N_19495,N_19496,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19912,N_19913,N_19914,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19936,N_19938,N_19939,N_19941,N_19942,N_19943,N_19945,N_19946,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20105,N_20106,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20147,N_20148,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20281,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20304,N_20305,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20341,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20352,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20371,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20635,N_20636,N_20637,N_20638,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20692,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20938,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21153,N_21154,N_21155,N_21156,N_21157,N_21159,N_21160,N_21161,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21203,N_21204,N_21205,N_21206,N_21207,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21367,N_21368,N_21369,N_21370,N_21371,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21620,N_21621,N_21622,N_21623,N_21624,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21771,N_21772,N_21773,N_21774,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22134,N_22135,N_22136,N_22137,N_22138,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22247,N_22248,N_22249,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22512,N_22513,N_22514,N_22515,N_22516,N_22518,N_22519,N_22521,N_22522,N_22523,N_22524,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22549,N_22550,N_22551,N_22552,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22724,N_22725,N_22726,N_22727,N_22728,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22953,N_22954,N_22955,N_22956,N_22957,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23048,N_23049,N_23050,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23413,N_23414,N_23415,N_23416,N_23417,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23631,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23872,N_23873,N_23874,N_23875,N_23876,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23908,N_23909,N_23910,N_23911,N_23912,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24214,N_24215,N_24216,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24293,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24340,N_24341,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24397,N_24398,N_24399,N_24400,N_24401,N_24403,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24452,N_24453,N_24454,N_24455,N_24456,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24491,N_24492,N_24493,N_24494,N_24495,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24567,N_24568,N_24569,N_24570,N_24571,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24600,N_24601,N_24602,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
or U0 (N_0,In_2146,In_638);
xnor U1 (N_1,In_2098,In_230);
xnor U2 (N_2,In_2412,In_2390);
nor U3 (N_3,In_2393,In_1537);
nor U4 (N_4,In_288,In_1736);
nor U5 (N_5,In_2421,In_1487);
nand U6 (N_6,In_300,In_624);
xor U7 (N_7,In_1006,In_1353);
or U8 (N_8,In_2008,In_2044);
and U9 (N_9,In_1044,In_970);
xnor U10 (N_10,In_1381,In_1358);
xnor U11 (N_11,In_2038,In_1627);
nor U12 (N_12,In_2492,In_155);
xnor U13 (N_13,In_485,In_2275);
or U14 (N_14,In_1757,In_2017);
nor U15 (N_15,In_980,In_2201);
nand U16 (N_16,In_2378,In_14);
xor U17 (N_17,In_34,In_109);
nor U18 (N_18,In_2141,In_1216);
xor U19 (N_19,In_771,In_252);
xor U20 (N_20,In_23,In_878);
nand U21 (N_21,In_1441,In_2488);
xor U22 (N_22,In_700,In_661);
xnor U23 (N_23,In_2490,In_956);
and U24 (N_24,In_2135,In_2221);
nand U25 (N_25,In_482,In_1470);
and U26 (N_26,In_398,In_951);
and U27 (N_27,In_1316,In_1984);
nand U28 (N_28,In_1869,In_2065);
or U29 (N_29,In_394,In_90);
xor U30 (N_30,In_1934,In_2450);
or U31 (N_31,In_198,In_815);
nor U32 (N_32,In_646,In_1489);
xor U33 (N_33,In_1564,In_1442);
xor U34 (N_34,In_967,In_1900);
and U35 (N_35,In_32,In_535);
and U36 (N_36,In_206,In_1720);
nand U37 (N_37,In_420,In_526);
xor U38 (N_38,In_1348,In_98);
xnor U39 (N_39,In_1172,In_2013);
xor U40 (N_40,In_1961,In_100);
nand U41 (N_41,In_1229,In_1948);
or U42 (N_42,In_2445,In_345);
or U43 (N_43,In_1037,In_774);
or U44 (N_44,In_701,In_118);
nor U45 (N_45,In_217,In_78);
or U46 (N_46,In_278,In_1086);
nand U47 (N_47,In_812,In_2039);
nand U48 (N_48,In_1885,In_1818);
nor U49 (N_49,In_1262,In_1458);
or U50 (N_50,In_1933,In_2430);
or U51 (N_51,In_1577,In_1892);
nor U52 (N_52,In_2410,In_2010);
nand U53 (N_53,In_455,In_645);
nor U54 (N_54,In_1614,In_1824);
nor U55 (N_55,In_226,In_938);
or U56 (N_56,In_193,In_2079);
nand U57 (N_57,In_2387,In_124);
or U58 (N_58,In_2391,In_1372);
xnor U59 (N_59,In_1499,In_1060);
nor U60 (N_60,In_486,In_857);
and U61 (N_61,In_1950,In_448);
nand U62 (N_62,In_1000,In_96);
nand U63 (N_63,In_196,In_1619);
nand U64 (N_64,In_2369,In_122);
nand U65 (N_65,In_1920,In_881);
and U66 (N_66,In_170,In_2380);
nor U67 (N_67,In_407,In_768);
nand U68 (N_68,In_93,In_619);
nor U69 (N_69,In_213,In_2286);
and U70 (N_70,In_593,In_2491);
or U71 (N_71,In_59,In_1019);
or U72 (N_72,In_322,In_2381);
nor U73 (N_73,In_1500,In_149);
nor U74 (N_74,In_373,In_2164);
nor U75 (N_75,In_549,In_1245);
and U76 (N_76,In_1980,In_1699);
xnor U77 (N_77,In_1547,In_2243);
and U78 (N_78,In_1194,In_130);
and U79 (N_79,In_1586,In_2396);
and U80 (N_80,In_859,In_1280);
nand U81 (N_81,In_2230,In_242);
and U82 (N_82,In_806,In_2249);
and U83 (N_83,In_1707,In_657);
nand U84 (N_84,In_802,In_1007);
nor U85 (N_85,In_357,In_1518);
and U86 (N_86,In_215,In_917);
or U87 (N_87,In_2311,In_1072);
or U88 (N_88,In_1297,In_2261);
or U89 (N_89,In_840,In_1015);
xor U90 (N_90,In_386,In_1616);
nand U91 (N_91,In_2106,In_18);
nand U92 (N_92,In_1403,In_1395);
and U93 (N_93,In_1485,In_319);
or U94 (N_94,In_1105,In_1288);
and U95 (N_95,In_1362,In_957);
and U96 (N_96,In_1452,In_2171);
nor U97 (N_97,In_1163,In_668);
and U98 (N_98,In_1561,In_247);
nand U99 (N_99,In_2365,In_1324);
and U100 (N_100,In_123,In_898);
nor U101 (N_101,In_1842,In_129);
xor U102 (N_102,In_2295,In_1067);
nand U103 (N_103,In_1415,In_1625);
or U104 (N_104,In_2478,In_2138);
and U105 (N_105,In_150,In_1643);
nor U106 (N_106,In_998,In_1726);
or U107 (N_107,In_1445,In_530);
nand U108 (N_108,In_1633,In_2428);
or U109 (N_109,In_566,In_2288);
xor U110 (N_110,In_1122,In_2251);
or U111 (N_111,In_2464,In_1941);
nor U112 (N_112,In_1755,In_1543);
nor U113 (N_113,In_2315,In_2499);
nand U114 (N_114,In_902,In_348);
nand U115 (N_115,In_311,In_2271);
and U116 (N_116,In_105,In_991);
nand U117 (N_117,In_906,In_552);
xor U118 (N_118,In_2375,In_1135);
xor U119 (N_119,In_2257,In_2136);
and U120 (N_120,In_2234,In_2110);
nor U121 (N_121,In_505,In_457);
xnor U122 (N_122,In_2468,In_1253);
and U123 (N_123,In_2133,In_1190);
and U124 (N_124,In_1361,In_1530);
and U125 (N_125,In_297,In_2435);
nand U126 (N_126,In_697,In_1460);
and U127 (N_127,In_2349,In_2006);
nand U128 (N_128,In_2120,In_2258);
nor U129 (N_129,In_167,In_1220);
or U130 (N_130,In_875,In_1123);
xor U131 (N_131,In_1375,In_703);
xor U132 (N_132,In_2190,In_243);
nand U133 (N_133,In_1569,In_2077);
nand U134 (N_134,In_825,In_1205);
or U135 (N_135,In_1888,In_1651);
nor U136 (N_136,In_212,In_396);
nand U137 (N_137,In_2188,In_2183);
xnor U138 (N_138,In_1713,In_112);
xnor U139 (N_139,In_423,In_1531);
xor U140 (N_140,In_1256,In_71);
and U141 (N_141,In_2448,In_251);
nor U142 (N_142,In_1680,In_2075);
xnor U143 (N_143,In_393,In_1812);
nor U144 (N_144,In_1865,In_1769);
nor U145 (N_145,In_1302,In_1159);
or U146 (N_146,In_735,In_419);
and U147 (N_147,In_679,In_2312);
nand U148 (N_148,In_2057,In_2111);
nand U149 (N_149,In_2350,In_846);
and U150 (N_150,In_673,In_576);
and U151 (N_151,In_1807,In_2329);
xor U152 (N_152,In_1343,In_1878);
nor U153 (N_153,In_949,In_1921);
and U154 (N_154,In_1797,In_2404);
and U155 (N_155,In_381,In_2415);
nand U156 (N_156,In_727,In_2336);
nand U157 (N_157,In_450,In_965);
or U158 (N_158,In_598,In_926);
or U159 (N_159,In_1847,In_1609);
and U160 (N_160,In_851,In_1438);
xor U161 (N_161,In_1212,In_959);
or U162 (N_162,In_1925,In_1868);
and U163 (N_163,In_1556,In_1404);
and U164 (N_164,In_1239,In_209);
and U165 (N_165,In_1018,In_1772);
nand U166 (N_166,In_21,In_2025);
nand U167 (N_167,In_563,In_1636);
xnor U168 (N_168,In_1834,In_940);
xnor U169 (N_169,In_1174,In_1965);
and U170 (N_170,In_1638,In_2370);
or U171 (N_171,In_777,In_635);
or U172 (N_172,In_974,In_1191);
nand U173 (N_173,In_1615,In_2262);
nand U174 (N_174,In_1778,In_1486);
xor U175 (N_175,In_1055,In_1221);
or U176 (N_176,In_931,In_1117);
nand U177 (N_177,In_293,In_820);
nor U178 (N_178,In_568,In_211);
nand U179 (N_179,In_2156,In_1150);
nand U180 (N_180,In_308,In_264);
nand U181 (N_181,In_403,In_480);
and U182 (N_182,In_0,In_775);
nand U183 (N_183,In_1606,In_350);
nor U184 (N_184,In_1915,In_41);
nand U185 (N_185,In_428,In_1623);
and U186 (N_186,In_1550,In_1644);
and U187 (N_187,In_192,In_2062);
xnor U188 (N_188,In_2093,In_66);
xor U189 (N_189,In_1581,In_539);
xnor U190 (N_190,In_928,In_1701);
or U191 (N_191,In_341,In_546);
xor U192 (N_192,In_440,In_558);
nor U193 (N_193,In_1990,In_1048);
nand U194 (N_194,In_445,In_498);
nor U195 (N_195,In_501,In_2260);
xnor U196 (N_196,In_3,In_818);
nor U197 (N_197,In_157,In_2245);
xor U198 (N_198,In_483,In_923);
or U199 (N_199,In_2352,In_1168);
and U200 (N_200,In_783,In_767);
and U201 (N_201,In_271,In_2240);
nand U202 (N_202,In_1151,In_2317);
nand U203 (N_203,In_2455,In_1099);
or U204 (N_204,In_1494,In_1815);
nand U205 (N_205,In_559,In_726);
or U206 (N_206,In_2267,In_1466);
and U207 (N_207,In_1991,In_1856);
nand U208 (N_208,In_1794,In_444);
nand U209 (N_209,In_92,In_391);
or U210 (N_210,In_1735,In_1440);
xnor U211 (N_211,In_933,In_347);
and U212 (N_212,In_612,In_402);
or U213 (N_213,In_1679,In_352);
nand U214 (N_214,In_146,In_459);
nand U215 (N_215,In_2265,In_338);
xor U216 (N_216,In_382,In_979);
xnor U217 (N_217,In_1337,In_1066);
nor U218 (N_218,In_1383,In_695);
and U219 (N_219,In_588,In_314);
and U220 (N_220,In_2224,In_2047);
and U221 (N_221,In_801,In_1836);
or U222 (N_222,In_2268,In_312);
nor U223 (N_223,In_2328,In_94);
nand U224 (N_224,In_2151,In_354);
or U225 (N_225,In_323,In_1250);
or U226 (N_226,In_1765,In_169);
and U227 (N_227,In_704,In_686);
or U228 (N_228,In_2345,In_597);
nor U229 (N_229,In_143,In_1109);
xor U230 (N_230,In_874,In_596);
or U231 (N_231,In_97,In_379);
nand U232 (N_232,In_2117,In_1088);
nor U233 (N_233,In_1901,In_2229);
nand U234 (N_234,In_664,In_1821);
nand U235 (N_235,In_2419,In_833);
and U236 (N_236,In_222,In_1913);
xnor U237 (N_237,In_538,In_1234);
or U238 (N_238,In_1505,In_2073);
and U239 (N_239,In_758,In_1761);
and U240 (N_240,In_698,In_1396);
or U241 (N_241,In_1671,In_1424);
xor U242 (N_242,In_1905,In_1448);
or U243 (N_243,In_454,In_1808);
and U244 (N_244,In_748,In_1800);
nor U245 (N_245,In_2424,In_1594);
nor U246 (N_246,In_375,In_1937);
or U247 (N_247,In_1180,In_1331);
or U248 (N_248,In_134,In_2332);
xor U249 (N_249,In_153,In_2359);
xor U250 (N_250,In_1228,In_893);
xnor U251 (N_251,In_863,In_299);
nand U252 (N_252,In_2300,In_1685);
nand U253 (N_253,In_1003,In_1598);
xnor U254 (N_254,In_218,In_2443);
or U255 (N_255,In_2320,In_1585);
and U256 (N_256,In_358,In_102);
or U257 (N_257,In_1804,In_1977);
nor U258 (N_258,In_1226,In_852);
and U259 (N_259,In_632,In_88);
or U260 (N_260,In_603,In_68);
and U261 (N_261,In_1779,In_1389);
nand U262 (N_262,In_33,In_834);
xnor U263 (N_263,In_2423,In_426);
and U264 (N_264,In_1575,In_1282);
or U265 (N_265,In_1972,In_2154);
or U266 (N_266,In_1070,In_1249);
xor U267 (N_267,In_1944,In_2326);
or U268 (N_268,In_674,In_1512);
xor U269 (N_269,In_1597,In_858);
and U270 (N_270,In_2383,In_714);
xnor U271 (N_271,In_2322,In_276);
and U272 (N_272,In_2399,In_1176);
nor U273 (N_273,In_2347,In_565);
nand U274 (N_274,In_1277,In_1144);
and U275 (N_275,In_2395,In_821);
xor U276 (N_276,In_1673,In_751);
nor U277 (N_277,In_717,In_1468);
and U278 (N_278,In_995,In_1371);
nand U279 (N_279,In_1162,In_1380);
or U280 (N_280,In_569,In_660);
and U281 (N_281,In_1539,In_2078);
and U282 (N_282,In_1542,In_2167);
nand U283 (N_283,In_2088,In_378);
nand U284 (N_284,In_219,In_1241);
xor U285 (N_285,In_912,In_1121);
nand U286 (N_286,In_377,In_1813);
xor U287 (N_287,In_656,In_1570);
and U288 (N_288,In_461,In_861);
xor U289 (N_289,In_2179,In_1873);
nor U290 (N_290,In_1654,In_2244);
or U291 (N_291,In_282,In_1902);
nand U292 (N_292,In_1085,In_2163);
nand U293 (N_293,In_1391,In_1126);
nor U294 (N_294,In_1491,In_966);
nand U295 (N_295,In_2247,In_1106);
and U296 (N_296,In_2192,In_1098);
or U297 (N_297,In_262,In_1566);
nor U298 (N_298,In_1762,In_1611);
nor U299 (N_299,In_2114,In_329);
or U300 (N_300,In_1766,In_1);
nand U301 (N_301,In_2469,In_127);
or U302 (N_302,In_895,In_1456);
or U303 (N_303,In_315,In_1823);
nor U304 (N_304,In_1718,In_927);
and U305 (N_305,In_356,In_2398);
xnor U306 (N_306,In_1447,In_647);
and U307 (N_307,In_1140,In_1014);
nor U308 (N_308,In_361,In_1173);
nand U309 (N_309,In_2087,In_2427);
or U310 (N_310,In_1822,In_185);
or U311 (N_311,In_533,In_2474);
and U312 (N_312,In_332,In_1536);
nand U313 (N_313,In_1269,In_214);
and U314 (N_314,In_1666,In_616);
nor U315 (N_315,In_788,In_793);
nand U316 (N_316,In_633,In_829);
xor U317 (N_317,In_1789,In_1509);
xor U318 (N_318,In_1112,In_1613);
xnor U319 (N_319,In_1087,In_947);
and U320 (N_320,In_231,In_2382);
and U321 (N_321,In_1867,In_866);
nand U322 (N_322,In_1744,In_2220);
and U323 (N_323,In_798,In_1439);
or U324 (N_324,In_1405,In_1672);
nand U325 (N_325,In_2132,In_914);
or U326 (N_326,In_1764,In_1544);
or U327 (N_327,In_813,In_1454);
nor U328 (N_328,In_888,In_696);
nand U329 (N_329,In_2162,In_1023);
and U330 (N_330,In_578,In_710);
nand U331 (N_331,In_383,In_1053);
and U332 (N_332,In_1747,In_805);
xnor U333 (N_333,In_1785,In_823);
xor U334 (N_334,In_1783,In_236);
or U335 (N_335,In_1711,In_665);
nand U336 (N_336,In_191,In_982);
and U337 (N_337,In_1540,In_2290);
xor U338 (N_338,In_1266,In_760);
or U339 (N_339,In_745,In_1700);
nand U340 (N_340,In_891,In_1605);
nor U341 (N_341,In_1376,In_1310);
xnor U342 (N_342,In_1394,In_611);
nand U343 (N_343,In_470,In_766);
xnor U344 (N_344,In_1929,In_958);
or U345 (N_345,In_631,In_1198);
and U346 (N_346,In_283,In_17);
or U347 (N_347,In_1094,In_2401);
xor U348 (N_348,In_1278,In_2123);
nand U349 (N_349,In_2457,In_1706);
nor U350 (N_350,In_26,In_853);
xor U351 (N_351,In_1942,In_2321);
xor U352 (N_352,In_25,In_2494);
or U353 (N_353,In_1155,In_437);
nor U354 (N_354,In_1659,In_2134);
and U355 (N_355,In_1422,In_2496);
nand U356 (N_356,In_73,In_1091);
or U357 (N_357,In_1386,In_595);
or U358 (N_358,In_113,In_1252);
and U359 (N_359,In_1457,In_1165);
or U360 (N_360,In_1774,In_1628);
or U361 (N_361,In_2480,In_487);
nand U362 (N_362,In_1898,In_2296);
nand U363 (N_363,In_2035,In_363);
nor U364 (N_364,In_415,In_2465);
xnor U365 (N_365,In_1683,In_1805);
or U366 (N_366,In_1525,In_1336);
and U367 (N_367,In_2071,In_1263);
xnor U368 (N_368,In_261,In_2191);
nor U369 (N_369,In_1062,In_1914);
xor U370 (N_370,In_884,In_2068);
nand U371 (N_371,In_2231,In_1399);
and U372 (N_372,In_1368,In_628);
xnor U373 (N_373,In_16,In_582);
and U374 (N_374,In_1129,In_892);
and U375 (N_375,In_1634,In_762);
nor U376 (N_376,In_2341,In_1884);
xnor U377 (N_377,In_210,In_909);
xnor U378 (N_378,In_1420,In_179);
nor U379 (N_379,In_605,In_2318);
xor U380 (N_380,In_2413,In_2446);
or U381 (N_381,In_1662,In_746);
nor U382 (N_382,In_2096,In_2099);
nand U383 (N_383,In_1649,In_843);
xnor U384 (N_384,In_2218,In_65);
nand U385 (N_385,In_1255,In_870);
nand U386 (N_386,In_776,In_1039);
nor U387 (N_387,In_610,In_1244);
nor U388 (N_388,In_1891,In_592);
xnor U389 (N_389,In_61,In_1164);
or U390 (N_390,In_1945,In_241);
and U391 (N_391,In_2314,In_1258);
and U392 (N_392,In_413,In_625);
or U393 (N_393,In_2449,In_2129);
and U394 (N_394,In_2386,In_886);
or U395 (N_395,In_1493,In_1741);
nor U396 (N_396,In_2287,In_1203);
xnor U397 (N_397,In_2487,In_2305);
xor U398 (N_398,In_1831,In_1477);
or U399 (N_399,In_2211,In_2225);
nor U400 (N_400,In_1142,In_687);
nor U401 (N_401,In_1705,In_2086);
nand U402 (N_402,In_2361,In_2473);
or U403 (N_403,In_2041,In_1935);
and U404 (N_404,In_1599,In_2178);
xnor U405 (N_405,In_694,In_1689);
or U406 (N_406,In_2127,In_1011);
and U407 (N_407,In_2301,In_1450);
nor U408 (N_408,In_1854,In_81);
and U409 (N_409,In_741,In_266);
nor U410 (N_410,In_997,In_234);
nor U411 (N_411,In_666,In_1926);
xnor U412 (N_412,In_856,In_1274);
xor U413 (N_413,In_1461,In_284);
nor U414 (N_414,In_56,In_331);
xor U415 (N_415,In_2475,In_216);
and U416 (N_416,In_877,In_371);
nand U417 (N_417,In_955,In_1588);
nand U418 (N_418,In_1517,In_1732);
or U419 (N_419,In_640,In_369);
xor U420 (N_420,In_2187,In_2357);
nand U421 (N_421,In_1286,In_1046);
and U422 (N_422,In_1809,In_543);
nand U423 (N_423,In_87,In_879);
and U424 (N_424,In_1025,In_709);
xnor U425 (N_425,In_901,In_882);
or U426 (N_426,In_934,In_1043);
and U427 (N_427,In_1077,In_1835);
or U428 (N_428,In_1279,In_2344);
or U429 (N_429,In_1896,In_2107);
nor U430 (N_430,In_328,In_964);
nor U431 (N_431,In_490,In_2012);
nor U432 (N_432,In_835,In_1031);
nand U433 (N_433,In_2219,In_988);
and U434 (N_434,In_2108,In_2097);
nand U435 (N_435,In_63,In_2397);
xnor U436 (N_436,In_2203,In_194);
nand U437 (N_437,In_1918,In_721);
or U438 (N_438,In_1572,In_1607);
nor U439 (N_439,In_2054,In_2340);
xnor U440 (N_440,In_1960,In_1786);
and U441 (N_441,In_2254,In_606);
xnor U442 (N_442,In_1602,In_1322);
nor U443 (N_443,In_2403,In_1412);
nor U444 (N_444,In_2283,In_446);
and U445 (N_445,In_1907,In_492);
and U446 (N_446,In_2130,In_1125);
or U447 (N_447,In_95,In_529);
nand U448 (N_448,In_1748,In_683);
xor U449 (N_449,In_156,In_838);
or U450 (N_450,In_36,In_1579);
nand U451 (N_451,In_313,In_2333);
and U452 (N_452,In_1318,In_1811);
and U453 (N_453,In_165,In_1475);
or U454 (N_454,In_983,In_702);
and U455 (N_455,In_1474,In_681);
or U456 (N_456,In_1083,In_1411);
and U457 (N_457,In_691,In_1521);
nand U458 (N_458,In_1733,In_2463);
nor U459 (N_459,In_1344,In_1759);
nand U460 (N_460,In_35,In_430);
nand U461 (N_461,In_132,In_1170);
nand U462 (N_462,In_1894,In_1848);
or U463 (N_463,In_280,In_1708);
nand U464 (N_464,In_1365,In_1946);
xor U465 (N_465,In_1149,In_725);
xnor U466 (N_466,In_567,In_1305);
and U467 (N_467,In_2368,In_525);
xnor U468 (N_468,In_2092,In_921);
nand U469 (N_469,In_722,In_1116);
and U470 (N_470,In_15,In_1975);
xnor U471 (N_471,In_1480,In_1035);
xor U472 (N_472,In_2418,In_2155);
xor U473 (N_473,In_924,In_1058);
or U474 (N_474,In_1970,In_2128);
or U475 (N_475,In_2072,In_309);
xnor U476 (N_476,In_855,In_519);
xnor U477 (N_477,In_1090,In_1791);
xor U478 (N_478,In_359,In_1511);
xor U479 (N_479,In_1538,In_1136);
and U480 (N_480,In_1535,In_1879);
xor U481 (N_481,In_2207,In_2238);
nand U482 (N_482,In_749,In_1985);
xor U483 (N_483,In_981,In_521);
nand U484 (N_484,In_589,In_978);
nor U485 (N_485,In_2009,In_765);
and U486 (N_486,In_1496,In_1604);
nand U487 (N_487,In_976,In_2023);
xnor U488 (N_488,In_2113,In_2067);
and U489 (N_489,In_1632,In_600);
and U490 (N_490,In_239,In_899);
or U491 (N_491,In_667,In_1739);
or U492 (N_492,In_996,In_992);
xnor U493 (N_493,In_946,In_142);
and U494 (N_494,In_307,In_1179);
xor U495 (N_495,In_1027,In_1382);
xor U496 (N_496,In_699,In_335);
and U497 (N_497,In_800,In_1068);
nor U498 (N_498,In_101,In_2241);
xnor U499 (N_499,In_677,In_1479);
nor U500 (N_500,In_1690,In_1178);
or U501 (N_501,In_1005,In_2353);
nand U502 (N_502,In_2331,In_4);
nor U503 (N_503,In_189,In_2157);
nor U504 (N_504,In_507,In_1810);
xor U505 (N_505,In_1233,In_913);
nand U506 (N_506,In_249,In_2213);
or U507 (N_507,In_466,In_1858);
xnor U508 (N_508,In_761,In_1026);
or U509 (N_509,In_12,In_1908);
nand U510 (N_510,In_658,In_1209);
xnor U511 (N_511,In_1940,In_560);
or U512 (N_512,In_2158,In_1160);
xnor U513 (N_513,In_1268,In_684);
or U514 (N_514,In_1276,In_1698);
xor U515 (N_515,In_1265,In_832);
or U516 (N_516,In_680,In_786);
or U517 (N_517,In_1267,In_42);
xor U518 (N_518,In_575,In_237);
nor U519 (N_519,In_465,In_2307);
nor U520 (N_520,In_1045,In_494);
nor U521 (N_521,In_2441,In_401);
and U522 (N_522,In_1377,In_1731);
xnor U523 (N_523,In_1428,In_2034);
xor U524 (N_524,In_1443,In_839);
or U525 (N_525,In_876,In_108);
nor U526 (N_526,In_75,In_1912);
nor U527 (N_527,In_463,In_2454);
nand U528 (N_528,In_1319,In_1294);
nor U529 (N_529,In_1421,In_462);
xnor U530 (N_530,In_1557,In_2066);
xnor U531 (N_531,In_1398,In_2440);
and U532 (N_532,In_1702,In_1568);
xnor U533 (N_533,In_2055,In_1334);
xor U534 (N_534,In_1860,In_993);
nor U535 (N_535,In_1110,In_48);
nor U536 (N_536,In_864,In_1646);
nand U537 (N_537,In_2103,In_1639);
and U538 (N_538,In_962,In_2497);
and U539 (N_539,In_493,In_431);
nand U540 (N_540,In_57,In_298);
or U541 (N_541,In_1749,In_670);
xnor U542 (N_542,In_1819,In_1855);
or U543 (N_543,In_1427,In_2002);
nand U544 (N_544,In_1040,In_2040);
nor U545 (N_545,In_1119,In_1603);
xnor U546 (N_546,In_1534,In_1021);
and U547 (N_547,In_1760,In_2367);
nand U548 (N_548,In_523,In_104);
or U549 (N_549,In_1520,In_570);
xor U550 (N_550,In_2362,In_1979);
and U551 (N_551,In_2313,In_238);
or U552 (N_552,In_1838,In_1664);
xnor U553 (N_553,In_2202,In_1281);
and U554 (N_554,In_52,In_2235);
nor U555 (N_555,In_1145,In_182);
nand U556 (N_556,In_2027,In_2292);
nand U557 (N_557,In_1754,In_1532);
or U558 (N_558,In_508,In_1924);
nand U559 (N_559,In_2263,In_67);
nor U560 (N_560,In_764,In_1473);
and U561 (N_561,In_827,In_7);
or U562 (N_562,In_432,In_294);
and U563 (N_563,In_400,In_1938);
xor U564 (N_564,In_414,In_269);
nor U565 (N_565,In_1153,In_807);
xor U566 (N_566,In_890,In_1097);
or U567 (N_567,In_19,In_1200);
and U568 (N_568,In_724,In_2181);
and U569 (N_569,In_1595,In_2118);
or U570 (N_570,In_433,In_439);
and U571 (N_571,In_1307,In_803);
or U572 (N_572,In_141,In_860);
nor U573 (N_573,In_2121,In_1184);
or U574 (N_574,In_1552,In_1682);
and U575 (N_575,In_2411,In_693);
nand U576 (N_576,In_2015,In_2425);
nor U577 (N_577,In_2364,In_794);
xnor U578 (N_578,In_1224,In_1910);
nor U579 (N_579,In_1844,In_1657);
or U580 (N_580,In_362,In_2289);
xor U581 (N_581,In_2070,In_828);
nand U582 (N_582,In_609,In_705);
xnor U583 (N_583,In_2436,In_232);
nor U584 (N_584,In_763,In_1752);
or U585 (N_585,In_471,In_1571);
nor U586 (N_586,In_139,In_908);
and U587 (N_587,In_1799,In_1236);
nor U588 (N_588,In_1642,In_1357);
or U589 (N_589,In_541,In_1326);
and U590 (N_590,In_1061,In_644);
nand U591 (N_591,In_1546,In_708);
or U592 (N_592,In_1272,In_1751);
or U593 (N_593,In_1936,In_1750);
or U594 (N_594,In_1877,In_1009);
nor U595 (N_595,In_1141,In_2405);
nor U596 (N_596,In_642,In_954);
nor U597 (N_597,In_2147,In_1528);
and U598 (N_598,In_757,In_1188);
and U599 (N_599,In_2385,In_2105);
nor U600 (N_600,In_1904,In_1994);
and U601 (N_601,In_2302,In_2316);
xor U602 (N_602,In_1373,In_2082);
xnor U603 (N_603,In_110,In_738);
nor U604 (N_604,In_1788,In_2193);
and U605 (N_605,In_1222,In_581);
xnor U606 (N_606,In_637,In_1770);
or U607 (N_607,In_1966,In_2479);
xnor U608 (N_608,In_2186,In_527);
and U609 (N_609,In_528,In_2447);
nor U610 (N_610,In_79,In_1010);
xor U611 (N_611,In_343,In_443);
xor U612 (N_612,In_1522,In_1541);
and U613 (N_613,In_810,In_1299);
nor U614 (N_614,In_1529,In_1364);
nand U615 (N_615,In_1618,In_973);
nand U616 (N_616,In_791,In_587);
xor U617 (N_617,In_1971,In_190);
nand U618 (N_618,In_119,In_1533);
and U619 (N_619,In_557,In_275);
and U620 (N_620,In_1650,In_1432);
and U621 (N_621,In_49,In_2074);
or U622 (N_622,In_968,In_1782);
xnor U623 (N_623,In_259,In_836);
nand U624 (N_624,In_116,In_1453);
or U625 (N_625,In_1560,In_518);
nand U626 (N_626,In_235,In_2028);
nand U627 (N_627,In_1196,In_2217);
and U628 (N_628,In_1124,In_942);
xnor U629 (N_629,In_1296,In_1455);
nand U630 (N_630,In_1075,In_2180);
xor U631 (N_631,In_1880,In_1465);
xor U632 (N_632,In_349,In_2481);
xor U633 (N_633,In_1631,In_1724);
nor U634 (N_634,In_2061,In_2145);
xnor U635 (N_635,In_317,In_573);
and U636 (N_636,In_346,In_1137);
xor U637 (N_637,In_1192,In_1670);
nor U638 (N_638,In_1211,In_1676);
nor U639 (N_639,In_86,In_1128);
and U640 (N_640,In_1346,In_2053);
nand U641 (N_641,In_187,In_2366);
nor U642 (N_642,In_2392,In_706);
nor U643 (N_643,In_1092,In_1899);
xor U644 (N_644,In_91,In_1347);
or U645 (N_645,In_1207,In_1030);
xor U646 (N_646,In_404,In_2298);
or U647 (N_647,In_145,In_1059);
or U648 (N_648,In_1600,In_295);
and U649 (N_649,In_1050,In_1327);
nor U650 (N_650,In_1519,In_1490);
or U651 (N_651,In_344,In_520);
or U652 (N_652,In_385,In_421);
and U653 (N_653,In_2477,In_137);
nor U654 (N_654,In_1622,In_254);
nor U655 (N_655,In_2222,In_1660);
nor U656 (N_656,In_2407,In_310);
nor U657 (N_657,In_630,In_225);
and U658 (N_658,In_952,In_1317);
and U659 (N_659,In_1729,In_1710);
or U660 (N_660,In_614,In_824);
or U661 (N_661,In_1413,In_685);
and U662 (N_662,In_248,In_2204);
xnor U663 (N_663,In_1674,In_2299);
nor U664 (N_664,In_999,In_1974);
nor U665 (N_665,In_496,In_1082);
and U666 (N_666,In_1507,In_532);
xor U667 (N_667,In_903,In_1290);
nor U668 (N_668,In_773,In_2310);
and U669 (N_669,In_1523,In_574);
nor U670 (N_670,In_1177,In_2050);
or U671 (N_671,In_713,In_910);
and U672 (N_672,In_1459,In_2471);
xnor U673 (N_673,In_1251,In_326);
nand U674 (N_674,In_1503,In_1687);
nand U675 (N_675,In_2356,In_469);
nor U676 (N_676,In_1516,In_1897);
xor U677 (N_677,In_918,In_636);
or U678 (N_678,In_781,In_939);
nand U679 (N_679,In_2306,In_731);
nand U680 (N_680,In_1064,In_617);
or U681 (N_681,In_1978,In_1032);
or U682 (N_682,In_1147,In_1369);
and U683 (N_683,In_1218,In_641);
or U684 (N_684,In_453,In_1437);
xnor U685 (N_685,In_1330,In_1758);
or U686 (N_686,In_1020,In_2426);
nand U687 (N_687,In_663,In_2032);
or U688 (N_688,In_1333,In_868);
and U689 (N_689,In_1968,In_174);
xnor U690 (N_690,In_2052,In_422);
nor U691 (N_691,In_1957,In_204);
nor U692 (N_692,In_31,In_1514);
xnor U693 (N_693,In_2456,In_1781);
nor U694 (N_694,In_907,In_1645);
and U695 (N_695,In_841,In_106);
and U696 (N_696,In_481,In_896);
nor U697 (N_697,In_1118,In_2277);
xnor U698 (N_698,In_2173,In_114);
or U699 (N_699,In_365,In_2294);
nor U700 (N_700,In_1089,In_905);
nand U701 (N_701,In_1423,In_590);
nor U702 (N_702,In_692,In_1235);
and U703 (N_703,In_1551,In_467);
or U704 (N_704,In_302,In_553);
nand U705 (N_705,In_1678,In_2021);
nor U706 (N_706,In_289,In_1193);
nor U707 (N_707,In_1621,In_2131);
nand U708 (N_708,In_1080,In_1833);
nand U709 (N_709,In_904,In_1029);
or U710 (N_710,In_449,In_1753);
nand U711 (N_711,In_1355,In_2215);
and U712 (N_712,In_1969,In_1104);
xnor U713 (N_713,In_1467,In_1951);
and U714 (N_714,In_1237,In_417);
nand U715 (N_715,In_2432,In_1261);
or U716 (N_716,In_2014,In_51);
and U717 (N_717,In_1034,In_1962);
and U718 (N_718,In_1492,In_883);
nand U719 (N_719,In_1352,In_941);
xor U720 (N_720,In_1583,In_2374);
or U721 (N_721,In_1304,In_2274);
or U722 (N_722,In_221,In_1275);
xnor U723 (N_723,In_975,In_577);
nor U724 (N_724,In_39,In_399);
nand U725 (N_725,In_1495,In_2102);
xnor U726 (N_726,In_943,In_1555);
xnor U727 (N_727,In_1861,In_1215);
and U728 (N_728,In_1806,In_1054);
and U729 (N_729,In_390,In_2308);
and U730 (N_730,In_1911,In_564);
nand U731 (N_731,In_1400,In_1360);
nand U732 (N_732,In_515,In_1576);
nand U733 (N_733,In_85,In_1895);
nor U734 (N_734,In_2206,In_2309);
xnor U735 (N_735,In_1004,In_862);
and U736 (N_736,In_2085,In_2182);
nand U737 (N_737,In_1704,In_916);
or U738 (N_738,In_1987,In_897);
xor U739 (N_739,In_2269,In_408);
or U740 (N_740,In_930,In_1169);
xnor U741 (N_741,In_1675,In_2384);
or U742 (N_742,In_1102,In_796);
nor U743 (N_743,In_2007,In_627);
or U744 (N_744,In_2051,In_1506);
nor U745 (N_745,In_623,In_1242);
xor U746 (N_746,In_1875,In_2429);
nor U747 (N_747,In_1964,In_822);
nor U748 (N_748,In_608,In_244);
and U749 (N_749,In_1709,In_2414);
xor U750 (N_750,In_971,In_2081);
nand U751 (N_751,In_171,In_1407);
nor U752 (N_752,In_2323,In_126);
xor U753 (N_753,In_2233,In_255);
and U754 (N_754,In_1798,In_1589);
xnor U755 (N_755,In_2153,In_1033);
xnor U756 (N_756,In_2214,In_45);
and U757 (N_757,In_2272,In_919);
nand U758 (N_758,In_1139,In_1728);
nor U759 (N_759,In_120,In_2291);
and U760 (N_760,In_1610,In_1309);
xor U761 (N_761,In_945,In_1953);
and U762 (N_762,In_2094,In_258);
nand U763 (N_763,In_562,In_1189);
nand U764 (N_764,In_545,In_342);
xnor U765 (N_765,In_994,In_1202);
or U766 (N_766,In_756,In_2355);
xor U767 (N_767,In_555,In_534);
and U768 (N_768,In_316,In_2459);
or U769 (N_769,In_474,In_138);
and U770 (N_770,In_1850,In_1183);
nand U771 (N_771,In_183,In_613);
nor U772 (N_772,In_2438,In_1038);
or U773 (N_773,In_250,In_1338);
nand U774 (N_774,In_55,In_1996);
and U775 (N_775,In_672,In_2461);
xnor U776 (N_776,In_1841,In_730);
nor U777 (N_777,In_1740,In_2408);
nand U778 (N_778,In_911,In_131);
xnor U779 (N_779,In_2377,In_1832);
xor U780 (N_780,In_1982,In_488);
or U781 (N_781,In_47,In_787);
nor U782 (N_782,In_1157,In_2325);
nand U783 (N_783,In_889,In_53);
xnor U784 (N_784,In_1199,In_599);
nand U785 (N_785,In_1008,In_1356);
and U786 (N_786,In_1429,In_296);
and U787 (N_787,In_2409,In_2101);
xnor U788 (N_788,In_1526,In_339);
nand U789 (N_789,In_1872,In_84);
xor U790 (N_790,In_1730,In_948);
nand U791 (N_791,In_1719,In_715);
and U792 (N_792,In_1321,In_1243);
xor U793 (N_793,In_2248,In_1069);
nor U794 (N_794,In_1792,In_1775);
nand U795 (N_795,In_1667,In_1208);
nand U796 (N_796,In_531,In_1665);
nand U797 (N_797,In_1093,In_1545);
and U798 (N_798,In_584,In_816);
nand U799 (N_799,In_2170,In_1016);
xnor U800 (N_800,In_2137,In_944);
or U801 (N_801,In_22,In_1283);
and U802 (N_802,In_2372,In_1156);
nor U803 (N_803,In_2029,In_144);
xor U804 (N_804,In_2184,In_1851);
nand U805 (N_805,In_152,In_1451);
and U806 (N_806,In_406,In_1989);
and U807 (N_807,In_188,In_1132);
nand U808 (N_808,In_1481,In_1745);
xor U809 (N_809,In_223,In_1515);
nand U810 (N_810,In_460,In_2281);
or U811 (N_811,In_2116,In_5);
nor U812 (N_812,In_1182,In_1909);
or U813 (N_813,In_671,In_50);
or U814 (N_814,In_1852,In_1484);
and U815 (N_815,In_1303,In_2);
nor U816 (N_816,In_1051,In_1954);
and U817 (N_817,In_1214,In_2165);
xnor U818 (N_818,In_1691,In_1469);
nand U819 (N_819,In_2037,In_1133);
and U820 (N_820,In_2388,In_1311);
nor U821 (N_821,In_580,In_291);
nand U822 (N_822,In_166,In_1247);
or U823 (N_823,In_953,In_1363);
nand U824 (N_824,In_848,In_220);
nand U825 (N_825,In_778,In_384);
and U826 (N_826,In_780,In_960);
nand U827 (N_827,In_1414,In_797);
or U828 (N_828,In_452,In_1367);
xor U829 (N_829,In_497,In_353);
nor U830 (N_830,In_1697,In_438);
nand U831 (N_831,In_814,In_629);
and U832 (N_832,In_2223,In_1341);
xnor U833 (N_833,In_2185,In_887);
or U834 (N_834,In_1186,In_2200);
nand U835 (N_835,In_1187,In_178);
nand U836 (N_836,In_1776,In_1108);
nand U837 (N_837,In_1686,In_2379);
nor U838 (N_838,In_2402,In_1881);
and U839 (N_839,In_2482,In_1669);
xor U840 (N_840,In_2467,In_159);
xnor U841 (N_841,In_925,In_2036);
nand U842 (N_842,In_1308,In_651);
nor U843 (N_843,In_405,In_1287);
or U844 (N_844,In_46,In_2140);
or U845 (N_845,In_733,In_1152);
xnor U846 (N_846,In_477,In_1114);
and U847 (N_847,In_1839,In_643);
and U848 (N_848,In_233,In_1359);
or U849 (N_849,In_1185,In_172);
nand U850 (N_850,In_854,In_1175);
and U851 (N_851,In_318,In_1997);
xnor U852 (N_852,In_1387,In_473);
nor U853 (N_853,In_894,In_2330);
xor U854 (N_854,In_561,In_2161);
nor U855 (N_855,In_826,In_475);
nor U856 (N_856,In_789,In_2453);
xor U857 (N_857,In_1870,In_2084);
xor U858 (N_858,In_1559,In_754);
nor U859 (N_859,In_28,In_1134);
nand U860 (N_860,In_591,In_542);
nand U861 (N_861,In_689,In_1065);
nand U862 (N_862,In_1342,In_1462);
xnor U863 (N_863,In_2216,In_1397);
xor U864 (N_864,In_799,In_1264);
nand U865 (N_865,In_186,In_412);
and U866 (N_866,In_1976,In_1553);
nand U867 (N_867,In_2159,In_1693);
xnor U868 (N_868,In_69,In_871);
nor U869 (N_869,In_265,In_60);
nand U870 (N_870,In_2486,In_1204);
or U871 (N_871,In_76,In_1148);
nor U872 (N_872,In_1408,In_1626);
nor U873 (N_873,In_1167,In_425);
and U874 (N_874,In_1620,In_2003);
nand U875 (N_875,In_1714,In_1927);
nor U876 (N_876,In_655,In_1074);
nor U877 (N_877,In_544,In_2060);
nor U878 (N_878,In_1231,In_2285);
nand U879 (N_879,In_484,In_2334);
and U880 (N_880,In_1640,In_2125);
nand U881 (N_881,In_1435,In_1416);
or U882 (N_882,In_747,In_935);
or U883 (N_883,In_1254,In_1889);
or U884 (N_884,In_1928,In_2342);
and U885 (N_885,In_1743,In_1939);
and U886 (N_886,In_1350,In_550);
nand U887 (N_887,In_932,In_162);
nand U888 (N_888,In_2212,In_301);
and U889 (N_889,In_1629,In_972);
xor U890 (N_890,In_1574,In_662);
nand U891 (N_891,In_817,In_1508);
xnor U892 (N_892,In_2360,In_447);
and U893 (N_893,In_2466,In_2444);
xnor U894 (N_894,In_1981,In_1593);
nor U895 (N_895,In_2227,In_2174);
xnor U896 (N_896,In_117,In_1763);
or U897 (N_897,In_729,In_6);
nand U898 (N_898,In_1887,In_1238);
and U899 (N_899,In_334,In_1213);
xnor U900 (N_900,In_2139,In_1883);
or U901 (N_901,In_125,In_1430);
nand U902 (N_902,In_202,In_2437);
nor U903 (N_903,In_240,In_1201);
and U904 (N_904,In_1314,In_2458);
and U905 (N_905,In_937,In_1052);
xnor U906 (N_906,In_1871,In_1291);
or U907 (N_907,In_873,In_1930);
and U908 (N_908,In_2371,In_2337);
nor U909 (N_909,In_1608,In_324);
xor U910 (N_910,In_1715,In_849);
and U911 (N_911,In_1246,In_389);
nand U912 (N_912,In_847,In_652);
or U913 (N_913,In_2439,In_2276);
nand U914 (N_914,In_963,In_495);
and U915 (N_915,In_1738,In_1079);
or U916 (N_916,In_1573,In_1784);
and U917 (N_917,In_1315,In_1830);
nor U918 (N_918,In_451,In_367);
or U919 (N_919,In_1482,In_984);
nand U920 (N_920,In_2452,In_522);
xnor U921 (N_921,In_175,In_1476);
or U922 (N_922,In_2175,In_1345);
and U923 (N_923,In_1295,In_554);
and U924 (N_924,In_1210,In_1384);
and U925 (N_925,In_2104,In_977);
nor U926 (N_926,In_1859,In_2246);
nor U927 (N_927,In_579,In_410);
nand U928 (N_928,In_245,In_1993);
nor U929 (N_929,In_615,In_424);
nor U930 (N_930,In_759,In_2476);
nor U931 (N_931,In_173,In_304);
and U932 (N_932,In_207,In_1115);
and U933 (N_933,In_479,In_1527);
xor U934 (N_934,In_121,In_2279);
xor U935 (N_935,In_1712,In_1260);
nor U936 (N_936,In_1095,In_989);
nor U937 (N_937,In_2080,In_654);
or U938 (N_938,In_990,In_458);
nor U939 (N_939,In_1433,In_2030);
and U940 (N_940,In_325,In_2063);
nor U941 (N_941,In_2327,In_2210);
nand U942 (N_942,In_1154,In_1692);
xor U943 (N_943,In_1773,In_24);
nor U944 (N_944,In_1992,In_2033);
and U945 (N_945,In_2284,In_70);
and U946 (N_946,In_1312,In_830);
and U947 (N_947,In_1410,In_1617);
or U948 (N_948,In_1013,In_506);
and U949 (N_949,In_1036,In_622);
nor U950 (N_950,In_1906,In_333);
xnor U951 (N_951,In_180,In_1012);
nor U952 (N_952,In_2049,In_1328);
xnor U953 (N_953,In_1298,In_1285);
xor U954 (N_954,In_712,In_1825);
or U955 (N_955,In_737,In_2339);
nor U956 (N_956,In_1668,In_513);
nand U957 (N_957,In_37,In_1017);
or U958 (N_958,In_1259,In_1502);
nor U959 (N_959,In_1524,In_2297);
nor U960 (N_960,In_845,In_1232);
and U961 (N_961,In_1329,In_2460);
and U962 (N_962,In_2019,In_1001);
and U963 (N_963,In_1721,In_1803);
nor U964 (N_964,In_1426,In_360);
nor U965 (N_965,In_2149,In_1041);
and U966 (N_966,In_1677,In_1999);
and U967 (N_967,In_1171,In_1446);
and U968 (N_968,In_1513,In_2177);
nand U969 (N_969,In_517,In_1379);
nand U970 (N_970,In_2226,In_1684);
or U971 (N_971,In_585,In_2400);
and U972 (N_972,In_1846,In_742);
nor U973 (N_973,In_2208,In_639);
and U974 (N_974,In_536,In_181);
xor U975 (N_975,In_551,In_2018);
xor U976 (N_976,In_2169,In_1890);
xnor U977 (N_977,In_290,In_772);
xor U978 (N_978,In_2270,In_1084);
xor U979 (N_979,In_2250,In_1876);
nand U980 (N_980,In_1717,In_2280);
xnor U981 (N_981,In_1002,In_602);
or U982 (N_982,In_1681,In_434);
nand U983 (N_983,In_986,In_2242);
nand U984 (N_984,In_1565,In_1409);
and U985 (N_985,In_2237,In_2143);
or U986 (N_986,In_164,In_650);
nand U987 (N_987,In_1138,In_1292);
nand U988 (N_988,In_718,In_272);
xnor U989 (N_989,In_2304,In_2124);
or U990 (N_990,In_376,In_1146);
and U991 (N_991,In_184,In_2259);
xor U992 (N_992,In_1653,In_922);
xnor U993 (N_993,In_1340,In_489);
or U994 (N_994,In_1917,In_808);
xnor U995 (N_995,In_1931,In_1648);
and U996 (N_996,In_556,In_950);
nand U997 (N_997,In_1828,In_2004);
nor U998 (N_998,In_500,In_128);
xor U999 (N_999,In_43,In_77);
nor U1000 (N_1000,In_2433,In_427);
nand U1001 (N_1001,In_257,In_418);
or U1002 (N_1002,In_2470,In_2489);
nand U1003 (N_1003,In_734,In_1725);
xor U1004 (N_1004,In_690,In_1922);
or U1005 (N_1005,In_1388,In_368);
xor U1006 (N_1006,In_1548,In_1955);
or U1007 (N_1007,In_1248,In_1431);
nor U1008 (N_1008,In_395,In_464);
and U1009 (N_1009,In_2434,In_2348);
and U1010 (N_1010,In_267,In_327);
xnor U1011 (N_1011,In_1580,In_1300);
and U1012 (N_1012,In_2354,In_1795);
nor U1013 (N_1013,In_1284,In_736);
nor U1014 (N_1014,In_831,In_770);
xnor U1015 (N_1015,In_1874,In_511);
nor U1016 (N_1016,In_2042,In_1802);
xor U1017 (N_1017,In_1956,In_2031);
xnor U1018 (N_1018,In_620,In_355);
and U1019 (N_1019,In_2232,In_540);
nor U1020 (N_1020,In_1103,In_160);
nand U1021 (N_1021,In_40,In_273);
nor U1022 (N_1022,In_653,In_2293);
xor U1023 (N_1023,In_2016,In_626);
nor U1024 (N_1024,In_10,In_1986);
or U1025 (N_1025,In_2485,In_987);
xnor U1026 (N_1026,In_744,In_1592);
xnor U1027 (N_1027,In_1351,In_1843);
or U1028 (N_1028,In_915,In_1780);
nor U1029 (N_1029,In_1113,In_1661);
or U1030 (N_1030,In_472,In_1130);
nor U1031 (N_1031,In_1845,In_429);
or U1032 (N_1032,In_1998,In_1313);
xor U1033 (N_1033,In_227,In_442);
or U1034 (N_1034,In_253,In_1230);
xor U1035 (N_1035,In_844,In_2236);
or U1036 (N_1036,In_1866,In_900);
and U1037 (N_1037,In_621,In_1049);
xor U1038 (N_1038,In_416,In_2043);
and U1039 (N_1039,In_634,In_2000);
nand U1040 (N_1040,In_1501,In_1270);
nor U1041 (N_1041,In_2022,In_1161);
nand U1042 (N_1042,In_719,In_197);
xnor U1043 (N_1043,In_38,In_961);
or U1044 (N_1044,In_1549,In_601);
nor U1045 (N_1045,In_1746,In_1181);
or U1046 (N_1046,In_478,In_785);
and U1047 (N_1047,In_2144,In_1301);
xnor U1048 (N_1048,In_27,In_2253);
xor U1049 (N_1049,In_286,In_1325);
and U1050 (N_1050,In_83,In_147);
nand U1051 (N_1051,In_246,In_659);
nand U1052 (N_1052,In_1320,In_682);
xor U1053 (N_1053,In_842,In_2406);
or U1054 (N_1054,In_2493,In_2324);
and U1055 (N_1055,In_277,In_1829);
and U1056 (N_1056,In_571,In_707);
and U1057 (N_1057,In_456,In_2090);
nand U1058 (N_1058,In_268,In_502);
or U1059 (N_1059,In_2126,In_2091);
or U1060 (N_1060,In_200,In_1947);
xnor U1061 (N_1061,In_303,In_1988);
nand U1062 (N_1062,In_1406,In_594);
or U1063 (N_1063,In_1596,In_2172);
xor U1064 (N_1064,In_199,In_158);
or U1065 (N_1065,In_2160,In_1227);
nor U1066 (N_1066,In_321,In_548);
nand U1067 (N_1067,In_2083,In_1219);
nand U1068 (N_1068,In_743,In_2056);
nor U1069 (N_1069,In_1641,In_2196);
nand U1070 (N_1070,In_969,In_1827);
nor U1071 (N_1071,In_2483,In_1554);
nor U1072 (N_1072,In_2059,In_648);
or U1073 (N_1073,In_1464,In_499);
or U1074 (N_1074,In_1107,In_739);
nand U1075 (N_1075,In_711,In_920);
nand U1076 (N_1076,In_2319,In_1419);
nand U1077 (N_1077,In_380,In_688);
xor U1078 (N_1078,In_1195,In_867);
and U1079 (N_1079,In_2048,In_2373);
nand U1080 (N_1080,In_1582,In_2122);
nor U1081 (N_1081,In_435,In_1801);
nor U1082 (N_1082,In_936,In_274);
nand U1083 (N_1083,In_1081,In_1793);
nor U1084 (N_1084,In_1335,In_1096);
or U1085 (N_1085,In_2194,In_279);
or U1086 (N_1086,In_790,In_154);
nand U1087 (N_1087,In_2303,In_1893);
and U1088 (N_1088,In_1127,In_1332);
nor U1089 (N_1089,In_649,In_1716);
nand U1090 (N_1090,In_1444,In_2422);
or U1091 (N_1091,In_1923,In_2266);
xnor U1092 (N_1092,In_716,In_1385);
xnor U1093 (N_1093,In_2239,In_819);
or U1094 (N_1094,In_388,In_1498);
or U1095 (N_1095,In_99,In_62);
and U1096 (N_1096,In_1073,In_2376);
nand U1097 (N_1097,In_1703,In_161);
nor U1098 (N_1098,In_1952,In_133);
or U1099 (N_1099,In_1767,In_320);
nor U1100 (N_1100,In_2358,In_1402);
nand U1101 (N_1101,In_1056,In_1558);
nor U1102 (N_1102,In_491,In_2255);
or U1103 (N_1103,In_1028,In_1562);
nand U1104 (N_1104,In_1063,In_880);
nor U1105 (N_1105,In_1293,In_1722);
and U1106 (N_1106,In_1635,In_1472);
xor U1107 (N_1107,In_1727,In_1737);
nor U1108 (N_1108,In_1612,In_752);
xor U1109 (N_1109,In_2431,In_1366);
and U1110 (N_1110,In_2076,In_583);
and U1111 (N_1111,In_1434,In_1271);
xor U1112 (N_1112,In_2189,In_1624);
nand U1113 (N_1113,In_2451,In_1688);
nor U1114 (N_1114,In_1225,In_2389);
and U1115 (N_1115,In_2198,In_782);
or U1116 (N_1116,In_929,In_2197);
nor U1117 (N_1117,In_1078,In_2273);
xnor U1118 (N_1118,In_509,In_2089);
nand U1119 (N_1119,In_336,In_1787);
nand U1120 (N_1120,In_1647,In_89);
or U1121 (N_1121,In_229,In_397);
nor U1122 (N_1122,In_1071,In_1240);
nand U1123 (N_1123,In_176,In_9);
xnor U1124 (N_1124,In_1567,In_1949);
or U1125 (N_1125,In_1658,In_270);
and U1126 (N_1126,In_2256,In_723);
nand U1127 (N_1127,In_292,In_516);
xnor U1128 (N_1128,In_2420,In_224);
xnor U1129 (N_1129,In_2195,In_1401);
and U1130 (N_1130,In_1817,In_1886);
or U1131 (N_1131,In_364,In_228);
and U1132 (N_1132,In_1374,In_1995);
nor U1133 (N_1133,In_1392,In_2495);
xor U1134 (N_1134,In_13,In_1916);
nor U1135 (N_1135,In_30,In_1471);
nor U1136 (N_1136,In_809,In_1849);
or U1137 (N_1137,In_728,In_2338);
nor U1138 (N_1138,In_2024,In_392);
nor U1139 (N_1139,In_1131,In_1497);
and U1140 (N_1140,In_1024,In_1820);
or U1141 (N_1141,In_1663,In_547);
nor U1142 (N_1142,In_177,In_20);
nor U1143 (N_1143,In_1563,In_1853);
nor U1144 (N_1144,In_2020,In_11);
nor U1145 (N_1145,In_58,In_305);
nand U1146 (N_1146,In_804,In_510);
and U1147 (N_1147,In_503,In_135);
and U1148 (N_1148,In_1197,In_2026);
or U1149 (N_1149,In_1587,In_2112);
and U1150 (N_1150,In_2064,In_1591);
nor U1151 (N_1151,In_163,In_779);
nor U1152 (N_1152,In_2228,In_1425);
and U1153 (N_1153,In_678,In_676);
nand U1154 (N_1154,In_337,In_2150);
nor U1155 (N_1155,In_2152,In_512);
nor U1156 (N_1156,In_1101,In_1390);
xnor U1157 (N_1157,In_1696,In_2442);
nor U1158 (N_1158,In_1306,In_372);
nand U1159 (N_1159,In_1223,In_260);
and U1160 (N_1160,In_811,In_1656);
nand U1161 (N_1161,In_151,In_1919);
xor U1162 (N_1162,In_1417,In_2005);
and U1163 (N_1163,In_285,In_795);
nand U1164 (N_1164,In_1734,In_1742);
and U1165 (N_1165,In_1418,In_1637);
xor U1166 (N_1166,In_374,In_2346);
nor U1167 (N_1167,In_1488,In_2343);
nand U1168 (N_1168,In_1959,In_64);
nand U1169 (N_1169,In_203,In_168);
or U1170 (N_1170,In_537,In_351);
and U1171 (N_1171,In_8,In_1349);
nand U1172 (N_1172,In_107,In_205);
and U1173 (N_1173,In_1601,In_1323);
nand U1174 (N_1174,In_985,In_136);
or U1175 (N_1175,In_2363,In_769);
xnor U1176 (N_1176,In_1076,In_1370);
nor U1177 (N_1177,In_2001,In_1393);
nand U1178 (N_1178,In_2095,In_750);
xor U1179 (N_1179,In_2264,In_1771);
xnor U1180 (N_1180,In_2282,In_441);
nor U1181 (N_1181,In_2462,In_1449);
nand U1182 (N_1182,In_1695,In_330);
and U1183 (N_1183,In_148,In_1436);
xnor U1184 (N_1184,In_1864,In_2209);
or U1185 (N_1185,In_2166,In_111);
and U1186 (N_1186,In_1816,In_2046);
nor U1187 (N_1187,In_281,In_1166);
nand U1188 (N_1188,In_1378,In_2416);
xnor U1189 (N_1189,In_1047,In_2058);
nand U1190 (N_1190,In_850,In_1120);
and U1191 (N_1191,In_732,In_409);
xor U1192 (N_1192,In_80,In_74);
nand U1193 (N_1193,In_784,In_1463);
nor U1194 (N_1194,In_1022,In_468);
or U1195 (N_1195,In_208,In_2100);
nor U1196 (N_1196,In_2142,In_865);
xnor U1197 (N_1197,In_2045,In_370);
xnor U1198 (N_1198,In_1768,In_1983);
and U1199 (N_1199,In_524,In_869);
or U1200 (N_1200,In_1504,In_1143);
and U1201 (N_1201,In_514,In_1584);
nand U1202 (N_1202,In_792,In_872);
nor U1203 (N_1203,In_1973,In_1111);
and U1204 (N_1204,In_1790,In_1882);
and U1205 (N_1205,In_2472,In_1273);
or U1206 (N_1206,In_2115,In_1826);
xnor U1207 (N_1207,In_201,In_2069);
and U1208 (N_1208,In_1158,In_837);
nand U1209 (N_1209,In_1796,In_476);
and U1210 (N_1210,In_1257,In_618);
or U1211 (N_1211,In_1042,In_1857);
or U1212 (N_1212,In_82,In_1339);
nand U1213 (N_1213,In_1814,In_753);
nor U1214 (N_1214,In_115,In_1840);
nand U1215 (N_1215,In_1590,In_195);
and U1216 (N_1216,In_1289,In_669);
nor U1217 (N_1217,In_2168,In_1963);
or U1218 (N_1218,In_2417,In_1057);
and U1219 (N_1219,In_504,In_586);
nand U1220 (N_1220,In_1478,In_607);
nand U1221 (N_1221,In_2278,In_1354);
nor U1222 (N_1222,In_1903,In_1100);
and U1223 (N_1223,In_54,In_44);
or U1224 (N_1224,In_740,In_1206);
and U1225 (N_1225,In_1694,In_2335);
xnor U1226 (N_1226,In_1967,In_306);
nand U1227 (N_1227,In_1652,In_1217);
nand U1228 (N_1228,In_755,In_1958);
and U1229 (N_1229,In_1777,In_1932);
nand U1230 (N_1230,In_1723,In_2252);
or U1231 (N_1231,In_2176,In_340);
or U1232 (N_1232,In_263,In_1510);
or U1233 (N_1233,In_29,In_436);
or U1234 (N_1234,In_103,In_1483);
xor U1235 (N_1235,In_2498,In_572);
and U1236 (N_1236,In_72,In_287);
nor U1237 (N_1237,In_366,In_2205);
or U1238 (N_1238,In_1837,In_2109);
nor U1239 (N_1239,In_885,In_720);
or U1240 (N_1240,In_1630,In_387);
or U1241 (N_1241,In_411,In_675);
or U1242 (N_1242,In_2351,In_2394);
nand U1243 (N_1243,In_1756,In_2011);
xnor U1244 (N_1244,In_140,In_1863);
nand U1245 (N_1245,In_2484,In_1862);
nor U1246 (N_1246,In_256,In_1578);
or U1247 (N_1247,In_1943,In_604);
nor U1248 (N_1248,In_2119,In_1655);
and U1249 (N_1249,In_2199,In_2148);
nor U1250 (N_1250,In_2301,In_384);
nand U1251 (N_1251,In_1698,In_994);
or U1252 (N_1252,In_1665,In_2269);
and U1253 (N_1253,In_795,In_1111);
nand U1254 (N_1254,In_1237,In_1759);
or U1255 (N_1255,In_2379,In_365);
xor U1256 (N_1256,In_954,In_1134);
nor U1257 (N_1257,In_1454,In_1437);
xor U1258 (N_1258,In_612,In_752);
and U1259 (N_1259,In_1041,In_2338);
and U1260 (N_1260,In_120,In_8);
xor U1261 (N_1261,In_292,In_1779);
xor U1262 (N_1262,In_814,In_215);
or U1263 (N_1263,In_173,In_674);
nor U1264 (N_1264,In_834,In_2370);
nor U1265 (N_1265,In_319,In_1475);
and U1266 (N_1266,In_1999,In_1445);
or U1267 (N_1267,In_1274,In_1219);
or U1268 (N_1268,In_977,In_219);
and U1269 (N_1269,In_2288,In_648);
nor U1270 (N_1270,In_1906,In_1247);
or U1271 (N_1271,In_601,In_1868);
nor U1272 (N_1272,In_1164,In_2088);
and U1273 (N_1273,In_2,In_1777);
nand U1274 (N_1274,In_2250,In_326);
nor U1275 (N_1275,In_472,In_2429);
xor U1276 (N_1276,In_1283,In_1435);
xnor U1277 (N_1277,In_508,In_1117);
and U1278 (N_1278,In_2387,In_1375);
or U1279 (N_1279,In_1783,In_1772);
xnor U1280 (N_1280,In_2253,In_2164);
xor U1281 (N_1281,In_801,In_1355);
nor U1282 (N_1282,In_1496,In_2102);
or U1283 (N_1283,In_1947,In_2071);
and U1284 (N_1284,In_730,In_1655);
nor U1285 (N_1285,In_1584,In_931);
nor U1286 (N_1286,In_531,In_2481);
xnor U1287 (N_1287,In_849,In_281);
nor U1288 (N_1288,In_599,In_2024);
xnor U1289 (N_1289,In_1842,In_21);
or U1290 (N_1290,In_1071,In_520);
nand U1291 (N_1291,In_408,In_1105);
nor U1292 (N_1292,In_2349,In_779);
and U1293 (N_1293,In_1486,In_1635);
xnor U1294 (N_1294,In_1581,In_548);
xor U1295 (N_1295,In_929,In_1835);
or U1296 (N_1296,In_1636,In_132);
nand U1297 (N_1297,In_322,In_2449);
nand U1298 (N_1298,In_426,In_1494);
nor U1299 (N_1299,In_1690,In_1517);
nor U1300 (N_1300,In_1379,In_209);
and U1301 (N_1301,In_1347,In_967);
and U1302 (N_1302,In_161,In_1760);
xor U1303 (N_1303,In_470,In_1290);
or U1304 (N_1304,In_401,In_583);
xor U1305 (N_1305,In_420,In_1545);
xor U1306 (N_1306,In_495,In_1805);
nor U1307 (N_1307,In_1575,In_456);
and U1308 (N_1308,In_817,In_886);
xor U1309 (N_1309,In_274,In_1521);
nand U1310 (N_1310,In_132,In_792);
or U1311 (N_1311,In_1849,In_2327);
nor U1312 (N_1312,In_1489,In_17);
nand U1313 (N_1313,In_1194,In_754);
nor U1314 (N_1314,In_2486,In_536);
nand U1315 (N_1315,In_382,In_794);
xor U1316 (N_1316,In_1432,In_1443);
or U1317 (N_1317,In_908,In_2105);
and U1318 (N_1318,In_647,In_889);
nand U1319 (N_1319,In_106,In_504);
xnor U1320 (N_1320,In_1900,In_94);
or U1321 (N_1321,In_2294,In_2038);
and U1322 (N_1322,In_1404,In_1631);
nand U1323 (N_1323,In_2126,In_1678);
xor U1324 (N_1324,In_1848,In_1785);
or U1325 (N_1325,In_1172,In_2317);
or U1326 (N_1326,In_515,In_1589);
nor U1327 (N_1327,In_965,In_1279);
or U1328 (N_1328,In_1035,In_1526);
or U1329 (N_1329,In_1558,In_1326);
or U1330 (N_1330,In_976,In_1055);
and U1331 (N_1331,In_837,In_1796);
nor U1332 (N_1332,In_1904,In_2273);
nand U1333 (N_1333,In_704,In_17);
and U1334 (N_1334,In_2432,In_1558);
nand U1335 (N_1335,In_1514,In_2344);
nor U1336 (N_1336,In_2221,In_2337);
nand U1337 (N_1337,In_1784,In_51);
nor U1338 (N_1338,In_1597,In_0);
nand U1339 (N_1339,In_755,In_2269);
or U1340 (N_1340,In_1373,In_885);
and U1341 (N_1341,In_1625,In_2412);
nand U1342 (N_1342,In_319,In_683);
or U1343 (N_1343,In_2381,In_963);
nand U1344 (N_1344,In_657,In_2430);
xnor U1345 (N_1345,In_969,In_106);
xnor U1346 (N_1346,In_2425,In_2248);
nor U1347 (N_1347,In_1098,In_1385);
xnor U1348 (N_1348,In_181,In_1774);
nand U1349 (N_1349,In_1276,In_612);
nand U1350 (N_1350,In_493,In_1777);
nand U1351 (N_1351,In_1840,In_1920);
and U1352 (N_1352,In_881,In_618);
and U1353 (N_1353,In_89,In_1794);
nor U1354 (N_1354,In_2435,In_371);
nor U1355 (N_1355,In_7,In_1971);
xor U1356 (N_1356,In_1077,In_2144);
nor U1357 (N_1357,In_1313,In_78);
xnor U1358 (N_1358,In_569,In_1083);
and U1359 (N_1359,In_1302,In_1080);
or U1360 (N_1360,In_581,In_1844);
nor U1361 (N_1361,In_2400,In_2270);
nand U1362 (N_1362,In_1627,In_1940);
xor U1363 (N_1363,In_2114,In_606);
xnor U1364 (N_1364,In_2344,In_2407);
or U1365 (N_1365,In_45,In_847);
and U1366 (N_1366,In_571,In_90);
and U1367 (N_1367,In_2224,In_1010);
nor U1368 (N_1368,In_1582,In_1492);
or U1369 (N_1369,In_1191,In_152);
and U1370 (N_1370,In_1884,In_439);
xor U1371 (N_1371,In_1668,In_1864);
xor U1372 (N_1372,In_548,In_172);
nor U1373 (N_1373,In_2159,In_952);
xor U1374 (N_1374,In_2346,In_1662);
and U1375 (N_1375,In_1543,In_42);
or U1376 (N_1376,In_992,In_2293);
nor U1377 (N_1377,In_1027,In_968);
nand U1378 (N_1378,In_2214,In_1064);
xor U1379 (N_1379,In_2094,In_2349);
nand U1380 (N_1380,In_387,In_2298);
or U1381 (N_1381,In_729,In_194);
nor U1382 (N_1382,In_494,In_607);
nor U1383 (N_1383,In_692,In_145);
or U1384 (N_1384,In_1974,In_289);
or U1385 (N_1385,In_1396,In_2469);
nand U1386 (N_1386,In_2494,In_481);
xor U1387 (N_1387,In_122,In_127);
nor U1388 (N_1388,In_1365,In_271);
and U1389 (N_1389,In_1357,In_1776);
xor U1390 (N_1390,In_1469,In_1006);
nand U1391 (N_1391,In_2286,In_2017);
and U1392 (N_1392,In_1569,In_1491);
nand U1393 (N_1393,In_1255,In_2147);
or U1394 (N_1394,In_26,In_2027);
xor U1395 (N_1395,In_561,In_1085);
nor U1396 (N_1396,In_223,In_1103);
xor U1397 (N_1397,In_913,In_2467);
or U1398 (N_1398,In_1430,In_503);
nor U1399 (N_1399,In_741,In_1310);
and U1400 (N_1400,In_256,In_261);
nand U1401 (N_1401,In_641,In_557);
or U1402 (N_1402,In_2329,In_2152);
and U1403 (N_1403,In_1724,In_1760);
and U1404 (N_1404,In_1419,In_125);
nor U1405 (N_1405,In_53,In_542);
nand U1406 (N_1406,In_2040,In_1528);
and U1407 (N_1407,In_1385,In_1075);
xnor U1408 (N_1408,In_1923,In_108);
nor U1409 (N_1409,In_1539,In_627);
nand U1410 (N_1410,In_2106,In_1258);
nand U1411 (N_1411,In_1223,In_2294);
and U1412 (N_1412,In_2268,In_342);
or U1413 (N_1413,In_2233,In_124);
or U1414 (N_1414,In_2437,In_59);
nand U1415 (N_1415,In_259,In_657);
and U1416 (N_1416,In_442,In_1523);
or U1417 (N_1417,In_347,In_1549);
nand U1418 (N_1418,In_2019,In_725);
and U1419 (N_1419,In_882,In_436);
and U1420 (N_1420,In_2163,In_1190);
nor U1421 (N_1421,In_1133,In_1085);
or U1422 (N_1422,In_1942,In_771);
nor U1423 (N_1423,In_1948,In_559);
or U1424 (N_1424,In_672,In_1419);
nand U1425 (N_1425,In_1737,In_1349);
and U1426 (N_1426,In_1238,In_2336);
nand U1427 (N_1427,In_920,In_506);
xor U1428 (N_1428,In_2453,In_2180);
or U1429 (N_1429,In_870,In_1602);
nor U1430 (N_1430,In_466,In_1363);
and U1431 (N_1431,In_126,In_313);
nor U1432 (N_1432,In_892,In_1767);
nor U1433 (N_1433,In_791,In_933);
nor U1434 (N_1434,In_1877,In_2231);
or U1435 (N_1435,In_2453,In_2176);
nand U1436 (N_1436,In_2182,In_1106);
and U1437 (N_1437,In_1792,In_205);
nand U1438 (N_1438,In_1398,In_1297);
xnor U1439 (N_1439,In_1506,In_106);
or U1440 (N_1440,In_1024,In_1594);
nand U1441 (N_1441,In_2065,In_31);
or U1442 (N_1442,In_906,In_488);
or U1443 (N_1443,In_1222,In_86);
nand U1444 (N_1444,In_1510,In_2104);
nor U1445 (N_1445,In_1337,In_1134);
and U1446 (N_1446,In_1199,In_1053);
nand U1447 (N_1447,In_600,In_2491);
nand U1448 (N_1448,In_1301,In_972);
nor U1449 (N_1449,In_242,In_778);
nand U1450 (N_1450,In_983,In_786);
nor U1451 (N_1451,In_442,In_257);
nor U1452 (N_1452,In_101,In_435);
nand U1453 (N_1453,In_982,In_503);
nand U1454 (N_1454,In_143,In_1093);
xor U1455 (N_1455,In_1210,In_1887);
xnor U1456 (N_1456,In_62,In_1699);
and U1457 (N_1457,In_178,In_527);
or U1458 (N_1458,In_460,In_541);
xor U1459 (N_1459,In_1234,In_754);
nor U1460 (N_1460,In_912,In_2306);
nor U1461 (N_1461,In_2022,In_1450);
or U1462 (N_1462,In_1361,In_515);
and U1463 (N_1463,In_528,In_790);
or U1464 (N_1464,In_2101,In_503);
or U1465 (N_1465,In_2450,In_423);
or U1466 (N_1466,In_2083,In_153);
xor U1467 (N_1467,In_1034,In_741);
xnor U1468 (N_1468,In_390,In_1587);
or U1469 (N_1469,In_1212,In_1598);
xnor U1470 (N_1470,In_2259,In_1732);
and U1471 (N_1471,In_974,In_1293);
and U1472 (N_1472,In_1420,In_978);
and U1473 (N_1473,In_183,In_2312);
and U1474 (N_1474,In_517,In_731);
nor U1475 (N_1475,In_256,In_2436);
and U1476 (N_1476,In_1672,In_636);
nand U1477 (N_1477,In_2402,In_533);
and U1478 (N_1478,In_520,In_2404);
nand U1479 (N_1479,In_773,In_238);
nand U1480 (N_1480,In_1632,In_107);
or U1481 (N_1481,In_2277,In_424);
xnor U1482 (N_1482,In_1137,In_1406);
nor U1483 (N_1483,In_2376,In_170);
nand U1484 (N_1484,In_1224,In_1877);
and U1485 (N_1485,In_569,In_2363);
nand U1486 (N_1486,In_956,In_1865);
and U1487 (N_1487,In_1792,In_1169);
nand U1488 (N_1488,In_1580,In_1956);
xnor U1489 (N_1489,In_1836,In_1825);
xor U1490 (N_1490,In_1569,In_1589);
and U1491 (N_1491,In_97,In_24);
xnor U1492 (N_1492,In_2235,In_1723);
nor U1493 (N_1493,In_2322,In_1567);
nand U1494 (N_1494,In_547,In_694);
nor U1495 (N_1495,In_948,In_538);
xor U1496 (N_1496,In_624,In_59);
and U1497 (N_1497,In_2219,In_1208);
nand U1498 (N_1498,In_326,In_747);
or U1499 (N_1499,In_2397,In_1510);
and U1500 (N_1500,In_280,In_1172);
nor U1501 (N_1501,In_1026,In_276);
and U1502 (N_1502,In_3,In_502);
xnor U1503 (N_1503,In_1105,In_1920);
xor U1504 (N_1504,In_1539,In_2008);
nor U1505 (N_1505,In_564,In_668);
or U1506 (N_1506,In_608,In_2293);
and U1507 (N_1507,In_1550,In_282);
or U1508 (N_1508,In_637,In_442);
or U1509 (N_1509,In_1174,In_1622);
nand U1510 (N_1510,In_1953,In_1060);
xor U1511 (N_1511,In_1442,In_397);
and U1512 (N_1512,In_2349,In_1525);
nand U1513 (N_1513,In_1916,In_1688);
xor U1514 (N_1514,In_2391,In_65);
and U1515 (N_1515,In_45,In_1510);
nor U1516 (N_1516,In_1978,In_1775);
nor U1517 (N_1517,In_2159,In_13);
and U1518 (N_1518,In_1214,In_190);
nand U1519 (N_1519,In_1317,In_629);
nor U1520 (N_1520,In_1083,In_2228);
or U1521 (N_1521,In_243,In_1956);
xor U1522 (N_1522,In_441,In_2101);
nor U1523 (N_1523,In_973,In_130);
and U1524 (N_1524,In_2063,In_982);
or U1525 (N_1525,In_2020,In_635);
xor U1526 (N_1526,In_1552,In_2241);
and U1527 (N_1527,In_470,In_2351);
nor U1528 (N_1528,In_1462,In_2282);
nand U1529 (N_1529,In_644,In_722);
nand U1530 (N_1530,In_629,In_1042);
and U1531 (N_1531,In_1203,In_1903);
nor U1532 (N_1532,In_1718,In_1432);
nand U1533 (N_1533,In_2195,In_2241);
or U1534 (N_1534,In_1014,In_957);
or U1535 (N_1535,In_2081,In_330);
or U1536 (N_1536,In_852,In_1246);
nor U1537 (N_1537,In_244,In_548);
or U1538 (N_1538,In_558,In_2317);
nor U1539 (N_1539,In_1820,In_1324);
and U1540 (N_1540,In_1666,In_318);
xor U1541 (N_1541,In_2204,In_651);
xnor U1542 (N_1542,In_2305,In_2194);
or U1543 (N_1543,In_1717,In_28);
nand U1544 (N_1544,In_315,In_2466);
nor U1545 (N_1545,In_1483,In_672);
or U1546 (N_1546,In_2389,In_1688);
nand U1547 (N_1547,In_2345,In_2237);
and U1548 (N_1548,In_2112,In_969);
nand U1549 (N_1549,In_1353,In_2345);
or U1550 (N_1550,In_1296,In_2182);
and U1551 (N_1551,In_1495,In_1997);
xnor U1552 (N_1552,In_369,In_2388);
nand U1553 (N_1553,In_1504,In_1219);
xnor U1554 (N_1554,In_2349,In_139);
nand U1555 (N_1555,In_143,In_634);
and U1556 (N_1556,In_1014,In_846);
nor U1557 (N_1557,In_2240,In_506);
nor U1558 (N_1558,In_2357,In_1224);
or U1559 (N_1559,In_1845,In_2115);
or U1560 (N_1560,In_723,In_1204);
or U1561 (N_1561,In_1676,In_551);
nand U1562 (N_1562,In_1774,In_1160);
xor U1563 (N_1563,In_2423,In_1231);
or U1564 (N_1564,In_1054,In_1986);
and U1565 (N_1565,In_11,In_2416);
nor U1566 (N_1566,In_1395,In_21);
nor U1567 (N_1567,In_488,In_945);
nand U1568 (N_1568,In_414,In_1027);
or U1569 (N_1569,In_1445,In_1341);
xor U1570 (N_1570,In_381,In_1221);
and U1571 (N_1571,In_1665,In_2319);
nand U1572 (N_1572,In_1790,In_1852);
nand U1573 (N_1573,In_676,In_910);
xor U1574 (N_1574,In_1752,In_2058);
and U1575 (N_1575,In_481,In_1277);
and U1576 (N_1576,In_795,In_1033);
nand U1577 (N_1577,In_5,In_1208);
nand U1578 (N_1578,In_2278,In_55);
nand U1579 (N_1579,In_517,In_1766);
nor U1580 (N_1580,In_153,In_1790);
xnor U1581 (N_1581,In_2110,In_2036);
nand U1582 (N_1582,In_1796,In_2229);
and U1583 (N_1583,In_1425,In_612);
and U1584 (N_1584,In_2044,In_1742);
and U1585 (N_1585,In_295,In_374);
or U1586 (N_1586,In_1758,In_423);
or U1587 (N_1587,In_680,In_451);
or U1588 (N_1588,In_2066,In_1755);
nand U1589 (N_1589,In_2275,In_1890);
and U1590 (N_1590,In_1659,In_385);
xnor U1591 (N_1591,In_1163,In_1621);
nand U1592 (N_1592,In_1619,In_780);
nand U1593 (N_1593,In_1086,In_337);
xor U1594 (N_1594,In_475,In_505);
xnor U1595 (N_1595,In_2236,In_2444);
nand U1596 (N_1596,In_1830,In_620);
or U1597 (N_1597,In_1351,In_1240);
nor U1598 (N_1598,In_870,In_198);
nand U1599 (N_1599,In_1416,In_522);
nand U1600 (N_1600,In_2207,In_423);
or U1601 (N_1601,In_255,In_939);
nor U1602 (N_1602,In_1661,In_2036);
nand U1603 (N_1603,In_1974,In_222);
nor U1604 (N_1604,In_23,In_1628);
nor U1605 (N_1605,In_100,In_1078);
xnor U1606 (N_1606,In_1621,In_2419);
nand U1607 (N_1607,In_2248,In_1089);
or U1608 (N_1608,In_266,In_2172);
or U1609 (N_1609,In_1168,In_1506);
or U1610 (N_1610,In_2244,In_2441);
xor U1611 (N_1611,In_2264,In_2188);
or U1612 (N_1612,In_681,In_163);
nand U1613 (N_1613,In_2180,In_2242);
nor U1614 (N_1614,In_587,In_1441);
nor U1615 (N_1615,In_1087,In_118);
or U1616 (N_1616,In_1305,In_1336);
and U1617 (N_1617,In_837,In_1331);
xor U1618 (N_1618,In_1821,In_322);
and U1619 (N_1619,In_601,In_796);
and U1620 (N_1620,In_1422,In_1);
or U1621 (N_1621,In_311,In_1425);
nor U1622 (N_1622,In_1008,In_1210);
and U1623 (N_1623,In_1769,In_1701);
and U1624 (N_1624,In_2162,In_849);
xor U1625 (N_1625,In_1292,In_534);
nor U1626 (N_1626,In_1944,In_2159);
xor U1627 (N_1627,In_500,In_2477);
or U1628 (N_1628,In_754,In_2103);
xor U1629 (N_1629,In_2315,In_1800);
xnor U1630 (N_1630,In_2384,In_1896);
or U1631 (N_1631,In_2090,In_198);
nand U1632 (N_1632,In_1695,In_1857);
or U1633 (N_1633,In_2369,In_1873);
nand U1634 (N_1634,In_367,In_109);
nor U1635 (N_1635,In_1215,In_212);
nand U1636 (N_1636,In_1256,In_256);
and U1637 (N_1637,In_1311,In_2112);
and U1638 (N_1638,In_2229,In_873);
nor U1639 (N_1639,In_1460,In_1195);
xor U1640 (N_1640,In_2168,In_1478);
or U1641 (N_1641,In_759,In_177);
nor U1642 (N_1642,In_1124,In_2188);
nor U1643 (N_1643,In_1262,In_1655);
xnor U1644 (N_1644,In_176,In_1728);
xnor U1645 (N_1645,In_1105,In_379);
nand U1646 (N_1646,In_397,In_571);
or U1647 (N_1647,In_1046,In_262);
and U1648 (N_1648,In_1181,In_794);
or U1649 (N_1649,In_2198,In_2174);
xnor U1650 (N_1650,In_1253,In_57);
or U1651 (N_1651,In_2376,In_410);
nor U1652 (N_1652,In_507,In_1600);
nand U1653 (N_1653,In_1169,In_2403);
and U1654 (N_1654,In_1770,In_1160);
or U1655 (N_1655,In_821,In_1905);
nand U1656 (N_1656,In_152,In_1972);
xnor U1657 (N_1657,In_2123,In_124);
xnor U1658 (N_1658,In_974,In_297);
or U1659 (N_1659,In_1702,In_713);
or U1660 (N_1660,In_1673,In_2439);
xnor U1661 (N_1661,In_2430,In_2495);
or U1662 (N_1662,In_45,In_1151);
nor U1663 (N_1663,In_69,In_1068);
and U1664 (N_1664,In_315,In_1436);
xor U1665 (N_1665,In_409,In_824);
nor U1666 (N_1666,In_1281,In_1235);
and U1667 (N_1667,In_1843,In_2048);
nor U1668 (N_1668,In_1261,In_871);
nand U1669 (N_1669,In_2335,In_519);
xor U1670 (N_1670,In_2333,In_2087);
nand U1671 (N_1671,In_1279,In_2414);
nand U1672 (N_1672,In_405,In_149);
or U1673 (N_1673,In_444,In_1677);
and U1674 (N_1674,In_729,In_2089);
nand U1675 (N_1675,In_1877,In_1330);
nor U1676 (N_1676,In_1167,In_1214);
nand U1677 (N_1677,In_2214,In_2295);
and U1678 (N_1678,In_176,In_2310);
or U1679 (N_1679,In_1743,In_1081);
or U1680 (N_1680,In_837,In_1814);
xor U1681 (N_1681,In_1284,In_1888);
nand U1682 (N_1682,In_1941,In_2308);
nor U1683 (N_1683,In_629,In_556);
and U1684 (N_1684,In_1099,In_1907);
or U1685 (N_1685,In_256,In_1510);
or U1686 (N_1686,In_2252,In_2193);
nand U1687 (N_1687,In_1186,In_1727);
and U1688 (N_1688,In_172,In_1578);
and U1689 (N_1689,In_1992,In_1765);
and U1690 (N_1690,In_516,In_1589);
nand U1691 (N_1691,In_128,In_1574);
nand U1692 (N_1692,In_1960,In_1592);
nand U1693 (N_1693,In_920,In_2279);
and U1694 (N_1694,In_631,In_2242);
xnor U1695 (N_1695,In_469,In_1212);
xnor U1696 (N_1696,In_2278,In_1169);
xor U1697 (N_1697,In_827,In_1164);
or U1698 (N_1698,In_691,In_39);
and U1699 (N_1699,In_638,In_612);
or U1700 (N_1700,In_2035,In_1626);
and U1701 (N_1701,In_144,In_2402);
xnor U1702 (N_1702,In_352,In_2318);
nor U1703 (N_1703,In_995,In_971);
xor U1704 (N_1704,In_1872,In_992);
or U1705 (N_1705,In_767,In_1644);
nand U1706 (N_1706,In_911,In_2168);
nor U1707 (N_1707,In_412,In_1995);
nand U1708 (N_1708,In_342,In_659);
or U1709 (N_1709,In_1183,In_2136);
nor U1710 (N_1710,In_2338,In_297);
nand U1711 (N_1711,In_2432,In_695);
xnor U1712 (N_1712,In_436,In_584);
xor U1713 (N_1713,In_1231,In_1533);
nor U1714 (N_1714,In_634,In_237);
nand U1715 (N_1715,In_1085,In_76);
xnor U1716 (N_1716,In_1803,In_1102);
xnor U1717 (N_1717,In_830,In_2467);
nand U1718 (N_1718,In_2090,In_1367);
and U1719 (N_1719,In_1516,In_1119);
nor U1720 (N_1720,In_815,In_531);
nor U1721 (N_1721,In_733,In_198);
xor U1722 (N_1722,In_1359,In_622);
nand U1723 (N_1723,In_2457,In_240);
and U1724 (N_1724,In_2370,In_724);
and U1725 (N_1725,In_671,In_2110);
xor U1726 (N_1726,In_621,In_451);
and U1727 (N_1727,In_2278,In_2036);
nor U1728 (N_1728,In_2065,In_2097);
xor U1729 (N_1729,In_1902,In_1995);
nor U1730 (N_1730,In_2110,In_1472);
nor U1731 (N_1731,In_1584,In_2426);
nand U1732 (N_1732,In_163,In_1611);
nand U1733 (N_1733,In_1728,In_1930);
nor U1734 (N_1734,In_2243,In_2253);
and U1735 (N_1735,In_2298,In_1895);
nor U1736 (N_1736,In_851,In_1602);
xor U1737 (N_1737,In_830,In_295);
and U1738 (N_1738,In_1408,In_2104);
nor U1739 (N_1739,In_266,In_1169);
xor U1740 (N_1740,In_944,In_2020);
nand U1741 (N_1741,In_977,In_601);
or U1742 (N_1742,In_1914,In_2155);
nor U1743 (N_1743,In_1417,In_861);
or U1744 (N_1744,In_4,In_1367);
or U1745 (N_1745,In_699,In_442);
and U1746 (N_1746,In_2094,In_719);
nor U1747 (N_1747,In_1593,In_1905);
nand U1748 (N_1748,In_2417,In_1203);
nor U1749 (N_1749,In_2140,In_2067);
nor U1750 (N_1750,In_1439,In_1974);
nand U1751 (N_1751,In_2379,In_2097);
and U1752 (N_1752,In_466,In_2302);
nor U1753 (N_1753,In_1718,In_1974);
nor U1754 (N_1754,In_1178,In_1335);
and U1755 (N_1755,In_2280,In_584);
xnor U1756 (N_1756,In_1294,In_1564);
and U1757 (N_1757,In_2013,In_352);
and U1758 (N_1758,In_271,In_2315);
nor U1759 (N_1759,In_846,In_181);
or U1760 (N_1760,In_1020,In_1220);
or U1761 (N_1761,In_289,In_1961);
nand U1762 (N_1762,In_1193,In_2287);
or U1763 (N_1763,In_1967,In_217);
nor U1764 (N_1764,In_231,In_1038);
and U1765 (N_1765,In_2467,In_856);
nor U1766 (N_1766,In_1592,In_1981);
or U1767 (N_1767,In_317,In_665);
or U1768 (N_1768,In_1003,In_516);
and U1769 (N_1769,In_2437,In_2074);
xnor U1770 (N_1770,In_1437,In_1926);
nand U1771 (N_1771,In_1104,In_1757);
nand U1772 (N_1772,In_1376,In_1194);
nor U1773 (N_1773,In_2178,In_2272);
xor U1774 (N_1774,In_1775,In_1700);
nor U1775 (N_1775,In_439,In_2129);
nand U1776 (N_1776,In_583,In_2032);
and U1777 (N_1777,In_391,In_801);
and U1778 (N_1778,In_1294,In_1796);
or U1779 (N_1779,In_2380,In_1369);
and U1780 (N_1780,In_748,In_135);
nor U1781 (N_1781,In_585,In_602);
and U1782 (N_1782,In_1777,In_2293);
or U1783 (N_1783,In_1330,In_911);
nand U1784 (N_1784,In_576,In_2452);
nand U1785 (N_1785,In_2452,In_44);
nor U1786 (N_1786,In_2405,In_2145);
or U1787 (N_1787,In_1628,In_4);
or U1788 (N_1788,In_1562,In_283);
nor U1789 (N_1789,In_384,In_1855);
xnor U1790 (N_1790,In_286,In_149);
or U1791 (N_1791,In_785,In_1135);
or U1792 (N_1792,In_2370,In_2129);
nor U1793 (N_1793,In_191,In_1018);
nor U1794 (N_1794,In_252,In_1677);
nor U1795 (N_1795,In_2060,In_523);
xor U1796 (N_1796,In_2476,In_2190);
or U1797 (N_1797,In_1486,In_731);
and U1798 (N_1798,In_1135,In_1741);
or U1799 (N_1799,In_1416,In_2026);
or U1800 (N_1800,In_1905,In_1321);
and U1801 (N_1801,In_892,In_1194);
and U1802 (N_1802,In_1043,In_2484);
and U1803 (N_1803,In_1554,In_790);
nor U1804 (N_1804,In_1523,In_2268);
nand U1805 (N_1805,In_1349,In_1486);
and U1806 (N_1806,In_1150,In_1397);
nor U1807 (N_1807,In_1478,In_1005);
and U1808 (N_1808,In_347,In_867);
xnor U1809 (N_1809,In_2176,In_1240);
nor U1810 (N_1810,In_1040,In_2042);
nor U1811 (N_1811,In_795,In_1081);
xnor U1812 (N_1812,In_886,In_497);
and U1813 (N_1813,In_377,In_767);
and U1814 (N_1814,In_2109,In_2341);
nor U1815 (N_1815,In_909,In_1270);
xor U1816 (N_1816,In_1379,In_1016);
nor U1817 (N_1817,In_178,In_717);
or U1818 (N_1818,In_2422,In_612);
nor U1819 (N_1819,In_471,In_2104);
and U1820 (N_1820,In_1082,In_388);
nand U1821 (N_1821,In_1206,In_2126);
xnor U1822 (N_1822,In_1659,In_247);
and U1823 (N_1823,In_1175,In_342);
xor U1824 (N_1824,In_903,In_2102);
nand U1825 (N_1825,In_1796,In_1225);
nor U1826 (N_1826,In_61,In_1364);
and U1827 (N_1827,In_1514,In_588);
nand U1828 (N_1828,In_681,In_877);
and U1829 (N_1829,In_533,In_50);
and U1830 (N_1830,In_2021,In_332);
nand U1831 (N_1831,In_1973,In_227);
nand U1832 (N_1832,In_1412,In_2177);
nor U1833 (N_1833,In_1983,In_1947);
nor U1834 (N_1834,In_802,In_729);
nand U1835 (N_1835,In_1746,In_819);
and U1836 (N_1836,In_941,In_764);
xnor U1837 (N_1837,In_2351,In_2005);
nor U1838 (N_1838,In_1962,In_2062);
or U1839 (N_1839,In_1945,In_932);
nand U1840 (N_1840,In_2329,In_1979);
or U1841 (N_1841,In_671,In_744);
nand U1842 (N_1842,In_815,In_1722);
or U1843 (N_1843,In_882,In_1156);
nor U1844 (N_1844,In_710,In_1922);
and U1845 (N_1845,In_2134,In_2408);
nor U1846 (N_1846,In_915,In_414);
nor U1847 (N_1847,In_125,In_2408);
xor U1848 (N_1848,In_1805,In_1536);
xnor U1849 (N_1849,In_2299,In_1264);
nand U1850 (N_1850,In_1390,In_1324);
or U1851 (N_1851,In_1519,In_1089);
nand U1852 (N_1852,In_969,In_883);
nand U1853 (N_1853,In_798,In_1853);
or U1854 (N_1854,In_1049,In_1202);
xor U1855 (N_1855,In_2159,In_1636);
xnor U1856 (N_1856,In_1600,In_971);
or U1857 (N_1857,In_1133,In_834);
and U1858 (N_1858,In_1380,In_1848);
and U1859 (N_1859,In_1310,In_536);
and U1860 (N_1860,In_2311,In_150);
nand U1861 (N_1861,In_1402,In_1220);
nor U1862 (N_1862,In_2140,In_1970);
and U1863 (N_1863,In_50,In_235);
or U1864 (N_1864,In_43,In_1565);
nand U1865 (N_1865,In_2341,In_190);
or U1866 (N_1866,In_1127,In_2127);
nand U1867 (N_1867,In_661,In_1822);
or U1868 (N_1868,In_32,In_1102);
nor U1869 (N_1869,In_856,In_767);
or U1870 (N_1870,In_1463,In_2222);
and U1871 (N_1871,In_412,In_864);
and U1872 (N_1872,In_2053,In_2314);
and U1873 (N_1873,In_412,In_1274);
nand U1874 (N_1874,In_828,In_2368);
or U1875 (N_1875,In_2301,In_353);
xor U1876 (N_1876,In_1500,In_2383);
or U1877 (N_1877,In_2180,In_1760);
and U1878 (N_1878,In_1121,In_630);
nand U1879 (N_1879,In_878,In_1310);
or U1880 (N_1880,In_2373,In_1381);
nor U1881 (N_1881,In_2033,In_1876);
xor U1882 (N_1882,In_714,In_1831);
nor U1883 (N_1883,In_1271,In_1221);
nor U1884 (N_1884,In_2050,In_1037);
and U1885 (N_1885,In_643,In_1857);
nand U1886 (N_1886,In_1188,In_1168);
nor U1887 (N_1887,In_1890,In_1402);
xnor U1888 (N_1888,In_1266,In_1512);
or U1889 (N_1889,In_1813,In_1658);
or U1890 (N_1890,In_1766,In_1852);
nand U1891 (N_1891,In_617,In_2453);
or U1892 (N_1892,In_518,In_1206);
xor U1893 (N_1893,In_752,In_525);
xor U1894 (N_1894,In_56,In_2240);
and U1895 (N_1895,In_1694,In_2012);
and U1896 (N_1896,In_1968,In_2466);
or U1897 (N_1897,In_688,In_236);
and U1898 (N_1898,In_2138,In_2330);
and U1899 (N_1899,In_490,In_131);
and U1900 (N_1900,In_261,In_1255);
or U1901 (N_1901,In_352,In_1614);
xnor U1902 (N_1902,In_1093,In_1727);
nor U1903 (N_1903,In_1925,In_2099);
or U1904 (N_1904,In_942,In_463);
and U1905 (N_1905,In_1640,In_1688);
nand U1906 (N_1906,In_2403,In_1425);
nor U1907 (N_1907,In_1571,In_2425);
nand U1908 (N_1908,In_2065,In_71);
xor U1909 (N_1909,In_1772,In_2052);
and U1910 (N_1910,In_2278,In_2022);
xor U1911 (N_1911,In_419,In_186);
nor U1912 (N_1912,In_655,In_946);
and U1913 (N_1913,In_2259,In_1573);
and U1914 (N_1914,In_104,In_1723);
nor U1915 (N_1915,In_2098,In_1104);
nor U1916 (N_1916,In_583,In_800);
and U1917 (N_1917,In_442,In_769);
xor U1918 (N_1918,In_472,In_1072);
nand U1919 (N_1919,In_442,In_1398);
nor U1920 (N_1920,In_274,In_899);
nand U1921 (N_1921,In_2334,In_63);
xor U1922 (N_1922,In_2347,In_2433);
and U1923 (N_1923,In_1673,In_1576);
xor U1924 (N_1924,In_186,In_2410);
xor U1925 (N_1925,In_1073,In_2130);
nor U1926 (N_1926,In_673,In_1445);
xnor U1927 (N_1927,In_964,In_595);
xor U1928 (N_1928,In_1026,In_907);
or U1929 (N_1929,In_1192,In_865);
and U1930 (N_1930,In_319,In_1637);
xnor U1931 (N_1931,In_1884,In_2002);
nand U1932 (N_1932,In_1453,In_294);
or U1933 (N_1933,In_1999,In_1353);
nand U1934 (N_1934,In_1116,In_122);
nor U1935 (N_1935,In_288,In_1712);
and U1936 (N_1936,In_441,In_2363);
nor U1937 (N_1937,In_552,In_1693);
and U1938 (N_1938,In_1708,In_1502);
nor U1939 (N_1939,In_151,In_1557);
and U1940 (N_1940,In_2469,In_2169);
nor U1941 (N_1941,In_879,In_2125);
xor U1942 (N_1942,In_72,In_484);
xor U1943 (N_1943,In_2258,In_2178);
nor U1944 (N_1944,In_358,In_1517);
and U1945 (N_1945,In_1537,In_764);
and U1946 (N_1946,In_552,In_917);
nand U1947 (N_1947,In_239,In_292);
nor U1948 (N_1948,In_1857,In_340);
nand U1949 (N_1949,In_339,In_2248);
nor U1950 (N_1950,In_841,In_2361);
nor U1951 (N_1951,In_548,In_2432);
xnor U1952 (N_1952,In_345,In_1177);
or U1953 (N_1953,In_1726,In_1961);
and U1954 (N_1954,In_1266,In_1327);
or U1955 (N_1955,In_2390,In_1617);
nand U1956 (N_1956,In_2144,In_2165);
nor U1957 (N_1957,In_46,In_743);
or U1958 (N_1958,In_1882,In_1511);
and U1959 (N_1959,In_2284,In_1587);
nand U1960 (N_1960,In_1208,In_1593);
nor U1961 (N_1961,In_2245,In_1721);
nand U1962 (N_1962,In_229,In_1511);
nand U1963 (N_1963,In_1513,In_67);
and U1964 (N_1964,In_2270,In_2377);
or U1965 (N_1965,In_899,In_961);
and U1966 (N_1966,In_1663,In_951);
or U1967 (N_1967,In_45,In_865);
nand U1968 (N_1968,In_38,In_1508);
or U1969 (N_1969,In_1658,In_1995);
or U1970 (N_1970,In_1412,In_1163);
and U1971 (N_1971,In_2180,In_312);
nor U1972 (N_1972,In_750,In_2100);
nand U1973 (N_1973,In_701,In_2406);
xnor U1974 (N_1974,In_1411,In_1250);
nand U1975 (N_1975,In_355,In_892);
xnor U1976 (N_1976,In_404,In_1315);
nor U1977 (N_1977,In_1994,In_1525);
nor U1978 (N_1978,In_1051,In_1877);
nand U1979 (N_1979,In_34,In_236);
and U1980 (N_1980,In_1241,In_842);
nor U1981 (N_1981,In_2194,In_1581);
and U1982 (N_1982,In_1473,In_1299);
or U1983 (N_1983,In_283,In_1308);
xor U1984 (N_1984,In_2022,In_195);
nand U1985 (N_1985,In_1196,In_228);
nand U1986 (N_1986,In_1862,In_2004);
and U1987 (N_1987,In_1433,In_1595);
xnor U1988 (N_1988,In_2403,In_1992);
nor U1989 (N_1989,In_1286,In_1693);
nand U1990 (N_1990,In_1001,In_1387);
xnor U1991 (N_1991,In_1572,In_305);
and U1992 (N_1992,In_2369,In_802);
nor U1993 (N_1993,In_1477,In_2342);
and U1994 (N_1994,In_1966,In_2196);
nand U1995 (N_1995,In_504,In_1300);
xnor U1996 (N_1996,In_2093,In_1764);
and U1997 (N_1997,In_2430,In_1717);
xnor U1998 (N_1998,In_1506,In_1014);
nor U1999 (N_1999,In_118,In_540);
nor U2000 (N_2000,In_724,In_803);
nand U2001 (N_2001,In_2457,In_528);
and U2002 (N_2002,In_1737,In_570);
nand U2003 (N_2003,In_1846,In_1147);
and U2004 (N_2004,In_291,In_1039);
nand U2005 (N_2005,In_1078,In_2323);
and U2006 (N_2006,In_1818,In_43);
or U2007 (N_2007,In_586,In_1057);
nand U2008 (N_2008,In_541,In_82);
and U2009 (N_2009,In_93,In_21);
or U2010 (N_2010,In_629,In_646);
and U2011 (N_2011,In_857,In_1941);
and U2012 (N_2012,In_83,In_1554);
and U2013 (N_2013,In_2375,In_1087);
nor U2014 (N_2014,In_2148,In_2413);
xnor U2015 (N_2015,In_139,In_1097);
or U2016 (N_2016,In_1527,In_128);
nor U2017 (N_2017,In_298,In_2166);
or U2018 (N_2018,In_1468,In_2213);
nor U2019 (N_2019,In_906,In_2234);
nand U2020 (N_2020,In_2492,In_612);
nor U2021 (N_2021,In_184,In_2473);
xnor U2022 (N_2022,In_1975,In_528);
or U2023 (N_2023,In_2217,In_2464);
xor U2024 (N_2024,In_271,In_272);
xnor U2025 (N_2025,In_1436,In_2410);
nor U2026 (N_2026,In_1909,In_517);
or U2027 (N_2027,In_2066,In_2347);
and U2028 (N_2028,In_764,In_341);
xor U2029 (N_2029,In_1198,In_2073);
nor U2030 (N_2030,In_238,In_2359);
and U2031 (N_2031,In_1322,In_2252);
xnor U2032 (N_2032,In_1446,In_121);
xor U2033 (N_2033,In_1029,In_812);
nor U2034 (N_2034,In_1083,In_1505);
nand U2035 (N_2035,In_2341,In_1137);
xor U2036 (N_2036,In_1354,In_1117);
or U2037 (N_2037,In_139,In_1987);
and U2038 (N_2038,In_1703,In_929);
nor U2039 (N_2039,In_2422,In_703);
nor U2040 (N_2040,In_2314,In_171);
nor U2041 (N_2041,In_1826,In_1487);
and U2042 (N_2042,In_2164,In_1409);
or U2043 (N_2043,In_1603,In_1543);
nand U2044 (N_2044,In_795,In_1945);
or U2045 (N_2045,In_238,In_1161);
or U2046 (N_2046,In_141,In_1121);
or U2047 (N_2047,In_1164,In_187);
and U2048 (N_2048,In_877,In_1792);
nor U2049 (N_2049,In_174,In_674);
or U2050 (N_2050,In_1021,In_998);
and U2051 (N_2051,In_1259,In_568);
or U2052 (N_2052,In_1998,In_2326);
xor U2053 (N_2053,In_2211,In_1061);
or U2054 (N_2054,In_119,In_1530);
or U2055 (N_2055,In_1879,In_2187);
or U2056 (N_2056,In_1761,In_1963);
nor U2057 (N_2057,In_83,In_2441);
nor U2058 (N_2058,In_1345,In_502);
or U2059 (N_2059,In_1002,In_2177);
or U2060 (N_2060,In_2354,In_2369);
xor U2061 (N_2061,In_1008,In_1433);
nand U2062 (N_2062,In_2480,In_1626);
nor U2063 (N_2063,In_745,In_511);
nand U2064 (N_2064,In_863,In_22);
nand U2065 (N_2065,In_1802,In_90);
xnor U2066 (N_2066,In_304,In_1930);
or U2067 (N_2067,In_2372,In_803);
nor U2068 (N_2068,In_2255,In_1322);
or U2069 (N_2069,In_1299,In_2461);
and U2070 (N_2070,In_1095,In_1991);
and U2071 (N_2071,In_849,In_1618);
or U2072 (N_2072,In_864,In_243);
nand U2073 (N_2073,In_2112,In_1917);
nor U2074 (N_2074,In_1125,In_542);
nor U2075 (N_2075,In_1362,In_1724);
or U2076 (N_2076,In_1344,In_2174);
nor U2077 (N_2077,In_2114,In_716);
nand U2078 (N_2078,In_1253,In_2302);
xnor U2079 (N_2079,In_695,In_956);
xnor U2080 (N_2080,In_1820,In_1844);
and U2081 (N_2081,In_1773,In_2266);
nand U2082 (N_2082,In_1145,In_1101);
and U2083 (N_2083,In_425,In_1902);
and U2084 (N_2084,In_774,In_1303);
and U2085 (N_2085,In_788,In_1143);
nor U2086 (N_2086,In_688,In_1694);
nor U2087 (N_2087,In_1313,In_1988);
or U2088 (N_2088,In_2227,In_937);
nor U2089 (N_2089,In_2301,In_637);
nor U2090 (N_2090,In_1301,In_1745);
or U2091 (N_2091,In_1628,In_764);
xnor U2092 (N_2092,In_1292,In_2431);
nor U2093 (N_2093,In_2219,In_1218);
xnor U2094 (N_2094,In_289,In_2252);
xnor U2095 (N_2095,In_2257,In_244);
and U2096 (N_2096,In_871,In_254);
or U2097 (N_2097,In_149,In_2377);
nand U2098 (N_2098,In_94,In_539);
or U2099 (N_2099,In_1985,In_1835);
nor U2100 (N_2100,In_2455,In_1342);
and U2101 (N_2101,In_1628,In_1533);
nand U2102 (N_2102,In_1894,In_1880);
or U2103 (N_2103,In_1247,In_1829);
xnor U2104 (N_2104,In_959,In_252);
and U2105 (N_2105,In_862,In_808);
and U2106 (N_2106,In_1388,In_1357);
or U2107 (N_2107,In_25,In_1816);
and U2108 (N_2108,In_1424,In_159);
nand U2109 (N_2109,In_857,In_116);
xnor U2110 (N_2110,In_175,In_1812);
nor U2111 (N_2111,In_1073,In_1879);
and U2112 (N_2112,In_1815,In_1816);
or U2113 (N_2113,In_897,In_2378);
xnor U2114 (N_2114,In_904,In_1149);
nor U2115 (N_2115,In_1999,In_449);
xnor U2116 (N_2116,In_808,In_1278);
nand U2117 (N_2117,In_496,In_730);
or U2118 (N_2118,In_1208,In_796);
and U2119 (N_2119,In_1872,In_89);
and U2120 (N_2120,In_1599,In_1465);
and U2121 (N_2121,In_1208,In_801);
nand U2122 (N_2122,In_1104,In_796);
or U2123 (N_2123,In_836,In_853);
nor U2124 (N_2124,In_550,In_517);
xor U2125 (N_2125,In_1961,In_420);
and U2126 (N_2126,In_1193,In_1599);
and U2127 (N_2127,In_1540,In_782);
nor U2128 (N_2128,In_368,In_649);
or U2129 (N_2129,In_1153,In_2198);
nor U2130 (N_2130,In_245,In_1889);
nand U2131 (N_2131,In_1372,In_19);
nand U2132 (N_2132,In_3,In_1045);
nor U2133 (N_2133,In_2280,In_2354);
or U2134 (N_2134,In_989,In_1710);
or U2135 (N_2135,In_2303,In_2269);
xnor U2136 (N_2136,In_1427,In_944);
nor U2137 (N_2137,In_2487,In_2007);
xnor U2138 (N_2138,In_1780,In_639);
and U2139 (N_2139,In_1432,In_1200);
nand U2140 (N_2140,In_396,In_1175);
and U2141 (N_2141,In_2157,In_472);
nand U2142 (N_2142,In_909,In_2032);
nor U2143 (N_2143,In_1552,In_1439);
nor U2144 (N_2144,In_375,In_783);
nand U2145 (N_2145,In_952,In_1403);
nand U2146 (N_2146,In_2064,In_2190);
xor U2147 (N_2147,In_15,In_1076);
or U2148 (N_2148,In_2196,In_1650);
nand U2149 (N_2149,In_1179,In_83);
xor U2150 (N_2150,In_1861,In_1800);
or U2151 (N_2151,In_246,In_2201);
and U2152 (N_2152,In_2479,In_1230);
nor U2153 (N_2153,In_1767,In_1286);
nand U2154 (N_2154,In_198,In_683);
xor U2155 (N_2155,In_1034,In_105);
and U2156 (N_2156,In_1410,In_2044);
and U2157 (N_2157,In_1433,In_153);
and U2158 (N_2158,In_2149,In_473);
or U2159 (N_2159,In_1272,In_2275);
nand U2160 (N_2160,In_2376,In_532);
nand U2161 (N_2161,In_2287,In_945);
xnor U2162 (N_2162,In_43,In_379);
nand U2163 (N_2163,In_467,In_181);
nand U2164 (N_2164,In_181,In_1910);
or U2165 (N_2165,In_1533,In_1778);
nand U2166 (N_2166,In_1095,In_2279);
nand U2167 (N_2167,In_1467,In_1075);
nor U2168 (N_2168,In_2331,In_1014);
xor U2169 (N_2169,In_173,In_1671);
xor U2170 (N_2170,In_1517,In_1062);
nand U2171 (N_2171,In_1784,In_1123);
xnor U2172 (N_2172,In_1372,In_2302);
xor U2173 (N_2173,In_1055,In_1752);
xnor U2174 (N_2174,In_1852,In_1659);
or U2175 (N_2175,In_995,In_1120);
nand U2176 (N_2176,In_2029,In_1689);
nor U2177 (N_2177,In_1520,In_2207);
nor U2178 (N_2178,In_1775,In_1813);
nor U2179 (N_2179,In_1817,In_2375);
xor U2180 (N_2180,In_374,In_857);
xor U2181 (N_2181,In_476,In_1844);
or U2182 (N_2182,In_1410,In_1134);
and U2183 (N_2183,In_1876,In_1496);
or U2184 (N_2184,In_2184,In_2234);
or U2185 (N_2185,In_1960,In_325);
or U2186 (N_2186,In_631,In_1786);
and U2187 (N_2187,In_2180,In_1644);
and U2188 (N_2188,In_1321,In_1582);
nand U2189 (N_2189,In_670,In_339);
nor U2190 (N_2190,In_1199,In_1770);
nor U2191 (N_2191,In_1698,In_1077);
and U2192 (N_2192,In_510,In_186);
xnor U2193 (N_2193,In_1008,In_180);
nor U2194 (N_2194,In_1697,In_2101);
nand U2195 (N_2195,In_1906,In_358);
xor U2196 (N_2196,In_673,In_1915);
xnor U2197 (N_2197,In_1600,In_491);
xor U2198 (N_2198,In_1374,In_630);
and U2199 (N_2199,In_1323,In_439);
and U2200 (N_2200,In_1100,In_2335);
nor U2201 (N_2201,In_876,In_2099);
nor U2202 (N_2202,In_136,In_1552);
xnor U2203 (N_2203,In_93,In_1711);
and U2204 (N_2204,In_2116,In_1890);
nand U2205 (N_2205,In_946,In_2093);
xnor U2206 (N_2206,In_1169,In_2053);
or U2207 (N_2207,In_1156,In_1830);
xnor U2208 (N_2208,In_2476,In_1898);
nor U2209 (N_2209,In_1929,In_1920);
nand U2210 (N_2210,In_1809,In_1851);
nand U2211 (N_2211,In_1215,In_208);
and U2212 (N_2212,In_1376,In_2095);
or U2213 (N_2213,In_2210,In_831);
and U2214 (N_2214,In_1216,In_1191);
xnor U2215 (N_2215,In_65,In_1362);
and U2216 (N_2216,In_475,In_1864);
or U2217 (N_2217,In_1433,In_1280);
xnor U2218 (N_2218,In_619,In_2060);
and U2219 (N_2219,In_1760,In_669);
nand U2220 (N_2220,In_246,In_1968);
nor U2221 (N_2221,In_1274,In_925);
nor U2222 (N_2222,In_1885,In_1089);
nor U2223 (N_2223,In_1872,In_2062);
nand U2224 (N_2224,In_582,In_2335);
or U2225 (N_2225,In_1115,In_2107);
nor U2226 (N_2226,In_1014,In_384);
nor U2227 (N_2227,In_846,In_1249);
nor U2228 (N_2228,In_44,In_1835);
and U2229 (N_2229,In_1452,In_1183);
nand U2230 (N_2230,In_1913,In_1769);
nor U2231 (N_2231,In_391,In_1691);
or U2232 (N_2232,In_2244,In_1037);
or U2233 (N_2233,In_2338,In_1138);
nor U2234 (N_2234,In_642,In_488);
and U2235 (N_2235,In_1036,In_2021);
xor U2236 (N_2236,In_14,In_1711);
nor U2237 (N_2237,In_1528,In_718);
and U2238 (N_2238,In_1226,In_363);
xnor U2239 (N_2239,In_1428,In_928);
or U2240 (N_2240,In_1066,In_1344);
or U2241 (N_2241,In_1092,In_863);
nand U2242 (N_2242,In_2302,In_1795);
or U2243 (N_2243,In_121,In_2163);
and U2244 (N_2244,In_1980,In_852);
or U2245 (N_2245,In_135,In_49);
or U2246 (N_2246,In_868,In_497);
or U2247 (N_2247,In_1995,In_833);
nand U2248 (N_2248,In_2304,In_2455);
nor U2249 (N_2249,In_1641,In_2386);
nand U2250 (N_2250,In_281,In_1957);
and U2251 (N_2251,In_134,In_975);
xnor U2252 (N_2252,In_998,In_1036);
or U2253 (N_2253,In_1004,In_430);
or U2254 (N_2254,In_81,In_2360);
and U2255 (N_2255,In_1968,In_621);
and U2256 (N_2256,In_854,In_326);
or U2257 (N_2257,In_1352,In_1178);
or U2258 (N_2258,In_2378,In_2145);
xor U2259 (N_2259,In_522,In_1837);
xor U2260 (N_2260,In_1631,In_600);
nand U2261 (N_2261,In_1384,In_2478);
and U2262 (N_2262,In_666,In_1801);
or U2263 (N_2263,In_1576,In_866);
nand U2264 (N_2264,In_2376,In_430);
nand U2265 (N_2265,In_2209,In_1369);
nor U2266 (N_2266,In_326,In_1207);
nor U2267 (N_2267,In_2142,In_2405);
xnor U2268 (N_2268,In_283,In_1028);
or U2269 (N_2269,In_990,In_1129);
nor U2270 (N_2270,In_673,In_1662);
or U2271 (N_2271,In_1619,In_504);
xor U2272 (N_2272,In_1398,In_1999);
or U2273 (N_2273,In_92,In_2404);
xnor U2274 (N_2274,In_1367,In_1007);
and U2275 (N_2275,In_1673,In_691);
xnor U2276 (N_2276,In_2497,In_1828);
and U2277 (N_2277,In_801,In_1934);
xnor U2278 (N_2278,In_613,In_2335);
and U2279 (N_2279,In_624,In_2344);
xor U2280 (N_2280,In_710,In_2012);
nand U2281 (N_2281,In_1471,In_3);
or U2282 (N_2282,In_844,In_517);
xnor U2283 (N_2283,In_791,In_1953);
and U2284 (N_2284,In_1966,In_301);
xnor U2285 (N_2285,In_1178,In_580);
and U2286 (N_2286,In_2058,In_639);
nand U2287 (N_2287,In_1645,In_1917);
xor U2288 (N_2288,In_2408,In_907);
or U2289 (N_2289,In_344,In_555);
nor U2290 (N_2290,In_2434,In_1585);
or U2291 (N_2291,In_409,In_144);
nor U2292 (N_2292,In_1030,In_1918);
or U2293 (N_2293,In_661,In_2377);
xor U2294 (N_2294,In_2175,In_346);
xnor U2295 (N_2295,In_794,In_331);
nand U2296 (N_2296,In_805,In_2217);
and U2297 (N_2297,In_2187,In_2004);
or U2298 (N_2298,In_2028,In_2412);
and U2299 (N_2299,In_1943,In_539);
nor U2300 (N_2300,In_1973,In_191);
or U2301 (N_2301,In_494,In_55);
and U2302 (N_2302,In_164,In_1341);
xnor U2303 (N_2303,In_1208,In_713);
and U2304 (N_2304,In_1493,In_1400);
nand U2305 (N_2305,In_1091,In_1574);
nor U2306 (N_2306,In_2104,In_2397);
nand U2307 (N_2307,In_250,In_1387);
and U2308 (N_2308,In_765,In_2192);
and U2309 (N_2309,In_104,In_405);
nand U2310 (N_2310,In_80,In_1990);
or U2311 (N_2311,In_1686,In_116);
nand U2312 (N_2312,In_683,In_671);
and U2313 (N_2313,In_1488,In_1285);
nand U2314 (N_2314,In_20,In_858);
xor U2315 (N_2315,In_1762,In_1441);
and U2316 (N_2316,In_490,In_1614);
and U2317 (N_2317,In_373,In_1510);
xor U2318 (N_2318,In_1350,In_2261);
nand U2319 (N_2319,In_186,In_301);
nor U2320 (N_2320,In_332,In_1712);
xnor U2321 (N_2321,In_1390,In_454);
nor U2322 (N_2322,In_227,In_310);
nor U2323 (N_2323,In_1185,In_1906);
or U2324 (N_2324,In_783,In_955);
and U2325 (N_2325,In_792,In_660);
and U2326 (N_2326,In_660,In_1899);
or U2327 (N_2327,In_275,In_443);
and U2328 (N_2328,In_187,In_961);
and U2329 (N_2329,In_352,In_2211);
xnor U2330 (N_2330,In_2213,In_1487);
and U2331 (N_2331,In_1469,In_140);
nor U2332 (N_2332,In_381,In_2106);
nor U2333 (N_2333,In_1350,In_1464);
nor U2334 (N_2334,In_1919,In_2256);
nor U2335 (N_2335,In_1615,In_1223);
xnor U2336 (N_2336,In_2188,In_1649);
and U2337 (N_2337,In_481,In_622);
nand U2338 (N_2338,In_901,In_2172);
or U2339 (N_2339,In_1393,In_1659);
nand U2340 (N_2340,In_1337,In_2107);
or U2341 (N_2341,In_156,In_878);
and U2342 (N_2342,In_970,In_1566);
xnor U2343 (N_2343,In_1990,In_954);
nand U2344 (N_2344,In_2453,In_2211);
xnor U2345 (N_2345,In_1942,In_1544);
nor U2346 (N_2346,In_327,In_376);
xor U2347 (N_2347,In_1641,In_313);
nand U2348 (N_2348,In_1627,In_1531);
nor U2349 (N_2349,In_352,In_1054);
or U2350 (N_2350,In_885,In_942);
nand U2351 (N_2351,In_437,In_398);
nand U2352 (N_2352,In_1057,In_1063);
xnor U2353 (N_2353,In_731,In_1062);
xnor U2354 (N_2354,In_136,In_1795);
nor U2355 (N_2355,In_1765,In_459);
nand U2356 (N_2356,In_868,In_552);
nor U2357 (N_2357,In_2018,In_1284);
or U2358 (N_2358,In_509,In_221);
and U2359 (N_2359,In_895,In_1201);
nor U2360 (N_2360,In_2085,In_1972);
xnor U2361 (N_2361,In_1375,In_1955);
nand U2362 (N_2362,In_510,In_1073);
xor U2363 (N_2363,In_2379,In_1252);
nor U2364 (N_2364,In_2361,In_1046);
or U2365 (N_2365,In_1481,In_1393);
and U2366 (N_2366,In_331,In_1143);
xnor U2367 (N_2367,In_2108,In_360);
or U2368 (N_2368,In_949,In_1256);
nor U2369 (N_2369,In_730,In_1200);
nor U2370 (N_2370,In_1029,In_2162);
and U2371 (N_2371,In_2187,In_867);
xnor U2372 (N_2372,In_1753,In_1247);
nor U2373 (N_2373,In_1605,In_1003);
and U2374 (N_2374,In_476,In_231);
nand U2375 (N_2375,In_159,In_59);
xnor U2376 (N_2376,In_912,In_1980);
nor U2377 (N_2377,In_390,In_1627);
nor U2378 (N_2378,In_1385,In_1384);
or U2379 (N_2379,In_50,In_1323);
xor U2380 (N_2380,In_946,In_2416);
or U2381 (N_2381,In_2317,In_147);
xor U2382 (N_2382,In_1220,In_472);
nand U2383 (N_2383,In_2111,In_1712);
nand U2384 (N_2384,In_747,In_107);
nor U2385 (N_2385,In_107,In_2335);
or U2386 (N_2386,In_779,In_560);
or U2387 (N_2387,In_611,In_921);
or U2388 (N_2388,In_838,In_1813);
xor U2389 (N_2389,In_512,In_1657);
or U2390 (N_2390,In_1404,In_85);
and U2391 (N_2391,In_1337,In_2130);
nand U2392 (N_2392,In_1867,In_1656);
nand U2393 (N_2393,In_1209,In_67);
nor U2394 (N_2394,In_125,In_2470);
or U2395 (N_2395,In_2417,In_306);
or U2396 (N_2396,In_1807,In_344);
nand U2397 (N_2397,In_55,In_653);
or U2398 (N_2398,In_1246,In_2303);
or U2399 (N_2399,In_726,In_1673);
or U2400 (N_2400,In_755,In_1459);
and U2401 (N_2401,In_57,In_42);
nor U2402 (N_2402,In_1484,In_1707);
xor U2403 (N_2403,In_393,In_2482);
or U2404 (N_2404,In_2097,In_336);
xor U2405 (N_2405,In_419,In_26);
and U2406 (N_2406,In_2052,In_1331);
nand U2407 (N_2407,In_251,In_1772);
nand U2408 (N_2408,In_503,In_245);
xnor U2409 (N_2409,In_1293,In_1667);
nor U2410 (N_2410,In_45,In_2053);
xor U2411 (N_2411,In_1574,In_464);
xnor U2412 (N_2412,In_19,In_1214);
and U2413 (N_2413,In_1330,In_173);
and U2414 (N_2414,In_1556,In_1152);
and U2415 (N_2415,In_1924,In_511);
and U2416 (N_2416,In_1948,In_455);
and U2417 (N_2417,In_1821,In_2230);
nand U2418 (N_2418,In_915,In_2474);
nor U2419 (N_2419,In_810,In_1495);
nor U2420 (N_2420,In_2259,In_2425);
or U2421 (N_2421,In_2419,In_59);
or U2422 (N_2422,In_522,In_132);
xor U2423 (N_2423,In_327,In_2221);
and U2424 (N_2424,In_1635,In_1239);
nand U2425 (N_2425,In_1509,In_2412);
nor U2426 (N_2426,In_903,In_1854);
xnor U2427 (N_2427,In_486,In_2206);
and U2428 (N_2428,In_2079,In_535);
nor U2429 (N_2429,In_2211,In_491);
nand U2430 (N_2430,In_1,In_1546);
and U2431 (N_2431,In_530,In_1344);
or U2432 (N_2432,In_1300,In_1390);
xor U2433 (N_2433,In_2067,In_516);
and U2434 (N_2434,In_1796,In_371);
or U2435 (N_2435,In_108,In_1946);
and U2436 (N_2436,In_2138,In_2042);
nand U2437 (N_2437,In_986,In_2132);
nand U2438 (N_2438,In_369,In_232);
or U2439 (N_2439,In_731,In_2428);
nor U2440 (N_2440,In_149,In_667);
xnor U2441 (N_2441,In_2348,In_2266);
and U2442 (N_2442,In_1388,In_869);
and U2443 (N_2443,In_1547,In_281);
or U2444 (N_2444,In_883,In_1452);
nor U2445 (N_2445,In_2055,In_1224);
nand U2446 (N_2446,In_1121,In_1867);
nor U2447 (N_2447,In_114,In_450);
nand U2448 (N_2448,In_724,In_871);
nand U2449 (N_2449,In_810,In_273);
xor U2450 (N_2450,In_2039,In_2219);
xnor U2451 (N_2451,In_2468,In_958);
nand U2452 (N_2452,In_2413,In_756);
xnor U2453 (N_2453,In_1300,In_1915);
or U2454 (N_2454,In_163,In_2279);
and U2455 (N_2455,In_358,In_296);
nor U2456 (N_2456,In_119,In_807);
and U2457 (N_2457,In_182,In_721);
or U2458 (N_2458,In_2189,In_1149);
and U2459 (N_2459,In_361,In_415);
nor U2460 (N_2460,In_1598,In_323);
and U2461 (N_2461,In_2303,In_2066);
nand U2462 (N_2462,In_439,In_91);
and U2463 (N_2463,In_753,In_2477);
xnor U2464 (N_2464,In_918,In_497);
xor U2465 (N_2465,In_820,In_2020);
nand U2466 (N_2466,In_886,In_1509);
xnor U2467 (N_2467,In_1126,In_918);
nor U2468 (N_2468,In_1760,In_867);
or U2469 (N_2469,In_744,In_2345);
nand U2470 (N_2470,In_335,In_2473);
nand U2471 (N_2471,In_1337,In_489);
and U2472 (N_2472,In_2178,In_602);
nand U2473 (N_2473,In_1544,In_111);
or U2474 (N_2474,In_430,In_709);
nor U2475 (N_2475,In_1362,In_108);
nand U2476 (N_2476,In_1891,In_589);
or U2477 (N_2477,In_766,In_101);
nor U2478 (N_2478,In_40,In_1105);
nand U2479 (N_2479,In_831,In_2425);
or U2480 (N_2480,In_2411,In_1259);
nand U2481 (N_2481,In_2091,In_1637);
or U2482 (N_2482,In_983,In_840);
nand U2483 (N_2483,In_1641,In_1548);
nor U2484 (N_2484,In_110,In_949);
nor U2485 (N_2485,In_2186,In_1072);
and U2486 (N_2486,In_406,In_60);
nand U2487 (N_2487,In_1913,In_585);
and U2488 (N_2488,In_661,In_1941);
or U2489 (N_2489,In_543,In_1168);
xnor U2490 (N_2490,In_2184,In_692);
nand U2491 (N_2491,In_1774,In_652);
and U2492 (N_2492,In_942,In_1667);
nand U2493 (N_2493,In_1032,In_1627);
and U2494 (N_2494,In_1852,In_1819);
nand U2495 (N_2495,In_1211,In_1831);
xor U2496 (N_2496,In_750,In_805);
or U2497 (N_2497,In_1181,In_2475);
nor U2498 (N_2498,In_1280,In_117);
or U2499 (N_2499,In_2183,In_776);
nor U2500 (N_2500,In_1802,In_453);
or U2501 (N_2501,In_768,In_1338);
or U2502 (N_2502,In_2181,In_710);
xnor U2503 (N_2503,In_2115,In_506);
and U2504 (N_2504,In_943,In_1376);
or U2505 (N_2505,In_2080,In_161);
and U2506 (N_2506,In_2009,In_617);
nand U2507 (N_2507,In_1056,In_1818);
and U2508 (N_2508,In_2294,In_1474);
nor U2509 (N_2509,In_883,In_619);
xnor U2510 (N_2510,In_40,In_2298);
nor U2511 (N_2511,In_89,In_789);
and U2512 (N_2512,In_646,In_624);
xnor U2513 (N_2513,In_642,In_535);
nand U2514 (N_2514,In_1963,In_1033);
and U2515 (N_2515,In_2227,In_1452);
xor U2516 (N_2516,In_1455,In_276);
or U2517 (N_2517,In_1955,In_710);
or U2518 (N_2518,In_159,In_245);
nor U2519 (N_2519,In_1358,In_331);
or U2520 (N_2520,In_1495,In_2350);
and U2521 (N_2521,In_2006,In_22);
and U2522 (N_2522,In_2016,In_527);
or U2523 (N_2523,In_624,In_1727);
or U2524 (N_2524,In_539,In_2392);
xor U2525 (N_2525,In_1393,In_1022);
or U2526 (N_2526,In_2450,In_767);
xnor U2527 (N_2527,In_1990,In_1995);
nand U2528 (N_2528,In_1600,In_2249);
xor U2529 (N_2529,In_607,In_1934);
and U2530 (N_2530,In_2400,In_405);
nor U2531 (N_2531,In_2242,In_1753);
nor U2532 (N_2532,In_1987,In_1526);
nand U2533 (N_2533,In_2162,In_1043);
and U2534 (N_2534,In_2379,In_56);
or U2535 (N_2535,In_691,In_528);
or U2536 (N_2536,In_770,In_2470);
nor U2537 (N_2537,In_2369,In_2193);
or U2538 (N_2538,In_201,In_921);
nand U2539 (N_2539,In_2107,In_307);
and U2540 (N_2540,In_1106,In_1524);
or U2541 (N_2541,In_2491,In_1759);
nand U2542 (N_2542,In_1516,In_1822);
and U2543 (N_2543,In_668,In_1108);
nand U2544 (N_2544,In_56,In_1857);
xnor U2545 (N_2545,In_412,In_1286);
and U2546 (N_2546,In_62,In_1134);
or U2547 (N_2547,In_1292,In_1178);
or U2548 (N_2548,In_2494,In_2495);
or U2549 (N_2549,In_2331,In_2148);
and U2550 (N_2550,In_117,In_1781);
nand U2551 (N_2551,In_1527,In_313);
and U2552 (N_2552,In_2027,In_1901);
nand U2553 (N_2553,In_218,In_2033);
xnor U2554 (N_2554,In_1160,In_1564);
nor U2555 (N_2555,In_51,In_259);
xnor U2556 (N_2556,In_1586,In_538);
nand U2557 (N_2557,In_1951,In_1727);
nand U2558 (N_2558,In_7,In_278);
nand U2559 (N_2559,In_1528,In_417);
or U2560 (N_2560,In_2084,In_1206);
xor U2561 (N_2561,In_561,In_1150);
nand U2562 (N_2562,In_291,In_2009);
or U2563 (N_2563,In_249,In_83);
or U2564 (N_2564,In_1266,In_2289);
nor U2565 (N_2565,In_438,In_1353);
or U2566 (N_2566,In_1550,In_2118);
and U2567 (N_2567,In_1562,In_745);
nand U2568 (N_2568,In_606,In_1321);
or U2569 (N_2569,In_361,In_1597);
nand U2570 (N_2570,In_397,In_533);
xor U2571 (N_2571,In_423,In_77);
or U2572 (N_2572,In_1753,In_580);
nor U2573 (N_2573,In_2050,In_1727);
and U2574 (N_2574,In_435,In_1061);
or U2575 (N_2575,In_1866,In_627);
nor U2576 (N_2576,In_2213,In_1882);
and U2577 (N_2577,In_367,In_1900);
nor U2578 (N_2578,In_2009,In_503);
nor U2579 (N_2579,In_2365,In_773);
and U2580 (N_2580,In_93,In_2147);
nand U2581 (N_2581,In_1963,In_640);
nor U2582 (N_2582,In_191,In_66);
nor U2583 (N_2583,In_1573,In_809);
or U2584 (N_2584,In_10,In_2316);
nand U2585 (N_2585,In_1520,In_2300);
xnor U2586 (N_2586,In_831,In_390);
and U2587 (N_2587,In_1676,In_1054);
nand U2588 (N_2588,In_2302,In_2406);
nor U2589 (N_2589,In_438,In_2231);
nand U2590 (N_2590,In_2289,In_1209);
or U2591 (N_2591,In_1688,In_1468);
xor U2592 (N_2592,In_710,In_906);
and U2593 (N_2593,In_633,In_2162);
or U2594 (N_2594,In_1778,In_2431);
xor U2595 (N_2595,In_1922,In_791);
xor U2596 (N_2596,In_1004,In_1050);
xnor U2597 (N_2597,In_1230,In_81);
xnor U2598 (N_2598,In_864,In_2477);
or U2599 (N_2599,In_429,In_2305);
nor U2600 (N_2600,In_236,In_2278);
nor U2601 (N_2601,In_1184,In_811);
nor U2602 (N_2602,In_1709,In_2056);
nand U2603 (N_2603,In_1367,In_1657);
and U2604 (N_2604,In_771,In_1510);
xor U2605 (N_2605,In_2333,In_2118);
nor U2606 (N_2606,In_2320,In_440);
and U2607 (N_2607,In_607,In_1333);
and U2608 (N_2608,In_1085,In_2241);
nand U2609 (N_2609,In_1243,In_1274);
and U2610 (N_2610,In_1249,In_286);
and U2611 (N_2611,In_1060,In_1033);
xnor U2612 (N_2612,In_2277,In_2366);
nand U2613 (N_2613,In_590,In_1860);
nand U2614 (N_2614,In_964,In_2017);
xnor U2615 (N_2615,In_5,In_838);
nand U2616 (N_2616,In_1607,In_2437);
xor U2617 (N_2617,In_2151,In_2372);
nand U2618 (N_2618,In_1896,In_432);
nor U2619 (N_2619,In_1156,In_1288);
nor U2620 (N_2620,In_283,In_2146);
and U2621 (N_2621,In_1341,In_27);
or U2622 (N_2622,In_1227,In_1773);
xnor U2623 (N_2623,In_1573,In_1129);
and U2624 (N_2624,In_525,In_1201);
xnor U2625 (N_2625,In_1511,In_82);
xnor U2626 (N_2626,In_169,In_326);
nand U2627 (N_2627,In_1713,In_2286);
and U2628 (N_2628,In_2377,In_1291);
nand U2629 (N_2629,In_1531,In_528);
xnor U2630 (N_2630,In_1755,In_2275);
or U2631 (N_2631,In_2200,In_1619);
nor U2632 (N_2632,In_1885,In_2322);
nor U2633 (N_2633,In_695,In_2292);
or U2634 (N_2634,In_597,In_986);
xnor U2635 (N_2635,In_1909,In_2158);
nor U2636 (N_2636,In_1444,In_1455);
nor U2637 (N_2637,In_1818,In_2365);
nor U2638 (N_2638,In_1633,In_2409);
and U2639 (N_2639,In_1926,In_1022);
or U2640 (N_2640,In_518,In_1279);
xor U2641 (N_2641,In_1703,In_1286);
and U2642 (N_2642,In_2251,In_2480);
xnor U2643 (N_2643,In_196,In_1735);
xor U2644 (N_2644,In_985,In_244);
nor U2645 (N_2645,In_2460,In_2421);
nor U2646 (N_2646,In_629,In_2059);
and U2647 (N_2647,In_1763,In_1722);
and U2648 (N_2648,In_83,In_753);
and U2649 (N_2649,In_1071,In_1565);
nor U2650 (N_2650,In_2369,In_1322);
and U2651 (N_2651,In_1577,In_833);
nand U2652 (N_2652,In_1310,In_471);
and U2653 (N_2653,In_316,In_1854);
and U2654 (N_2654,In_1832,In_1393);
or U2655 (N_2655,In_1544,In_1079);
xnor U2656 (N_2656,In_2064,In_1878);
or U2657 (N_2657,In_937,In_1275);
xor U2658 (N_2658,In_950,In_134);
nor U2659 (N_2659,In_19,In_2365);
and U2660 (N_2660,In_1781,In_1428);
nor U2661 (N_2661,In_1728,In_870);
or U2662 (N_2662,In_1432,In_1562);
nor U2663 (N_2663,In_420,In_1231);
nor U2664 (N_2664,In_1392,In_1292);
nand U2665 (N_2665,In_1970,In_2105);
xor U2666 (N_2666,In_31,In_900);
nand U2667 (N_2667,In_1031,In_1470);
xnor U2668 (N_2668,In_1039,In_832);
or U2669 (N_2669,In_144,In_2436);
and U2670 (N_2670,In_1467,In_2167);
nand U2671 (N_2671,In_2106,In_2081);
and U2672 (N_2672,In_1726,In_1768);
or U2673 (N_2673,In_871,In_1664);
or U2674 (N_2674,In_540,In_1560);
nand U2675 (N_2675,In_98,In_567);
or U2676 (N_2676,In_2369,In_2462);
or U2677 (N_2677,In_1347,In_2314);
and U2678 (N_2678,In_470,In_2215);
or U2679 (N_2679,In_157,In_1835);
or U2680 (N_2680,In_776,In_262);
and U2681 (N_2681,In_513,In_969);
or U2682 (N_2682,In_2436,In_2060);
and U2683 (N_2683,In_643,In_1332);
or U2684 (N_2684,In_1431,In_512);
xor U2685 (N_2685,In_807,In_346);
and U2686 (N_2686,In_2010,In_110);
or U2687 (N_2687,In_1470,In_188);
and U2688 (N_2688,In_1145,In_102);
or U2689 (N_2689,In_2148,In_78);
or U2690 (N_2690,In_2496,In_928);
or U2691 (N_2691,In_2459,In_564);
nor U2692 (N_2692,In_2216,In_72);
nor U2693 (N_2693,In_1184,In_882);
or U2694 (N_2694,In_1761,In_2182);
and U2695 (N_2695,In_1351,In_703);
xnor U2696 (N_2696,In_240,In_1238);
or U2697 (N_2697,In_562,In_1456);
xor U2698 (N_2698,In_1121,In_1688);
nor U2699 (N_2699,In_452,In_2003);
nor U2700 (N_2700,In_458,In_560);
xor U2701 (N_2701,In_1349,In_236);
or U2702 (N_2702,In_817,In_2396);
nor U2703 (N_2703,In_1479,In_1628);
nor U2704 (N_2704,In_1635,In_1199);
nand U2705 (N_2705,In_1136,In_112);
and U2706 (N_2706,In_2282,In_454);
and U2707 (N_2707,In_1918,In_267);
xnor U2708 (N_2708,In_1556,In_1216);
xor U2709 (N_2709,In_2467,In_1283);
nand U2710 (N_2710,In_1019,In_2143);
or U2711 (N_2711,In_2401,In_669);
nor U2712 (N_2712,In_1679,In_1642);
nand U2713 (N_2713,In_431,In_1215);
or U2714 (N_2714,In_110,In_548);
and U2715 (N_2715,In_223,In_2084);
and U2716 (N_2716,In_1374,In_513);
nand U2717 (N_2717,In_767,In_1416);
and U2718 (N_2718,In_238,In_1380);
or U2719 (N_2719,In_412,In_165);
and U2720 (N_2720,In_958,In_1251);
or U2721 (N_2721,In_1914,In_2288);
and U2722 (N_2722,In_406,In_1306);
xor U2723 (N_2723,In_2403,In_1031);
nor U2724 (N_2724,In_1816,In_1018);
and U2725 (N_2725,In_596,In_1081);
or U2726 (N_2726,In_556,In_711);
and U2727 (N_2727,In_37,In_649);
xnor U2728 (N_2728,In_1083,In_2257);
and U2729 (N_2729,In_784,In_207);
xnor U2730 (N_2730,In_635,In_1406);
nand U2731 (N_2731,In_1867,In_2131);
nor U2732 (N_2732,In_997,In_753);
nor U2733 (N_2733,In_326,In_721);
nand U2734 (N_2734,In_32,In_1853);
or U2735 (N_2735,In_1577,In_2291);
nand U2736 (N_2736,In_619,In_2241);
nor U2737 (N_2737,In_315,In_2218);
xnor U2738 (N_2738,In_768,In_1512);
and U2739 (N_2739,In_1350,In_31);
and U2740 (N_2740,In_401,In_821);
and U2741 (N_2741,In_1137,In_133);
and U2742 (N_2742,In_717,In_1130);
nand U2743 (N_2743,In_957,In_2261);
xnor U2744 (N_2744,In_1524,In_307);
nand U2745 (N_2745,In_1676,In_868);
xor U2746 (N_2746,In_155,In_2338);
or U2747 (N_2747,In_471,In_2450);
xor U2748 (N_2748,In_2492,In_739);
or U2749 (N_2749,In_1735,In_956);
nor U2750 (N_2750,In_883,In_1998);
nand U2751 (N_2751,In_1291,In_856);
nand U2752 (N_2752,In_460,In_51);
or U2753 (N_2753,In_83,In_1109);
and U2754 (N_2754,In_795,In_1748);
and U2755 (N_2755,In_885,In_2309);
and U2756 (N_2756,In_781,In_2075);
nor U2757 (N_2757,In_108,In_938);
nand U2758 (N_2758,In_645,In_121);
or U2759 (N_2759,In_932,In_1586);
xor U2760 (N_2760,In_686,In_955);
or U2761 (N_2761,In_2096,In_780);
nor U2762 (N_2762,In_1904,In_390);
nand U2763 (N_2763,In_2349,In_1281);
or U2764 (N_2764,In_1377,In_126);
nand U2765 (N_2765,In_1459,In_1496);
nand U2766 (N_2766,In_1466,In_2063);
nand U2767 (N_2767,In_1769,In_1399);
and U2768 (N_2768,In_1622,In_800);
and U2769 (N_2769,In_32,In_513);
and U2770 (N_2770,In_620,In_2085);
and U2771 (N_2771,In_991,In_175);
nand U2772 (N_2772,In_1861,In_1976);
xor U2773 (N_2773,In_1122,In_2119);
or U2774 (N_2774,In_897,In_142);
and U2775 (N_2775,In_719,In_357);
nand U2776 (N_2776,In_1560,In_362);
and U2777 (N_2777,In_2437,In_2244);
nand U2778 (N_2778,In_1908,In_2489);
and U2779 (N_2779,In_779,In_589);
xor U2780 (N_2780,In_1329,In_1556);
nand U2781 (N_2781,In_1797,In_878);
nor U2782 (N_2782,In_845,In_66);
or U2783 (N_2783,In_1078,In_402);
xnor U2784 (N_2784,In_1814,In_2455);
nand U2785 (N_2785,In_842,In_420);
or U2786 (N_2786,In_83,In_1862);
nand U2787 (N_2787,In_248,In_1675);
xnor U2788 (N_2788,In_1682,In_1875);
nand U2789 (N_2789,In_2389,In_2083);
xor U2790 (N_2790,In_1368,In_2228);
or U2791 (N_2791,In_1266,In_323);
and U2792 (N_2792,In_373,In_2391);
nand U2793 (N_2793,In_398,In_2189);
nand U2794 (N_2794,In_755,In_1843);
or U2795 (N_2795,In_899,In_976);
nor U2796 (N_2796,In_325,In_886);
xor U2797 (N_2797,In_960,In_2401);
nand U2798 (N_2798,In_627,In_834);
nand U2799 (N_2799,In_1503,In_2295);
nor U2800 (N_2800,In_1854,In_2136);
nor U2801 (N_2801,In_1031,In_1646);
xnor U2802 (N_2802,In_2435,In_414);
xor U2803 (N_2803,In_1120,In_120);
nand U2804 (N_2804,In_653,In_2411);
and U2805 (N_2805,In_1288,In_794);
or U2806 (N_2806,In_832,In_2000);
and U2807 (N_2807,In_680,In_428);
xor U2808 (N_2808,In_1743,In_1400);
nor U2809 (N_2809,In_788,In_1371);
xor U2810 (N_2810,In_781,In_1271);
or U2811 (N_2811,In_1163,In_650);
and U2812 (N_2812,In_348,In_1008);
nor U2813 (N_2813,In_366,In_1924);
xor U2814 (N_2814,In_1,In_1080);
nor U2815 (N_2815,In_2424,In_699);
nand U2816 (N_2816,In_378,In_2139);
nand U2817 (N_2817,In_1624,In_2372);
or U2818 (N_2818,In_801,In_2116);
nand U2819 (N_2819,In_1454,In_735);
nand U2820 (N_2820,In_1758,In_1533);
nand U2821 (N_2821,In_1006,In_2456);
nor U2822 (N_2822,In_281,In_2354);
nor U2823 (N_2823,In_2183,In_2337);
and U2824 (N_2824,In_114,In_891);
nand U2825 (N_2825,In_1107,In_22);
or U2826 (N_2826,In_1985,In_2099);
nand U2827 (N_2827,In_135,In_1226);
or U2828 (N_2828,In_2090,In_1557);
nand U2829 (N_2829,In_979,In_1481);
and U2830 (N_2830,In_2243,In_113);
or U2831 (N_2831,In_1603,In_1068);
or U2832 (N_2832,In_539,In_2460);
nand U2833 (N_2833,In_315,In_1772);
nor U2834 (N_2834,In_1634,In_2495);
nand U2835 (N_2835,In_2388,In_1640);
or U2836 (N_2836,In_1769,In_1441);
and U2837 (N_2837,In_151,In_2048);
nor U2838 (N_2838,In_584,In_1540);
xor U2839 (N_2839,In_1384,In_9);
or U2840 (N_2840,In_2203,In_2413);
nor U2841 (N_2841,In_632,In_1043);
and U2842 (N_2842,In_1523,In_394);
xnor U2843 (N_2843,In_552,In_382);
or U2844 (N_2844,In_304,In_1953);
xor U2845 (N_2845,In_1702,In_1816);
xnor U2846 (N_2846,In_584,In_2412);
nand U2847 (N_2847,In_1957,In_1340);
nand U2848 (N_2848,In_1967,In_1367);
nand U2849 (N_2849,In_259,In_2200);
and U2850 (N_2850,In_2344,In_351);
xor U2851 (N_2851,In_1168,In_1124);
nor U2852 (N_2852,In_2367,In_1165);
xnor U2853 (N_2853,In_1695,In_530);
or U2854 (N_2854,In_201,In_1577);
and U2855 (N_2855,In_1599,In_1061);
nand U2856 (N_2856,In_1745,In_1059);
or U2857 (N_2857,In_2396,In_1062);
nor U2858 (N_2858,In_2459,In_1277);
nand U2859 (N_2859,In_344,In_998);
nor U2860 (N_2860,In_756,In_910);
nand U2861 (N_2861,In_2031,In_268);
nor U2862 (N_2862,In_2419,In_471);
xor U2863 (N_2863,In_1380,In_2259);
nand U2864 (N_2864,In_1753,In_1974);
or U2865 (N_2865,In_1377,In_1031);
xor U2866 (N_2866,In_2100,In_1125);
and U2867 (N_2867,In_1562,In_133);
nor U2868 (N_2868,In_1542,In_527);
nand U2869 (N_2869,In_881,In_1865);
nand U2870 (N_2870,In_1817,In_1884);
nand U2871 (N_2871,In_652,In_1904);
and U2872 (N_2872,In_1790,In_569);
and U2873 (N_2873,In_1749,In_1797);
xnor U2874 (N_2874,In_2230,In_116);
nand U2875 (N_2875,In_179,In_1424);
xnor U2876 (N_2876,In_2107,In_2083);
or U2877 (N_2877,In_935,In_1714);
nor U2878 (N_2878,In_397,In_1877);
or U2879 (N_2879,In_2031,In_474);
nand U2880 (N_2880,In_734,In_74);
or U2881 (N_2881,In_1527,In_698);
or U2882 (N_2882,In_1498,In_1282);
and U2883 (N_2883,In_300,In_1678);
and U2884 (N_2884,In_2195,In_1413);
or U2885 (N_2885,In_391,In_1134);
or U2886 (N_2886,In_1797,In_2413);
or U2887 (N_2887,In_287,In_417);
xor U2888 (N_2888,In_809,In_1154);
and U2889 (N_2889,In_672,In_1958);
nand U2890 (N_2890,In_983,In_1457);
xnor U2891 (N_2891,In_1350,In_476);
nand U2892 (N_2892,In_734,In_1058);
xnor U2893 (N_2893,In_163,In_363);
nor U2894 (N_2894,In_178,In_1863);
nor U2895 (N_2895,In_1084,In_1441);
nand U2896 (N_2896,In_2440,In_1826);
xnor U2897 (N_2897,In_1482,In_2416);
nor U2898 (N_2898,In_1839,In_673);
xnor U2899 (N_2899,In_2315,In_1296);
nand U2900 (N_2900,In_1232,In_1986);
and U2901 (N_2901,In_566,In_2262);
and U2902 (N_2902,In_2006,In_2189);
nor U2903 (N_2903,In_1400,In_210);
nand U2904 (N_2904,In_0,In_2050);
or U2905 (N_2905,In_1788,In_2107);
or U2906 (N_2906,In_2220,In_255);
xor U2907 (N_2907,In_2332,In_485);
nand U2908 (N_2908,In_1308,In_120);
xnor U2909 (N_2909,In_618,In_1067);
and U2910 (N_2910,In_1200,In_2129);
xor U2911 (N_2911,In_1374,In_1395);
nor U2912 (N_2912,In_704,In_2109);
or U2913 (N_2913,In_1535,In_1662);
nor U2914 (N_2914,In_1797,In_622);
xnor U2915 (N_2915,In_2403,In_2049);
nor U2916 (N_2916,In_1939,In_255);
or U2917 (N_2917,In_9,In_1498);
nand U2918 (N_2918,In_940,In_2380);
xnor U2919 (N_2919,In_2,In_1405);
and U2920 (N_2920,In_1252,In_364);
or U2921 (N_2921,In_2047,In_571);
nand U2922 (N_2922,In_1346,In_2028);
and U2923 (N_2923,In_1657,In_219);
nand U2924 (N_2924,In_1326,In_2144);
xor U2925 (N_2925,In_961,In_2447);
nand U2926 (N_2926,In_1926,In_1316);
xnor U2927 (N_2927,In_652,In_735);
nand U2928 (N_2928,In_270,In_934);
nor U2929 (N_2929,In_1416,In_1395);
nor U2930 (N_2930,In_2057,In_623);
or U2931 (N_2931,In_1406,In_1885);
nand U2932 (N_2932,In_2299,In_1226);
xor U2933 (N_2933,In_607,In_2386);
xor U2934 (N_2934,In_1830,In_431);
or U2935 (N_2935,In_1890,In_1772);
and U2936 (N_2936,In_549,In_890);
nor U2937 (N_2937,In_1140,In_367);
or U2938 (N_2938,In_288,In_129);
and U2939 (N_2939,In_176,In_1434);
nand U2940 (N_2940,In_1200,In_1779);
xor U2941 (N_2941,In_145,In_558);
xor U2942 (N_2942,In_365,In_348);
xor U2943 (N_2943,In_876,In_2201);
or U2944 (N_2944,In_1767,In_895);
or U2945 (N_2945,In_772,In_867);
xnor U2946 (N_2946,In_1221,In_1722);
nor U2947 (N_2947,In_1950,In_723);
nand U2948 (N_2948,In_95,In_538);
nor U2949 (N_2949,In_941,In_351);
or U2950 (N_2950,In_1326,In_44);
nand U2951 (N_2951,In_2316,In_1118);
and U2952 (N_2952,In_1103,In_1483);
or U2953 (N_2953,In_1733,In_1669);
xor U2954 (N_2954,In_308,In_2233);
nand U2955 (N_2955,In_1614,In_689);
xnor U2956 (N_2956,In_57,In_1871);
nor U2957 (N_2957,In_1807,In_833);
xor U2958 (N_2958,In_1912,In_1619);
nand U2959 (N_2959,In_281,In_1264);
or U2960 (N_2960,In_712,In_1044);
and U2961 (N_2961,In_964,In_2022);
and U2962 (N_2962,In_1191,In_219);
and U2963 (N_2963,In_652,In_214);
or U2964 (N_2964,In_1431,In_1718);
or U2965 (N_2965,In_959,In_1140);
nor U2966 (N_2966,In_1865,In_54);
xnor U2967 (N_2967,In_14,In_206);
xor U2968 (N_2968,In_328,In_1244);
nand U2969 (N_2969,In_1354,In_127);
xnor U2970 (N_2970,In_268,In_2064);
or U2971 (N_2971,In_167,In_601);
xor U2972 (N_2972,In_1457,In_641);
and U2973 (N_2973,In_1005,In_1666);
or U2974 (N_2974,In_1095,In_2173);
and U2975 (N_2975,In_1813,In_229);
xnor U2976 (N_2976,In_839,In_1938);
nor U2977 (N_2977,In_779,In_1226);
xor U2978 (N_2978,In_354,In_276);
or U2979 (N_2979,In_1193,In_1900);
and U2980 (N_2980,In_1115,In_910);
or U2981 (N_2981,In_1555,In_1330);
nand U2982 (N_2982,In_460,In_2330);
and U2983 (N_2983,In_486,In_1893);
and U2984 (N_2984,In_1644,In_2079);
nand U2985 (N_2985,In_1892,In_1733);
nand U2986 (N_2986,In_749,In_2247);
xor U2987 (N_2987,In_1382,In_2205);
and U2988 (N_2988,In_1955,In_1858);
nand U2989 (N_2989,In_2248,In_380);
xor U2990 (N_2990,In_1489,In_923);
and U2991 (N_2991,In_1916,In_806);
nor U2992 (N_2992,In_771,In_2119);
and U2993 (N_2993,In_1917,In_464);
or U2994 (N_2994,In_1680,In_1491);
and U2995 (N_2995,In_2187,In_153);
and U2996 (N_2996,In_98,In_1956);
xor U2997 (N_2997,In_2007,In_2318);
and U2998 (N_2998,In_224,In_1106);
xnor U2999 (N_2999,In_1718,In_313);
or U3000 (N_3000,In_650,In_2122);
xnor U3001 (N_3001,In_1238,In_311);
nand U3002 (N_3002,In_1147,In_2141);
and U3003 (N_3003,In_1458,In_940);
nor U3004 (N_3004,In_936,In_1120);
nand U3005 (N_3005,In_836,In_2016);
and U3006 (N_3006,In_115,In_302);
nand U3007 (N_3007,In_2444,In_955);
xor U3008 (N_3008,In_1536,In_1310);
and U3009 (N_3009,In_733,In_1320);
and U3010 (N_3010,In_1496,In_408);
and U3011 (N_3011,In_634,In_1811);
and U3012 (N_3012,In_1871,In_487);
and U3013 (N_3013,In_2222,In_1272);
xor U3014 (N_3014,In_1652,In_1236);
nor U3015 (N_3015,In_1042,In_1212);
nand U3016 (N_3016,In_293,In_624);
xnor U3017 (N_3017,In_2436,In_2491);
nand U3018 (N_3018,In_2095,In_669);
or U3019 (N_3019,In_1111,In_1681);
and U3020 (N_3020,In_740,In_93);
nand U3021 (N_3021,In_57,In_1059);
and U3022 (N_3022,In_1593,In_502);
or U3023 (N_3023,In_1087,In_1144);
nand U3024 (N_3024,In_654,In_561);
xnor U3025 (N_3025,In_1155,In_1441);
or U3026 (N_3026,In_1342,In_491);
and U3027 (N_3027,In_1821,In_1020);
or U3028 (N_3028,In_1552,In_493);
and U3029 (N_3029,In_799,In_2017);
and U3030 (N_3030,In_665,In_1769);
nor U3031 (N_3031,In_886,In_2168);
xor U3032 (N_3032,In_1588,In_1472);
nand U3033 (N_3033,In_536,In_1804);
nand U3034 (N_3034,In_2399,In_448);
and U3035 (N_3035,In_55,In_1597);
or U3036 (N_3036,In_1332,In_607);
xor U3037 (N_3037,In_1936,In_1959);
xnor U3038 (N_3038,In_705,In_1627);
and U3039 (N_3039,In_1627,In_1642);
nand U3040 (N_3040,In_465,In_1562);
or U3041 (N_3041,In_1373,In_1954);
and U3042 (N_3042,In_1125,In_1391);
nor U3043 (N_3043,In_2337,In_1994);
nand U3044 (N_3044,In_548,In_2145);
nand U3045 (N_3045,In_361,In_2109);
and U3046 (N_3046,In_229,In_1073);
xor U3047 (N_3047,In_278,In_1895);
nor U3048 (N_3048,In_696,In_512);
or U3049 (N_3049,In_1417,In_1736);
or U3050 (N_3050,In_2081,In_216);
nand U3051 (N_3051,In_1682,In_69);
and U3052 (N_3052,In_1973,In_1611);
nor U3053 (N_3053,In_538,In_603);
xnor U3054 (N_3054,In_1946,In_741);
and U3055 (N_3055,In_1276,In_1700);
and U3056 (N_3056,In_1146,In_1561);
or U3057 (N_3057,In_2056,In_1012);
xnor U3058 (N_3058,In_1051,In_1117);
or U3059 (N_3059,In_415,In_126);
nor U3060 (N_3060,In_849,In_715);
or U3061 (N_3061,In_2166,In_463);
or U3062 (N_3062,In_1243,In_899);
or U3063 (N_3063,In_1623,In_1795);
nor U3064 (N_3064,In_1053,In_772);
nand U3065 (N_3065,In_2419,In_1502);
nor U3066 (N_3066,In_1381,In_1426);
nand U3067 (N_3067,In_801,In_2199);
nor U3068 (N_3068,In_2150,In_973);
nor U3069 (N_3069,In_894,In_672);
nor U3070 (N_3070,In_305,In_527);
nor U3071 (N_3071,In_99,In_973);
xor U3072 (N_3072,In_2086,In_2123);
and U3073 (N_3073,In_1913,In_1015);
or U3074 (N_3074,In_1843,In_1002);
nand U3075 (N_3075,In_334,In_1072);
nand U3076 (N_3076,In_911,In_1758);
xor U3077 (N_3077,In_731,In_1002);
xor U3078 (N_3078,In_91,In_522);
or U3079 (N_3079,In_2033,In_357);
and U3080 (N_3080,In_1231,In_2018);
nor U3081 (N_3081,In_2138,In_2415);
nand U3082 (N_3082,In_2256,In_726);
or U3083 (N_3083,In_1292,In_1232);
nor U3084 (N_3084,In_1799,In_1271);
nor U3085 (N_3085,In_2089,In_2285);
or U3086 (N_3086,In_2339,In_1691);
and U3087 (N_3087,In_745,In_1685);
or U3088 (N_3088,In_868,In_2341);
or U3089 (N_3089,In_445,In_1084);
xnor U3090 (N_3090,In_777,In_1219);
xnor U3091 (N_3091,In_1495,In_2109);
nor U3092 (N_3092,In_1603,In_1713);
nor U3093 (N_3093,In_4,In_368);
or U3094 (N_3094,In_817,In_812);
or U3095 (N_3095,In_1228,In_46);
or U3096 (N_3096,In_1398,In_169);
xnor U3097 (N_3097,In_455,In_1422);
or U3098 (N_3098,In_2313,In_521);
and U3099 (N_3099,In_569,In_420);
and U3100 (N_3100,In_155,In_797);
nor U3101 (N_3101,In_1454,In_819);
xnor U3102 (N_3102,In_1447,In_1529);
nor U3103 (N_3103,In_1043,In_1285);
xnor U3104 (N_3104,In_1016,In_2059);
nand U3105 (N_3105,In_918,In_21);
nor U3106 (N_3106,In_2060,In_1910);
and U3107 (N_3107,In_1348,In_1911);
and U3108 (N_3108,In_1564,In_2421);
or U3109 (N_3109,In_2452,In_2027);
xor U3110 (N_3110,In_580,In_263);
nand U3111 (N_3111,In_1440,In_2172);
nor U3112 (N_3112,In_172,In_540);
xnor U3113 (N_3113,In_198,In_71);
xnor U3114 (N_3114,In_1553,In_1265);
or U3115 (N_3115,In_418,In_834);
nand U3116 (N_3116,In_1017,In_364);
and U3117 (N_3117,In_2104,In_1452);
and U3118 (N_3118,In_1622,In_2484);
or U3119 (N_3119,In_2434,In_1820);
nor U3120 (N_3120,In_330,In_1430);
xnor U3121 (N_3121,In_16,In_550);
and U3122 (N_3122,In_2352,In_1344);
nand U3123 (N_3123,In_2115,In_1391);
xnor U3124 (N_3124,In_2423,In_1587);
and U3125 (N_3125,In_337,In_606);
nor U3126 (N_3126,In_2305,In_395);
or U3127 (N_3127,In_2162,In_235);
and U3128 (N_3128,In_2497,In_100);
and U3129 (N_3129,In_1371,In_629);
nor U3130 (N_3130,In_2372,In_720);
and U3131 (N_3131,In_1917,In_835);
nand U3132 (N_3132,In_1537,In_1184);
nand U3133 (N_3133,In_1409,In_1815);
nand U3134 (N_3134,In_608,In_2418);
xor U3135 (N_3135,In_2110,In_2277);
nor U3136 (N_3136,In_31,In_1637);
or U3137 (N_3137,In_164,In_591);
xor U3138 (N_3138,In_1734,In_888);
xor U3139 (N_3139,In_2177,In_43);
or U3140 (N_3140,In_712,In_1173);
and U3141 (N_3141,In_1194,In_1623);
nand U3142 (N_3142,In_313,In_1673);
or U3143 (N_3143,In_174,In_813);
nor U3144 (N_3144,In_1877,In_453);
or U3145 (N_3145,In_165,In_1024);
xnor U3146 (N_3146,In_2147,In_940);
and U3147 (N_3147,In_1666,In_656);
and U3148 (N_3148,In_486,In_511);
xor U3149 (N_3149,In_860,In_1162);
or U3150 (N_3150,In_1572,In_752);
or U3151 (N_3151,In_1228,In_2250);
or U3152 (N_3152,In_986,In_1363);
or U3153 (N_3153,In_2233,In_1634);
or U3154 (N_3154,In_829,In_344);
xnor U3155 (N_3155,In_2409,In_1317);
and U3156 (N_3156,In_275,In_2045);
nor U3157 (N_3157,In_2296,In_199);
xor U3158 (N_3158,In_358,In_1113);
nor U3159 (N_3159,In_2097,In_1907);
xor U3160 (N_3160,In_754,In_698);
or U3161 (N_3161,In_1662,In_1749);
nand U3162 (N_3162,In_1541,In_1613);
nand U3163 (N_3163,In_2101,In_1946);
or U3164 (N_3164,In_1434,In_149);
and U3165 (N_3165,In_1127,In_227);
and U3166 (N_3166,In_48,In_516);
and U3167 (N_3167,In_1369,In_1545);
nor U3168 (N_3168,In_1479,In_1544);
nand U3169 (N_3169,In_533,In_10);
nand U3170 (N_3170,In_244,In_1238);
nor U3171 (N_3171,In_1973,In_2304);
and U3172 (N_3172,In_1916,In_1516);
nor U3173 (N_3173,In_1180,In_1197);
nand U3174 (N_3174,In_2002,In_684);
nor U3175 (N_3175,In_1342,In_2103);
or U3176 (N_3176,In_1797,In_2071);
nor U3177 (N_3177,In_815,In_2453);
nor U3178 (N_3178,In_1428,In_1659);
nand U3179 (N_3179,In_431,In_1435);
nand U3180 (N_3180,In_970,In_1262);
nand U3181 (N_3181,In_1160,In_1039);
xor U3182 (N_3182,In_929,In_377);
and U3183 (N_3183,In_1206,In_226);
xor U3184 (N_3184,In_1051,In_1687);
nor U3185 (N_3185,In_1931,In_67);
nand U3186 (N_3186,In_511,In_675);
nand U3187 (N_3187,In_772,In_559);
nor U3188 (N_3188,In_298,In_1625);
and U3189 (N_3189,In_412,In_1355);
nand U3190 (N_3190,In_856,In_1735);
and U3191 (N_3191,In_654,In_1921);
xor U3192 (N_3192,In_1418,In_2460);
nand U3193 (N_3193,In_2112,In_1740);
and U3194 (N_3194,In_1245,In_1995);
and U3195 (N_3195,In_2141,In_718);
xor U3196 (N_3196,In_1010,In_579);
and U3197 (N_3197,In_1516,In_1121);
nor U3198 (N_3198,In_1873,In_2104);
xnor U3199 (N_3199,In_2136,In_826);
xnor U3200 (N_3200,In_1123,In_2100);
and U3201 (N_3201,In_713,In_1478);
nand U3202 (N_3202,In_1024,In_594);
nor U3203 (N_3203,In_957,In_1180);
or U3204 (N_3204,In_1725,In_954);
or U3205 (N_3205,In_2104,In_356);
and U3206 (N_3206,In_1025,In_866);
or U3207 (N_3207,In_6,In_2498);
nand U3208 (N_3208,In_2126,In_1207);
xnor U3209 (N_3209,In_1745,In_160);
nor U3210 (N_3210,In_694,In_894);
nand U3211 (N_3211,In_2017,In_80);
and U3212 (N_3212,In_970,In_2001);
nor U3213 (N_3213,In_1839,In_2307);
xnor U3214 (N_3214,In_2147,In_435);
xnor U3215 (N_3215,In_388,In_1773);
or U3216 (N_3216,In_2,In_865);
or U3217 (N_3217,In_893,In_2496);
nand U3218 (N_3218,In_922,In_1977);
or U3219 (N_3219,In_543,In_2163);
nor U3220 (N_3220,In_1278,In_190);
nand U3221 (N_3221,In_252,In_577);
and U3222 (N_3222,In_768,In_366);
or U3223 (N_3223,In_227,In_2150);
xnor U3224 (N_3224,In_1923,In_1019);
nand U3225 (N_3225,In_2188,In_251);
nand U3226 (N_3226,In_2014,In_234);
and U3227 (N_3227,In_930,In_1246);
xnor U3228 (N_3228,In_525,In_1296);
nand U3229 (N_3229,In_816,In_64);
or U3230 (N_3230,In_1673,In_677);
nand U3231 (N_3231,In_2249,In_1688);
and U3232 (N_3232,In_2146,In_2329);
and U3233 (N_3233,In_1394,In_1352);
and U3234 (N_3234,In_737,In_162);
or U3235 (N_3235,In_2346,In_585);
nand U3236 (N_3236,In_1876,In_2022);
xor U3237 (N_3237,In_2181,In_311);
and U3238 (N_3238,In_1507,In_1861);
or U3239 (N_3239,In_167,In_13);
nor U3240 (N_3240,In_144,In_1387);
nand U3241 (N_3241,In_1994,In_1760);
nor U3242 (N_3242,In_772,In_1656);
and U3243 (N_3243,In_144,In_578);
xnor U3244 (N_3244,In_1194,In_2169);
or U3245 (N_3245,In_720,In_1813);
nand U3246 (N_3246,In_759,In_1021);
nand U3247 (N_3247,In_1174,In_1138);
nor U3248 (N_3248,In_1494,In_827);
nand U3249 (N_3249,In_912,In_1748);
or U3250 (N_3250,In_1548,In_443);
and U3251 (N_3251,In_1759,In_2281);
or U3252 (N_3252,In_199,In_781);
nand U3253 (N_3253,In_2306,In_1851);
nand U3254 (N_3254,In_1456,In_1416);
nand U3255 (N_3255,In_71,In_557);
nor U3256 (N_3256,In_887,In_395);
nand U3257 (N_3257,In_625,In_1134);
or U3258 (N_3258,In_925,In_1161);
and U3259 (N_3259,In_2285,In_2481);
and U3260 (N_3260,In_1489,In_378);
and U3261 (N_3261,In_1203,In_1345);
nand U3262 (N_3262,In_2244,In_2084);
nor U3263 (N_3263,In_1369,In_1011);
and U3264 (N_3264,In_1435,In_708);
xor U3265 (N_3265,In_2134,In_2086);
and U3266 (N_3266,In_937,In_1750);
nor U3267 (N_3267,In_1315,In_1528);
and U3268 (N_3268,In_2027,In_1839);
nor U3269 (N_3269,In_1545,In_575);
or U3270 (N_3270,In_1215,In_1810);
or U3271 (N_3271,In_116,In_649);
xnor U3272 (N_3272,In_982,In_1902);
and U3273 (N_3273,In_38,In_185);
nand U3274 (N_3274,In_2417,In_1891);
nand U3275 (N_3275,In_773,In_1816);
xnor U3276 (N_3276,In_1031,In_1034);
nor U3277 (N_3277,In_911,In_1419);
xor U3278 (N_3278,In_1575,In_2191);
or U3279 (N_3279,In_1802,In_1052);
and U3280 (N_3280,In_2124,In_205);
xnor U3281 (N_3281,In_1067,In_897);
and U3282 (N_3282,In_561,In_1421);
nand U3283 (N_3283,In_1324,In_1453);
and U3284 (N_3284,In_392,In_1713);
xor U3285 (N_3285,In_1546,In_1556);
or U3286 (N_3286,In_117,In_600);
or U3287 (N_3287,In_1132,In_1392);
nor U3288 (N_3288,In_2240,In_2449);
xor U3289 (N_3289,In_321,In_137);
nor U3290 (N_3290,In_1816,In_2361);
or U3291 (N_3291,In_127,In_2374);
or U3292 (N_3292,In_1161,In_112);
nand U3293 (N_3293,In_1696,In_1);
xnor U3294 (N_3294,In_667,In_2159);
nor U3295 (N_3295,In_1681,In_804);
and U3296 (N_3296,In_792,In_177);
and U3297 (N_3297,In_562,In_1321);
or U3298 (N_3298,In_321,In_647);
and U3299 (N_3299,In_1349,In_96);
and U3300 (N_3300,In_1990,In_1538);
nand U3301 (N_3301,In_1992,In_172);
and U3302 (N_3302,In_1061,In_757);
xnor U3303 (N_3303,In_807,In_1737);
and U3304 (N_3304,In_2491,In_1507);
nand U3305 (N_3305,In_1990,In_2180);
xnor U3306 (N_3306,In_2311,In_631);
or U3307 (N_3307,In_226,In_385);
nand U3308 (N_3308,In_749,In_2120);
xnor U3309 (N_3309,In_1581,In_600);
nor U3310 (N_3310,In_2154,In_883);
nor U3311 (N_3311,In_1455,In_367);
nand U3312 (N_3312,In_1076,In_2146);
or U3313 (N_3313,In_1412,In_2258);
nand U3314 (N_3314,In_420,In_1202);
or U3315 (N_3315,In_1849,In_1034);
and U3316 (N_3316,In_529,In_1227);
nand U3317 (N_3317,In_719,In_118);
nor U3318 (N_3318,In_1661,In_1018);
nand U3319 (N_3319,In_235,In_1264);
xnor U3320 (N_3320,In_1549,In_1506);
or U3321 (N_3321,In_658,In_1185);
xor U3322 (N_3322,In_119,In_1994);
nor U3323 (N_3323,In_498,In_512);
or U3324 (N_3324,In_527,In_2358);
or U3325 (N_3325,In_1063,In_1597);
or U3326 (N_3326,In_1570,In_1149);
nor U3327 (N_3327,In_563,In_727);
nor U3328 (N_3328,In_351,In_764);
xor U3329 (N_3329,In_1442,In_2119);
nand U3330 (N_3330,In_589,In_1453);
nor U3331 (N_3331,In_321,In_1761);
xor U3332 (N_3332,In_1354,In_2289);
nand U3333 (N_3333,In_601,In_2276);
xor U3334 (N_3334,In_214,In_1900);
xor U3335 (N_3335,In_1380,In_1452);
and U3336 (N_3336,In_2274,In_1689);
nor U3337 (N_3337,In_2465,In_910);
nor U3338 (N_3338,In_897,In_1162);
nand U3339 (N_3339,In_2205,In_573);
or U3340 (N_3340,In_1331,In_2413);
xnor U3341 (N_3341,In_587,In_2036);
nor U3342 (N_3342,In_2022,In_561);
nand U3343 (N_3343,In_356,In_2384);
xnor U3344 (N_3344,In_174,In_1698);
or U3345 (N_3345,In_821,In_957);
or U3346 (N_3346,In_1872,In_71);
or U3347 (N_3347,In_1331,In_2255);
nand U3348 (N_3348,In_1709,In_1797);
and U3349 (N_3349,In_655,In_1983);
or U3350 (N_3350,In_2470,In_1287);
nor U3351 (N_3351,In_846,In_620);
or U3352 (N_3352,In_1168,In_1907);
xnor U3353 (N_3353,In_187,In_1798);
xor U3354 (N_3354,In_2182,In_2295);
or U3355 (N_3355,In_2195,In_1898);
xor U3356 (N_3356,In_1929,In_1948);
nor U3357 (N_3357,In_753,In_1341);
nand U3358 (N_3358,In_521,In_595);
or U3359 (N_3359,In_795,In_579);
xor U3360 (N_3360,In_1508,In_454);
nor U3361 (N_3361,In_1404,In_1976);
or U3362 (N_3362,In_2303,In_1295);
and U3363 (N_3363,In_1033,In_1808);
nor U3364 (N_3364,In_1336,In_759);
or U3365 (N_3365,In_698,In_2472);
or U3366 (N_3366,In_1821,In_283);
xnor U3367 (N_3367,In_1396,In_942);
nand U3368 (N_3368,In_1035,In_2485);
nand U3369 (N_3369,In_2402,In_455);
nand U3370 (N_3370,In_202,In_180);
or U3371 (N_3371,In_2305,In_1237);
nor U3372 (N_3372,In_1510,In_1593);
nor U3373 (N_3373,In_1792,In_1857);
and U3374 (N_3374,In_1039,In_1471);
and U3375 (N_3375,In_1815,In_213);
nand U3376 (N_3376,In_2046,In_860);
xnor U3377 (N_3377,In_629,In_339);
xnor U3378 (N_3378,In_2127,In_2174);
nor U3379 (N_3379,In_32,In_510);
and U3380 (N_3380,In_1974,In_1429);
or U3381 (N_3381,In_2376,In_64);
and U3382 (N_3382,In_1633,In_2124);
or U3383 (N_3383,In_755,In_1868);
and U3384 (N_3384,In_109,In_927);
xor U3385 (N_3385,In_1537,In_1036);
nand U3386 (N_3386,In_1991,In_1858);
nand U3387 (N_3387,In_1938,In_720);
nand U3388 (N_3388,In_474,In_2149);
nor U3389 (N_3389,In_1109,In_2202);
or U3390 (N_3390,In_1692,In_2483);
nand U3391 (N_3391,In_402,In_2059);
nand U3392 (N_3392,In_932,In_550);
nand U3393 (N_3393,In_1157,In_382);
nand U3394 (N_3394,In_1803,In_1828);
and U3395 (N_3395,In_1474,In_1972);
or U3396 (N_3396,In_917,In_1246);
xnor U3397 (N_3397,In_1911,In_100);
or U3398 (N_3398,In_1632,In_1182);
and U3399 (N_3399,In_1516,In_2269);
xor U3400 (N_3400,In_702,In_1260);
xnor U3401 (N_3401,In_726,In_531);
nand U3402 (N_3402,In_687,In_752);
nor U3403 (N_3403,In_350,In_2220);
nor U3404 (N_3404,In_1094,In_2331);
xor U3405 (N_3405,In_1150,In_2465);
nand U3406 (N_3406,In_2284,In_530);
and U3407 (N_3407,In_98,In_938);
and U3408 (N_3408,In_1160,In_2437);
xnor U3409 (N_3409,In_764,In_103);
or U3410 (N_3410,In_538,In_206);
nor U3411 (N_3411,In_1539,In_1188);
or U3412 (N_3412,In_1820,In_5);
nand U3413 (N_3413,In_1132,In_2256);
and U3414 (N_3414,In_626,In_1428);
and U3415 (N_3415,In_1232,In_2009);
or U3416 (N_3416,In_841,In_1510);
xnor U3417 (N_3417,In_1814,In_1666);
nor U3418 (N_3418,In_2181,In_1500);
nand U3419 (N_3419,In_2160,In_357);
xnor U3420 (N_3420,In_2062,In_1458);
and U3421 (N_3421,In_1762,In_1853);
xnor U3422 (N_3422,In_968,In_1626);
and U3423 (N_3423,In_2455,In_1058);
and U3424 (N_3424,In_1432,In_1469);
nand U3425 (N_3425,In_121,In_1144);
xor U3426 (N_3426,In_1794,In_1561);
or U3427 (N_3427,In_2212,In_374);
or U3428 (N_3428,In_784,In_268);
xor U3429 (N_3429,In_1787,In_1322);
and U3430 (N_3430,In_1380,In_2219);
nand U3431 (N_3431,In_2025,In_1953);
nor U3432 (N_3432,In_564,In_1569);
xnor U3433 (N_3433,In_1042,In_22);
nand U3434 (N_3434,In_1022,In_2275);
nor U3435 (N_3435,In_738,In_1589);
or U3436 (N_3436,In_1739,In_2145);
or U3437 (N_3437,In_1504,In_1023);
nand U3438 (N_3438,In_2478,In_222);
and U3439 (N_3439,In_1759,In_1737);
nor U3440 (N_3440,In_5,In_1037);
nand U3441 (N_3441,In_2339,In_768);
nand U3442 (N_3442,In_2486,In_2321);
nor U3443 (N_3443,In_952,In_2470);
or U3444 (N_3444,In_529,In_1165);
xnor U3445 (N_3445,In_1005,In_360);
and U3446 (N_3446,In_1567,In_2021);
nand U3447 (N_3447,In_1404,In_992);
nor U3448 (N_3448,In_377,In_1821);
nand U3449 (N_3449,In_78,In_1705);
nor U3450 (N_3450,In_345,In_2411);
nand U3451 (N_3451,In_2093,In_2442);
or U3452 (N_3452,In_1659,In_579);
and U3453 (N_3453,In_350,In_1632);
xor U3454 (N_3454,In_1303,In_148);
or U3455 (N_3455,In_2480,In_1392);
nand U3456 (N_3456,In_356,In_1342);
nor U3457 (N_3457,In_1794,In_805);
and U3458 (N_3458,In_1025,In_411);
and U3459 (N_3459,In_1459,In_1527);
nor U3460 (N_3460,In_618,In_2184);
and U3461 (N_3461,In_159,In_670);
xnor U3462 (N_3462,In_2372,In_2306);
and U3463 (N_3463,In_1936,In_1543);
and U3464 (N_3464,In_611,In_2410);
or U3465 (N_3465,In_901,In_663);
nor U3466 (N_3466,In_30,In_1355);
and U3467 (N_3467,In_1785,In_1464);
nor U3468 (N_3468,In_117,In_1076);
nor U3469 (N_3469,In_1765,In_857);
nand U3470 (N_3470,In_1875,In_1912);
nor U3471 (N_3471,In_1462,In_1880);
nor U3472 (N_3472,In_2117,In_774);
and U3473 (N_3473,In_1860,In_1258);
nand U3474 (N_3474,In_1793,In_780);
nor U3475 (N_3475,In_1475,In_1588);
nor U3476 (N_3476,In_508,In_839);
nor U3477 (N_3477,In_855,In_2417);
and U3478 (N_3478,In_2432,In_1844);
nor U3479 (N_3479,In_1779,In_2126);
and U3480 (N_3480,In_2442,In_2241);
nor U3481 (N_3481,In_1160,In_1715);
and U3482 (N_3482,In_1535,In_2128);
and U3483 (N_3483,In_2421,In_962);
xnor U3484 (N_3484,In_94,In_1945);
or U3485 (N_3485,In_1458,In_542);
nor U3486 (N_3486,In_1863,In_1015);
nand U3487 (N_3487,In_938,In_2348);
nor U3488 (N_3488,In_1647,In_1213);
or U3489 (N_3489,In_2100,In_2432);
or U3490 (N_3490,In_2118,In_2279);
or U3491 (N_3491,In_1372,In_526);
nor U3492 (N_3492,In_1996,In_597);
or U3493 (N_3493,In_509,In_1494);
nor U3494 (N_3494,In_2011,In_707);
nand U3495 (N_3495,In_426,In_1957);
nand U3496 (N_3496,In_899,In_1678);
nand U3497 (N_3497,In_1490,In_2097);
or U3498 (N_3498,In_698,In_499);
xor U3499 (N_3499,In_2249,In_1987);
xor U3500 (N_3500,In_832,In_688);
or U3501 (N_3501,In_2486,In_1455);
and U3502 (N_3502,In_1582,In_569);
nor U3503 (N_3503,In_1399,In_1527);
or U3504 (N_3504,In_1906,In_1565);
xnor U3505 (N_3505,In_332,In_786);
and U3506 (N_3506,In_1606,In_1138);
xnor U3507 (N_3507,In_998,In_1854);
nor U3508 (N_3508,In_186,In_732);
nand U3509 (N_3509,In_2303,In_2220);
nor U3510 (N_3510,In_2061,In_1246);
nor U3511 (N_3511,In_505,In_813);
xnor U3512 (N_3512,In_2323,In_1707);
and U3513 (N_3513,In_1026,In_2128);
or U3514 (N_3514,In_2353,In_2274);
nor U3515 (N_3515,In_2318,In_1067);
and U3516 (N_3516,In_1297,In_1625);
nand U3517 (N_3517,In_1866,In_282);
xor U3518 (N_3518,In_304,In_807);
nor U3519 (N_3519,In_1644,In_1346);
nand U3520 (N_3520,In_177,In_123);
or U3521 (N_3521,In_2439,In_2070);
and U3522 (N_3522,In_586,In_1434);
and U3523 (N_3523,In_1342,In_1732);
or U3524 (N_3524,In_916,In_752);
nor U3525 (N_3525,In_249,In_46);
and U3526 (N_3526,In_1149,In_1720);
nor U3527 (N_3527,In_77,In_501);
nand U3528 (N_3528,In_956,In_1450);
nor U3529 (N_3529,In_770,In_1836);
xnor U3530 (N_3530,In_635,In_1957);
nand U3531 (N_3531,In_33,In_297);
nor U3532 (N_3532,In_331,In_1537);
nor U3533 (N_3533,In_1035,In_167);
xor U3534 (N_3534,In_950,In_386);
and U3535 (N_3535,In_2483,In_1605);
and U3536 (N_3536,In_2293,In_4);
and U3537 (N_3537,In_2435,In_410);
nor U3538 (N_3538,In_449,In_1954);
or U3539 (N_3539,In_222,In_2345);
and U3540 (N_3540,In_2203,In_25);
nand U3541 (N_3541,In_726,In_1841);
nor U3542 (N_3542,In_1249,In_2065);
or U3543 (N_3543,In_319,In_1292);
nor U3544 (N_3544,In_1365,In_68);
xor U3545 (N_3545,In_2198,In_2027);
nand U3546 (N_3546,In_1758,In_190);
or U3547 (N_3547,In_2338,In_1128);
nand U3548 (N_3548,In_1246,In_1927);
or U3549 (N_3549,In_2439,In_2152);
nor U3550 (N_3550,In_2438,In_754);
nor U3551 (N_3551,In_1576,In_753);
and U3552 (N_3552,In_234,In_2060);
nand U3553 (N_3553,In_931,In_1819);
xor U3554 (N_3554,In_433,In_180);
nand U3555 (N_3555,In_1513,In_1194);
nand U3556 (N_3556,In_206,In_2355);
nand U3557 (N_3557,In_2165,In_143);
and U3558 (N_3558,In_2474,In_424);
or U3559 (N_3559,In_256,In_2143);
nand U3560 (N_3560,In_75,In_764);
or U3561 (N_3561,In_1589,In_2462);
and U3562 (N_3562,In_340,In_2439);
or U3563 (N_3563,In_1711,In_1938);
nor U3564 (N_3564,In_1541,In_1273);
xnor U3565 (N_3565,In_1696,In_287);
nand U3566 (N_3566,In_177,In_1881);
nor U3567 (N_3567,In_1761,In_784);
or U3568 (N_3568,In_470,In_2268);
nor U3569 (N_3569,In_214,In_519);
nor U3570 (N_3570,In_657,In_1782);
and U3571 (N_3571,In_1504,In_2406);
and U3572 (N_3572,In_1814,In_385);
nand U3573 (N_3573,In_87,In_209);
nand U3574 (N_3574,In_2052,In_2365);
nor U3575 (N_3575,In_232,In_355);
and U3576 (N_3576,In_2453,In_1131);
xor U3577 (N_3577,In_723,In_2209);
nor U3578 (N_3578,In_3,In_1587);
nand U3579 (N_3579,In_441,In_2499);
nand U3580 (N_3580,In_1038,In_1160);
or U3581 (N_3581,In_1794,In_2130);
xnor U3582 (N_3582,In_1486,In_728);
nand U3583 (N_3583,In_2035,In_1652);
nand U3584 (N_3584,In_429,In_1918);
xor U3585 (N_3585,In_962,In_1223);
nand U3586 (N_3586,In_1462,In_1124);
nor U3587 (N_3587,In_1860,In_1666);
nand U3588 (N_3588,In_1141,In_2172);
nor U3589 (N_3589,In_1005,In_1958);
and U3590 (N_3590,In_1430,In_1852);
nor U3591 (N_3591,In_1052,In_371);
xnor U3592 (N_3592,In_1691,In_845);
xnor U3593 (N_3593,In_1697,In_33);
nand U3594 (N_3594,In_2428,In_1901);
and U3595 (N_3595,In_2442,In_2355);
nand U3596 (N_3596,In_875,In_454);
nand U3597 (N_3597,In_1045,In_2246);
and U3598 (N_3598,In_429,In_443);
and U3599 (N_3599,In_1005,In_1233);
nor U3600 (N_3600,In_2087,In_2121);
nor U3601 (N_3601,In_1092,In_1355);
nor U3602 (N_3602,In_2331,In_1012);
and U3603 (N_3603,In_401,In_423);
or U3604 (N_3604,In_2345,In_1562);
nand U3605 (N_3605,In_669,In_523);
nand U3606 (N_3606,In_2411,In_1933);
and U3607 (N_3607,In_1635,In_1145);
or U3608 (N_3608,In_632,In_1167);
nand U3609 (N_3609,In_1995,In_2152);
nand U3610 (N_3610,In_1322,In_477);
xor U3611 (N_3611,In_196,In_1626);
nand U3612 (N_3612,In_2301,In_999);
nor U3613 (N_3613,In_1032,In_1368);
xor U3614 (N_3614,In_1077,In_1043);
nand U3615 (N_3615,In_393,In_438);
xnor U3616 (N_3616,In_519,In_1620);
xnor U3617 (N_3617,In_1693,In_433);
xnor U3618 (N_3618,In_1142,In_1482);
nor U3619 (N_3619,In_408,In_2068);
or U3620 (N_3620,In_748,In_989);
xor U3621 (N_3621,In_1990,In_381);
or U3622 (N_3622,In_1585,In_1446);
and U3623 (N_3623,In_1986,In_1673);
and U3624 (N_3624,In_853,In_2477);
nor U3625 (N_3625,In_990,In_1822);
and U3626 (N_3626,In_843,In_1686);
xnor U3627 (N_3627,In_1652,In_1059);
nor U3628 (N_3628,In_2231,In_1362);
nand U3629 (N_3629,In_2130,In_2171);
xor U3630 (N_3630,In_1226,In_1191);
and U3631 (N_3631,In_1687,In_1599);
nand U3632 (N_3632,In_642,In_1993);
nand U3633 (N_3633,In_476,In_247);
xor U3634 (N_3634,In_1003,In_2286);
nand U3635 (N_3635,In_1436,In_2074);
nand U3636 (N_3636,In_1466,In_443);
nand U3637 (N_3637,In_962,In_120);
and U3638 (N_3638,In_608,In_112);
nor U3639 (N_3639,In_2456,In_1952);
or U3640 (N_3640,In_46,In_586);
nor U3641 (N_3641,In_1414,In_2487);
xor U3642 (N_3642,In_733,In_1656);
xor U3643 (N_3643,In_447,In_1004);
xnor U3644 (N_3644,In_557,In_1375);
and U3645 (N_3645,In_1900,In_1057);
nor U3646 (N_3646,In_2244,In_1510);
and U3647 (N_3647,In_441,In_637);
nand U3648 (N_3648,In_473,In_892);
and U3649 (N_3649,In_1541,In_1925);
and U3650 (N_3650,In_1949,In_144);
or U3651 (N_3651,In_2190,In_2425);
and U3652 (N_3652,In_544,In_135);
nor U3653 (N_3653,In_2304,In_2137);
nand U3654 (N_3654,In_1400,In_2027);
xnor U3655 (N_3655,In_1267,In_2407);
nand U3656 (N_3656,In_1400,In_1675);
and U3657 (N_3657,In_990,In_1859);
and U3658 (N_3658,In_942,In_334);
or U3659 (N_3659,In_846,In_810);
xnor U3660 (N_3660,In_1907,In_194);
or U3661 (N_3661,In_161,In_218);
xnor U3662 (N_3662,In_1360,In_2296);
and U3663 (N_3663,In_602,In_1734);
xnor U3664 (N_3664,In_1283,In_591);
or U3665 (N_3665,In_1503,In_616);
nand U3666 (N_3666,In_1862,In_1334);
or U3667 (N_3667,In_755,In_2249);
nand U3668 (N_3668,In_18,In_963);
or U3669 (N_3669,In_1728,In_174);
and U3670 (N_3670,In_730,In_2269);
nor U3671 (N_3671,In_1896,In_251);
nor U3672 (N_3672,In_676,In_183);
xor U3673 (N_3673,In_446,In_771);
nor U3674 (N_3674,In_786,In_2484);
nand U3675 (N_3675,In_352,In_2489);
or U3676 (N_3676,In_1929,In_1153);
nand U3677 (N_3677,In_681,In_2239);
xnor U3678 (N_3678,In_1955,In_943);
nand U3679 (N_3679,In_1855,In_1866);
nor U3680 (N_3680,In_2498,In_839);
or U3681 (N_3681,In_215,In_468);
or U3682 (N_3682,In_1554,In_2406);
or U3683 (N_3683,In_119,In_623);
or U3684 (N_3684,In_327,In_102);
nor U3685 (N_3685,In_1245,In_1058);
xor U3686 (N_3686,In_460,In_1798);
nand U3687 (N_3687,In_488,In_1220);
nand U3688 (N_3688,In_577,In_1500);
xnor U3689 (N_3689,In_2176,In_757);
nor U3690 (N_3690,In_115,In_1118);
nand U3691 (N_3691,In_2126,In_235);
and U3692 (N_3692,In_273,In_2296);
nor U3693 (N_3693,In_1689,In_2309);
nand U3694 (N_3694,In_1845,In_35);
or U3695 (N_3695,In_1675,In_1808);
or U3696 (N_3696,In_1265,In_31);
nand U3697 (N_3697,In_1644,In_1278);
and U3698 (N_3698,In_52,In_2349);
or U3699 (N_3699,In_1073,In_1253);
nor U3700 (N_3700,In_1977,In_39);
nand U3701 (N_3701,In_1404,In_2472);
and U3702 (N_3702,In_1398,In_138);
or U3703 (N_3703,In_2480,In_1343);
nand U3704 (N_3704,In_526,In_1844);
or U3705 (N_3705,In_418,In_894);
xor U3706 (N_3706,In_817,In_1819);
nand U3707 (N_3707,In_1020,In_807);
nand U3708 (N_3708,In_332,In_1520);
xor U3709 (N_3709,In_846,In_1051);
or U3710 (N_3710,In_1202,In_1496);
and U3711 (N_3711,In_1813,In_56);
nor U3712 (N_3712,In_1815,In_420);
or U3713 (N_3713,In_983,In_219);
or U3714 (N_3714,In_940,In_1376);
xor U3715 (N_3715,In_43,In_1952);
or U3716 (N_3716,In_1177,In_1309);
xnor U3717 (N_3717,In_995,In_14);
nand U3718 (N_3718,In_1625,In_209);
and U3719 (N_3719,In_523,In_1506);
and U3720 (N_3720,In_1120,In_2022);
or U3721 (N_3721,In_1330,In_662);
or U3722 (N_3722,In_1230,In_1845);
xor U3723 (N_3723,In_498,In_490);
nand U3724 (N_3724,In_1833,In_1502);
or U3725 (N_3725,In_1812,In_303);
nor U3726 (N_3726,In_2418,In_171);
and U3727 (N_3727,In_1740,In_1363);
nand U3728 (N_3728,In_2399,In_1738);
xor U3729 (N_3729,In_1677,In_1808);
nand U3730 (N_3730,In_1013,In_987);
nor U3731 (N_3731,In_2316,In_2444);
xor U3732 (N_3732,In_1117,In_1659);
nor U3733 (N_3733,In_1015,In_749);
and U3734 (N_3734,In_677,In_2377);
xnor U3735 (N_3735,In_270,In_2308);
xor U3736 (N_3736,In_97,In_2110);
and U3737 (N_3737,In_1236,In_132);
xor U3738 (N_3738,In_462,In_583);
or U3739 (N_3739,In_1960,In_826);
and U3740 (N_3740,In_2258,In_1700);
nand U3741 (N_3741,In_481,In_2202);
xor U3742 (N_3742,In_1257,In_2180);
nand U3743 (N_3743,In_683,In_968);
xor U3744 (N_3744,In_1760,In_776);
or U3745 (N_3745,In_1441,In_1926);
nor U3746 (N_3746,In_797,In_392);
nand U3747 (N_3747,In_718,In_698);
nand U3748 (N_3748,In_2371,In_368);
xor U3749 (N_3749,In_705,In_1377);
or U3750 (N_3750,In_792,In_1122);
and U3751 (N_3751,In_1648,In_1637);
xnor U3752 (N_3752,In_970,In_214);
and U3753 (N_3753,In_1256,In_2194);
nor U3754 (N_3754,In_2045,In_130);
nand U3755 (N_3755,In_343,In_244);
nor U3756 (N_3756,In_1740,In_1357);
or U3757 (N_3757,In_2422,In_1505);
nor U3758 (N_3758,In_56,In_1811);
xor U3759 (N_3759,In_2453,In_1723);
and U3760 (N_3760,In_1236,In_1826);
and U3761 (N_3761,In_508,In_1686);
xnor U3762 (N_3762,In_1396,In_1483);
and U3763 (N_3763,In_812,In_1713);
or U3764 (N_3764,In_2207,In_1983);
nand U3765 (N_3765,In_153,In_2085);
nor U3766 (N_3766,In_2482,In_127);
and U3767 (N_3767,In_1304,In_1536);
nand U3768 (N_3768,In_754,In_2174);
nand U3769 (N_3769,In_156,In_1453);
nor U3770 (N_3770,In_889,In_1526);
xnor U3771 (N_3771,In_818,In_561);
xnor U3772 (N_3772,In_2433,In_2239);
xor U3773 (N_3773,In_308,In_2438);
nand U3774 (N_3774,In_2125,In_603);
xnor U3775 (N_3775,In_1716,In_533);
and U3776 (N_3776,In_1190,In_861);
and U3777 (N_3777,In_2294,In_2307);
and U3778 (N_3778,In_1161,In_123);
nor U3779 (N_3779,In_2382,In_1898);
xor U3780 (N_3780,In_858,In_1311);
nand U3781 (N_3781,In_209,In_1496);
nor U3782 (N_3782,In_1400,In_402);
or U3783 (N_3783,In_526,In_161);
nor U3784 (N_3784,In_1923,In_1268);
and U3785 (N_3785,In_552,In_1155);
and U3786 (N_3786,In_142,In_1166);
nor U3787 (N_3787,In_2415,In_1766);
xnor U3788 (N_3788,In_2037,In_1472);
nor U3789 (N_3789,In_347,In_700);
nand U3790 (N_3790,In_201,In_174);
nor U3791 (N_3791,In_1465,In_168);
nand U3792 (N_3792,In_1408,In_1448);
xor U3793 (N_3793,In_1206,In_1299);
xnor U3794 (N_3794,In_2321,In_2172);
nor U3795 (N_3795,In_1235,In_34);
nor U3796 (N_3796,In_2321,In_891);
or U3797 (N_3797,In_1486,In_1505);
nor U3798 (N_3798,In_92,In_82);
nor U3799 (N_3799,In_1839,In_1971);
and U3800 (N_3800,In_1446,In_201);
xor U3801 (N_3801,In_1970,In_943);
or U3802 (N_3802,In_2403,In_1703);
nor U3803 (N_3803,In_1279,In_1518);
and U3804 (N_3804,In_1265,In_257);
nor U3805 (N_3805,In_2473,In_539);
and U3806 (N_3806,In_1443,In_311);
or U3807 (N_3807,In_2035,In_1080);
nor U3808 (N_3808,In_759,In_2468);
nor U3809 (N_3809,In_2357,In_2179);
nor U3810 (N_3810,In_2232,In_1970);
and U3811 (N_3811,In_2150,In_1221);
and U3812 (N_3812,In_381,In_616);
and U3813 (N_3813,In_756,In_1298);
nand U3814 (N_3814,In_2064,In_1873);
or U3815 (N_3815,In_1640,In_2383);
and U3816 (N_3816,In_550,In_497);
or U3817 (N_3817,In_1525,In_2319);
and U3818 (N_3818,In_2306,In_1286);
and U3819 (N_3819,In_1288,In_1942);
and U3820 (N_3820,In_804,In_1438);
and U3821 (N_3821,In_985,In_182);
or U3822 (N_3822,In_1792,In_2325);
and U3823 (N_3823,In_2286,In_562);
nor U3824 (N_3824,In_1779,In_1086);
xor U3825 (N_3825,In_568,In_702);
nor U3826 (N_3826,In_1705,In_753);
and U3827 (N_3827,In_1795,In_1582);
or U3828 (N_3828,In_531,In_2483);
xor U3829 (N_3829,In_301,In_1335);
nor U3830 (N_3830,In_1881,In_416);
and U3831 (N_3831,In_823,In_722);
xor U3832 (N_3832,In_1162,In_1990);
nand U3833 (N_3833,In_1038,In_1667);
xnor U3834 (N_3834,In_619,In_2188);
nand U3835 (N_3835,In_2127,In_303);
nor U3836 (N_3836,In_1625,In_1486);
and U3837 (N_3837,In_114,In_1297);
or U3838 (N_3838,In_1905,In_2268);
nor U3839 (N_3839,In_1812,In_489);
xor U3840 (N_3840,In_398,In_1743);
or U3841 (N_3841,In_1479,In_2466);
nor U3842 (N_3842,In_1948,In_85);
xor U3843 (N_3843,In_1671,In_1820);
and U3844 (N_3844,In_286,In_1177);
and U3845 (N_3845,In_585,In_2371);
nor U3846 (N_3846,In_275,In_1303);
and U3847 (N_3847,In_1463,In_932);
and U3848 (N_3848,In_560,In_1463);
xor U3849 (N_3849,In_1170,In_2083);
nand U3850 (N_3850,In_2098,In_712);
nor U3851 (N_3851,In_2493,In_1833);
or U3852 (N_3852,In_1799,In_1759);
xor U3853 (N_3853,In_744,In_382);
nor U3854 (N_3854,In_1320,In_831);
or U3855 (N_3855,In_1840,In_451);
or U3856 (N_3856,In_981,In_1023);
or U3857 (N_3857,In_1956,In_633);
xnor U3858 (N_3858,In_940,In_1971);
and U3859 (N_3859,In_1381,In_1394);
xor U3860 (N_3860,In_1535,In_388);
xnor U3861 (N_3861,In_2035,In_2255);
xnor U3862 (N_3862,In_667,In_2061);
nand U3863 (N_3863,In_1313,In_1144);
or U3864 (N_3864,In_1952,In_878);
xnor U3865 (N_3865,In_1721,In_580);
nand U3866 (N_3866,In_1702,In_454);
or U3867 (N_3867,In_1527,In_1740);
or U3868 (N_3868,In_659,In_499);
and U3869 (N_3869,In_329,In_648);
xnor U3870 (N_3870,In_1491,In_638);
or U3871 (N_3871,In_1273,In_966);
xor U3872 (N_3872,In_848,In_763);
nor U3873 (N_3873,In_2366,In_1118);
nor U3874 (N_3874,In_1485,In_1249);
and U3875 (N_3875,In_2382,In_1374);
and U3876 (N_3876,In_515,In_2353);
nor U3877 (N_3877,In_489,In_1781);
nor U3878 (N_3878,In_1762,In_1959);
or U3879 (N_3879,In_538,In_1793);
nand U3880 (N_3880,In_73,In_991);
and U3881 (N_3881,In_1090,In_870);
nor U3882 (N_3882,In_2416,In_94);
nor U3883 (N_3883,In_1079,In_2197);
nand U3884 (N_3884,In_498,In_672);
xor U3885 (N_3885,In_262,In_70);
xnor U3886 (N_3886,In_1954,In_58);
xor U3887 (N_3887,In_199,In_589);
xnor U3888 (N_3888,In_1800,In_475);
nor U3889 (N_3889,In_1201,In_1705);
or U3890 (N_3890,In_2261,In_1611);
nor U3891 (N_3891,In_1915,In_901);
xnor U3892 (N_3892,In_316,In_1125);
and U3893 (N_3893,In_1358,In_2105);
nor U3894 (N_3894,In_665,In_806);
nand U3895 (N_3895,In_1688,In_676);
or U3896 (N_3896,In_1625,In_942);
nand U3897 (N_3897,In_1029,In_1533);
and U3898 (N_3898,In_225,In_615);
xnor U3899 (N_3899,In_2039,In_129);
nor U3900 (N_3900,In_1245,In_1106);
xnor U3901 (N_3901,In_1758,In_170);
xnor U3902 (N_3902,In_876,In_1669);
nor U3903 (N_3903,In_1802,In_1371);
nand U3904 (N_3904,In_2297,In_2359);
and U3905 (N_3905,In_2252,In_2448);
nand U3906 (N_3906,In_89,In_184);
nand U3907 (N_3907,In_1600,In_458);
xor U3908 (N_3908,In_1390,In_83);
and U3909 (N_3909,In_2221,In_888);
or U3910 (N_3910,In_2408,In_1176);
and U3911 (N_3911,In_834,In_1367);
xnor U3912 (N_3912,In_622,In_2467);
nor U3913 (N_3913,In_1627,In_75);
nor U3914 (N_3914,In_1227,In_380);
and U3915 (N_3915,In_800,In_73);
or U3916 (N_3916,In_67,In_165);
and U3917 (N_3917,In_205,In_2152);
and U3918 (N_3918,In_207,In_1381);
and U3919 (N_3919,In_1296,In_197);
nor U3920 (N_3920,In_554,In_298);
nor U3921 (N_3921,In_2192,In_129);
xor U3922 (N_3922,In_964,In_1486);
nand U3923 (N_3923,In_1684,In_1853);
xor U3924 (N_3924,In_1681,In_1488);
nor U3925 (N_3925,In_724,In_2202);
xor U3926 (N_3926,In_513,In_885);
nor U3927 (N_3927,In_696,In_1381);
nor U3928 (N_3928,In_439,In_1934);
xor U3929 (N_3929,In_1041,In_1226);
nor U3930 (N_3930,In_2460,In_2240);
nand U3931 (N_3931,In_1287,In_490);
xnor U3932 (N_3932,In_1940,In_2417);
and U3933 (N_3933,In_342,In_1835);
xnor U3934 (N_3934,In_2343,In_2272);
or U3935 (N_3935,In_1998,In_1116);
nand U3936 (N_3936,In_46,In_2);
nor U3937 (N_3937,In_775,In_347);
xnor U3938 (N_3938,In_639,In_2041);
nand U3939 (N_3939,In_2198,In_547);
or U3940 (N_3940,In_618,In_847);
and U3941 (N_3941,In_2313,In_118);
nor U3942 (N_3942,In_457,In_836);
and U3943 (N_3943,In_256,In_1377);
and U3944 (N_3944,In_1082,In_756);
or U3945 (N_3945,In_2436,In_546);
and U3946 (N_3946,In_1737,In_320);
or U3947 (N_3947,In_459,In_1665);
xor U3948 (N_3948,In_1905,In_1374);
nor U3949 (N_3949,In_539,In_430);
and U3950 (N_3950,In_1415,In_517);
nor U3951 (N_3951,In_2489,In_985);
nor U3952 (N_3952,In_2013,In_511);
or U3953 (N_3953,In_2106,In_678);
nand U3954 (N_3954,In_815,In_1017);
or U3955 (N_3955,In_796,In_2007);
and U3956 (N_3956,In_620,In_324);
xnor U3957 (N_3957,In_36,In_2163);
xor U3958 (N_3958,In_421,In_758);
nand U3959 (N_3959,In_2219,In_2285);
or U3960 (N_3960,In_1451,In_1603);
nor U3961 (N_3961,In_1809,In_855);
xnor U3962 (N_3962,In_1417,In_2004);
and U3963 (N_3963,In_1918,In_1626);
and U3964 (N_3964,In_1177,In_720);
nand U3965 (N_3965,In_2079,In_1454);
nor U3966 (N_3966,In_571,In_1589);
xor U3967 (N_3967,In_2003,In_1581);
nand U3968 (N_3968,In_1485,In_1595);
nand U3969 (N_3969,In_1959,In_216);
xnor U3970 (N_3970,In_1631,In_2061);
nand U3971 (N_3971,In_1867,In_664);
nand U3972 (N_3972,In_907,In_1770);
xnor U3973 (N_3973,In_2383,In_119);
xor U3974 (N_3974,In_1961,In_2377);
xor U3975 (N_3975,In_1015,In_1374);
xnor U3976 (N_3976,In_2477,In_2108);
and U3977 (N_3977,In_424,In_1268);
xnor U3978 (N_3978,In_1368,In_590);
nand U3979 (N_3979,In_421,In_2191);
nand U3980 (N_3980,In_1786,In_72);
xor U3981 (N_3981,In_1699,In_1918);
or U3982 (N_3982,In_1748,In_2145);
xor U3983 (N_3983,In_1265,In_1228);
nor U3984 (N_3984,In_40,In_1466);
xnor U3985 (N_3985,In_1614,In_118);
nand U3986 (N_3986,In_260,In_464);
and U3987 (N_3987,In_1830,In_1033);
nand U3988 (N_3988,In_2168,In_1269);
or U3989 (N_3989,In_640,In_202);
or U3990 (N_3990,In_1882,In_333);
or U3991 (N_3991,In_1533,In_1178);
and U3992 (N_3992,In_1249,In_814);
and U3993 (N_3993,In_1349,In_115);
or U3994 (N_3994,In_2095,In_1541);
xor U3995 (N_3995,In_1975,In_2126);
and U3996 (N_3996,In_1589,In_607);
xor U3997 (N_3997,In_984,In_802);
or U3998 (N_3998,In_1801,In_1903);
or U3999 (N_3999,In_568,In_971);
or U4000 (N_4000,In_1135,In_885);
nor U4001 (N_4001,In_402,In_2395);
xnor U4002 (N_4002,In_322,In_1931);
nand U4003 (N_4003,In_690,In_975);
or U4004 (N_4004,In_59,In_1772);
nand U4005 (N_4005,In_55,In_712);
nand U4006 (N_4006,In_515,In_933);
and U4007 (N_4007,In_178,In_285);
and U4008 (N_4008,In_268,In_2095);
or U4009 (N_4009,In_71,In_368);
and U4010 (N_4010,In_2493,In_648);
xnor U4011 (N_4011,In_50,In_97);
or U4012 (N_4012,In_1383,In_25);
or U4013 (N_4013,In_2350,In_2333);
nand U4014 (N_4014,In_66,In_1173);
nand U4015 (N_4015,In_93,In_2106);
nor U4016 (N_4016,In_42,In_2409);
nand U4017 (N_4017,In_1708,In_104);
or U4018 (N_4018,In_2094,In_1974);
xor U4019 (N_4019,In_2470,In_1036);
and U4020 (N_4020,In_1595,In_2278);
xnor U4021 (N_4021,In_1147,In_1351);
or U4022 (N_4022,In_1330,In_1297);
xor U4023 (N_4023,In_645,In_958);
nand U4024 (N_4024,In_186,In_2203);
nor U4025 (N_4025,In_674,In_1924);
nor U4026 (N_4026,In_2074,In_302);
and U4027 (N_4027,In_1176,In_1511);
nor U4028 (N_4028,In_1638,In_566);
xnor U4029 (N_4029,In_2032,In_2340);
and U4030 (N_4030,In_1796,In_2393);
or U4031 (N_4031,In_2084,In_1819);
or U4032 (N_4032,In_2255,In_846);
nor U4033 (N_4033,In_1680,In_2323);
nor U4034 (N_4034,In_1462,In_804);
and U4035 (N_4035,In_1052,In_1585);
nor U4036 (N_4036,In_1335,In_1005);
and U4037 (N_4037,In_1838,In_2389);
nand U4038 (N_4038,In_177,In_2229);
nor U4039 (N_4039,In_526,In_2029);
nand U4040 (N_4040,In_1975,In_127);
nand U4041 (N_4041,In_536,In_1826);
or U4042 (N_4042,In_564,In_1895);
and U4043 (N_4043,In_690,In_1476);
nor U4044 (N_4044,In_735,In_985);
xnor U4045 (N_4045,In_1479,In_2484);
xnor U4046 (N_4046,In_48,In_76);
or U4047 (N_4047,In_1326,In_1034);
xnor U4048 (N_4048,In_41,In_1315);
and U4049 (N_4049,In_1544,In_2267);
nor U4050 (N_4050,In_2247,In_721);
nand U4051 (N_4051,In_1750,In_1360);
xor U4052 (N_4052,In_753,In_2331);
nand U4053 (N_4053,In_682,In_719);
nand U4054 (N_4054,In_557,In_1097);
nor U4055 (N_4055,In_1005,In_826);
and U4056 (N_4056,In_2134,In_505);
xnor U4057 (N_4057,In_1708,In_180);
xor U4058 (N_4058,In_1119,In_975);
xnor U4059 (N_4059,In_918,In_993);
and U4060 (N_4060,In_581,In_1941);
xor U4061 (N_4061,In_2230,In_1019);
and U4062 (N_4062,In_2162,In_2165);
xor U4063 (N_4063,In_1772,In_1698);
nor U4064 (N_4064,In_1562,In_1012);
xnor U4065 (N_4065,In_1510,In_1925);
nand U4066 (N_4066,In_834,In_2044);
xnor U4067 (N_4067,In_2062,In_875);
or U4068 (N_4068,In_692,In_1295);
xnor U4069 (N_4069,In_1578,In_1507);
nand U4070 (N_4070,In_202,In_874);
xor U4071 (N_4071,In_302,In_1610);
or U4072 (N_4072,In_1735,In_743);
and U4073 (N_4073,In_733,In_721);
nor U4074 (N_4074,In_2229,In_724);
nand U4075 (N_4075,In_1178,In_35);
and U4076 (N_4076,In_2420,In_2168);
nor U4077 (N_4077,In_2447,In_1575);
or U4078 (N_4078,In_2000,In_2397);
nor U4079 (N_4079,In_1992,In_1416);
nor U4080 (N_4080,In_137,In_752);
nor U4081 (N_4081,In_172,In_1054);
or U4082 (N_4082,In_389,In_1934);
xor U4083 (N_4083,In_1195,In_70);
nor U4084 (N_4084,In_1772,In_241);
nor U4085 (N_4085,In_1556,In_1003);
nor U4086 (N_4086,In_1392,In_1653);
nand U4087 (N_4087,In_1913,In_2422);
nand U4088 (N_4088,In_1088,In_1585);
xor U4089 (N_4089,In_1976,In_713);
xor U4090 (N_4090,In_582,In_2442);
or U4091 (N_4091,In_2080,In_1946);
nor U4092 (N_4092,In_1455,In_874);
xnor U4093 (N_4093,In_630,In_1538);
nor U4094 (N_4094,In_1402,In_1079);
or U4095 (N_4095,In_508,In_218);
and U4096 (N_4096,In_2412,In_497);
and U4097 (N_4097,In_1389,In_886);
nor U4098 (N_4098,In_98,In_298);
and U4099 (N_4099,In_267,In_2224);
or U4100 (N_4100,In_1228,In_968);
nand U4101 (N_4101,In_1063,In_186);
and U4102 (N_4102,In_154,In_512);
nand U4103 (N_4103,In_595,In_1022);
or U4104 (N_4104,In_779,In_556);
and U4105 (N_4105,In_2083,In_416);
xnor U4106 (N_4106,In_2365,In_921);
nand U4107 (N_4107,In_361,In_247);
nand U4108 (N_4108,In_334,In_53);
xor U4109 (N_4109,In_1077,In_2172);
nand U4110 (N_4110,In_453,In_614);
and U4111 (N_4111,In_1038,In_564);
nand U4112 (N_4112,In_1434,In_175);
nand U4113 (N_4113,In_410,In_1329);
nor U4114 (N_4114,In_1618,In_1696);
nand U4115 (N_4115,In_2189,In_287);
or U4116 (N_4116,In_1208,In_143);
xor U4117 (N_4117,In_1814,In_398);
or U4118 (N_4118,In_2345,In_1896);
and U4119 (N_4119,In_2181,In_2459);
and U4120 (N_4120,In_1588,In_1956);
nor U4121 (N_4121,In_2391,In_1602);
and U4122 (N_4122,In_1423,In_2273);
xnor U4123 (N_4123,In_1168,In_2338);
xnor U4124 (N_4124,In_243,In_589);
xor U4125 (N_4125,In_600,In_1565);
and U4126 (N_4126,In_876,In_1973);
and U4127 (N_4127,In_1884,In_229);
nor U4128 (N_4128,In_2109,In_739);
xor U4129 (N_4129,In_1213,In_8);
nor U4130 (N_4130,In_1815,In_162);
or U4131 (N_4131,In_960,In_100);
xnor U4132 (N_4132,In_527,In_1177);
or U4133 (N_4133,In_132,In_821);
or U4134 (N_4134,In_23,In_1084);
xnor U4135 (N_4135,In_261,In_584);
and U4136 (N_4136,In_54,In_596);
nor U4137 (N_4137,In_436,In_136);
nand U4138 (N_4138,In_856,In_176);
and U4139 (N_4139,In_1110,In_1487);
nand U4140 (N_4140,In_1287,In_2473);
nand U4141 (N_4141,In_944,In_819);
nor U4142 (N_4142,In_278,In_2436);
nor U4143 (N_4143,In_1559,In_1169);
nor U4144 (N_4144,In_2133,In_2094);
and U4145 (N_4145,In_681,In_1645);
or U4146 (N_4146,In_1713,In_751);
and U4147 (N_4147,In_1479,In_321);
xor U4148 (N_4148,In_296,In_215);
nand U4149 (N_4149,In_1245,In_1505);
and U4150 (N_4150,In_1612,In_386);
nand U4151 (N_4151,In_1234,In_2279);
or U4152 (N_4152,In_658,In_2174);
nand U4153 (N_4153,In_875,In_1477);
nand U4154 (N_4154,In_2223,In_1171);
or U4155 (N_4155,In_1880,In_432);
nand U4156 (N_4156,In_663,In_249);
nor U4157 (N_4157,In_1370,In_2245);
nor U4158 (N_4158,In_2165,In_680);
nor U4159 (N_4159,In_1162,In_527);
or U4160 (N_4160,In_695,In_1509);
nand U4161 (N_4161,In_970,In_60);
or U4162 (N_4162,In_1167,In_974);
nor U4163 (N_4163,In_945,In_391);
nor U4164 (N_4164,In_1296,In_77);
nor U4165 (N_4165,In_1692,In_112);
and U4166 (N_4166,In_293,In_1570);
xnor U4167 (N_4167,In_2280,In_435);
xnor U4168 (N_4168,In_1261,In_1096);
xnor U4169 (N_4169,In_193,In_86);
nor U4170 (N_4170,In_828,In_743);
or U4171 (N_4171,In_2152,In_458);
or U4172 (N_4172,In_1903,In_724);
or U4173 (N_4173,In_659,In_379);
or U4174 (N_4174,In_690,In_1756);
nand U4175 (N_4175,In_1177,In_419);
nor U4176 (N_4176,In_1510,In_1644);
and U4177 (N_4177,In_2431,In_1248);
and U4178 (N_4178,In_2171,In_1788);
nor U4179 (N_4179,In_293,In_1979);
xor U4180 (N_4180,In_1756,In_708);
and U4181 (N_4181,In_2389,In_494);
and U4182 (N_4182,In_1749,In_973);
and U4183 (N_4183,In_1409,In_2339);
and U4184 (N_4184,In_9,In_1943);
nor U4185 (N_4185,In_831,In_1288);
nor U4186 (N_4186,In_2087,In_2227);
and U4187 (N_4187,In_397,In_1233);
and U4188 (N_4188,In_1442,In_2335);
and U4189 (N_4189,In_1664,In_2439);
nand U4190 (N_4190,In_306,In_251);
nand U4191 (N_4191,In_326,In_2405);
nor U4192 (N_4192,In_561,In_1580);
and U4193 (N_4193,In_1623,In_1596);
and U4194 (N_4194,In_603,In_2223);
nand U4195 (N_4195,In_2158,In_1150);
nor U4196 (N_4196,In_2472,In_2020);
or U4197 (N_4197,In_339,In_1058);
nor U4198 (N_4198,In_414,In_1352);
or U4199 (N_4199,In_2467,In_1459);
nand U4200 (N_4200,In_1731,In_804);
or U4201 (N_4201,In_1450,In_1883);
nor U4202 (N_4202,In_1914,In_1233);
xor U4203 (N_4203,In_1850,In_2297);
nor U4204 (N_4204,In_527,In_2118);
or U4205 (N_4205,In_2058,In_105);
nor U4206 (N_4206,In_386,In_1333);
xnor U4207 (N_4207,In_2109,In_437);
nand U4208 (N_4208,In_1125,In_1613);
nor U4209 (N_4209,In_629,In_2307);
or U4210 (N_4210,In_1297,In_1544);
or U4211 (N_4211,In_2266,In_611);
nand U4212 (N_4212,In_196,In_1526);
and U4213 (N_4213,In_1883,In_772);
xnor U4214 (N_4214,In_1952,In_269);
and U4215 (N_4215,In_589,In_1954);
or U4216 (N_4216,In_2360,In_1040);
or U4217 (N_4217,In_1040,In_2100);
nand U4218 (N_4218,In_1636,In_335);
nand U4219 (N_4219,In_2237,In_696);
nand U4220 (N_4220,In_565,In_806);
nor U4221 (N_4221,In_161,In_814);
nor U4222 (N_4222,In_458,In_456);
nor U4223 (N_4223,In_2101,In_450);
or U4224 (N_4224,In_2200,In_406);
xnor U4225 (N_4225,In_1141,In_441);
or U4226 (N_4226,In_2450,In_2051);
nand U4227 (N_4227,In_889,In_1584);
nand U4228 (N_4228,In_2278,In_1914);
or U4229 (N_4229,In_473,In_2442);
xor U4230 (N_4230,In_1876,In_2315);
and U4231 (N_4231,In_2365,In_1336);
xor U4232 (N_4232,In_554,In_1433);
and U4233 (N_4233,In_2377,In_195);
nor U4234 (N_4234,In_364,In_1052);
and U4235 (N_4235,In_1326,In_72);
or U4236 (N_4236,In_1990,In_327);
xor U4237 (N_4237,In_872,In_824);
xnor U4238 (N_4238,In_2069,In_1916);
and U4239 (N_4239,In_2028,In_1466);
and U4240 (N_4240,In_628,In_932);
nand U4241 (N_4241,In_352,In_1081);
nor U4242 (N_4242,In_1035,In_1991);
xor U4243 (N_4243,In_2384,In_424);
or U4244 (N_4244,In_1876,In_1823);
xor U4245 (N_4245,In_1067,In_499);
nor U4246 (N_4246,In_1631,In_1539);
or U4247 (N_4247,In_720,In_1148);
and U4248 (N_4248,In_2331,In_891);
nor U4249 (N_4249,In_2108,In_2134);
nor U4250 (N_4250,In_1684,In_730);
xor U4251 (N_4251,In_1681,In_123);
xor U4252 (N_4252,In_1916,In_298);
nor U4253 (N_4253,In_1031,In_2343);
or U4254 (N_4254,In_288,In_2434);
xor U4255 (N_4255,In_1300,In_1758);
and U4256 (N_4256,In_1012,In_2421);
and U4257 (N_4257,In_1172,In_967);
or U4258 (N_4258,In_813,In_1182);
and U4259 (N_4259,In_19,In_703);
or U4260 (N_4260,In_305,In_1868);
or U4261 (N_4261,In_869,In_1937);
nand U4262 (N_4262,In_311,In_984);
and U4263 (N_4263,In_1460,In_1100);
or U4264 (N_4264,In_11,In_311);
nand U4265 (N_4265,In_1071,In_1179);
xnor U4266 (N_4266,In_2266,In_911);
and U4267 (N_4267,In_1914,In_1344);
xnor U4268 (N_4268,In_751,In_2485);
xor U4269 (N_4269,In_274,In_1539);
or U4270 (N_4270,In_553,In_2220);
and U4271 (N_4271,In_1473,In_1521);
xor U4272 (N_4272,In_930,In_324);
or U4273 (N_4273,In_882,In_965);
or U4274 (N_4274,In_182,In_2489);
nor U4275 (N_4275,In_1137,In_1409);
and U4276 (N_4276,In_1279,In_19);
and U4277 (N_4277,In_884,In_2393);
nand U4278 (N_4278,In_134,In_420);
nand U4279 (N_4279,In_1668,In_717);
or U4280 (N_4280,In_2192,In_534);
and U4281 (N_4281,In_1761,In_1191);
or U4282 (N_4282,In_274,In_1646);
nand U4283 (N_4283,In_1586,In_2065);
or U4284 (N_4284,In_1773,In_101);
or U4285 (N_4285,In_1998,In_2329);
or U4286 (N_4286,In_1108,In_736);
and U4287 (N_4287,In_2289,In_1809);
nor U4288 (N_4288,In_2198,In_1971);
xor U4289 (N_4289,In_136,In_1894);
nor U4290 (N_4290,In_1309,In_328);
and U4291 (N_4291,In_2452,In_1379);
and U4292 (N_4292,In_936,In_588);
xnor U4293 (N_4293,In_2221,In_1607);
nand U4294 (N_4294,In_1098,In_418);
and U4295 (N_4295,In_458,In_2211);
or U4296 (N_4296,In_1904,In_128);
and U4297 (N_4297,In_546,In_64);
xor U4298 (N_4298,In_2494,In_1869);
and U4299 (N_4299,In_884,In_450);
xnor U4300 (N_4300,In_1004,In_1896);
or U4301 (N_4301,In_1756,In_1240);
or U4302 (N_4302,In_872,In_820);
nand U4303 (N_4303,In_1532,In_796);
xor U4304 (N_4304,In_976,In_643);
xnor U4305 (N_4305,In_18,In_2033);
xnor U4306 (N_4306,In_824,In_1097);
nor U4307 (N_4307,In_930,In_1770);
or U4308 (N_4308,In_1676,In_53);
and U4309 (N_4309,In_960,In_860);
nor U4310 (N_4310,In_863,In_1445);
xnor U4311 (N_4311,In_1706,In_2090);
and U4312 (N_4312,In_1924,In_1096);
xnor U4313 (N_4313,In_1887,In_2233);
xor U4314 (N_4314,In_44,In_429);
or U4315 (N_4315,In_1033,In_2385);
xor U4316 (N_4316,In_880,In_1411);
and U4317 (N_4317,In_2022,In_1506);
xnor U4318 (N_4318,In_1046,In_2115);
and U4319 (N_4319,In_129,In_1620);
or U4320 (N_4320,In_715,In_1634);
nand U4321 (N_4321,In_116,In_615);
or U4322 (N_4322,In_150,In_1161);
nand U4323 (N_4323,In_633,In_2227);
xor U4324 (N_4324,In_1396,In_2088);
or U4325 (N_4325,In_1928,In_1112);
nand U4326 (N_4326,In_2485,In_1961);
xor U4327 (N_4327,In_1661,In_2245);
nand U4328 (N_4328,In_1692,In_2444);
and U4329 (N_4329,In_9,In_1597);
or U4330 (N_4330,In_1,In_2430);
and U4331 (N_4331,In_653,In_1865);
and U4332 (N_4332,In_1283,In_801);
and U4333 (N_4333,In_220,In_2320);
nor U4334 (N_4334,In_759,In_432);
nor U4335 (N_4335,In_1171,In_785);
nand U4336 (N_4336,In_250,In_1678);
nand U4337 (N_4337,In_856,In_1509);
nor U4338 (N_4338,In_169,In_1601);
xnor U4339 (N_4339,In_1827,In_1057);
nand U4340 (N_4340,In_2110,In_133);
nor U4341 (N_4341,In_691,In_1391);
xnor U4342 (N_4342,In_1418,In_1779);
and U4343 (N_4343,In_1632,In_2208);
nand U4344 (N_4344,In_1008,In_271);
or U4345 (N_4345,In_2063,In_390);
nor U4346 (N_4346,In_1325,In_1062);
and U4347 (N_4347,In_1873,In_1672);
xnor U4348 (N_4348,In_1767,In_2068);
xnor U4349 (N_4349,In_1694,In_1975);
and U4350 (N_4350,In_1407,In_1479);
or U4351 (N_4351,In_1759,In_1292);
nand U4352 (N_4352,In_296,In_198);
xnor U4353 (N_4353,In_1003,In_2071);
or U4354 (N_4354,In_1666,In_1800);
xnor U4355 (N_4355,In_1427,In_1830);
nor U4356 (N_4356,In_1033,In_1130);
or U4357 (N_4357,In_1069,In_1309);
nand U4358 (N_4358,In_217,In_1455);
or U4359 (N_4359,In_1287,In_58);
xnor U4360 (N_4360,In_1867,In_1922);
nor U4361 (N_4361,In_621,In_2327);
xnor U4362 (N_4362,In_1787,In_63);
nand U4363 (N_4363,In_1798,In_2261);
nor U4364 (N_4364,In_2348,In_92);
nor U4365 (N_4365,In_686,In_2062);
nand U4366 (N_4366,In_742,In_602);
nor U4367 (N_4367,In_1132,In_583);
or U4368 (N_4368,In_945,In_2331);
or U4369 (N_4369,In_1728,In_1900);
and U4370 (N_4370,In_2021,In_1937);
nand U4371 (N_4371,In_813,In_548);
or U4372 (N_4372,In_957,In_0);
or U4373 (N_4373,In_1896,In_1578);
xnor U4374 (N_4374,In_262,In_1159);
nand U4375 (N_4375,In_528,In_2209);
nor U4376 (N_4376,In_1747,In_1944);
and U4377 (N_4377,In_1525,In_1104);
or U4378 (N_4378,In_1174,In_1368);
nor U4379 (N_4379,In_404,In_130);
and U4380 (N_4380,In_1674,In_588);
and U4381 (N_4381,In_1207,In_2316);
xor U4382 (N_4382,In_707,In_545);
xor U4383 (N_4383,In_224,In_106);
nand U4384 (N_4384,In_401,In_1699);
nand U4385 (N_4385,In_1677,In_886);
nand U4386 (N_4386,In_161,In_700);
xnor U4387 (N_4387,In_321,In_1856);
and U4388 (N_4388,In_2325,In_516);
nand U4389 (N_4389,In_45,In_1705);
and U4390 (N_4390,In_1329,In_1545);
nor U4391 (N_4391,In_1319,In_102);
and U4392 (N_4392,In_1176,In_1275);
nor U4393 (N_4393,In_831,In_1796);
and U4394 (N_4394,In_1264,In_22);
nor U4395 (N_4395,In_2277,In_1664);
nor U4396 (N_4396,In_2458,In_1598);
or U4397 (N_4397,In_1314,In_2426);
nor U4398 (N_4398,In_1272,In_195);
xnor U4399 (N_4399,In_857,In_1262);
nand U4400 (N_4400,In_346,In_228);
and U4401 (N_4401,In_914,In_1363);
xor U4402 (N_4402,In_1860,In_454);
or U4403 (N_4403,In_1712,In_1592);
nor U4404 (N_4404,In_330,In_1046);
xor U4405 (N_4405,In_2460,In_1955);
nand U4406 (N_4406,In_1653,In_791);
or U4407 (N_4407,In_1552,In_720);
nand U4408 (N_4408,In_695,In_1419);
nor U4409 (N_4409,In_1811,In_2120);
xor U4410 (N_4410,In_2473,In_998);
nor U4411 (N_4411,In_1991,In_1290);
or U4412 (N_4412,In_1717,In_1377);
nor U4413 (N_4413,In_646,In_184);
nor U4414 (N_4414,In_1445,In_2255);
nor U4415 (N_4415,In_1508,In_2347);
xnor U4416 (N_4416,In_1970,In_1750);
and U4417 (N_4417,In_1489,In_2321);
nand U4418 (N_4418,In_359,In_2049);
and U4419 (N_4419,In_1181,In_1800);
nand U4420 (N_4420,In_2257,In_659);
nor U4421 (N_4421,In_617,In_755);
nand U4422 (N_4422,In_2257,In_2143);
xnor U4423 (N_4423,In_772,In_616);
or U4424 (N_4424,In_1676,In_908);
nor U4425 (N_4425,In_2395,In_838);
xor U4426 (N_4426,In_1974,In_1916);
nor U4427 (N_4427,In_378,In_708);
nand U4428 (N_4428,In_2301,In_1181);
xor U4429 (N_4429,In_1226,In_2146);
xnor U4430 (N_4430,In_977,In_1400);
and U4431 (N_4431,In_1833,In_653);
nor U4432 (N_4432,In_1712,In_1466);
nor U4433 (N_4433,In_215,In_1137);
or U4434 (N_4434,In_216,In_1404);
and U4435 (N_4435,In_155,In_2148);
nand U4436 (N_4436,In_1681,In_1708);
nand U4437 (N_4437,In_1119,In_1116);
and U4438 (N_4438,In_1578,In_2016);
and U4439 (N_4439,In_1171,In_1479);
nand U4440 (N_4440,In_310,In_1139);
and U4441 (N_4441,In_67,In_1795);
or U4442 (N_4442,In_201,In_237);
nand U4443 (N_4443,In_530,In_1399);
nand U4444 (N_4444,In_653,In_1427);
nor U4445 (N_4445,In_2487,In_304);
or U4446 (N_4446,In_1348,In_787);
xnor U4447 (N_4447,In_2346,In_318);
nand U4448 (N_4448,In_303,In_1290);
and U4449 (N_4449,In_0,In_1031);
nor U4450 (N_4450,In_2279,In_210);
and U4451 (N_4451,In_2180,In_558);
and U4452 (N_4452,In_2203,In_1240);
or U4453 (N_4453,In_1140,In_2349);
nand U4454 (N_4454,In_702,In_1683);
nand U4455 (N_4455,In_1773,In_2335);
and U4456 (N_4456,In_1943,In_1484);
or U4457 (N_4457,In_1245,In_670);
xor U4458 (N_4458,In_1891,In_1075);
nor U4459 (N_4459,In_1287,In_1195);
or U4460 (N_4460,In_943,In_1770);
nor U4461 (N_4461,In_1401,In_1029);
or U4462 (N_4462,In_2489,In_669);
nor U4463 (N_4463,In_1104,In_2039);
nor U4464 (N_4464,In_2084,In_1308);
nor U4465 (N_4465,In_254,In_1906);
nor U4466 (N_4466,In_305,In_1158);
xnor U4467 (N_4467,In_718,In_2468);
xor U4468 (N_4468,In_380,In_583);
xnor U4469 (N_4469,In_559,In_1082);
xnor U4470 (N_4470,In_1226,In_54);
nor U4471 (N_4471,In_636,In_2147);
xnor U4472 (N_4472,In_649,In_1670);
nand U4473 (N_4473,In_749,In_1456);
and U4474 (N_4474,In_902,In_2152);
or U4475 (N_4475,In_1125,In_2099);
nand U4476 (N_4476,In_1713,In_2241);
and U4477 (N_4477,In_1334,In_767);
nor U4478 (N_4478,In_1261,In_115);
xnor U4479 (N_4479,In_2053,In_1588);
or U4480 (N_4480,In_2164,In_2347);
and U4481 (N_4481,In_2407,In_2010);
or U4482 (N_4482,In_1923,In_1475);
nand U4483 (N_4483,In_2265,In_705);
xnor U4484 (N_4484,In_1701,In_1735);
nor U4485 (N_4485,In_743,In_560);
and U4486 (N_4486,In_1077,In_2488);
and U4487 (N_4487,In_713,In_2404);
and U4488 (N_4488,In_903,In_156);
xnor U4489 (N_4489,In_813,In_2253);
or U4490 (N_4490,In_1570,In_459);
nor U4491 (N_4491,In_1281,In_1612);
xnor U4492 (N_4492,In_2052,In_770);
and U4493 (N_4493,In_177,In_826);
and U4494 (N_4494,In_128,In_424);
and U4495 (N_4495,In_2261,In_1202);
and U4496 (N_4496,In_2061,In_2266);
nand U4497 (N_4497,In_1874,In_1834);
nand U4498 (N_4498,In_865,In_2435);
nand U4499 (N_4499,In_1058,In_1476);
nor U4500 (N_4500,In_2244,In_2476);
nor U4501 (N_4501,In_1060,In_771);
nor U4502 (N_4502,In_913,In_1191);
and U4503 (N_4503,In_956,In_1711);
nand U4504 (N_4504,In_213,In_853);
nor U4505 (N_4505,In_660,In_1514);
xor U4506 (N_4506,In_224,In_685);
nor U4507 (N_4507,In_2496,In_1375);
nand U4508 (N_4508,In_1434,In_124);
and U4509 (N_4509,In_1400,In_511);
xor U4510 (N_4510,In_2204,In_2184);
nand U4511 (N_4511,In_852,In_710);
and U4512 (N_4512,In_706,In_1292);
nand U4513 (N_4513,In_1833,In_1285);
and U4514 (N_4514,In_1062,In_272);
and U4515 (N_4515,In_2129,In_235);
nand U4516 (N_4516,In_310,In_2412);
nand U4517 (N_4517,In_1015,In_2332);
or U4518 (N_4518,In_1323,In_1890);
and U4519 (N_4519,In_864,In_1698);
or U4520 (N_4520,In_630,In_2411);
and U4521 (N_4521,In_1908,In_2062);
or U4522 (N_4522,In_1354,In_794);
nand U4523 (N_4523,In_682,In_698);
nand U4524 (N_4524,In_121,In_945);
nand U4525 (N_4525,In_1761,In_286);
nand U4526 (N_4526,In_1155,In_803);
and U4527 (N_4527,In_1159,In_46);
xor U4528 (N_4528,In_1995,In_1042);
or U4529 (N_4529,In_613,In_2309);
nand U4530 (N_4530,In_976,In_1350);
or U4531 (N_4531,In_333,In_2193);
and U4532 (N_4532,In_1133,In_1346);
xnor U4533 (N_4533,In_1174,In_1546);
nor U4534 (N_4534,In_1302,In_2204);
nor U4535 (N_4535,In_1154,In_791);
nor U4536 (N_4536,In_2311,In_243);
nand U4537 (N_4537,In_72,In_1256);
nor U4538 (N_4538,In_2071,In_383);
and U4539 (N_4539,In_1192,In_1485);
nand U4540 (N_4540,In_566,In_247);
and U4541 (N_4541,In_1082,In_2263);
or U4542 (N_4542,In_2099,In_1253);
and U4543 (N_4543,In_981,In_1487);
or U4544 (N_4544,In_921,In_2023);
and U4545 (N_4545,In_826,In_1718);
nor U4546 (N_4546,In_337,In_1981);
or U4547 (N_4547,In_1606,In_686);
xnor U4548 (N_4548,In_683,In_251);
nand U4549 (N_4549,In_1742,In_2240);
nand U4550 (N_4550,In_333,In_1128);
xor U4551 (N_4551,In_1956,In_1960);
nand U4552 (N_4552,In_536,In_1977);
xor U4553 (N_4553,In_33,In_2056);
xnor U4554 (N_4554,In_220,In_1318);
nand U4555 (N_4555,In_656,In_753);
and U4556 (N_4556,In_2094,In_853);
nand U4557 (N_4557,In_2485,In_2488);
nor U4558 (N_4558,In_1233,In_1435);
or U4559 (N_4559,In_1221,In_1064);
nor U4560 (N_4560,In_611,In_309);
or U4561 (N_4561,In_2325,In_1670);
and U4562 (N_4562,In_2493,In_1247);
and U4563 (N_4563,In_1307,In_1477);
nand U4564 (N_4564,In_1507,In_2270);
nand U4565 (N_4565,In_817,In_1964);
and U4566 (N_4566,In_1832,In_979);
xnor U4567 (N_4567,In_1150,In_1990);
nand U4568 (N_4568,In_2256,In_696);
and U4569 (N_4569,In_1755,In_1262);
xnor U4570 (N_4570,In_1118,In_1081);
nand U4571 (N_4571,In_827,In_1058);
and U4572 (N_4572,In_1312,In_284);
and U4573 (N_4573,In_2247,In_1471);
or U4574 (N_4574,In_1327,In_2382);
or U4575 (N_4575,In_1898,In_1694);
xor U4576 (N_4576,In_2096,In_312);
nand U4577 (N_4577,In_1847,In_2498);
nor U4578 (N_4578,In_621,In_553);
xnor U4579 (N_4579,In_1150,In_342);
nand U4580 (N_4580,In_652,In_208);
xnor U4581 (N_4581,In_2135,In_30);
nor U4582 (N_4582,In_475,In_722);
and U4583 (N_4583,In_976,In_1121);
and U4584 (N_4584,In_199,In_322);
nor U4585 (N_4585,In_2405,In_41);
or U4586 (N_4586,In_2498,In_1164);
xnor U4587 (N_4587,In_410,In_1591);
nor U4588 (N_4588,In_587,In_1236);
and U4589 (N_4589,In_1868,In_260);
and U4590 (N_4590,In_660,In_702);
or U4591 (N_4591,In_485,In_396);
nand U4592 (N_4592,In_24,In_704);
or U4593 (N_4593,In_522,In_1456);
or U4594 (N_4594,In_1495,In_1255);
and U4595 (N_4595,In_2308,In_1025);
nor U4596 (N_4596,In_1884,In_904);
xnor U4597 (N_4597,In_899,In_2293);
and U4598 (N_4598,In_926,In_1760);
xnor U4599 (N_4599,In_1267,In_1704);
nor U4600 (N_4600,In_1782,In_137);
nor U4601 (N_4601,In_2243,In_1429);
and U4602 (N_4602,In_652,In_61);
nor U4603 (N_4603,In_673,In_2387);
or U4604 (N_4604,In_46,In_1541);
and U4605 (N_4605,In_1823,In_52);
and U4606 (N_4606,In_588,In_1161);
nor U4607 (N_4607,In_1858,In_969);
xor U4608 (N_4608,In_700,In_1880);
xnor U4609 (N_4609,In_101,In_1894);
or U4610 (N_4610,In_2104,In_1728);
nand U4611 (N_4611,In_1630,In_2028);
xnor U4612 (N_4612,In_1130,In_1465);
and U4613 (N_4613,In_2074,In_854);
nand U4614 (N_4614,In_1061,In_2484);
nor U4615 (N_4615,In_429,In_523);
and U4616 (N_4616,In_1561,In_2192);
and U4617 (N_4617,In_488,In_703);
nor U4618 (N_4618,In_1596,In_1583);
xnor U4619 (N_4619,In_1010,In_1926);
or U4620 (N_4620,In_804,In_1234);
nand U4621 (N_4621,In_2186,In_2084);
nand U4622 (N_4622,In_569,In_2494);
nand U4623 (N_4623,In_340,In_1185);
xor U4624 (N_4624,In_1451,In_1033);
nand U4625 (N_4625,In_1906,In_1329);
nor U4626 (N_4626,In_1507,In_1834);
or U4627 (N_4627,In_1044,In_2117);
and U4628 (N_4628,In_226,In_1559);
and U4629 (N_4629,In_649,In_1756);
nand U4630 (N_4630,In_1337,In_238);
and U4631 (N_4631,In_179,In_517);
and U4632 (N_4632,In_969,In_489);
and U4633 (N_4633,In_2412,In_462);
nor U4634 (N_4634,In_577,In_2398);
nand U4635 (N_4635,In_2495,In_438);
nor U4636 (N_4636,In_2060,In_1294);
or U4637 (N_4637,In_1800,In_1904);
and U4638 (N_4638,In_714,In_1754);
xnor U4639 (N_4639,In_830,In_1648);
xnor U4640 (N_4640,In_2242,In_457);
nor U4641 (N_4641,In_1995,In_1642);
nand U4642 (N_4642,In_1196,In_712);
xor U4643 (N_4643,In_2153,In_1633);
nand U4644 (N_4644,In_2499,In_1638);
nor U4645 (N_4645,In_2135,In_1073);
and U4646 (N_4646,In_484,In_1372);
xnor U4647 (N_4647,In_1673,In_2368);
or U4648 (N_4648,In_1996,In_1603);
or U4649 (N_4649,In_2254,In_1851);
or U4650 (N_4650,In_586,In_1170);
and U4651 (N_4651,In_708,In_2081);
nor U4652 (N_4652,In_2155,In_855);
or U4653 (N_4653,In_1522,In_1425);
and U4654 (N_4654,In_1512,In_2181);
or U4655 (N_4655,In_684,In_1093);
nor U4656 (N_4656,In_2483,In_875);
xor U4657 (N_4657,In_859,In_1691);
or U4658 (N_4658,In_678,In_63);
xnor U4659 (N_4659,In_1905,In_537);
or U4660 (N_4660,In_12,In_703);
nor U4661 (N_4661,In_236,In_1006);
nor U4662 (N_4662,In_1524,In_2024);
nor U4663 (N_4663,In_627,In_560);
xnor U4664 (N_4664,In_282,In_2105);
nor U4665 (N_4665,In_433,In_2156);
xnor U4666 (N_4666,In_1314,In_760);
or U4667 (N_4667,In_171,In_1373);
nand U4668 (N_4668,In_221,In_1908);
xor U4669 (N_4669,In_1892,In_2034);
nand U4670 (N_4670,In_2004,In_956);
and U4671 (N_4671,In_1076,In_1887);
nand U4672 (N_4672,In_1668,In_1182);
and U4673 (N_4673,In_460,In_803);
nor U4674 (N_4674,In_2468,In_880);
xnor U4675 (N_4675,In_705,In_1700);
nand U4676 (N_4676,In_2347,In_926);
xor U4677 (N_4677,In_1832,In_499);
or U4678 (N_4678,In_2073,In_1520);
or U4679 (N_4679,In_1208,In_2197);
or U4680 (N_4680,In_1848,In_763);
or U4681 (N_4681,In_1188,In_291);
nor U4682 (N_4682,In_1479,In_798);
or U4683 (N_4683,In_317,In_1607);
nand U4684 (N_4684,In_1366,In_722);
nand U4685 (N_4685,In_820,In_887);
nor U4686 (N_4686,In_1573,In_748);
or U4687 (N_4687,In_1641,In_2322);
xor U4688 (N_4688,In_422,In_1537);
nor U4689 (N_4689,In_154,In_517);
xnor U4690 (N_4690,In_890,In_786);
xnor U4691 (N_4691,In_2112,In_1683);
or U4692 (N_4692,In_1787,In_1136);
or U4693 (N_4693,In_2021,In_35);
or U4694 (N_4694,In_2301,In_1151);
and U4695 (N_4695,In_950,In_193);
or U4696 (N_4696,In_22,In_880);
nand U4697 (N_4697,In_1435,In_145);
or U4698 (N_4698,In_364,In_1853);
and U4699 (N_4699,In_1298,In_1754);
nor U4700 (N_4700,In_549,In_257);
and U4701 (N_4701,In_997,In_724);
xor U4702 (N_4702,In_343,In_772);
and U4703 (N_4703,In_1688,In_2159);
xor U4704 (N_4704,In_201,In_1519);
and U4705 (N_4705,In_1645,In_578);
xnor U4706 (N_4706,In_1396,In_32);
and U4707 (N_4707,In_1344,In_1778);
nor U4708 (N_4708,In_1917,In_1661);
and U4709 (N_4709,In_1510,In_1009);
nor U4710 (N_4710,In_537,In_954);
xor U4711 (N_4711,In_2455,In_1493);
and U4712 (N_4712,In_778,In_504);
or U4713 (N_4713,In_11,In_2266);
nor U4714 (N_4714,In_471,In_1508);
xor U4715 (N_4715,In_481,In_1768);
xor U4716 (N_4716,In_2330,In_2031);
nor U4717 (N_4717,In_1114,In_923);
nand U4718 (N_4718,In_1860,In_890);
or U4719 (N_4719,In_1260,In_1437);
nor U4720 (N_4720,In_2390,In_2417);
or U4721 (N_4721,In_1122,In_1504);
xnor U4722 (N_4722,In_523,In_2310);
nor U4723 (N_4723,In_2462,In_1077);
nor U4724 (N_4724,In_1682,In_98);
or U4725 (N_4725,In_427,In_1741);
or U4726 (N_4726,In_1551,In_2017);
nand U4727 (N_4727,In_2285,In_2229);
and U4728 (N_4728,In_1720,In_826);
and U4729 (N_4729,In_484,In_525);
nor U4730 (N_4730,In_709,In_244);
nor U4731 (N_4731,In_1404,In_2330);
nand U4732 (N_4732,In_911,In_1188);
nor U4733 (N_4733,In_1563,In_1977);
nor U4734 (N_4734,In_477,In_1390);
or U4735 (N_4735,In_2353,In_2016);
nand U4736 (N_4736,In_2228,In_1750);
xnor U4737 (N_4737,In_2182,In_1885);
xnor U4738 (N_4738,In_495,In_919);
nor U4739 (N_4739,In_1892,In_240);
xnor U4740 (N_4740,In_2320,In_2276);
nand U4741 (N_4741,In_919,In_1864);
or U4742 (N_4742,In_2210,In_108);
nand U4743 (N_4743,In_72,In_164);
xor U4744 (N_4744,In_853,In_1779);
nor U4745 (N_4745,In_1865,In_1051);
nand U4746 (N_4746,In_788,In_2002);
nor U4747 (N_4747,In_1236,In_270);
nand U4748 (N_4748,In_872,In_712);
or U4749 (N_4749,In_68,In_1918);
nor U4750 (N_4750,In_1854,In_1463);
nand U4751 (N_4751,In_1934,In_996);
xnor U4752 (N_4752,In_1625,In_557);
or U4753 (N_4753,In_2097,In_1245);
xnor U4754 (N_4754,In_762,In_1424);
nand U4755 (N_4755,In_1264,In_1565);
or U4756 (N_4756,In_2174,In_1509);
xor U4757 (N_4757,In_840,In_1863);
or U4758 (N_4758,In_1588,In_1695);
nand U4759 (N_4759,In_1551,In_1556);
xnor U4760 (N_4760,In_2093,In_2103);
nor U4761 (N_4761,In_917,In_1903);
nand U4762 (N_4762,In_501,In_300);
and U4763 (N_4763,In_1132,In_422);
or U4764 (N_4764,In_2440,In_2367);
nand U4765 (N_4765,In_1419,In_452);
xor U4766 (N_4766,In_1671,In_247);
xnor U4767 (N_4767,In_2345,In_2417);
or U4768 (N_4768,In_1519,In_1856);
xnor U4769 (N_4769,In_1294,In_73);
and U4770 (N_4770,In_211,In_1806);
nor U4771 (N_4771,In_1440,In_997);
nand U4772 (N_4772,In_374,In_935);
xor U4773 (N_4773,In_1687,In_1686);
and U4774 (N_4774,In_2015,In_317);
or U4775 (N_4775,In_1151,In_2354);
nor U4776 (N_4776,In_781,In_320);
nand U4777 (N_4777,In_84,In_1199);
or U4778 (N_4778,In_468,In_1670);
or U4779 (N_4779,In_1974,In_34);
nor U4780 (N_4780,In_1593,In_1591);
or U4781 (N_4781,In_87,In_453);
or U4782 (N_4782,In_1037,In_94);
xnor U4783 (N_4783,In_1609,In_934);
nor U4784 (N_4784,In_2282,In_2175);
nand U4785 (N_4785,In_1990,In_1116);
or U4786 (N_4786,In_1184,In_1985);
and U4787 (N_4787,In_1155,In_1541);
and U4788 (N_4788,In_1967,In_1053);
xor U4789 (N_4789,In_2130,In_824);
nor U4790 (N_4790,In_1719,In_1008);
nand U4791 (N_4791,In_167,In_2053);
and U4792 (N_4792,In_420,In_19);
nand U4793 (N_4793,In_2294,In_2002);
and U4794 (N_4794,In_2346,In_955);
nor U4795 (N_4795,In_138,In_422);
nor U4796 (N_4796,In_2055,In_1480);
nor U4797 (N_4797,In_2294,In_86);
xor U4798 (N_4798,In_556,In_1855);
xnor U4799 (N_4799,In_714,In_753);
xor U4800 (N_4800,In_1922,In_2385);
nor U4801 (N_4801,In_1270,In_1371);
nor U4802 (N_4802,In_2471,In_498);
and U4803 (N_4803,In_826,In_1627);
nand U4804 (N_4804,In_54,In_1711);
nand U4805 (N_4805,In_751,In_1347);
or U4806 (N_4806,In_1065,In_2239);
and U4807 (N_4807,In_485,In_1891);
xor U4808 (N_4808,In_2260,In_2231);
nor U4809 (N_4809,In_216,In_1646);
nor U4810 (N_4810,In_2437,In_1625);
or U4811 (N_4811,In_204,In_1285);
xor U4812 (N_4812,In_1931,In_1471);
xnor U4813 (N_4813,In_2051,In_2387);
and U4814 (N_4814,In_704,In_173);
or U4815 (N_4815,In_2343,In_1429);
or U4816 (N_4816,In_1886,In_1200);
and U4817 (N_4817,In_1035,In_34);
nor U4818 (N_4818,In_63,In_82);
xnor U4819 (N_4819,In_1116,In_2210);
and U4820 (N_4820,In_68,In_1088);
xnor U4821 (N_4821,In_2194,In_2142);
or U4822 (N_4822,In_2270,In_937);
xor U4823 (N_4823,In_416,In_252);
xor U4824 (N_4824,In_2191,In_1394);
nor U4825 (N_4825,In_799,In_1528);
xor U4826 (N_4826,In_1504,In_11);
and U4827 (N_4827,In_1753,In_1097);
or U4828 (N_4828,In_1986,In_834);
and U4829 (N_4829,In_2263,In_1222);
nand U4830 (N_4830,In_1330,In_695);
nor U4831 (N_4831,In_2129,In_1681);
nand U4832 (N_4832,In_1821,In_1684);
xor U4833 (N_4833,In_1186,In_1010);
and U4834 (N_4834,In_2031,In_670);
or U4835 (N_4835,In_503,In_865);
nand U4836 (N_4836,In_1615,In_27);
nand U4837 (N_4837,In_616,In_1984);
and U4838 (N_4838,In_1071,In_1289);
or U4839 (N_4839,In_969,In_1925);
xnor U4840 (N_4840,In_2358,In_1171);
or U4841 (N_4841,In_890,In_1684);
xnor U4842 (N_4842,In_2198,In_1729);
nand U4843 (N_4843,In_488,In_954);
nand U4844 (N_4844,In_124,In_939);
and U4845 (N_4845,In_2448,In_1321);
nor U4846 (N_4846,In_1120,In_1020);
and U4847 (N_4847,In_2178,In_814);
and U4848 (N_4848,In_1969,In_645);
and U4849 (N_4849,In_1073,In_1232);
or U4850 (N_4850,In_1344,In_209);
nor U4851 (N_4851,In_1382,In_742);
nor U4852 (N_4852,In_484,In_2398);
xor U4853 (N_4853,In_131,In_1595);
xor U4854 (N_4854,In_727,In_1489);
and U4855 (N_4855,In_568,In_869);
nand U4856 (N_4856,In_772,In_1477);
or U4857 (N_4857,In_2272,In_768);
or U4858 (N_4858,In_1492,In_2471);
xor U4859 (N_4859,In_2468,In_324);
and U4860 (N_4860,In_382,In_1412);
or U4861 (N_4861,In_2227,In_1905);
nand U4862 (N_4862,In_2425,In_214);
xnor U4863 (N_4863,In_1086,In_2039);
or U4864 (N_4864,In_82,In_238);
or U4865 (N_4865,In_1450,In_2461);
xnor U4866 (N_4866,In_672,In_1999);
xor U4867 (N_4867,In_1379,In_138);
nor U4868 (N_4868,In_1815,In_2078);
and U4869 (N_4869,In_1237,In_162);
or U4870 (N_4870,In_1477,In_1095);
xor U4871 (N_4871,In_1469,In_989);
nor U4872 (N_4872,In_446,In_998);
and U4873 (N_4873,In_1640,In_2008);
and U4874 (N_4874,In_1855,In_1119);
or U4875 (N_4875,In_2493,In_292);
or U4876 (N_4876,In_44,In_1494);
nor U4877 (N_4877,In_372,In_849);
nand U4878 (N_4878,In_2261,In_2177);
and U4879 (N_4879,In_1850,In_1988);
nand U4880 (N_4880,In_1106,In_1214);
xor U4881 (N_4881,In_16,In_1588);
nand U4882 (N_4882,In_2357,In_823);
and U4883 (N_4883,In_829,In_1486);
nand U4884 (N_4884,In_1383,In_39);
nor U4885 (N_4885,In_1016,In_1072);
nand U4886 (N_4886,In_1297,In_1153);
and U4887 (N_4887,In_2091,In_1968);
nand U4888 (N_4888,In_2329,In_1104);
or U4889 (N_4889,In_967,In_997);
nor U4890 (N_4890,In_316,In_673);
and U4891 (N_4891,In_2066,In_803);
and U4892 (N_4892,In_2381,In_2287);
nand U4893 (N_4893,In_196,In_1386);
nand U4894 (N_4894,In_1944,In_1278);
nor U4895 (N_4895,In_844,In_2159);
nor U4896 (N_4896,In_1639,In_180);
nand U4897 (N_4897,In_618,In_1169);
nand U4898 (N_4898,In_1472,In_106);
and U4899 (N_4899,In_1546,In_1405);
and U4900 (N_4900,In_674,In_616);
xnor U4901 (N_4901,In_1628,In_1281);
and U4902 (N_4902,In_1738,In_1334);
and U4903 (N_4903,In_261,In_1826);
xor U4904 (N_4904,In_566,In_421);
xnor U4905 (N_4905,In_2132,In_2306);
nand U4906 (N_4906,In_349,In_1491);
xor U4907 (N_4907,In_663,In_2386);
nand U4908 (N_4908,In_1463,In_296);
or U4909 (N_4909,In_1111,In_439);
nand U4910 (N_4910,In_1416,In_1245);
xnor U4911 (N_4911,In_1712,In_1029);
nand U4912 (N_4912,In_851,In_2167);
and U4913 (N_4913,In_1728,In_658);
nor U4914 (N_4914,In_957,In_1759);
or U4915 (N_4915,In_1938,In_363);
nand U4916 (N_4916,In_91,In_515);
xor U4917 (N_4917,In_2419,In_1986);
and U4918 (N_4918,In_1354,In_1088);
xor U4919 (N_4919,In_570,In_1844);
nor U4920 (N_4920,In_517,In_507);
or U4921 (N_4921,In_830,In_1065);
xnor U4922 (N_4922,In_558,In_1287);
nor U4923 (N_4923,In_880,In_1050);
and U4924 (N_4924,In_922,In_1394);
and U4925 (N_4925,In_447,In_1745);
or U4926 (N_4926,In_38,In_1943);
xnor U4927 (N_4927,In_1975,In_1150);
xor U4928 (N_4928,In_942,In_1740);
nor U4929 (N_4929,In_2484,In_1607);
nor U4930 (N_4930,In_1595,In_1033);
nor U4931 (N_4931,In_126,In_2472);
or U4932 (N_4932,In_1434,In_1755);
xor U4933 (N_4933,In_382,In_2285);
nor U4934 (N_4934,In_489,In_2384);
nand U4935 (N_4935,In_862,In_1851);
and U4936 (N_4936,In_33,In_35);
nand U4937 (N_4937,In_1208,In_447);
nand U4938 (N_4938,In_1094,In_378);
and U4939 (N_4939,In_1991,In_291);
nand U4940 (N_4940,In_726,In_867);
or U4941 (N_4941,In_950,In_279);
and U4942 (N_4942,In_1063,In_1532);
or U4943 (N_4943,In_1959,In_2163);
nor U4944 (N_4944,In_1075,In_685);
or U4945 (N_4945,In_552,In_1446);
or U4946 (N_4946,In_1649,In_2094);
or U4947 (N_4947,In_1851,In_673);
nand U4948 (N_4948,In_2448,In_1563);
and U4949 (N_4949,In_1311,In_2124);
nand U4950 (N_4950,In_1376,In_1691);
nor U4951 (N_4951,In_1661,In_1094);
xor U4952 (N_4952,In_1183,In_2275);
or U4953 (N_4953,In_1170,In_828);
and U4954 (N_4954,In_505,In_1022);
nor U4955 (N_4955,In_2349,In_117);
and U4956 (N_4956,In_748,In_2215);
nand U4957 (N_4957,In_686,In_722);
nor U4958 (N_4958,In_163,In_1602);
and U4959 (N_4959,In_1374,In_2022);
xor U4960 (N_4960,In_563,In_725);
nand U4961 (N_4961,In_1462,In_1067);
nand U4962 (N_4962,In_1832,In_1551);
and U4963 (N_4963,In_587,In_933);
and U4964 (N_4964,In_911,In_1707);
or U4965 (N_4965,In_66,In_2148);
and U4966 (N_4966,In_1680,In_565);
and U4967 (N_4967,In_1349,In_503);
nor U4968 (N_4968,In_1203,In_1086);
xor U4969 (N_4969,In_2051,In_156);
nand U4970 (N_4970,In_544,In_754);
or U4971 (N_4971,In_1270,In_1871);
nor U4972 (N_4972,In_1421,In_1345);
or U4973 (N_4973,In_1144,In_1840);
and U4974 (N_4974,In_1229,In_2210);
or U4975 (N_4975,In_2346,In_782);
nand U4976 (N_4976,In_259,In_457);
nor U4977 (N_4977,In_1125,In_1354);
nand U4978 (N_4978,In_1017,In_2403);
nor U4979 (N_4979,In_699,In_149);
xor U4980 (N_4980,In_1428,In_273);
nor U4981 (N_4981,In_811,In_643);
nand U4982 (N_4982,In_1695,In_2161);
xor U4983 (N_4983,In_1313,In_2072);
xor U4984 (N_4984,In_121,In_2272);
nand U4985 (N_4985,In_1896,In_483);
and U4986 (N_4986,In_982,In_843);
or U4987 (N_4987,In_635,In_1028);
xnor U4988 (N_4988,In_1040,In_1011);
nor U4989 (N_4989,In_268,In_451);
or U4990 (N_4990,In_1949,In_1844);
or U4991 (N_4991,In_470,In_2287);
nor U4992 (N_4992,In_1027,In_2342);
and U4993 (N_4993,In_693,In_2428);
and U4994 (N_4994,In_129,In_983);
and U4995 (N_4995,In_708,In_626);
and U4996 (N_4996,In_1930,In_15);
xnor U4997 (N_4997,In_1051,In_1921);
nand U4998 (N_4998,In_2470,In_1294);
xor U4999 (N_4999,In_649,In_1036);
nand U5000 (N_5000,In_133,In_136);
or U5001 (N_5001,In_1503,In_898);
or U5002 (N_5002,In_2224,In_1753);
nand U5003 (N_5003,In_604,In_642);
or U5004 (N_5004,In_1354,In_413);
and U5005 (N_5005,In_1879,In_1026);
or U5006 (N_5006,In_709,In_492);
or U5007 (N_5007,In_1847,In_285);
nand U5008 (N_5008,In_1421,In_2408);
or U5009 (N_5009,In_2120,In_2216);
nor U5010 (N_5010,In_716,In_1567);
and U5011 (N_5011,In_2121,In_128);
nand U5012 (N_5012,In_740,In_1435);
xnor U5013 (N_5013,In_1358,In_2403);
and U5014 (N_5014,In_722,In_1486);
or U5015 (N_5015,In_1886,In_2030);
nor U5016 (N_5016,In_1801,In_567);
and U5017 (N_5017,In_1591,In_1124);
or U5018 (N_5018,In_1988,In_1929);
xnor U5019 (N_5019,In_2209,In_23);
and U5020 (N_5020,In_440,In_2142);
and U5021 (N_5021,In_548,In_1746);
nand U5022 (N_5022,In_866,In_651);
and U5023 (N_5023,In_2270,In_2417);
or U5024 (N_5024,In_1933,In_1611);
nor U5025 (N_5025,In_2093,In_1435);
xnor U5026 (N_5026,In_2475,In_454);
nor U5027 (N_5027,In_1207,In_2480);
and U5028 (N_5028,In_873,In_74);
nand U5029 (N_5029,In_1537,In_1327);
or U5030 (N_5030,In_475,In_603);
xor U5031 (N_5031,In_386,In_137);
xor U5032 (N_5032,In_866,In_863);
xor U5033 (N_5033,In_979,In_1398);
and U5034 (N_5034,In_1821,In_2439);
and U5035 (N_5035,In_1113,In_1229);
and U5036 (N_5036,In_282,In_377);
and U5037 (N_5037,In_679,In_1836);
xor U5038 (N_5038,In_2236,In_670);
nand U5039 (N_5039,In_1337,In_709);
nor U5040 (N_5040,In_552,In_1300);
nand U5041 (N_5041,In_628,In_741);
nor U5042 (N_5042,In_1305,In_793);
or U5043 (N_5043,In_2053,In_2293);
and U5044 (N_5044,In_1385,In_1249);
and U5045 (N_5045,In_804,In_1076);
or U5046 (N_5046,In_494,In_1157);
nor U5047 (N_5047,In_1921,In_2408);
or U5048 (N_5048,In_1132,In_2031);
and U5049 (N_5049,In_1078,In_1566);
nand U5050 (N_5050,In_1579,In_1316);
and U5051 (N_5051,In_1798,In_242);
nor U5052 (N_5052,In_1185,In_503);
nor U5053 (N_5053,In_1003,In_1582);
or U5054 (N_5054,In_1947,In_1139);
xnor U5055 (N_5055,In_1637,In_882);
or U5056 (N_5056,In_1732,In_208);
nor U5057 (N_5057,In_315,In_401);
nor U5058 (N_5058,In_333,In_266);
and U5059 (N_5059,In_750,In_771);
nor U5060 (N_5060,In_467,In_1379);
and U5061 (N_5061,In_1209,In_2479);
nor U5062 (N_5062,In_985,In_1875);
xnor U5063 (N_5063,In_1936,In_2146);
and U5064 (N_5064,In_1321,In_480);
or U5065 (N_5065,In_564,In_1130);
nor U5066 (N_5066,In_2333,In_1474);
nand U5067 (N_5067,In_1316,In_143);
nor U5068 (N_5068,In_2298,In_1080);
nor U5069 (N_5069,In_324,In_543);
or U5070 (N_5070,In_747,In_764);
or U5071 (N_5071,In_322,In_1902);
nor U5072 (N_5072,In_244,In_2197);
nand U5073 (N_5073,In_821,In_419);
nor U5074 (N_5074,In_932,In_2291);
and U5075 (N_5075,In_2388,In_1630);
or U5076 (N_5076,In_15,In_1565);
nand U5077 (N_5077,In_490,In_2377);
or U5078 (N_5078,In_1533,In_1235);
nand U5079 (N_5079,In_1095,In_2157);
nand U5080 (N_5080,In_603,In_1363);
nand U5081 (N_5081,In_171,In_711);
xnor U5082 (N_5082,In_2393,In_1991);
xor U5083 (N_5083,In_1744,In_1169);
nand U5084 (N_5084,In_1526,In_144);
and U5085 (N_5085,In_1495,In_1632);
xor U5086 (N_5086,In_991,In_2291);
or U5087 (N_5087,In_1226,In_102);
nor U5088 (N_5088,In_269,In_661);
and U5089 (N_5089,In_289,In_2276);
and U5090 (N_5090,In_2094,In_913);
nor U5091 (N_5091,In_1027,In_445);
nand U5092 (N_5092,In_620,In_2240);
and U5093 (N_5093,In_1319,In_1035);
nand U5094 (N_5094,In_671,In_1386);
xnor U5095 (N_5095,In_734,In_458);
and U5096 (N_5096,In_1388,In_1036);
nor U5097 (N_5097,In_414,In_1381);
nor U5098 (N_5098,In_1868,In_607);
xnor U5099 (N_5099,In_2482,In_121);
nand U5100 (N_5100,In_2106,In_681);
or U5101 (N_5101,In_68,In_374);
and U5102 (N_5102,In_950,In_1875);
nand U5103 (N_5103,In_1460,In_371);
and U5104 (N_5104,In_1079,In_17);
nor U5105 (N_5105,In_1150,In_1647);
nand U5106 (N_5106,In_2284,In_1785);
or U5107 (N_5107,In_2285,In_2338);
and U5108 (N_5108,In_1335,In_2219);
nand U5109 (N_5109,In_776,In_1409);
or U5110 (N_5110,In_562,In_1956);
nor U5111 (N_5111,In_297,In_959);
nand U5112 (N_5112,In_2485,In_378);
xnor U5113 (N_5113,In_320,In_606);
xnor U5114 (N_5114,In_8,In_778);
and U5115 (N_5115,In_484,In_1267);
xor U5116 (N_5116,In_981,In_2043);
and U5117 (N_5117,In_2317,In_2421);
and U5118 (N_5118,In_1211,In_1105);
and U5119 (N_5119,In_413,In_1848);
or U5120 (N_5120,In_2194,In_490);
or U5121 (N_5121,In_929,In_2456);
xnor U5122 (N_5122,In_848,In_178);
and U5123 (N_5123,In_132,In_1153);
nand U5124 (N_5124,In_562,In_2471);
nand U5125 (N_5125,In_2426,In_1);
or U5126 (N_5126,In_2399,In_583);
xnor U5127 (N_5127,In_1924,In_2423);
xnor U5128 (N_5128,In_1190,In_2273);
nor U5129 (N_5129,In_560,In_1641);
xnor U5130 (N_5130,In_1641,In_1517);
xor U5131 (N_5131,In_729,In_335);
nor U5132 (N_5132,In_729,In_2380);
nor U5133 (N_5133,In_1279,In_2324);
xnor U5134 (N_5134,In_2226,In_1308);
nand U5135 (N_5135,In_664,In_2369);
nand U5136 (N_5136,In_29,In_1801);
or U5137 (N_5137,In_2124,In_1351);
or U5138 (N_5138,In_2289,In_1065);
and U5139 (N_5139,In_2366,In_1565);
nor U5140 (N_5140,In_2256,In_38);
nor U5141 (N_5141,In_857,In_1107);
nand U5142 (N_5142,In_1570,In_785);
nand U5143 (N_5143,In_2052,In_630);
or U5144 (N_5144,In_2091,In_1101);
nor U5145 (N_5145,In_2471,In_2310);
xor U5146 (N_5146,In_745,In_2448);
or U5147 (N_5147,In_2000,In_518);
and U5148 (N_5148,In_330,In_2496);
and U5149 (N_5149,In_69,In_1475);
or U5150 (N_5150,In_1851,In_1411);
nor U5151 (N_5151,In_2468,In_1079);
xnor U5152 (N_5152,In_2389,In_705);
or U5153 (N_5153,In_143,In_1971);
nand U5154 (N_5154,In_911,In_2214);
or U5155 (N_5155,In_1054,In_2176);
nand U5156 (N_5156,In_1079,In_621);
and U5157 (N_5157,In_784,In_2161);
nand U5158 (N_5158,In_1242,In_1672);
xnor U5159 (N_5159,In_1611,In_700);
or U5160 (N_5160,In_1966,In_1363);
nand U5161 (N_5161,In_628,In_2472);
xor U5162 (N_5162,In_2235,In_1575);
or U5163 (N_5163,In_252,In_934);
and U5164 (N_5164,In_494,In_1038);
or U5165 (N_5165,In_1630,In_1260);
nor U5166 (N_5166,In_1329,In_1747);
nand U5167 (N_5167,In_1910,In_782);
nor U5168 (N_5168,In_2249,In_1097);
and U5169 (N_5169,In_2379,In_1755);
nor U5170 (N_5170,In_490,In_2079);
xnor U5171 (N_5171,In_1139,In_560);
xnor U5172 (N_5172,In_470,In_1803);
and U5173 (N_5173,In_988,In_1014);
nand U5174 (N_5174,In_1360,In_732);
nor U5175 (N_5175,In_87,In_756);
nor U5176 (N_5176,In_301,In_629);
xnor U5177 (N_5177,In_1910,In_1280);
or U5178 (N_5178,In_70,In_1298);
nand U5179 (N_5179,In_2009,In_1859);
or U5180 (N_5180,In_1489,In_851);
or U5181 (N_5181,In_908,In_1799);
nor U5182 (N_5182,In_1216,In_889);
nand U5183 (N_5183,In_409,In_2157);
nand U5184 (N_5184,In_1566,In_1035);
nand U5185 (N_5185,In_1196,In_676);
and U5186 (N_5186,In_1954,In_291);
and U5187 (N_5187,In_1532,In_555);
nor U5188 (N_5188,In_891,In_1533);
xor U5189 (N_5189,In_527,In_1074);
nor U5190 (N_5190,In_398,In_2101);
or U5191 (N_5191,In_1737,In_1953);
nor U5192 (N_5192,In_888,In_1841);
nand U5193 (N_5193,In_362,In_1615);
nor U5194 (N_5194,In_2413,In_325);
nand U5195 (N_5195,In_1218,In_214);
and U5196 (N_5196,In_2149,In_1541);
nor U5197 (N_5197,In_1834,In_1629);
or U5198 (N_5198,In_1980,In_377);
xor U5199 (N_5199,In_42,In_1082);
xor U5200 (N_5200,In_1506,In_599);
or U5201 (N_5201,In_1381,In_2455);
nand U5202 (N_5202,In_765,In_789);
and U5203 (N_5203,In_1406,In_1118);
and U5204 (N_5204,In_1253,In_1421);
xor U5205 (N_5205,In_1330,In_831);
xnor U5206 (N_5206,In_588,In_896);
and U5207 (N_5207,In_2076,In_312);
xor U5208 (N_5208,In_1393,In_55);
nand U5209 (N_5209,In_862,In_692);
nand U5210 (N_5210,In_1297,In_778);
or U5211 (N_5211,In_476,In_90);
or U5212 (N_5212,In_2381,In_420);
nor U5213 (N_5213,In_273,In_1334);
nor U5214 (N_5214,In_2107,In_1472);
xnor U5215 (N_5215,In_1445,In_2486);
and U5216 (N_5216,In_288,In_1243);
nand U5217 (N_5217,In_1368,In_1443);
nor U5218 (N_5218,In_1234,In_2317);
and U5219 (N_5219,In_816,In_680);
or U5220 (N_5220,In_1717,In_2320);
nor U5221 (N_5221,In_1356,In_2020);
or U5222 (N_5222,In_1787,In_2374);
nor U5223 (N_5223,In_913,In_1189);
nor U5224 (N_5224,In_2491,In_2477);
or U5225 (N_5225,In_1648,In_1091);
nor U5226 (N_5226,In_1640,In_530);
and U5227 (N_5227,In_270,In_1919);
xor U5228 (N_5228,In_1720,In_879);
xor U5229 (N_5229,In_920,In_1969);
or U5230 (N_5230,In_902,In_1961);
nor U5231 (N_5231,In_868,In_1974);
or U5232 (N_5232,In_2216,In_1572);
nand U5233 (N_5233,In_746,In_596);
xor U5234 (N_5234,In_506,In_2187);
and U5235 (N_5235,In_619,In_2460);
nand U5236 (N_5236,In_1788,In_749);
or U5237 (N_5237,In_2411,In_799);
xnor U5238 (N_5238,In_941,In_456);
or U5239 (N_5239,In_2386,In_2356);
and U5240 (N_5240,In_1678,In_2461);
or U5241 (N_5241,In_920,In_1795);
nor U5242 (N_5242,In_2497,In_145);
and U5243 (N_5243,In_1055,In_1371);
nor U5244 (N_5244,In_3,In_1481);
xor U5245 (N_5245,In_378,In_1938);
nand U5246 (N_5246,In_495,In_2018);
and U5247 (N_5247,In_2231,In_1089);
and U5248 (N_5248,In_2109,In_2046);
and U5249 (N_5249,In_2033,In_1771);
or U5250 (N_5250,In_406,In_1069);
or U5251 (N_5251,In_1331,In_488);
nand U5252 (N_5252,In_1318,In_1599);
nor U5253 (N_5253,In_505,In_1541);
nor U5254 (N_5254,In_668,In_114);
or U5255 (N_5255,In_531,In_333);
xnor U5256 (N_5256,In_1730,In_1446);
nor U5257 (N_5257,In_872,In_161);
xnor U5258 (N_5258,In_174,In_735);
nor U5259 (N_5259,In_748,In_1451);
nand U5260 (N_5260,In_2448,In_163);
and U5261 (N_5261,In_351,In_74);
xor U5262 (N_5262,In_535,In_1442);
and U5263 (N_5263,In_738,In_846);
nand U5264 (N_5264,In_114,In_1941);
nor U5265 (N_5265,In_1430,In_910);
or U5266 (N_5266,In_1805,In_950);
and U5267 (N_5267,In_2374,In_1134);
and U5268 (N_5268,In_2099,In_837);
and U5269 (N_5269,In_1831,In_1363);
and U5270 (N_5270,In_1445,In_187);
nor U5271 (N_5271,In_1230,In_1893);
xor U5272 (N_5272,In_1162,In_934);
nand U5273 (N_5273,In_1843,In_2295);
or U5274 (N_5274,In_2105,In_1944);
or U5275 (N_5275,In_1072,In_366);
and U5276 (N_5276,In_971,In_144);
and U5277 (N_5277,In_1766,In_461);
nor U5278 (N_5278,In_1002,In_198);
xnor U5279 (N_5279,In_796,In_1305);
and U5280 (N_5280,In_854,In_1978);
and U5281 (N_5281,In_691,In_2145);
and U5282 (N_5282,In_1745,In_1435);
nor U5283 (N_5283,In_1193,In_112);
or U5284 (N_5284,In_82,In_1579);
nor U5285 (N_5285,In_342,In_1628);
nor U5286 (N_5286,In_1575,In_884);
and U5287 (N_5287,In_563,In_1246);
and U5288 (N_5288,In_2390,In_2101);
nand U5289 (N_5289,In_1798,In_2100);
nand U5290 (N_5290,In_473,In_1754);
nor U5291 (N_5291,In_1064,In_51);
xnor U5292 (N_5292,In_810,In_1376);
nor U5293 (N_5293,In_1600,In_1375);
nand U5294 (N_5294,In_404,In_298);
xnor U5295 (N_5295,In_1407,In_674);
nand U5296 (N_5296,In_1494,In_503);
nand U5297 (N_5297,In_763,In_50);
and U5298 (N_5298,In_2118,In_1654);
and U5299 (N_5299,In_539,In_1596);
nand U5300 (N_5300,In_1563,In_1771);
nor U5301 (N_5301,In_89,In_2133);
or U5302 (N_5302,In_1258,In_2169);
or U5303 (N_5303,In_2481,In_1631);
or U5304 (N_5304,In_1362,In_378);
or U5305 (N_5305,In_505,In_1773);
xor U5306 (N_5306,In_1536,In_818);
and U5307 (N_5307,In_1740,In_1546);
nor U5308 (N_5308,In_996,In_2458);
or U5309 (N_5309,In_2091,In_2079);
xor U5310 (N_5310,In_475,In_2230);
nor U5311 (N_5311,In_782,In_265);
and U5312 (N_5312,In_563,In_221);
and U5313 (N_5313,In_794,In_1509);
nor U5314 (N_5314,In_37,In_2086);
and U5315 (N_5315,In_1177,In_1439);
and U5316 (N_5316,In_874,In_1632);
nor U5317 (N_5317,In_2381,In_2208);
nor U5318 (N_5318,In_528,In_459);
xnor U5319 (N_5319,In_2238,In_1258);
or U5320 (N_5320,In_1522,In_2049);
nor U5321 (N_5321,In_2421,In_782);
xnor U5322 (N_5322,In_1575,In_670);
nand U5323 (N_5323,In_723,In_1767);
and U5324 (N_5324,In_187,In_1611);
xor U5325 (N_5325,In_1086,In_329);
and U5326 (N_5326,In_1716,In_1961);
and U5327 (N_5327,In_1074,In_2330);
nor U5328 (N_5328,In_2311,In_1576);
nand U5329 (N_5329,In_905,In_2174);
or U5330 (N_5330,In_682,In_1300);
and U5331 (N_5331,In_844,In_1474);
xnor U5332 (N_5332,In_2261,In_121);
or U5333 (N_5333,In_216,In_2336);
or U5334 (N_5334,In_773,In_671);
nand U5335 (N_5335,In_2359,In_178);
or U5336 (N_5336,In_1096,In_165);
and U5337 (N_5337,In_805,In_2463);
nand U5338 (N_5338,In_319,In_1633);
and U5339 (N_5339,In_1682,In_1747);
nor U5340 (N_5340,In_1473,In_359);
or U5341 (N_5341,In_2041,In_1027);
nor U5342 (N_5342,In_2113,In_2213);
and U5343 (N_5343,In_2330,In_2112);
xor U5344 (N_5344,In_1004,In_1626);
xnor U5345 (N_5345,In_2471,In_2011);
nand U5346 (N_5346,In_288,In_1205);
nand U5347 (N_5347,In_946,In_1787);
and U5348 (N_5348,In_997,In_1950);
xnor U5349 (N_5349,In_1314,In_1787);
or U5350 (N_5350,In_1610,In_1186);
or U5351 (N_5351,In_250,In_1047);
nor U5352 (N_5352,In_487,In_1402);
nand U5353 (N_5353,In_527,In_1220);
and U5354 (N_5354,In_2250,In_1121);
and U5355 (N_5355,In_666,In_783);
xnor U5356 (N_5356,In_1646,In_968);
and U5357 (N_5357,In_2254,In_1052);
or U5358 (N_5358,In_790,In_137);
nor U5359 (N_5359,In_510,In_1658);
xnor U5360 (N_5360,In_17,In_1319);
nor U5361 (N_5361,In_480,In_2345);
xor U5362 (N_5362,In_432,In_1916);
xnor U5363 (N_5363,In_744,In_1914);
nor U5364 (N_5364,In_1292,In_1396);
xor U5365 (N_5365,In_489,In_1923);
or U5366 (N_5366,In_2335,In_2341);
and U5367 (N_5367,In_578,In_1914);
nor U5368 (N_5368,In_1694,In_1193);
nor U5369 (N_5369,In_1828,In_1990);
nor U5370 (N_5370,In_1811,In_1186);
nor U5371 (N_5371,In_802,In_1167);
or U5372 (N_5372,In_1095,In_1089);
nor U5373 (N_5373,In_571,In_901);
nand U5374 (N_5374,In_2067,In_1959);
xnor U5375 (N_5375,In_346,In_1270);
nand U5376 (N_5376,In_695,In_736);
xor U5377 (N_5377,In_1263,In_888);
or U5378 (N_5378,In_1964,In_195);
and U5379 (N_5379,In_2347,In_1804);
or U5380 (N_5380,In_199,In_1972);
nand U5381 (N_5381,In_1688,In_904);
or U5382 (N_5382,In_1497,In_1217);
xor U5383 (N_5383,In_1886,In_1943);
or U5384 (N_5384,In_677,In_1478);
xnor U5385 (N_5385,In_363,In_1353);
nor U5386 (N_5386,In_2097,In_1222);
or U5387 (N_5387,In_1919,In_1763);
nor U5388 (N_5388,In_352,In_1360);
nor U5389 (N_5389,In_2383,In_666);
or U5390 (N_5390,In_1352,In_2039);
nor U5391 (N_5391,In_2339,In_826);
xnor U5392 (N_5392,In_1763,In_1080);
nand U5393 (N_5393,In_1208,In_261);
and U5394 (N_5394,In_566,In_1422);
xor U5395 (N_5395,In_721,In_1841);
nor U5396 (N_5396,In_228,In_2261);
xnor U5397 (N_5397,In_163,In_1515);
xnor U5398 (N_5398,In_114,In_327);
nor U5399 (N_5399,In_772,In_521);
and U5400 (N_5400,In_835,In_1764);
or U5401 (N_5401,In_2283,In_240);
and U5402 (N_5402,In_922,In_340);
and U5403 (N_5403,In_2336,In_2160);
xor U5404 (N_5404,In_1475,In_2370);
or U5405 (N_5405,In_1568,In_694);
nand U5406 (N_5406,In_1262,In_2002);
nor U5407 (N_5407,In_246,In_2449);
and U5408 (N_5408,In_692,In_666);
or U5409 (N_5409,In_2074,In_1347);
xnor U5410 (N_5410,In_523,In_263);
and U5411 (N_5411,In_550,In_492);
and U5412 (N_5412,In_1561,In_496);
or U5413 (N_5413,In_1214,In_1034);
and U5414 (N_5414,In_2015,In_1137);
nand U5415 (N_5415,In_274,In_441);
and U5416 (N_5416,In_1644,In_2067);
nor U5417 (N_5417,In_868,In_2067);
xnor U5418 (N_5418,In_452,In_37);
nand U5419 (N_5419,In_954,In_103);
or U5420 (N_5420,In_2217,In_324);
xor U5421 (N_5421,In_48,In_598);
nor U5422 (N_5422,In_1670,In_284);
nand U5423 (N_5423,In_663,In_2160);
or U5424 (N_5424,In_856,In_348);
nor U5425 (N_5425,In_2281,In_451);
and U5426 (N_5426,In_2240,In_1965);
nand U5427 (N_5427,In_970,In_1823);
or U5428 (N_5428,In_917,In_1267);
nor U5429 (N_5429,In_1779,In_1553);
nor U5430 (N_5430,In_1169,In_1694);
xor U5431 (N_5431,In_2410,In_1588);
or U5432 (N_5432,In_2393,In_1258);
nor U5433 (N_5433,In_485,In_1256);
xor U5434 (N_5434,In_1777,In_2308);
xor U5435 (N_5435,In_815,In_2455);
nand U5436 (N_5436,In_281,In_2305);
nand U5437 (N_5437,In_799,In_66);
xor U5438 (N_5438,In_2335,In_324);
and U5439 (N_5439,In_1511,In_41);
nand U5440 (N_5440,In_1293,In_1009);
or U5441 (N_5441,In_1931,In_337);
nand U5442 (N_5442,In_1982,In_0);
and U5443 (N_5443,In_231,In_2373);
and U5444 (N_5444,In_1766,In_1629);
xnor U5445 (N_5445,In_1491,In_2090);
nor U5446 (N_5446,In_1281,In_1347);
nand U5447 (N_5447,In_1945,In_1504);
or U5448 (N_5448,In_276,In_692);
nor U5449 (N_5449,In_231,In_1630);
nand U5450 (N_5450,In_1104,In_1968);
nand U5451 (N_5451,In_1698,In_1002);
nor U5452 (N_5452,In_2098,In_1363);
xnor U5453 (N_5453,In_2165,In_2347);
or U5454 (N_5454,In_1694,In_203);
nor U5455 (N_5455,In_608,In_904);
or U5456 (N_5456,In_819,In_1679);
or U5457 (N_5457,In_1597,In_2274);
xnor U5458 (N_5458,In_1050,In_1869);
nand U5459 (N_5459,In_1282,In_1897);
nor U5460 (N_5460,In_253,In_921);
or U5461 (N_5461,In_36,In_2322);
nor U5462 (N_5462,In_1813,In_1831);
nand U5463 (N_5463,In_1283,In_315);
xnor U5464 (N_5464,In_2307,In_1557);
nor U5465 (N_5465,In_2412,In_2375);
and U5466 (N_5466,In_719,In_98);
and U5467 (N_5467,In_71,In_1238);
xnor U5468 (N_5468,In_298,In_2169);
and U5469 (N_5469,In_2432,In_1544);
or U5470 (N_5470,In_2067,In_1979);
nor U5471 (N_5471,In_140,In_556);
nand U5472 (N_5472,In_334,In_1222);
or U5473 (N_5473,In_1377,In_448);
and U5474 (N_5474,In_1283,In_1457);
nand U5475 (N_5475,In_2070,In_1579);
xnor U5476 (N_5476,In_1253,In_2062);
and U5477 (N_5477,In_351,In_1922);
nand U5478 (N_5478,In_1614,In_144);
and U5479 (N_5479,In_1781,In_1618);
and U5480 (N_5480,In_1504,In_800);
xor U5481 (N_5481,In_664,In_927);
nand U5482 (N_5482,In_2247,In_2131);
xnor U5483 (N_5483,In_995,In_777);
xnor U5484 (N_5484,In_127,In_1872);
xnor U5485 (N_5485,In_181,In_2424);
xnor U5486 (N_5486,In_2295,In_1105);
and U5487 (N_5487,In_2219,In_660);
nor U5488 (N_5488,In_775,In_301);
nand U5489 (N_5489,In_76,In_802);
nand U5490 (N_5490,In_2202,In_76);
xor U5491 (N_5491,In_1079,In_2114);
nor U5492 (N_5492,In_2404,In_1604);
or U5493 (N_5493,In_1870,In_1392);
nor U5494 (N_5494,In_294,In_1175);
or U5495 (N_5495,In_1903,In_1571);
xnor U5496 (N_5496,In_117,In_509);
nor U5497 (N_5497,In_1957,In_1449);
xnor U5498 (N_5498,In_2276,In_2096);
nor U5499 (N_5499,In_172,In_1919);
xor U5500 (N_5500,In_1858,In_664);
or U5501 (N_5501,In_1687,In_2328);
nor U5502 (N_5502,In_1758,In_1678);
nor U5503 (N_5503,In_376,In_505);
and U5504 (N_5504,In_713,In_2117);
nor U5505 (N_5505,In_1741,In_1073);
or U5506 (N_5506,In_1660,In_108);
nor U5507 (N_5507,In_1877,In_889);
xor U5508 (N_5508,In_947,In_886);
or U5509 (N_5509,In_450,In_1392);
or U5510 (N_5510,In_751,In_616);
nor U5511 (N_5511,In_1615,In_1275);
xnor U5512 (N_5512,In_656,In_1822);
and U5513 (N_5513,In_1262,In_1531);
nand U5514 (N_5514,In_56,In_2282);
and U5515 (N_5515,In_1243,In_1103);
nor U5516 (N_5516,In_402,In_195);
and U5517 (N_5517,In_2496,In_680);
and U5518 (N_5518,In_2182,In_1438);
and U5519 (N_5519,In_1801,In_874);
nor U5520 (N_5520,In_465,In_1603);
and U5521 (N_5521,In_2176,In_37);
nor U5522 (N_5522,In_2010,In_1692);
and U5523 (N_5523,In_1205,In_1985);
or U5524 (N_5524,In_915,In_1496);
xor U5525 (N_5525,In_793,In_1098);
nor U5526 (N_5526,In_566,In_2321);
nand U5527 (N_5527,In_1633,In_791);
nor U5528 (N_5528,In_725,In_2018);
nand U5529 (N_5529,In_808,In_1393);
nor U5530 (N_5530,In_1865,In_66);
or U5531 (N_5531,In_100,In_305);
or U5532 (N_5532,In_1869,In_218);
or U5533 (N_5533,In_1,In_2277);
and U5534 (N_5534,In_993,In_483);
nand U5535 (N_5535,In_1657,In_1765);
nand U5536 (N_5536,In_1013,In_1762);
nand U5537 (N_5537,In_1549,In_547);
nor U5538 (N_5538,In_512,In_608);
xor U5539 (N_5539,In_1580,In_419);
nor U5540 (N_5540,In_1502,In_1302);
xor U5541 (N_5541,In_2042,In_1429);
xor U5542 (N_5542,In_744,In_1060);
or U5543 (N_5543,In_747,In_2038);
and U5544 (N_5544,In_100,In_542);
and U5545 (N_5545,In_2016,In_1457);
or U5546 (N_5546,In_547,In_976);
xnor U5547 (N_5547,In_207,In_971);
or U5548 (N_5548,In_2396,In_656);
xor U5549 (N_5549,In_551,In_55);
and U5550 (N_5550,In_103,In_1111);
nand U5551 (N_5551,In_2231,In_2364);
xnor U5552 (N_5552,In_999,In_1697);
and U5553 (N_5553,In_2389,In_1110);
or U5554 (N_5554,In_1061,In_2002);
xor U5555 (N_5555,In_215,In_629);
or U5556 (N_5556,In_916,In_1559);
nand U5557 (N_5557,In_1749,In_728);
or U5558 (N_5558,In_2276,In_465);
nand U5559 (N_5559,In_1963,In_1730);
xnor U5560 (N_5560,In_1896,In_126);
nor U5561 (N_5561,In_2052,In_18);
or U5562 (N_5562,In_1334,In_1203);
nand U5563 (N_5563,In_1706,In_817);
and U5564 (N_5564,In_462,In_2034);
and U5565 (N_5565,In_1411,In_1700);
nor U5566 (N_5566,In_2072,In_808);
nand U5567 (N_5567,In_1398,In_853);
nand U5568 (N_5568,In_2171,In_1009);
or U5569 (N_5569,In_253,In_2340);
and U5570 (N_5570,In_1682,In_972);
xor U5571 (N_5571,In_1708,In_507);
or U5572 (N_5572,In_1688,In_783);
and U5573 (N_5573,In_1263,In_353);
or U5574 (N_5574,In_1453,In_529);
xnor U5575 (N_5575,In_286,In_2186);
and U5576 (N_5576,In_1272,In_2159);
or U5577 (N_5577,In_1501,In_643);
xnor U5578 (N_5578,In_1787,In_158);
nor U5579 (N_5579,In_1946,In_2498);
nor U5580 (N_5580,In_1617,In_807);
nand U5581 (N_5581,In_2349,In_188);
and U5582 (N_5582,In_1213,In_424);
and U5583 (N_5583,In_1442,In_1080);
xor U5584 (N_5584,In_395,In_2464);
nand U5585 (N_5585,In_1700,In_887);
nor U5586 (N_5586,In_1161,In_1175);
nand U5587 (N_5587,In_1502,In_1070);
or U5588 (N_5588,In_1397,In_1231);
xnor U5589 (N_5589,In_1505,In_1063);
nor U5590 (N_5590,In_2325,In_1386);
and U5591 (N_5591,In_1233,In_876);
xnor U5592 (N_5592,In_875,In_341);
or U5593 (N_5593,In_2463,In_2259);
xor U5594 (N_5594,In_1553,In_1717);
xor U5595 (N_5595,In_823,In_413);
nand U5596 (N_5596,In_2048,In_2388);
or U5597 (N_5597,In_398,In_2250);
xor U5598 (N_5598,In_1434,In_1680);
nand U5599 (N_5599,In_1542,In_2008);
and U5600 (N_5600,In_1847,In_379);
nor U5601 (N_5601,In_1163,In_778);
xnor U5602 (N_5602,In_772,In_598);
xnor U5603 (N_5603,In_411,In_2270);
or U5604 (N_5604,In_2485,In_1284);
or U5605 (N_5605,In_1966,In_1579);
xnor U5606 (N_5606,In_1805,In_2);
nor U5607 (N_5607,In_931,In_2324);
nor U5608 (N_5608,In_594,In_914);
nor U5609 (N_5609,In_1452,In_2225);
or U5610 (N_5610,In_1577,In_1894);
xor U5611 (N_5611,In_1352,In_12);
nand U5612 (N_5612,In_1852,In_509);
and U5613 (N_5613,In_2073,In_2442);
xnor U5614 (N_5614,In_508,In_2450);
xor U5615 (N_5615,In_2159,In_1699);
and U5616 (N_5616,In_1338,In_2416);
xnor U5617 (N_5617,In_2160,In_563);
or U5618 (N_5618,In_2267,In_1677);
nand U5619 (N_5619,In_56,In_2395);
xor U5620 (N_5620,In_935,In_2257);
xnor U5621 (N_5621,In_2380,In_1568);
xnor U5622 (N_5622,In_884,In_2336);
nor U5623 (N_5623,In_447,In_2423);
nor U5624 (N_5624,In_738,In_812);
xor U5625 (N_5625,In_1619,In_2248);
or U5626 (N_5626,In_2202,In_2446);
or U5627 (N_5627,In_184,In_1584);
xor U5628 (N_5628,In_1047,In_2060);
xnor U5629 (N_5629,In_428,In_1918);
xor U5630 (N_5630,In_200,In_1352);
and U5631 (N_5631,In_325,In_1689);
nor U5632 (N_5632,In_1919,In_2357);
xor U5633 (N_5633,In_632,In_652);
and U5634 (N_5634,In_2326,In_364);
or U5635 (N_5635,In_560,In_778);
or U5636 (N_5636,In_1574,In_790);
or U5637 (N_5637,In_210,In_361);
nor U5638 (N_5638,In_908,In_2207);
or U5639 (N_5639,In_2294,In_619);
and U5640 (N_5640,In_815,In_607);
xnor U5641 (N_5641,In_2049,In_2193);
and U5642 (N_5642,In_908,In_61);
or U5643 (N_5643,In_1260,In_80);
and U5644 (N_5644,In_2199,In_427);
xor U5645 (N_5645,In_1822,In_72);
nand U5646 (N_5646,In_2482,In_2480);
nand U5647 (N_5647,In_1069,In_2431);
nor U5648 (N_5648,In_818,In_500);
xor U5649 (N_5649,In_168,In_2463);
nor U5650 (N_5650,In_2371,In_2077);
or U5651 (N_5651,In_1312,In_2178);
xor U5652 (N_5652,In_891,In_1369);
and U5653 (N_5653,In_779,In_1476);
and U5654 (N_5654,In_200,In_1673);
and U5655 (N_5655,In_1857,In_58);
and U5656 (N_5656,In_1876,In_1267);
and U5657 (N_5657,In_789,In_1256);
nor U5658 (N_5658,In_1067,In_1695);
nor U5659 (N_5659,In_1919,In_1368);
nor U5660 (N_5660,In_63,In_568);
and U5661 (N_5661,In_674,In_1535);
or U5662 (N_5662,In_1677,In_737);
and U5663 (N_5663,In_538,In_798);
nor U5664 (N_5664,In_2093,In_1560);
or U5665 (N_5665,In_85,In_52);
nand U5666 (N_5666,In_693,In_38);
or U5667 (N_5667,In_1778,In_1275);
nor U5668 (N_5668,In_1981,In_2337);
xnor U5669 (N_5669,In_2309,In_273);
and U5670 (N_5670,In_1734,In_1954);
or U5671 (N_5671,In_1001,In_2332);
and U5672 (N_5672,In_912,In_697);
xnor U5673 (N_5673,In_962,In_2245);
nand U5674 (N_5674,In_2080,In_1721);
and U5675 (N_5675,In_397,In_841);
xor U5676 (N_5676,In_545,In_611);
and U5677 (N_5677,In_650,In_175);
nand U5678 (N_5678,In_2319,In_2429);
nor U5679 (N_5679,In_1525,In_1605);
and U5680 (N_5680,In_1212,In_1245);
or U5681 (N_5681,In_1280,In_486);
or U5682 (N_5682,In_1650,In_2309);
xor U5683 (N_5683,In_2250,In_1756);
and U5684 (N_5684,In_486,In_1694);
nor U5685 (N_5685,In_1613,In_1072);
nand U5686 (N_5686,In_1414,In_1369);
nand U5687 (N_5687,In_635,In_626);
xor U5688 (N_5688,In_1163,In_353);
nor U5689 (N_5689,In_26,In_391);
and U5690 (N_5690,In_1067,In_1383);
nor U5691 (N_5691,In_858,In_1021);
nand U5692 (N_5692,In_275,In_2148);
nand U5693 (N_5693,In_1901,In_365);
and U5694 (N_5694,In_2335,In_1428);
or U5695 (N_5695,In_4,In_332);
and U5696 (N_5696,In_422,In_116);
nor U5697 (N_5697,In_516,In_1349);
nand U5698 (N_5698,In_1270,In_2389);
nor U5699 (N_5699,In_1961,In_851);
nand U5700 (N_5700,In_2414,In_74);
xnor U5701 (N_5701,In_1623,In_237);
and U5702 (N_5702,In_1177,In_261);
nand U5703 (N_5703,In_956,In_2157);
nor U5704 (N_5704,In_1159,In_303);
or U5705 (N_5705,In_1767,In_1954);
or U5706 (N_5706,In_434,In_812);
nor U5707 (N_5707,In_783,In_1780);
and U5708 (N_5708,In_1271,In_1792);
nor U5709 (N_5709,In_162,In_179);
xnor U5710 (N_5710,In_728,In_1179);
or U5711 (N_5711,In_1890,In_2186);
or U5712 (N_5712,In_567,In_640);
nor U5713 (N_5713,In_1489,In_2134);
nor U5714 (N_5714,In_696,In_2236);
or U5715 (N_5715,In_2104,In_2495);
nor U5716 (N_5716,In_2215,In_391);
nand U5717 (N_5717,In_166,In_1442);
and U5718 (N_5718,In_824,In_1865);
and U5719 (N_5719,In_1832,In_1209);
nand U5720 (N_5720,In_1754,In_1015);
xnor U5721 (N_5721,In_1666,In_1975);
nor U5722 (N_5722,In_294,In_128);
nand U5723 (N_5723,In_2290,In_1301);
nand U5724 (N_5724,In_126,In_1653);
xnor U5725 (N_5725,In_1161,In_1638);
nor U5726 (N_5726,In_2105,In_624);
nor U5727 (N_5727,In_417,In_700);
xnor U5728 (N_5728,In_156,In_1984);
nand U5729 (N_5729,In_1979,In_1414);
and U5730 (N_5730,In_1024,In_1758);
nor U5731 (N_5731,In_200,In_1369);
or U5732 (N_5732,In_959,In_2197);
nor U5733 (N_5733,In_113,In_1861);
or U5734 (N_5734,In_533,In_460);
nand U5735 (N_5735,In_1079,In_972);
nand U5736 (N_5736,In_2484,In_1000);
and U5737 (N_5737,In_118,In_838);
and U5738 (N_5738,In_851,In_2356);
and U5739 (N_5739,In_1473,In_1127);
or U5740 (N_5740,In_171,In_1941);
nor U5741 (N_5741,In_2119,In_2188);
nand U5742 (N_5742,In_1354,In_1599);
xnor U5743 (N_5743,In_1943,In_450);
nand U5744 (N_5744,In_368,In_739);
and U5745 (N_5745,In_1987,In_1813);
xnor U5746 (N_5746,In_88,In_506);
nor U5747 (N_5747,In_1759,In_1528);
nor U5748 (N_5748,In_190,In_2384);
or U5749 (N_5749,In_1210,In_458);
xor U5750 (N_5750,In_695,In_711);
nand U5751 (N_5751,In_277,In_2316);
nand U5752 (N_5752,In_276,In_318);
nor U5753 (N_5753,In_1651,In_558);
nor U5754 (N_5754,In_2172,In_2451);
nand U5755 (N_5755,In_61,In_1946);
nand U5756 (N_5756,In_281,In_433);
nand U5757 (N_5757,In_1641,In_2041);
nor U5758 (N_5758,In_657,In_600);
nand U5759 (N_5759,In_597,In_2);
nor U5760 (N_5760,In_2177,In_1195);
and U5761 (N_5761,In_774,In_1916);
and U5762 (N_5762,In_1457,In_690);
or U5763 (N_5763,In_2160,In_151);
xnor U5764 (N_5764,In_1372,In_2269);
nand U5765 (N_5765,In_382,In_2134);
xor U5766 (N_5766,In_2254,In_1612);
nor U5767 (N_5767,In_1282,In_306);
nor U5768 (N_5768,In_215,In_715);
nand U5769 (N_5769,In_59,In_1964);
nor U5770 (N_5770,In_705,In_1151);
xnor U5771 (N_5771,In_2147,In_680);
and U5772 (N_5772,In_2418,In_612);
xor U5773 (N_5773,In_1418,In_2449);
xor U5774 (N_5774,In_2248,In_2063);
or U5775 (N_5775,In_2356,In_1191);
xor U5776 (N_5776,In_1440,In_47);
and U5777 (N_5777,In_2348,In_2322);
nor U5778 (N_5778,In_329,In_999);
nand U5779 (N_5779,In_1854,In_2263);
and U5780 (N_5780,In_1865,In_2074);
xor U5781 (N_5781,In_526,In_1680);
nor U5782 (N_5782,In_1568,In_1129);
nand U5783 (N_5783,In_1498,In_1856);
xnor U5784 (N_5784,In_1994,In_2410);
xor U5785 (N_5785,In_395,In_648);
and U5786 (N_5786,In_1010,In_1191);
or U5787 (N_5787,In_1622,In_131);
or U5788 (N_5788,In_2091,In_2397);
xnor U5789 (N_5789,In_954,In_2195);
and U5790 (N_5790,In_1495,In_2017);
and U5791 (N_5791,In_1132,In_65);
nand U5792 (N_5792,In_258,In_1046);
or U5793 (N_5793,In_274,In_1569);
or U5794 (N_5794,In_837,In_1705);
or U5795 (N_5795,In_0,In_2255);
or U5796 (N_5796,In_52,In_1589);
nand U5797 (N_5797,In_1079,In_1891);
and U5798 (N_5798,In_1770,In_93);
nand U5799 (N_5799,In_1403,In_184);
nor U5800 (N_5800,In_152,In_1881);
nand U5801 (N_5801,In_1569,In_1321);
nor U5802 (N_5802,In_1488,In_965);
nor U5803 (N_5803,In_472,In_679);
or U5804 (N_5804,In_17,In_361);
xor U5805 (N_5805,In_617,In_1365);
or U5806 (N_5806,In_287,In_898);
and U5807 (N_5807,In_2069,In_859);
or U5808 (N_5808,In_637,In_73);
nand U5809 (N_5809,In_1349,In_1347);
nor U5810 (N_5810,In_867,In_687);
nand U5811 (N_5811,In_2072,In_1776);
and U5812 (N_5812,In_1407,In_16);
xor U5813 (N_5813,In_875,In_1660);
nand U5814 (N_5814,In_1638,In_1690);
nor U5815 (N_5815,In_214,In_108);
nand U5816 (N_5816,In_2107,In_1001);
xnor U5817 (N_5817,In_216,In_1106);
and U5818 (N_5818,In_1568,In_1978);
and U5819 (N_5819,In_957,In_2255);
nor U5820 (N_5820,In_2269,In_1140);
and U5821 (N_5821,In_1140,In_2311);
nor U5822 (N_5822,In_629,In_1048);
nand U5823 (N_5823,In_296,In_71);
nor U5824 (N_5824,In_520,In_1188);
and U5825 (N_5825,In_1273,In_361);
and U5826 (N_5826,In_1306,In_2272);
or U5827 (N_5827,In_1301,In_1665);
or U5828 (N_5828,In_1985,In_196);
and U5829 (N_5829,In_490,In_440);
nand U5830 (N_5830,In_2165,In_1943);
nor U5831 (N_5831,In_1483,In_924);
nand U5832 (N_5832,In_692,In_979);
xor U5833 (N_5833,In_650,In_2464);
nand U5834 (N_5834,In_1657,In_1382);
nor U5835 (N_5835,In_2319,In_378);
or U5836 (N_5836,In_1241,In_2113);
and U5837 (N_5837,In_1818,In_128);
or U5838 (N_5838,In_137,In_1502);
nand U5839 (N_5839,In_143,In_2327);
xor U5840 (N_5840,In_347,In_1);
or U5841 (N_5841,In_1578,In_1977);
nand U5842 (N_5842,In_717,In_905);
xor U5843 (N_5843,In_723,In_1770);
and U5844 (N_5844,In_1015,In_1293);
and U5845 (N_5845,In_1943,In_260);
nor U5846 (N_5846,In_1504,In_2251);
or U5847 (N_5847,In_104,In_809);
nor U5848 (N_5848,In_1238,In_1853);
and U5849 (N_5849,In_1312,In_2094);
and U5850 (N_5850,In_1256,In_611);
nor U5851 (N_5851,In_475,In_1129);
xor U5852 (N_5852,In_1800,In_1753);
and U5853 (N_5853,In_1282,In_1808);
xor U5854 (N_5854,In_1325,In_1478);
nor U5855 (N_5855,In_1520,In_2017);
xnor U5856 (N_5856,In_1911,In_1523);
and U5857 (N_5857,In_457,In_1293);
or U5858 (N_5858,In_2430,In_1320);
nor U5859 (N_5859,In_1504,In_1041);
and U5860 (N_5860,In_583,In_841);
and U5861 (N_5861,In_505,In_1196);
nand U5862 (N_5862,In_1997,In_1705);
nor U5863 (N_5863,In_528,In_170);
or U5864 (N_5864,In_1223,In_1114);
and U5865 (N_5865,In_2265,In_2393);
nor U5866 (N_5866,In_1824,In_2152);
xor U5867 (N_5867,In_2480,In_412);
or U5868 (N_5868,In_280,In_257);
or U5869 (N_5869,In_805,In_1990);
nand U5870 (N_5870,In_967,In_1199);
nand U5871 (N_5871,In_838,In_249);
or U5872 (N_5872,In_1573,In_457);
nand U5873 (N_5873,In_1318,In_2039);
or U5874 (N_5874,In_1956,In_1105);
and U5875 (N_5875,In_2472,In_402);
nand U5876 (N_5876,In_2272,In_762);
or U5877 (N_5877,In_1545,In_839);
nor U5878 (N_5878,In_2279,In_384);
or U5879 (N_5879,In_499,In_2283);
nand U5880 (N_5880,In_2210,In_1359);
xor U5881 (N_5881,In_359,In_350);
nor U5882 (N_5882,In_1928,In_2428);
and U5883 (N_5883,In_298,In_1717);
nand U5884 (N_5884,In_1177,In_75);
xnor U5885 (N_5885,In_1762,In_1027);
xor U5886 (N_5886,In_1804,In_478);
nand U5887 (N_5887,In_647,In_1646);
nand U5888 (N_5888,In_681,In_2310);
or U5889 (N_5889,In_298,In_486);
or U5890 (N_5890,In_1294,In_1747);
nor U5891 (N_5891,In_2286,In_2218);
nand U5892 (N_5892,In_120,In_520);
nand U5893 (N_5893,In_763,In_1822);
nor U5894 (N_5894,In_844,In_2363);
and U5895 (N_5895,In_1357,In_1484);
xnor U5896 (N_5896,In_1522,In_473);
nor U5897 (N_5897,In_2078,In_595);
and U5898 (N_5898,In_1285,In_2088);
nand U5899 (N_5899,In_1272,In_575);
nor U5900 (N_5900,In_252,In_2403);
and U5901 (N_5901,In_1966,In_1613);
and U5902 (N_5902,In_271,In_605);
or U5903 (N_5903,In_1337,In_1945);
and U5904 (N_5904,In_2092,In_628);
xnor U5905 (N_5905,In_1066,In_1918);
or U5906 (N_5906,In_2357,In_63);
and U5907 (N_5907,In_620,In_751);
or U5908 (N_5908,In_372,In_2121);
nand U5909 (N_5909,In_2272,In_1959);
and U5910 (N_5910,In_1448,In_529);
xor U5911 (N_5911,In_309,In_1444);
nand U5912 (N_5912,In_1943,In_172);
or U5913 (N_5913,In_312,In_1423);
nand U5914 (N_5914,In_2001,In_2291);
and U5915 (N_5915,In_1950,In_2491);
nor U5916 (N_5916,In_496,In_1936);
or U5917 (N_5917,In_60,In_951);
nand U5918 (N_5918,In_1667,In_608);
xor U5919 (N_5919,In_1072,In_1280);
nand U5920 (N_5920,In_1452,In_534);
or U5921 (N_5921,In_999,In_41);
or U5922 (N_5922,In_1275,In_2119);
nor U5923 (N_5923,In_1416,In_656);
or U5924 (N_5924,In_1071,In_720);
and U5925 (N_5925,In_527,In_1030);
and U5926 (N_5926,In_2391,In_1981);
xnor U5927 (N_5927,In_122,In_1918);
nand U5928 (N_5928,In_2393,In_888);
or U5929 (N_5929,In_1969,In_705);
and U5930 (N_5930,In_2096,In_1477);
xor U5931 (N_5931,In_1733,In_1812);
xnor U5932 (N_5932,In_147,In_1253);
nand U5933 (N_5933,In_1948,In_1804);
and U5934 (N_5934,In_66,In_358);
xnor U5935 (N_5935,In_2178,In_2137);
nand U5936 (N_5936,In_819,In_1284);
xnor U5937 (N_5937,In_1212,In_285);
xnor U5938 (N_5938,In_1678,In_773);
and U5939 (N_5939,In_378,In_1281);
and U5940 (N_5940,In_1591,In_143);
or U5941 (N_5941,In_979,In_961);
or U5942 (N_5942,In_288,In_1097);
nand U5943 (N_5943,In_64,In_2276);
and U5944 (N_5944,In_1387,In_331);
xor U5945 (N_5945,In_902,In_703);
or U5946 (N_5946,In_1833,In_1581);
nor U5947 (N_5947,In_1753,In_262);
nor U5948 (N_5948,In_73,In_1757);
xnor U5949 (N_5949,In_2233,In_1995);
and U5950 (N_5950,In_2276,In_1635);
or U5951 (N_5951,In_1758,In_2054);
nand U5952 (N_5952,In_1539,In_973);
nand U5953 (N_5953,In_2466,In_1554);
nor U5954 (N_5954,In_1087,In_1378);
xnor U5955 (N_5955,In_2316,In_280);
nand U5956 (N_5956,In_1507,In_1781);
nor U5957 (N_5957,In_1172,In_1031);
nor U5958 (N_5958,In_1756,In_1558);
xor U5959 (N_5959,In_119,In_236);
xnor U5960 (N_5960,In_24,In_805);
or U5961 (N_5961,In_173,In_1459);
xnor U5962 (N_5962,In_109,In_2);
nor U5963 (N_5963,In_898,In_1322);
xnor U5964 (N_5964,In_152,In_1168);
nor U5965 (N_5965,In_31,In_1878);
or U5966 (N_5966,In_1633,In_2043);
nor U5967 (N_5967,In_1094,In_619);
nor U5968 (N_5968,In_1210,In_8);
and U5969 (N_5969,In_2037,In_1711);
nor U5970 (N_5970,In_1486,In_1715);
or U5971 (N_5971,In_310,In_2144);
nand U5972 (N_5972,In_769,In_1760);
or U5973 (N_5973,In_2056,In_1404);
xnor U5974 (N_5974,In_596,In_587);
or U5975 (N_5975,In_690,In_1761);
xnor U5976 (N_5976,In_2373,In_2452);
nand U5977 (N_5977,In_116,In_622);
or U5978 (N_5978,In_2043,In_298);
nor U5979 (N_5979,In_1960,In_707);
nor U5980 (N_5980,In_302,In_1159);
and U5981 (N_5981,In_1763,In_21);
xnor U5982 (N_5982,In_1079,In_1629);
nor U5983 (N_5983,In_657,In_164);
or U5984 (N_5984,In_726,In_566);
xnor U5985 (N_5985,In_1917,In_485);
xnor U5986 (N_5986,In_884,In_440);
xor U5987 (N_5987,In_1880,In_720);
or U5988 (N_5988,In_2115,In_1718);
and U5989 (N_5989,In_416,In_1879);
and U5990 (N_5990,In_2186,In_535);
nand U5991 (N_5991,In_1793,In_1640);
or U5992 (N_5992,In_757,In_400);
and U5993 (N_5993,In_457,In_1152);
xnor U5994 (N_5994,In_399,In_1193);
nand U5995 (N_5995,In_1798,In_1611);
nand U5996 (N_5996,In_1422,In_924);
or U5997 (N_5997,In_1133,In_881);
or U5998 (N_5998,In_2365,In_2161);
or U5999 (N_5999,In_346,In_852);
or U6000 (N_6000,In_692,In_1495);
nand U6001 (N_6001,In_276,In_1077);
and U6002 (N_6002,In_1575,In_694);
nand U6003 (N_6003,In_698,In_496);
nand U6004 (N_6004,In_2426,In_1066);
nor U6005 (N_6005,In_207,In_1214);
nor U6006 (N_6006,In_362,In_1419);
xnor U6007 (N_6007,In_1478,In_488);
or U6008 (N_6008,In_321,In_1302);
and U6009 (N_6009,In_1797,In_1620);
or U6010 (N_6010,In_1366,In_1819);
and U6011 (N_6011,In_2354,In_483);
xor U6012 (N_6012,In_1222,In_1690);
xor U6013 (N_6013,In_1536,In_1663);
xnor U6014 (N_6014,In_711,In_1260);
or U6015 (N_6015,In_117,In_1068);
nand U6016 (N_6016,In_2247,In_2164);
or U6017 (N_6017,In_1933,In_447);
xnor U6018 (N_6018,In_1684,In_317);
nand U6019 (N_6019,In_1669,In_1335);
xor U6020 (N_6020,In_2406,In_360);
or U6021 (N_6021,In_2486,In_1461);
or U6022 (N_6022,In_611,In_2295);
or U6023 (N_6023,In_1796,In_1691);
or U6024 (N_6024,In_2223,In_1266);
nand U6025 (N_6025,In_1192,In_1625);
nand U6026 (N_6026,In_2305,In_728);
nand U6027 (N_6027,In_624,In_2333);
and U6028 (N_6028,In_1568,In_821);
or U6029 (N_6029,In_1516,In_192);
nand U6030 (N_6030,In_80,In_98);
nand U6031 (N_6031,In_171,In_726);
xor U6032 (N_6032,In_2078,In_1302);
nand U6033 (N_6033,In_905,In_2107);
nand U6034 (N_6034,In_1599,In_930);
or U6035 (N_6035,In_1474,In_1406);
nor U6036 (N_6036,In_1745,In_776);
nor U6037 (N_6037,In_198,In_2363);
nor U6038 (N_6038,In_497,In_1902);
nand U6039 (N_6039,In_474,In_589);
or U6040 (N_6040,In_1551,In_1101);
or U6041 (N_6041,In_1075,In_1672);
nor U6042 (N_6042,In_1240,In_1930);
nand U6043 (N_6043,In_1392,In_988);
or U6044 (N_6044,In_687,In_2330);
nand U6045 (N_6045,In_1327,In_979);
nand U6046 (N_6046,In_754,In_1754);
nand U6047 (N_6047,In_2455,In_583);
or U6048 (N_6048,In_282,In_1108);
xnor U6049 (N_6049,In_2016,In_2471);
xnor U6050 (N_6050,In_1231,In_388);
nand U6051 (N_6051,In_246,In_829);
nand U6052 (N_6052,In_438,In_468);
and U6053 (N_6053,In_181,In_2318);
and U6054 (N_6054,In_1425,In_924);
and U6055 (N_6055,In_1610,In_2468);
xor U6056 (N_6056,In_1163,In_656);
and U6057 (N_6057,In_1552,In_395);
nand U6058 (N_6058,In_1242,In_1011);
xor U6059 (N_6059,In_1674,In_1258);
nor U6060 (N_6060,In_54,In_2398);
or U6061 (N_6061,In_412,In_496);
nand U6062 (N_6062,In_2175,In_1972);
xor U6063 (N_6063,In_1251,In_427);
xnor U6064 (N_6064,In_1601,In_1092);
or U6065 (N_6065,In_267,In_161);
nand U6066 (N_6066,In_1255,In_2112);
xor U6067 (N_6067,In_1293,In_1883);
xor U6068 (N_6068,In_1800,In_1051);
nand U6069 (N_6069,In_1374,In_2353);
xnor U6070 (N_6070,In_1514,In_2126);
nor U6071 (N_6071,In_2269,In_1428);
nand U6072 (N_6072,In_54,In_2323);
nand U6073 (N_6073,In_980,In_1229);
nor U6074 (N_6074,In_734,In_2452);
nand U6075 (N_6075,In_850,In_1092);
and U6076 (N_6076,In_2231,In_1110);
nor U6077 (N_6077,In_1629,In_209);
xnor U6078 (N_6078,In_2416,In_827);
nor U6079 (N_6079,In_1409,In_1363);
xnor U6080 (N_6080,In_463,In_2199);
nor U6081 (N_6081,In_649,In_1018);
xnor U6082 (N_6082,In_203,In_1061);
nand U6083 (N_6083,In_536,In_84);
nand U6084 (N_6084,In_600,In_2487);
and U6085 (N_6085,In_1138,In_2262);
or U6086 (N_6086,In_1356,In_458);
or U6087 (N_6087,In_526,In_586);
nand U6088 (N_6088,In_2262,In_205);
xor U6089 (N_6089,In_2489,In_309);
or U6090 (N_6090,In_2166,In_1454);
xor U6091 (N_6091,In_1006,In_96);
nor U6092 (N_6092,In_1700,In_2197);
nand U6093 (N_6093,In_728,In_274);
nand U6094 (N_6094,In_1053,In_222);
nor U6095 (N_6095,In_970,In_1409);
nor U6096 (N_6096,In_305,In_184);
nand U6097 (N_6097,In_1229,In_954);
and U6098 (N_6098,In_1149,In_2058);
xor U6099 (N_6099,In_1778,In_2374);
nand U6100 (N_6100,In_1053,In_694);
or U6101 (N_6101,In_1929,In_914);
xor U6102 (N_6102,In_2118,In_1121);
nor U6103 (N_6103,In_1480,In_690);
xor U6104 (N_6104,In_1978,In_305);
or U6105 (N_6105,In_648,In_1562);
nand U6106 (N_6106,In_1279,In_103);
nor U6107 (N_6107,In_1367,In_120);
and U6108 (N_6108,In_2498,In_974);
xor U6109 (N_6109,In_112,In_1004);
nand U6110 (N_6110,In_2432,In_2042);
nand U6111 (N_6111,In_319,In_1991);
or U6112 (N_6112,In_322,In_292);
and U6113 (N_6113,In_110,In_2336);
nor U6114 (N_6114,In_2431,In_896);
xnor U6115 (N_6115,In_1950,In_278);
xnor U6116 (N_6116,In_650,In_2194);
xnor U6117 (N_6117,In_896,In_1109);
or U6118 (N_6118,In_318,In_1611);
xnor U6119 (N_6119,In_1876,In_1903);
or U6120 (N_6120,In_98,In_1781);
nand U6121 (N_6121,In_2246,In_341);
or U6122 (N_6122,In_1029,In_1789);
or U6123 (N_6123,In_338,In_1006);
nand U6124 (N_6124,In_1754,In_2105);
and U6125 (N_6125,In_913,In_1352);
nor U6126 (N_6126,In_1997,In_1731);
or U6127 (N_6127,In_2223,In_2093);
nand U6128 (N_6128,In_2458,In_2410);
or U6129 (N_6129,In_692,In_495);
nand U6130 (N_6130,In_1922,In_39);
and U6131 (N_6131,In_853,In_1489);
xor U6132 (N_6132,In_1746,In_330);
nand U6133 (N_6133,In_2073,In_985);
nand U6134 (N_6134,In_1055,In_1593);
nand U6135 (N_6135,In_1907,In_460);
nor U6136 (N_6136,In_856,In_2244);
xnor U6137 (N_6137,In_1439,In_1707);
xor U6138 (N_6138,In_2233,In_1008);
or U6139 (N_6139,In_2147,In_2449);
and U6140 (N_6140,In_1056,In_807);
xnor U6141 (N_6141,In_1492,In_2143);
nand U6142 (N_6142,In_2344,In_1321);
or U6143 (N_6143,In_398,In_995);
and U6144 (N_6144,In_2091,In_1347);
nand U6145 (N_6145,In_1164,In_2329);
nand U6146 (N_6146,In_1457,In_2419);
or U6147 (N_6147,In_2449,In_1467);
xor U6148 (N_6148,In_665,In_2090);
and U6149 (N_6149,In_586,In_280);
xor U6150 (N_6150,In_2261,In_2485);
nor U6151 (N_6151,In_1769,In_2345);
nand U6152 (N_6152,In_866,In_111);
or U6153 (N_6153,In_2181,In_1232);
or U6154 (N_6154,In_284,In_636);
nor U6155 (N_6155,In_1497,In_1749);
or U6156 (N_6156,In_775,In_2051);
xor U6157 (N_6157,In_1360,In_1934);
nor U6158 (N_6158,In_1439,In_1146);
or U6159 (N_6159,In_1257,In_144);
and U6160 (N_6160,In_2398,In_1938);
and U6161 (N_6161,In_2211,In_6);
and U6162 (N_6162,In_1308,In_740);
xnor U6163 (N_6163,In_942,In_709);
and U6164 (N_6164,In_623,In_477);
xnor U6165 (N_6165,In_1971,In_2249);
nand U6166 (N_6166,In_2390,In_2208);
nand U6167 (N_6167,In_175,In_2315);
nor U6168 (N_6168,In_370,In_1358);
xor U6169 (N_6169,In_2370,In_2419);
or U6170 (N_6170,In_2218,In_1296);
nand U6171 (N_6171,In_1946,In_1291);
or U6172 (N_6172,In_175,In_351);
nand U6173 (N_6173,In_1099,In_1204);
and U6174 (N_6174,In_1145,In_1620);
and U6175 (N_6175,In_2300,In_2310);
or U6176 (N_6176,In_2248,In_2104);
nor U6177 (N_6177,In_303,In_1430);
xnor U6178 (N_6178,In_89,In_2482);
xnor U6179 (N_6179,In_174,In_1284);
nand U6180 (N_6180,In_106,In_887);
nand U6181 (N_6181,In_288,In_1371);
nor U6182 (N_6182,In_89,In_76);
xnor U6183 (N_6183,In_2267,In_1832);
nand U6184 (N_6184,In_53,In_372);
xnor U6185 (N_6185,In_1325,In_1474);
and U6186 (N_6186,In_552,In_623);
nand U6187 (N_6187,In_1595,In_2446);
and U6188 (N_6188,In_2100,In_1998);
and U6189 (N_6189,In_426,In_1881);
or U6190 (N_6190,In_2267,In_499);
xnor U6191 (N_6191,In_778,In_356);
and U6192 (N_6192,In_126,In_1505);
or U6193 (N_6193,In_848,In_2488);
or U6194 (N_6194,In_474,In_436);
and U6195 (N_6195,In_154,In_2167);
nand U6196 (N_6196,In_790,In_840);
and U6197 (N_6197,In_520,In_1245);
nor U6198 (N_6198,In_2325,In_966);
and U6199 (N_6199,In_465,In_1683);
xor U6200 (N_6200,In_549,In_1899);
xor U6201 (N_6201,In_1234,In_1937);
xor U6202 (N_6202,In_2365,In_1493);
or U6203 (N_6203,In_857,In_849);
and U6204 (N_6204,In_1941,In_34);
and U6205 (N_6205,In_836,In_13);
xnor U6206 (N_6206,In_255,In_1350);
or U6207 (N_6207,In_217,In_349);
and U6208 (N_6208,In_1843,In_152);
nand U6209 (N_6209,In_940,In_1264);
or U6210 (N_6210,In_2478,In_2106);
xor U6211 (N_6211,In_2181,In_742);
nor U6212 (N_6212,In_318,In_1883);
xnor U6213 (N_6213,In_1085,In_2382);
nand U6214 (N_6214,In_1950,In_847);
nor U6215 (N_6215,In_2161,In_174);
or U6216 (N_6216,In_1872,In_726);
or U6217 (N_6217,In_648,In_441);
nor U6218 (N_6218,In_1822,In_1837);
nor U6219 (N_6219,In_487,In_573);
nand U6220 (N_6220,In_2437,In_581);
nor U6221 (N_6221,In_2100,In_830);
nand U6222 (N_6222,In_880,In_1102);
or U6223 (N_6223,In_268,In_1485);
and U6224 (N_6224,In_1727,In_1073);
or U6225 (N_6225,In_1226,In_146);
nor U6226 (N_6226,In_2105,In_1017);
xnor U6227 (N_6227,In_587,In_2001);
nor U6228 (N_6228,In_1498,In_966);
and U6229 (N_6229,In_220,In_1151);
or U6230 (N_6230,In_2087,In_676);
xnor U6231 (N_6231,In_537,In_776);
and U6232 (N_6232,In_1636,In_2455);
or U6233 (N_6233,In_521,In_221);
nor U6234 (N_6234,In_1119,In_2381);
and U6235 (N_6235,In_2046,In_1607);
nor U6236 (N_6236,In_1274,In_129);
nand U6237 (N_6237,In_336,In_563);
and U6238 (N_6238,In_1146,In_763);
nand U6239 (N_6239,In_900,In_1948);
xnor U6240 (N_6240,In_1448,In_1413);
nor U6241 (N_6241,In_526,In_2197);
and U6242 (N_6242,In_2,In_847);
and U6243 (N_6243,In_126,In_906);
and U6244 (N_6244,In_1132,In_1216);
or U6245 (N_6245,In_721,In_2225);
xor U6246 (N_6246,In_724,In_1439);
xnor U6247 (N_6247,In_1571,In_7);
xnor U6248 (N_6248,In_1526,In_736);
and U6249 (N_6249,In_306,In_1753);
nand U6250 (N_6250,N_4685,N_1823);
or U6251 (N_6251,N_5493,N_2364);
and U6252 (N_6252,N_3381,N_5681);
nor U6253 (N_6253,N_4851,N_5355);
nor U6254 (N_6254,N_5755,N_2654);
nand U6255 (N_6255,N_5986,N_6115);
nand U6256 (N_6256,N_1713,N_413);
nor U6257 (N_6257,N_4937,N_362);
nor U6258 (N_6258,N_4087,N_5226);
and U6259 (N_6259,N_2342,N_981);
nor U6260 (N_6260,N_406,N_3225);
or U6261 (N_6261,N_3441,N_1492);
or U6262 (N_6262,N_146,N_1202);
and U6263 (N_6263,N_2737,N_3097);
nor U6264 (N_6264,N_5813,N_493);
nand U6265 (N_6265,N_1047,N_4025);
xor U6266 (N_6266,N_6097,N_2754);
nand U6267 (N_6267,N_6125,N_1976);
and U6268 (N_6268,N_4178,N_1053);
and U6269 (N_6269,N_3801,N_6246);
xor U6270 (N_6270,N_5034,N_5603);
xor U6271 (N_6271,N_4397,N_5770);
nor U6272 (N_6272,N_5531,N_3330);
nand U6273 (N_6273,N_4664,N_6021);
or U6274 (N_6274,N_5463,N_573);
nand U6275 (N_6275,N_5663,N_3004);
xor U6276 (N_6276,N_4272,N_2302);
nor U6277 (N_6277,N_4845,N_1716);
and U6278 (N_6278,N_5162,N_2917);
nor U6279 (N_6279,N_6018,N_81);
xnor U6280 (N_6280,N_3933,N_5227);
and U6281 (N_6281,N_1003,N_3333);
nor U6282 (N_6282,N_1511,N_2515);
nand U6283 (N_6283,N_1841,N_2106);
nor U6284 (N_6284,N_4719,N_3064);
nor U6285 (N_6285,N_3204,N_6088);
or U6286 (N_6286,N_746,N_3835);
nor U6287 (N_6287,N_5348,N_291);
or U6288 (N_6288,N_2058,N_2794);
nor U6289 (N_6289,N_3453,N_2994);
nor U6290 (N_6290,N_2714,N_5680);
and U6291 (N_6291,N_3949,N_2743);
xor U6292 (N_6292,N_6071,N_5840);
or U6293 (N_6293,N_145,N_4654);
nor U6294 (N_6294,N_214,N_1617);
xnor U6295 (N_6295,N_4760,N_4809);
nor U6296 (N_6296,N_3559,N_2059);
or U6297 (N_6297,N_722,N_1778);
xnor U6298 (N_6298,N_4779,N_4256);
nand U6299 (N_6299,N_2474,N_1870);
nor U6300 (N_6300,N_5653,N_800);
nand U6301 (N_6301,N_4278,N_969);
or U6302 (N_6302,N_1142,N_477);
xor U6303 (N_6303,N_1443,N_433);
and U6304 (N_6304,N_5931,N_4544);
or U6305 (N_6305,N_3399,N_1735);
and U6306 (N_6306,N_3943,N_4449);
and U6307 (N_6307,N_3880,N_4606);
nor U6308 (N_6308,N_875,N_2121);
nand U6309 (N_6309,N_5209,N_1149);
or U6310 (N_6310,N_683,N_961);
and U6311 (N_6311,N_4669,N_5554);
nor U6312 (N_6312,N_872,N_5989);
nand U6313 (N_6313,N_3718,N_5578);
nor U6314 (N_6314,N_3270,N_3211);
or U6315 (N_6315,N_5788,N_5023);
nand U6316 (N_6316,N_2362,N_5766);
and U6317 (N_6317,N_218,N_3557);
or U6318 (N_6318,N_1738,N_2128);
xnor U6319 (N_6319,N_6038,N_2397);
nor U6320 (N_6320,N_1324,N_4808);
nor U6321 (N_6321,N_3051,N_3793);
and U6322 (N_6322,N_3572,N_3058);
nand U6323 (N_6323,N_1311,N_2719);
or U6324 (N_6324,N_2579,N_6064);
and U6325 (N_6325,N_5735,N_3057);
or U6326 (N_6326,N_93,N_1117);
nor U6327 (N_6327,N_417,N_4240);
or U6328 (N_6328,N_5979,N_4900);
xor U6329 (N_6329,N_495,N_6230);
nand U6330 (N_6330,N_5937,N_3605);
xnor U6331 (N_6331,N_1669,N_494);
nor U6332 (N_6332,N_4612,N_2844);
nand U6333 (N_6333,N_3872,N_730);
nand U6334 (N_6334,N_45,N_4550);
nand U6335 (N_6335,N_1152,N_2210);
xnor U6336 (N_6336,N_4890,N_2735);
nor U6337 (N_6337,N_5389,N_5095);
or U6338 (N_6338,N_2919,N_3767);
nand U6339 (N_6339,N_445,N_2442);
or U6340 (N_6340,N_2260,N_6106);
nor U6341 (N_6341,N_4530,N_904);
and U6342 (N_6342,N_1074,N_2586);
and U6343 (N_6343,N_6191,N_2452);
xor U6344 (N_6344,N_3878,N_1515);
xor U6345 (N_6345,N_2407,N_2079);
and U6346 (N_6346,N_6089,N_6155);
or U6347 (N_6347,N_850,N_4261);
nor U6348 (N_6348,N_1840,N_1925);
nand U6349 (N_6349,N_5777,N_2825);
nand U6350 (N_6350,N_4827,N_3323);
and U6351 (N_6351,N_5909,N_5829);
and U6352 (N_6352,N_325,N_91);
or U6353 (N_6353,N_1508,N_3296);
nor U6354 (N_6354,N_1328,N_398);
xor U6355 (N_6355,N_1245,N_2701);
nand U6356 (N_6356,N_88,N_6);
nand U6357 (N_6357,N_4994,N_3839);
nor U6358 (N_6358,N_3674,N_2665);
or U6359 (N_6359,N_2390,N_348);
and U6360 (N_6360,N_6236,N_1795);
and U6361 (N_6361,N_1058,N_1538);
nor U6362 (N_6362,N_536,N_4614);
and U6363 (N_6363,N_2114,N_1908);
and U6364 (N_6364,N_375,N_963);
or U6365 (N_6365,N_2771,N_828);
and U6366 (N_6366,N_2975,N_6219);
nand U6367 (N_6367,N_4535,N_5070);
or U6368 (N_6368,N_2140,N_2959);
nand U6369 (N_6369,N_617,N_3998);
and U6370 (N_6370,N_6004,N_2011);
nor U6371 (N_6371,N_2125,N_1471);
nand U6372 (N_6372,N_684,N_3581);
or U6373 (N_6373,N_2633,N_2045);
or U6374 (N_6374,N_3575,N_3929);
nand U6375 (N_6375,N_6133,N_1869);
xor U6376 (N_6376,N_5089,N_133);
xor U6377 (N_6377,N_932,N_6249);
nor U6378 (N_6378,N_5573,N_3950);
xnor U6379 (N_6379,N_3926,N_1213);
xor U6380 (N_6380,N_3957,N_4354);
nand U6381 (N_6381,N_4643,N_2532);
nor U6382 (N_6382,N_868,N_4842);
xnor U6383 (N_6383,N_4466,N_2672);
and U6384 (N_6384,N_4062,N_1051);
or U6385 (N_6385,N_3707,N_3053);
or U6386 (N_6386,N_3639,N_4181);
nand U6387 (N_6387,N_1276,N_5193);
nand U6388 (N_6388,N_639,N_2393);
xnor U6389 (N_6389,N_4621,N_2257);
and U6390 (N_6390,N_2187,N_1323);
nand U6391 (N_6391,N_2884,N_4149);
or U6392 (N_6392,N_566,N_5361);
nor U6393 (N_6393,N_387,N_1235);
nor U6394 (N_6394,N_2043,N_1846);
xor U6395 (N_6395,N_4444,N_4468);
or U6396 (N_6396,N_5006,N_1940);
xor U6397 (N_6397,N_2836,N_4784);
xor U6398 (N_6398,N_1601,N_570);
nand U6399 (N_6399,N_2376,N_4789);
nand U6400 (N_6400,N_2280,N_4419);
xnor U6401 (N_6401,N_5948,N_6218);
or U6402 (N_6402,N_905,N_708);
and U6403 (N_6403,N_2296,N_163);
or U6404 (N_6404,N_4145,N_4484);
or U6405 (N_6405,N_5163,N_3494);
and U6406 (N_6406,N_5700,N_1594);
and U6407 (N_6407,N_3744,N_4655);
nor U6408 (N_6408,N_1250,N_5907);
xnor U6409 (N_6409,N_4184,N_4716);
xnor U6410 (N_6410,N_3106,N_1688);
nor U6411 (N_6411,N_3711,N_3772);
or U6412 (N_6412,N_4213,N_3466);
or U6413 (N_6413,N_4035,N_3840);
nand U6414 (N_6414,N_578,N_2469);
nand U6415 (N_6415,N_4895,N_5819);
nor U6416 (N_6416,N_2887,N_2698);
and U6417 (N_6417,N_5599,N_1584);
xor U6418 (N_6418,N_6077,N_4101);
nand U6419 (N_6419,N_1698,N_436);
nor U6420 (N_6420,N_5543,N_5094);
and U6421 (N_6421,N_2731,N_4347);
xor U6422 (N_6422,N_5188,N_6035);
or U6423 (N_6423,N_3791,N_3411);
or U6424 (N_6424,N_1804,N_1364);
and U6425 (N_6425,N_5113,N_3721);
nor U6426 (N_6426,N_2823,N_948);
nor U6427 (N_6427,N_174,N_5678);
and U6428 (N_6428,N_4099,N_129);
nor U6429 (N_6429,N_4751,N_3329);
xor U6430 (N_6430,N_3511,N_4266);
or U6431 (N_6431,N_4799,N_4316);
nand U6432 (N_6432,N_5849,N_3003);
and U6433 (N_6433,N_1434,N_6027);
and U6434 (N_6434,N_3770,N_4399);
nand U6435 (N_6435,N_333,N_2635);
nand U6436 (N_6436,N_2668,N_2160);
nand U6437 (N_6437,N_3101,N_350);
and U6438 (N_6438,N_3126,N_2749);
nand U6439 (N_6439,N_4408,N_8);
xor U6440 (N_6440,N_4246,N_3351);
xor U6441 (N_6441,N_3592,N_2688);
nand U6442 (N_6442,N_5311,N_1215);
and U6443 (N_6443,N_4858,N_4407);
xor U6444 (N_6444,N_5154,N_86);
xor U6445 (N_6445,N_3577,N_2873);
or U6446 (N_6446,N_3188,N_2645);
xnor U6447 (N_6447,N_1307,N_3060);
nor U6448 (N_6448,N_2261,N_2923);
xor U6449 (N_6449,N_4877,N_2632);
nand U6450 (N_6450,N_720,N_3017);
and U6451 (N_6451,N_267,N_6130);
nand U6452 (N_6452,N_3022,N_3606);
nand U6453 (N_6453,N_2153,N_3964);
nand U6454 (N_6454,N_478,N_3334);
xnor U6455 (N_6455,N_1251,N_2175);
xor U6456 (N_6456,N_733,N_5468);
and U6457 (N_6457,N_5148,N_6135);
or U6458 (N_6458,N_1334,N_5642);
nor U6459 (N_6459,N_35,N_2109);
nor U6460 (N_6460,N_5858,N_5533);
xnor U6461 (N_6461,N_4392,N_5269);
nor U6462 (N_6462,N_3205,N_1168);
or U6463 (N_6463,N_701,N_4624);
nor U6464 (N_6464,N_1977,N_5494);
nor U6465 (N_6465,N_560,N_839);
nor U6466 (N_6466,N_4817,N_3692);
nand U6467 (N_6467,N_3966,N_4514);
and U6468 (N_6468,N_1270,N_3139);
xor U6469 (N_6469,N_6151,N_51);
nand U6470 (N_6470,N_313,N_2792);
nand U6471 (N_6471,N_4462,N_1791);
nand U6472 (N_6472,N_4322,N_5080);
and U6473 (N_6473,N_4837,N_5575);
nand U6474 (N_6474,N_463,N_1773);
xnor U6475 (N_6475,N_3815,N_724);
or U6476 (N_6476,N_4772,N_5496);
nand U6477 (N_6477,N_5536,N_4192);
nor U6478 (N_6478,N_4375,N_5305);
nand U6479 (N_6479,N_4095,N_6205);
and U6480 (N_6480,N_3916,N_6190);
nor U6481 (N_6481,N_3128,N_1026);
and U6482 (N_6482,N_4790,N_3183);
xnor U6483 (N_6483,N_1563,N_212);
xnor U6484 (N_6484,N_728,N_3102);
nor U6485 (N_6485,N_2584,N_6170);
nand U6486 (N_6486,N_3138,N_5697);
and U6487 (N_6487,N_4430,N_1847);
xor U6488 (N_6488,N_6059,N_4414);
and U6489 (N_6489,N_6046,N_512);
nor U6490 (N_6490,N_202,N_4455);
nand U6491 (N_6491,N_625,N_2608);
or U6492 (N_6492,N_3987,N_44);
or U6493 (N_6493,N_4584,N_518);
or U6494 (N_6494,N_6194,N_565);
nand U6495 (N_6495,N_5122,N_42);
and U6496 (N_6496,N_1579,N_274);
nor U6497 (N_6497,N_5143,N_2101);
or U6498 (N_6498,N_4488,N_2269);
nand U6499 (N_6499,N_4166,N_2639);
and U6500 (N_6500,N_1017,N_3990);
nand U6501 (N_6501,N_4954,N_6026);
or U6502 (N_6502,N_4541,N_5545);
and U6503 (N_6503,N_3873,N_378);
xnor U6504 (N_6504,N_702,N_2640);
or U6505 (N_6505,N_806,N_1640);
nor U6506 (N_6506,N_879,N_5888);
xnor U6507 (N_6507,N_5033,N_510);
xnor U6508 (N_6508,N_5927,N_38);
nor U6509 (N_6509,N_216,N_2458);
nand U6510 (N_6510,N_3985,N_4296);
xnor U6511 (N_6511,N_1595,N_1268);
nor U6512 (N_6512,N_2089,N_551);
and U6513 (N_6513,N_3626,N_4824);
nor U6514 (N_6514,N_5624,N_4565);
and U6515 (N_6515,N_1062,N_1897);
and U6516 (N_6516,N_1257,N_393);
nor U6517 (N_6517,N_5067,N_2065);
xor U6518 (N_6518,N_5489,N_1691);
and U6519 (N_6519,N_5881,N_4745);
nand U6520 (N_6520,N_4313,N_2829);
xnor U6521 (N_6521,N_863,N_4485);
nand U6522 (N_6522,N_3689,N_3306);
or U6523 (N_6523,N_6043,N_3221);
xnor U6524 (N_6524,N_237,N_658);
or U6525 (N_6525,N_3005,N_4801);
nand U6526 (N_6526,N_2624,N_4008);
nor U6527 (N_6527,N_1483,N_401);
xor U6528 (N_6528,N_1126,N_3912);
nand U6529 (N_6529,N_5445,N_1302);
nand U6530 (N_6530,N_2961,N_46);
nand U6531 (N_6531,N_5619,N_5180);
or U6532 (N_6532,N_1566,N_2807);
or U6533 (N_6533,N_3960,N_3182);
nand U6534 (N_6534,N_5201,N_469);
nor U6535 (N_6535,N_2508,N_1242);
nand U6536 (N_6536,N_1796,N_1551);
or U6537 (N_6537,N_2497,N_1442);
nand U6538 (N_6538,N_1934,N_287);
nor U6539 (N_6539,N_833,N_2834);
xor U6540 (N_6540,N_3226,N_5977);
nand U6541 (N_6541,N_226,N_6212);
or U6542 (N_6542,N_1346,N_688);
nand U6543 (N_6543,N_1024,N_3380);
and U6544 (N_6544,N_3391,N_444);
nand U6545 (N_6545,N_990,N_2385);
or U6546 (N_6546,N_3341,N_190);
nor U6547 (N_6547,N_4668,N_592);
and U6548 (N_6548,N_1936,N_4021);
nor U6549 (N_6549,N_4766,N_1468);
or U6550 (N_6550,N_4497,N_6148);
nand U6551 (N_6551,N_2185,N_1931);
nand U6552 (N_6552,N_2682,N_2530);
xor U6553 (N_6553,N_3970,N_2411);
xor U6554 (N_6554,N_5257,N_2055);
or U6555 (N_6555,N_2309,N_3473);
or U6556 (N_6556,N_4627,N_4412);
and U6557 (N_6557,N_4415,N_2386);
or U6558 (N_6558,N_2226,N_5669);
xnor U6559 (N_6559,N_3385,N_4041);
and U6560 (N_6560,N_2343,N_4786);
nor U6561 (N_6561,N_3922,N_3851);
and U6562 (N_6562,N_3162,N_2400);
or U6563 (N_6563,N_3170,N_4956);
xor U6564 (N_6564,N_3039,N_2194);
nand U6565 (N_6565,N_4733,N_5921);
xor U6566 (N_6566,N_6163,N_3779);
nand U6567 (N_6567,N_3075,N_4540);
nand U6568 (N_6568,N_703,N_845);
and U6569 (N_6569,N_2980,N_5260);
and U6570 (N_6570,N_2694,N_968);
or U6571 (N_6571,N_5827,N_5808);
nor U6572 (N_6572,N_3663,N_4708);
xnor U6573 (N_6573,N_5996,N_6181);
xor U6574 (N_6574,N_1389,N_6006);
xnor U6575 (N_6575,N_751,N_5346);
nand U6576 (N_6576,N_647,N_3078);
xor U6577 (N_6577,N_5694,N_4335);
and U6578 (N_6578,N_3971,N_4486);
xor U6579 (N_6579,N_514,N_747);
nor U6580 (N_6580,N_3734,N_768);
or U6581 (N_6581,N_1297,N_5385);
and U6582 (N_6582,N_232,N_5394);
nand U6583 (N_6583,N_4102,N_3690);
xnor U6584 (N_6584,N_2818,N_3681);
nor U6585 (N_6585,N_2489,N_2828);
and U6586 (N_6586,N_5276,N_2705);
xnor U6587 (N_6587,N_1793,N_3703);
and U6588 (N_6588,N_1040,N_2435);
and U6589 (N_6589,N_5284,N_1306);
and U6590 (N_6590,N_4359,N_2144);
nand U6591 (N_6591,N_4290,N_4253);
or U6592 (N_6592,N_3216,N_5894);
nand U6593 (N_6593,N_2889,N_540);
xor U6594 (N_6594,N_3091,N_5606);
nor U6595 (N_6595,N_4024,N_3918);
nand U6596 (N_6596,N_4918,N_1955);
xnor U6597 (N_6597,N_5842,N_3315);
nor U6598 (N_6598,N_3065,N_1777);
or U6599 (N_6599,N_3623,N_5147);
xor U6600 (N_6600,N_1507,N_4252);
and U6601 (N_6601,N_1304,N_458);
nor U6602 (N_6602,N_2237,N_4969);
and U6603 (N_6603,N_4961,N_3273);
and U6604 (N_6604,N_454,N_5843);
and U6605 (N_6605,N_5851,N_4351);
xor U6606 (N_6606,N_5453,N_3742);
and U6607 (N_6607,N_4276,N_157);
or U6608 (N_6608,N_4919,N_3253);
nor U6609 (N_6609,N_685,N_5923);
and U6610 (N_6610,N_5865,N_1537);
nand U6611 (N_6611,N_5446,N_4736);
or U6612 (N_6612,N_3968,N_158);
nand U6613 (N_6613,N_5214,N_546);
or U6614 (N_6614,N_4601,N_2084);
nor U6615 (N_6615,N_2326,N_669);
xnor U6616 (N_6616,N_6174,N_3601);
nand U6617 (N_6617,N_1922,N_1899);
xor U6618 (N_6618,N_439,N_3917);
nor U6619 (N_6619,N_2293,N_2760);
nand U6620 (N_6620,N_3762,N_3165);
nor U6621 (N_6621,N_3999,N_2088);
nand U6622 (N_6622,N_310,N_3530);
xnor U6623 (N_6623,N_1676,N_2547);
nand U6624 (N_6624,N_3092,N_3665);
nand U6625 (N_6625,N_2858,N_5086);
xnor U6626 (N_6626,N_4150,N_553);
nand U6627 (N_6627,N_502,N_6114);
nor U6628 (N_6628,N_3321,N_4834);
nand U6629 (N_6629,N_1065,N_2942);
nand U6630 (N_6630,N_4060,N_3508);
nand U6631 (N_6631,N_4479,N_4501);
nand U6632 (N_6632,N_6060,N_3836);
nor U6633 (N_6633,N_552,N_98);
xnor U6634 (N_6634,N_5875,N_5487);
nand U6635 (N_6635,N_1907,N_2747);
or U6636 (N_6636,N_1265,N_3140);
and U6637 (N_6637,N_1813,N_180);
and U6638 (N_6638,N_5130,N_5885);
or U6639 (N_6639,N_2085,N_1190);
nor U6640 (N_6640,N_3594,N_3865);
xor U6641 (N_6641,N_3485,N_5010);
nand U6642 (N_6642,N_6072,N_194);
nor U6643 (N_6643,N_5457,N_2073);
and U6644 (N_6644,N_5149,N_5863);
nand U6645 (N_6645,N_3090,N_3370);
nand U6646 (N_6646,N_723,N_4314);
or U6647 (N_6647,N_418,N_3729);
and U6648 (N_6648,N_3234,N_1606);
xnor U6649 (N_6649,N_1219,N_1423);
nand U6650 (N_6650,N_2596,N_140);
xnor U6651 (N_6651,N_4570,N_5435);
or U6652 (N_6652,N_3849,N_6104);
nor U6653 (N_6653,N_4810,N_5527);
xor U6654 (N_6654,N_6134,N_1231);
xnor U6655 (N_6655,N_5768,N_4717);
or U6656 (N_6656,N_3363,N_4475);
nand U6657 (N_6657,N_49,N_317);
nor U6658 (N_6658,N_646,N_320);
nor U6659 (N_6659,N_3108,N_1920);
nand U6660 (N_6660,N_2851,N_1638);
or U6661 (N_6661,N_2231,N_118);
nor U6662 (N_6662,N_4720,N_2782);
nand U6663 (N_6663,N_3266,N_1352);
or U6664 (N_6664,N_4338,N_1968);
or U6665 (N_6665,N_917,N_2205);
and U6666 (N_6666,N_3967,N_80);
xor U6667 (N_6667,N_4306,N_3656);
nor U6668 (N_6668,N_5383,N_54);
nand U6669 (N_6669,N_1919,N_742);
and U6670 (N_6670,N_4863,N_753);
and U6671 (N_6671,N_4925,N_1137);
nand U6672 (N_6672,N_588,N_3);
xnor U6673 (N_6673,N_865,N_1914);
nor U6674 (N_6674,N_985,N_5776);
or U6675 (N_6675,N_27,N_4406);
xnor U6676 (N_6676,N_4000,N_2690);
and U6677 (N_6677,N_18,N_687);
nor U6678 (N_6678,N_824,N_5739);
nor U6679 (N_6679,N_1808,N_5144);
xnor U6680 (N_6680,N_5549,N_3227);
xnor U6681 (N_6681,N_1371,N_979);
and U6682 (N_6682,N_3921,N_4762);
or U6683 (N_6683,N_5483,N_6164);
or U6684 (N_6684,N_3730,N_6075);
and U6685 (N_6685,N_1170,N_4050);
or U6686 (N_6686,N_3580,N_2607);
xor U6687 (N_6687,N_1435,N_1391);
nand U6688 (N_6688,N_5124,N_1178);
and U6689 (N_6689,N_1417,N_823);
and U6690 (N_6690,N_5454,N_1432);
and U6691 (N_6691,N_6162,N_4388);
and U6692 (N_6692,N_258,N_4704);
nand U6693 (N_6693,N_5207,N_3959);
xor U6694 (N_6694,N_6031,N_5357);
xor U6695 (N_6695,N_3129,N_2693);
nand U6696 (N_6696,N_5568,N_4830);
nor U6697 (N_6697,N_4951,N_3994);
xnor U6698 (N_6698,N_3379,N_3350);
or U6699 (N_6699,N_2796,N_2835);
and U6700 (N_6700,N_3159,N_5956);
or U6701 (N_6701,N_1412,N_860);
nand U6702 (N_6702,N_4500,N_1995);
xor U6703 (N_6703,N_2591,N_2475);
nor U6704 (N_6704,N_1605,N_2173);
and U6705 (N_6705,N_4134,N_446);
or U6706 (N_6706,N_1779,N_246);
nand U6707 (N_6707,N_4334,N_2812);
and U6708 (N_6708,N_2049,N_4543);
nor U6709 (N_6709,N_931,N_988);
nor U6710 (N_6710,N_206,N_4121);
nand U6711 (N_6711,N_3651,N_4431);
nand U6712 (N_6712,N_2500,N_481);
xnor U6713 (N_6713,N_4363,N_2778);
and U6714 (N_6714,N_2966,N_5289);
nand U6715 (N_6715,N_3624,N_4761);
and U6716 (N_6716,N_5484,N_6098);
and U6717 (N_6717,N_5957,N_1743);
and U6718 (N_6718,N_1335,N_2786);
or U6719 (N_6719,N_4265,N_2263);
nand U6720 (N_6720,N_1536,N_4694);
nand U6721 (N_6721,N_852,N_4288);
nand U6722 (N_6722,N_5516,N_4771);
nand U6723 (N_6723,N_910,N_5192);
nand U6724 (N_6724,N_3517,N_6017);
xnor U6725 (N_6725,N_4896,N_2396);
nand U6726 (N_6726,N_816,N_5174);
and U6727 (N_6727,N_3802,N_2227);
xnor U6728 (N_6728,N_5358,N_5797);
and U6729 (N_6729,N_2042,N_727);
nor U6730 (N_6730,N_3208,N_3757);
and U6731 (N_6731,N_5281,N_2466);
nor U6732 (N_6732,N_1624,N_5199);
and U6733 (N_6733,N_2888,N_4516);
or U6734 (N_6734,N_5093,N_1263);
nand U6735 (N_6735,N_5791,N_4273);
or U6736 (N_6736,N_5076,N_2667);
and U6737 (N_6737,N_2282,N_4742);
xnor U6738 (N_6738,N_4110,N_5313);
nand U6739 (N_6739,N_353,N_1657);
nor U6740 (N_6740,N_5521,N_2854);
or U6741 (N_6741,N_256,N_1971);
and U6742 (N_6742,N_3903,N_1121);
nand U6743 (N_6743,N_5138,N_4057);
xor U6744 (N_6744,N_1809,N_641);
nand U6745 (N_6745,N_228,N_1923);
and U6746 (N_6746,N_2992,N_5469);
nand U6747 (N_6747,N_2075,N_1556);
nand U6748 (N_6748,N_2820,N_4985);
nand U6749 (N_6749,N_1771,N_2300);
nor U6750 (N_6750,N_1542,N_4237);
and U6751 (N_6751,N_4702,N_3586);
nor U6752 (N_6752,N_3297,N_3176);
and U6753 (N_6753,N_5727,N_4165);
nor U6754 (N_6754,N_1646,N_3324);
nand U6755 (N_6755,N_3955,N_5475);
or U6756 (N_6756,N_3790,N_1812);
and U6757 (N_6757,N_4836,N_268);
nor U6758 (N_6758,N_2787,N_3547);
or U6759 (N_6759,N_3355,N_3748);
or U6760 (N_6760,N_6223,N_3212);
xor U6761 (N_6761,N_986,N_4828);
or U6762 (N_6762,N_4864,N_4053);
and U6763 (N_6763,N_3392,N_1761);
nor U6764 (N_6764,N_3817,N_2151);
or U6765 (N_6765,N_4190,N_3897);
and U6766 (N_6766,N_5003,N_3218);
and U6767 (N_6767,N_3736,N_3595);
and U6768 (N_6768,N_4673,N_798);
nor U6769 (N_6769,N_3054,N_5765);
or U6770 (N_6770,N_1012,N_4170);
nor U6771 (N_6771,N_2870,N_5430);
nand U6772 (N_6772,N_389,N_3625);
and U6773 (N_6773,N_453,N_4083);
nor U6774 (N_6774,N_2881,N_2236);
nand U6775 (N_6775,N_1588,N_4039);
xor U6776 (N_6776,N_4079,N_515);
and U6777 (N_6777,N_572,N_2158);
nand U6778 (N_6778,N_197,N_5171);
nor U6779 (N_6779,N_1757,N_241);
or U6780 (N_6780,N_5682,N_848);
and U6781 (N_6781,N_5798,N_1034);
or U6782 (N_6782,N_3864,N_2927);
xnor U6783 (N_6783,N_221,N_5510);
xor U6784 (N_6784,N_3134,N_4802);
or U6785 (N_6785,N_1203,N_2802);
or U6786 (N_6786,N_490,N_5823);
xor U6787 (N_6787,N_2074,N_1221);
or U6788 (N_6788,N_152,N_5161);
nand U6789 (N_6789,N_4054,N_5359);
nand U6790 (N_6790,N_5395,N_4474);
nor U6791 (N_6791,N_2278,N_3755);
or U6792 (N_6792,N_3010,N_2230);
and U6793 (N_6793,N_596,N_5751);
and U6794 (N_6794,N_5784,N_1820);
nand U6795 (N_6795,N_4357,N_126);
nand U6796 (N_6796,N_4141,N_1156);
xor U6797 (N_6797,N_2611,N_5304);
nor U6798 (N_6798,N_5477,N_2081);
nor U6799 (N_6799,N_956,N_5179);
and U6800 (N_6800,N_324,N_1684);
nor U6801 (N_6801,N_5438,N_5139);
xor U6802 (N_6802,N_4775,N_3496);
nand U6803 (N_6803,N_5614,N_2208);
xor U6804 (N_6804,N_497,N_900);
nand U6805 (N_6805,N_576,N_5638);
nand U6806 (N_6806,N_2543,N_4732);
nor U6807 (N_6807,N_3224,N_4746);
nand U6808 (N_6808,N_748,N_4542);
nand U6809 (N_6809,N_3209,N_1751);
nor U6810 (N_6810,N_5861,N_5690);
or U6811 (N_6811,N_5995,N_1455);
xnor U6812 (N_6812,N_2190,N_3495);
nor U6813 (N_6813,N_5352,N_1187);
xor U6814 (N_6814,N_4861,N_815);
and U6815 (N_6815,N_6067,N_3307);
xnor U6816 (N_6816,N_2509,N_3766);
or U6817 (N_6817,N_2327,N_6201);
xnor U6818 (N_6818,N_2447,N_6048);
or U6819 (N_6819,N_5115,N_6193);
xnor U6820 (N_6820,N_1446,N_2978);
xor U6821 (N_6821,N_2921,N_1873);
or U6822 (N_6822,N_3468,N_5373);
and U6823 (N_6823,N_365,N_3410);
or U6824 (N_6824,N_1007,N_3353);
nand U6825 (N_6825,N_4257,N_4280);
nor U6826 (N_6826,N_6167,N_5712);
or U6827 (N_6827,N_4119,N_4015);
and U6828 (N_6828,N_4546,N_456);
nand U6829 (N_6829,N_3710,N_2815);
nor U6830 (N_6830,N_3672,N_5743);
and U6831 (N_6831,N_2365,N_6231);
and U6832 (N_6832,N_600,N_2948);
or U6833 (N_6833,N_4293,N_2289);
and U6834 (N_6834,N_3756,N_1411);
xnor U6835 (N_6835,N_773,N_1072);
nand U6836 (N_6836,N_5341,N_196);
nand U6837 (N_6837,N_4040,N_4097);
or U6838 (N_6838,N_1127,N_4232);
xnor U6839 (N_6839,N_332,N_4966);
nand U6840 (N_6840,N_674,N_3318);
and U6841 (N_6841,N_262,N_110);
or U6842 (N_6842,N_4349,N_3232);
and U6843 (N_6843,N_2294,N_1672);
and U6844 (N_6844,N_1036,N_5431);
nor U6845 (N_6845,N_4855,N_2761);
or U6846 (N_6846,N_4684,N_999);
or U6847 (N_6847,N_2361,N_71);
and U6848 (N_6848,N_1081,N_1294);
xnor U6849 (N_6849,N_1524,N_4976);
or U6850 (N_6850,N_2029,N_2572);
nand U6851 (N_6851,N_826,N_2661);
xor U6852 (N_6852,N_2072,N_4867);
or U6853 (N_6853,N_5228,N_1658);
or U6854 (N_6854,N_3367,N_5525);
or U6855 (N_6855,N_84,N_5325);
xor U6856 (N_6856,N_1063,N_2568);
nor U6857 (N_6857,N_5805,N_1656);
nor U6858 (N_6858,N_1293,N_635);
nor U6859 (N_6859,N_5736,N_539);
nor U6860 (N_6860,N_4934,N_1504);
or U6861 (N_6861,N_425,N_5471);
nor U6862 (N_6862,N_1548,N_179);
and U6863 (N_6863,N_3015,N_1359);
xnor U6864 (N_6864,N_891,N_3923);
nand U6865 (N_6865,N_41,N_6022);
or U6866 (N_6866,N_1898,N_2307);
or U6867 (N_6867,N_304,N_1912);
nand U6868 (N_6868,N_4756,N_5215);
or U6869 (N_6869,N_2170,N_2984);
and U6870 (N_6870,N_3469,N_3257);
nand U6871 (N_6871,N_3346,N_5030);
nor U6872 (N_6872,N_6100,N_4904);
or U6873 (N_6873,N_2060,N_3844);
xnor U6874 (N_6874,N_4857,N_4251);
and U6875 (N_6875,N_2996,N_5345);
and U6876 (N_6876,N_780,N_2482);
and U6877 (N_6877,N_4064,N_3582);
nand U6878 (N_6878,N_2649,N_3049);
xor U6879 (N_6879,N_1816,N_4868);
or U6880 (N_6880,N_2244,N_5608);
or U6881 (N_6881,N_5836,N_1223);
xnor U6882 (N_6882,N_4782,N_3488);
nand U6883 (N_6883,N_4318,N_6138);
nor U6884 (N_6884,N_4077,N_3609);
or U6885 (N_6885,N_4312,N_370);
or U6886 (N_6886,N_2115,N_5443);
nor U6887 (N_6887,N_5561,N_4561);
nand U6888 (N_6888,N_5272,N_5191);
xor U6889 (N_6889,N_599,N_5418);
nor U6890 (N_6890,N_3322,N_3475);
nor U6891 (N_6891,N_6168,N_4777);
xnor U6892 (N_6892,N_4350,N_4693);
nand U6893 (N_6893,N_3404,N_2181);
or U6894 (N_6894,N_4111,N_40);
or U6895 (N_6895,N_346,N_4944);
or U6896 (N_6896,N_5892,N_2039);
and U6897 (N_6897,N_1406,N_1150);
nand U6898 (N_6898,N_4814,N_210);
nor U6899 (N_6899,N_4058,N_2800);
and U6900 (N_6900,N_4608,N_4045);
nor U6901 (N_6901,N_4681,N_423);
and U6902 (N_6902,N_4203,N_6210);
xnor U6903 (N_6903,N_5296,N_5022);
and U6904 (N_6904,N_4030,N_1558);
nand U6905 (N_6905,N_2773,N_5617);
nor U6906 (N_6906,N_4453,N_6126);
xnor U6907 (N_6907,N_175,N_6082);
or U6908 (N_6908,N_2052,N_4886);
or U6909 (N_6909,N_2589,N_4622);
or U6910 (N_6910,N_4176,N_2646);
nor U6911 (N_6911,N_159,N_1806);
nand U6912 (N_6912,N_3939,N_5787);
nor U6913 (N_6913,N_3310,N_2528);
or U6914 (N_6914,N_2687,N_2511);
nor U6915 (N_6915,N_4426,N_1539);
nand U6916 (N_6916,N_5990,N_2233);
nand U6917 (N_6917,N_1564,N_2879);
and U6918 (N_6918,N_1158,N_134);
nand U6919 (N_6919,N_2179,N_4876);
nand U6920 (N_6920,N_3210,N_5542);
xor U6921 (N_6921,N_5860,N_2673);
and U6922 (N_6922,N_3478,N_2795);
and U6923 (N_6923,N_2006,N_3285);
xnor U6924 (N_6924,N_1102,N_880);
xnor U6925 (N_6925,N_3349,N_1830);
nor U6926 (N_6926,N_5558,N_1801);
xnor U6927 (N_6927,N_1844,N_4109);
nor U6928 (N_6928,N_3133,N_3506);
nor U6929 (N_6929,N_987,N_5998);
nor U6930 (N_6930,N_789,N_473);
or U6931 (N_6931,N_1146,N_5592);
nand U6932 (N_6932,N_5922,N_4436);
nor U6933 (N_6933,N_4358,N_5962);
nand U6934 (N_6934,N_3910,N_4859);
or U6935 (N_6935,N_4072,N_5105);
nor U6936 (N_6936,N_3570,N_3490);
nor U6937 (N_6937,N_3121,N_2862);
and U6938 (N_6938,N_3439,N_1106);
and U6939 (N_6939,N_6206,N_1500);
nor U6940 (N_6940,N_3298,N_6076);
or U6941 (N_6941,N_754,N_737);
xor U6942 (N_6942,N_2392,N_3785);
nand U6943 (N_6943,N_279,N_989);
xnor U6944 (N_6944,N_250,N_5025);
xor U6945 (N_6945,N_5248,N_2195);
nand U6946 (N_6946,N_3445,N_4225);
nor U6947 (N_6947,N_4471,N_2883);
nor U6948 (N_6948,N_5718,N_5703);
nand U6949 (N_6949,N_2838,N_2720);
or U6950 (N_6950,N_3825,N_5462);
nor U6951 (N_6951,N_4052,N_1009);
nor U6952 (N_6952,N_2325,N_4469);
nor U6953 (N_6953,N_3154,N_5371);
nand U6954 (N_6954,N_3026,N_5046);
nor U6955 (N_6955,N_1287,N_3397);
and U6956 (N_6956,N_273,N_342);
and U6957 (N_6957,N_1394,N_655);
and U6958 (N_6958,N_695,N_116);
or U6959 (N_6959,N_5643,N_52);
nor U6960 (N_6960,N_5795,N_1192);
or U6961 (N_6961,N_1365,N_1132);
and U6962 (N_6962,N_2997,N_2650);
nand U6963 (N_6963,N_311,N_4180);
nand U6964 (N_6964,N_507,N_5704);
or U6965 (N_6965,N_1573,N_484);
and U6966 (N_6966,N_3032,N_2371);
nor U6967 (N_6967,N_1629,N_5263);
or U6968 (N_6968,N_4194,N_942);
or U6969 (N_6969,N_26,N_1831);
or U6970 (N_6970,N_3962,N_2165);
or U6971 (N_6971,N_4942,N_3144);
nand U6972 (N_6972,N_1236,N_2002);
and U6973 (N_6973,N_3002,N_4187);
nor U6974 (N_6974,N_360,N_367);
and U6975 (N_6975,N_2156,N_5203);
and U6976 (N_6976,N_1661,N_3720);
or U6977 (N_6977,N_62,N_1998);
xor U6978 (N_6978,N_541,N_3464);
nor U6979 (N_6979,N_1754,N_6142);
or U6980 (N_6980,N_4210,N_3452);
xor U6981 (N_6981,N_1341,N_3783);
or U6982 (N_6982,N_4476,N_2592);
and U6983 (N_6983,N_5409,N_2986);
nor U6984 (N_6984,N_1490,N_1402);
nand U6985 (N_6985,N_1860,N_5992);
nor U6986 (N_6986,N_1965,N_5650);
and U6987 (N_6987,N_4393,N_3531);
nor U6988 (N_6988,N_5635,N_4262);
nand U6989 (N_6989,N_70,N_6220);
nand U6990 (N_6990,N_4764,N_1670);
nor U6991 (N_6991,N_1641,N_225);
nand U6992 (N_6992,N_4880,N_3598);
nor U6993 (N_6993,N_2843,N_1596);
xnor U6994 (N_6994,N_611,N_3338);
and U6995 (N_6995,N_5685,N_4418);
nor U6996 (N_6996,N_4229,N_25);
and U6997 (N_6997,N_2212,N_6215);
nand U6998 (N_6998,N_6242,N_1032);
xnor U6999 (N_6999,N_4490,N_488);
and U7000 (N_7000,N_219,N_1875);
xnor U7001 (N_7001,N_1719,N_2911);
xor U7002 (N_7002,N_5073,N_3294);
and U7003 (N_7003,N_5440,N_2335);
and U7004 (N_7004,N_5854,N_43);
and U7005 (N_7005,N_4676,N_2806);
xnor U7006 (N_7006,N_2845,N_5478);
xnor U7007 (N_7007,N_443,N_2318);
or U7008 (N_7008,N_5056,N_1401);
nand U7009 (N_7009,N_2492,N_10);
nand U7010 (N_7010,N_5981,N_918);
or U7011 (N_7011,N_3231,N_709);
nand U7012 (N_7012,N_1855,N_3527);
nand U7013 (N_7013,N_4098,N_1296);
xnor U7014 (N_7014,N_1357,N_2644);
and U7015 (N_7015,N_1138,N_459);
xnor U7016 (N_7016,N_3797,N_4623);
nor U7017 (N_7017,N_2653,N_2131);
nand U7018 (N_7018,N_2022,N_245);
nor U7019 (N_7019,N_1703,N_2880);
xnor U7020 (N_7020,N_90,N_721);
nand U7021 (N_7021,N_4520,N_1397);
xor U7022 (N_7022,N_6226,N_532);
nor U7023 (N_7023,N_1039,N_1439);
nor U7024 (N_7024,N_3145,N_5833);
or U7025 (N_7025,N_95,N_2833);
or U7026 (N_7026,N_2330,N_6131);
or U7027 (N_7027,N_3124,N_3412);
xnor U7028 (N_7028,N_1607,N_5078);
xnor U7029 (N_7029,N_4588,N_3821);
nor U7030 (N_7030,N_5559,N_5960);
or U7031 (N_7031,N_5967,N_2061);
or U7032 (N_7032,N_3504,N_1631);
xnor U7033 (N_7033,N_3207,N_376);
nand U7034 (N_7034,N_2198,N_677);
nand U7035 (N_7035,N_1289,N_781);
and U7036 (N_7036,N_3171,N_4589);
nand U7037 (N_7037,N_1896,N_3284);
xor U7038 (N_7038,N_2803,N_1718);
nand U7039 (N_7039,N_1290,N_1503);
and U7040 (N_7040,N_6019,N_247);
nor U7041 (N_7041,N_2062,N_5785);
xor U7042 (N_7042,N_36,N_2004);
nor U7043 (N_7043,N_700,N_3826);
nor U7044 (N_7044,N_1929,N_4289);
or U7045 (N_7045,N_345,N_76);
and U7046 (N_7046,N_5109,N_830);
nor U7047 (N_7047,N_1112,N_1788);
or U7048 (N_7048,N_3633,N_1859);
nand U7049 (N_7049,N_6189,N_4999);
xor U7050 (N_7050,N_2582,N_5585);
and U7051 (N_7051,N_1247,N_3275);
or U7052 (N_7052,N_558,N_5249);
and U7053 (N_7053,N_2174,N_5319);
or U7054 (N_7054,N_4882,N_4967);
nand U7055 (N_7055,N_5740,N_527);
or U7056 (N_7056,N_5604,N_3558);
or U7057 (N_7057,N_4818,N_4188);
and U7058 (N_7058,N_2259,N_4364);
nor U7059 (N_7059,N_2077,N_1482);
xnor U7060 (N_7060,N_2359,N_544);
nand U7061 (N_7061,N_5384,N_992);
nor U7062 (N_7062,N_504,N_2464);
and U7063 (N_7063,N_170,N_5541);
nand U7064 (N_7064,N_1781,N_4955);
or U7065 (N_7065,N_4629,N_411);
and U7066 (N_7066,N_3348,N_1969);
xnor U7067 (N_7067,N_1616,N_50);
or U7068 (N_7068,N_2775,N_1622);
nor U7069 (N_7069,N_3891,N_3549);
nand U7070 (N_7070,N_1619,N_4648);
xor U7071 (N_7071,N_2926,N_3319);
and U7072 (N_7072,N_5153,N_303);
and U7073 (N_7073,N_3942,N_5150);
and U7074 (N_7074,N_2938,N_1838);
and U7075 (N_7075,N_2674,N_2550);
xnor U7076 (N_7076,N_537,N_5673);
and U7077 (N_7077,N_452,N_4286);
and U7078 (N_7078,N_1732,N_4164);
nand U7079 (N_7079,N_199,N_4454);
xor U7080 (N_7080,N_3143,N_3087);
xor U7081 (N_7081,N_817,N_3537);
nor U7082 (N_7082,N_2962,N_1165);
xor U7083 (N_7083,N_2934,N_2904);
and U7084 (N_7084,N_4387,N_2420);
nand U7085 (N_7085,N_3716,N_122);
nor U7086 (N_7086,N_1366,N_1494);
nor U7087 (N_7087,N_832,N_4930);
nand U7088 (N_7088,N_3637,N_5702);
nor U7089 (N_7089,N_4642,N_4012);
or U7090 (N_7090,N_1826,N_4508);
or U7091 (N_7091,N_1882,N_4743);
and U7092 (N_7092,N_466,N_2946);
nor U7093 (N_7093,N_281,N_127);
and U7094 (N_7094,N_4483,N_3551);
nor U7095 (N_7095,N_2824,N_4282);
nor U7096 (N_7096,N_4104,N_4195);
or U7097 (N_7097,N_920,N_5323);
or U7098 (N_7098,N_2370,N_4581);
nand U7099 (N_7099,N_2382,N_972);
or U7100 (N_7100,N_4329,N_2506);
xor U7101 (N_7101,N_2619,N_1682);
nor U7102 (N_7102,N_5600,N_4798);
and U7103 (N_7103,N_344,N_3077);
xor U7104 (N_7104,N_2000,N_740);
nor U7105 (N_7105,N_1461,N_5952);
nand U7106 (N_7106,N_4848,N_6050);
nand U7107 (N_7107,N_739,N_5621);
and U7108 (N_7108,N_5636,N_1336);
nand U7109 (N_7109,N_5451,N_6102);
and U7110 (N_7110,N_3727,N_671);
or U7111 (N_7111,N_1999,N_4191);
or U7112 (N_7112,N_1225,N_5221);
nand U7113 (N_7113,N_16,N_4441);
nor U7114 (N_7114,N_2213,N_260);
nand U7115 (N_7115,N_5647,N_2143);
nand U7116 (N_7116,N_2580,N_5202);
and U7117 (N_7117,N_3117,N_4360);
xor U7118 (N_7118,N_6025,N_2537);
and U7119 (N_7119,N_1183,N_2161);
xnor U7120 (N_7120,N_1222,N_2186);
or U7121 (N_7121,N_5889,N_1748);
or U7122 (N_7122,N_4554,N_3646);
or U7123 (N_7123,N_5299,N_2922);
and U7124 (N_7124,N_593,N_1721);
and U7125 (N_7125,N_1330,N_4505);
xor U7126 (N_7126,N_5966,N_2790);
nor U7127 (N_7127,N_2265,N_3548);
nand U7128 (N_7128,N_2527,N_4797);
xnor U7129 (N_7129,N_1140,N_3300);
nand U7130 (N_7130,N_4979,N_2047);
and U7131 (N_7131,N_912,N_5292);
nor U7132 (N_7132,N_4394,N_4935);
and U7133 (N_7133,N_2757,N_1160);
xor U7134 (N_7134,N_2718,N_4617);
nand U7135 (N_7135,N_4413,N_3116);
nand U7136 (N_7136,N_5364,N_5051);
nand U7137 (N_7137,N_5676,N_103);
xnor U7138 (N_7138,N_1637,N_784);
and U7139 (N_7139,N_2675,N_2799);
or U7140 (N_7140,N_764,N_4380);
xnor U7141 (N_7141,N_5537,N_2254);
nor U7142 (N_7142,N_138,N_1534);
nand U7143 (N_7143,N_2615,N_399);
xnor U7144 (N_7144,N_640,N_4302);
or U7145 (N_7145,N_4142,N_2235);
and U7146 (N_7146,N_161,N_1319);
or U7147 (N_7147,N_4920,N_545);
nor U7148 (N_7148,N_4712,N_6195);
or U7149 (N_7149,N_524,N_1978);
nor U7150 (N_7150,N_1600,N_1636);
nand U7151 (N_7151,N_5567,N_3746);
and U7152 (N_7152,N_6129,N_2030);
nor U7153 (N_7153,N_5645,N_4963);
xnor U7154 (N_7154,N_6234,N_4429);
nor U7155 (N_7155,N_4506,N_4911);
nor U7156 (N_7156,N_4171,N_1232);
or U7157 (N_7157,N_2856,N_1680);
and U7158 (N_7158,N_4804,N_5556);
and U7159 (N_7159,N_1484,N_5728);
nor U7160 (N_7160,N_3365,N_1994);
xnor U7161 (N_7161,N_2478,N_2739);
nand U7162 (N_7162,N_4793,N_1762);
nor U7163 (N_7163,N_2462,N_5884);
nor U7164 (N_7164,N_3948,N_2699);
xnor U7165 (N_7165,N_3983,N_5891);
xnor U7166 (N_7166,N_2781,N_3024);
or U7167 (N_7167,N_4872,N_5103);
or U7168 (N_7168,N_1667,N_424);
nand U7169 (N_7169,N_4710,N_2292);
xor U7170 (N_7170,N_945,N_3856);
or U7171 (N_7171,N_4078,N_1466);
or U7172 (N_7172,N_3500,N_4913);
nand U7173 (N_7173,N_5729,N_4037);
or U7174 (N_7174,N_5707,N_3156);
nor U7175 (N_7175,N_5792,N_694);
nand U7176 (N_7176,N_5734,N_4869);
nand U7177 (N_7177,N_3568,N_3137);
and U7178 (N_7178,N_4231,N_2009);
and U7179 (N_7179,N_5753,N_4433);
or U7180 (N_7180,N_1066,N_1042);
or U7181 (N_7181,N_4879,N_2998);
and U7182 (N_7182,N_3364,N_272);
nand U7183 (N_7183,N_1829,N_99);
nand U7184 (N_7184,N_811,N_2041);
xnor U7185 (N_7185,N_5566,N_5668);
and U7186 (N_7186,N_533,N_4823);
nand U7187 (N_7187,N_1753,N_5955);
or U7188 (N_7188,N_2438,N_2496);
and U7189 (N_7189,N_1333,N_2855);
xor U7190 (N_7190,N_2430,N_1161);
nor U7191 (N_7191,N_2981,N_5064);
or U7192 (N_7192,N_616,N_6156);
nand U7193 (N_7193,N_5002,N_5301);
nor U7194 (N_7194,N_1387,N_20);
nand U7195 (N_7195,N_1464,N_1530);
xor U7196 (N_7196,N_293,N_1509);
nor U7197 (N_7197,N_1706,N_4090);
and U7198 (N_7198,N_3040,N_2340);
xnor U7199 (N_7199,N_5926,N_5242);
and U7200 (N_7200,N_1520,N_6204);
nand U7201 (N_7201,N_5111,N_3614);
and U7202 (N_7202,N_3486,N_5005);
nand U7203 (N_7203,N_738,N_4674);
xnor U7204 (N_7204,N_3331,N_5632);
xnor U7205 (N_7205,N_810,N_4167);
nand U7206 (N_7206,N_3080,N_2053);
or U7207 (N_7207,N_3980,N_2183);
nor U7208 (N_7208,N_2886,N_543);
xor U7209 (N_7209,N_2416,N_3657);
and U7210 (N_7210,N_5767,N_6117);
or U7211 (N_7211,N_750,N_4997);
nor U7212 (N_7212,N_355,N_5231);
and U7213 (N_7213,N_2982,N_2839);
and U7214 (N_7214,N_1428,N_1750);
nand U7215 (N_7215,N_4339,N_4279);
nor U7216 (N_7216,N_3458,N_1679);
and U7217 (N_7217,N_178,N_5369);
nand U7218 (N_7218,N_1105,N_1692);
nor U7219 (N_7219,N_487,N_559);
and U7220 (N_7220,N_4326,N_1737);
or U7221 (N_7221,N_5273,N_4437);
nor U7222 (N_7222,N_3429,N_5530);
nand U7223 (N_7223,N_3023,N_4410);
xor U7224 (N_7224,N_363,N_4785);
nand U7225 (N_7225,N_2991,N_5847);
nor U7226 (N_7226,N_960,N_898);
nor U7227 (N_7227,N_3775,N_5773);
and U7228 (N_7228,N_1045,N_581);
or U7229 (N_7229,N_2603,N_925);
nand U7230 (N_7230,N_6095,N_5332);
xor U7231 (N_7231,N_628,N_5243);
or U7232 (N_7232,N_5450,N_2239);
nand U7233 (N_7233,N_976,N_927);
xnor U7234 (N_7234,N_3786,N_2918);
or U7235 (N_7235,N_4082,N_1089);
nor U7236 (N_7236,N_1973,N_1495);
xnor U7237 (N_7237,N_2192,N_909);
and U7238 (N_7238,N_4737,N_3578);
nand U7239 (N_7239,N_2306,N_5674);
nor U7240 (N_7240,N_3986,N_11);
or U7241 (N_7241,N_5244,N_779);
nand U7242 (N_7242,N_2063,N_4593);
or U7243 (N_7243,N_4852,N_2388);
and U7244 (N_7244,N_4248,N_2605);
and U7245 (N_7245,N_888,N_2630);
nor U7246 (N_7246,N_3167,N_2381);
or U7247 (N_7247,N_5250,N_5811);
nand U7248 (N_7248,N_2551,N_2627);
xor U7249 (N_7249,N_4939,N_2995);
nor U7250 (N_7250,N_6118,N_682);
and U7251 (N_7251,N_4644,N_2567);
and U7252 (N_7252,N_3027,N_3118);
and U7253 (N_7253,N_5333,N_2512);
or U7254 (N_7254,N_1076,N_3514);
or U7255 (N_7255,N_4832,N_4552);
xor U7256 (N_7256,N_5020,N_827);
xnor U7257 (N_7257,N_1856,N_1362);
nand U7258 (N_7258,N_4971,N_3669);
nor U7259 (N_7259,N_3426,N_4656);
xnor U7260 (N_7260,N_6090,N_2005);
xor U7261 (N_7261,N_1256,N_967);
xnor U7262 (N_7262,N_3553,N_1759);
nand U7263 (N_7263,N_3189,N_5769);
and U7264 (N_7264,N_4618,N_1398);
nand U7265 (N_7265,N_5131,N_4820);
or U7266 (N_7266,N_4592,N_2091);
xnor U7267 (N_7267,N_2521,N_5098);
or U7268 (N_7268,N_249,N_5013);
nor U7269 (N_7269,N_5081,N_2138);
nand U7270 (N_7270,N_3723,N_1612);
and U7271 (N_7271,N_2202,N_4330);
nor U7272 (N_7272,N_4816,N_3642);
xor U7273 (N_7273,N_4613,N_211);
and U7274 (N_7274,N_5127,N_5742);
nand U7275 (N_7275,N_2658,N_2877);
nand U7276 (N_7276,N_5055,N_3951);
nor U7277 (N_7277,N_4416,N_2955);
xnor U7278 (N_7278,N_4023,N_5997);
or U7279 (N_7279,N_4871,N_5087);
nand U7280 (N_7280,N_2557,N_4502);
or U7281 (N_7281,N_4321,N_6202);
xor U7282 (N_7282,N_5505,N_2320);
and U7283 (N_7283,N_2864,N_3761);
nand U7284 (N_7284,N_3541,N_4368);
or U7285 (N_7285,N_2436,N_5481);
and U7286 (N_7286,N_4127,N_4547);
and U7287 (N_7287,N_2740,N_1238);
nor U7288 (N_7288,N_5251,N_4549);
and U7289 (N_7289,N_3683,N_3571);
nand U7290 (N_7290,N_2324,N_4605);
nor U7291 (N_7291,N_6180,N_615);
nor U7292 (N_7292,N_5701,N_1653);
or U7293 (N_7293,N_2200,N_4049);
and U7294 (N_7294,N_1854,N_3089);
nor U7295 (N_7295,N_83,N_3336);
and U7296 (N_7296,N_1050,N_3976);
or U7297 (N_7297,N_4700,N_1452);
nor U7298 (N_7298,N_5400,N_5611);
xor U7299 (N_7299,N_5261,N_1400);
xor U7300 (N_7300,N_265,N_959);
and U7301 (N_7301,N_3898,N_4063);
or U7302 (N_7302,N_3995,N_4154);
or U7303 (N_7303,N_3837,N_5342);
nand U7304 (N_7304,N_429,N_2431);
nand U7305 (N_7305,N_5000,N_1145);
and U7306 (N_7306,N_2336,N_1124);
xnor U7307 (N_7307,N_1957,N_4438);
nand U7308 (N_7308,N_77,N_5597);
nand U7309 (N_7309,N_92,N_5890);
nand U7310 (N_7310,N_6140,N_4228);
xnor U7311 (N_7311,N_2711,N_121);
xnor U7312 (N_7312,N_4009,N_3011);
or U7313 (N_7313,N_5945,N_4796);
or U7314 (N_7314,N_4821,N_5309);
xor U7315 (N_7315,N_4328,N_6149);
xnor U7316 (N_7316,N_6159,N_2348);
or U7317 (N_7317,N_2214,N_3299);
nand U7318 (N_7318,N_3436,N_1008);
nor U7319 (N_7319,N_886,N_6196);
and U7320 (N_7320,N_2216,N_3597);
nor U7321 (N_7321,N_4690,N_5259);
nand U7322 (N_7322,N_5378,N_2641);
xor U7323 (N_7323,N_5156,N_1704);
or U7324 (N_7324,N_2372,N_4193);
nor U7325 (N_7325,N_5899,N_954);
xnor U7326 (N_7326,N_3928,N_5239);
and U7327 (N_7327,N_4432,N_3523);
xor U7328 (N_7328,N_349,N_3934);
xor U7329 (N_7329,N_4718,N_5984);
nor U7330 (N_7330,N_2598,N_1634);
and U7331 (N_7331,N_2271,N_836);
xnor U7332 (N_7332,N_5572,N_1368);
or U7333 (N_7333,N_5264,N_308);
or U7334 (N_7334,N_1518,N_4978);
or U7335 (N_7335,N_4341,N_2941);
and U7336 (N_7336,N_6023,N_2752);
xnor U7337 (N_7337,N_1675,N_5662);
and U7338 (N_7338,N_1061,N_5711);
nor U7339 (N_7339,N_183,N_2516);
or U7340 (N_7340,N_330,N_191);
and U7341 (N_7341,N_2098,N_1707);
nor U7342 (N_7342,N_1437,N_793);
nand U7343 (N_7343,N_79,N_4566);
xor U7344 (N_7344,N_2467,N_5790);
or U7345 (N_7345,N_160,N_2670);
nor U7346 (N_7346,N_2847,N_430);
nor U7347 (N_7347,N_2990,N_1689);
or U7348 (N_7348,N_531,N_5774);
xor U7349 (N_7349,N_3745,N_5039);
nand U7350 (N_7350,N_1070,N_3279);
nor U7351 (N_7351,N_2374,N_5310);
or U7352 (N_7352,N_5503,N_1205);
nor U7353 (N_7353,N_2520,N_4591);
nor U7354 (N_7354,N_2765,N_3396);
nand U7355 (N_7355,N_1733,N_1316);
or U7356 (N_7356,N_1674,N_3213);
nand U7357 (N_7357,N_5630,N_3701);
or U7358 (N_7358,N_5396,N_2176);
and U7359 (N_7359,N_2965,N_5532);
and U7360 (N_7360,N_1372,N_3248);
nand U7361 (N_7361,N_6065,N_2628);
and U7362 (N_7362,N_519,N_5278);
or U7363 (N_7363,N_1917,N_1960);
xor U7364 (N_7364,N_4214,N_3421);
nor U7365 (N_7365,N_56,N_3670);
and U7366 (N_7366,N_2756,N_4428);
or U7367 (N_7367,N_4532,N_4587);
xor U7368 (N_7368,N_5402,N_3862);
nand U7369 (N_7369,N_902,N_4791);
or U7370 (N_7370,N_3352,N_334);
nand U7371 (N_7371,N_2051,N_3398);
nor U7372 (N_7372,N_4204,N_254);
nor U7373 (N_7373,N_953,N_1932);
nor U7374 (N_7374,N_5758,N_2910);
xor U7375 (N_7375,N_1299,N_3402);
or U7376 (N_7376,N_5804,N_5771);
nor U7377 (N_7377,N_2410,N_1625);
xnor U7378 (N_7378,N_785,N_579);
xor U7379 (N_7379,N_3206,N_4492);
nor U7380 (N_7380,N_306,N_3155);
xnor U7381 (N_7381,N_5235,N_3706);
nand U7382 (N_7382,N_4239,N_2534);
or U7383 (N_7383,N_3070,N_5607);
and U7384 (N_7384,N_4778,N_2940);
xnor U7385 (N_7385,N_449,N_1006);
nand U7386 (N_7386,N_4092,N_2678);
and U7387 (N_7387,N_5155,N_4151);
or U7388 (N_7388,N_2207,N_1722);
nor U7389 (N_7389,N_620,N_1308);
or U7390 (N_7390,N_1278,N_629);
and U7391 (N_7391,N_4281,N_3052);
nand U7392 (N_7392,N_648,N_1935);
and U7393 (N_7393,N_5972,N_1647);
nand U7394 (N_7394,N_289,N_643);
and U7395 (N_7395,N_548,N_5938);
or U7396 (N_7396,N_4553,N_5303);
xor U7397 (N_7397,N_5211,N_1493);
xor U7398 (N_7398,N_962,N_803);
xnor U7399 (N_7399,N_2274,N_1369);
nor U7400 (N_7400,N_1874,N_660);
and U7401 (N_7401,N_3141,N_4576);
xor U7402 (N_7402,N_3325,N_2751);
nor U7403 (N_7403,N_1094,N_5501);
xnor U7404 (N_7404,N_427,N_2529);
xor U7405 (N_7405,N_2867,N_177);
xor U7406 (N_7406,N_2841,N_4284);
xor U7407 (N_7407,N_3648,N_147);
nor U7408 (N_7408,N_4776,N_2936);
xor U7409 (N_7409,N_3191,N_6009);
or U7410 (N_7410,N_4124,N_4287);
nor U7411 (N_7411,N_280,N_2590);
xnor U7412 (N_7412,N_2903,N_4988);
nor U7413 (N_7413,N_3259,N_3263);
xnor U7414 (N_7414,N_1470,N_3940);
nor U7415 (N_7415,N_2931,N_106);
or U7416 (N_7416,N_5037,N_4986);
nand U7417 (N_7417,N_3104,N_1528);
nor U7418 (N_7418,N_2552,N_5637);
and U7419 (N_7419,N_930,N_3749);
xnor U7420 (N_7420,N_3773,N_3184);
nand U7421 (N_7421,N_154,N_2305);
nand U7422 (N_7422,N_3747,N_4011);
xor U7423 (N_7423,N_523,N_1367);
or U7424 (N_7424,N_1900,N_4263);
or U7425 (N_7425,N_2945,N_906);
and U7426 (N_7426,N_3413,N_5158);
nor U7427 (N_7427,N_3460,N_991);
nor U7428 (N_7428,N_5300,N_4750);
and U7429 (N_7429,N_1084,N_3702);
nand U7430 (N_7430,N_6207,N_4269);
xnor U7431 (N_7431,N_2314,N_6139);
nand U7432 (N_7432,N_6010,N_5879);
or U7433 (N_7433,N_1513,N_7);
xor U7434 (N_7434,N_6020,N_3827);
nor U7435 (N_7435,N_1832,N_4551);
nor U7436 (N_7436,N_462,N_3843);
xor U7437 (N_7437,N_2346,N_1154);
nand U7438 (N_7438,N_2526,N_2023);
and U7439 (N_7439,N_1162,N_998);
and U7440 (N_7440,N_171,N_15);
nor U7441 (N_7441,N_1321,N_4117);
or U7442 (N_7442,N_2924,N_1186);
or U7443 (N_7443,N_4603,N_3935);
nor U7444 (N_7444,N_1343,N_4657);
or U7445 (N_7445,N_2616,N_681);
nand U7446 (N_7446,N_1902,N_534);
nor U7447 (N_7447,N_520,N_2709);
xor U7448 (N_7448,N_4033,N_2816);
nor U7449 (N_7449,N_2610,N_3416);
nand U7450 (N_7450,N_5746,N_1553);
nand U7451 (N_7451,N_2007,N_1021);
nor U7452 (N_7452,N_4885,N_5622);
and U7453 (N_7453,N_3585,N_2240);
and U7454 (N_7454,N_1545,N_5318);
nor U7455 (N_7455,N_234,N_829);
nor U7456 (N_7456,N_1469,N_68);
and U7457 (N_7457,N_1519,N_5411);
nand U7458 (N_7458,N_4596,N_3066);
or U7459 (N_7459,N_1821,N_1488);
or U7460 (N_7460,N_3719,N_3197);
and U7461 (N_7461,N_3893,N_1155);
nor U7462 (N_7462,N_3518,N_4639);
nor U7463 (N_7463,N_3383,N_2479);
xor U7464 (N_7464,N_1191,N_5038);
nor U7465 (N_7465,N_1073,N_2869);
xnor U7466 (N_7466,N_5052,N_5285);
nor U7467 (N_7467,N_4675,N_1475);
xnor U7468 (N_7468,N_3414,N_1966);
xnor U7469 (N_7469,N_2448,N_2142);
nor U7470 (N_7470,N_5044,N_5490);
xnor U7471 (N_7471,N_2360,N_2270);
xnor U7472 (N_7472,N_1910,N_5029);
or U7473 (N_7473,N_82,N_1849);
xor U7474 (N_7474,N_1059,N_6182);
or U7475 (N_7475,N_1379,N_5594);
or U7476 (N_7476,N_563,N_264);
nor U7477 (N_7477,N_3774,N_4405);
nand U7478 (N_7478,N_575,N_3459);
or U7479 (N_7479,N_4903,N_1560);
nand U7480 (N_7480,N_4123,N_5666);
or U7481 (N_7481,N_3389,N_5427);
xnor U7482 (N_7482,N_3937,N_4822);
nand U7483 (N_7483,N_5216,N_1416);
nand U7484 (N_7484,N_3524,N_642);
xor U7485 (N_7485,N_4333,N_4856);
nor U7486 (N_7486,N_3697,N_5982);
nor U7487 (N_7487,N_5110,N_5266);
nand U7488 (N_7488,N_2768,N_6185);
nor U7489 (N_7489,N_3366,N_3522);
nand U7490 (N_7490,N_1496,N_2112);
nor U7491 (N_7491,N_6176,N_1642);
and U7492 (N_7492,N_3620,N_1104);
or U7493 (N_7493,N_3973,N_2762);
and U7494 (N_7494,N_5381,N_4395);
nor U7495 (N_7495,N_877,N_6229);
nor U7496 (N_7496,N_4992,N_3119);
nand U7497 (N_7497,N_1450,N_2974);
nor U7498 (N_7498,N_5733,N_5552);
xor U7499 (N_7499,N_3735,N_2920);
nand U7500 (N_7500,N_3991,N_3602);
and U7501 (N_7501,N_867,N_4032);
nand U7502 (N_7502,N_4735,N_4369);
and U7503 (N_7503,N_3305,N_266);
or U7504 (N_7504,N_503,N_2745);
xnor U7505 (N_7505,N_1613,N_2283);
xnor U7506 (N_7506,N_678,N_1345);
xnor U7507 (N_7507,N_59,N_5200);
nand U7508 (N_7508,N_5677,N_2460);
nor U7509 (N_7509,N_1157,N_1755);
or U7510 (N_7510,N_4991,N_1033);
or U7511 (N_7511,N_2159,N_5961);
nor U7512 (N_7512,N_3782,N_5101);
nand U7513 (N_7513,N_1390,N_2373);
xnor U7514 (N_7514,N_4143,N_3289);
and U7515 (N_7515,N_337,N_719);
and U7516 (N_7516,N_5959,N_2951);
and U7517 (N_7517,N_1822,N_1312);
nor U7518 (N_7518,N_4147,N_1720);
or U7519 (N_7519,N_124,N_3984);
nor U7520 (N_7520,N_690,N_5031);
and U7521 (N_7521,N_2971,N_3874);
xnor U7522 (N_7522,N_3387,N_352);
xnor U7523 (N_7523,N_3679,N_4107);
or U7524 (N_7524,N_3956,N_3433);
and U7525 (N_7525,N_2949,N_3456);
and U7526 (N_7526,N_4112,N_1173);
and U7527 (N_7527,N_1385,N_4371);
xnor U7528 (N_7528,N_2334,N_5422);
nor U7529 (N_7529,N_2338,N_1038);
and U7530 (N_7530,N_4813,N_3678);
nor U7531 (N_7531,N_3214,N_5837);
nor U7532 (N_7532,N_4179,N_2166);
or U7533 (N_7533,N_1583,N_2315);
and U7534 (N_7534,N_1758,N_4381);
and U7535 (N_7535,N_821,N_5908);
xor U7536 (N_7536,N_1666,N_111);
or U7537 (N_7537,N_661,N_4342);
nand U7538 (N_7538,N_4701,N_4002);
nor U7539 (N_7539,N_5782,N_2914);
xnor U7540 (N_7540,N_3645,N_6084);
nand U7541 (N_7541,N_4336,N_2444);
nor U7542 (N_7542,N_693,N_4975);
and U7543 (N_7543,N_5710,N_6187);
nand U7544 (N_7544,N_1615,N_1800);
xor U7545 (N_7545,N_1279,N_34);
and U7546 (N_7546,N_4044,N_5497);
nand U7547 (N_7547,N_3538,N_338);
or U7548 (N_7548,N_2067,N_3809);
nand U7549 (N_7549,N_6120,N_6203);
xnor U7550 (N_7550,N_4767,N_5126);
nor U7551 (N_7551,N_3345,N_4899);
nand U7552 (N_7552,N_2969,N_3151);
nor U7553 (N_7553,N_5096,N_1031);
and U7554 (N_7554,N_5695,N_6214);
nor U7555 (N_7555,N_2726,N_5353);
nor U7556 (N_7556,N_4470,N_3301);
and U7557 (N_7557,N_3741,N_5448);
nand U7558 (N_7558,N_2037,N_4572);
and U7559 (N_7559,N_1853,N_1410);
or U7560 (N_7560,N_3981,N_2150);
xor U7561 (N_7561,N_1164,N_4384);
nor U7562 (N_7562,N_4707,N_3853);
nor U7563 (N_7563,N_4970,N_2057);
and U7564 (N_7564,N_2602,N_4683);
and U7565 (N_7565,N_731,N_1456);
and U7566 (N_7566,N_4367,N_5780);
or U7567 (N_7567,N_1760,N_28);
nand U7568 (N_7568,N_716,N_2008);
and U7569 (N_7569,N_4048,N_5343);
xnor U7570 (N_7570,N_4374,N_5041);
and U7571 (N_7571,N_2033,N_5413);
and U7572 (N_7572,N_4510,N_2491);
and U7573 (N_7573,N_654,N_5053);
or U7574 (N_7574,N_3483,N_862);
xor U7575 (N_7575,N_3634,N_1426);
or U7576 (N_7576,N_5946,N_3822);
or U7577 (N_7577,N_2531,N_3400);
and U7578 (N_7578,N_39,N_3062);
nor U7579 (N_7579,N_1477,N_1581);
xnor U7580 (N_7580,N_5404,N_5933);
or U7581 (N_7581,N_5692,N_21);
xnor U7582 (N_7582,N_1742,N_2449);
and U7583 (N_7583,N_2963,N_4960);
and U7584 (N_7584,N_3229,N_193);
nand U7585 (N_7585,N_3911,N_5437);
nand U7586 (N_7586,N_1313,N_4538);
and U7587 (N_7587,N_1533,N_5321);
nand U7588 (N_7588,N_277,N_3047);
and U7589 (N_7589,N_2399,N_1614);
and U7590 (N_7590,N_1204,N_5372);
nor U7591 (N_7591,N_4715,N_1098);
xnor U7592 (N_7592,N_1309,N_148);
xor U7593 (N_7593,N_169,N_2659);
xnor U7594 (N_7594,N_185,N_3477);
or U7595 (N_7595,N_3274,N_608);
nor U7596 (N_7596,N_2721,N_2126);
nand U7597 (N_7597,N_613,N_675);
nand U7598 (N_7598,N_4493,N_1582);
xor U7599 (N_7599,N_4660,N_1122);
or U7600 (N_7600,N_5184,N_5106);
xor U7601 (N_7601,N_831,N_4575);
xnor U7602 (N_7602,N_5116,N_2548);
and U7603 (N_7603,N_5008,N_5817);
nor U7604 (N_7604,N_5656,N_2660);
or U7605 (N_7605,N_6211,N_3892);
nor U7606 (N_7606,N_1430,N_3789);
and U7607 (N_7607,N_450,N_6198);
nand U7608 (N_7608,N_6056,N_1229);
xnor U7609 (N_7609,N_4795,N_5730);
xnor U7610 (N_7610,N_3709,N_2723);
nor U7611 (N_7611,N_2220,N_1188);
nand U7612 (N_7612,N_5670,N_4385);
nand U7613 (N_7613,N_2199,N_4067);
nand U7614 (N_7614,N_706,N_480);
xor U7615 (N_7615,N_6008,N_1206);
or U7616 (N_7616,N_4299,N_1353);
nor U7617 (N_7617,N_5968,N_496);
nand U7618 (N_7618,N_4144,N_386);
nand U7619 (N_7619,N_5818,N_555);
or U7620 (N_7620,N_5750,N_382);
or U7621 (N_7621,N_5978,N_4034);
xor U7622 (N_7622,N_361,N_3977);
xor U7623 (N_7623,N_335,N_1694);
nand U7624 (N_7624,N_1429,N_670);
nand U7625 (N_7625,N_5725,N_354);
nand U7626 (N_7626,N_1603,N_2954);
or U7627 (N_7627,N_1453,N_3492);
or U7628 (N_7628,N_4533,N_1180);
and U7629 (N_7629,N_1198,N_1239);
nand U7630 (N_7630,N_4202,N_1610);
and U7631 (N_7631,N_1837,N_672);
or U7632 (N_7632,N_3193,N_6241);
or U7633 (N_7633,N_3340,N_1567);
nand U7634 (N_7634,N_5088,N_4297);
nand U7635 (N_7635,N_181,N_4697);
nand U7636 (N_7636,N_5832,N_2811);
nor U7637 (N_7637,N_6029,N_2892);
and U7638 (N_7638,N_4812,N_1415);
nor U7639 (N_7639,N_4120,N_4105);
xnor U7640 (N_7640,N_698,N_4917);
and U7641 (N_7641,N_4625,N_3220);
and U7642 (N_7642,N_528,N_3031);
nor U7643 (N_7643,N_3590,N_1123);
and U7644 (N_7644,N_464,N_5206);
nand U7645 (N_7645,N_5595,N_5204);
nand U7646 (N_7646,N_1114,N_1041);
xor U7647 (N_7647,N_2291,N_820);
xor U7648 (N_7648,N_6132,N_1233);
nor U7649 (N_7649,N_4590,N_4346);
or U7650 (N_7650,N_2623,N_3894);
and U7651 (N_7651,N_2014,N_4445);
nor U7652 (N_7652,N_4968,N_476);
nor U7653 (N_7653,N_5399,N_243);
or U7654 (N_7654,N_5810,N_5099);
nor U7655 (N_7655,N_2247,N_5405);
nor U7656 (N_7656,N_5100,N_2027);
or U7657 (N_7657,N_150,N_5141);
xor U7658 (N_7658,N_5864,N_3552);
or U7659 (N_7659,N_5613,N_623);
nor U7660 (N_7660,N_2132,N_5511);
nand U7661 (N_7661,N_2456,N_3907);
nand U7662 (N_7662,N_1980,N_4854);
or U7663 (N_7663,N_4730,N_5444);
nand U7664 (N_7664,N_3750,N_1315);
nand U7665 (N_7665,N_292,N_4753);
or U7666 (N_7666,N_2172,N_4650);
xor U7667 (N_7667,N_3408,N_5274);
xnor U7668 (N_7668,N_1941,N_5134);
and U7669 (N_7669,N_5626,N_871);
or U7670 (N_7670,N_108,N_679);
nor U7671 (N_7671,N_2742,N_5958);
nor U7672 (N_7672,N_2036,N_5255);
and U7673 (N_7673,N_23,N_4853);
nor U7674 (N_7674,N_1201,N_6209);
xor U7675 (N_7675,N_3082,N_542);
nand U7676 (N_7676,N_4241,N_2313);
xor U7677 (N_7677,N_769,N_973);
or U7678 (N_7678,N_5387,N_2298);
nor U7679 (N_7679,N_2357,N_2064);
or U7680 (N_7680,N_1529,N_673);
or U7681 (N_7681,N_5175,N_1909);
or U7682 (N_7682,N_5057,N_1139);
and U7683 (N_7683,N_1850,N_3619);
nand U7684 (N_7684,N_5236,N_5983);
nor U7685 (N_7685,N_951,N_2730);
or U7686 (N_7686,N_5456,N_4993);
nand U7687 (N_7687,N_6178,N_2565);
nand U7688 (N_7688,N_359,N_5380);
nor U7689 (N_7689,N_2137,N_4713);
or U7690 (N_7690,N_5664,N_4815);
nor U7691 (N_7691,N_3498,N_64);
or U7692 (N_7692,N_2406,N_3431);
xor U7693 (N_7693,N_1687,N_5132);
and U7694 (N_7694,N_4595,N_4773);
and U7695 (N_7695,N_1608,N_1079);
or U7696 (N_7696,N_6003,N_1329);
or U7697 (N_7697,N_2184,N_2849);
xnor U7698 (N_7698,N_1723,N_5189);
or U7699 (N_7699,N_4463,N_3632);
or U7700 (N_7700,N_2290,N_5252);
nand U7701 (N_7701,N_1532,N_316);
nor U7702 (N_7702,N_4560,N_2120);
nor U7703 (N_7703,N_6062,N_1901);
or U7704 (N_7704,N_5565,N_4671);
and U7705 (N_7705,N_3831,N_788);
nand U7706 (N_7706,N_319,N_1340);
or U7707 (N_7707,N_3450,N_950);
nor U7708 (N_7708,N_5551,N_607);
or U7709 (N_7709,N_1292,N_1877);
and U7710 (N_7710,N_1618,N_1237);
or U7711 (N_7711,N_4638,N_4883);
or U7712 (N_7712,N_5834,N_5855);
and U7713 (N_7713,N_2459,N_663);
nand U7714 (N_7714,N_151,N_407);
nor U7715 (N_7715,N_2746,N_2127);
or U7716 (N_7716,N_3394,N_4687);
xnor U7717 (N_7717,N_3666,N_2238);
nand U7718 (N_7718,N_5047,N_3271);
and U7719 (N_7719,N_223,N_4780);
nor U7720 (N_7720,N_1944,N_73);
or U7721 (N_7721,N_5950,N_4558);
xor U7722 (N_7722,N_4711,N_1399);
nor U7723 (N_7723,N_5874,N_631);
or U7724 (N_7724,N_3919,N_4511);
nand U7725 (N_7725,N_3638,N_4378);
or U7726 (N_7726,N_755,N_856);
nand U7727 (N_7727,N_2016,N_2606);
xor U7728 (N_7728,N_2119,N_1275);
nor U7729 (N_7729,N_5136,N_5893);
and U7730 (N_7730,N_2,N_5623);
nand U7731 (N_7731,N_5495,N_5112);
nand U7732 (N_7732,N_2331,N_847);
or U7733 (N_7733,N_2732,N_4362);
nand U7734 (N_7734,N_5609,N_3969);
nor U7735 (N_7735,N_652,N_1449);
nand U7736 (N_7736,N_4391,N_5142);
nand U7737 (N_7737,N_3326,N_3854);
or U7738 (N_7738,N_2221,N_2798);
nand U7739 (N_7739,N_5793,N_5083);
nand U7740 (N_7740,N_4616,N_5234);
xor U7741 (N_7741,N_482,N_6224);
xor U7742 (N_7742,N_3142,N_5026);
nand U7743 (N_7743,N_1937,N_1911);
or U7744 (N_7744,N_2837,N_1787);
nand U7745 (N_7745,N_5386,N_113);
xor U7746 (N_7746,N_4303,N_4026);
nand U7747 (N_7747,N_6005,N_4014);
nor U7748 (N_7748,N_2560,N_5356);
nand U7749 (N_7749,N_3997,N_2525);
and U7750 (N_7750,N_1085,N_634);
or U7751 (N_7751,N_5071,N_248);
and U7752 (N_7752,N_5128,N_4157);
xnor U7753 (N_7753,N_1996,N_4115);
or U7754 (N_7754,N_5140,N_656);
or U7755 (N_7755,N_1576,N_1243);
nor U7756 (N_7756,N_5523,N_1982);
nand U7757 (N_7757,N_3608,N_2141);
nor U7758 (N_7758,N_3149,N_1288);
nand U7759 (N_7759,N_6103,N_1918);
and U7760 (N_7760,N_5198,N_5065);
and U7761 (N_7761,N_4931,N_1705);
nand U7762 (N_7762,N_2408,N_6037);
nand U7763 (N_7763,N_6154,N_1505);
nand U7764 (N_7764,N_2094,N_384);
xnor U7765 (N_7765,N_5197,N_1260);
xor U7766 (N_7766,N_5756,N_5224);
nor U7767 (N_7767,N_3555,N_5911);
nor U7768 (N_7768,N_2976,N_3357);
nand U7769 (N_7769,N_2394,N_5268);
or U7770 (N_7770,N_4196,N_3252);
nor U7771 (N_7771,N_3830,N_6028);
nand U7772 (N_7772,N_5856,N_5107);
xnor U7773 (N_7773,N_4215,N_5738);
or U7774 (N_7774,N_808,N_878);
or U7775 (N_7775,N_1696,N_4461);
or U7776 (N_7776,N_5627,N_2902);
xor U7777 (N_7777,N_6200,N_3451);
and U7778 (N_7778,N_2956,N_275);
nor U7779 (N_7779,N_3848,N_1951);
nor U7780 (N_7780,N_1067,N_1905);
and U7781 (N_7781,N_4169,N_6116);
nor U7782 (N_7782,N_4372,N_4435);
and U7783 (N_7783,N_1460,N_5018);
nor U7784 (N_7784,N_4352,N_1906);
xnor U7785 (N_7785,N_3630,N_3953);
nor U7786 (N_7786,N_5640,N_2111);
nor U7787 (N_7787,N_3328,N_1096);
and U7788 (N_7788,N_3979,N_2777);
nand U7789 (N_7789,N_5828,N_4206);
and U7790 (N_7790,N_5421,N_1876);
nand U7791 (N_7791,N_4396,N_5282);
xnor U7792 (N_7792,N_5806,N_3810);
xor U7793 (N_7793,N_6232,N_2860);
nand U7794 (N_7794,N_696,N_5876);
and U7795 (N_7795,N_2717,N_4130);
or U7796 (N_7796,N_437,N_3812);
or U7797 (N_7797,N_294,N_2123);
xnor U7798 (N_7798,N_569,N_4983);
or U7799 (N_7799,N_6073,N_5288);
and U7800 (N_7800,N_3316,N_1866);
xnor U7801 (N_7801,N_4482,N_3202);
or U7802 (N_7802,N_167,N_144);
xor U7803 (N_7803,N_3260,N_1763);
and U7804 (N_7804,N_2366,N_602);
and U7805 (N_7805,N_5910,N_2339);
or U7806 (N_7806,N_5715,N_4610);
or U7807 (N_7807,N_5721,N_3196);
xor U7808 (N_7808,N_6074,N_5151);
or U7809 (N_7809,N_6111,N_222);
or U7810 (N_7810,N_1593,N_2907);
nor U7811 (N_7811,N_1904,N_4140);
xor U7812 (N_7812,N_1768,N_4116);
nand U7813 (N_7813,N_4709,N_2866);
nor U7814 (N_7814,N_5486,N_3042);
xnor U7815 (N_7815,N_1664,N_2433);
nor U7816 (N_7816,N_805,N_840);
nand U7817 (N_7817,N_3249,N_4781);
nor U7818 (N_7818,N_1380,N_3675);
nand U7819 (N_7819,N_5011,N_2648);
and U7820 (N_7820,N_2432,N_3869);
nand U7821 (N_7821,N_4155,N_4106);
or U7822 (N_7822,N_455,N_323);
xnor U7823 (N_7823,N_4774,N_1383);
xnor U7824 (N_7824,N_4769,N_3760);
xnor U7825 (N_7825,N_3607,N_1868);
xnor U7826 (N_7826,N_1961,N_6001);
nand U7827 (N_7827,N_448,N_189);
or U7828 (N_7828,N_1339,N_2713);
nand U7829 (N_7829,N_1729,N_3824);
and U7830 (N_7830,N_4420,N_3164);
xnor U7831 (N_7831,N_58,N_4758);
xor U7832 (N_7832,N_1772,N_420);
nor U7833 (N_7833,N_3838,N_622);
xor U7834 (N_7834,N_396,N_4295);
and U7835 (N_7835,N_1785,N_1374);
or U7836 (N_7836,N_1986,N_3513);
or U7837 (N_7837,N_1997,N_3180);
or U7838 (N_7838,N_6107,N_2445);
and U7839 (N_7839,N_1467,N_5918);
nand U7840 (N_7840,N_4224,N_1592);
or U7841 (N_7841,N_5222,N_5706);
or U7842 (N_7842,N_1002,N_5591);
and U7843 (N_7843,N_5287,N_3074);
nand U7844 (N_7844,N_207,N_412);
or U7845 (N_7845,N_3235,N_5349);
or U7846 (N_7846,N_3407,N_3562);
nand U7847 (N_7847,N_5476,N_4498);
xnor U7848 (N_7848,N_4292,N_882);
nand U7849 (N_7849,N_5040,N_3313);
or U7850 (N_7850,N_1967,N_6041);
nand U7851 (N_7851,N_1701,N_1792);
xor U7852 (N_7852,N_4460,N_668);
and U7853 (N_7853,N_1375,N_4953);
nand U7854 (N_7854,N_3076,N_271);
or U7855 (N_7855,N_3603,N_188);
nor U7856 (N_7856,N_4100,N_5121);
or U7857 (N_7857,N_2631,N_6158);
or U7858 (N_7858,N_4404,N_4223);
and U7859 (N_7859,N_4421,N_1354);
or U7860 (N_7860,N_3818,N_4464);
or U7861 (N_7861,N_5460,N_1090);
nand U7862 (N_7862,N_3777,N_4692);
and U7863 (N_7863,N_1970,N_5839);
or U7864 (N_7864,N_5869,N_6124);
xnor U7865 (N_7865,N_3860,N_5015);
nand U7866 (N_7866,N_5277,N_2329);
or U7867 (N_7867,N_166,N_402);
xor U7868 (N_7868,N_4521,N_3650);
and U7869 (N_7869,N_3705,N_3616);
nor U7870 (N_7870,N_2929,N_419);
xor U7871 (N_7871,N_5297,N_5724);
nor U7872 (N_7872,N_4740,N_2620);
nand U7873 (N_7873,N_2100,N_5867);
xnor U7874 (N_7874,N_5267,N_2536);
nand U7875 (N_7875,N_3794,N_2495);
xor U7876 (N_7876,N_735,N_3647);
nand U7877 (N_7877,N_3667,N_5835);
xnor U7878 (N_7878,N_2383,N_4477);
xnor U7879 (N_7879,N_2715,N_3813);
nor U7880 (N_7880,N_1195,N_5935);
and U7881 (N_7881,N_1550,N_109);
or U7882 (N_7882,N_4448,N_630);
xor U7883 (N_7883,N_6011,N_4662);
or U7884 (N_7884,N_4211,N_1056);
xnor U7885 (N_7885,N_2908,N_5212);
xnor U7886 (N_7886,N_5815,N_6237);
or U7887 (N_7887,N_5294,N_3811);
and U7888 (N_7888,N_1013,N_5326);
nor U7889 (N_7889,N_1487,N_3282);
nand U7890 (N_7890,N_5137,N_939);
nor U7891 (N_7891,N_5698,N_5166);
xnor U7892 (N_7892,N_5133,N_3596);
or U7893 (N_7893,N_2080,N_3099);
or U7894 (N_7894,N_101,N_3417);
nor U7895 (N_7895,N_1209,N_2333);
and U7896 (N_7896,N_5555,N_4323);
or U7897 (N_7897,N_5170,N_4850);
or U7898 (N_7898,N_5275,N_5293);
xnor U7899 (N_7899,N_3662,N_4331);
nor U7900 (N_7900,N_5118,N_3166);
and U7901 (N_7901,N_5245,N_3448);
xor U7902 (N_7902,N_2676,N_2599);
or U7903 (N_7903,N_371,N_421);
nor U7904 (N_7904,N_4456,N_1166);
xnor U7905 (N_7905,N_4923,N_2171);
nand U7906 (N_7906,N_996,N_3769);
nand U7907 (N_7907,N_1060,N_4013);
nor U7908 (N_7908,N_5233,N_4829);
xnor U7909 (N_7909,N_3909,N_1848);
xnor U7910 (N_7910,N_2154,N_5123);
nor U7911 (N_7911,N_1407,N_235);
nand U7912 (N_7912,N_4897,N_2677);
and U7913 (N_7913,N_1988,N_3161);
or U7914 (N_7914,N_1210,N_605);
nand U7915 (N_7915,N_1438,N_4921);
xor U7916 (N_7916,N_6141,N_2310);
or U7917 (N_7917,N_614,N_2684);
nor U7918 (N_7918,N_5370,N_4699);
nand U7919 (N_7919,N_119,N_3474);
nand U7920 (N_7920,N_2068,N_3247);
xor U7921 (N_7921,N_4559,N_6049);
nand U7922 (N_7922,N_4129,N_4457);
xnor U7923 (N_7923,N_441,N_2337);
nand U7924 (N_7924,N_4653,N_982);
and U7925 (N_7925,N_1803,N_295);
xor U7926 (N_7926,N_4838,N_5538);
or U7927 (N_7927,N_1388,N_853);
nor U7928 (N_7928,N_2262,N_1648);
and U7929 (N_7929,N_4724,N_426);
nand U7930 (N_7930,N_5563,N_5382);
nor U7931 (N_7931,N_2865,N_4125);
or U7932 (N_7932,N_3764,N_3536);
nor U7933 (N_7933,N_5825,N_6188);
and U7934 (N_7934,N_1517,N_2395);
or U7935 (N_7935,N_1478,N_6245);
nor U7936 (N_7936,N_3591,N_2483);
and U7937 (N_7937,N_2209,N_5157);
nor U7938 (N_7938,N_3563,N_2750);
nor U7939 (N_7939,N_5528,N_714);
nor U7940 (N_7940,N_4964,N_5949);
nor U7941 (N_7941,N_3800,N_1325);
nand U7942 (N_7942,N_3371,N_0);
xor U7943 (N_7943,N_4958,N_4515);
or U7944 (N_7944,N_1424,N_5390);
and U7945 (N_7945,N_1590,N_3503);
nor U7946 (N_7946,N_1780,N_4936);
and U7947 (N_7947,N_2652,N_3726);
and U7948 (N_7948,N_1797,N_3733);
nand U7949 (N_7949,N_3061,N_2774);
nand U7950 (N_7950,N_3765,N_5761);
and U7951 (N_7951,N_3265,N_2258);
nand U7952 (N_7952,N_5914,N_2031);
nor U7953 (N_7953,N_3560,N_5314);
xnor U7954 (N_7954,N_3081,N_601);
xor U7955 (N_7955,N_5716,N_5091);
or U7956 (N_7956,N_2822,N_257);
nor U7957 (N_7957,N_1510,N_3712);
and U7958 (N_7958,N_1148,N_2744);
and U7959 (N_7959,N_2979,N_3308);
nand U7960 (N_7960,N_4884,N_916);
xnor U7961 (N_7961,N_3185,N_198);
xor U7962 (N_7962,N_3699,N_3035);
xor U7963 (N_7963,N_4422,N_3203);
or U7964 (N_7964,N_666,N_5433);
or U7965 (N_7965,N_4646,N_1320);
or U7966 (N_7966,N_1349,N_2696);
or U7967 (N_7967,N_2519,N_3148);
and U7968 (N_7968,N_4442,N_550);
nand U7969 (N_7969,N_1827,N_5414);
nor U7970 (N_7970,N_1975,N_2012);
xor U7971 (N_7971,N_4599,N_2428);
nand U7972 (N_7972,N_3519,N_5331);
nor U7973 (N_7973,N_491,N_5017);
nand U7974 (N_7974,N_4310,N_1632);
or U7975 (N_7975,N_5699,N_5167);
nor U7976 (N_7976,N_5419,N_2662);
and U7977 (N_7977,N_3888,N_3241);
nand U7978 (N_7978,N_2626,N_2070);
or U7979 (N_7979,N_2272,N_3550);
nand U7980 (N_7980,N_964,N_892);
nand U7981 (N_7981,N_3828,N_4452);
and U7982 (N_7982,N_3534,N_1972);
xnor U7983 (N_7983,N_4234,N_5550);
xnor U7984 (N_7984,N_513,N_1200);
xnor U7985 (N_7985,N_595,N_2422);
or U7986 (N_7986,N_2960,N_2897);
or U7987 (N_7987,N_298,N_2893);
nor U7988 (N_7988,N_3152,N_1651);
and U7989 (N_7989,N_2405,N_589);
or U7990 (N_7990,N_1043,N_204);
nand U7991 (N_7991,N_4424,N_4714);
xnor U7992 (N_7992,N_2763,N_1169);
or U7993 (N_7993,N_1418,N_415);
or U7994 (N_7994,N_937,N_1943);
xnor U7995 (N_7995,N_6119,N_4965);
xnor U7996 (N_7996,N_1030,N_5920);
and U7997 (N_7997,N_1258,N_4243);
xor U7998 (N_7998,N_603,N_5229);
nand U7999 (N_7999,N_4658,N_4626);
or U8000 (N_8000,N_1734,N_4843);
or U8001 (N_8001,N_774,N_1824);
or U8002 (N_8002,N_3704,N_3136);
xor U8003 (N_8003,N_5529,N_2412);
or U8004 (N_8004,N_6080,N_3941);
nand U8005 (N_8005,N_1699,N_2999);
nor U8006 (N_8006,N_6040,N_3858);
and U8007 (N_8007,N_5524,N_483);
or U8008 (N_8008,N_874,N_6007);
nand U8009 (N_8009,N_1413,N_4332);
nor U8010 (N_8010,N_465,N_5286);
nor U8011 (N_8011,N_2912,N_4425);
and U8012 (N_8012,N_1014,N_1131);
nor U8013 (N_8013,N_255,N_1473);
xor U8014 (N_8014,N_993,N_1317);
nand U8015 (N_8015,N_4208,N_2285);
nand U8016 (N_8016,N_1655,N_2471);
and U8017 (N_8017,N_1097,N_3846);
xnor U8018 (N_8018,N_5644,N_5853);
xor U8019 (N_8019,N_983,N_5987);
xnor U8020 (N_8020,N_2124,N_3302);
nand U8021 (N_8021,N_5745,N_1395);
and U8022 (N_8022,N_3611,N_3931);
xnor U8023 (N_8023,N_5075,N_5976);
or U8024 (N_8024,N_2398,N_322);
xor U8025 (N_8025,N_3158,N_2157);
xnor U8026 (N_8026,N_936,N_583);
and U8027 (N_8027,N_2561,N_3217);
xnor U8028 (N_8028,N_2708,N_2741);
xnor U8029 (N_8029,N_435,N_3085);
nand U8030 (N_8030,N_3327,N_3795);
or U8031 (N_8031,N_3512,N_72);
xnor U8032 (N_8032,N_5904,N_1663);
and U8033 (N_8033,N_172,N_2453);
nand U8034 (N_8034,N_1963,N_762);
nor U8035 (N_8035,N_5407,N_3362);
and U8036 (N_8036,N_1811,N_5870);
and U8037 (N_8037,N_5362,N_6083);
nor U8038 (N_8038,N_5408,N_4759);
xnor U8039 (N_8039,N_5794,N_3573);
nor U8040 (N_8040,N_4071,N_5993);
nor U8041 (N_8041,N_2575,N_366);
nand U8042 (N_8042,N_4089,N_4122);
nor U8043 (N_8043,N_851,N_4345);
and U8044 (N_8044,N_4787,N_2032);
nor U8045 (N_8045,N_5213,N_5429);
nor U8046 (N_8046,N_1927,N_5425);
and U8047 (N_8047,N_74,N_3925);
xor U8048 (N_8048,N_4907,N_2553);
nand U8049 (N_8049,N_2423,N_156);
xor U8050 (N_8050,N_2875,N_5069);
nand U8051 (N_8051,N_1885,N_2001);
and U8052 (N_8052,N_4465,N_2691);
or U8053 (N_8053,N_1269,N_2095);
or U8054 (N_8054,N_1481,N_1093);
or U8055 (N_8055,N_5974,N_3018);
nand U8056 (N_8056,N_2852,N_5254);
xnor U8057 (N_8057,N_3664,N_3068);
or U8058 (N_8058,N_6085,N_3014);
xor U8059 (N_8059,N_5312,N_4255);
or U8060 (N_8060,N_6042,N_4632);
xor U8061 (N_8061,N_3261,N_3115);
or U8062 (N_8062,N_885,N_5223);
nor U8063 (N_8063,N_5672,N_309);
nor U8064 (N_8064,N_1255,N_1028);
nor U8065 (N_8065,N_4337,N_2703);
xnor U8066 (N_8066,N_4373,N_2219);
nand U8067 (N_8067,N_2663,N_2358);
nand U8068 (N_8068,N_1029,N_3635);
or U8069 (N_8069,N_2722,N_4888);
nor U8070 (N_8070,N_4849,N_3280);
nand U8071 (N_8071,N_3012,N_2403);
or U8072 (N_8072,N_4489,N_2578);
xnor U8073 (N_8073,N_1422,N_5994);
nand U8074 (N_8074,N_1136,N_1884);
xnor U8075 (N_8075,N_3420,N_3510);
or U8076 (N_8076,N_5298,N_2539);
or U8077 (N_8077,N_4526,N_1678);
and U8078 (N_8078,N_3677,N_6233);
or U8079 (N_8079,N_651,N_3899);
xnor U8080 (N_8080,N_2697,N_1671);
nand U8081 (N_8081,N_4989,N_4128);
and U8082 (N_8082,N_1683,N_5208);
nor U8083 (N_8083,N_1677,N_1715);
and U8084 (N_8084,N_5919,N_1774);
and U8085 (N_8085,N_4800,N_2010);
nor U8086 (N_8086,N_5778,N_825);
nand U8087 (N_8087,N_6143,N_1916);
and U8088 (N_8088,N_3579,N_4556);
and U8089 (N_8089,N_3722,N_705);
xnor U8090 (N_8090,N_4974,N_849);
nand U8091 (N_8091,N_5570,N_1020);
and U8092 (N_8092,N_3001,N_5569);
xor U8093 (N_8093,N_2809,N_5308);
and U8094 (N_8094,N_5651,N_4757);
or U8095 (N_8095,N_1585,N_1851);
or U8096 (N_8096,N_2323,N_562);
xnor U8097 (N_8097,N_6240,N_5007);
or U8098 (N_8098,N_1048,N_4725);
nor U8099 (N_8099,N_1322,N_2204);
nand U8100 (N_8100,N_4051,N_4440);
or U8101 (N_8101,N_6101,N_3343);
or U8102 (N_8102,N_772,N_3147);
nor U8103 (N_8103,N_302,N_5172);
xor U8104 (N_8104,N_5633,N_1554);
nor U8105 (N_8105,N_5334,N_3238);
nor U8106 (N_8106,N_388,N_2078);
or U8107 (N_8107,N_1128,N_1396);
nor U8108 (N_8108,N_299,N_2347);
nor U8109 (N_8109,N_4602,N_1752);
and U8110 (N_8110,N_745,N_585);
nor U8111 (N_8111,N_5705,N_5634);
or U8112 (N_8112,N_1602,N_4731);
nor U8113 (N_8113,N_1099,N_5176);
nor U8114 (N_8114,N_1644,N_5393);
nor U8115 (N_8115,N_1557,N_286);
and U8116 (N_8116,N_5330,N_2245);
and U8117 (N_8117,N_4682,N_5036);
and U8118 (N_8118,N_5612,N_1834);
nand U8119 (N_8119,N_4186,N_3859);
nor U8120 (N_8120,N_3175,N_940);
nand U8121 (N_8121,N_3418,N_1044);
and U8122 (N_8122,N_3419,N_1790);
or U8123 (N_8123,N_5683,N_1930);
xnor U8124 (N_8124,N_3868,N_2554);
or U8125 (N_8125,N_3393,N_3653);
nor U8126 (N_8126,N_2558,N_1984);
nand U8127 (N_8127,N_296,N_1802);
nor U8128 (N_8128,N_4862,N_5615);
nand U8129 (N_8129,N_1189,N_2861);
xnor U8130 (N_8130,N_3463,N_4881);
nand U8131 (N_8131,N_506,N_6239);
nor U8132 (N_8132,N_3290,N_5913);
nor U8133 (N_8133,N_3447,N_4788);
and U8134 (N_8134,N_5783,N_1108);
and U8135 (N_8135,N_5210,N_3556);
xor U8136 (N_8136,N_841,N_5912);
and U8137 (N_8137,N_1945,N_2169);
nor U8138 (N_8138,N_975,N_5625);
xor U8139 (N_8139,N_949,N_14);
or U8140 (N_8140,N_2253,N_4076);
nand U8141 (N_8141,N_4831,N_5660);
nor U8142 (N_8142,N_4446,N_3025);
and U8143 (N_8143,N_5649,N_2267);
xnor U8144 (N_8144,N_5723,N_797);
nand U8145 (N_8145,N_57,N_5693);
nor U8146 (N_8146,N_3179,N_2384);
xor U8147 (N_8147,N_485,N_4748);
and U8148 (N_8148,N_4103,N_239);
and U8149 (N_8149,N_5726,N_736);
nand U8150 (N_8150,N_4055,N_3696);
xnor U8151 (N_8151,N_977,N_3731);
xnor U8152 (N_8152,N_2766,N_3629);
xor U8153 (N_8153,N_6057,N_3172);
nor U8154 (N_8154,N_1645,N_115);
xnor U8155 (N_8155,N_941,N_1569);
or U8156 (N_8156,N_4929,N_4846);
or U8157 (N_8157,N_6014,N_1810);
nand U8158 (N_8158,N_5001,N_5502);
nor U8159 (N_8159,N_1068,N_5317);
nand U8160 (N_8160,N_2540,N_5237);
nand U8161 (N_8161,N_4198,N_89);
xor U8162 (N_8162,N_2281,N_5991);
and U8163 (N_8163,N_5410,N_934);
xnor U8164 (N_8164,N_6039,N_6016);
nor U8165 (N_8165,N_2136,N_1115);
xnor U8166 (N_8166,N_2564,N_2344);
and U8167 (N_8167,N_409,N_1337);
nor U8168 (N_8168,N_5696,N_1628);
nor U8169 (N_8169,N_300,N_4564);
nand U8170 (N_8170,N_5571,N_3879);
xnor U8171 (N_8171,N_3996,N_3110);
nor U8172 (N_8172,N_3528,N_2099);
nor U8173 (N_8173,N_1420,N_6094);
nand U8174 (N_8174,N_60,N_3621);
nand U8175 (N_8175,N_5152,N_3130);
and U8176 (N_8176,N_3472,N_4004);
or U8177 (N_8177,N_4227,N_489);
nor U8178 (N_8178,N_132,N_2086);
nand U8179 (N_8179,N_1078,N_3444);
xnor U8180 (N_8180,N_1949,N_3465);
nand U8181 (N_8181,N_3462,N_618);
or U8182 (N_8182,N_3262,N_3636);
nand U8183 (N_8183,N_6054,N_2759);
nor U8184 (N_8184,N_3649,N_4927);
nor U8185 (N_8185,N_2201,N_3875);
or U8186 (N_8186,N_5631,N_1301);
xor U8187 (N_8187,N_908,N_1486);
nand U8188 (N_8188,N_2930,N_6093);
nand U8189 (N_8189,N_3063,N_3866);
or U8190 (N_8190,N_3258,N_3160);
xnor U8191 (N_8191,N_1825,N_1668);
nand U8192 (N_8192,N_1459,N_2050);
xor U8193 (N_8193,N_1083,N_1522);
or U8194 (N_8194,N_1747,N_2647);
xnor U8195 (N_8195,N_1591,N_3045);
nand U8196 (N_8196,N_1071,N_2287);
nor U8197 (N_8197,N_5526,N_4806);
nor U8198 (N_8198,N_5327,N_5492);
nand U8199 (N_8199,N_3832,N_5392);
xnor U8200 (N_8200,N_783,N_947);
nand U8201 (N_8201,N_2522,N_2524);
nand U8202 (N_8202,N_4235,N_6150);
xnor U8203 (N_8203,N_3000,N_1141);
xor U8204 (N_8204,N_5939,N_5964);
xor U8205 (N_8205,N_1531,N_2570);
nand U8206 (N_8206,N_1643,N_2401);
xor U8207 (N_8207,N_5196,N_184);
xor U8208 (N_8208,N_1756,N_3067);
nor U8209 (N_8209,N_5350,N_405);
and U8210 (N_8210,N_4734,N_2791);
and U8211 (N_8211,N_1749,N_1474);
nor U8212 (N_8212,N_1782,N_356);
nand U8213 (N_8213,N_2102,N_4747);
nor U8214 (N_8214,N_3255,N_505);
xor U8215 (N_8215,N_1836,N_3244);
or U8216 (N_8216,N_2443,N_4647);
or U8217 (N_8217,N_2321,N_2484);
nor U8218 (N_8218,N_4611,N_3583);
or U8219 (N_8219,N_2015,N_2148);
nor U8220 (N_8220,N_3759,N_5965);
nand U8221 (N_8221,N_1794,N_66);
nand U8222 (N_8222,N_1134,N_3028);
and U8223 (N_8223,N_3505,N_2669);
xor U8224 (N_8224,N_5388,N_2437);
or U8225 (N_8225,N_5336,N_3938);
nor U8226 (N_8226,N_4022,N_2480);
nand U8227 (N_8227,N_2223,N_1730);
xnor U8228 (N_8228,N_3542,N_1887);
nand U8229 (N_8229,N_4185,N_2349);
and U8230 (N_8230,N_1246,N_5814);
xor U8231 (N_8231,N_5467,N_530);
nor U8232 (N_8232,N_5406,N_5539);
xnor U8233 (N_8233,N_1082,N_1207);
nand U8234 (N_8234,N_778,N_1274);
nand U8235 (N_8235,N_2686,N_3673);
and U8236 (N_8236,N_763,N_4984);
nand U8237 (N_8237,N_3833,N_926);
xor U8238 (N_8238,N_2970,N_2905);
and U8239 (N_8239,N_1404,N_2859);
and U8240 (N_8240,N_2574,N_3952);
and U8241 (N_8241,N_392,N_5466);
and U8242 (N_8242,N_3515,N_4126);
nand U8243 (N_8243,N_5760,N_4563);
or U8244 (N_8244,N_3545,N_686);
xnor U8245 (N_8245,N_895,N_2028);
xnor U8246 (N_8246,N_4207,N_2545);
nor U8247 (N_8247,N_556,N_3628);
or U8248 (N_8248,N_5973,N_3753);
xnor U8249 (N_8249,N_4665,N_5789);
nand U8250 (N_8250,N_522,N_3008);
nand U8251 (N_8251,N_468,N_3376);
xor U8252 (N_8252,N_3157,N_5066);
or U8253 (N_8253,N_1845,N_343);
nand U8254 (N_8254,N_5367,N_1057);
nor U8255 (N_8255,N_4029,N_231);
or U8256 (N_8256,N_3083,N_5903);
and U8257 (N_8257,N_6047,N_2273);
nand U8258 (N_8258,N_4005,N_2706);
xor U8259 (N_8259,N_4258,N_6227);
or U8260 (N_8260,N_1928,N_6244);
or U8261 (N_8261,N_691,N_1770);
nand U8262 (N_8262,N_3780,N_3358);
and U8263 (N_8263,N_5580,N_2518);
xnor U8264 (N_8264,N_117,N_4135);
or U8265 (N_8265,N_4728,N_2069);
or U8266 (N_8266,N_1431,N_1597);
nor U8267 (N_8267,N_6034,N_5042);
xor U8268 (N_8268,N_1295,N_3600);
or U8269 (N_8269,N_5799,N_4870);
xor U8270 (N_8270,N_1709,N_4585);
xor U8271 (N_8271,N_4069,N_5424);
and U8272 (N_8272,N_3112,N_3020);
and U8273 (N_8273,N_5898,N_5062);
nor U8274 (N_8274,N_3584,N_846);
xor U8275 (N_8275,N_5807,N_5488);
nand U8276 (N_8276,N_2035,N_4197);
and U8277 (N_8277,N_3479,N_2700);
or U8278 (N_8278,N_3484,N_6053);
nor U8279 (N_8279,N_913,N_1842);
nand U8280 (N_8280,N_796,N_1281);
or U8281 (N_8281,N_3963,N_4131);
xor U8282 (N_8282,N_2470,N_1436);
or U8283 (N_8283,N_2651,N_78);
or U8284 (N_8284,N_3725,N_903);
or U8285 (N_8285,N_5074,N_381);
nor U8286 (N_8286,N_3269,N_5709);
nand U8287 (N_8287,N_5596,N_4439);
nor U8288 (N_8288,N_4689,N_2666);
nand U8289 (N_8289,N_358,N_4909);
or U8290 (N_8290,N_1179,N_4847);
nand U8291 (N_8291,N_894,N_5498);
xor U8292 (N_8292,N_4691,N_2789);
nand U8293 (N_8293,N_4133,N_3455);
xnor U8294 (N_8294,N_261,N_1880);
nor U8295 (N_8295,N_357,N_2118);
nand U8296 (N_8296,N_5181,N_3982);
nand U8297 (N_8297,N_4177,N_2450);
nor U8298 (N_8298,N_5217,N_883);
and U8299 (N_8299,N_5027,N_1019);
nand U8300 (N_8300,N_1580,N_2311);
nand U8301 (N_8301,N_1861,N_2913);
nand U8302 (N_8302,N_2256,N_4389);
or U8303 (N_8303,N_3186,N_1253);
and U8304 (N_8304,N_168,N_4525);
or U8305 (N_8305,N_612,N_5458);
xor U8306 (N_8306,N_1857,N_3033);
xnor U8307 (N_8307,N_61,N_2164);
and U8308 (N_8308,N_1208,N_2003);
nand U8309 (N_8309,N_4752,N_1291);
xor U8310 (N_8310,N_3737,N_2776);
and U8311 (N_8311,N_2943,N_1266);
nand U8312 (N_8312,N_1457,N_5841);
xnor U8313 (N_8313,N_312,N_2404);
or U8314 (N_8314,N_4959,N_1516);
xnor U8315 (N_8315,N_2502,N_3902);
nand U8316 (N_8316,N_347,N_1261);
and U8317 (N_8317,N_4765,N_4686);
nor U8318 (N_8318,N_3533,N_6105);
nand U8319 (N_8319,N_1217,N_3120);
and U8320 (N_8320,N_4325,N_4950);
or U8321 (N_8321,N_5513,N_1027);
or U8322 (N_8322,N_2736,N_236);
nor U8323 (N_8323,N_1283,N_4327);
xnor U8324 (N_8324,N_3798,N_4770);
xnor U8325 (N_8325,N_582,N_1331);
and U8326 (N_8326,N_6177,N_5436);
or U8327 (N_8327,N_4390,N_952);
nor U8328 (N_8328,N_1805,N_3317);
and U8329 (N_8329,N_2350,N_1833);
nor U8330 (N_8330,N_1103,N_2772);
and U8331 (N_8331,N_1571,N_5218);
nand U8332 (N_8332,N_3095,N_4887);
nor U8333 (N_8333,N_1865,N_6015);
nand U8334 (N_8334,N_1979,N_2504);
nor U8335 (N_8335,N_227,N_1559);
nor U8336 (N_8336,N_1171,N_1305);
xor U8337 (N_8337,N_5054,N_4630);
xnor U8338 (N_8338,N_3823,N_4301);
nor U8339 (N_8339,N_4628,N_5205);
nor U8340 (N_8340,N_3059,N_717);
nor U8341 (N_8341,N_854,N_2284);
nor U8342 (N_8342,N_4275,N_259);
xnor U8343 (N_8343,N_5415,N_4916);
xnor U8344 (N_8344,N_4982,N_4320);
nand U8345 (N_8345,N_3654,N_2167);
or U8346 (N_8346,N_3491,N_5717);
or U8347 (N_8347,N_5646,N_4866);
nor U8348 (N_8348,N_1552,N_2853);
nor U8349 (N_8349,N_3043,N_3109);
and U8350 (N_8350,N_5924,N_4889);
nor U8351 (N_8351,N_3286,N_787);
and U8352 (N_8352,N_4283,N_689);
nand U8353 (N_8353,N_1621,N_470);
or U8354 (N_8354,N_2222,N_791);
and U8355 (N_8355,N_3847,N_1088);
or U8356 (N_8356,N_5661,N_5980);
or U8357 (N_8357,N_5562,N_2113);
nor U8358 (N_8358,N_4027,N_4518);
and U8359 (N_8359,N_1598,N_2234);
nor U8360 (N_8360,N_2972,N_2490);
nand U8361 (N_8361,N_203,N_141);
nand U8362 (N_8362,N_2925,N_4153);
or U8363 (N_8363,N_3240,N_3292);
and U8364 (N_8364,N_3254,N_120);
nand U8365 (N_8365,N_776,N_3415);
nand U8366 (N_8366,N_5713,N_3691);
nor U8367 (N_8367,N_2896,N_4230);
nor U8368 (N_8368,N_2505,N_1241);
nor U8369 (N_8369,N_282,N_1959);
or U8370 (N_8370,N_5942,N_5953);
nand U8371 (N_8371,N_321,N_3009);
nand U8372 (N_8372,N_162,N_4749);
and U8373 (N_8373,N_4472,N_5752);
and U8374 (N_8374,N_5574,N_2417);
nand U8375 (N_8375,N_3724,N_4878);
or U8376 (N_8376,N_4259,N_5708);
nand U8377 (N_8377,N_2425,N_1727);
or U8378 (N_8378,N_2692,N_2468);
nor U8379 (N_8379,N_5940,N_4311);
nand U8380 (N_8380,N_3913,N_6199);
nand U8381 (N_8381,N_2277,N_329);
nand U8382 (N_8382,N_67,N_2964);
and U8383 (N_8383,N_467,N_2135);
or U8384 (N_8384,N_3251,N_2279);
nor U8385 (N_8385,N_3438,N_859);
and U8386 (N_8386,N_2379,N_5160);
or U8387 (N_8387,N_2026,N_4938);
nand U8388 (N_8388,N_6144,N_5507);
nand U8389 (N_8389,N_3127,N_5831);
nor U8390 (N_8390,N_2612,N_2197);
xor U8391 (N_8391,N_609,N_1947);
nor U8392 (N_8392,N_4524,N_4523);
xor U8393 (N_8393,N_1211,N_6152);
or U8394 (N_8394,N_3819,N_2577);
xnor U8395 (N_8395,N_3631,N_3264);
nand U8396 (N_8396,N_4531,N_2177);
and U8397 (N_8397,N_587,N_1686);
xor U8398 (N_8398,N_1163,N_5868);
nor U8399 (N_8399,N_3618,N_2299);
nor U8400 (N_8400,N_4633,N_3884);
nand U8401 (N_8401,N_1393,N_2133);
nand U8402 (N_8402,N_1377,N_5845);
nand U8403 (N_8403,N_2147,N_4094);
xnor U8404 (N_8404,N_1765,N_6086);
or U8405 (N_8405,N_3867,N_2783);
nand U8406 (N_8406,N_3293,N_2770);
or U8407 (N_8407,N_4409,N_4043);
nand U8408 (N_8408,N_5732,N_4138);
and U8409 (N_8409,N_743,N_3882);
xor U8410 (N_8410,N_3610,N_4031);
and U8411 (N_8411,N_1193,N_4943);
and U8412 (N_8412,N_5906,N_2090);
xor U8413 (N_8413,N_1992,N_5930);
and U8414 (N_8414,N_2727,N_2637);
or U8415 (N_8415,N_3174,N_6238);
xnor U8416 (N_8416,N_4744,N_644);
and U8417 (N_8417,N_3954,N_3700);
or U8418 (N_8418,N_2413,N_341);
nor U8419 (N_8419,N_4260,N_2813);
xnor U8420 (N_8420,N_2712,N_2457);
or U8421 (N_8421,N_5464,N_3520);
or U8422 (N_8422,N_3714,N_2891);
nor U8423 (N_8423,N_1506,N_3693);
nand U8424 (N_8424,N_5934,N_1035);
or U8425 (N_8425,N_1310,N_3684);
nor U8426 (N_8426,N_5534,N_5238);
nand U8427 (N_8427,N_3242,N_5629);
nor U8428 (N_8428,N_5522,N_538);
nand U8429 (N_8429,N_3792,N_3131);
xnor U8430 (N_8430,N_3885,N_4977);
and U8431 (N_8431,N_4663,N_4152);
nand U8432 (N_8432,N_2785,N_6165);
xnor U8433 (N_8433,N_5772,N_2206);
xnor U8434 (N_8434,N_5461,N_3502);
or U8435 (N_8435,N_2755,N_2046);
and U8436 (N_8436,N_5295,N_1318);
nand U8437 (N_8437,N_4819,N_3529);
nor U8438 (N_8438,N_4513,N_3168);
nand U8439 (N_8439,N_461,N_5821);
and U8440 (N_8440,N_1194,N_2477);
nor U8441 (N_8441,N_149,N_5655);
and U8442 (N_8442,N_1069,N_3493);
nor U8443 (N_8443,N_3713,N_9);
nor U8444 (N_8444,N_1373,N_568);
xor U8445 (N_8445,N_2593,N_2562);
xor U8446 (N_8446,N_5085,N_2332);
xor U8447 (N_8447,N_662,N_1086);
nand U8448 (N_8448,N_4891,N_2671);
xor U8449 (N_8449,N_5194,N_3088);
and U8450 (N_8450,N_2753,N_2129);
nor U8451 (N_8451,N_3430,N_500);
or U8452 (N_8452,N_4417,N_3715);
or U8453 (N_8453,N_1182,N_209);
and U8454 (N_8454,N_397,N_4998);
or U8455 (N_8455,N_5781,N_2241);
and U8456 (N_8456,N_921,N_1714);
xor U8457 (N_8457,N_624,N_5886);
nor U8458 (N_8458,N_4597,N_3332);
nor U8459 (N_8459,N_970,N_1893);
or U8460 (N_8460,N_5786,N_3471);
or U8461 (N_8461,N_2389,N_2724);
xnor U8462 (N_8462,N_1561,N_3038);
or U8463 (N_8463,N_1125,N_4536);
nor U8464 (N_8464,N_3680,N_3771);
or U8465 (N_8465,N_2251,N_5291);
and U8466 (N_8466,N_4496,N_2725);
nand U8467 (N_8467,N_6161,N_1630);
or U8468 (N_8468,N_3272,N_5077);
or U8469 (N_8469,N_577,N_842);
nand U8470 (N_8470,N_1280,N_3222);
nor U8471 (N_8471,N_5975,N_3369);
and U8472 (N_8472,N_5420,N_2542);
nor U8473 (N_8473,N_4137,N_3643);
or U8474 (N_8474,N_5589,N_5895);
nand U8475 (N_8475,N_3752,N_4001);
nor U8476 (N_8476,N_3564,N_263);
xnor U8477 (N_8477,N_5936,N_2576);
and U8478 (N_8478,N_3481,N_2968);
nand U8479 (N_8479,N_1220,N_3507);
and U8480 (N_8480,N_307,N_2264);
xnor U8481 (N_8481,N_4370,N_6096);
nor U8482 (N_8482,N_5480,N_1448);
xor U8483 (N_8483,N_767,N_2618);
or U8484 (N_8484,N_726,N_5657);
nor U8485 (N_8485,N_3671,N_3644);
and U8486 (N_8486,N_1479,N_2391);
xnor U8487 (N_8487,N_3877,N_1526);
nor U8488 (N_8488,N_3246,N_2901);
xnor U8489 (N_8489,N_1858,N_1462);
and U8490 (N_8490,N_1993,N_645);
or U8491 (N_8491,N_2898,N_6175);
xnor U8492 (N_8492,N_697,N_3382);
and U8493 (N_8493,N_1633,N_580);
and U8494 (N_8494,N_3589,N_2276);
and U8495 (N_8495,N_3201,N_3356);
and U8496 (N_8496,N_3423,N_2957);
or U8497 (N_8497,N_2071,N_6012);
and U8498 (N_8498,N_4309,N_2486);
nor U8499 (N_8499,N_1843,N_2510);
nand U8500 (N_8500,N_5159,N_4670);
or U8501 (N_8501,N_2679,N_5230);
and U8502 (N_8502,N_1541,N_5754);
nor U8503 (N_8503,N_2215,N_326);
nor U8504 (N_8504,N_5862,N_2600);
nand U8505 (N_8505,N_1784,N_1728);
and U8506 (N_8506,N_4038,N_1408);
nor U8507 (N_8507,N_5012,N_5971);
and U8508 (N_8508,N_3857,N_4132);
or U8509 (N_8509,N_638,N_4635);
xor U8510 (N_8510,N_3036,N_758);
nand U8511 (N_8511,N_923,N_4562);
nor U8512 (N_8512,N_4028,N_3852);
nand U8513 (N_8513,N_5068,N_876);
nor U8514 (N_8514,N_1798,N_1445);
and U8515 (N_8515,N_1361,N_1023);
or U8516 (N_8516,N_3287,N_3449);
xor U8517 (N_8517,N_3497,N_759);
xor U8518 (N_8518,N_1710,N_984);
and U8519 (N_8519,N_5090,N_5747);
or U8520 (N_8520,N_2832,N_3915);
nand U8521 (N_8521,N_2182,N_4902);
xor U8522 (N_8522,N_3655,N_508);
nor U8523 (N_8523,N_5665,N_4987);
or U8524 (N_8524,N_1228,N_5117);
xor U8525 (N_8525,N_6066,N_1472);
and U8526 (N_8526,N_971,N_858);
nand U8527 (N_8527,N_6183,N_1326);
nor U8528 (N_8528,N_3808,N_2817);
nand U8529 (N_8529,N_626,N_1799);
or U8530 (N_8530,N_3975,N_1892);
xor U8531 (N_8531,N_5816,N_2409);
or U8532 (N_8532,N_2024,N_5877);
xnor U8533 (N_8533,N_1565,N_4361);
nand U8534 (N_8534,N_4901,N_5280);
and U8535 (N_8535,N_3187,N_5482);
xnor U8536 (N_8536,N_3016,N_440);
nand U8537 (N_8537,N_6217,N_431);
and U8538 (N_8538,N_4583,N_1386);
xor U8539 (N_8539,N_125,N_5514);
nand U8540 (N_8540,N_351,N_6058);
nor U8541 (N_8541,N_938,N_5465);
nand U8542 (N_8542,N_2831,N_4221);
and U8543 (N_8543,N_4825,N_6145);
nand U8544 (N_8544,N_3659,N_85);
xnor U8545 (N_8545,N_653,N_3820);
and U8546 (N_8546,N_2286,N_1954);
xnor U8547 (N_8547,N_4924,N_6013);
nand U8548 (N_8548,N_2915,N_5459);
nor U8549 (N_8549,N_2868,N_69);
or U8550 (N_8550,N_4754,N_557);
nand U8551 (N_8551,N_3215,N_5506);
nor U8552 (N_8552,N_1441,N_3992);
xor U8553 (N_8553,N_5553,N_2523);
and U8554 (N_8554,N_65,N_4006);
nand U8555 (N_8555,N_5063,N_4019);
or U8556 (N_8556,N_5639,N_3695);
xnor U8557 (N_8557,N_529,N_5691);
nand U8558 (N_8558,N_6228,N_1881);
xnor U8559 (N_8559,N_2048,N_128);
nor U8560 (N_8560,N_1214,N_2797);
nand U8561 (N_8561,N_1000,N_1409);
nand U8562 (N_8562,N_2544,N_4865);
or U8563 (N_8563,N_4451,N_3930);
nor U8564 (N_8564,N_451,N_4990);
xor U8565 (N_8565,N_4304,N_2356);
and U8566 (N_8566,N_2681,N_1234);
and U8567 (N_8567,N_2134,N_4061);
and U8568 (N_8568,N_4047,N_1262);
or U8569 (N_8569,N_2826,N_2076);
xnor U8570 (N_8570,N_318,N_899);
or U8571 (N_8571,N_1491,N_3816);
and U8572 (N_8572,N_2685,N_5165);
and U8573 (N_8573,N_2044,N_2189);
xor U8574 (N_8574,N_3535,N_3501);
nor U8575 (N_8575,N_2248,N_5262);
nand U8576 (N_8576,N_775,N_2308);
and U8577 (N_8577,N_2909,N_525);
or U8578 (N_8578,N_1489,N_3378);
xor U8579 (N_8579,N_901,N_2473);
xnor U8580 (N_8580,N_5583,N_5988);
nand U8581 (N_8581,N_5518,N_3660);
nor U8582 (N_8582,N_4659,N_2935);
or U8583 (N_8583,N_1298,N_1933);
xor U8584 (N_8584,N_3658,N_2092);
xor U8585 (N_8585,N_3763,N_3432);
nand U8586 (N_8586,N_233,N_4096);
nor U8587 (N_8587,N_6172,N_3861);
xor U8588 (N_8588,N_408,N_2228);
nor U8589 (N_8589,N_1347,N_3784);
nand U8590 (N_8590,N_3424,N_1724);
nor U8591 (N_8591,N_757,N_3098);
nand U8592 (N_8592,N_471,N_5014);
nand U8593 (N_8593,N_3668,N_4695);
or U8594 (N_8594,N_6108,N_1697);
and U8595 (N_8595,N_3945,N_1872);
nor U8596 (N_8596,N_4582,N_5021);
and U8597 (N_8597,N_770,N_5449);
nand U8598 (N_8598,N_5120,N_1370);
or U8599 (N_8599,N_6081,N_4962);
nor U8600 (N_8600,N_3359,N_2656);
xnor U8601 (N_8601,N_2728,N_4480);
nand U8602 (N_8602,N_2018,N_3230);
or U8603 (N_8603,N_1891,N_3652);
and U8604 (N_8604,N_2634,N_6109);
nand U8605 (N_8605,N_1864,N_3895);
nand U8606 (N_8606,N_1218,N_4952);
or U8607 (N_8607,N_4161,N_3546);
or U8608 (N_8608,N_4300,N_887);
and U8609 (N_8609,N_1116,N_2427);
nand U8610 (N_8610,N_2625,N_873);
nor U8611 (N_8611,N_3805,N_4666);
xor U8612 (N_8612,N_1650,N_97);
and U8613 (N_8613,N_2168,N_391);
and U8614 (N_8614,N_6087,N_4305);
or U8615 (N_8615,N_4400,N_4481);
nor U8616 (N_8616,N_479,N_590);
nand U8617 (N_8617,N_3435,N_5328);
xnor U8618 (N_8618,N_48,N_2295);
nand U8619 (N_8619,N_6213,N_4458);
nor U8620 (N_8620,N_4487,N_6070);
and U8621 (N_8621,N_4567,N_2581);
xnor U8622 (N_8622,N_240,N_1077);
nor U8623 (N_8623,N_1075,N_4036);
nor U8624 (N_8624,N_3122,N_5048);
xor U8625 (N_8625,N_1543,N_136);
nand U8626 (N_8626,N_3177,N_4366);
nor U8627 (N_8627,N_3457,N_3972);
and U8628 (N_8628,N_6045,N_3440);
and U8629 (N_8629,N_4839,N_1924);
nand U8630 (N_8630,N_13,N_4447);
nor U8631 (N_8631,N_3050,N_5882);
and U8632 (N_8632,N_889,N_5749);
nand U8633 (N_8633,N_4245,N_2642);
and U8634 (N_8634,N_2163,N_2034);
nand U8635 (N_8635,N_794,N_3401);
nor U8636 (N_8636,N_5581,N_2352);
and U8637 (N_8637,N_1514,N_1852);
and U8638 (N_8638,N_2096,N_229);
xor U8639 (N_8639,N_2288,N_1376);
nand U8640 (N_8640,N_3863,N_1958);
xnor U8641 (N_8641,N_5426,N_4573);
nor U8642 (N_8642,N_1143,N_3169);
or U8643 (N_8643,N_5618,N_597);
nand U8644 (N_8644,N_2617,N_946);
and U8645 (N_8645,N_5519,N_4512);
or U8646 (N_8646,N_2988,N_2481);
nand U8647 (N_8647,N_4619,N_416);
xor U8648 (N_8648,N_4578,N_621);
nand U8649 (N_8649,N_4317,N_4270);
xor U8650 (N_8650,N_1665,N_5043);
or U8651 (N_8651,N_4324,N_253);
xnor U8652 (N_8652,N_2380,N_3787);
xor U8653 (N_8653,N_5173,N_447);
and U8654 (N_8654,N_5363,N_4478);
nand U8655 (N_8655,N_978,N_2377);
nand U8656 (N_8656,N_4277,N_3314);
nand U8657 (N_8657,N_822,N_1101);
nor U8658 (N_8658,N_4434,N_3406);
nand U8659 (N_8659,N_3073,N_3245);
nand U8660 (N_8660,N_5586,N_4146);
nor U8661 (N_8661,N_3694,N_792);
and U8662 (N_8662,N_6030,N_2107);
nand U8663 (N_8663,N_4254,N_1740);
and U8664 (N_8664,N_2446,N_5351);
nand U8665 (N_8665,N_1662,N_6146);
and U8666 (N_8666,N_3768,N_4244);
nor U8667 (N_8667,N_3686,N_4308);
nor U8668 (N_8668,N_3905,N_3914);
or U8669 (N_8669,N_834,N_217);
xor U8670 (N_8670,N_4411,N_2601);
or U8671 (N_8671,N_3037,N_4174);
nor U8672 (N_8672,N_368,N_1839);
nand U8673 (N_8673,N_1878,N_5439);
nor U8674 (N_8674,N_2546,N_5830);
nand U8675 (N_8675,N_2152,N_1087);
xnor U8676 (N_8676,N_2556,N_2419);
nand U8677 (N_8677,N_1983,N_5324);
xnor U8678 (N_8678,N_3521,N_1952);
or U8679 (N_8679,N_3132,N_2993);
xor U8680 (N_8680,N_6127,N_6235);
xor U8681 (N_8681,N_619,N_4494);
and U8682 (N_8682,N_3781,N_3509);
nand U8683 (N_8683,N_1991,N_3107);
nand U8684 (N_8684,N_442,N_4537);
and U8685 (N_8685,N_1433,N_1224);
and U8686 (N_8686,N_112,N_3375);
nor U8687 (N_8687,N_400,N_974);
nand U8688 (N_8688,N_4020,N_1176);
nand U8689 (N_8689,N_5397,N_4534);
xnor U8690 (N_8690,N_2894,N_3395);
xnor U8691 (N_8691,N_1153,N_94);
xor U8692 (N_8692,N_2840,N_633);
nand U8693 (N_8693,N_2899,N_4113);
nor U8694 (N_8694,N_919,N_3958);
nand U8695 (N_8695,N_5826,N_3814);
xnor U8696 (N_8696,N_4598,N_5452);
xnor U8697 (N_8697,N_4376,N_1314);
nor U8698 (N_8698,N_1981,N_4427);
or U8699 (N_8699,N_1107,N_5929);
nand U8700 (N_8700,N_297,N_4640);
or U8701 (N_8701,N_5114,N_4860);
nand U8702 (N_8702,N_5963,N_3219);
or U8703 (N_8703,N_5035,N_766);
nor U8704 (N_8704,N_5654,N_2878);
xor U8705 (N_8705,N_2764,N_1570);
or U8706 (N_8706,N_5271,N_2367);
nor U8707 (N_8707,N_2533,N_935);
nand U8708 (N_8708,N_5560,N_3055);
and U8709 (N_8709,N_6243,N_1889);
or U8710 (N_8710,N_5943,N_955);
nor U8711 (N_8711,N_1046,N_1695);
xor U8712 (N_8712,N_328,N_3988);
nor U8713 (N_8713,N_5535,N_4233);
or U8714 (N_8714,N_3946,N_2583);
and U8715 (N_8715,N_2476,N_1264);
and U8716 (N_8716,N_2748,N_1011);
and U8717 (N_8717,N_2871,N_4348);
or U8718 (N_8718,N_5925,N_1227);
and U8719 (N_8719,N_4003,N_3291);
nor U8720 (N_8720,N_6036,N_4236);
or U8721 (N_8721,N_3454,N_1054);
and U8722 (N_8722,N_5401,N_5762);
and U8723 (N_8723,N_2895,N_3163);
nor U8724 (N_8724,N_2985,N_3687);
and U8725 (N_8725,N_305,N_1037);
and U8726 (N_8726,N_55,N_4291);
and U8727 (N_8727,N_4307,N_107);
nand U8728 (N_8728,N_269,N_3567);
and U8729 (N_8729,N_5164,N_2145);
or U8730 (N_8730,N_1819,N_3480);
or U8731 (N_8731,N_3807,N_5028);
nand U8732 (N_8732,N_1252,N_6248);
xnor U8733 (N_8733,N_5582,N_17);
nor U8734 (N_8734,N_4698,N_6091);
xor U8735 (N_8735,N_3965,N_220);
or U8736 (N_8736,N_5667,N_2354);
xor U8737 (N_8737,N_627,N_2702);
nor U8738 (N_8738,N_4794,N_5379);
nand U8739 (N_8739,N_3084,N_4114);
nand U8740 (N_8740,N_2493,N_5391);
nand U8741 (N_8741,N_6186,N_285);
or U8742 (N_8742,N_4522,N_5335);
nand U8743 (N_8743,N_3422,N_4688);
nand U8744 (N_8744,N_5265,N_6147);
and U8745 (N_8745,N_2322,N_301);
and U8746 (N_8746,N_1867,N_933);
xor U8747 (N_8747,N_5376,N_5544);
xor U8748 (N_8748,N_561,N_2217);
or U8749 (N_8749,N_5247,N_3855);
and U8750 (N_8750,N_4680,N_2268);
and U8751 (N_8751,N_457,N_4199);
nor U8752 (N_8752,N_1381,N_2103);
nor U8753 (N_8753,N_4519,N_2733);
xor U8754 (N_8754,N_5004,N_4892);
nor U8755 (N_8755,N_5985,N_2569);
or U8756 (N_8756,N_6136,N_1378);
and U8757 (N_8757,N_5225,N_4356);
and U8758 (N_8758,N_586,N_6033);
xnor U8759 (N_8759,N_1562,N_4569);
nor U8760 (N_8760,N_1119,N_4841);
nor U8761 (N_8761,N_2498,N_3311);
xor U8762 (N_8762,N_4928,N_2604);
nor U8763 (N_8763,N_364,N_5145);
nand U8764 (N_8764,N_6184,N_3372);
and U8765 (N_8765,N_3021,N_4403);
xor U8766 (N_8766,N_3593,N_3283);
xnor U8767 (N_8767,N_1895,N_4898);
or U8768 (N_8768,N_535,N_5195);
and U8769 (N_8769,N_2105,N_1974);
nor U8770 (N_8770,N_3617,N_1174);
and U8771 (N_8771,N_2368,N_2541);
xor U8772 (N_8772,N_1129,N_914);
and U8773 (N_8773,N_2629,N_5741);
nor U8774 (N_8774,N_385,N_251);
and U8775 (N_8775,N_1903,N_1463);
nor U8776 (N_8776,N_2117,N_2566);
nand U8777 (N_8777,N_2937,N_2808);
and U8778 (N_8778,N_2555,N_5290);
or U8779 (N_8779,N_2613,N_4066);
nand U8780 (N_8780,N_5932,N_380);
nor U8781 (N_8781,N_1578,N_438);
xnor U8782 (N_8782,N_4088,N_3526);
xor U8783 (N_8783,N_5432,N_5901);
and U8784 (N_8784,N_492,N_3100);
nor U8785 (N_8785,N_6216,N_2054);
nand U8786 (N_8786,N_2415,N_5809);
xnor U8787 (N_8787,N_2252,N_5564);
nor U8788 (N_8788,N_5169,N_511);
nand U8789 (N_8789,N_761,N_5779);
nor U8790 (N_8790,N_5315,N_5024);
and U8791 (N_8791,N_123,N_554);
or U8792 (N_8792,N_4216,N_2454);
nand U8793 (N_8793,N_4017,N_1458);
nor U8794 (N_8794,N_2013,N_907);
or U8795 (N_8795,N_24,N_472);
or U8796 (N_8796,N_5820,N_3434);
xor U8797 (N_8797,N_6069,N_870);
and U8798 (N_8798,N_3881,N_1702);
xor U8799 (N_8799,N_4940,N_1693);
nor U8800 (N_8800,N_1338,N_741);
or U8801 (N_8801,N_3030,N_1151);
or U8802 (N_8802,N_1022,N_4651);
nand U8803 (N_8803,N_1092,N_1890);
and U8804 (N_8804,N_4580,N_5009);
nand U8805 (N_8805,N_5338,N_1725);
xor U8806 (N_8806,N_2928,N_4528);
nor U8807 (N_8807,N_3237,N_6068);
or U8808 (N_8808,N_517,N_5061);
and U8809 (N_8809,N_2573,N_3007);
and U8810 (N_8810,N_3153,N_5548);
or U8811 (N_8811,N_105,N_4355);
nand U8812 (N_8812,N_3883,N_1599);
nand U8813 (N_8813,N_732,N_1080);
nor U8814 (N_8814,N_3554,N_1197);
nor U8815 (N_8815,N_4340,N_2351);
nand U8816 (N_8816,N_1185,N_2549);
nor U8817 (N_8817,N_201,N_2538);
and U8818 (N_8818,N_5186,N_4600);
nor U8819 (N_8819,N_3304,N_665);
nand U8820 (N_8820,N_4949,N_3079);
or U8821 (N_8821,N_3288,N_5442);
or U8822 (N_8822,N_3233,N_5423);
and U8823 (N_8823,N_2664,N_966);
nor U8824 (N_8824,N_4755,N_837);
nand U8825 (N_8825,N_835,N_2821);
nand U8826 (N_8826,N_2082,N_3640);
nand U8827 (N_8827,N_4826,N_3041);
xor U8828 (N_8828,N_3086,N_3377);
xnor U8829 (N_8829,N_2188,N_2638);
nand U8830 (N_8830,N_5801,N_2983);
xnor U8831 (N_8831,N_1611,N_4238);
and U8832 (N_8832,N_4068,N_1789);
nor U8833 (N_8833,N_142,N_4807);
and U8834 (N_8834,N_3829,N_5084);
xnor U8835 (N_8835,N_5177,N_838);
nand U8836 (N_8836,N_3239,N_1863);
nand U8837 (N_8837,N_2225,N_744);
nand U8838 (N_8838,N_4495,N_4763);
nor U8839 (N_8839,N_725,N_29);
nor U8840 (N_8840,N_4705,N_4926);
and U8841 (N_8841,N_5365,N_5577);
xnor U8842 (N_8842,N_866,N_3758);
or U8843 (N_8843,N_4914,N_2429);
or U8844 (N_8844,N_1273,N_6002);
xor U8845 (N_8845,N_5850,N_5347);
xor U8846 (N_8846,N_4739,N_5759);
nor U8847 (N_8847,N_756,N_137);
nor U8848 (N_8848,N_1948,N_2780);
nor U8849 (N_8849,N_6166,N_4586);
nor U8850 (N_8850,N_4264,N_5473);
or U8851 (N_8851,N_1259,N_3295);
xnor U8852 (N_8852,N_102,N_4081);
nor U8853 (N_8853,N_377,N_1712);
and U8854 (N_8854,N_3228,N_943);
and U8855 (N_8855,N_5416,N_37);
xnor U8856 (N_8856,N_884,N_2614);
nand U8857 (N_8857,N_3425,N_591);
nand U8858 (N_8858,N_1392,N_4980);
nor U8859 (N_8859,N_224,N_760);
nor U8860 (N_8860,N_1015,N_929);
or U8861 (N_8861,N_3135,N_5720);
and U8862 (N_8862,N_6099,N_2369);
nor U8863 (N_8863,N_2243,N_4401);
xor U8864 (N_8864,N_2439,N_1285);
nor U8865 (N_8865,N_5620,N_4285);
and U8866 (N_8866,N_4912,N_5641);
and U8867 (N_8867,N_4948,N_807);
or U8868 (N_8868,N_5129,N_3944);
nand U8869 (N_8869,N_5954,N_1879);
or U8870 (N_8870,N_1199,N_4661);
nor U8871 (N_8871,N_3337,N_2162);
xor U8872 (N_8872,N_6110,N_1745);
xnor U8873 (N_8873,N_1574,N_1244);
nor U8874 (N_8874,N_5320,N_3904);
xor U8875 (N_8875,N_5059,N_2872);
nand U8876 (N_8876,N_208,N_3804);
nor U8877 (N_8877,N_2387,N_4108);
nor U8878 (N_8878,N_1447,N_4604);
or U8879 (N_8879,N_5344,N_410);
nor U8880 (N_8880,N_270,N_4016);
and U8881 (N_8881,N_3841,N_22);
nand U8882 (N_8882,N_276,N_75);
xor U8883 (N_8883,N_1956,N_3013);
or U8884 (N_8884,N_6024,N_1175);
xor U8885 (N_8885,N_1741,N_4894);
nor U8886 (N_8886,N_2402,N_164);
nor U8887 (N_8887,N_2178,N_4579);
nand U8888 (N_8888,N_4652,N_2779);
or U8889 (N_8889,N_3034,N_1444);
nor U8890 (N_8890,N_4609,N_1144);
nand U8891 (N_8891,N_1786,N_4182);
or U8892 (N_8892,N_474,N_3543);
xor U8893 (N_8893,N_6128,N_1271);
nor U8894 (N_8894,N_1230,N_1133);
or U8895 (N_8895,N_284,N_4209);
xnor U8896 (N_8896,N_3574,N_3740);
nand U8897 (N_8897,N_4548,N_818);
xnor U8898 (N_8898,N_2139,N_1130);
nor U8899 (N_8899,N_3093,N_4557);
or U8900 (N_8900,N_1440,N_4377);
and U8901 (N_8901,N_3056,N_5941);
or U8902 (N_8902,N_2906,N_5366);
or U8903 (N_8903,N_5258,N_3947);
xnor U8904 (N_8904,N_4607,N_114);
nor U8905 (N_8905,N_1167,N_636);
nor U8906 (N_8906,N_3900,N_4667);
nand U8907 (N_8907,N_5857,N_4945);
or U8908 (N_8908,N_3974,N_327);
nor U8909 (N_8909,N_53,N_2414);
xnor U8910 (N_8910,N_2621,N_1348);
and U8911 (N_8911,N_1454,N_1871);
or U8912 (N_8912,N_165,N_5368);
xor U8913 (N_8913,N_2890,N_819);
or U8914 (N_8914,N_2655,N_3103);
xnor U8915 (N_8915,N_230,N_6160);
nor U8916 (N_8916,N_5905,N_2609);
nand U8917 (N_8917,N_3803,N_2683);
and U8918 (N_8918,N_4723,N_4620);
and U8919 (N_8919,N_2793,N_1216);
nand U8920 (N_8920,N_782,N_31);
or U8921 (N_8921,N_1118,N_139);
nand U8922 (N_8922,N_4386,N_804);
nand U8923 (N_8923,N_1427,N_4379);
xnor U8924 (N_8924,N_3173,N_5846);
nor U8925 (N_8925,N_428,N_5504);
and U8926 (N_8926,N_3114,N_5097);
or U8927 (N_8927,N_2242,N_3685);
and U8928 (N_8928,N_4467,N_2967);
xnor U8929 (N_8929,N_2932,N_5900);
and U8930 (N_8930,N_4172,N_4768);
xnor U8931 (N_8931,N_5302,N_2116);
nor U8932 (N_8932,N_1950,N_5675);
xnor U8933 (N_8933,N_3612,N_1775);
nand U8934 (N_8934,N_6112,N_3256);
and U8935 (N_8935,N_6052,N_5428);
xnor U8936 (N_8936,N_1064,N_4727);
nand U8937 (N_8937,N_2695,N_3532);
nand U8938 (N_8938,N_1546,N_47);
nand U8939 (N_8939,N_5802,N_1277);
xor U8940 (N_8940,N_2180,N_6000);
and U8941 (N_8941,N_3048,N_915);
nand U8942 (N_8942,N_1111,N_3743);
or U8943 (N_8943,N_1303,N_2363);
or U8944 (N_8944,N_2814,N_5045);
or U8945 (N_8945,N_2947,N_1685);
or U8946 (N_8946,N_153,N_1731);
nand U8947 (N_8947,N_713,N_5763);
nand U8948 (N_8948,N_3739,N_4018);
nand U8949 (N_8949,N_3708,N_2461);
xor U8950 (N_8950,N_1776,N_5916);
and U8951 (N_8951,N_205,N_2421);
nand U8952 (N_8952,N_1681,N_2689);
nor U8953 (N_8953,N_2846,N_1990);
and U8954 (N_8954,N_1049,N_567);
nand U8955 (N_8955,N_2810,N_1332);
or U8956 (N_8956,N_1527,N_2588);
nor U8957 (N_8957,N_5270,N_1783);
xnor U8958 (N_8958,N_1913,N_3192);
nor U8959 (N_8959,N_659,N_4568);
and U8960 (N_8960,N_104,N_4093);
nand U8961 (N_8961,N_2571,N_1985);
or U8962 (N_8962,N_1018,N_1240);
and U8963 (N_8963,N_1521,N_5125);
and U8964 (N_8964,N_4504,N_5479);
nor U8965 (N_8965,N_1926,N_4729);
or U8966 (N_8966,N_1555,N_2989);
xor U8967 (N_8967,N_1815,N_5256);
and U8968 (N_8968,N_5219,N_2019);
xnor U8969 (N_8969,N_3125,N_422);
and U8970 (N_8970,N_1883,N_186);
or U8971 (N_8971,N_5686,N_6208);
xor U8972 (N_8972,N_288,N_1300);
or U8973 (N_8973,N_4677,N_2485);
and U8974 (N_8974,N_667,N_734);
and U8975 (N_8975,N_3373,N_4893);
or U8976 (N_8976,N_1384,N_2585);
nor U8977 (N_8977,N_3516,N_2487);
xor U8978 (N_8978,N_1690,N_3281);
and U8979 (N_8979,N_2848,N_2297);
xnor U8980 (N_8980,N_2595,N_1419);
nor U8981 (N_8981,N_4220,N_958);
and U8982 (N_8982,N_2465,N_5576);
xor U8983 (N_8983,N_3303,N_5119);
or U8984 (N_8984,N_1627,N_1177);
and U8985 (N_8985,N_32,N_4160);
xor U8986 (N_8986,N_143,N_4649);
nand U8987 (N_8987,N_5848,N_3806);
nand U8988 (N_8988,N_5253,N_5354);
xnor U8989 (N_8989,N_4594,N_5616);
xor U8990 (N_8990,N_4212,N_3482);
and U8991 (N_8991,N_4383,N_2083);
xnor U8992 (N_8992,N_1147,N_3796);
and U8993 (N_8993,N_3006,N_1184);
and U8994 (N_8994,N_5859,N_4555);
nor U8995 (N_8995,N_2863,N_699);
and U8996 (N_8996,N_5398,N_131);
nand U8997 (N_8997,N_3223,N_1327);
xnor U8998 (N_8998,N_521,N_4906);
nor U8999 (N_8999,N_4343,N_3243);
nand U9000 (N_9000,N_610,N_2434);
and U9001 (N_9001,N_1766,N_2769);
and U9002 (N_9002,N_598,N_5);
xor U9003 (N_9003,N_5019,N_5902);
xor U9004 (N_9004,N_6173,N_2093);
and U9005 (N_9005,N_3178,N_2378);
nor U9006 (N_9006,N_2680,N_4084);
nand U9007 (N_9007,N_3403,N_3113);
nor U9008 (N_9008,N_3470,N_19);
and U9009 (N_9009,N_5866,N_710);
and U9010 (N_9010,N_1589,N_3717);
nor U9011 (N_9011,N_5092,N_4545);
or U9012 (N_9012,N_2108,N_5731);
or U9013 (N_9013,N_5687,N_4158);
nor U9014 (N_9014,N_594,N_711);
xor U9015 (N_9015,N_995,N_4085);
nor U9016 (N_9016,N_1609,N_1886);
nand U9017 (N_9017,N_5339,N_2874);
and U9018 (N_9018,N_5517,N_3889);
and U9019 (N_9019,N_3046,N_5880);
xor U9020 (N_9020,N_680,N_5307);
nor U9021 (N_9021,N_5182,N_574);
xnor U9022 (N_9022,N_3309,N_3476);
nor U9023 (N_9023,N_2563,N_1726);
or U9024 (N_9024,N_4571,N_516);
or U9025 (N_9025,N_3354,N_718);
nor U9026 (N_9026,N_2304,N_5183);
nor U9027 (N_9027,N_1342,N_1540);
or U9028 (N_9028,N_3932,N_3405);
nand U9029 (N_9029,N_3561,N_5719);
nor U9030 (N_9030,N_4075,N_3676);
xor U9031 (N_9031,N_4933,N_5883);
or U9032 (N_9032,N_1987,N_5748);
or U9033 (N_9033,N_4091,N_1512);
and U9034 (N_9034,N_2643,N_1649);
xnor U9035 (N_9035,N_1660,N_4249);
xor U9036 (N_9036,N_2463,N_5279);
nand U9037 (N_9037,N_1267,N_379);
xor U9038 (N_9038,N_2345,N_100);
nor U9039 (N_9039,N_5016,N_1005);
nand U9040 (N_9040,N_4010,N_3029);
nand U9041 (N_9041,N_5412,N_5878);
and U9042 (N_9042,N_707,N_242);
nand U9043 (N_9043,N_403,N_5050);
nor U9044 (N_9044,N_4162,N_2636);
nor U9045 (N_9045,N_4222,N_2266);
xnor U9046 (N_9046,N_1739,N_4218);
nand U9047 (N_9047,N_6247,N_3044);
or U9048 (N_9048,N_3236,N_3428);
and U9049 (N_9049,N_1016,N_3072);
and U9050 (N_9050,N_1249,N_564);
and U9051 (N_9051,N_1915,N_3569);
or U9052 (N_9052,N_6157,N_2784);
nand U9053 (N_9053,N_4811,N_5584);
and U9054 (N_9054,N_1654,N_604);
and U9055 (N_9055,N_339,N_3267);
nor U9056 (N_9056,N_373,N_4835);
nand U9057 (N_9057,N_2316,N_4267);
and U9058 (N_9058,N_2950,N_3525);
nor U9059 (N_9059,N_1673,N_3181);
and U9060 (N_9060,N_4840,N_2328);
nor U9061 (N_9061,N_861,N_5340);
and U9062 (N_9062,N_5737,N_2353);
xnor U9063 (N_9063,N_383,N_3361);
nor U9064 (N_9064,N_5509,N_2418);
xor U9065 (N_9065,N_278,N_3901);
and U9066 (N_9066,N_4268,N_1989);
nand U9067 (N_9067,N_1226,N_4226);
nand U9068 (N_9068,N_4183,N_4803);
nor U9069 (N_9069,N_4271,N_195);
xnor U9070 (N_9070,N_3924,N_173);
or U9071 (N_9071,N_3788,N_5360);
xnor U9072 (N_9072,N_4539,N_2218);
and U9073 (N_9073,N_5316,N_3390);
xor U9074 (N_9074,N_1414,N_3887);
nor U9075 (N_9075,N_3870,N_1544);
nand U9076 (N_9076,N_1835,N_3499);
and U9077 (N_9077,N_5072,N_3698);
or U9078 (N_9078,N_1575,N_1351);
xor U9079 (N_9079,N_3437,N_2758);
nand U9080 (N_9080,N_2517,N_4175);
and U9081 (N_9081,N_1272,N_1356);
nor U9082 (N_9082,N_5800,N_844);
or U9083 (N_9083,N_3200,N_394);
or U9084 (N_9084,N_4353,N_1586);
and U9085 (N_9085,N_6061,N_2355);
nand U9086 (N_9086,N_2657,N_4148);
and U9087 (N_9087,N_5947,N_1172);
xnor U9088 (N_9088,N_314,N_372);
xor U9089 (N_9089,N_1502,N_3347);
xnor U9090 (N_9090,N_3871,N_657);
xnor U9091 (N_9091,N_2501,N_486);
or U9092 (N_9092,N_813,N_5944);
and U9093 (N_9093,N_3920,N_5512);
nand U9094 (N_9094,N_3360,N_5824);
and U9095 (N_9095,N_3732,N_2424);
and U9096 (N_9096,N_12,N_2255);
nor U9097 (N_9097,N_526,N_3540);
or U9098 (N_9098,N_6192,N_2191);
nand U9099 (N_9099,N_1888,N_2710);
and U9100 (N_9100,N_1964,N_3190);
xnor U9101 (N_9101,N_4645,N_2857);
nor U9102 (N_9102,N_4577,N_5520);
xor U9103 (N_9103,N_1091,N_331);
or U9104 (N_9104,N_3565,N_340);
nand U9105 (N_9105,N_2876,N_2017);
nor U9106 (N_9106,N_3961,N_87);
nand U9107 (N_9107,N_3312,N_4294);
xnor U9108 (N_9108,N_6121,N_3845);
or U9109 (N_9109,N_5491,N_4517);
nand U9110 (N_9110,N_1700,N_4189);
nand U9111 (N_9111,N_252,N_2716);
xor U9112 (N_9112,N_3268,N_632);
nand U9113 (N_9113,N_777,N_6122);
nor U9114 (N_9114,N_2196,N_3604);
xnor U9115 (N_9115,N_1,N_1764);
or U9116 (N_9116,N_676,N_5557);
or U9117 (N_9117,N_315,N_5871);
or U9118 (N_9118,N_5764,N_3388);
and U9119 (N_9119,N_4726,N_1711);
or U9120 (N_9120,N_4631,N_4792);
or U9121 (N_9121,N_2958,N_2275);
nand U9122 (N_9122,N_1623,N_2882);
nand U9123 (N_9123,N_765,N_3906);
or U9124 (N_9124,N_1109,N_1652);
nand U9125 (N_9125,N_498,N_1525);
and U9126 (N_9126,N_6078,N_6179);
xnor U9127 (N_9127,N_4678,N_432);
xnor U9128 (N_9128,N_4874,N_3622);
nor U9129 (N_9129,N_3442,N_1358);
nand U9130 (N_9130,N_1159,N_6197);
nor U9131 (N_9131,N_5970,N_96);
nor U9132 (N_9132,N_571,N_244);
xnor U9133 (N_9133,N_2738,N_2977);
and U9134 (N_9134,N_404,N_6063);
nand U9135 (N_9135,N_4637,N_1282);
xnor U9136 (N_9136,N_215,N_890);
xnor U9137 (N_9137,N_2850,N_5441);
nor U9138 (N_9138,N_5887,N_4947);
xor U9139 (N_9139,N_5104,N_649);
nand U9140 (N_9140,N_4402,N_1212);
nand U9141 (N_9141,N_4382,N_1620);
and U9142 (N_9142,N_5803,N_5108);
and U9143 (N_9143,N_5684,N_2025);
nor U9144 (N_9144,N_2939,N_4738);
xor U9145 (N_9145,N_5844,N_1286);
nand U9146 (N_9146,N_499,N_5688);
xnor U9147 (N_9147,N_5593,N_3487);
nand U9148 (N_9148,N_4344,N_1828);
or U9149 (N_9149,N_922,N_1344);
nand U9150 (N_9150,N_5872,N_2830);
nor U9151 (N_9151,N_650,N_5232);
nor U9152 (N_9152,N_4080,N_5757);
and U9153 (N_9153,N_2514,N_5283);
and U9154 (N_9154,N_1181,N_1421);
nand U9155 (N_9155,N_3936,N_5322);
xor U9156 (N_9156,N_2513,N_3339);
xor U9157 (N_9157,N_5775,N_4042);
nor U9158 (N_9158,N_855,N_5812);
and U9159 (N_9159,N_4274,N_475);
and U9160 (N_9160,N_509,N_5417);
xnor U9161 (N_9161,N_664,N_5241);
and U9162 (N_9162,N_4509,N_1501);
nand U9163 (N_9163,N_5102,N_3335);
nor U9164 (N_9164,N_4,N_2249);
nand U9165 (N_9165,N_2488,N_4139);
nor U9166 (N_9166,N_994,N_1284);
nor U9167 (N_9167,N_2704,N_5679);
and U9168 (N_9168,N_1451,N_5403);
or U9169 (N_9169,N_3539,N_3250);
and U9170 (N_9170,N_1360,N_2056);
or U9171 (N_9171,N_5434,N_5337);
nor U9172 (N_9172,N_5999,N_390);
nor U9173 (N_9173,N_5187,N_187);
xor U9174 (N_9174,N_2952,N_2472);
nand U9175 (N_9175,N_4783,N_2426);
nor U9176 (N_9176,N_3276,N_5602);
nor U9177 (N_9177,N_1535,N_1604);
and U9178 (N_9178,N_1480,N_1572);
nand U9179 (N_9179,N_3277,N_5185);
and U9180 (N_9180,N_5722,N_584);
or U9181 (N_9181,N_3588,N_5540);
nor U9182 (N_9182,N_2155,N_5659);
nor U9183 (N_9183,N_5796,N_3682);
xnor U9184 (N_9184,N_3627,N_4641);
nand U9185 (N_9185,N_1498,N_3661);
xnor U9186 (N_9186,N_1465,N_4007);
or U9187 (N_9187,N_501,N_5897);
nand U9188 (N_9188,N_3778,N_1894);
nor U9189 (N_9189,N_4159,N_1639);
nand U9190 (N_9190,N_4873,N_5060);
or U9191 (N_9191,N_4615,N_6044);
and U9192 (N_9192,N_6032,N_4219);
nor U9193 (N_9193,N_3842,N_752);
xor U9194 (N_9194,N_2503,N_812);
nand U9195 (N_9195,N_30,N_2559);
xor U9196 (N_9196,N_4499,N_2193);
or U9197 (N_9197,N_5579,N_1355);
or U9198 (N_9198,N_893,N_799);
and U9199 (N_9199,N_5648,N_1248);
and U9200 (N_9200,N_5306,N_5508);
or U9201 (N_9201,N_2097,N_4247);
and U9202 (N_9202,N_1746,N_1095);
nand U9203 (N_9203,N_1862,N_3427);
xnor U9204 (N_9204,N_1405,N_1744);
and U9205 (N_9205,N_2104,N_5146);
xnor U9206 (N_9206,N_5689,N_3071);
xnor U9207 (N_9207,N_4056,N_5896);
and U9208 (N_9208,N_3576,N_5852);
xor U9209 (N_9209,N_814,N_2130);
xnor U9210 (N_9210,N_3096,N_2341);
nand U9211 (N_9211,N_980,N_5928);
xor U9212 (N_9212,N_1708,N_4450);
xnor U9213 (N_9213,N_2842,N_729);
nor U9214 (N_9214,N_2597,N_5377);
and U9215 (N_9215,N_5220,N_414);
nand U9216 (N_9216,N_1110,N_795);
xnor U9217 (N_9217,N_1025,N_4086);
and U9218 (N_9218,N_1635,N_3123);
nor U9219 (N_9219,N_1942,N_4242);
or U9220 (N_9220,N_2707,N_434);
or U9221 (N_9221,N_5547,N_4981);
nor U9222 (N_9222,N_5628,N_1052);
and U9223 (N_9223,N_4672,N_1769);
xnor U9224 (N_9224,N_2232,N_2535);
xnor U9225 (N_9225,N_897,N_4365);
nor U9226 (N_9226,N_5714,N_5658);
nor U9227 (N_9227,N_4168,N_2819);
or U9228 (N_9228,N_2122,N_6051);
nor U9229 (N_9229,N_843,N_1254);
nand U9230 (N_9230,N_5951,N_6092);
xnor U9231 (N_9231,N_1499,N_4315);
or U9232 (N_9232,N_957,N_2804);
xnor U9233 (N_9233,N_4721,N_1736);
nand U9234 (N_9234,N_4634,N_4046);
nor U9235 (N_9235,N_2319,N_1587);
and U9236 (N_9236,N_4679,N_1403);
nand U9237 (N_9237,N_3198,N_3566);
nand U9238 (N_9238,N_4833,N_4922);
nand U9239 (N_9239,N_2953,N_715);
nor U9240 (N_9240,N_3278,N_3194);
or U9241 (N_9241,N_5601,N_3446);
or U9242 (N_9242,N_4706,N_4319);
xnor U9243 (N_9243,N_2788,N_4995);
xor U9244 (N_9244,N_5049,N_1350);
or U9245 (N_9245,N_2246,N_2767);
or U9246 (N_9246,N_5374,N_1921);
or U9247 (N_9247,N_5470,N_1382);
xor U9248 (N_9248,N_771,N_869);
nand U9249 (N_9249,N_1717,N_944);
nor U9250 (N_9250,N_3146,N_2827);
or U9251 (N_9251,N_155,N_3754);
xor U9252 (N_9252,N_2933,N_4696);
nand U9253 (N_9253,N_749,N_4932);
xnor U9254 (N_9254,N_1004,N_2451);
or U9255 (N_9255,N_5485,N_4741);
nand U9256 (N_9256,N_4905,N_3443);
or U9257 (N_9257,N_4473,N_790);
xor U9258 (N_9258,N_336,N_2944);
and U9259 (N_9259,N_4957,N_4875);
xor U9260 (N_9260,N_4527,N_4908);
and U9261 (N_9261,N_5915,N_3320);
nor U9262 (N_9262,N_1807,N_2317);
xnor U9263 (N_9263,N_801,N_606);
xor U9264 (N_9264,N_4298,N_3896);
nor U9265 (N_9265,N_5671,N_63);
and U9266 (N_9266,N_5744,N_5472);
xor U9267 (N_9267,N_1363,N_809);
nor U9268 (N_9268,N_4805,N_2301);
and U9269 (N_9269,N_2973,N_5246);
and U9270 (N_9270,N_5082,N_2499);
or U9271 (N_9271,N_6169,N_4136);
or U9272 (N_9272,N_1626,N_4996);
nor U9273 (N_9273,N_2303,N_3111);
nand U9274 (N_9274,N_4459,N_3344);
and U9275 (N_9275,N_5168,N_5610);
and U9276 (N_9276,N_3544,N_4910);
and U9277 (N_9277,N_2594,N_4941);
xnor U9278 (N_9278,N_1953,N_2110);
xor U9279 (N_9279,N_2455,N_4201);
nor U9280 (N_9280,N_1425,N_135);
xor U9281 (N_9281,N_3489,N_4946);
xnor U9282 (N_9282,N_3587,N_3688);
nand U9283 (N_9283,N_928,N_1659);
and U9284 (N_9284,N_3386,N_3776);
nand U9285 (N_9285,N_4703,N_4156);
and U9286 (N_9286,N_2900,N_283);
or U9287 (N_9287,N_2066,N_864);
and U9288 (N_9288,N_6137,N_2229);
nand U9289 (N_9289,N_5822,N_2020);
and U9290 (N_9290,N_1939,N_6221);
and U9291 (N_9291,N_2885,N_5873);
nand U9292 (N_9292,N_704,N_395);
or U9293 (N_9293,N_547,N_33);
nand U9294 (N_9294,N_4065,N_4722);
nand U9295 (N_9295,N_5455,N_3890);
nand U9296 (N_9296,N_1577,N_3069);
and U9297 (N_9297,N_2801,N_3886);
and U9298 (N_9298,N_3342,N_5447);
nor U9299 (N_9299,N_4205,N_213);
nand U9300 (N_9300,N_1767,N_1001);
and U9301 (N_9301,N_911,N_5588);
nor U9302 (N_9302,N_6222,N_2622);
nand U9303 (N_9303,N_182,N_5499);
or U9304 (N_9304,N_1938,N_4503);
or U9305 (N_9305,N_2087,N_6153);
or U9306 (N_9306,N_176,N_4073);
nand U9307 (N_9307,N_3150,N_3019);
nor U9308 (N_9308,N_4972,N_1135);
or U9309 (N_9309,N_5605,N_5546);
and U9310 (N_9310,N_2146,N_1010);
nor U9311 (N_9311,N_2211,N_2224);
xor U9312 (N_9312,N_1196,N_2250);
nor U9313 (N_9313,N_712,N_2916);
nand U9314 (N_9314,N_2587,N_4973);
nor U9315 (N_9315,N_2987,N_6079);
or U9316 (N_9316,N_6171,N_1549);
nand U9317 (N_9317,N_6225,N_5838);
or U9318 (N_9318,N_4529,N_3989);
nand U9319 (N_9319,N_5178,N_4173);
xnor U9320 (N_9320,N_3799,N_4507);
and U9321 (N_9321,N_2729,N_1962);
xnor U9322 (N_9322,N_2038,N_374);
and U9323 (N_9323,N_3368,N_881);
nor U9324 (N_9324,N_857,N_2441);
nor U9325 (N_9325,N_2312,N_1818);
nor U9326 (N_9326,N_1946,N_3105);
nand U9327 (N_9327,N_1055,N_3199);
nor U9328 (N_9328,N_5652,N_1814);
nor U9329 (N_9329,N_2149,N_1497);
nand U9330 (N_9330,N_3461,N_549);
nand U9331 (N_9331,N_130,N_5079);
or U9332 (N_9332,N_6113,N_4915);
xor U9333 (N_9333,N_3728,N_786);
or U9334 (N_9334,N_5474,N_3467);
xor U9335 (N_9335,N_4200,N_2440);
and U9336 (N_9336,N_3738,N_4163);
xnor U9337 (N_9337,N_896,N_802);
nand U9338 (N_9338,N_3374,N_997);
nand U9339 (N_9339,N_4070,N_1120);
or U9340 (N_9340,N_637,N_6123);
nand U9341 (N_9341,N_5190,N_5329);
xor U9342 (N_9342,N_3195,N_4423);
nor U9343 (N_9343,N_460,N_4074);
xor U9344 (N_9344,N_1113,N_3094);
nor U9345 (N_9345,N_3615,N_3384);
nand U9346 (N_9346,N_2494,N_5515);
and U9347 (N_9347,N_2805,N_238);
nand U9348 (N_9348,N_4059,N_1485);
and U9349 (N_9349,N_3876,N_290);
or U9350 (N_9350,N_1568,N_3908);
nand U9351 (N_9351,N_2040,N_5590);
or U9352 (N_9352,N_1476,N_3751);
nand U9353 (N_9353,N_4443,N_5500);
and U9354 (N_9354,N_5598,N_4574);
xor U9355 (N_9355,N_3641,N_5917);
nor U9356 (N_9356,N_5375,N_200);
or U9357 (N_9357,N_5587,N_1523);
and U9358 (N_9358,N_4491,N_2507);
and U9359 (N_9359,N_3409,N_2375);
nand U9360 (N_9360,N_924,N_5969);
xnor U9361 (N_9361,N_3993,N_1100);
and U9362 (N_9362,N_4250,N_5135);
nor U9363 (N_9363,N_2021,N_3599);
nand U9364 (N_9364,N_5058,N_5032);
or U9365 (N_9365,N_2734,N_1547);
xor U9366 (N_9366,N_3834,N_965);
nor U9367 (N_9367,N_3978,N_4118);
or U9368 (N_9368,N_4636,N_3613);
and U9369 (N_9369,N_192,N_4844);
and U9370 (N_9370,N_3927,N_5240);
and U9371 (N_9371,N_4217,N_2203);
nor U9372 (N_9372,N_3850,N_4398);
or U9373 (N_9373,N_369,N_1817);
nor U9374 (N_9374,N_6055,N_692);
and U9375 (N_9375,N_860,N_2966);
nand U9376 (N_9376,N_3809,N_715);
nor U9377 (N_9377,N_2090,N_859);
xor U9378 (N_9378,N_5644,N_5778);
nand U9379 (N_9379,N_273,N_4330);
nor U9380 (N_9380,N_4686,N_5475);
xor U9381 (N_9381,N_743,N_241);
nand U9382 (N_9382,N_673,N_2023);
nand U9383 (N_9383,N_4678,N_1349);
nand U9384 (N_9384,N_626,N_3012);
nand U9385 (N_9385,N_1406,N_864);
xor U9386 (N_9386,N_4710,N_3104);
or U9387 (N_9387,N_3466,N_46);
xor U9388 (N_9388,N_4457,N_295);
nor U9389 (N_9389,N_4891,N_1675);
nor U9390 (N_9390,N_3923,N_6207);
xnor U9391 (N_9391,N_387,N_3735);
nand U9392 (N_9392,N_554,N_4548);
nor U9393 (N_9393,N_553,N_3531);
or U9394 (N_9394,N_3884,N_5590);
nand U9395 (N_9395,N_593,N_581);
or U9396 (N_9396,N_1196,N_5126);
nand U9397 (N_9397,N_2077,N_5311);
xnor U9398 (N_9398,N_1898,N_4906);
nor U9399 (N_9399,N_5661,N_3023);
xnor U9400 (N_9400,N_5113,N_595);
and U9401 (N_9401,N_5770,N_118);
xor U9402 (N_9402,N_3531,N_4443);
nand U9403 (N_9403,N_3943,N_675);
or U9404 (N_9404,N_3595,N_247);
nor U9405 (N_9405,N_1136,N_498);
and U9406 (N_9406,N_953,N_1595);
or U9407 (N_9407,N_1184,N_5108);
or U9408 (N_9408,N_5889,N_5991);
nor U9409 (N_9409,N_2428,N_5269);
xnor U9410 (N_9410,N_2149,N_1745);
or U9411 (N_9411,N_1639,N_300);
nand U9412 (N_9412,N_4025,N_1691);
xnor U9413 (N_9413,N_5466,N_214);
nor U9414 (N_9414,N_3277,N_3049);
and U9415 (N_9415,N_1795,N_1283);
and U9416 (N_9416,N_2301,N_1219);
xor U9417 (N_9417,N_136,N_4983);
nor U9418 (N_9418,N_2057,N_4330);
or U9419 (N_9419,N_4158,N_3489);
and U9420 (N_9420,N_2380,N_4937);
or U9421 (N_9421,N_5764,N_3544);
or U9422 (N_9422,N_3373,N_3556);
xnor U9423 (N_9423,N_5873,N_4411);
xnor U9424 (N_9424,N_3149,N_5907);
or U9425 (N_9425,N_1687,N_1058);
or U9426 (N_9426,N_26,N_5580);
nand U9427 (N_9427,N_1941,N_4408);
or U9428 (N_9428,N_546,N_2995);
nand U9429 (N_9429,N_4806,N_1463);
nand U9430 (N_9430,N_2257,N_3783);
xor U9431 (N_9431,N_4458,N_1844);
xor U9432 (N_9432,N_30,N_4265);
and U9433 (N_9433,N_5041,N_4387);
or U9434 (N_9434,N_4514,N_1221);
or U9435 (N_9435,N_2866,N_2311);
nor U9436 (N_9436,N_3873,N_2454);
and U9437 (N_9437,N_967,N_1039);
or U9438 (N_9438,N_4490,N_1303);
nand U9439 (N_9439,N_5711,N_951);
or U9440 (N_9440,N_5225,N_6193);
xnor U9441 (N_9441,N_6047,N_5541);
xor U9442 (N_9442,N_4838,N_1671);
nor U9443 (N_9443,N_700,N_102);
nand U9444 (N_9444,N_1179,N_4027);
nor U9445 (N_9445,N_2602,N_4154);
and U9446 (N_9446,N_5261,N_5910);
and U9447 (N_9447,N_1545,N_2108);
nand U9448 (N_9448,N_1003,N_5633);
nand U9449 (N_9449,N_207,N_5051);
or U9450 (N_9450,N_1683,N_2849);
or U9451 (N_9451,N_98,N_1109);
and U9452 (N_9452,N_5081,N_2385);
or U9453 (N_9453,N_3974,N_111);
and U9454 (N_9454,N_3743,N_4020);
nor U9455 (N_9455,N_4956,N_505);
or U9456 (N_9456,N_5156,N_2564);
or U9457 (N_9457,N_3160,N_1150);
nand U9458 (N_9458,N_4142,N_3928);
and U9459 (N_9459,N_3502,N_2549);
nor U9460 (N_9460,N_3229,N_2908);
or U9461 (N_9461,N_4695,N_4129);
xor U9462 (N_9462,N_4418,N_2432);
nand U9463 (N_9463,N_1622,N_1112);
nand U9464 (N_9464,N_3590,N_1058);
and U9465 (N_9465,N_5797,N_145);
xor U9466 (N_9466,N_4854,N_4920);
xor U9467 (N_9467,N_6052,N_5002);
nor U9468 (N_9468,N_5864,N_3903);
and U9469 (N_9469,N_4984,N_1336);
or U9470 (N_9470,N_6074,N_3810);
and U9471 (N_9471,N_4806,N_5849);
nand U9472 (N_9472,N_4962,N_5522);
and U9473 (N_9473,N_2567,N_1012);
nor U9474 (N_9474,N_5549,N_2491);
or U9475 (N_9475,N_4214,N_747);
or U9476 (N_9476,N_863,N_5638);
nor U9477 (N_9477,N_5566,N_1478);
nand U9478 (N_9478,N_3233,N_4697);
or U9479 (N_9479,N_1051,N_3655);
nand U9480 (N_9480,N_1581,N_2506);
or U9481 (N_9481,N_1224,N_3662);
xor U9482 (N_9482,N_5395,N_2303);
nor U9483 (N_9483,N_3654,N_3965);
or U9484 (N_9484,N_5912,N_2244);
and U9485 (N_9485,N_4343,N_2464);
nand U9486 (N_9486,N_1282,N_2322);
nor U9487 (N_9487,N_1066,N_87);
nor U9488 (N_9488,N_1996,N_4173);
or U9489 (N_9489,N_1422,N_3200);
xor U9490 (N_9490,N_109,N_1262);
or U9491 (N_9491,N_4394,N_5096);
xor U9492 (N_9492,N_3577,N_3742);
xor U9493 (N_9493,N_1725,N_537);
nor U9494 (N_9494,N_2833,N_5040);
nand U9495 (N_9495,N_5642,N_1982);
and U9496 (N_9496,N_1222,N_3256);
or U9497 (N_9497,N_2766,N_1167);
nand U9498 (N_9498,N_382,N_4557);
nand U9499 (N_9499,N_1015,N_714);
and U9500 (N_9500,N_771,N_5521);
and U9501 (N_9501,N_3961,N_5209);
xor U9502 (N_9502,N_2747,N_2553);
xnor U9503 (N_9503,N_4744,N_1548);
xnor U9504 (N_9504,N_1386,N_3944);
xor U9505 (N_9505,N_6210,N_1013);
nand U9506 (N_9506,N_3234,N_1311);
xor U9507 (N_9507,N_874,N_1893);
or U9508 (N_9508,N_755,N_1123);
and U9509 (N_9509,N_6201,N_1103);
xor U9510 (N_9510,N_502,N_4179);
nor U9511 (N_9511,N_3519,N_258);
nand U9512 (N_9512,N_4973,N_4907);
or U9513 (N_9513,N_1276,N_2300);
nand U9514 (N_9514,N_724,N_2971);
xnor U9515 (N_9515,N_6138,N_5702);
xnor U9516 (N_9516,N_6052,N_6144);
or U9517 (N_9517,N_4630,N_2371);
or U9518 (N_9518,N_4195,N_945);
or U9519 (N_9519,N_3367,N_2888);
nor U9520 (N_9520,N_4138,N_5039);
and U9521 (N_9521,N_4828,N_4469);
nand U9522 (N_9522,N_959,N_3245);
and U9523 (N_9523,N_4462,N_4044);
and U9524 (N_9524,N_5473,N_3868);
or U9525 (N_9525,N_2288,N_135);
nor U9526 (N_9526,N_2703,N_2675);
nand U9527 (N_9527,N_2702,N_2298);
nand U9528 (N_9528,N_2251,N_1349);
nor U9529 (N_9529,N_4609,N_3411);
xor U9530 (N_9530,N_1257,N_1743);
xor U9531 (N_9531,N_4917,N_1992);
and U9532 (N_9532,N_6014,N_5713);
nor U9533 (N_9533,N_6057,N_278);
and U9534 (N_9534,N_251,N_2819);
xor U9535 (N_9535,N_4476,N_3138);
xor U9536 (N_9536,N_4555,N_4256);
xnor U9537 (N_9537,N_2510,N_3766);
nor U9538 (N_9538,N_558,N_1593);
and U9539 (N_9539,N_3290,N_5930);
xor U9540 (N_9540,N_4737,N_2237);
and U9541 (N_9541,N_3719,N_2395);
nand U9542 (N_9542,N_957,N_3049);
nor U9543 (N_9543,N_4759,N_3465);
nand U9544 (N_9544,N_4489,N_3376);
and U9545 (N_9545,N_5876,N_5978);
nand U9546 (N_9546,N_614,N_3478);
xnor U9547 (N_9547,N_2919,N_2422);
nand U9548 (N_9548,N_2623,N_1797);
and U9549 (N_9549,N_1787,N_173);
nor U9550 (N_9550,N_1786,N_3529);
or U9551 (N_9551,N_5887,N_939);
nand U9552 (N_9552,N_1891,N_4658);
nor U9553 (N_9553,N_253,N_3197);
nand U9554 (N_9554,N_3584,N_4981);
and U9555 (N_9555,N_1811,N_1059);
xor U9556 (N_9556,N_3112,N_2431);
and U9557 (N_9557,N_4669,N_4928);
nor U9558 (N_9558,N_6243,N_3804);
xnor U9559 (N_9559,N_3756,N_2036);
nand U9560 (N_9560,N_596,N_1598);
nand U9561 (N_9561,N_1154,N_2213);
and U9562 (N_9562,N_1857,N_1337);
nand U9563 (N_9563,N_2675,N_928);
and U9564 (N_9564,N_2983,N_272);
xor U9565 (N_9565,N_3913,N_2187);
or U9566 (N_9566,N_4634,N_1766);
nor U9567 (N_9567,N_4295,N_2643);
xor U9568 (N_9568,N_1076,N_5202);
or U9569 (N_9569,N_4851,N_4068);
nand U9570 (N_9570,N_144,N_1761);
and U9571 (N_9571,N_2654,N_3379);
or U9572 (N_9572,N_228,N_3721);
or U9573 (N_9573,N_4386,N_435);
nor U9574 (N_9574,N_4381,N_1575);
nand U9575 (N_9575,N_277,N_6041);
nor U9576 (N_9576,N_2684,N_5739);
nor U9577 (N_9577,N_5076,N_1122);
nor U9578 (N_9578,N_4651,N_980);
or U9579 (N_9579,N_5252,N_4715);
or U9580 (N_9580,N_1584,N_3818);
nor U9581 (N_9581,N_2527,N_3609);
or U9582 (N_9582,N_2448,N_5470);
and U9583 (N_9583,N_3901,N_480);
xnor U9584 (N_9584,N_523,N_5186);
nor U9585 (N_9585,N_1915,N_679);
nand U9586 (N_9586,N_228,N_884);
or U9587 (N_9587,N_4541,N_3893);
nor U9588 (N_9588,N_2745,N_1157);
or U9589 (N_9589,N_5822,N_5336);
xnor U9590 (N_9590,N_3626,N_2204);
and U9591 (N_9591,N_4219,N_1138);
xnor U9592 (N_9592,N_85,N_5759);
xor U9593 (N_9593,N_1126,N_1358);
nor U9594 (N_9594,N_135,N_1079);
xor U9595 (N_9595,N_5613,N_2487);
nand U9596 (N_9596,N_3481,N_3293);
nand U9597 (N_9597,N_1821,N_1300);
or U9598 (N_9598,N_1067,N_2570);
nand U9599 (N_9599,N_2097,N_1063);
nor U9600 (N_9600,N_3291,N_1989);
nor U9601 (N_9601,N_2098,N_3512);
or U9602 (N_9602,N_6097,N_2415);
xor U9603 (N_9603,N_3440,N_6119);
or U9604 (N_9604,N_2167,N_4622);
nor U9605 (N_9605,N_1365,N_2765);
or U9606 (N_9606,N_1932,N_1940);
or U9607 (N_9607,N_1647,N_3985);
or U9608 (N_9608,N_1501,N_3068);
xor U9609 (N_9609,N_2966,N_3305);
xor U9610 (N_9610,N_3828,N_1449);
xor U9611 (N_9611,N_3586,N_5282);
nor U9612 (N_9612,N_2847,N_2541);
and U9613 (N_9613,N_2789,N_384);
and U9614 (N_9614,N_5150,N_5485);
nand U9615 (N_9615,N_2916,N_3297);
or U9616 (N_9616,N_2194,N_1391);
xnor U9617 (N_9617,N_5712,N_977);
and U9618 (N_9618,N_4072,N_1603);
nor U9619 (N_9619,N_2206,N_5659);
and U9620 (N_9620,N_4158,N_1083);
nor U9621 (N_9621,N_5700,N_5579);
or U9622 (N_9622,N_2486,N_4766);
or U9623 (N_9623,N_3689,N_4530);
and U9624 (N_9624,N_3195,N_1319);
nor U9625 (N_9625,N_753,N_940);
nor U9626 (N_9626,N_3498,N_14);
and U9627 (N_9627,N_1958,N_1156);
and U9628 (N_9628,N_1402,N_2946);
and U9629 (N_9629,N_1108,N_53);
and U9630 (N_9630,N_6001,N_5749);
nor U9631 (N_9631,N_177,N_4386);
or U9632 (N_9632,N_5610,N_1191);
xor U9633 (N_9633,N_1904,N_3316);
and U9634 (N_9634,N_5168,N_1097);
or U9635 (N_9635,N_5647,N_2553);
nor U9636 (N_9636,N_392,N_3492);
and U9637 (N_9637,N_2398,N_3689);
nor U9638 (N_9638,N_967,N_843);
and U9639 (N_9639,N_3630,N_4669);
or U9640 (N_9640,N_2057,N_5283);
and U9641 (N_9641,N_1296,N_1470);
and U9642 (N_9642,N_5696,N_2666);
xnor U9643 (N_9643,N_2339,N_5850);
nor U9644 (N_9644,N_6081,N_4212);
nor U9645 (N_9645,N_2497,N_2437);
xnor U9646 (N_9646,N_4835,N_5135);
nand U9647 (N_9647,N_5845,N_373);
nor U9648 (N_9648,N_3608,N_4933);
and U9649 (N_9649,N_4981,N_4215);
nand U9650 (N_9650,N_3117,N_2400);
xnor U9651 (N_9651,N_163,N_5335);
nor U9652 (N_9652,N_1339,N_1842);
and U9653 (N_9653,N_5407,N_2002);
and U9654 (N_9654,N_564,N_4479);
or U9655 (N_9655,N_1730,N_1450);
xor U9656 (N_9656,N_6133,N_5766);
or U9657 (N_9657,N_272,N_2881);
nor U9658 (N_9658,N_3233,N_2067);
nor U9659 (N_9659,N_685,N_319);
nor U9660 (N_9660,N_736,N_5406);
and U9661 (N_9661,N_3829,N_2974);
nor U9662 (N_9662,N_348,N_2993);
nor U9663 (N_9663,N_3742,N_1704);
and U9664 (N_9664,N_5717,N_833);
and U9665 (N_9665,N_3539,N_2199);
xor U9666 (N_9666,N_3792,N_1627);
nand U9667 (N_9667,N_693,N_1670);
nor U9668 (N_9668,N_2310,N_2756);
xnor U9669 (N_9669,N_5307,N_4113);
or U9670 (N_9670,N_2115,N_5612);
or U9671 (N_9671,N_4576,N_4823);
and U9672 (N_9672,N_449,N_4186);
nor U9673 (N_9673,N_744,N_1716);
xor U9674 (N_9674,N_1872,N_1624);
nand U9675 (N_9675,N_5551,N_463);
nand U9676 (N_9676,N_83,N_1409);
nor U9677 (N_9677,N_4656,N_443);
xnor U9678 (N_9678,N_2355,N_643);
xnor U9679 (N_9679,N_4609,N_5448);
or U9680 (N_9680,N_5437,N_1465);
nand U9681 (N_9681,N_3176,N_2044);
xnor U9682 (N_9682,N_5887,N_641);
xnor U9683 (N_9683,N_4771,N_2941);
xnor U9684 (N_9684,N_587,N_5774);
and U9685 (N_9685,N_2929,N_5664);
xor U9686 (N_9686,N_5464,N_5087);
and U9687 (N_9687,N_5852,N_4488);
or U9688 (N_9688,N_3530,N_6238);
xnor U9689 (N_9689,N_4328,N_1478);
xor U9690 (N_9690,N_5202,N_2413);
nand U9691 (N_9691,N_2540,N_307);
or U9692 (N_9692,N_6130,N_537);
and U9693 (N_9693,N_4537,N_59);
and U9694 (N_9694,N_3611,N_4696);
nor U9695 (N_9695,N_3822,N_5949);
xnor U9696 (N_9696,N_3288,N_5961);
xnor U9697 (N_9697,N_5689,N_5596);
nor U9698 (N_9698,N_190,N_2915);
and U9699 (N_9699,N_5419,N_3388);
and U9700 (N_9700,N_3982,N_3788);
or U9701 (N_9701,N_3735,N_3201);
nand U9702 (N_9702,N_4410,N_2539);
nor U9703 (N_9703,N_735,N_1730);
or U9704 (N_9704,N_6084,N_1614);
xor U9705 (N_9705,N_2899,N_1848);
nor U9706 (N_9706,N_5321,N_5490);
and U9707 (N_9707,N_5655,N_4832);
and U9708 (N_9708,N_1528,N_2866);
and U9709 (N_9709,N_436,N_3820);
or U9710 (N_9710,N_6115,N_642);
or U9711 (N_9711,N_1745,N_5985);
xnor U9712 (N_9712,N_5847,N_239);
and U9713 (N_9713,N_472,N_4886);
nor U9714 (N_9714,N_3196,N_4847);
nand U9715 (N_9715,N_2093,N_280);
or U9716 (N_9716,N_3009,N_5431);
nor U9717 (N_9717,N_2514,N_3918);
or U9718 (N_9718,N_2337,N_1684);
and U9719 (N_9719,N_3737,N_5385);
xor U9720 (N_9720,N_6039,N_1912);
xor U9721 (N_9721,N_596,N_1941);
and U9722 (N_9722,N_236,N_2195);
and U9723 (N_9723,N_4610,N_2577);
nor U9724 (N_9724,N_3813,N_6086);
nand U9725 (N_9725,N_3147,N_3064);
nor U9726 (N_9726,N_4193,N_4234);
nor U9727 (N_9727,N_90,N_5325);
xnor U9728 (N_9728,N_4108,N_6162);
and U9729 (N_9729,N_6159,N_1402);
xor U9730 (N_9730,N_3310,N_3434);
nand U9731 (N_9731,N_651,N_5097);
nand U9732 (N_9732,N_4619,N_4609);
nor U9733 (N_9733,N_3912,N_3469);
and U9734 (N_9734,N_4174,N_905);
xnor U9735 (N_9735,N_4615,N_4026);
nor U9736 (N_9736,N_1616,N_2655);
nor U9737 (N_9737,N_1865,N_5704);
or U9738 (N_9738,N_2249,N_2996);
nor U9739 (N_9739,N_1247,N_5242);
xnor U9740 (N_9740,N_686,N_1741);
nand U9741 (N_9741,N_5252,N_2365);
nor U9742 (N_9742,N_2550,N_5528);
nand U9743 (N_9743,N_1100,N_1812);
and U9744 (N_9744,N_6017,N_3514);
nand U9745 (N_9745,N_1453,N_2817);
nor U9746 (N_9746,N_2598,N_6140);
nor U9747 (N_9747,N_3456,N_3647);
nor U9748 (N_9748,N_314,N_4837);
nor U9749 (N_9749,N_6022,N_374);
or U9750 (N_9750,N_5604,N_4679);
nor U9751 (N_9751,N_2846,N_4838);
or U9752 (N_9752,N_2546,N_3244);
or U9753 (N_9753,N_3014,N_2396);
nand U9754 (N_9754,N_5066,N_3686);
and U9755 (N_9755,N_3280,N_99);
or U9756 (N_9756,N_3114,N_3000);
xor U9757 (N_9757,N_5791,N_5258);
xor U9758 (N_9758,N_2878,N_1707);
or U9759 (N_9759,N_1707,N_5401);
xnor U9760 (N_9760,N_55,N_4946);
and U9761 (N_9761,N_3779,N_5585);
nor U9762 (N_9762,N_2241,N_5200);
nor U9763 (N_9763,N_5461,N_1020);
nand U9764 (N_9764,N_5000,N_1421);
or U9765 (N_9765,N_3085,N_2037);
nor U9766 (N_9766,N_5938,N_3989);
xnor U9767 (N_9767,N_5050,N_1099);
and U9768 (N_9768,N_2189,N_2938);
or U9769 (N_9769,N_5868,N_4277);
nand U9770 (N_9770,N_104,N_5090);
or U9771 (N_9771,N_5384,N_2711);
nand U9772 (N_9772,N_2688,N_5542);
nand U9773 (N_9773,N_500,N_2384);
and U9774 (N_9774,N_5302,N_3429);
nand U9775 (N_9775,N_1747,N_3757);
nor U9776 (N_9776,N_5175,N_4150);
xor U9777 (N_9777,N_2364,N_4655);
or U9778 (N_9778,N_3852,N_5194);
and U9779 (N_9779,N_409,N_5444);
xor U9780 (N_9780,N_2239,N_5630);
xor U9781 (N_9781,N_226,N_4323);
and U9782 (N_9782,N_1815,N_1244);
nor U9783 (N_9783,N_3301,N_6000);
or U9784 (N_9784,N_1907,N_1414);
nor U9785 (N_9785,N_2216,N_2349);
or U9786 (N_9786,N_1416,N_3797);
nand U9787 (N_9787,N_473,N_3846);
xnor U9788 (N_9788,N_4033,N_3446);
xor U9789 (N_9789,N_1718,N_1353);
nor U9790 (N_9790,N_3666,N_11);
and U9791 (N_9791,N_2602,N_5938);
or U9792 (N_9792,N_5341,N_2839);
and U9793 (N_9793,N_596,N_2531);
nand U9794 (N_9794,N_1613,N_1868);
xnor U9795 (N_9795,N_5852,N_2787);
or U9796 (N_9796,N_5608,N_3403);
and U9797 (N_9797,N_3985,N_6131);
or U9798 (N_9798,N_4621,N_2911);
and U9799 (N_9799,N_4433,N_2376);
xor U9800 (N_9800,N_6206,N_5389);
xor U9801 (N_9801,N_5737,N_3616);
nand U9802 (N_9802,N_5122,N_2256);
and U9803 (N_9803,N_5295,N_5677);
nor U9804 (N_9804,N_2329,N_2224);
nor U9805 (N_9805,N_181,N_4326);
or U9806 (N_9806,N_2581,N_4872);
and U9807 (N_9807,N_3033,N_3699);
xnor U9808 (N_9808,N_1957,N_5632);
and U9809 (N_9809,N_5238,N_5666);
xnor U9810 (N_9810,N_3048,N_5464);
nand U9811 (N_9811,N_2346,N_2527);
nand U9812 (N_9812,N_4031,N_5432);
nand U9813 (N_9813,N_820,N_3497);
or U9814 (N_9814,N_1885,N_1901);
nand U9815 (N_9815,N_4812,N_6214);
or U9816 (N_9816,N_140,N_2997);
nand U9817 (N_9817,N_6086,N_5819);
nand U9818 (N_9818,N_4666,N_4556);
nand U9819 (N_9819,N_4287,N_1781);
nor U9820 (N_9820,N_5106,N_228);
nand U9821 (N_9821,N_3619,N_5752);
xor U9822 (N_9822,N_2007,N_2838);
and U9823 (N_9823,N_317,N_4392);
and U9824 (N_9824,N_3719,N_5452);
nand U9825 (N_9825,N_1431,N_5601);
xor U9826 (N_9826,N_568,N_812);
nand U9827 (N_9827,N_4071,N_4965);
nand U9828 (N_9828,N_1480,N_772);
and U9829 (N_9829,N_5182,N_5472);
nor U9830 (N_9830,N_5587,N_1441);
or U9831 (N_9831,N_3649,N_4412);
nor U9832 (N_9832,N_6067,N_4017);
nor U9833 (N_9833,N_1401,N_5219);
or U9834 (N_9834,N_410,N_3518);
xnor U9835 (N_9835,N_3173,N_3910);
and U9836 (N_9836,N_3107,N_3361);
nand U9837 (N_9837,N_2439,N_121);
and U9838 (N_9838,N_2659,N_272);
and U9839 (N_9839,N_2322,N_417);
xor U9840 (N_9840,N_5783,N_2537);
and U9841 (N_9841,N_6213,N_1318);
or U9842 (N_9842,N_1653,N_3811);
xor U9843 (N_9843,N_4052,N_5059);
nand U9844 (N_9844,N_482,N_5046);
nor U9845 (N_9845,N_5646,N_2518);
or U9846 (N_9846,N_3044,N_1090);
and U9847 (N_9847,N_719,N_1527);
nor U9848 (N_9848,N_2968,N_1563);
and U9849 (N_9849,N_2852,N_1935);
nor U9850 (N_9850,N_5060,N_5507);
xor U9851 (N_9851,N_1388,N_3489);
or U9852 (N_9852,N_2002,N_3045);
nor U9853 (N_9853,N_5969,N_2540);
nand U9854 (N_9854,N_4963,N_273);
or U9855 (N_9855,N_3580,N_4209);
nor U9856 (N_9856,N_2284,N_4874);
nand U9857 (N_9857,N_661,N_2874);
and U9858 (N_9858,N_3752,N_4465);
xor U9859 (N_9859,N_2215,N_662);
or U9860 (N_9860,N_504,N_5247);
nor U9861 (N_9861,N_3168,N_844);
or U9862 (N_9862,N_1106,N_2544);
xnor U9863 (N_9863,N_1461,N_2790);
and U9864 (N_9864,N_1772,N_2329);
xor U9865 (N_9865,N_4648,N_5617);
nand U9866 (N_9866,N_1752,N_3181);
and U9867 (N_9867,N_4393,N_2196);
or U9868 (N_9868,N_1981,N_3730);
xnor U9869 (N_9869,N_3739,N_2533);
or U9870 (N_9870,N_807,N_1682);
nand U9871 (N_9871,N_4096,N_1906);
nor U9872 (N_9872,N_3169,N_5855);
or U9873 (N_9873,N_2791,N_4834);
nand U9874 (N_9874,N_3997,N_1648);
or U9875 (N_9875,N_3346,N_1333);
and U9876 (N_9876,N_4326,N_2265);
or U9877 (N_9877,N_1942,N_6070);
nor U9878 (N_9878,N_4595,N_5017);
xor U9879 (N_9879,N_4877,N_4096);
and U9880 (N_9880,N_80,N_5607);
nor U9881 (N_9881,N_774,N_2375);
nor U9882 (N_9882,N_1621,N_1354);
or U9883 (N_9883,N_1050,N_615);
and U9884 (N_9884,N_5729,N_3059);
and U9885 (N_9885,N_2588,N_4684);
or U9886 (N_9886,N_3496,N_4945);
xor U9887 (N_9887,N_3933,N_145);
nand U9888 (N_9888,N_4114,N_5851);
xor U9889 (N_9889,N_3193,N_4561);
nand U9890 (N_9890,N_4599,N_4212);
or U9891 (N_9891,N_5813,N_3016);
xor U9892 (N_9892,N_1488,N_844);
nor U9893 (N_9893,N_1601,N_2819);
or U9894 (N_9894,N_5386,N_5408);
nand U9895 (N_9895,N_4378,N_5302);
or U9896 (N_9896,N_3046,N_3527);
and U9897 (N_9897,N_3293,N_2891);
xor U9898 (N_9898,N_3152,N_2054);
nor U9899 (N_9899,N_4895,N_3326);
nor U9900 (N_9900,N_1635,N_2440);
nand U9901 (N_9901,N_4602,N_4332);
nand U9902 (N_9902,N_5492,N_4480);
or U9903 (N_9903,N_516,N_4615);
and U9904 (N_9904,N_661,N_4009);
nand U9905 (N_9905,N_3766,N_4220);
nand U9906 (N_9906,N_5808,N_3517);
nor U9907 (N_9907,N_3993,N_1497);
nor U9908 (N_9908,N_556,N_1937);
nor U9909 (N_9909,N_5591,N_4566);
or U9910 (N_9910,N_4153,N_982);
and U9911 (N_9911,N_491,N_650);
nor U9912 (N_9912,N_2545,N_3564);
nor U9913 (N_9913,N_3042,N_3261);
nand U9914 (N_9914,N_3046,N_3161);
xnor U9915 (N_9915,N_997,N_449);
and U9916 (N_9916,N_4570,N_3295);
nand U9917 (N_9917,N_5454,N_1388);
nand U9918 (N_9918,N_2267,N_5720);
nor U9919 (N_9919,N_552,N_3907);
nand U9920 (N_9920,N_507,N_1111);
or U9921 (N_9921,N_4515,N_5764);
and U9922 (N_9922,N_1718,N_3766);
or U9923 (N_9923,N_5848,N_5572);
nand U9924 (N_9924,N_2472,N_5310);
xnor U9925 (N_9925,N_810,N_3459);
xor U9926 (N_9926,N_3976,N_2330);
xnor U9927 (N_9927,N_14,N_4791);
and U9928 (N_9928,N_2636,N_989);
and U9929 (N_9929,N_6080,N_3061);
or U9930 (N_9930,N_117,N_1718);
and U9931 (N_9931,N_1578,N_4904);
nor U9932 (N_9932,N_3599,N_1395);
or U9933 (N_9933,N_5704,N_1790);
nand U9934 (N_9934,N_6008,N_182);
and U9935 (N_9935,N_1243,N_4736);
and U9936 (N_9936,N_1078,N_456);
and U9937 (N_9937,N_659,N_1236);
and U9938 (N_9938,N_409,N_4942);
nand U9939 (N_9939,N_1002,N_5059);
nand U9940 (N_9940,N_2086,N_3266);
and U9941 (N_9941,N_2996,N_3825);
nand U9942 (N_9942,N_686,N_4665);
and U9943 (N_9943,N_2039,N_2395);
nand U9944 (N_9944,N_2567,N_5654);
and U9945 (N_9945,N_5107,N_4182);
xor U9946 (N_9946,N_1947,N_753);
and U9947 (N_9947,N_3988,N_477);
nand U9948 (N_9948,N_215,N_965);
or U9949 (N_9949,N_5701,N_846);
nand U9950 (N_9950,N_2063,N_5232);
nor U9951 (N_9951,N_1151,N_1870);
xor U9952 (N_9952,N_3759,N_4754);
xor U9953 (N_9953,N_1641,N_2755);
and U9954 (N_9954,N_6029,N_3404);
and U9955 (N_9955,N_1794,N_5597);
and U9956 (N_9956,N_2853,N_4371);
nand U9957 (N_9957,N_1670,N_3551);
nor U9958 (N_9958,N_3631,N_2556);
xnor U9959 (N_9959,N_4729,N_171);
nand U9960 (N_9960,N_1216,N_2404);
or U9961 (N_9961,N_5826,N_3457);
nor U9962 (N_9962,N_2894,N_3953);
and U9963 (N_9963,N_170,N_943);
and U9964 (N_9964,N_6199,N_4026);
and U9965 (N_9965,N_1651,N_5890);
nand U9966 (N_9966,N_242,N_1680);
or U9967 (N_9967,N_4332,N_2172);
nand U9968 (N_9968,N_541,N_4954);
nor U9969 (N_9969,N_5727,N_1966);
and U9970 (N_9970,N_1608,N_1021);
or U9971 (N_9971,N_2299,N_5892);
nand U9972 (N_9972,N_1987,N_4694);
or U9973 (N_9973,N_270,N_1794);
nand U9974 (N_9974,N_2154,N_4617);
xnor U9975 (N_9975,N_469,N_3747);
and U9976 (N_9976,N_338,N_5714);
or U9977 (N_9977,N_5964,N_2894);
or U9978 (N_9978,N_1974,N_2300);
nor U9979 (N_9979,N_5488,N_2973);
nor U9980 (N_9980,N_3301,N_4405);
and U9981 (N_9981,N_2733,N_46);
or U9982 (N_9982,N_5475,N_4488);
nor U9983 (N_9983,N_4324,N_2462);
nor U9984 (N_9984,N_1922,N_1738);
xor U9985 (N_9985,N_2384,N_125);
or U9986 (N_9986,N_2527,N_26);
nor U9987 (N_9987,N_3978,N_3765);
nor U9988 (N_9988,N_4449,N_5789);
nor U9989 (N_9989,N_1742,N_6246);
xor U9990 (N_9990,N_4030,N_2820);
and U9991 (N_9991,N_4951,N_4235);
or U9992 (N_9992,N_288,N_5654);
xor U9993 (N_9993,N_4092,N_5600);
nand U9994 (N_9994,N_3213,N_2950);
xnor U9995 (N_9995,N_1319,N_483);
nor U9996 (N_9996,N_5002,N_3881);
and U9997 (N_9997,N_4389,N_4022);
nand U9998 (N_9998,N_4389,N_1440);
xor U9999 (N_9999,N_2909,N_2328);
nand U10000 (N_10000,N_1134,N_342);
nand U10001 (N_10001,N_4007,N_2191);
nand U10002 (N_10002,N_3331,N_2494);
xnor U10003 (N_10003,N_4747,N_5241);
nor U10004 (N_10004,N_3158,N_2082);
or U10005 (N_10005,N_3234,N_2174);
nand U10006 (N_10006,N_4653,N_52);
nor U10007 (N_10007,N_1067,N_4250);
nand U10008 (N_10008,N_556,N_1527);
and U10009 (N_10009,N_3850,N_3880);
or U10010 (N_10010,N_2003,N_4978);
xnor U10011 (N_10011,N_4031,N_1435);
and U10012 (N_10012,N_3793,N_3460);
xnor U10013 (N_10013,N_5877,N_4572);
xnor U10014 (N_10014,N_1530,N_3992);
and U10015 (N_10015,N_370,N_1312);
nand U10016 (N_10016,N_4471,N_1971);
xor U10017 (N_10017,N_1009,N_3846);
or U10018 (N_10018,N_2882,N_3620);
nor U10019 (N_10019,N_5175,N_1576);
xor U10020 (N_10020,N_3061,N_1740);
nand U10021 (N_10021,N_516,N_3160);
nor U10022 (N_10022,N_4495,N_4695);
or U10023 (N_10023,N_66,N_5706);
nor U10024 (N_10024,N_2062,N_802);
and U10025 (N_10025,N_6155,N_3542);
nor U10026 (N_10026,N_4788,N_2800);
xnor U10027 (N_10027,N_5741,N_3401);
nand U10028 (N_10028,N_6080,N_1294);
nand U10029 (N_10029,N_744,N_4146);
nor U10030 (N_10030,N_5826,N_1843);
xor U10031 (N_10031,N_2238,N_5299);
nand U10032 (N_10032,N_72,N_3623);
or U10033 (N_10033,N_4841,N_2255);
xnor U10034 (N_10034,N_5476,N_286);
or U10035 (N_10035,N_2783,N_4106);
and U10036 (N_10036,N_562,N_1279);
or U10037 (N_10037,N_6161,N_2097);
nor U10038 (N_10038,N_1413,N_3898);
nor U10039 (N_10039,N_1779,N_4203);
or U10040 (N_10040,N_2182,N_2154);
or U10041 (N_10041,N_4247,N_2514);
nor U10042 (N_10042,N_5289,N_4048);
or U10043 (N_10043,N_1578,N_4152);
and U10044 (N_10044,N_258,N_4670);
or U10045 (N_10045,N_685,N_6212);
nand U10046 (N_10046,N_5053,N_3243);
and U10047 (N_10047,N_1687,N_4288);
and U10048 (N_10048,N_3380,N_3778);
nand U10049 (N_10049,N_4118,N_2983);
xnor U10050 (N_10050,N_3020,N_5979);
nor U10051 (N_10051,N_3787,N_2734);
and U10052 (N_10052,N_4675,N_3284);
nand U10053 (N_10053,N_4481,N_744);
and U10054 (N_10054,N_1799,N_1138);
nor U10055 (N_10055,N_3020,N_3779);
and U10056 (N_10056,N_4150,N_4088);
xor U10057 (N_10057,N_1018,N_2994);
or U10058 (N_10058,N_5713,N_3615);
and U10059 (N_10059,N_2885,N_2020);
xor U10060 (N_10060,N_5449,N_5504);
xor U10061 (N_10061,N_1110,N_869);
nor U10062 (N_10062,N_4653,N_4595);
or U10063 (N_10063,N_979,N_3703);
nor U10064 (N_10064,N_1875,N_4363);
nand U10065 (N_10065,N_553,N_4659);
nor U10066 (N_10066,N_5881,N_562);
or U10067 (N_10067,N_3227,N_1842);
xor U10068 (N_10068,N_224,N_3436);
nor U10069 (N_10069,N_2435,N_5357);
xor U10070 (N_10070,N_997,N_2300);
nand U10071 (N_10071,N_1951,N_1731);
nor U10072 (N_10072,N_6110,N_881);
xor U10073 (N_10073,N_5112,N_6152);
or U10074 (N_10074,N_2156,N_6244);
xor U10075 (N_10075,N_6228,N_2143);
xor U10076 (N_10076,N_4757,N_3746);
and U10077 (N_10077,N_3483,N_3636);
nor U10078 (N_10078,N_2197,N_3208);
nand U10079 (N_10079,N_5089,N_5444);
xnor U10080 (N_10080,N_1306,N_2564);
nor U10081 (N_10081,N_5921,N_2975);
nor U10082 (N_10082,N_5883,N_653);
nor U10083 (N_10083,N_1351,N_2380);
xnor U10084 (N_10084,N_2186,N_5342);
or U10085 (N_10085,N_1144,N_3863);
and U10086 (N_10086,N_5945,N_1870);
and U10087 (N_10087,N_140,N_2330);
nand U10088 (N_10088,N_3786,N_3584);
and U10089 (N_10089,N_3973,N_5279);
nand U10090 (N_10090,N_4780,N_4064);
and U10091 (N_10091,N_4746,N_3494);
and U10092 (N_10092,N_2539,N_4202);
or U10093 (N_10093,N_3263,N_875);
and U10094 (N_10094,N_3892,N_3727);
or U10095 (N_10095,N_5670,N_3952);
and U10096 (N_10096,N_2708,N_4611);
or U10097 (N_10097,N_5245,N_962);
or U10098 (N_10098,N_51,N_6128);
nand U10099 (N_10099,N_1248,N_3662);
xnor U10100 (N_10100,N_3383,N_251);
nand U10101 (N_10101,N_2193,N_4502);
xor U10102 (N_10102,N_563,N_2979);
and U10103 (N_10103,N_589,N_3920);
and U10104 (N_10104,N_5922,N_3351);
nor U10105 (N_10105,N_509,N_3033);
or U10106 (N_10106,N_594,N_75);
nor U10107 (N_10107,N_3014,N_1769);
nand U10108 (N_10108,N_1139,N_3670);
nand U10109 (N_10109,N_2976,N_4549);
nand U10110 (N_10110,N_5828,N_4777);
and U10111 (N_10111,N_1328,N_838);
xnor U10112 (N_10112,N_5431,N_5637);
and U10113 (N_10113,N_2850,N_515);
nor U10114 (N_10114,N_4394,N_6059);
and U10115 (N_10115,N_650,N_5306);
and U10116 (N_10116,N_6035,N_3103);
or U10117 (N_10117,N_4621,N_853);
nor U10118 (N_10118,N_3534,N_5347);
or U10119 (N_10119,N_1079,N_2239);
nand U10120 (N_10120,N_1541,N_3351);
or U10121 (N_10121,N_1101,N_5862);
nand U10122 (N_10122,N_2887,N_2809);
xor U10123 (N_10123,N_5265,N_3344);
xnor U10124 (N_10124,N_5289,N_5549);
or U10125 (N_10125,N_3433,N_2796);
or U10126 (N_10126,N_5909,N_506);
or U10127 (N_10127,N_2199,N_627);
nand U10128 (N_10128,N_3513,N_2550);
and U10129 (N_10129,N_3187,N_4172);
nor U10130 (N_10130,N_1209,N_1571);
nand U10131 (N_10131,N_2154,N_766);
nor U10132 (N_10132,N_275,N_6100);
nand U10133 (N_10133,N_5228,N_2624);
xnor U10134 (N_10134,N_3161,N_664);
nand U10135 (N_10135,N_1094,N_4801);
and U10136 (N_10136,N_2989,N_1354);
nor U10137 (N_10137,N_2987,N_3241);
and U10138 (N_10138,N_2360,N_680);
or U10139 (N_10139,N_4532,N_2519);
nor U10140 (N_10140,N_391,N_4683);
nand U10141 (N_10141,N_1462,N_1269);
xnor U10142 (N_10142,N_2637,N_2567);
nor U10143 (N_10143,N_3418,N_1091);
or U10144 (N_10144,N_3546,N_3171);
nor U10145 (N_10145,N_470,N_2264);
nor U10146 (N_10146,N_3513,N_1849);
and U10147 (N_10147,N_1932,N_2480);
nor U10148 (N_10148,N_925,N_1577);
nor U10149 (N_10149,N_5303,N_3021);
and U10150 (N_10150,N_2208,N_271);
xnor U10151 (N_10151,N_2443,N_252);
and U10152 (N_10152,N_5216,N_842);
nand U10153 (N_10153,N_3908,N_3229);
and U10154 (N_10154,N_1013,N_6048);
and U10155 (N_10155,N_1824,N_4348);
and U10156 (N_10156,N_6106,N_2942);
and U10157 (N_10157,N_3320,N_4884);
or U10158 (N_10158,N_3405,N_3209);
or U10159 (N_10159,N_4464,N_4258);
xor U10160 (N_10160,N_2095,N_4913);
nand U10161 (N_10161,N_2005,N_32);
and U10162 (N_10162,N_489,N_2352);
nand U10163 (N_10163,N_4048,N_653);
and U10164 (N_10164,N_798,N_892);
nor U10165 (N_10165,N_744,N_2467);
nor U10166 (N_10166,N_2247,N_618);
xor U10167 (N_10167,N_2297,N_3744);
and U10168 (N_10168,N_2574,N_3361);
nand U10169 (N_10169,N_1130,N_2722);
nand U10170 (N_10170,N_4299,N_3426);
or U10171 (N_10171,N_1840,N_1056);
or U10172 (N_10172,N_1850,N_3692);
xnor U10173 (N_10173,N_3755,N_5916);
or U10174 (N_10174,N_2423,N_4309);
nor U10175 (N_10175,N_3466,N_4406);
nand U10176 (N_10176,N_3098,N_4259);
nand U10177 (N_10177,N_3400,N_2010);
xor U10178 (N_10178,N_5670,N_4364);
or U10179 (N_10179,N_2392,N_2965);
xnor U10180 (N_10180,N_2794,N_3042);
and U10181 (N_10181,N_2823,N_637);
nand U10182 (N_10182,N_3198,N_4855);
xnor U10183 (N_10183,N_1355,N_3613);
nor U10184 (N_10184,N_5088,N_1872);
nand U10185 (N_10185,N_1007,N_1321);
nor U10186 (N_10186,N_956,N_2740);
nand U10187 (N_10187,N_1640,N_4649);
nand U10188 (N_10188,N_1300,N_1207);
nor U10189 (N_10189,N_3117,N_4266);
and U10190 (N_10190,N_4302,N_5728);
and U10191 (N_10191,N_146,N_2231);
and U10192 (N_10192,N_3625,N_3348);
nor U10193 (N_10193,N_3211,N_4112);
or U10194 (N_10194,N_2990,N_2613);
and U10195 (N_10195,N_720,N_2253);
nand U10196 (N_10196,N_1957,N_2984);
and U10197 (N_10197,N_404,N_6182);
xnor U10198 (N_10198,N_2527,N_1987);
or U10199 (N_10199,N_3304,N_394);
or U10200 (N_10200,N_471,N_6);
xor U10201 (N_10201,N_5233,N_3612);
xor U10202 (N_10202,N_1850,N_3503);
nand U10203 (N_10203,N_3298,N_2623);
nor U10204 (N_10204,N_3447,N_1562);
xnor U10205 (N_10205,N_2062,N_4594);
nor U10206 (N_10206,N_1632,N_509);
nand U10207 (N_10207,N_696,N_1089);
xnor U10208 (N_10208,N_4273,N_2370);
or U10209 (N_10209,N_1906,N_1218);
xor U10210 (N_10210,N_819,N_4167);
nand U10211 (N_10211,N_4251,N_940);
and U10212 (N_10212,N_1218,N_3696);
nand U10213 (N_10213,N_437,N_720);
and U10214 (N_10214,N_538,N_776);
or U10215 (N_10215,N_1083,N_1542);
or U10216 (N_10216,N_431,N_3122);
nand U10217 (N_10217,N_3102,N_1965);
nand U10218 (N_10218,N_2997,N_5310);
nor U10219 (N_10219,N_4659,N_1239);
or U10220 (N_10220,N_3385,N_3975);
nand U10221 (N_10221,N_2716,N_2961);
and U10222 (N_10222,N_885,N_2782);
nor U10223 (N_10223,N_3647,N_5214);
nand U10224 (N_10224,N_4772,N_690);
xor U10225 (N_10225,N_3200,N_5980);
or U10226 (N_10226,N_5391,N_3294);
and U10227 (N_10227,N_2085,N_4308);
nand U10228 (N_10228,N_5246,N_4993);
or U10229 (N_10229,N_4362,N_1124);
nor U10230 (N_10230,N_1348,N_175);
nand U10231 (N_10231,N_1337,N_6175);
xnor U10232 (N_10232,N_1155,N_1060);
or U10233 (N_10233,N_992,N_4061);
or U10234 (N_10234,N_3818,N_1444);
and U10235 (N_10235,N_5393,N_2043);
and U10236 (N_10236,N_2612,N_1729);
nor U10237 (N_10237,N_1481,N_6221);
xor U10238 (N_10238,N_4343,N_2763);
nand U10239 (N_10239,N_4403,N_5639);
or U10240 (N_10240,N_2960,N_3504);
xnor U10241 (N_10241,N_910,N_530);
nor U10242 (N_10242,N_3322,N_3061);
nand U10243 (N_10243,N_2573,N_1648);
xor U10244 (N_10244,N_4878,N_2524);
xor U10245 (N_10245,N_1598,N_3605);
or U10246 (N_10246,N_6064,N_5998);
or U10247 (N_10247,N_4246,N_1873);
nand U10248 (N_10248,N_882,N_1533);
nand U10249 (N_10249,N_3400,N_4315);
nand U10250 (N_10250,N_2450,N_2693);
or U10251 (N_10251,N_6151,N_3992);
nand U10252 (N_10252,N_464,N_4828);
and U10253 (N_10253,N_2119,N_1685);
or U10254 (N_10254,N_4505,N_4732);
and U10255 (N_10255,N_3913,N_3039);
xnor U10256 (N_10256,N_4228,N_1862);
xor U10257 (N_10257,N_2376,N_4462);
nand U10258 (N_10258,N_3257,N_625);
nand U10259 (N_10259,N_348,N_4097);
nor U10260 (N_10260,N_3246,N_5930);
nor U10261 (N_10261,N_3432,N_1866);
nor U10262 (N_10262,N_645,N_1747);
and U10263 (N_10263,N_5705,N_3776);
nor U10264 (N_10264,N_3973,N_1919);
or U10265 (N_10265,N_2939,N_1542);
nor U10266 (N_10266,N_2268,N_4699);
nand U10267 (N_10267,N_4994,N_4303);
nand U10268 (N_10268,N_2373,N_4601);
nor U10269 (N_10269,N_5050,N_5036);
nor U10270 (N_10270,N_4259,N_5377);
xnor U10271 (N_10271,N_700,N_5280);
xnor U10272 (N_10272,N_2248,N_626);
or U10273 (N_10273,N_3236,N_931);
or U10274 (N_10274,N_1854,N_2288);
nand U10275 (N_10275,N_701,N_753);
nand U10276 (N_10276,N_809,N_2173);
nand U10277 (N_10277,N_4534,N_4209);
and U10278 (N_10278,N_2679,N_3193);
or U10279 (N_10279,N_356,N_2845);
nor U10280 (N_10280,N_5970,N_5177);
or U10281 (N_10281,N_4957,N_985);
or U10282 (N_10282,N_1423,N_6070);
xnor U10283 (N_10283,N_4764,N_4076);
and U10284 (N_10284,N_2168,N_12);
or U10285 (N_10285,N_3111,N_4471);
xnor U10286 (N_10286,N_4928,N_2256);
and U10287 (N_10287,N_4460,N_5529);
nor U10288 (N_10288,N_5279,N_3219);
and U10289 (N_10289,N_1024,N_2957);
xnor U10290 (N_10290,N_1922,N_1446);
nor U10291 (N_10291,N_5563,N_1991);
xor U10292 (N_10292,N_4993,N_2886);
nand U10293 (N_10293,N_3407,N_2309);
xor U10294 (N_10294,N_1484,N_1357);
or U10295 (N_10295,N_2783,N_2213);
or U10296 (N_10296,N_1110,N_4799);
and U10297 (N_10297,N_2044,N_1389);
xnor U10298 (N_10298,N_1695,N_2129);
nand U10299 (N_10299,N_1877,N_99);
nor U10300 (N_10300,N_4443,N_557);
xor U10301 (N_10301,N_3255,N_5024);
and U10302 (N_10302,N_33,N_1454);
nor U10303 (N_10303,N_56,N_462);
xnor U10304 (N_10304,N_4322,N_62);
or U10305 (N_10305,N_4425,N_5941);
nand U10306 (N_10306,N_2137,N_3304);
or U10307 (N_10307,N_4242,N_2552);
or U10308 (N_10308,N_3661,N_234);
and U10309 (N_10309,N_2228,N_4720);
xor U10310 (N_10310,N_5951,N_774);
nand U10311 (N_10311,N_5043,N_1889);
and U10312 (N_10312,N_2881,N_3916);
nand U10313 (N_10313,N_3087,N_3941);
nand U10314 (N_10314,N_5447,N_4996);
or U10315 (N_10315,N_5547,N_328);
nand U10316 (N_10316,N_267,N_4514);
nand U10317 (N_10317,N_389,N_4357);
or U10318 (N_10318,N_3884,N_3340);
nor U10319 (N_10319,N_1201,N_3309);
nand U10320 (N_10320,N_419,N_6038);
or U10321 (N_10321,N_4965,N_354);
nor U10322 (N_10322,N_2529,N_2317);
nand U10323 (N_10323,N_1825,N_2454);
xnor U10324 (N_10324,N_1472,N_4417);
nand U10325 (N_10325,N_5288,N_340);
xor U10326 (N_10326,N_3179,N_2318);
nor U10327 (N_10327,N_3828,N_4717);
nand U10328 (N_10328,N_5364,N_4457);
nand U10329 (N_10329,N_1841,N_2416);
or U10330 (N_10330,N_4704,N_4994);
xnor U10331 (N_10331,N_6133,N_1461);
nor U10332 (N_10332,N_5538,N_4592);
xor U10333 (N_10333,N_5723,N_2696);
and U10334 (N_10334,N_6152,N_3501);
nor U10335 (N_10335,N_1097,N_1417);
nand U10336 (N_10336,N_511,N_1739);
and U10337 (N_10337,N_4202,N_5551);
xnor U10338 (N_10338,N_3638,N_3659);
nor U10339 (N_10339,N_5238,N_1265);
nand U10340 (N_10340,N_3263,N_3171);
nand U10341 (N_10341,N_4573,N_3904);
xnor U10342 (N_10342,N_3268,N_1301);
nor U10343 (N_10343,N_5599,N_5423);
or U10344 (N_10344,N_96,N_3678);
nor U10345 (N_10345,N_2838,N_4821);
nor U10346 (N_10346,N_5667,N_110);
nand U10347 (N_10347,N_1303,N_5501);
nand U10348 (N_10348,N_3930,N_694);
nor U10349 (N_10349,N_5661,N_5906);
nor U10350 (N_10350,N_1395,N_4604);
and U10351 (N_10351,N_408,N_3075);
nor U10352 (N_10352,N_3388,N_5200);
or U10353 (N_10353,N_5734,N_4101);
nand U10354 (N_10354,N_1343,N_4298);
or U10355 (N_10355,N_2766,N_3238);
xnor U10356 (N_10356,N_3299,N_1754);
xnor U10357 (N_10357,N_1174,N_1192);
nor U10358 (N_10358,N_5994,N_2155);
nor U10359 (N_10359,N_4739,N_2314);
nand U10360 (N_10360,N_3301,N_1415);
or U10361 (N_10361,N_5943,N_5565);
and U10362 (N_10362,N_5317,N_348);
and U10363 (N_10363,N_678,N_1205);
nor U10364 (N_10364,N_1027,N_2471);
nand U10365 (N_10365,N_4028,N_3344);
or U10366 (N_10366,N_1671,N_2105);
or U10367 (N_10367,N_3023,N_670);
xnor U10368 (N_10368,N_4165,N_3694);
and U10369 (N_10369,N_5390,N_5308);
xor U10370 (N_10370,N_690,N_2057);
or U10371 (N_10371,N_295,N_1909);
xnor U10372 (N_10372,N_5551,N_508);
xor U10373 (N_10373,N_968,N_2810);
or U10374 (N_10374,N_5338,N_1056);
or U10375 (N_10375,N_5903,N_6098);
and U10376 (N_10376,N_3530,N_3404);
nand U10377 (N_10377,N_3727,N_4455);
xnor U10378 (N_10378,N_1452,N_2255);
xor U10379 (N_10379,N_3452,N_511);
and U10380 (N_10380,N_4102,N_5936);
or U10381 (N_10381,N_5594,N_944);
nor U10382 (N_10382,N_2426,N_4919);
nand U10383 (N_10383,N_3254,N_3661);
or U10384 (N_10384,N_5234,N_5103);
nor U10385 (N_10385,N_3293,N_2061);
nand U10386 (N_10386,N_5213,N_2472);
xor U10387 (N_10387,N_6086,N_5479);
nand U10388 (N_10388,N_2110,N_816);
nand U10389 (N_10389,N_2346,N_3858);
and U10390 (N_10390,N_3190,N_2287);
xnor U10391 (N_10391,N_429,N_1351);
xor U10392 (N_10392,N_1000,N_408);
or U10393 (N_10393,N_1635,N_1034);
xnor U10394 (N_10394,N_3509,N_4436);
nor U10395 (N_10395,N_1802,N_6076);
nand U10396 (N_10396,N_4227,N_2409);
nor U10397 (N_10397,N_5861,N_829);
nor U10398 (N_10398,N_1804,N_993);
and U10399 (N_10399,N_3930,N_6108);
and U10400 (N_10400,N_3527,N_2297);
xor U10401 (N_10401,N_213,N_5689);
nand U10402 (N_10402,N_4863,N_4086);
or U10403 (N_10403,N_5682,N_5639);
nand U10404 (N_10404,N_5534,N_5621);
nor U10405 (N_10405,N_5117,N_3785);
or U10406 (N_10406,N_1142,N_1592);
xor U10407 (N_10407,N_2311,N_2255);
or U10408 (N_10408,N_4164,N_1956);
xnor U10409 (N_10409,N_771,N_1340);
nor U10410 (N_10410,N_3253,N_3669);
xor U10411 (N_10411,N_2862,N_4361);
or U10412 (N_10412,N_4236,N_593);
nor U10413 (N_10413,N_5612,N_1109);
nor U10414 (N_10414,N_4249,N_5629);
xnor U10415 (N_10415,N_3435,N_1711);
or U10416 (N_10416,N_3281,N_15);
or U10417 (N_10417,N_1125,N_2730);
xor U10418 (N_10418,N_1025,N_960);
nor U10419 (N_10419,N_3276,N_1865);
nand U10420 (N_10420,N_1666,N_3913);
and U10421 (N_10421,N_2530,N_4810);
xor U10422 (N_10422,N_3589,N_4819);
nand U10423 (N_10423,N_5669,N_5515);
xnor U10424 (N_10424,N_3403,N_3717);
nand U10425 (N_10425,N_5550,N_3495);
and U10426 (N_10426,N_6214,N_6224);
or U10427 (N_10427,N_1580,N_1651);
xor U10428 (N_10428,N_1023,N_1200);
and U10429 (N_10429,N_4212,N_221);
nor U10430 (N_10430,N_5784,N_1964);
and U10431 (N_10431,N_1681,N_3046);
xnor U10432 (N_10432,N_325,N_3902);
nor U10433 (N_10433,N_2316,N_4308);
xor U10434 (N_10434,N_3305,N_494);
nor U10435 (N_10435,N_2701,N_3122);
nor U10436 (N_10436,N_4574,N_1493);
nor U10437 (N_10437,N_5572,N_4335);
or U10438 (N_10438,N_4518,N_2984);
or U10439 (N_10439,N_1293,N_854);
nand U10440 (N_10440,N_3772,N_3463);
or U10441 (N_10441,N_1331,N_6134);
nor U10442 (N_10442,N_5907,N_2215);
nor U10443 (N_10443,N_4239,N_700);
nor U10444 (N_10444,N_6095,N_5324);
and U10445 (N_10445,N_5214,N_3818);
nor U10446 (N_10446,N_2863,N_4591);
nor U10447 (N_10447,N_2820,N_4061);
or U10448 (N_10448,N_2256,N_2525);
and U10449 (N_10449,N_33,N_4905);
nor U10450 (N_10450,N_2083,N_3390);
nand U10451 (N_10451,N_4967,N_2377);
xor U10452 (N_10452,N_282,N_1436);
and U10453 (N_10453,N_2344,N_5941);
or U10454 (N_10454,N_2083,N_5413);
nand U10455 (N_10455,N_2578,N_155);
nand U10456 (N_10456,N_4689,N_2837);
xor U10457 (N_10457,N_5793,N_1680);
nand U10458 (N_10458,N_868,N_5588);
nor U10459 (N_10459,N_5312,N_5358);
xor U10460 (N_10460,N_3571,N_2653);
nor U10461 (N_10461,N_1143,N_162);
xnor U10462 (N_10462,N_3877,N_3441);
and U10463 (N_10463,N_5246,N_176);
or U10464 (N_10464,N_5737,N_3925);
nand U10465 (N_10465,N_5669,N_184);
and U10466 (N_10466,N_5303,N_2065);
nor U10467 (N_10467,N_3604,N_3379);
or U10468 (N_10468,N_3944,N_4146);
nor U10469 (N_10469,N_734,N_4513);
nor U10470 (N_10470,N_4692,N_6052);
nand U10471 (N_10471,N_5415,N_1347);
and U10472 (N_10472,N_5202,N_4095);
nand U10473 (N_10473,N_887,N_747);
and U10474 (N_10474,N_2505,N_3902);
nand U10475 (N_10475,N_2049,N_722);
nand U10476 (N_10476,N_5884,N_5211);
nand U10477 (N_10477,N_690,N_1146);
or U10478 (N_10478,N_2960,N_3663);
nor U10479 (N_10479,N_2703,N_1857);
or U10480 (N_10480,N_3106,N_4036);
nand U10481 (N_10481,N_5584,N_508);
nor U10482 (N_10482,N_2025,N_3833);
xor U10483 (N_10483,N_744,N_2601);
and U10484 (N_10484,N_713,N_2508);
or U10485 (N_10485,N_1812,N_2560);
nor U10486 (N_10486,N_6147,N_5391);
nor U10487 (N_10487,N_1560,N_5176);
or U10488 (N_10488,N_180,N_68);
or U10489 (N_10489,N_2523,N_3812);
or U10490 (N_10490,N_2335,N_5379);
nor U10491 (N_10491,N_4880,N_4281);
nor U10492 (N_10492,N_5351,N_1563);
xor U10493 (N_10493,N_2995,N_6080);
and U10494 (N_10494,N_2962,N_5260);
or U10495 (N_10495,N_3999,N_771);
and U10496 (N_10496,N_5666,N_1188);
nor U10497 (N_10497,N_2738,N_5635);
nor U10498 (N_10498,N_4720,N_2950);
and U10499 (N_10499,N_194,N_1383);
nor U10500 (N_10500,N_1917,N_5559);
or U10501 (N_10501,N_1081,N_3907);
nor U10502 (N_10502,N_2928,N_6142);
nor U10503 (N_10503,N_3408,N_279);
or U10504 (N_10504,N_4743,N_5864);
nor U10505 (N_10505,N_3681,N_4018);
and U10506 (N_10506,N_4415,N_3592);
or U10507 (N_10507,N_3894,N_2988);
xor U10508 (N_10508,N_2409,N_3483);
or U10509 (N_10509,N_4683,N_1144);
or U10510 (N_10510,N_2379,N_766);
and U10511 (N_10511,N_691,N_6055);
nand U10512 (N_10512,N_5111,N_3405);
nor U10513 (N_10513,N_2730,N_4953);
nand U10514 (N_10514,N_322,N_2753);
nand U10515 (N_10515,N_1715,N_3403);
nor U10516 (N_10516,N_1871,N_198);
nor U10517 (N_10517,N_5994,N_3993);
nor U10518 (N_10518,N_5386,N_4759);
xor U10519 (N_10519,N_2547,N_2153);
xor U10520 (N_10520,N_1254,N_3926);
nand U10521 (N_10521,N_5112,N_2970);
or U10522 (N_10522,N_4968,N_76);
nand U10523 (N_10523,N_4311,N_5938);
nor U10524 (N_10524,N_800,N_5467);
nor U10525 (N_10525,N_5270,N_933);
xor U10526 (N_10526,N_4948,N_706);
nor U10527 (N_10527,N_2182,N_3065);
xor U10528 (N_10528,N_6081,N_3080);
and U10529 (N_10529,N_639,N_4719);
xnor U10530 (N_10530,N_1622,N_4630);
and U10531 (N_10531,N_5848,N_1887);
nand U10532 (N_10532,N_2556,N_5397);
nand U10533 (N_10533,N_283,N_2263);
nand U10534 (N_10534,N_4596,N_4828);
nor U10535 (N_10535,N_5067,N_3338);
nor U10536 (N_10536,N_3598,N_292);
nand U10537 (N_10537,N_3405,N_2888);
or U10538 (N_10538,N_4695,N_2018);
or U10539 (N_10539,N_818,N_5513);
or U10540 (N_10540,N_4530,N_562);
nor U10541 (N_10541,N_5857,N_5572);
xnor U10542 (N_10542,N_1983,N_4455);
xor U10543 (N_10543,N_6067,N_3678);
nor U10544 (N_10544,N_4546,N_2717);
xor U10545 (N_10545,N_664,N_1830);
nand U10546 (N_10546,N_5329,N_4054);
and U10547 (N_10547,N_5311,N_4962);
or U10548 (N_10548,N_1177,N_1496);
or U10549 (N_10549,N_3263,N_3363);
nor U10550 (N_10550,N_627,N_3584);
and U10551 (N_10551,N_1097,N_4669);
and U10552 (N_10552,N_611,N_4237);
nand U10553 (N_10553,N_2610,N_4245);
nand U10554 (N_10554,N_1991,N_1902);
xor U10555 (N_10555,N_1004,N_71);
nand U10556 (N_10556,N_1337,N_4171);
or U10557 (N_10557,N_3479,N_796);
nand U10558 (N_10558,N_130,N_3361);
or U10559 (N_10559,N_3347,N_444);
and U10560 (N_10560,N_1670,N_988);
or U10561 (N_10561,N_2634,N_1269);
nand U10562 (N_10562,N_4559,N_1339);
nor U10563 (N_10563,N_2163,N_493);
nand U10564 (N_10564,N_3905,N_5714);
and U10565 (N_10565,N_197,N_2814);
nand U10566 (N_10566,N_5290,N_5605);
or U10567 (N_10567,N_2160,N_1492);
xor U10568 (N_10568,N_5337,N_6225);
nor U10569 (N_10569,N_876,N_5448);
xnor U10570 (N_10570,N_3784,N_3319);
or U10571 (N_10571,N_3874,N_15);
nor U10572 (N_10572,N_1195,N_2881);
or U10573 (N_10573,N_3865,N_5545);
nor U10574 (N_10574,N_510,N_4769);
or U10575 (N_10575,N_1643,N_4812);
and U10576 (N_10576,N_2103,N_5892);
nand U10577 (N_10577,N_2943,N_2335);
xor U10578 (N_10578,N_5955,N_3216);
nand U10579 (N_10579,N_6211,N_5947);
nor U10580 (N_10580,N_5152,N_1310);
nor U10581 (N_10581,N_5596,N_2708);
nor U10582 (N_10582,N_5742,N_4903);
xnor U10583 (N_10583,N_5337,N_4024);
or U10584 (N_10584,N_4512,N_2305);
or U10585 (N_10585,N_4415,N_5180);
or U10586 (N_10586,N_4660,N_1782);
xnor U10587 (N_10587,N_3679,N_5071);
xor U10588 (N_10588,N_4274,N_1597);
and U10589 (N_10589,N_2825,N_2234);
xor U10590 (N_10590,N_475,N_1963);
xnor U10591 (N_10591,N_2920,N_4613);
nor U10592 (N_10592,N_5255,N_2574);
and U10593 (N_10593,N_3633,N_5026);
and U10594 (N_10594,N_5600,N_641);
nand U10595 (N_10595,N_768,N_4879);
and U10596 (N_10596,N_1741,N_2197);
or U10597 (N_10597,N_2214,N_2659);
and U10598 (N_10598,N_671,N_5385);
or U10599 (N_10599,N_3552,N_2545);
xnor U10600 (N_10600,N_5703,N_1635);
nor U10601 (N_10601,N_2585,N_231);
or U10602 (N_10602,N_2563,N_5305);
nor U10603 (N_10603,N_3555,N_4036);
nor U10604 (N_10604,N_2235,N_4374);
xnor U10605 (N_10605,N_3108,N_5546);
nor U10606 (N_10606,N_1741,N_3281);
and U10607 (N_10607,N_2936,N_2265);
and U10608 (N_10608,N_5357,N_673);
nand U10609 (N_10609,N_5384,N_1184);
nand U10610 (N_10610,N_6141,N_2214);
and U10611 (N_10611,N_2677,N_2896);
and U10612 (N_10612,N_2935,N_2502);
nor U10613 (N_10613,N_4200,N_2976);
xor U10614 (N_10614,N_285,N_4953);
nor U10615 (N_10615,N_2828,N_2015);
or U10616 (N_10616,N_1578,N_3300);
or U10617 (N_10617,N_2996,N_5512);
xnor U10618 (N_10618,N_5642,N_5098);
or U10619 (N_10619,N_5499,N_1122);
xor U10620 (N_10620,N_2322,N_269);
nor U10621 (N_10621,N_4327,N_3852);
xnor U10622 (N_10622,N_4538,N_5918);
or U10623 (N_10623,N_2233,N_4998);
xnor U10624 (N_10624,N_2678,N_1522);
nor U10625 (N_10625,N_1019,N_4212);
or U10626 (N_10626,N_2220,N_3646);
and U10627 (N_10627,N_311,N_946);
nor U10628 (N_10628,N_5549,N_5109);
and U10629 (N_10629,N_6057,N_1169);
xor U10630 (N_10630,N_819,N_1496);
and U10631 (N_10631,N_2320,N_5166);
nor U10632 (N_10632,N_2643,N_4400);
or U10633 (N_10633,N_3956,N_3627);
xnor U10634 (N_10634,N_2656,N_2165);
nor U10635 (N_10635,N_5264,N_422);
and U10636 (N_10636,N_362,N_5212);
or U10637 (N_10637,N_4636,N_4552);
nor U10638 (N_10638,N_3877,N_2771);
and U10639 (N_10639,N_902,N_2903);
xnor U10640 (N_10640,N_1535,N_5020);
or U10641 (N_10641,N_184,N_5584);
and U10642 (N_10642,N_1932,N_3657);
or U10643 (N_10643,N_4060,N_4031);
and U10644 (N_10644,N_3241,N_3469);
and U10645 (N_10645,N_1949,N_6186);
xnor U10646 (N_10646,N_5158,N_4351);
and U10647 (N_10647,N_472,N_2543);
xnor U10648 (N_10648,N_3468,N_992);
xnor U10649 (N_10649,N_3849,N_4719);
and U10650 (N_10650,N_3522,N_2491);
nand U10651 (N_10651,N_5948,N_4513);
or U10652 (N_10652,N_1620,N_6219);
xor U10653 (N_10653,N_3573,N_6217);
nor U10654 (N_10654,N_2161,N_3062);
or U10655 (N_10655,N_2126,N_2036);
xor U10656 (N_10656,N_4909,N_6088);
nor U10657 (N_10657,N_5447,N_1391);
xnor U10658 (N_10658,N_2258,N_4);
and U10659 (N_10659,N_989,N_1488);
nand U10660 (N_10660,N_2494,N_1618);
and U10661 (N_10661,N_4924,N_3075);
and U10662 (N_10662,N_2755,N_4044);
nor U10663 (N_10663,N_1612,N_2375);
or U10664 (N_10664,N_1156,N_1669);
nand U10665 (N_10665,N_2863,N_3439);
xnor U10666 (N_10666,N_961,N_556);
xor U10667 (N_10667,N_5996,N_1017);
nor U10668 (N_10668,N_5659,N_428);
nand U10669 (N_10669,N_1985,N_5857);
xnor U10670 (N_10670,N_1579,N_3442);
or U10671 (N_10671,N_3931,N_1564);
nor U10672 (N_10672,N_5610,N_3478);
xnor U10673 (N_10673,N_5462,N_5472);
nand U10674 (N_10674,N_2211,N_5648);
and U10675 (N_10675,N_340,N_3647);
nand U10676 (N_10676,N_5234,N_4369);
nor U10677 (N_10677,N_4966,N_3506);
xor U10678 (N_10678,N_5465,N_5572);
nor U10679 (N_10679,N_5795,N_2825);
and U10680 (N_10680,N_5151,N_815);
nor U10681 (N_10681,N_3734,N_3514);
nor U10682 (N_10682,N_736,N_5709);
xor U10683 (N_10683,N_754,N_2469);
nand U10684 (N_10684,N_1530,N_1225);
and U10685 (N_10685,N_3966,N_972);
or U10686 (N_10686,N_5664,N_5399);
nor U10687 (N_10687,N_4916,N_2656);
nor U10688 (N_10688,N_3642,N_3057);
and U10689 (N_10689,N_2711,N_2736);
nor U10690 (N_10690,N_4051,N_4383);
nor U10691 (N_10691,N_3464,N_4723);
xnor U10692 (N_10692,N_3064,N_653);
xor U10693 (N_10693,N_3887,N_4229);
nor U10694 (N_10694,N_2503,N_1511);
nor U10695 (N_10695,N_121,N_389);
nand U10696 (N_10696,N_3771,N_495);
and U10697 (N_10697,N_4535,N_4465);
nand U10698 (N_10698,N_1059,N_5482);
and U10699 (N_10699,N_3477,N_2210);
xnor U10700 (N_10700,N_264,N_3516);
nor U10701 (N_10701,N_301,N_1337);
nand U10702 (N_10702,N_4527,N_4359);
nor U10703 (N_10703,N_473,N_1991);
and U10704 (N_10704,N_166,N_930);
and U10705 (N_10705,N_1335,N_2300);
nor U10706 (N_10706,N_496,N_2593);
nand U10707 (N_10707,N_6158,N_4255);
nor U10708 (N_10708,N_5711,N_557);
or U10709 (N_10709,N_2802,N_4347);
xnor U10710 (N_10710,N_3152,N_4291);
xnor U10711 (N_10711,N_3782,N_3162);
xor U10712 (N_10712,N_161,N_2337);
nor U10713 (N_10713,N_2409,N_6066);
and U10714 (N_10714,N_4707,N_2020);
or U10715 (N_10715,N_5589,N_3528);
nor U10716 (N_10716,N_5399,N_4747);
or U10717 (N_10717,N_3645,N_1953);
xor U10718 (N_10718,N_1606,N_3069);
or U10719 (N_10719,N_2742,N_1031);
or U10720 (N_10720,N_2347,N_3310);
nor U10721 (N_10721,N_2433,N_463);
or U10722 (N_10722,N_922,N_2390);
nand U10723 (N_10723,N_3839,N_3596);
and U10724 (N_10724,N_4924,N_5468);
nor U10725 (N_10725,N_1001,N_4672);
and U10726 (N_10726,N_5258,N_890);
nor U10727 (N_10727,N_3864,N_3779);
nor U10728 (N_10728,N_81,N_1664);
and U10729 (N_10729,N_2646,N_1720);
nor U10730 (N_10730,N_6043,N_5093);
or U10731 (N_10731,N_2061,N_1410);
nor U10732 (N_10732,N_4662,N_2461);
and U10733 (N_10733,N_2232,N_821);
or U10734 (N_10734,N_5066,N_2360);
and U10735 (N_10735,N_4130,N_167);
or U10736 (N_10736,N_3404,N_5929);
nand U10737 (N_10737,N_2703,N_2326);
or U10738 (N_10738,N_484,N_728);
xor U10739 (N_10739,N_5850,N_2357);
and U10740 (N_10740,N_1368,N_2278);
or U10741 (N_10741,N_4104,N_213);
and U10742 (N_10742,N_46,N_5881);
and U10743 (N_10743,N_828,N_4864);
and U10744 (N_10744,N_1536,N_953);
nand U10745 (N_10745,N_3203,N_2682);
nand U10746 (N_10746,N_1378,N_6073);
nor U10747 (N_10747,N_2993,N_485);
or U10748 (N_10748,N_3600,N_4180);
nor U10749 (N_10749,N_1139,N_351);
nand U10750 (N_10750,N_1955,N_5802);
xor U10751 (N_10751,N_1107,N_4177);
or U10752 (N_10752,N_4928,N_1853);
nand U10753 (N_10753,N_5101,N_3454);
and U10754 (N_10754,N_135,N_3743);
or U10755 (N_10755,N_5403,N_4330);
and U10756 (N_10756,N_5643,N_3818);
nand U10757 (N_10757,N_5498,N_3024);
nand U10758 (N_10758,N_2315,N_5028);
and U10759 (N_10759,N_4595,N_1404);
or U10760 (N_10760,N_1253,N_6015);
and U10761 (N_10761,N_3637,N_4130);
nor U10762 (N_10762,N_4203,N_5247);
nand U10763 (N_10763,N_2012,N_1342);
or U10764 (N_10764,N_4933,N_269);
or U10765 (N_10765,N_396,N_3069);
nor U10766 (N_10766,N_4740,N_1586);
nand U10767 (N_10767,N_3385,N_5517);
or U10768 (N_10768,N_12,N_4759);
nand U10769 (N_10769,N_5845,N_2328);
xor U10770 (N_10770,N_4913,N_2251);
nand U10771 (N_10771,N_4664,N_4213);
or U10772 (N_10772,N_2475,N_4389);
or U10773 (N_10773,N_52,N_1194);
xnor U10774 (N_10774,N_3054,N_138);
or U10775 (N_10775,N_645,N_5486);
xnor U10776 (N_10776,N_3199,N_428);
nand U10777 (N_10777,N_920,N_3534);
nor U10778 (N_10778,N_3568,N_4528);
nor U10779 (N_10779,N_3556,N_2588);
xnor U10780 (N_10780,N_4906,N_6132);
or U10781 (N_10781,N_2131,N_1957);
nor U10782 (N_10782,N_779,N_1438);
or U10783 (N_10783,N_1224,N_4393);
nand U10784 (N_10784,N_3799,N_5290);
xor U10785 (N_10785,N_4816,N_4035);
nand U10786 (N_10786,N_1633,N_1063);
nor U10787 (N_10787,N_1450,N_759);
nand U10788 (N_10788,N_5280,N_1032);
nand U10789 (N_10789,N_5135,N_5109);
nand U10790 (N_10790,N_3234,N_5144);
and U10791 (N_10791,N_3995,N_2004);
nand U10792 (N_10792,N_5977,N_4808);
nor U10793 (N_10793,N_3149,N_3099);
nand U10794 (N_10794,N_441,N_3604);
and U10795 (N_10795,N_769,N_3597);
and U10796 (N_10796,N_5544,N_5963);
nand U10797 (N_10797,N_6205,N_5927);
nand U10798 (N_10798,N_2732,N_3736);
nand U10799 (N_10799,N_724,N_3837);
and U10800 (N_10800,N_4474,N_3258);
and U10801 (N_10801,N_4304,N_4032);
nand U10802 (N_10802,N_5927,N_4267);
xor U10803 (N_10803,N_873,N_825);
xor U10804 (N_10804,N_2205,N_350);
or U10805 (N_10805,N_2211,N_862);
or U10806 (N_10806,N_78,N_4366);
nand U10807 (N_10807,N_470,N_3860);
xnor U10808 (N_10808,N_299,N_4832);
nand U10809 (N_10809,N_3246,N_5132);
nor U10810 (N_10810,N_3885,N_4935);
and U10811 (N_10811,N_2095,N_5050);
nand U10812 (N_10812,N_5055,N_2307);
or U10813 (N_10813,N_961,N_261);
nand U10814 (N_10814,N_1634,N_1934);
or U10815 (N_10815,N_5680,N_5225);
nor U10816 (N_10816,N_1078,N_313);
nand U10817 (N_10817,N_1106,N_1671);
or U10818 (N_10818,N_3384,N_5188);
and U10819 (N_10819,N_2102,N_453);
nor U10820 (N_10820,N_4949,N_4057);
and U10821 (N_10821,N_1550,N_640);
xor U10822 (N_10822,N_3097,N_5923);
nor U10823 (N_10823,N_4040,N_5515);
nand U10824 (N_10824,N_1176,N_4850);
xor U10825 (N_10825,N_530,N_3532);
xor U10826 (N_10826,N_3102,N_4901);
or U10827 (N_10827,N_5170,N_3244);
or U10828 (N_10828,N_5368,N_3587);
or U10829 (N_10829,N_4633,N_6078);
or U10830 (N_10830,N_4852,N_2258);
and U10831 (N_10831,N_388,N_2643);
or U10832 (N_10832,N_4317,N_1170);
and U10833 (N_10833,N_1794,N_3045);
and U10834 (N_10834,N_74,N_4435);
nor U10835 (N_10835,N_932,N_2261);
and U10836 (N_10836,N_3033,N_761);
and U10837 (N_10837,N_3353,N_5731);
nor U10838 (N_10838,N_3125,N_6113);
nor U10839 (N_10839,N_4259,N_2032);
and U10840 (N_10840,N_175,N_4863);
and U10841 (N_10841,N_1426,N_334);
nand U10842 (N_10842,N_2487,N_3697);
or U10843 (N_10843,N_301,N_4686);
and U10844 (N_10844,N_1702,N_4802);
nor U10845 (N_10845,N_527,N_279);
and U10846 (N_10846,N_613,N_5944);
nor U10847 (N_10847,N_3454,N_4235);
nand U10848 (N_10848,N_1137,N_1910);
or U10849 (N_10849,N_161,N_3488);
nor U10850 (N_10850,N_4525,N_206);
nor U10851 (N_10851,N_3762,N_5981);
xnor U10852 (N_10852,N_1809,N_4337);
xnor U10853 (N_10853,N_2585,N_5959);
xor U10854 (N_10854,N_6237,N_4138);
nor U10855 (N_10855,N_5974,N_1003);
or U10856 (N_10856,N_4378,N_131);
nor U10857 (N_10857,N_3060,N_514);
xor U10858 (N_10858,N_1721,N_3443);
or U10859 (N_10859,N_4899,N_1354);
nand U10860 (N_10860,N_5843,N_250);
xnor U10861 (N_10861,N_1592,N_4471);
nand U10862 (N_10862,N_4733,N_4325);
and U10863 (N_10863,N_1741,N_1421);
or U10864 (N_10864,N_3789,N_5472);
nand U10865 (N_10865,N_1555,N_1631);
and U10866 (N_10866,N_4996,N_1388);
nand U10867 (N_10867,N_5466,N_4949);
and U10868 (N_10868,N_3097,N_4983);
and U10869 (N_10869,N_5237,N_3946);
or U10870 (N_10870,N_5879,N_5289);
and U10871 (N_10871,N_1340,N_3875);
nor U10872 (N_10872,N_4209,N_4893);
or U10873 (N_10873,N_3934,N_1613);
nand U10874 (N_10874,N_3036,N_5677);
and U10875 (N_10875,N_1904,N_6053);
nand U10876 (N_10876,N_2335,N_1279);
nor U10877 (N_10877,N_383,N_3005);
nor U10878 (N_10878,N_1618,N_11);
xnor U10879 (N_10879,N_3327,N_154);
nand U10880 (N_10880,N_1687,N_2155);
or U10881 (N_10881,N_4697,N_571);
and U10882 (N_10882,N_508,N_4806);
nand U10883 (N_10883,N_2090,N_3391);
xor U10884 (N_10884,N_2158,N_6200);
nand U10885 (N_10885,N_5566,N_4724);
xor U10886 (N_10886,N_5275,N_5985);
or U10887 (N_10887,N_3815,N_1750);
nor U10888 (N_10888,N_3014,N_3631);
nor U10889 (N_10889,N_6077,N_4705);
or U10890 (N_10890,N_5426,N_1405);
nand U10891 (N_10891,N_5602,N_465);
nand U10892 (N_10892,N_3252,N_5478);
and U10893 (N_10893,N_2531,N_5397);
xnor U10894 (N_10894,N_4213,N_2351);
and U10895 (N_10895,N_4358,N_5438);
nand U10896 (N_10896,N_2659,N_5783);
xnor U10897 (N_10897,N_5194,N_5623);
xor U10898 (N_10898,N_4490,N_4051);
and U10899 (N_10899,N_6015,N_5368);
and U10900 (N_10900,N_4882,N_3935);
nor U10901 (N_10901,N_259,N_2130);
xnor U10902 (N_10902,N_1956,N_3031);
nor U10903 (N_10903,N_4744,N_5924);
nand U10904 (N_10904,N_2507,N_1967);
xor U10905 (N_10905,N_293,N_3357);
and U10906 (N_10906,N_2194,N_5364);
or U10907 (N_10907,N_1269,N_4055);
nor U10908 (N_10908,N_467,N_4596);
nand U10909 (N_10909,N_1794,N_4072);
nor U10910 (N_10910,N_5408,N_3344);
nor U10911 (N_10911,N_4459,N_3698);
nor U10912 (N_10912,N_856,N_2457);
and U10913 (N_10913,N_768,N_2706);
nor U10914 (N_10914,N_2799,N_2877);
nor U10915 (N_10915,N_3730,N_1116);
and U10916 (N_10916,N_5166,N_4180);
or U10917 (N_10917,N_830,N_4348);
nor U10918 (N_10918,N_4715,N_1949);
nor U10919 (N_10919,N_4627,N_5838);
and U10920 (N_10920,N_2421,N_2331);
or U10921 (N_10921,N_1227,N_5902);
xor U10922 (N_10922,N_3654,N_5025);
or U10923 (N_10923,N_907,N_1409);
nand U10924 (N_10924,N_3353,N_302);
or U10925 (N_10925,N_2147,N_1437);
and U10926 (N_10926,N_4753,N_4863);
or U10927 (N_10927,N_5655,N_789);
nor U10928 (N_10928,N_293,N_4983);
or U10929 (N_10929,N_1712,N_4255);
xnor U10930 (N_10930,N_106,N_3779);
or U10931 (N_10931,N_2586,N_1028);
nor U10932 (N_10932,N_2490,N_3469);
and U10933 (N_10933,N_2865,N_6027);
and U10934 (N_10934,N_892,N_3716);
xnor U10935 (N_10935,N_3754,N_2600);
nor U10936 (N_10936,N_2440,N_3024);
nand U10937 (N_10937,N_4806,N_1942);
or U10938 (N_10938,N_2017,N_1587);
nand U10939 (N_10939,N_1501,N_5063);
or U10940 (N_10940,N_4659,N_4902);
and U10941 (N_10941,N_4175,N_5335);
and U10942 (N_10942,N_2796,N_4589);
and U10943 (N_10943,N_5886,N_4633);
xor U10944 (N_10944,N_5946,N_719);
nor U10945 (N_10945,N_1536,N_447);
and U10946 (N_10946,N_633,N_5707);
or U10947 (N_10947,N_6017,N_3062);
xnor U10948 (N_10948,N_2693,N_2738);
nor U10949 (N_10949,N_2992,N_2776);
or U10950 (N_10950,N_5848,N_3277);
nor U10951 (N_10951,N_3651,N_2142);
xor U10952 (N_10952,N_1393,N_6233);
nand U10953 (N_10953,N_5511,N_5412);
and U10954 (N_10954,N_3735,N_3187);
or U10955 (N_10955,N_710,N_190);
nand U10956 (N_10956,N_3284,N_2799);
xnor U10957 (N_10957,N_4169,N_672);
nand U10958 (N_10958,N_2832,N_4267);
nand U10959 (N_10959,N_5632,N_4125);
nor U10960 (N_10960,N_3131,N_936);
nand U10961 (N_10961,N_142,N_6177);
nand U10962 (N_10962,N_5436,N_1014);
xnor U10963 (N_10963,N_1372,N_3005);
or U10964 (N_10964,N_2170,N_4382);
nand U10965 (N_10965,N_103,N_190);
xor U10966 (N_10966,N_5074,N_4496);
nor U10967 (N_10967,N_4271,N_2741);
nor U10968 (N_10968,N_4988,N_4802);
nand U10969 (N_10969,N_2500,N_1707);
xor U10970 (N_10970,N_4672,N_3040);
nor U10971 (N_10971,N_3418,N_2773);
and U10972 (N_10972,N_3448,N_4714);
or U10973 (N_10973,N_6054,N_2447);
and U10974 (N_10974,N_3083,N_1934);
nor U10975 (N_10975,N_5382,N_5657);
nand U10976 (N_10976,N_2014,N_2875);
and U10977 (N_10977,N_3515,N_1505);
xor U10978 (N_10978,N_1701,N_890);
and U10979 (N_10979,N_14,N_2691);
xor U10980 (N_10980,N_1428,N_3161);
or U10981 (N_10981,N_3546,N_843);
xor U10982 (N_10982,N_4413,N_3133);
and U10983 (N_10983,N_4622,N_5861);
nor U10984 (N_10984,N_2717,N_4704);
or U10985 (N_10985,N_430,N_2504);
and U10986 (N_10986,N_5235,N_3801);
xnor U10987 (N_10987,N_6132,N_4225);
or U10988 (N_10988,N_3791,N_1158);
xor U10989 (N_10989,N_4687,N_1306);
nand U10990 (N_10990,N_4882,N_2339);
nor U10991 (N_10991,N_4458,N_2110);
nand U10992 (N_10992,N_3891,N_3711);
nor U10993 (N_10993,N_4426,N_2538);
xor U10994 (N_10994,N_4512,N_3717);
or U10995 (N_10995,N_4521,N_5595);
nand U10996 (N_10996,N_4313,N_2105);
nand U10997 (N_10997,N_3300,N_3357);
and U10998 (N_10998,N_1004,N_2081);
nand U10999 (N_10999,N_6196,N_6156);
nor U11000 (N_11000,N_4929,N_3503);
or U11001 (N_11001,N_4380,N_5591);
nor U11002 (N_11002,N_3309,N_3934);
and U11003 (N_11003,N_1304,N_2243);
nor U11004 (N_11004,N_80,N_4801);
and U11005 (N_11005,N_4640,N_745);
xor U11006 (N_11006,N_1316,N_4902);
xnor U11007 (N_11007,N_4555,N_395);
or U11008 (N_11008,N_2154,N_1226);
nor U11009 (N_11009,N_2153,N_1841);
nand U11010 (N_11010,N_2929,N_4067);
xnor U11011 (N_11011,N_2044,N_2399);
and U11012 (N_11012,N_2584,N_3307);
xnor U11013 (N_11013,N_3088,N_2264);
nor U11014 (N_11014,N_35,N_2174);
and U11015 (N_11015,N_608,N_1502);
or U11016 (N_11016,N_3336,N_3176);
nor U11017 (N_11017,N_2082,N_3302);
xnor U11018 (N_11018,N_5606,N_1479);
nand U11019 (N_11019,N_1726,N_2753);
and U11020 (N_11020,N_5507,N_1229);
nand U11021 (N_11021,N_5674,N_4161);
xor U11022 (N_11022,N_1035,N_4605);
nor U11023 (N_11023,N_5962,N_3728);
xnor U11024 (N_11024,N_4160,N_3599);
xor U11025 (N_11025,N_2339,N_1372);
nand U11026 (N_11026,N_3823,N_2005);
and U11027 (N_11027,N_2672,N_1020);
nand U11028 (N_11028,N_928,N_179);
xnor U11029 (N_11029,N_2451,N_6045);
and U11030 (N_11030,N_4910,N_2867);
nor U11031 (N_11031,N_41,N_3948);
xor U11032 (N_11032,N_5749,N_71);
nor U11033 (N_11033,N_3410,N_5009);
nor U11034 (N_11034,N_3907,N_2267);
and U11035 (N_11035,N_4626,N_1463);
nand U11036 (N_11036,N_2883,N_3952);
and U11037 (N_11037,N_1792,N_4137);
nor U11038 (N_11038,N_3794,N_4485);
nor U11039 (N_11039,N_4292,N_15);
and U11040 (N_11040,N_3052,N_5165);
nor U11041 (N_11041,N_4,N_3889);
nand U11042 (N_11042,N_6027,N_3689);
or U11043 (N_11043,N_4409,N_3633);
xor U11044 (N_11044,N_4176,N_5895);
nand U11045 (N_11045,N_884,N_220);
nand U11046 (N_11046,N_3241,N_2168);
nand U11047 (N_11047,N_793,N_2959);
xnor U11048 (N_11048,N_2645,N_5992);
nand U11049 (N_11049,N_4588,N_119);
xnor U11050 (N_11050,N_788,N_5095);
nand U11051 (N_11051,N_2998,N_6200);
nor U11052 (N_11052,N_4250,N_5470);
nand U11053 (N_11053,N_459,N_8);
and U11054 (N_11054,N_5207,N_1439);
or U11055 (N_11055,N_3126,N_2513);
nor U11056 (N_11056,N_6088,N_3509);
nor U11057 (N_11057,N_77,N_394);
nand U11058 (N_11058,N_43,N_856);
nand U11059 (N_11059,N_1318,N_2176);
xor U11060 (N_11060,N_5408,N_604);
and U11061 (N_11061,N_4914,N_2156);
or U11062 (N_11062,N_3818,N_3667);
nand U11063 (N_11063,N_5349,N_745);
nand U11064 (N_11064,N_290,N_1180);
nor U11065 (N_11065,N_4558,N_1370);
and U11066 (N_11066,N_1618,N_2542);
nor U11067 (N_11067,N_5772,N_3944);
or U11068 (N_11068,N_3292,N_4381);
nand U11069 (N_11069,N_4271,N_6169);
xor U11070 (N_11070,N_328,N_3708);
xnor U11071 (N_11071,N_4130,N_4792);
nand U11072 (N_11072,N_4319,N_3987);
and U11073 (N_11073,N_3043,N_2070);
or U11074 (N_11074,N_3713,N_2212);
or U11075 (N_11075,N_5694,N_4965);
or U11076 (N_11076,N_3825,N_5290);
and U11077 (N_11077,N_2755,N_3369);
or U11078 (N_11078,N_2882,N_1133);
nand U11079 (N_11079,N_945,N_1454);
nor U11080 (N_11080,N_3252,N_3282);
xnor U11081 (N_11081,N_2735,N_5469);
or U11082 (N_11082,N_2752,N_2320);
xnor U11083 (N_11083,N_432,N_1696);
nand U11084 (N_11084,N_3162,N_1354);
and U11085 (N_11085,N_4210,N_3449);
or U11086 (N_11086,N_4702,N_1757);
xor U11087 (N_11087,N_2071,N_2578);
nor U11088 (N_11088,N_4053,N_1416);
nor U11089 (N_11089,N_3854,N_2247);
xor U11090 (N_11090,N_4630,N_6013);
and U11091 (N_11091,N_1251,N_4335);
nor U11092 (N_11092,N_5914,N_3338);
nor U11093 (N_11093,N_2222,N_4078);
nor U11094 (N_11094,N_716,N_4163);
and U11095 (N_11095,N_3136,N_1427);
nor U11096 (N_11096,N_4614,N_5342);
nor U11097 (N_11097,N_4074,N_5470);
nor U11098 (N_11098,N_3920,N_4572);
nor U11099 (N_11099,N_811,N_5226);
nor U11100 (N_11100,N_592,N_270);
or U11101 (N_11101,N_1504,N_3245);
or U11102 (N_11102,N_6021,N_3042);
and U11103 (N_11103,N_4752,N_4755);
or U11104 (N_11104,N_1178,N_4418);
xnor U11105 (N_11105,N_6107,N_4117);
or U11106 (N_11106,N_5891,N_6203);
or U11107 (N_11107,N_5073,N_1726);
or U11108 (N_11108,N_5328,N_2146);
nand U11109 (N_11109,N_5665,N_2623);
nand U11110 (N_11110,N_2315,N_4326);
nand U11111 (N_11111,N_1465,N_5262);
or U11112 (N_11112,N_3608,N_6046);
nand U11113 (N_11113,N_4054,N_4994);
nand U11114 (N_11114,N_4487,N_2237);
nor U11115 (N_11115,N_2800,N_1211);
nand U11116 (N_11116,N_3713,N_2195);
nand U11117 (N_11117,N_4183,N_4733);
or U11118 (N_11118,N_4790,N_3893);
xor U11119 (N_11119,N_2906,N_4222);
nand U11120 (N_11120,N_3345,N_4557);
and U11121 (N_11121,N_1004,N_2628);
and U11122 (N_11122,N_2364,N_2469);
nor U11123 (N_11123,N_4449,N_1111);
or U11124 (N_11124,N_3936,N_6015);
nand U11125 (N_11125,N_2583,N_5180);
or U11126 (N_11126,N_6116,N_1177);
and U11127 (N_11127,N_899,N_5748);
and U11128 (N_11128,N_2632,N_1215);
and U11129 (N_11129,N_5348,N_2714);
nand U11130 (N_11130,N_648,N_911);
nor U11131 (N_11131,N_1742,N_3925);
nor U11132 (N_11132,N_1032,N_892);
xnor U11133 (N_11133,N_5443,N_2070);
and U11134 (N_11134,N_3104,N_3358);
and U11135 (N_11135,N_1435,N_1652);
nor U11136 (N_11136,N_5162,N_590);
xnor U11137 (N_11137,N_3287,N_4444);
and U11138 (N_11138,N_2362,N_4903);
nor U11139 (N_11139,N_3974,N_3820);
and U11140 (N_11140,N_2777,N_3836);
xor U11141 (N_11141,N_69,N_3112);
nor U11142 (N_11142,N_696,N_2832);
nand U11143 (N_11143,N_1981,N_2639);
nand U11144 (N_11144,N_6179,N_3330);
xor U11145 (N_11145,N_1751,N_1159);
and U11146 (N_11146,N_5845,N_5629);
or U11147 (N_11147,N_433,N_2627);
nor U11148 (N_11148,N_2270,N_830);
nand U11149 (N_11149,N_835,N_1853);
xnor U11150 (N_11150,N_4717,N_4841);
and U11151 (N_11151,N_1832,N_3178);
nand U11152 (N_11152,N_3662,N_5742);
or U11153 (N_11153,N_1621,N_4798);
or U11154 (N_11154,N_2450,N_5854);
nand U11155 (N_11155,N_1775,N_2965);
nor U11156 (N_11156,N_5563,N_980);
xnor U11157 (N_11157,N_1182,N_2559);
nand U11158 (N_11158,N_716,N_1167);
nand U11159 (N_11159,N_4014,N_2290);
xor U11160 (N_11160,N_6083,N_5405);
and U11161 (N_11161,N_549,N_5060);
xnor U11162 (N_11162,N_635,N_5623);
nand U11163 (N_11163,N_342,N_3183);
nand U11164 (N_11164,N_2293,N_4812);
or U11165 (N_11165,N_3146,N_4030);
nand U11166 (N_11166,N_2572,N_4826);
and U11167 (N_11167,N_2806,N_5890);
and U11168 (N_11168,N_428,N_1983);
nor U11169 (N_11169,N_859,N_4199);
nand U11170 (N_11170,N_500,N_5267);
xnor U11171 (N_11171,N_1053,N_2849);
or U11172 (N_11172,N_4208,N_1393);
and U11173 (N_11173,N_1676,N_742);
nor U11174 (N_11174,N_5718,N_3312);
or U11175 (N_11175,N_783,N_3793);
nor U11176 (N_11176,N_5406,N_5919);
nand U11177 (N_11177,N_5915,N_3953);
nand U11178 (N_11178,N_4016,N_212);
and U11179 (N_11179,N_5201,N_3513);
or U11180 (N_11180,N_4726,N_2484);
nand U11181 (N_11181,N_2666,N_377);
nor U11182 (N_11182,N_2763,N_2588);
nand U11183 (N_11183,N_262,N_3679);
nand U11184 (N_11184,N_2035,N_5598);
or U11185 (N_11185,N_5393,N_2133);
or U11186 (N_11186,N_2737,N_5146);
nor U11187 (N_11187,N_5366,N_6084);
or U11188 (N_11188,N_6169,N_658);
and U11189 (N_11189,N_2952,N_1050);
nand U11190 (N_11190,N_6216,N_1973);
nand U11191 (N_11191,N_5069,N_1085);
xor U11192 (N_11192,N_490,N_1868);
and U11193 (N_11193,N_5979,N_1951);
xor U11194 (N_11194,N_1471,N_2150);
nand U11195 (N_11195,N_4038,N_3133);
or U11196 (N_11196,N_1362,N_671);
nor U11197 (N_11197,N_3291,N_6078);
and U11198 (N_11198,N_907,N_3066);
and U11199 (N_11199,N_4723,N_5923);
nor U11200 (N_11200,N_1114,N_2980);
or U11201 (N_11201,N_3573,N_4303);
and U11202 (N_11202,N_2927,N_3605);
nor U11203 (N_11203,N_4770,N_1923);
xnor U11204 (N_11204,N_3135,N_4844);
nor U11205 (N_11205,N_1890,N_3330);
nand U11206 (N_11206,N_1365,N_4888);
xnor U11207 (N_11207,N_4901,N_1995);
xor U11208 (N_11208,N_6196,N_5184);
or U11209 (N_11209,N_3172,N_1458);
nor U11210 (N_11210,N_4097,N_2504);
xor U11211 (N_11211,N_3086,N_6186);
xnor U11212 (N_11212,N_4595,N_2435);
xnor U11213 (N_11213,N_878,N_411);
nor U11214 (N_11214,N_5815,N_4970);
or U11215 (N_11215,N_6237,N_1582);
nor U11216 (N_11216,N_2078,N_3032);
and U11217 (N_11217,N_6066,N_6242);
and U11218 (N_11218,N_3513,N_2417);
or U11219 (N_11219,N_5770,N_4545);
or U11220 (N_11220,N_2760,N_4693);
xnor U11221 (N_11221,N_9,N_1164);
and U11222 (N_11222,N_2217,N_52);
nor U11223 (N_11223,N_5167,N_4581);
nand U11224 (N_11224,N_1900,N_3076);
or U11225 (N_11225,N_251,N_5229);
nor U11226 (N_11226,N_1284,N_1633);
or U11227 (N_11227,N_4118,N_563);
or U11228 (N_11228,N_1863,N_3538);
nand U11229 (N_11229,N_6070,N_1350);
and U11230 (N_11230,N_5045,N_3046);
nand U11231 (N_11231,N_2692,N_1691);
nand U11232 (N_11232,N_418,N_2878);
or U11233 (N_11233,N_327,N_5359);
nor U11234 (N_11234,N_2571,N_4477);
xor U11235 (N_11235,N_6181,N_804);
or U11236 (N_11236,N_4727,N_3818);
xnor U11237 (N_11237,N_328,N_2707);
nor U11238 (N_11238,N_458,N_2194);
and U11239 (N_11239,N_5671,N_5217);
xnor U11240 (N_11240,N_4448,N_506);
xnor U11241 (N_11241,N_1057,N_574);
nand U11242 (N_11242,N_5794,N_3109);
nand U11243 (N_11243,N_2648,N_1921);
and U11244 (N_11244,N_3185,N_1643);
nor U11245 (N_11245,N_3873,N_4949);
xnor U11246 (N_11246,N_5130,N_874);
nor U11247 (N_11247,N_3320,N_3964);
nor U11248 (N_11248,N_5050,N_598);
or U11249 (N_11249,N_4477,N_3483);
nand U11250 (N_11250,N_308,N_5072);
and U11251 (N_11251,N_144,N_3591);
xnor U11252 (N_11252,N_2186,N_1377);
nor U11253 (N_11253,N_2215,N_2664);
nand U11254 (N_11254,N_507,N_5394);
or U11255 (N_11255,N_6189,N_2153);
nand U11256 (N_11256,N_2067,N_1713);
xor U11257 (N_11257,N_749,N_1493);
nand U11258 (N_11258,N_855,N_2549);
and U11259 (N_11259,N_5983,N_796);
and U11260 (N_11260,N_2262,N_366);
nor U11261 (N_11261,N_5105,N_5938);
nand U11262 (N_11262,N_1769,N_1130);
or U11263 (N_11263,N_6055,N_4591);
nand U11264 (N_11264,N_3342,N_2261);
xor U11265 (N_11265,N_385,N_5520);
or U11266 (N_11266,N_5116,N_3896);
xor U11267 (N_11267,N_1175,N_2520);
and U11268 (N_11268,N_3995,N_2519);
xor U11269 (N_11269,N_2348,N_5043);
xor U11270 (N_11270,N_3376,N_5442);
or U11271 (N_11271,N_5604,N_2747);
nor U11272 (N_11272,N_6069,N_1103);
or U11273 (N_11273,N_895,N_2615);
nand U11274 (N_11274,N_3414,N_4055);
and U11275 (N_11275,N_3780,N_4978);
or U11276 (N_11276,N_5514,N_4969);
nand U11277 (N_11277,N_1539,N_1996);
nand U11278 (N_11278,N_403,N_2466);
nor U11279 (N_11279,N_587,N_121);
and U11280 (N_11280,N_3233,N_1083);
nand U11281 (N_11281,N_3547,N_5778);
xnor U11282 (N_11282,N_4281,N_6186);
xor U11283 (N_11283,N_846,N_4743);
and U11284 (N_11284,N_5352,N_5939);
or U11285 (N_11285,N_3728,N_2648);
nand U11286 (N_11286,N_2368,N_4721);
xnor U11287 (N_11287,N_1863,N_4277);
nor U11288 (N_11288,N_168,N_6226);
nand U11289 (N_11289,N_1512,N_6240);
or U11290 (N_11290,N_3564,N_6223);
nor U11291 (N_11291,N_4977,N_1883);
and U11292 (N_11292,N_1654,N_3021);
and U11293 (N_11293,N_156,N_5833);
xor U11294 (N_11294,N_5071,N_647);
nand U11295 (N_11295,N_662,N_1291);
nand U11296 (N_11296,N_4965,N_5424);
xnor U11297 (N_11297,N_2838,N_5616);
xnor U11298 (N_11298,N_3809,N_1231);
nand U11299 (N_11299,N_1409,N_3340);
or U11300 (N_11300,N_4600,N_3100);
or U11301 (N_11301,N_5777,N_764);
nor U11302 (N_11302,N_3111,N_1751);
and U11303 (N_11303,N_4657,N_3602);
xor U11304 (N_11304,N_1395,N_1775);
nand U11305 (N_11305,N_4495,N_1116);
and U11306 (N_11306,N_4551,N_1819);
or U11307 (N_11307,N_1014,N_2351);
nand U11308 (N_11308,N_1258,N_3862);
and U11309 (N_11309,N_3579,N_4981);
nand U11310 (N_11310,N_5924,N_1306);
nor U11311 (N_11311,N_1244,N_394);
or U11312 (N_11312,N_3023,N_4176);
or U11313 (N_11313,N_2443,N_4676);
nand U11314 (N_11314,N_6211,N_2243);
nor U11315 (N_11315,N_1733,N_6246);
nor U11316 (N_11316,N_3155,N_3319);
nor U11317 (N_11317,N_681,N_2314);
or U11318 (N_11318,N_1449,N_2814);
and U11319 (N_11319,N_2183,N_3125);
and U11320 (N_11320,N_1338,N_4027);
or U11321 (N_11321,N_1596,N_823);
and U11322 (N_11322,N_3650,N_945);
or U11323 (N_11323,N_3704,N_5035);
nor U11324 (N_11324,N_5135,N_1556);
and U11325 (N_11325,N_908,N_486);
or U11326 (N_11326,N_790,N_1111);
xor U11327 (N_11327,N_1863,N_2575);
or U11328 (N_11328,N_1046,N_2684);
xor U11329 (N_11329,N_4685,N_5446);
and U11330 (N_11330,N_4052,N_5988);
xor U11331 (N_11331,N_1616,N_5262);
nand U11332 (N_11332,N_5096,N_3957);
nor U11333 (N_11333,N_450,N_2078);
or U11334 (N_11334,N_1227,N_1032);
nand U11335 (N_11335,N_2290,N_4499);
nor U11336 (N_11336,N_3811,N_5009);
xnor U11337 (N_11337,N_3802,N_2847);
and U11338 (N_11338,N_578,N_215);
xor U11339 (N_11339,N_5929,N_3835);
nor U11340 (N_11340,N_5361,N_2624);
xnor U11341 (N_11341,N_3322,N_922);
nor U11342 (N_11342,N_1529,N_3236);
nand U11343 (N_11343,N_1111,N_3456);
and U11344 (N_11344,N_5817,N_1493);
nand U11345 (N_11345,N_2740,N_4270);
and U11346 (N_11346,N_1095,N_5231);
and U11347 (N_11347,N_3042,N_700);
nor U11348 (N_11348,N_2994,N_3147);
xnor U11349 (N_11349,N_2172,N_1112);
and U11350 (N_11350,N_415,N_1130);
xnor U11351 (N_11351,N_2573,N_3990);
or U11352 (N_11352,N_1586,N_4402);
xor U11353 (N_11353,N_503,N_1712);
nor U11354 (N_11354,N_2,N_2490);
nor U11355 (N_11355,N_2824,N_3482);
nor U11356 (N_11356,N_5331,N_5575);
nand U11357 (N_11357,N_3254,N_6137);
xnor U11358 (N_11358,N_820,N_4928);
or U11359 (N_11359,N_3027,N_5401);
xnor U11360 (N_11360,N_1799,N_2225);
xnor U11361 (N_11361,N_133,N_748);
and U11362 (N_11362,N_2590,N_2230);
xnor U11363 (N_11363,N_1688,N_3912);
and U11364 (N_11364,N_3273,N_1257);
xnor U11365 (N_11365,N_6164,N_2921);
or U11366 (N_11366,N_3674,N_366);
nand U11367 (N_11367,N_5514,N_4757);
and U11368 (N_11368,N_2061,N_335);
or U11369 (N_11369,N_4051,N_5086);
or U11370 (N_11370,N_3423,N_5520);
nand U11371 (N_11371,N_5117,N_4664);
nand U11372 (N_11372,N_3820,N_4834);
nand U11373 (N_11373,N_811,N_5611);
and U11374 (N_11374,N_720,N_1688);
or U11375 (N_11375,N_1119,N_86);
or U11376 (N_11376,N_3206,N_3633);
xor U11377 (N_11377,N_1212,N_552);
nand U11378 (N_11378,N_3090,N_833);
xor U11379 (N_11379,N_1884,N_18);
nor U11380 (N_11380,N_3909,N_3328);
and U11381 (N_11381,N_687,N_5051);
nand U11382 (N_11382,N_979,N_2806);
xor U11383 (N_11383,N_4366,N_5957);
or U11384 (N_11384,N_1537,N_1752);
nor U11385 (N_11385,N_1455,N_2677);
xor U11386 (N_11386,N_4819,N_3654);
nor U11387 (N_11387,N_4078,N_2839);
xor U11388 (N_11388,N_4860,N_3040);
nor U11389 (N_11389,N_1113,N_1269);
or U11390 (N_11390,N_5093,N_1273);
xor U11391 (N_11391,N_2336,N_1386);
xnor U11392 (N_11392,N_2012,N_2387);
or U11393 (N_11393,N_2904,N_5006);
and U11394 (N_11394,N_4957,N_1845);
or U11395 (N_11395,N_5234,N_257);
nand U11396 (N_11396,N_3938,N_413);
xnor U11397 (N_11397,N_5813,N_5388);
nor U11398 (N_11398,N_2434,N_4231);
or U11399 (N_11399,N_4208,N_3915);
xnor U11400 (N_11400,N_4899,N_6113);
nor U11401 (N_11401,N_5609,N_1453);
nand U11402 (N_11402,N_3237,N_2898);
nor U11403 (N_11403,N_3643,N_4023);
xnor U11404 (N_11404,N_4055,N_1510);
nand U11405 (N_11405,N_6241,N_5902);
nand U11406 (N_11406,N_4388,N_4525);
and U11407 (N_11407,N_5424,N_4819);
or U11408 (N_11408,N_5513,N_6175);
xnor U11409 (N_11409,N_2612,N_338);
or U11410 (N_11410,N_1070,N_1507);
xnor U11411 (N_11411,N_3229,N_5916);
and U11412 (N_11412,N_703,N_6138);
nor U11413 (N_11413,N_3238,N_798);
nand U11414 (N_11414,N_4828,N_5676);
xor U11415 (N_11415,N_2894,N_1731);
nand U11416 (N_11416,N_2289,N_596);
or U11417 (N_11417,N_2830,N_3745);
nor U11418 (N_11418,N_1309,N_4227);
xnor U11419 (N_11419,N_3723,N_5351);
nand U11420 (N_11420,N_6199,N_6230);
or U11421 (N_11421,N_5030,N_2811);
nand U11422 (N_11422,N_5457,N_2931);
nor U11423 (N_11423,N_469,N_200);
xor U11424 (N_11424,N_5478,N_723);
and U11425 (N_11425,N_2990,N_6178);
or U11426 (N_11426,N_3309,N_613);
nand U11427 (N_11427,N_5423,N_2597);
and U11428 (N_11428,N_5515,N_2899);
xor U11429 (N_11429,N_3182,N_5265);
nand U11430 (N_11430,N_4766,N_2366);
xor U11431 (N_11431,N_5941,N_5918);
nor U11432 (N_11432,N_5201,N_4377);
nand U11433 (N_11433,N_213,N_5052);
and U11434 (N_11434,N_5315,N_1622);
and U11435 (N_11435,N_6236,N_5097);
xnor U11436 (N_11436,N_249,N_5355);
or U11437 (N_11437,N_1379,N_3828);
nor U11438 (N_11438,N_2022,N_3881);
xnor U11439 (N_11439,N_6117,N_5284);
xor U11440 (N_11440,N_455,N_5382);
nand U11441 (N_11441,N_2545,N_5676);
or U11442 (N_11442,N_5513,N_2305);
nand U11443 (N_11443,N_2143,N_85);
or U11444 (N_11444,N_4937,N_5740);
nor U11445 (N_11445,N_598,N_3348);
nor U11446 (N_11446,N_3740,N_3124);
nand U11447 (N_11447,N_167,N_1512);
and U11448 (N_11448,N_6052,N_5008);
or U11449 (N_11449,N_4025,N_5392);
xnor U11450 (N_11450,N_4402,N_4826);
and U11451 (N_11451,N_3100,N_6009);
or U11452 (N_11452,N_2126,N_5022);
and U11453 (N_11453,N_250,N_5474);
or U11454 (N_11454,N_4215,N_953);
xnor U11455 (N_11455,N_5850,N_4620);
nand U11456 (N_11456,N_2910,N_3771);
nand U11457 (N_11457,N_5729,N_2112);
xor U11458 (N_11458,N_2666,N_5933);
or U11459 (N_11459,N_2643,N_1810);
xor U11460 (N_11460,N_4209,N_2815);
nand U11461 (N_11461,N_2217,N_5142);
xnor U11462 (N_11462,N_2269,N_1649);
nor U11463 (N_11463,N_1990,N_302);
xor U11464 (N_11464,N_4399,N_4478);
xnor U11465 (N_11465,N_774,N_5279);
or U11466 (N_11466,N_5774,N_292);
and U11467 (N_11467,N_4470,N_3712);
or U11468 (N_11468,N_4767,N_5664);
nor U11469 (N_11469,N_4937,N_5244);
nor U11470 (N_11470,N_490,N_5770);
nand U11471 (N_11471,N_2381,N_2462);
nand U11472 (N_11472,N_3661,N_2508);
or U11473 (N_11473,N_2752,N_624);
nor U11474 (N_11474,N_6241,N_2674);
nand U11475 (N_11475,N_2998,N_5097);
and U11476 (N_11476,N_2197,N_5810);
or U11477 (N_11477,N_4810,N_4057);
nand U11478 (N_11478,N_428,N_4283);
nand U11479 (N_11479,N_556,N_3747);
and U11480 (N_11480,N_2912,N_538);
xnor U11481 (N_11481,N_1481,N_3170);
nor U11482 (N_11482,N_4851,N_1542);
xor U11483 (N_11483,N_5188,N_5100);
xnor U11484 (N_11484,N_4161,N_4656);
or U11485 (N_11485,N_1571,N_2486);
nand U11486 (N_11486,N_3305,N_2067);
nand U11487 (N_11487,N_1373,N_765);
and U11488 (N_11488,N_4826,N_3068);
nor U11489 (N_11489,N_5219,N_3834);
xnor U11490 (N_11490,N_1041,N_1537);
and U11491 (N_11491,N_4123,N_2049);
nand U11492 (N_11492,N_534,N_5979);
nand U11493 (N_11493,N_2841,N_215);
and U11494 (N_11494,N_1134,N_6064);
nand U11495 (N_11495,N_5410,N_138);
nand U11496 (N_11496,N_1758,N_6230);
and U11497 (N_11497,N_5058,N_5509);
nand U11498 (N_11498,N_4624,N_420);
or U11499 (N_11499,N_3570,N_334);
and U11500 (N_11500,N_1797,N_258);
nand U11501 (N_11501,N_1019,N_6011);
or U11502 (N_11502,N_5438,N_5915);
xor U11503 (N_11503,N_1829,N_588);
xnor U11504 (N_11504,N_144,N_5319);
or U11505 (N_11505,N_4254,N_5706);
nand U11506 (N_11506,N_3128,N_92);
xnor U11507 (N_11507,N_5088,N_2418);
xor U11508 (N_11508,N_2467,N_3501);
xor U11509 (N_11509,N_3472,N_3912);
and U11510 (N_11510,N_3991,N_3031);
xnor U11511 (N_11511,N_530,N_754);
xnor U11512 (N_11512,N_3719,N_5603);
or U11513 (N_11513,N_1684,N_1888);
nor U11514 (N_11514,N_4408,N_1802);
xnor U11515 (N_11515,N_2600,N_4378);
nor U11516 (N_11516,N_2219,N_3952);
nor U11517 (N_11517,N_1260,N_2608);
nand U11518 (N_11518,N_4226,N_5655);
xnor U11519 (N_11519,N_1539,N_3829);
nor U11520 (N_11520,N_462,N_1119);
and U11521 (N_11521,N_4771,N_4229);
or U11522 (N_11522,N_1720,N_857);
or U11523 (N_11523,N_2848,N_179);
nand U11524 (N_11524,N_3882,N_633);
nand U11525 (N_11525,N_3563,N_5528);
or U11526 (N_11526,N_5027,N_5327);
and U11527 (N_11527,N_1097,N_3049);
or U11528 (N_11528,N_1796,N_3401);
and U11529 (N_11529,N_2505,N_1603);
nand U11530 (N_11530,N_1516,N_2140);
or U11531 (N_11531,N_2401,N_2321);
xor U11532 (N_11532,N_3441,N_2895);
xnor U11533 (N_11533,N_2292,N_2868);
or U11534 (N_11534,N_299,N_2132);
or U11535 (N_11535,N_275,N_45);
and U11536 (N_11536,N_131,N_2337);
nand U11537 (N_11537,N_949,N_3973);
and U11538 (N_11538,N_4145,N_1294);
nor U11539 (N_11539,N_3616,N_5141);
xnor U11540 (N_11540,N_5342,N_4772);
nand U11541 (N_11541,N_606,N_5177);
or U11542 (N_11542,N_3149,N_1301);
xor U11543 (N_11543,N_3245,N_499);
or U11544 (N_11544,N_6038,N_3847);
and U11545 (N_11545,N_3852,N_6052);
nand U11546 (N_11546,N_103,N_2984);
nand U11547 (N_11547,N_1193,N_3728);
nor U11548 (N_11548,N_5376,N_6118);
and U11549 (N_11549,N_4134,N_3530);
nand U11550 (N_11550,N_4749,N_351);
and U11551 (N_11551,N_2015,N_93);
xor U11552 (N_11552,N_2408,N_3741);
xor U11553 (N_11553,N_1711,N_2716);
nor U11554 (N_11554,N_819,N_5412);
nand U11555 (N_11555,N_5611,N_3104);
and U11556 (N_11556,N_5291,N_5483);
and U11557 (N_11557,N_2964,N_1581);
nand U11558 (N_11558,N_537,N_5280);
or U11559 (N_11559,N_5308,N_4841);
and U11560 (N_11560,N_5367,N_1357);
and U11561 (N_11561,N_3684,N_3290);
nand U11562 (N_11562,N_6217,N_5225);
nor U11563 (N_11563,N_750,N_2378);
or U11564 (N_11564,N_2497,N_2315);
or U11565 (N_11565,N_5140,N_3008);
nand U11566 (N_11566,N_2931,N_4708);
nor U11567 (N_11567,N_5595,N_2834);
nand U11568 (N_11568,N_423,N_21);
or U11569 (N_11569,N_358,N_5124);
xor U11570 (N_11570,N_5783,N_2824);
xor U11571 (N_11571,N_4864,N_5315);
or U11572 (N_11572,N_1789,N_820);
or U11573 (N_11573,N_2832,N_1000);
and U11574 (N_11574,N_1390,N_5308);
xnor U11575 (N_11575,N_316,N_3610);
xnor U11576 (N_11576,N_5479,N_2541);
xnor U11577 (N_11577,N_1111,N_1581);
or U11578 (N_11578,N_1013,N_748);
or U11579 (N_11579,N_5743,N_3654);
xor U11580 (N_11580,N_1821,N_4133);
nor U11581 (N_11581,N_5435,N_2329);
nor U11582 (N_11582,N_2445,N_1847);
nor U11583 (N_11583,N_1257,N_4918);
nand U11584 (N_11584,N_2516,N_3895);
nor U11585 (N_11585,N_46,N_3649);
nor U11586 (N_11586,N_554,N_5293);
or U11587 (N_11587,N_3114,N_384);
xnor U11588 (N_11588,N_4611,N_4923);
xnor U11589 (N_11589,N_3154,N_2339);
or U11590 (N_11590,N_3591,N_5961);
and U11591 (N_11591,N_1286,N_1925);
or U11592 (N_11592,N_2874,N_3434);
and U11593 (N_11593,N_1939,N_3809);
nor U11594 (N_11594,N_2115,N_1192);
and U11595 (N_11595,N_3622,N_1121);
or U11596 (N_11596,N_5219,N_2096);
and U11597 (N_11597,N_1433,N_1424);
nor U11598 (N_11598,N_2644,N_4511);
or U11599 (N_11599,N_5773,N_807);
nand U11600 (N_11600,N_5034,N_5739);
nor U11601 (N_11601,N_6050,N_3015);
and U11602 (N_11602,N_2440,N_5386);
and U11603 (N_11603,N_5800,N_57);
or U11604 (N_11604,N_3738,N_3718);
and U11605 (N_11605,N_3258,N_2992);
and U11606 (N_11606,N_3809,N_3268);
and U11607 (N_11607,N_1251,N_1930);
and U11608 (N_11608,N_3783,N_4765);
or U11609 (N_11609,N_2643,N_3619);
and U11610 (N_11610,N_3463,N_638);
or U11611 (N_11611,N_2572,N_6069);
nor U11612 (N_11612,N_829,N_4709);
and U11613 (N_11613,N_4863,N_3687);
nand U11614 (N_11614,N_528,N_3105);
xor U11615 (N_11615,N_1338,N_6067);
and U11616 (N_11616,N_1341,N_1643);
nand U11617 (N_11617,N_2248,N_2293);
or U11618 (N_11618,N_5197,N_6173);
nand U11619 (N_11619,N_2170,N_6052);
xor U11620 (N_11620,N_4643,N_1613);
nand U11621 (N_11621,N_1330,N_2454);
nor U11622 (N_11622,N_4172,N_5686);
xnor U11623 (N_11623,N_3866,N_4422);
nand U11624 (N_11624,N_2937,N_3450);
or U11625 (N_11625,N_2745,N_2998);
nand U11626 (N_11626,N_3224,N_4139);
xor U11627 (N_11627,N_4251,N_5326);
or U11628 (N_11628,N_4013,N_2509);
nand U11629 (N_11629,N_540,N_2361);
xnor U11630 (N_11630,N_5884,N_5144);
xor U11631 (N_11631,N_890,N_4680);
xor U11632 (N_11632,N_2191,N_5840);
and U11633 (N_11633,N_4737,N_780);
and U11634 (N_11634,N_4678,N_1649);
and U11635 (N_11635,N_1120,N_3238);
nand U11636 (N_11636,N_2279,N_2780);
xnor U11637 (N_11637,N_3377,N_560);
and U11638 (N_11638,N_974,N_2627);
xor U11639 (N_11639,N_5481,N_2107);
and U11640 (N_11640,N_3970,N_2816);
and U11641 (N_11641,N_5607,N_5367);
nand U11642 (N_11642,N_5250,N_4708);
and U11643 (N_11643,N_4520,N_5389);
nand U11644 (N_11644,N_4025,N_4815);
and U11645 (N_11645,N_4423,N_671);
and U11646 (N_11646,N_1627,N_875);
nand U11647 (N_11647,N_4498,N_5885);
nor U11648 (N_11648,N_2134,N_2335);
nand U11649 (N_11649,N_4584,N_5165);
or U11650 (N_11650,N_5924,N_5649);
xnor U11651 (N_11651,N_1698,N_399);
or U11652 (N_11652,N_1244,N_5792);
xnor U11653 (N_11653,N_4039,N_373);
and U11654 (N_11654,N_2182,N_4513);
nor U11655 (N_11655,N_2592,N_3958);
or U11656 (N_11656,N_5031,N_2254);
or U11657 (N_11657,N_5365,N_1942);
xor U11658 (N_11658,N_6209,N_2482);
nand U11659 (N_11659,N_5410,N_533);
xnor U11660 (N_11660,N_4087,N_1673);
nand U11661 (N_11661,N_2939,N_202);
or U11662 (N_11662,N_290,N_2386);
xor U11663 (N_11663,N_525,N_3288);
or U11664 (N_11664,N_5583,N_3589);
or U11665 (N_11665,N_4937,N_5632);
or U11666 (N_11666,N_5474,N_420);
or U11667 (N_11667,N_3269,N_3011);
xor U11668 (N_11668,N_5661,N_6049);
xnor U11669 (N_11669,N_2316,N_6219);
and U11670 (N_11670,N_54,N_275);
or U11671 (N_11671,N_4654,N_5581);
nand U11672 (N_11672,N_4424,N_4360);
xor U11673 (N_11673,N_5781,N_2105);
and U11674 (N_11674,N_1156,N_5603);
nand U11675 (N_11675,N_5199,N_4717);
nand U11676 (N_11676,N_453,N_2462);
nand U11677 (N_11677,N_3324,N_5654);
nor U11678 (N_11678,N_5256,N_4563);
and U11679 (N_11679,N_3156,N_4948);
nor U11680 (N_11680,N_2440,N_1511);
nor U11681 (N_11681,N_4704,N_4754);
nor U11682 (N_11682,N_2295,N_9);
and U11683 (N_11683,N_2070,N_3261);
and U11684 (N_11684,N_1328,N_5131);
and U11685 (N_11685,N_460,N_2749);
or U11686 (N_11686,N_4993,N_3723);
and U11687 (N_11687,N_4401,N_5131);
xnor U11688 (N_11688,N_2747,N_4590);
nor U11689 (N_11689,N_571,N_707);
xor U11690 (N_11690,N_4397,N_1574);
xnor U11691 (N_11691,N_4413,N_1667);
and U11692 (N_11692,N_2479,N_927);
nor U11693 (N_11693,N_5906,N_4505);
or U11694 (N_11694,N_949,N_759);
nand U11695 (N_11695,N_5398,N_3695);
nor U11696 (N_11696,N_954,N_4574);
or U11697 (N_11697,N_3297,N_447);
xor U11698 (N_11698,N_982,N_3689);
and U11699 (N_11699,N_4570,N_2634);
xor U11700 (N_11700,N_4414,N_5378);
or U11701 (N_11701,N_2498,N_1029);
nand U11702 (N_11702,N_2215,N_3882);
xor U11703 (N_11703,N_1085,N_3729);
and U11704 (N_11704,N_6131,N_1743);
or U11705 (N_11705,N_4432,N_2595);
or U11706 (N_11706,N_2149,N_144);
nand U11707 (N_11707,N_5316,N_566);
xnor U11708 (N_11708,N_4520,N_2139);
xnor U11709 (N_11709,N_2355,N_2154);
nor U11710 (N_11710,N_2266,N_3298);
and U11711 (N_11711,N_2080,N_3344);
or U11712 (N_11712,N_3724,N_2280);
nor U11713 (N_11713,N_2042,N_3577);
nand U11714 (N_11714,N_487,N_5787);
or U11715 (N_11715,N_5235,N_3875);
xor U11716 (N_11716,N_1738,N_1);
nor U11717 (N_11717,N_4906,N_5491);
or U11718 (N_11718,N_4289,N_524);
nand U11719 (N_11719,N_978,N_997);
nand U11720 (N_11720,N_5319,N_3630);
and U11721 (N_11721,N_462,N_5635);
nor U11722 (N_11722,N_336,N_1893);
nand U11723 (N_11723,N_5780,N_4893);
xor U11724 (N_11724,N_4228,N_4299);
xnor U11725 (N_11725,N_1699,N_3270);
or U11726 (N_11726,N_6058,N_3247);
nand U11727 (N_11727,N_861,N_326);
and U11728 (N_11728,N_5427,N_5016);
nor U11729 (N_11729,N_2397,N_3737);
nor U11730 (N_11730,N_6113,N_2805);
xnor U11731 (N_11731,N_3182,N_3736);
or U11732 (N_11732,N_4448,N_3827);
and U11733 (N_11733,N_3739,N_5521);
xnor U11734 (N_11734,N_2731,N_1334);
nor U11735 (N_11735,N_993,N_4271);
nand U11736 (N_11736,N_1338,N_3995);
nand U11737 (N_11737,N_3042,N_5621);
and U11738 (N_11738,N_5261,N_3794);
nand U11739 (N_11739,N_1290,N_1903);
or U11740 (N_11740,N_1979,N_1562);
and U11741 (N_11741,N_348,N_5154);
nor U11742 (N_11742,N_5571,N_3250);
xor U11743 (N_11743,N_492,N_1627);
nor U11744 (N_11744,N_190,N_2474);
xnor U11745 (N_11745,N_4153,N_6070);
or U11746 (N_11746,N_1918,N_1553);
xor U11747 (N_11747,N_3499,N_2614);
or U11748 (N_11748,N_2711,N_5315);
nor U11749 (N_11749,N_4462,N_781);
or U11750 (N_11750,N_3994,N_302);
and U11751 (N_11751,N_2656,N_604);
nand U11752 (N_11752,N_5252,N_598);
or U11753 (N_11753,N_3169,N_4553);
xnor U11754 (N_11754,N_2945,N_5851);
and U11755 (N_11755,N_4336,N_5185);
nor U11756 (N_11756,N_418,N_38);
nor U11757 (N_11757,N_5642,N_1077);
xnor U11758 (N_11758,N_4863,N_4771);
nor U11759 (N_11759,N_2529,N_2951);
or U11760 (N_11760,N_1404,N_6093);
xnor U11761 (N_11761,N_1751,N_5414);
and U11762 (N_11762,N_3744,N_1534);
xnor U11763 (N_11763,N_2747,N_1666);
or U11764 (N_11764,N_371,N_1354);
nand U11765 (N_11765,N_1391,N_240);
nand U11766 (N_11766,N_340,N_1875);
or U11767 (N_11767,N_1470,N_356);
xnor U11768 (N_11768,N_457,N_2131);
nand U11769 (N_11769,N_5483,N_20);
and U11770 (N_11770,N_3373,N_5781);
and U11771 (N_11771,N_3734,N_4102);
or U11772 (N_11772,N_2388,N_1913);
nor U11773 (N_11773,N_5844,N_4460);
or U11774 (N_11774,N_3515,N_5020);
nor U11775 (N_11775,N_2907,N_3925);
nand U11776 (N_11776,N_1220,N_4549);
nand U11777 (N_11777,N_4637,N_4241);
xor U11778 (N_11778,N_10,N_1245);
xnor U11779 (N_11779,N_5301,N_3163);
xnor U11780 (N_11780,N_406,N_4810);
nand U11781 (N_11781,N_4337,N_4546);
nand U11782 (N_11782,N_2041,N_2115);
or U11783 (N_11783,N_4728,N_3547);
nor U11784 (N_11784,N_526,N_4828);
and U11785 (N_11785,N_3349,N_4955);
xnor U11786 (N_11786,N_5446,N_5597);
xnor U11787 (N_11787,N_2004,N_223);
and U11788 (N_11788,N_3785,N_1373);
nand U11789 (N_11789,N_1411,N_5423);
and U11790 (N_11790,N_4238,N_5935);
nor U11791 (N_11791,N_1875,N_2606);
xnor U11792 (N_11792,N_1147,N_972);
or U11793 (N_11793,N_5878,N_3751);
xnor U11794 (N_11794,N_4480,N_2554);
or U11795 (N_11795,N_5454,N_4455);
nor U11796 (N_11796,N_248,N_3849);
or U11797 (N_11797,N_4536,N_4131);
nor U11798 (N_11798,N_3751,N_1845);
nand U11799 (N_11799,N_3683,N_5175);
nand U11800 (N_11800,N_1278,N_3008);
and U11801 (N_11801,N_2203,N_6023);
nand U11802 (N_11802,N_5034,N_251);
or U11803 (N_11803,N_2753,N_121);
nor U11804 (N_11804,N_1451,N_1050);
nor U11805 (N_11805,N_1987,N_4118);
and U11806 (N_11806,N_2028,N_906);
nor U11807 (N_11807,N_4756,N_577);
nor U11808 (N_11808,N_241,N_440);
nor U11809 (N_11809,N_5226,N_5006);
nor U11810 (N_11810,N_585,N_361);
nand U11811 (N_11811,N_4267,N_5506);
nor U11812 (N_11812,N_1864,N_2692);
and U11813 (N_11813,N_5640,N_423);
and U11814 (N_11814,N_2336,N_214);
nand U11815 (N_11815,N_810,N_1837);
or U11816 (N_11816,N_5247,N_1762);
xor U11817 (N_11817,N_822,N_805);
nor U11818 (N_11818,N_2881,N_4572);
xor U11819 (N_11819,N_5300,N_5363);
and U11820 (N_11820,N_940,N_3736);
or U11821 (N_11821,N_5172,N_3915);
or U11822 (N_11822,N_2575,N_4072);
or U11823 (N_11823,N_3747,N_1624);
xor U11824 (N_11824,N_4810,N_1411);
and U11825 (N_11825,N_1277,N_3772);
nor U11826 (N_11826,N_595,N_6107);
or U11827 (N_11827,N_2661,N_747);
xnor U11828 (N_11828,N_1882,N_3246);
nand U11829 (N_11829,N_1625,N_3759);
nand U11830 (N_11830,N_4641,N_4645);
xor U11831 (N_11831,N_4512,N_400);
or U11832 (N_11832,N_979,N_4158);
or U11833 (N_11833,N_4285,N_3808);
nand U11834 (N_11834,N_4367,N_1688);
or U11835 (N_11835,N_4513,N_2439);
nand U11836 (N_11836,N_5353,N_751);
xnor U11837 (N_11837,N_4920,N_5330);
or U11838 (N_11838,N_164,N_1507);
nor U11839 (N_11839,N_4174,N_6153);
and U11840 (N_11840,N_3919,N_67);
nor U11841 (N_11841,N_37,N_1574);
nor U11842 (N_11842,N_528,N_2302);
nand U11843 (N_11843,N_3350,N_2074);
xor U11844 (N_11844,N_4832,N_4426);
or U11845 (N_11845,N_3925,N_2943);
nand U11846 (N_11846,N_4266,N_1967);
xnor U11847 (N_11847,N_4896,N_4472);
and U11848 (N_11848,N_5819,N_1147);
nor U11849 (N_11849,N_1339,N_2009);
and U11850 (N_11850,N_4156,N_4655);
nor U11851 (N_11851,N_267,N_5146);
nand U11852 (N_11852,N_2434,N_1237);
or U11853 (N_11853,N_180,N_5688);
and U11854 (N_11854,N_4754,N_90);
nand U11855 (N_11855,N_1212,N_525);
or U11856 (N_11856,N_2468,N_4816);
and U11857 (N_11857,N_4663,N_1751);
or U11858 (N_11858,N_5819,N_1301);
nand U11859 (N_11859,N_4200,N_2342);
or U11860 (N_11860,N_4447,N_2395);
nand U11861 (N_11861,N_3941,N_582);
or U11862 (N_11862,N_3540,N_4431);
or U11863 (N_11863,N_5866,N_5840);
nand U11864 (N_11864,N_2575,N_5060);
xnor U11865 (N_11865,N_3963,N_4618);
and U11866 (N_11866,N_5063,N_2212);
nor U11867 (N_11867,N_3547,N_6183);
or U11868 (N_11868,N_5908,N_2397);
and U11869 (N_11869,N_2427,N_3023);
nor U11870 (N_11870,N_755,N_6092);
or U11871 (N_11871,N_2602,N_1929);
or U11872 (N_11872,N_5536,N_3682);
xor U11873 (N_11873,N_2676,N_5957);
nor U11874 (N_11874,N_2190,N_3584);
nand U11875 (N_11875,N_3254,N_5096);
and U11876 (N_11876,N_5302,N_6221);
xnor U11877 (N_11877,N_5732,N_4866);
nor U11878 (N_11878,N_4715,N_404);
nand U11879 (N_11879,N_6208,N_2506);
and U11880 (N_11880,N_794,N_1870);
nor U11881 (N_11881,N_3725,N_4143);
xor U11882 (N_11882,N_3651,N_3950);
nand U11883 (N_11883,N_5514,N_4230);
and U11884 (N_11884,N_1735,N_2346);
or U11885 (N_11885,N_4139,N_2648);
xor U11886 (N_11886,N_1984,N_4267);
xor U11887 (N_11887,N_2388,N_2500);
and U11888 (N_11888,N_5997,N_2751);
nand U11889 (N_11889,N_6242,N_1978);
xnor U11890 (N_11890,N_5575,N_4139);
xnor U11891 (N_11891,N_6227,N_3770);
and U11892 (N_11892,N_1450,N_1462);
and U11893 (N_11893,N_4111,N_4424);
and U11894 (N_11894,N_4062,N_2846);
xor U11895 (N_11895,N_1887,N_2073);
nand U11896 (N_11896,N_1739,N_2432);
and U11897 (N_11897,N_2773,N_4277);
nor U11898 (N_11898,N_5253,N_2299);
nor U11899 (N_11899,N_5960,N_2627);
or U11900 (N_11900,N_1094,N_5680);
nor U11901 (N_11901,N_2736,N_3898);
nand U11902 (N_11902,N_4225,N_4166);
xor U11903 (N_11903,N_4424,N_1847);
xnor U11904 (N_11904,N_2561,N_657);
xor U11905 (N_11905,N_2152,N_5867);
nor U11906 (N_11906,N_1442,N_627);
nand U11907 (N_11907,N_3,N_4638);
or U11908 (N_11908,N_6152,N_4340);
xnor U11909 (N_11909,N_1368,N_5322);
xor U11910 (N_11910,N_5130,N_2068);
xnor U11911 (N_11911,N_1681,N_4022);
xor U11912 (N_11912,N_1254,N_5551);
and U11913 (N_11913,N_482,N_3415);
and U11914 (N_11914,N_4260,N_4750);
xor U11915 (N_11915,N_887,N_4158);
and U11916 (N_11916,N_2991,N_752);
and U11917 (N_11917,N_2224,N_1642);
nor U11918 (N_11918,N_1001,N_2951);
nor U11919 (N_11919,N_1891,N_1308);
nand U11920 (N_11920,N_2041,N_4110);
xnor U11921 (N_11921,N_3226,N_605);
nor U11922 (N_11922,N_5041,N_4527);
xnor U11923 (N_11923,N_2588,N_1548);
nor U11924 (N_11924,N_1308,N_1367);
nor U11925 (N_11925,N_2005,N_2828);
and U11926 (N_11926,N_3697,N_3506);
or U11927 (N_11927,N_1385,N_3600);
xnor U11928 (N_11928,N_1551,N_2847);
or U11929 (N_11929,N_578,N_5810);
and U11930 (N_11930,N_5025,N_3432);
and U11931 (N_11931,N_3147,N_2129);
or U11932 (N_11932,N_1804,N_2864);
nand U11933 (N_11933,N_5941,N_2957);
nand U11934 (N_11934,N_5306,N_4906);
nor U11935 (N_11935,N_4182,N_341);
or U11936 (N_11936,N_3257,N_5899);
nand U11937 (N_11937,N_254,N_3454);
nor U11938 (N_11938,N_1940,N_529);
and U11939 (N_11939,N_3772,N_117);
or U11940 (N_11940,N_5194,N_3649);
or U11941 (N_11941,N_1774,N_1631);
xnor U11942 (N_11942,N_4348,N_752);
or U11943 (N_11943,N_2960,N_1984);
nor U11944 (N_11944,N_3094,N_5155);
nand U11945 (N_11945,N_3423,N_1046);
nand U11946 (N_11946,N_292,N_3626);
nand U11947 (N_11947,N_4995,N_1894);
and U11948 (N_11948,N_3034,N_6082);
xor U11949 (N_11949,N_2661,N_4074);
nor U11950 (N_11950,N_5116,N_597);
nor U11951 (N_11951,N_5721,N_5493);
or U11952 (N_11952,N_1112,N_2592);
or U11953 (N_11953,N_3330,N_1775);
xnor U11954 (N_11954,N_188,N_3791);
xor U11955 (N_11955,N_3344,N_3836);
or U11956 (N_11956,N_5127,N_991);
and U11957 (N_11957,N_441,N_5774);
nor U11958 (N_11958,N_5484,N_3914);
nand U11959 (N_11959,N_2669,N_5220);
nor U11960 (N_11960,N_6023,N_3938);
or U11961 (N_11961,N_1485,N_2573);
nor U11962 (N_11962,N_1578,N_5644);
nand U11963 (N_11963,N_2651,N_6213);
or U11964 (N_11964,N_759,N_1595);
or U11965 (N_11965,N_1128,N_5716);
or U11966 (N_11966,N_237,N_5032);
nand U11967 (N_11967,N_4977,N_4110);
or U11968 (N_11968,N_133,N_5918);
nor U11969 (N_11969,N_771,N_448);
and U11970 (N_11970,N_6005,N_548);
nor U11971 (N_11971,N_2717,N_5714);
or U11972 (N_11972,N_5943,N_3162);
or U11973 (N_11973,N_1393,N_5525);
nand U11974 (N_11974,N_482,N_1365);
and U11975 (N_11975,N_1217,N_6113);
and U11976 (N_11976,N_308,N_4026);
xor U11977 (N_11977,N_1014,N_3890);
xnor U11978 (N_11978,N_493,N_4811);
and U11979 (N_11979,N_5694,N_4380);
and U11980 (N_11980,N_3248,N_5121);
nor U11981 (N_11981,N_3053,N_779);
xnor U11982 (N_11982,N_1499,N_1644);
nor U11983 (N_11983,N_677,N_2651);
and U11984 (N_11984,N_88,N_163);
or U11985 (N_11985,N_2176,N_272);
nand U11986 (N_11986,N_5757,N_3621);
nor U11987 (N_11987,N_3045,N_2371);
nor U11988 (N_11988,N_2750,N_310);
or U11989 (N_11989,N_1955,N_6105);
nor U11990 (N_11990,N_4014,N_3510);
nor U11991 (N_11991,N_1345,N_545);
nand U11992 (N_11992,N_1394,N_5248);
xor U11993 (N_11993,N_2137,N_6000);
or U11994 (N_11994,N_3734,N_3274);
nor U11995 (N_11995,N_2482,N_1508);
xnor U11996 (N_11996,N_820,N_3120);
nand U11997 (N_11997,N_3669,N_196);
and U11998 (N_11998,N_4666,N_957);
and U11999 (N_11999,N_3555,N_4156);
and U12000 (N_12000,N_4222,N_4841);
xnor U12001 (N_12001,N_227,N_3133);
xnor U12002 (N_12002,N_4391,N_584);
nor U12003 (N_12003,N_3404,N_5117);
xnor U12004 (N_12004,N_5724,N_2481);
nand U12005 (N_12005,N_1211,N_4484);
nor U12006 (N_12006,N_227,N_5747);
and U12007 (N_12007,N_4436,N_3343);
nor U12008 (N_12008,N_2956,N_5232);
xor U12009 (N_12009,N_3798,N_38);
xor U12010 (N_12010,N_1866,N_2836);
or U12011 (N_12011,N_4290,N_202);
xor U12012 (N_12012,N_5164,N_401);
xor U12013 (N_12013,N_2402,N_4155);
or U12014 (N_12014,N_2422,N_1112);
and U12015 (N_12015,N_2604,N_3459);
nand U12016 (N_12016,N_739,N_1522);
and U12017 (N_12017,N_147,N_5076);
nand U12018 (N_12018,N_4544,N_2295);
nor U12019 (N_12019,N_5460,N_999);
nor U12020 (N_12020,N_2814,N_2671);
xnor U12021 (N_12021,N_3224,N_4560);
or U12022 (N_12022,N_5816,N_4457);
nand U12023 (N_12023,N_4099,N_2139);
and U12024 (N_12024,N_4445,N_5901);
and U12025 (N_12025,N_2107,N_1145);
nand U12026 (N_12026,N_1716,N_2350);
nor U12027 (N_12027,N_2692,N_2218);
nor U12028 (N_12028,N_4645,N_6041);
nand U12029 (N_12029,N_5399,N_5050);
or U12030 (N_12030,N_3844,N_5217);
or U12031 (N_12031,N_561,N_3873);
xnor U12032 (N_12032,N_4695,N_5306);
nand U12033 (N_12033,N_104,N_1993);
nand U12034 (N_12034,N_2959,N_3836);
nand U12035 (N_12035,N_5332,N_5608);
and U12036 (N_12036,N_2118,N_4763);
xor U12037 (N_12037,N_18,N_2712);
nor U12038 (N_12038,N_1407,N_883);
nor U12039 (N_12039,N_548,N_234);
and U12040 (N_12040,N_3966,N_4169);
xor U12041 (N_12041,N_454,N_5788);
or U12042 (N_12042,N_282,N_4313);
and U12043 (N_12043,N_945,N_5768);
nand U12044 (N_12044,N_889,N_2000);
xnor U12045 (N_12045,N_1921,N_4361);
and U12046 (N_12046,N_1749,N_2165);
or U12047 (N_12047,N_1870,N_5350);
or U12048 (N_12048,N_330,N_2150);
or U12049 (N_12049,N_1467,N_1722);
or U12050 (N_12050,N_4377,N_3444);
or U12051 (N_12051,N_2877,N_2448);
and U12052 (N_12052,N_2028,N_1);
nor U12053 (N_12053,N_4142,N_2532);
or U12054 (N_12054,N_1668,N_6127);
nor U12055 (N_12055,N_3122,N_5274);
nor U12056 (N_12056,N_2222,N_2389);
or U12057 (N_12057,N_4959,N_4416);
and U12058 (N_12058,N_2677,N_1896);
or U12059 (N_12059,N_4342,N_995);
or U12060 (N_12060,N_2563,N_5778);
and U12061 (N_12061,N_3267,N_519);
nand U12062 (N_12062,N_1673,N_3451);
nand U12063 (N_12063,N_5721,N_793);
nand U12064 (N_12064,N_4924,N_156);
nand U12065 (N_12065,N_5178,N_6071);
and U12066 (N_12066,N_6118,N_4309);
or U12067 (N_12067,N_3153,N_6038);
nand U12068 (N_12068,N_2258,N_1548);
and U12069 (N_12069,N_5490,N_6126);
and U12070 (N_12070,N_5331,N_5240);
nand U12071 (N_12071,N_3919,N_4611);
or U12072 (N_12072,N_697,N_6087);
nand U12073 (N_12073,N_6064,N_779);
and U12074 (N_12074,N_5400,N_2677);
xor U12075 (N_12075,N_2649,N_2174);
and U12076 (N_12076,N_978,N_1871);
and U12077 (N_12077,N_2444,N_2121);
nand U12078 (N_12078,N_2086,N_5793);
and U12079 (N_12079,N_3010,N_2334);
nor U12080 (N_12080,N_3970,N_5134);
and U12081 (N_12081,N_1336,N_2470);
nor U12082 (N_12082,N_4196,N_2568);
xnor U12083 (N_12083,N_3403,N_3018);
or U12084 (N_12084,N_5073,N_4531);
xnor U12085 (N_12085,N_368,N_318);
or U12086 (N_12086,N_3534,N_807);
xor U12087 (N_12087,N_3418,N_5966);
nand U12088 (N_12088,N_3167,N_3531);
and U12089 (N_12089,N_4048,N_713);
xnor U12090 (N_12090,N_2883,N_5086);
nand U12091 (N_12091,N_5797,N_4499);
or U12092 (N_12092,N_5430,N_3088);
or U12093 (N_12093,N_6042,N_109);
nand U12094 (N_12094,N_4214,N_4712);
and U12095 (N_12095,N_3727,N_1849);
and U12096 (N_12096,N_3504,N_5667);
or U12097 (N_12097,N_3072,N_2735);
nand U12098 (N_12098,N_4262,N_563);
nand U12099 (N_12099,N_3142,N_2078);
xor U12100 (N_12100,N_5478,N_3849);
and U12101 (N_12101,N_1694,N_6063);
nor U12102 (N_12102,N_5250,N_309);
xor U12103 (N_12103,N_6119,N_5088);
and U12104 (N_12104,N_4471,N_916);
nor U12105 (N_12105,N_4114,N_1139);
and U12106 (N_12106,N_768,N_1060);
nor U12107 (N_12107,N_3227,N_5431);
xnor U12108 (N_12108,N_1446,N_136);
nand U12109 (N_12109,N_5615,N_1281);
xnor U12110 (N_12110,N_5535,N_5103);
nand U12111 (N_12111,N_5996,N_1364);
nor U12112 (N_12112,N_3300,N_857);
and U12113 (N_12113,N_4237,N_1391);
or U12114 (N_12114,N_4354,N_2874);
nand U12115 (N_12115,N_5670,N_3282);
xor U12116 (N_12116,N_5123,N_4364);
and U12117 (N_12117,N_4415,N_4934);
xnor U12118 (N_12118,N_2860,N_4276);
nor U12119 (N_12119,N_4044,N_5045);
nand U12120 (N_12120,N_1597,N_1526);
xnor U12121 (N_12121,N_3975,N_4718);
nor U12122 (N_12122,N_4474,N_5583);
or U12123 (N_12123,N_4555,N_2399);
nor U12124 (N_12124,N_5276,N_3737);
or U12125 (N_12125,N_466,N_2817);
nand U12126 (N_12126,N_5507,N_3479);
nor U12127 (N_12127,N_937,N_989);
or U12128 (N_12128,N_5360,N_2627);
nor U12129 (N_12129,N_3716,N_301);
and U12130 (N_12130,N_2695,N_2088);
nor U12131 (N_12131,N_3400,N_237);
nand U12132 (N_12132,N_5072,N_1879);
xor U12133 (N_12133,N_4121,N_5793);
xnor U12134 (N_12134,N_628,N_2460);
nor U12135 (N_12135,N_2323,N_5376);
nor U12136 (N_12136,N_5024,N_3757);
or U12137 (N_12137,N_2142,N_1314);
or U12138 (N_12138,N_3208,N_3417);
nand U12139 (N_12139,N_6228,N_4291);
nor U12140 (N_12140,N_280,N_555);
nor U12141 (N_12141,N_6212,N_3131);
nand U12142 (N_12142,N_5509,N_2868);
xor U12143 (N_12143,N_5391,N_72);
nor U12144 (N_12144,N_387,N_190);
nand U12145 (N_12145,N_303,N_4162);
nor U12146 (N_12146,N_5579,N_3921);
and U12147 (N_12147,N_4178,N_1403);
nor U12148 (N_12148,N_631,N_1659);
nor U12149 (N_12149,N_2970,N_2906);
nand U12150 (N_12150,N_3647,N_1016);
nand U12151 (N_12151,N_172,N_1534);
nor U12152 (N_12152,N_3137,N_6116);
nor U12153 (N_12153,N_1106,N_1631);
or U12154 (N_12154,N_3021,N_4024);
and U12155 (N_12155,N_1930,N_3456);
nand U12156 (N_12156,N_798,N_4506);
or U12157 (N_12157,N_2484,N_611);
xor U12158 (N_12158,N_836,N_316);
xor U12159 (N_12159,N_1807,N_4673);
and U12160 (N_12160,N_3285,N_5959);
nor U12161 (N_12161,N_2349,N_5915);
and U12162 (N_12162,N_5126,N_5776);
xor U12163 (N_12163,N_1914,N_3449);
xnor U12164 (N_12164,N_2111,N_1086);
and U12165 (N_12165,N_1405,N_4929);
or U12166 (N_12166,N_5560,N_5577);
nor U12167 (N_12167,N_1241,N_0);
or U12168 (N_12168,N_5325,N_4465);
or U12169 (N_12169,N_5644,N_52);
nand U12170 (N_12170,N_579,N_3217);
xnor U12171 (N_12171,N_257,N_5816);
or U12172 (N_12172,N_1776,N_921);
nor U12173 (N_12173,N_4678,N_2525);
nand U12174 (N_12174,N_4981,N_5590);
nand U12175 (N_12175,N_6062,N_4545);
nor U12176 (N_12176,N_3767,N_2791);
and U12177 (N_12177,N_5993,N_89);
xnor U12178 (N_12178,N_3393,N_4778);
nor U12179 (N_12179,N_4043,N_3984);
nor U12180 (N_12180,N_2668,N_841);
xor U12181 (N_12181,N_247,N_5075);
nor U12182 (N_12182,N_3575,N_6030);
or U12183 (N_12183,N_4395,N_1039);
or U12184 (N_12184,N_574,N_2136);
xor U12185 (N_12185,N_4428,N_46);
xor U12186 (N_12186,N_4693,N_4438);
xor U12187 (N_12187,N_6189,N_1220);
nor U12188 (N_12188,N_4428,N_1839);
and U12189 (N_12189,N_2073,N_2536);
nor U12190 (N_12190,N_714,N_2456);
xnor U12191 (N_12191,N_4563,N_4283);
xor U12192 (N_12192,N_3867,N_1861);
nand U12193 (N_12193,N_3182,N_1583);
or U12194 (N_12194,N_5831,N_200);
xor U12195 (N_12195,N_959,N_3845);
nand U12196 (N_12196,N_5044,N_4407);
and U12197 (N_12197,N_5144,N_3784);
xnor U12198 (N_12198,N_1330,N_3254);
or U12199 (N_12199,N_4231,N_324);
and U12200 (N_12200,N_3591,N_3705);
nor U12201 (N_12201,N_6064,N_2389);
and U12202 (N_12202,N_5996,N_3117);
and U12203 (N_12203,N_5912,N_3829);
and U12204 (N_12204,N_6004,N_5928);
nor U12205 (N_12205,N_3721,N_4752);
nor U12206 (N_12206,N_3810,N_3292);
xnor U12207 (N_12207,N_5114,N_1839);
or U12208 (N_12208,N_5544,N_937);
and U12209 (N_12209,N_5518,N_5317);
nor U12210 (N_12210,N_3709,N_3170);
or U12211 (N_12211,N_3372,N_748);
and U12212 (N_12212,N_6081,N_1731);
or U12213 (N_12213,N_4300,N_2238);
nand U12214 (N_12214,N_2078,N_6051);
xnor U12215 (N_12215,N_6238,N_5721);
nand U12216 (N_12216,N_6146,N_5580);
nor U12217 (N_12217,N_1914,N_4978);
and U12218 (N_12218,N_1107,N_4720);
xnor U12219 (N_12219,N_1516,N_1529);
nor U12220 (N_12220,N_5296,N_407);
nand U12221 (N_12221,N_4574,N_4331);
or U12222 (N_12222,N_3691,N_1682);
nand U12223 (N_12223,N_3454,N_3672);
or U12224 (N_12224,N_5279,N_5177);
nor U12225 (N_12225,N_3044,N_1397);
or U12226 (N_12226,N_4910,N_3513);
xnor U12227 (N_12227,N_938,N_1245);
and U12228 (N_12228,N_5440,N_4076);
nor U12229 (N_12229,N_6229,N_2155);
nand U12230 (N_12230,N_1641,N_4665);
or U12231 (N_12231,N_635,N_4980);
xor U12232 (N_12232,N_4693,N_1436);
nand U12233 (N_12233,N_3433,N_4042);
xor U12234 (N_12234,N_3789,N_5485);
or U12235 (N_12235,N_1256,N_5383);
nor U12236 (N_12236,N_5124,N_4361);
nand U12237 (N_12237,N_407,N_3787);
nand U12238 (N_12238,N_993,N_424);
and U12239 (N_12239,N_5717,N_1651);
or U12240 (N_12240,N_1082,N_2962);
and U12241 (N_12241,N_4951,N_5212);
nor U12242 (N_12242,N_5397,N_1464);
or U12243 (N_12243,N_3525,N_4511);
nor U12244 (N_12244,N_5833,N_39);
xnor U12245 (N_12245,N_2632,N_4704);
or U12246 (N_12246,N_1293,N_5159);
nand U12247 (N_12247,N_4707,N_1384);
nand U12248 (N_12248,N_2919,N_2870);
and U12249 (N_12249,N_4661,N_3543);
and U12250 (N_12250,N_6241,N_4134);
xnor U12251 (N_12251,N_2107,N_2923);
or U12252 (N_12252,N_2562,N_148);
nor U12253 (N_12253,N_5350,N_1160);
nand U12254 (N_12254,N_814,N_379);
or U12255 (N_12255,N_2136,N_5711);
nor U12256 (N_12256,N_2962,N_4414);
nand U12257 (N_12257,N_4577,N_5262);
nor U12258 (N_12258,N_3728,N_4829);
or U12259 (N_12259,N_1361,N_1567);
and U12260 (N_12260,N_2500,N_1706);
or U12261 (N_12261,N_5853,N_3990);
and U12262 (N_12262,N_99,N_6102);
or U12263 (N_12263,N_2538,N_595);
nand U12264 (N_12264,N_764,N_469);
nor U12265 (N_12265,N_1928,N_2883);
nand U12266 (N_12266,N_2784,N_440);
or U12267 (N_12267,N_1407,N_3640);
and U12268 (N_12268,N_3192,N_22);
nand U12269 (N_12269,N_3363,N_5461);
nor U12270 (N_12270,N_5320,N_4473);
xor U12271 (N_12271,N_5201,N_404);
nor U12272 (N_12272,N_155,N_5185);
and U12273 (N_12273,N_4014,N_5922);
and U12274 (N_12274,N_2482,N_747);
nor U12275 (N_12275,N_5617,N_4433);
and U12276 (N_12276,N_1736,N_5963);
xnor U12277 (N_12277,N_418,N_5412);
and U12278 (N_12278,N_4391,N_6181);
and U12279 (N_12279,N_1543,N_1738);
nor U12280 (N_12280,N_3722,N_3007);
or U12281 (N_12281,N_5700,N_4380);
or U12282 (N_12282,N_981,N_3093);
or U12283 (N_12283,N_6089,N_2759);
nor U12284 (N_12284,N_1658,N_2540);
xnor U12285 (N_12285,N_3474,N_2345);
or U12286 (N_12286,N_2820,N_2824);
xnor U12287 (N_12287,N_308,N_1392);
nand U12288 (N_12288,N_1656,N_4531);
nor U12289 (N_12289,N_461,N_4767);
nor U12290 (N_12290,N_4814,N_1725);
or U12291 (N_12291,N_3181,N_974);
nand U12292 (N_12292,N_4408,N_1994);
xor U12293 (N_12293,N_3695,N_768);
or U12294 (N_12294,N_1619,N_1882);
nand U12295 (N_12295,N_3453,N_3298);
or U12296 (N_12296,N_4860,N_480);
xor U12297 (N_12297,N_3959,N_4178);
and U12298 (N_12298,N_2711,N_1817);
nor U12299 (N_12299,N_5795,N_410);
or U12300 (N_12300,N_1795,N_2885);
nor U12301 (N_12301,N_5532,N_4008);
and U12302 (N_12302,N_52,N_5024);
nor U12303 (N_12303,N_1777,N_3132);
and U12304 (N_12304,N_4323,N_3760);
and U12305 (N_12305,N_5359,N_5707);
and U12306 (N_12306,N_3673,N_810);
and U12307 (N_12307,N_6096,N_6029);
nand U12308 (N_12308,N_1029,N_1054);
nand U12309 (N_12309,N_986,N_6148);
nor U12310 (N_12310,N_4069,N_3876);
or U12311 (N_12311,N_1879,N_4778);
and U12312 (N_12312,N_958,N_836);
nand U12313 (N_12313,N_2195,N_475);
nand U12314 (N_12314,N_4634,N_1129);
or U12315 (N_12315,N_3426,N_4797);
and U12316 (N_12316,N_1737,N_1849);
nand U12317 (N_12317,N_5147,N_5118);
nor U12318 (N_12318,N_3435,N_1129);
nand U12319 (N_12319,N_3278,N_4116);
xor U12320 (N_12320,N_1849,N_4353);
and U12321 (N_12321,N_5703,N_4123);
or U12322 (N_12322,N_2637,N_3240);
xor U12323 (N_12323,N_2095,N_6045);
xnor U12324 (N_12324,N_1365,N_661);
and U12325 (N_12325,N_1411,N_515);
nor U12326 (N_12326,N_4409,N_2907);
or U12327 (N_12327,N_2892,N_1162);
nor U12328 (N_12328,N_1340,N_1364);
xnor U12329 (N_12329,N_1515,N_4767);
and U12330 (N_12330,N_5574,N_2123);
or U12331 (N_12331,N_3299,N_3016);
and U12332 (N_12332,N_5706,N_3337);
nor U12333 (N_12333,N_3691,N_4918);
or U12334 (N_12334,N_2170,N_1862);
nor U12335 (N_12335,N_5342,N_1843);
xnor U12336 (N_12336,N_5992,N_2650);
xor U12337 (N_12337,N_3182,N_3142);
xnor U12338 (N_12338,N_1599,N_2879);
and U12339 (N_12339,N_4823,N_2173);
nand U12340 (N_12340,N_434,N_4115);
xnor U12341 (N_12341,N_2650,N_3389);
xnor U12342 (N_12342,N_1449,N_5301);
or U12343 (N_12343,N_4040,N_5338);
nand U12344 (N_12344,N_219,N_3854);
xnor U12345 (N_12345,N_5079,N_5850);
nand U12346 (N_12346,N_1842,N_1404);
nand U12347 (N_12347,N_531,N_4391);
or U12348 (N_12348,N_1187,N_173);
nor U12349 (N_12349,N_3909,N_5405);
nand U12350 (N_12350,N_1763,N_6220);
nor U12351 (N_12351,N_2135,N_6165);
nand U12352 (N_12352,N_1459,N_5475);
or U12353 (N_12353,N_6214,N_5685);
nand U12354 (N_12354,N_4615,N_1216);
and U12355 (N_12355,N_5913,N_4529);
and U12356 (N_12356,N_3259,N_1747);
nor U12357 (N_12357,N_5803,N_1862);
nand U12358 (N_12358,N_4407,N_1619);
xnor U12359 (N_12359,N_5740,N_1853);
xor U12360 (N_12360,N_3555,N_5999);
or U12361 (N_12361,N_597,N_3993);
nand U12362 (N_12362,N_5460,N_4705);
xor U12363 (N_12363,N_3513,N_1350);
nand U12364 (N_12364,N_3417,N_1039);
nand U12365 (N_12365,N_260,N_5644);
and U12366 (N_12366,N_6094,N_4871);
nor U12367 (N_12367,N_4000,N_3136);
nor U12368 (N_12368,N_4806,N_1390);
nand U12369 (N_12369,N_3574,N_6195);
nor U12370 (N_12370,N_4103,N_63);
and U12371 (N_12371,N_4365,N_339);
nand U12372 (N_12372,N_3205,N_4922);
and U12373 (N_12373,N_887,N_4949);
and U12374 (N_12374,N_3571,N_4640);
or U12375 (N_12375,N_119,N_2631);
nor U12376 (N_12376,N_4046,N_3882);
nor U12377 (N_12377,N_1603,N_1873);
nor U12378 (N_12378,N_895,N_5982);
or U12379 (N_12379,N_4084,N_1493);
nand U12380 (N_12380,N_980,N_4456);
nand U12381 (N_12381,N_2672,N_1882);
nor U12382 (N_12382,N_1242,N_1972);
and U12383 (N_12383,N_2679,N_541);
nor U12384 (N_12384,N_5425,N_61);
nor U12385 (N_12385,N_5793,N_3283);
or U12386 (N_12386,N_3923,N_4623);
nand U12387 (N_12387,N_39,N_5623);
or U12388 (N_12388,N_1014,N_5706);
and U12389 (N_12389,N_4288,N_3884);
and U12390 (N_12390,N_2652,N_181);
and U12391 (N_12391,N_4366,N_4670);
xnor U12392 (N_12392,N_6180,N_5030);
nor U12393 (N_12393,N_3565,N_3781);
nand U12394 (N_12394,N_5996,N_1292);
and U12395 (N_12395,N_1934,N_3125);
nor U12396 (N_12396,N_3314,N_5140);
xnor U12397 (N_12397,N_4072,N_2005);
xor U12398 (N_12398,N_3675,N_5749);
and U12399 (N_12399,N_3813,N_3229);
nor U12400 (N_12400,N_4125,N_1806);
xnor U12401 (N_12401,N_1374,N_1470);
and U12402 (N_12402,N_5374,N_3711);
and U12403 (N_12403,N_2532,N_3406);
xor U12404 (N_12404,N_1668,N_2565);
xnor U12405 (N_12405,N_1587,N_5087);
and U12406 (N_12406,N_680,N_2746);
nor U12407 (N_12407,N_3144,N_2298);
xor U12408 (N_12408,N_3661,N_3509);
or U12409 (N_12409,N_5119,N_2702);
and U12410 (N_12410,N_4130,N_113);
nand U12411 (N_12411,N_6008,N_1343);
or U12412 (N_12412,N_5916,N_5882);
nor U12413 (N_12413,N_4896,N_287);
and U12414 (N_12414,N_4990,N_1552);
or U12415 (N_12415,N_5711,N_1941);
nand U12416 (N_12416,N_5911,N_2210);
and U12417 (N_12417,N_6138,N_21);
nor U12418 (N_12418,N_1431,N_2335);
xor U12419 (N_12419,N_4150,N_2650);
nor U12420 (N_12420,N_4280,N_1327);
and U12421 (N_12421,N_2032,N_4422);
or U12422 (N_12422,N_809,N_2184);
and U12423 (N_12423,N_2606,N_1659);
nand U12424 (N_12424,N_2131,N_4194);
nand U12425 (N_12425,N_2313,N_3260);
and U12426 (N_12426,N_4187,N_5572);
nor U12427 (N_12427,N_4932,N_5598);
or U12428 (N_12428,N_779,N_932);
xnor U12429 (N_12429,N_5021,N_5699);
xnor U12430 (N_12430,N_400,N_1251);
nand U12431 (N_12431,N_630,N_6039);
or U12432 (N_12432,N_5936,N_3630);
or U12433 (N_12433,N_3210,N_1596);
nand U12434 (N_12434,N_4674,N_521);
nor U12435 (N_12435,N_1237,N_2404);
nand U12436 (N_12436,N_4499,N_5366);
or U12437 (N_12437,N_5969,N_1581);
or U12438 (N_12438,N_1148,N_899);
and U12439 (N_12439,N_1434,N_149);
and U12440 (N_12440,N_3761,N_2308);
or U12441 (N_12441,N_2424,N_4838);
or U12442 (N_12442,N_2200,N_3937);
xnor U12443 (N_12443,N_3038,N_5913);
or U12444 (N_12444,N_306,N_2511);
or U12445 (N_12445,N_2789,N_3737);
and U12446 (N_12446,N_6113,N_2696);
nor U12447 (N_12447,N_4850,N_669);
xor U12448 (N_12448,N_5314,N_168);
or U12449 (N_12449,N_6085,N_5619);
nor U12450 (N_12450,N_5160,N_362);
nor U12451 (N_12451,N_2789,N_4964);
nor U12452 (N_12452,N_3430,N_1942);
or U12453 (N_12453,N_1895,N_4854);
and U12454 (N_12454,N_4131,N_3459);
xnor U12455 (N_12455,N_2021,N_5928);
nor U12456 (N_12456,N_76,N_71);
and U12457 (N_12457,N_4422,N_6107);
nor U12458 (N_12458,N_498,N_945);
nor U12459 (N_12459,N_1678,N_3227);
or U12460 (N_12460,N_5012,N_3700);
or U12461 (N_12461,N_35,N_3317);
or U12462 (N_12462,N_5645,N_5582);
nand U12463 (N_12463,N_2978,N_2840);
or U12464 (N_12464,N_4850,N_6027);
xnor U12465 (N_12465,N_699,N_397);
nand U12466 (N_12466,N_4282,N_4914);
nor U12467 (N_12467,N_3771,N_1710);
and U12468 (N_12468,N_3986,N_2884);
and U12469 (N_12469,N_798,N_5562);
or U12470 (N_12470,N_2527,N_5074);
nand U12471 (N_12471,N_2745,N_2521);
xor U12472 (N_12472,N_4982,N_4594);
nor U12473 (N_12473,N_1251,N_3754);
nor U12474 (N_12474,N_5780,N_461);
or U12475 (N_12475,N_5441,N_2394);
nand U12476 (N_12476,N_4087,N_4290);
nand U12477 (N_12477,N_4400,N_3471);
nor U12478 (N_12478,N_5003,N_4985);
nand U12479 (N_12479,N_1747,N_859);
xor U12480 (N_12480,N_1111,N_3752);
nand U12481 (N_12481,N_5556,N_4032);
xor U12482 (N_12482,N_2900,N_212);
nand U12483 (N_12483,N_5530,N_3665);
or U12484 (N_12484,N_3696,N_6209);
and U12485 (N_12485,N_5027,N_627);
nand U12486 (N_12486,N_3936,N_126);
xor U12487 (N_12487,N_2874,N_6239);
and U12488 (N_12488,N_5178,N_961);
nand U12489 (N_12489,N_1348,N_4668);
nand U12490 (N_12490,N_5584,N_2431);
nand U12491 (N_12491,N_2521,N_425);
and U12492 (N_12492,N_2244,N_1030);
and U12493 (N_12493,N_5636,N_3939);
nand U12494 (N_12494,N_2355,N_2842);
nand U12495 (N_12495,N_684,N_4939);
nor U12496 (N_12496,N_1937,N_5249);
or U12497 (N_12497,N_2806,N_5342);
and U12498 (N_12498,N_3597,N_5779);
xor U12499 (N_12499,N_925,N_1555);
or U12500 (N_12500,N_11126,N_10508);
nand U12501 (N_12501,N_6647,N_8899);
and U12502 (N_12502,N_11141,N_9732);
xor U12503 (N_12503,N_9728,N_10283);
and U12504 (N_12504,N_12235,N_9001);
nand U12505 (N_12505,N_6493,N_9205);
xor U12506 (N_12506,N_11186,N_10081);
nand U12507 (N_12507,N_12195,N_12449);
nand U12508 (N_12508,N_8895,N_8516);
nand U12509 (N_12509,N_11779,N_9597);
nand U12510 (N_12510,N_7062,N_9570);
xnor U12511 (N_12511,N_8556,N_11272);
and U12512 (N_12512,N_10029,N_6847);
xor U12513 (N_12513,N_7970,N_7006);
or U12514 (N_12514,N_9095,N_8723);
and U12515 (N_12515,N_9510,N_10743);
nor U12516 (N_12516,N_12207,N_11408);
or U12517 (N_12517,N_6892,N_11856);
xnor U12518 (N_12518,N_6571,N_10308);
nor U12519 (N_12519,N_9514,N_7540);
and U12520 (N_12520,N_7881,N_11072);
xor U12521 (N_12521,N_11235,N_7903);
nand U12522 (N_12522,N_6548,N_10120);
or U12523 (N_12523,N_10864,N_9152);
nand U12524 (N_12524,N_6653,N_12476);
and U12525 (N_12525,N_8449,N_10357);
xnor U12526 (N_12526,N_9127,N_9981);
xor U12527 (N_12527,N_8925,N_8035);
or U12528 (N_12528,N_7964,N_11871);
and U12529 (N_12529,N_7063,N_10032);
nor U12530 (N_12530,N_8621,N_8459);
or U12531 (N_12531,N_9388,N_11417);
or U12532 (N_12532,N_6894,N_9947);
nor U12533 (N_12533,N_7913,N_7546);
and U12534 (N_12534,N_7982,N_7478);
and U12535 (N_12535,N_6725,N_9761);
nand U12536 (N_12536,N_12424,N_9929);
or U12537 (N_12537,N_11810,N_11735);
nand U12538 (N_12538,N_9557,N_6928);
xnor U12539 (N_12539,N_7604,N_8849);
and U12540 (N_12540,N_11113,N_8606);
nor U12541 (N_12541,N_7525,N_11159);
and U12542 (N_12542,N_7998,N_9181);
nor U12543 (N_12543,N_10822,N_10232);
and U12544 (N_12544,N_8773,N_6632);
nor U12545 (N_12545,N_11544,N_10644);
nor U12546 (N_12546,N_9771,N_9989);
or U12547 (N_12547,N_10615,N_11323);
nand U12548 (N_12548,N_7953,N_9183);
nand U12549 (N_12549,N_11898,N_7190);
xnor U12550 (N_12550,N_11382,N_7782);
or U12551 (N_12551,N_12233,N_11004);
nand U12552 (N_12552,N_11513,N_10141);
and U12553 (N_12553,N_12458,N_11669);
nand U12554 (N_12554,N_7298,N_6325);
or U12555 (N_12555,N_7343,N_11054);
xnor U12556 (N_12556,N_10038,N_10041);
and U12557 (N_12557,N_6413,N_7716);
xor U12558 (N_12558,N_9263,N_12145);
and U12559 (N_12559,N_8192,N_9889);
nor U12560 (N_12560,N_7284,N_12150);
nand U12561 (N_12561,N_11612,N_10335);
and U12562 (N_12562,N_9968,N_11028);
or U12563 (N_12563,N_6883,N_10079);
nand U12564 (N_12564,N_7196,N_9232);
xnor U12565 (N_12565,N_7025,N_10151);
and U12566 (N_12566,N_9290,N_7107);
and U12567 (N_12567,N_10467,N_6408);
nor U12568 (N_12568,N_7094,N_10218);
xor U12569 (N_12569,N_10778,N_11104);
or U12570 (N_12570,N_11070,N_10868);
xnor U12571 (N_12571,N_6474,N_6665);
nand U12572 (N_12572,N_7297,N_9223);
nand U12573 (N_12573,N_7395,N_6314);
nor U12574 (N_12574,N_8215,N_10674);
nand U12575 (N_12575,N_7447,N_9988);
nor U12576 (N_12576,N_9688,N_8846);
nand U12577 (N_12577,N_11430,N_11448);
xnor U12578 (N_12578,N_6902,N_12058);
xor U12579 (N_12579,N_9375,N_7558);
xnor U12580 (N_12580,N_10682,N_9116);
xor U12581 (N_12581,N_12399,N_7210);
nor U12582 (N_12582,N_7225,N_9666);
xor U12583 (N_12583,N_6843,N_10680);
xnor U12584 (N_12584,N_11158,N_9273);
nor U12585 (N_12585,N_8345,N_9569);
xnor U12586 (N_12586,N_11532,N_9540);
and U12587 (N_12587,N_9500,N_12271);
nor U12588 (N_12588,N_9280,N_11608);
xnor U12589 (N_12589,N_8826,N_11862);
xnor U12590 (N_12590,N_7130,N_6643);
and U12591 (N_12591,N_11212,N_7232);
and U12592 (N_12592,N_9114,N_8324);
and U12593 (N_12593,N_9503,N_9701);
and U12594 (N_12594,N_10803,N_7852);
or U12595 (N_12595,N_6719,N_10236);
and U12596 (N_12596,N_7317,N_9920);
or U12597 (N_12597,N_7383,N_10178);
and U12598 (N_12598,N_7844,N_7874);
xor U12599 (N_12599,N_10890,N_6924);
xnor U12600 (N_12600,N_9274,N_10581);
xor U12601 (N_12601,N_11986,N_6416);
nand U12602 (N_12602,N_8744,N_9966);
and U12603 (N_12603,N_7932,N_6874);
and U12604 (N_12604,N_10645,N_11407);
and U12605 (N_12605,N_9584,N_6779);
or U12606 (N_12606,N_10115,N_6385);
xor U12607 (N_12607,N_8398,N_7240);
xnor U12608 (N_12608,N_7472,N_6771);
nand U12609 (N_12609,N_10661,N_6401);
and U12610 (N_12610,N_9170,N_10769);
or U12611 (N_12611,N_11223,N_8778);
or U12612 (N_12612,N_8421,N_10612);
nor U12613 (N_12613,N_12358,N_7281);
xnor U12614 (N_12614,N_11746,N_10948);
xor U12615 (N_12615,N_11447,N_9367);
xor U12616 (N_12616,N_7060,N_6830);
or U12617 (N_12617,N_6618,N_7363);
and U12618 (N_12618,N_8876,N_9011);
xnor U12619 (N_12619,N_6681,N_9803);
xnor U12620 (N_12620,N_12492,N_10498);
or U12621 (N_12621,N_10731,N_10820);
nand U12622 (N_12622,N_8332,N_9348);
nand U12623 (N_12623,N_9305,N_7924);
nand U12624 (N_12624,N_12227,N_11869);
or U12625 (N_12625,N_6983,N_7526);
nand U12626 (N_12626,N_9511,N_7246);
or U12627 (N_12627,N_11795,N_12061);
and U12628 (N_12628,N_9296,N_12133);
or U12629 (N_12629,N_8133,N_6578);
nand U12630 (N_12630,N_9244,N_10251);
and U12631 (N_12631,N_6755,N_10815);
nor U12632 (N_12632,N_6270,N_11075);
xnor U12633 (N_12633,N_9617,N_11578);
xnor U12634 (N_12634,N_9864,N_7047);
nor U12635 (N_12635,N_9397,N_8143);
nand U12636 (N_12636,N_9137,N_11674);
or U12637 (N_12637,N_12077,N_7419);
and U12638 (N_12638,N_11432,N_8278);
xnor U12639 (N_12639,N_11250,N_9174);
and U12640 (N_12640,N_8205,N_6484);
and U12641 (N_12641,N_8637,N_9786);
and U12642 (N_12642,N_8063,N_11256);
or U12643 (N_12643,N_10920,N_9749);
nor U12644 (N_12644,N_7693,N_7099);
xor U12645 (N_12645,N_11482,N_11575);
or U12646 (N_12646,N_11248,N_12041);
nand U12647 (N_12647,N_8655,N_11917);
xor U12648 (N_12648,N_9319,N_10454);
xor U12649 (N_12649,N_12286,N_12373);
nor U12650 (N_12650,N_7128,N_8206);
or U12651 (N_12651,N_11894,N_6567);
and U12652 (N_12652,N_6595,N_7642);
xor U12653 (N_12653,N_10909,N_9381);
nand U12654 (N_12654,N_12276,N_11255);
and U12655 (N_12655,N_10771,N_10233);
xor U12656 (N_12656,N_8460,N_7274);
nor U12657 (N_12657,N_6423,N_10895);
xnor U12658 (N_12658,N_8738,N_9795);
xnor U12659 (N_12659,N_12438,N_7988);
or U12660 (N_12660,N_8557,N_7502);
nor U12661 (N_12661,N_9598,N_9055);
nand U12662 (N_12662,N_8707,N_6351);
xor U12663 (N_12663,N_7519,N_9379);
xnor U12664 (N_12664,N_12322,N_6251);
or U12665 (N_12665,N_10159,N_8817);
nand U12666 (N_12666,N_11355,N_10226);
or U12667 (N_12667,N_7905,N_10985);
and U12668 (N_12668,N_11463,N_10336);
nand U12669 (N_12669,N_10238,N_7591);
or U12670 (N_12670,N_10906,N_7077);
and U12671 (N_12671,N_9233,N_7795);
and U12672 (N_12672,N_8253,N_8720);
and U12673 (N_12673,N_10026,N_6706);
or U12674 (N_12674,N_6387,N_10254);
xor U12675 (N_12675,N_9671,N_8104);
nand U12676 (N_12676,N_11800,N_11787);
or U12677 (N_12677,N_9143,N_11650);
and U12678 (N_12678,N_8222,N_8670);
nand U12679 (N_12679,N_8545,N_9655);
and U12680 (N_12680,N_7338,N_9742);
nand U12681 (N_12681,N_7763,N_9428);
nand U12682 (N_12682,N_6391,N_10738);
xnor U12683 (N_12683,N_6508,N_7718);
nand U12684 (N_12684,N_12076,N_9533);
and U12685 (N_12685,N_8646,N_6613);
or U12686 (N_12686,N_9357,N_10714);
and U12687 (N_12687,N_7115,N_10175);
nand U12688 (N_12688,N_10973,N_8033);
nand U12689 (N_12689,N_11486,N_11279);
and U12690 (N_12690,N_9494,N_8737);
and U12691 (N_12691,N_8787,N_10307);
or U12692 (N_12692,N_10568,N_9365);
xor U12693 (N_12693,N_11540,N_9396);
and U12694 (N_12694,N_8057,N_7846);
xnor U12695 (N_12695,N_6935,N_10294);
or U12696 (N_12696,N_8942,N_7837);
nand U12697 (N_12697,N_7574,N_9960);
nor U12698 (N_12698,N_6263,N_11362);
nand U12699 (N_12699,N_11309,N_8704);
and U12700 (N_12700,N_6676,N_8464);
nand U12701 (N_12701,N_8923,N_9343);
nand U12702 (N_12702,N_9559,N_8082);
xor U12703 (N_12703,N_6357,N_6992);
xor U12704 (N_12704,N_12236,N_9142);
nand U12705 (N_12705,N_11844,N_6936);
and U12706 (N_12706,N_7646,N_8184);
and U12707 (N_12707,N_12383,N_10669);
xor U12708 (N_12708,N_9812,N_12436);
nor U12709 (N_12709,N_10514,N_7163);
or U12710 (N_12710,N_10284,N_10885);
or U12711 (N_12711,N_7984,N_6574);
and U12712 (N_12712,N_8496,N_8906);
or U12713 (N_12713,N_9391,N_9470);
nor U12714 (N_12714,N_7167,N_10882);
and U12715 (N_12715,N_11115,N_10225);
and U12716 (N_12716,N_12310,N_8197);
xor U12717 (N_12717,N_11500,N_8370);
nand U12718 (N_12718,N_7530,N_9899);
nor U12719 (N_12719,N_9302,N_9744);
xor U12720 (N_12720,N_7310,N_11767);
and U12721 (N_12721,N_8209,N_12388);
nor U12722 (N_12722,N_7853,N_7332);
and U12723 (N_12723,N_11994,N_6486);
nor U12724 (N_12724,N_9667,N_9188);
or U12725 (N_12725,N_7364,N_11055);
nor U12726 (N_12726,N_8589,N_6481);
nor U12727 (N_12727,N_10306,N_7076);
or U12728 (N_12728,N_7545,N_10595);
and U12729 (N_12729,N_10886,N_6887);
xor U12730 (N_12730,N_7926,N_10659);
nand U12731 (N_12731,N_7251,N_6916);
or U12732 (N_12732,N_11818,N_9478);
xor U12733 (N_12733,N_11556,N_9316);
nor U12734 (N_12734,N_12242,N_6603);
or U12735 (N_12735,N_10910,N_12452);
or U12736 (N_12736,N_10200,N_7208);
and U12737 (N_12737,N_9279,N_11858);
nand U12738 (N_12738,N_10795,N_9099);
and U12739 (N_12739,N_8991,N_7814);
xor U12740 (N_12740,N_9507,N_8513);
xor U12741 (N_12741,N_8062,N_7688);
xnor U12742 (N_12742,N_9271,N_10417);
and U12743 (N_12743,N_8588,N_10511);
and U12744 (N_12744,N_10340,N_10314);
or U12745 (N_12745,N_12109,N_10300);
or U12746 (N_12746,N_7972,N_6397);
or U12747 (N_12747,N_12071,N_11657);
xor U12748 (N_12748,N_11456,N_9860);
and U12749 (N_12749,N_7108,N_8664);
nand U12750 (N_12750,N_6298,N_11013);
nor U12751 (N_12751,N_11812,N_11849);
xnor U12752 (N_12752,N_10978,N_11438);
and U12753 (N_12753,N_7470,N_9096);
or U12754 (N_12754,N_10935,N_7566);
nand U12755 (N_12755,N_12244,N_7333);
nand U12756 (N_12756,N_9974,N_10875);
nand U12757 (N_12757,N_10927,N_11748);
xor U12758 (N_12758,N_12411,N_10524);
or U12759 (N_12759,N_6995,N_10360);
or U12760 (N_12760,N_9735,N_11506);
nor U12761 (N_12761,N_7304,N_11586);
nor U12762 (N_12762,N_8495,N_10222);
and U12763 (N_12763,N_9798,N_6480);
nand U12764 (N_12764,N_9878,N_7503);
nand U12765 (N_12765,N_8487,N_10916);
xor U12766 (N_12766,N_12090,N_7560);
xnor U12767 (N_12767,N_9684,N_10492);
and U12768 (N_12768,N_8970,N_10835);
xnor U12769 (N_12769,N_9841,N_6692);
nor U12770 (N_12770,N_10521,N_6309);
xor U12771 (N_12771,N_10441,N_9627);
nand U12772 (N_12772,N_11040,N_8125);
xor U12773 (N_12773,N_11496,N_11139);
xnor U12774 (N_12774,N_9487,N_9586);
nor U12775 (N_12775,N_8889,N_11807);
xor U12776 (N_12776,N_9562,N_11777);
or U12777 (N_12777,N_8090,N_7695);
nor U12778 (N_12778,N_7725,N_11985);
nor U12779 (N_12779,N_11332,N_10870);
xnor U12780 (N_12780,N_6592,N_10427);
nor U12781 (N_12781,N_11011,N_12444);
nand U12782 (N_12782,N_7028,N_9501);
nand U12783 (N_12783,N_8410,N_8521);
nor U12784 (N_12784,N_12191,N_8081);
xnor U12785 (N_12785,N_11225,N_6498);
xnor U12786 (N_12786,N_7501,N_11231);
nand U12787 (N_12787,N_9564,N_10326);
or U12788 (N_12788,N_8167,N_9431);
xor U12789 (N_12789,N_8186,N_10549);
nor U12790 (N_12790,N_7670,N_10630);
nor U12791 (N_12791,N_9252,N_7738);
and U12792 (N_12792,N_10000,N_8668);
nor U12793 (N_12793,N_6952,N_6475);
and U12794 (N_12794,N_9068,N_8187);
nand U12795 (N_12795,N_12105,N_10555);
nor U12796 (N_12796,N_8008,N_10031);
and U12797 (N_12797,N_8048,N_7969);
nor U12798 (N_12798,N_12184,N_7262);
or U12799 (N_12799,N_9956,N_11234);
or U12800 (N_12800,N_8853,N_10631);
nand U12801 (N_12801,N_7605,N_11038);
nor U12802 (N_12802,N_12282,N_12047);
nor U12803 (N_12803,N_11947,N_8497);
nand U12804 (N_12804,N_11281,N_8973);
and U12805 (N_12805,N_10312,N_7014);
xnor U12806 (N_12806,N_9896,N_11307);
nand U12807 (N_12807,N_8483,N_9577);
xnor U12808 (N_12808,N_6772,N_6739);
nor U12809 (N_12809,N_10107,N_8872);
nand U12810 (N_12810,N_8536,N_8602);
nor U12811 (N_12811,N_7171,N_8444);
xnor U12812 (N_12812,N_8198,N_11966);
and U12813 (N_12813,N_7942,N_8885);
xnor U12814 (N_12814,N_7404,N_11222);
and U12815 (N_12815,N_10628,N_10375);
nand U12816 (N_12816,N_10167,N_7160);
or U12817 (N_12817,N_12313,N_8266);
and U12818 (N_12818,N_7214,N_12367);
xnor U12819 (N_12819,N_9418,N_7151);
or U12820 (N_12820,N_6842,N_11048);
nor U12821 (N_12821,N_8023,N_6758);
or U12822 (N_12822,N_10535,N_9964);
nand U12823 (N_12823,N_11784,N_12381);
and U12824 (N_12824,N_7557,N_8013);
xor U12825 (N_12825,N_11446,N_6956);
and U12826 (N_12826,N_7911,N_9058);
nor U12827 (N_12827,N_8381,N_8979);
and U12828 (N_12828,N_10476,N_9179);
and U12829 (N_12829,N_10426,N_12481);
xnor U12830 (N_12830,N_8654,N_7097);
nor U12831 (N_12831,N_6683,N_11458);
and U12832 (N_12832,N_6748,N_8193);
nand U12833 (N_12833,N_9460,N_9619);
and U12834 (N_12834,N_10692,N_6732);
nor U12835 (N_12835,N_6811,N_6791);
xnor U12836 (N_12836,N_8331,N_10063);
or U12837 (N_12837,N_11983,N_9625);
xor U12838 (N_12838,N_7039,N_10364);
nand U12839 (N_12839,N_8477,N_6269);
nand U12840 (N_12840,N_8191,N_8501);
or U12841 (N_12841,N_10675,N_11488);
xnor U12842 (N_12842,N_12219,N_8056);
or U12843 (N_12843,N_10704,N_7631);
nor U12844 (N_12844,N_9685,N_11238);
and U12845 (N_12845,N_9282,N_7660);
xor U12846 (N_12846,N_12321,N_8416);
xor U12847 (N_12847,N_11991,N_10433);
and U12848 (N_12848,N_10030,N_11153);
xnor U12849 (N_12849,N_9306,N_11593);
and U12850 (N_12850,N_7464,N_11185);
nor U12851 (N_12851,N_8042,N_10726);
or U12852 (N_12852,N_10366,N_6318);
or U12853 (N_12853,N_11830,N_7860);
and U12854 (N_12854,N_9032,N_6875);
xor U12855 (N_12855,N_11814,N_8811);
xnor U12856 (N_12856,N_12098,N_6261);
nand U12857 (N_12857,N_11128,N_11919);
or U12858 (N_12858,N_12027,N_10527);
or U12859 (N_12859,N_10171,N_10515);
and U12860 (N_12860,N_11330,N_6967);
nor U12861 (N_12861,N_10878,N_8815);
and U12862 (N_12862,N_9024,N_8924);
and U12863 (N_12863,N_7523,N_7320);
nor U12864 (N_12864,N_11311,N_11009);
xnor U12865 (N_12865,N_7941,N_10755);
xor U12866 (N_12866,N_9030,N_7597);
nor U12867 (N_12867,N_8547,N_12176);
nor U12868 (N_12868,N_11706,N_12127);
or U12869 (N_12869,N_8369,N_6450);
nand U12870 (N_12870,N_8624,N_8856);
or U12871 (N_12871,N_10787,N_6795);
or U12872 (N_12872,N_12342,N_8433);
nand U12873 (N_12873,N_9107,N_7052);
xnor U12874 (N_12874,N_11228,N_9019);
nor U12875 (N_12875,N_10852,N_8659);
and U12876 (N_12876,N_6915,N_12249);
nand U12877 (N_12877,N_7778,N_7770);
nand U12878 (N_12878,N_8060,N_7512);
or U12879 (N_12879,N_10642,N_8880);
and U12880 (N_12880,N_8164,N_7682);
xor U12881 (N_12881,N_10610,N_10428);
or U12882 (N_12882,N_11123,N_9034);
nand U12883 (N_12883,N_8950,N_7544);
nand U12884 (N_12884,N_7368,N_7451);
nor U12885 (N_12885,N_8007,N_6579);
or U12886 (N_12886,N_7336,N_7956);
or U12887 (N_12887,N_9120,N_10707);
nor U12888 (N_12888,N_10474,N_10698);
nor U12889 (N_12889,N_7684,N_8219);
or U12890 (N_12890,N_8210,N_9243);
nand U12891 (N_12891,N_12314,N_12043);
and U12892 (N_12892,N_10809,N_10784);
nor U12893 (N_12893,N_8393,N_7069);
xnor U12894 (N_12894,N_10880,N_11956);
nand U12895 (N_12895,N_9637,N_6421);
nor U12896 (N_12896,N_11006,N_8458);
xnor U12897 (N_12897,N_9249,N_11628);
and U12898 (N_12898,N_10172,N_10046);
or U12899 (N_12899,N_11096,N_10083);
nand U12900 (N_12900,N_9547,N_7637);
nand U12901 (N_12901,N_9476,N_6328);
or U12902 (N_12902,N_9147,N_7263);
and U12903 (N_12903,N_10278,N_6855);
or U12904 (N_12904,N_8208,N_9502);
or U12905 (N_12905,N_11389,N_10737);
nor U12906 (N_12906,N_9884,N_10087);
nor U12907 (N_12907,N_11051,N_7068);
nor U12908 (N_12908,N_10520,N_11077);
nor U12909 (N_12909,N_8653,N_8328);
nand U12910 (N_12910,N_6953,N_12439);
xor U12911 (N_12911,N_8956,N_11258);
nand U12912 (N_12912,N_10440,N_10466);
nor U12913 (N_12913,N_8879,N_9387);
xor U12914 (N_12914,N_6642,N_7510);
and U12915 (N_12915,N_11662,N_6965);
xnor U12916 (N_12916,N_12395,N_11973);
nor U12917 (N_12917,N_12220,N_10398);
nand U12918 (N_12918,N_11783,N_9443);
nand U12919 (N_12919,N_7719,N_8128);
xnor U12920 (N_12920,N_11270,N_7830);
nor U12921 (N_12921,N_11673,N_6334);
nor U12922 (N_12922,N_6738,N_12084);
nand U12923 (N_12923,N_7840,N_10449);
or U12924 (N_12924,N_8179,N_8274);
or U12925 (N_12925,N_8947,N_9076);
nor U12926 (N_12926,N_6788,N_7629);
nand U12927 (N_12927,N_6551,N_8898);
xnor U12928 (N_12928,N_12026,N_9139);
nor U12929 (N_12929,N_10565,N_9285);
nor U12930 (N_12930,N_11184,N_11618);
nor U12931 (N_12931,N_11741,N_7593);
or U12932 (N_12932,N_10198,N_11291);
nor U12933 (N_12933,N_8200,N_11968);
nor U12934 (N_12934,N_10318,N_8714);
or U12935 (N_12935,N_8718,N_8298);
or U12936 (N_12936,N_7397,N_7382);
nor U12937 (N_12937,N_12122,N_6296);
or U12938 (N_12938,N_8524,N_7949);
nor U12939 (N_12939,N_7669,N_7974);
xnor U12940 (N_12940,N_10173,N_8795);
or U12941 (N_12941,N_10712,N_8339);
or U12942 (N_12942,N_8816,N_9260);
nor U12943 (N_12943,N_12432,N_9835);
xnor U12944 (N_12944,N_10597,N_8387);
or U12945 (N_12945,N_7437,N_9363);
nand U12946 (N_12946,N_8257,N_6422);
and U12947 (N_12947,N_11083,N_10324);
nand U12948 (N_12948,N_11473,N_6250);
nand U12949 (N_12949,N_8270,N_9031);
nor U12950 (N_12950,N_11630,N_6724);
nor U12951 (N_12951,N_9948,N_6289);
xor U12952 (N_12952,N_12232,N_6557);
nand U12953 (N_12953,N_11501,N_11824);
or U12954 (N_12954,N_6808,N_7549);
xnor U12955 (N_12955,N_10007,N_11899);
xor U12956 (N_12956,N_10673,N_9508);
nor U12957 (N_12957,N_8201,N_8835);
xnor U12958 (N_12958,N_8523,N_10656);
and U12959 (N_12959,N_8310,N_11672);
xnor U12960 (N_12960,N_10619,N_11404);
and U12961 (N_12961,N_10637,N_6654);
nor U12962 (N_12962,N_11731,N_7730);
or U12963 (N_12963,N_11663,N_7462);
nor U12964 (N_12964,N_7999,N_11419);
nor U12965 (N_12965,N_6737,N_10231);
nand U12966 (N_12966,N_12456,N_7564);
xnor U12967 (N_12967,N_7004,N_8202);
and U12968 (N_12968,N_10983,N_10451);
nor U12969 (N_12969,N_10846,N_6867);
nor U12970 (N_12970,N_10108,N_9103);
nand U12971 (N_12971,N_11635,N_11936);
and U12972 (N_12972,N_6945,N_7042);
and U12973 (N_12973,N_7319,N_7453);
nand U12974 (N_12974,N_11959,N_8805);
xnor U12975 (N_12975,N_12253,N_11464);
nor U12976 (N_12976,N_6369,N_6908);
nor U12977 (N_12977,N_7485,N_6346);
nor U12978 (N_12978,N_7239,N_9741);
or U12979 (N_12979,N_10177,N_9861);
and U12980 (N_12980,N_10235,N_9416);
and U12981 (N_12981,N_11656,N_8583);
xor U12982 (N_12982,N_8877,N_8156);
nand U12983 (N_12983,N_7012,N_6471);
nand U12984 (N_12984,N_11439,N_6671);
nand U12985 (N_12985,N_11740,N_8633);
nor U12986 (N_12986,N_11230,N_10827);
or U12987 (N_12987,N_10197,N_9925);
nand U12988 (N_12988,N_11308,N_9506);
nand U12989 (N_12989,N_8262,N_8550);
or U12990 (N_12990,N_9498,N_10034);
nor U12991 (N_12991,N_11970,N_8785);
xor U12992 (N_12992,N_7474,N_10599);
xnor U12993 (N_12993,N_12451,N_6761);
nor U12994 (N_12994,N_9373,N_9719);
nor U12995 (N_12995,N_12164,N_6439);
and U12996 (N_12996,N_7520,N_7231);
nor U12997 (N_12997,N_11387,N_12487);
nor U12998 (N_12998,N_7329,N_11088);
nor U12999 (N_12999,N_12437,N_6650);
and U13000 (N_13000,N_7638,N_6539);
or U13001 (N_13001,N_7165,N_11867);
xnor U13002 (N_13002,N_8951,N_10963);
nand U13003 (N_13003,N_6386,N_8406);
nand U13004 (N_13004,N_8995,N_7575);
nor U13005 (N_13005,N_8551,N_12094);
and U13006 (N_13006,N_6379,N_9286);
xor U13007 (N_13007,N_10329,N_7863);
nand U13008 (N_13008,N_7402,N_10588);
and U13009 (N_13009,N_12025,N_11529);
or U13010 (N_13010,N_10378,N_11512);
nand U13011 (N_13011,N_10700,N_7767);
and U13012 (N_13012,N_8093,N_8251);
nor U13013 (N_13013,N_12151,N_6291);
nor U13014 (N_13014,N_10240,N_6392);
xor U13015 (N_13015,N_8226,N_11493);
nor U13016 (N_13016,N_11197,N_12416);
xor U13017 (N_13017,N_9109,N_9295);
nand U13018 (N_13018,N_12407,N_6777);
or U13019 (N_13019,N_9405,N_7352);
and U13020 (N_13020,N_10718,N_8265);
and U13021 (N_13021,N_12425,N_7686);
nand U13022 (N_13022,N_9571,N_12199);
xnor U13023 (N_13023,N_7141,N_9199);
nor U13024 (N_13024,N_6774,N_8608);
and U13025 (N_13025,N_10723,N_11987);
or U13026 (N_13026,N_6868,N_6490);
and U13027 (N_13027,N_8442,N_10447);
xnor U13028 (N_13028,N_9880,N_10831);
and U13029 (N_13029,N_8452,N_8977);
nor U13030 (N_13030,N_11237,N_7040);
or U13031 (N_13031,N_12277,N_8552);
or U13032 (N_13032,N_9230,N_8404);
and U13033 (N_13033,N_10189,N_7921);
nand U13034 (N_13034,N_12472,N_10092);
xnor U13035 (N_13035,N_12108,N_8269);
nand U13036 (N_13036,N_6405,N_8250);
xnor U13037 (N_13037,N_8910,N_7418);
nand U13038 (N_13038,N_7901,N_7704);
nand U13039 (N_13039,N_11027,N_7715);
and U13040 (N_13040,N_11629,N_8825);
xor U13041 (N_13041,N_9862,N_9628);
xor U13042 (N_13042,N_7614,N_11350);
nor U13043 (N_13043,N_7993,N_10352);
nand U13044 (N_13044,N_7583,N_11162);
nor U13045 (N_13045,N_6871,N_10721);
nand U13046 (N_13046,N_6521,N_11356);
or U13047 (N_13047,N_11178,N_10613);
nand U13048 (N_13048,N_11964,N_6520);
xnor U13049 (N_13049,N_9594,N_12468);
nor U13050 (N_13050,N_9550,N_11091);
and U13051 (N_13051,N_12273,N_7005);
xnor U13052 (N_13052,N_9875,N_12017);
and U13053 (N_13053,N_10944,N_9954);
nand U13054 (N_13054,N_11560,N_6881);
or U13055 (N_13055,N_12318,N_10557);
xor U13056 (N_13056,N_10987,N_12185);
nor U13057 (N_13057,N_11286,N_8363);
nor U13058 (N_13058,N_12360,N_12116);
nor U13059 (N_13059,N_6382,N_7082);
and U13060 (N_13060,N_8508,N_8686);
or U13061 (N_13061,N_11978,N_9384);
nand U13062 (N_13062,N_8292,N_8688);
nand U13063 (N_13063,N_8358,N_9119);
and U13064 (N_13064,N_6646,N_10842);
xor U13065 (N_13065,N_9490,N_7493);
or U13066 (N_13066,N_12114,N_9612);
and U13067 (N_13067,N_12131,N_7341);
or U13068 (N_13068,N_10327,N_11246);
xor U13069 (N_13069,N_6470,N_11900);
nand U13070 (N_13070,N_9372,N_8935);
xnor U13071 (N_13071,N_7002,N_7586);
and U13072 (N_13072,N_12008,N_7156);
nand U13073 (N_13073,N_7027,N_11604);
and U13074 (N_13074,N_10372,N_9457);
nor U13075 (N_13075,N_8820,N_7460);
xor U13076 (N_13076,N_6449,N_8320);
xor U13077 (N_13077,N_12317,N_9410);
or U13078 (N_13078,N_11012,N_7973);
nand U13079 (N_13079,N_7408,N_7134);
nor U13080 (N_13080,N_11436,N_7906);
and U13081 (N_13081,N_10843,N_7954);
xnor U13082 (N_13082,N_9014,N_7439);
xor U13083 (N_13083,N_11887,N_10996);
xor U13084 (N_13084,N_10190,N_8985);
nor U13085 (N_13085,N_12368,N_9007);
nor U13086 (N_13086,N_9872,N_9876);
xnor U13087 (N_13087,N_8751,N_7979);
nor U13088 (N_13088,N_7757,N_9323);
xor U13089 (N_13089,N_6549,N_6476);
or U13090 (N_13090,N_7198,N_12409);
or U13091 (N_13091,N_9089,N_8595);
xnor U13092 (N_13092,N_7559,N_7031);
xnor U13093 (N_13093,N_9300,N_7087);
or U13094 (N_13094,N_6550,N_10664);
and U13095 (N_13095,N_7119,N_8518);
nand U13096 (N_13096,N_8634,N_9452);
and U13097 (N_13097,N_9950,N_8401);
or U13098 (N_13098,N_8706,N_7098);
nand U13099 (N_13099,N_10811,N_8175);
xor U13100 (N_13100,N_6922,N_8758);
nand U13101 (N_13101,N_10431,N_11846);
xor U13102 (N_13102,N_10657,N_9588);
or U13103 (N_13103,N_8453,N_7791);
and U13104 (N_13104,N_6509,N_7733);
and U13105 (N_13105,N_8323,N_7432);
nand U13106 (N_13106,N_7743,N_6785);
xnor U13107 (N_13107,N_8700,N_8380);
and U13108 (N_13108,N_7976,N_8859);
xnor U13109 (N_13109,N_7977,N_11349);
nand U13110 (N_13110,N_9662,N_8343);
nand U13111 (N_13111,N_8967,N_9814);
or U13112 (N_13112,N_7235,N_7102);
or U13113 (N_13113,N_7385,N_10291);
or U13114 (N_13114,N_10382,N_6865);
nor U13115 (N_13115,N_11980,N_10146);
nand U13116 (N_13116,N_6715,N_10814);
or U13117 (N_13117,N_7584,N_10564);
nor U13118 (N_13118,N_10725,N_10767);
nor U13119 (N_13119,N_7112,N_12413);
and U13120 (N_13120,N_12331,N_11333);
or U13121 (N_13121,N_9969,N_11817);
and U13122 (N_13122,N_6997,N_6821);
nor U13123 (N_13123,N_6819,N_6586);
nor U13124 (N_13124,N_7075,N_10857);
xnor U13125 (N_13125,N_6781,N_11049);
nor U13126 (N_13126,N_6456,N_10044);
nand U13127 (N_13127,N_11546,N_7659);
or U13128 (N_13128,N_8150,N_10179);
xnor U13129 (N_13129,N_12243,N_12394);
or U13130 (N_13130,N_11336,N_9400);
or U13131 (N_13131,N_7960,N_7289);
nor U13132 (N_13132,N_6398,N_10202);
and U13133 (N_13133,N_8632,N_7420);
xnor U13134 (N_13134,N_8256,N_8986);
nor U13135 (N_13135,N_6287,N_7789);
nor U13136 (N_13136,N_10261,N_6904);
or U13137 (N_13137,N_7030,N_9005);
and U13138 (N_13138,N_10269,N_9760);
or U13139 (N_13139,N_8867,N_9832);
nand U13140 (N_13140,N_7562,N_8617);
nand U13141 (N_13141,N_10429,N_10273);
xor U13142 (N_13142,N_7350,N_7433);
nand U13143 (N_13143,N_10489,N_11758);
nand U13144 (N_13144,N_8649,N_10914);
nand U13145 (N_13145,N_12324,N_6464);
or U13146 (N_13146,N_10883,N_7422);
xor U13147 (N_13147,N_7518,N_8540);
or U13148 (N_13148,N_11080,N_8020);
nor U13149 (N_13149,N_8884,N_9180);
nand U13150 (N_13150,N_9793,N_11569);
nor U13151 (N_13151,N_9646,N_11694);
or U13152 (N_13152,N_11392,N_9843);
nor U13153 (N_13153,N_11563,N_7554);
or U13154 (N_13154,N_6720,N_7816);
or U13155 (N_13155,N_10195,N_6624);
xnor U13156 (N_13156,N_9168,N_10539);
or U13157 (N_13157,N_10686,N_8172);
xor U13158 (N_13158,N_8018,N_8890);
or U13159 (N_13159,N_8851,N_6368);
or U13160 (N_13160,N_9926,N_7192);
xor U13161 (N_13161,N_9155,N_6656);
xor U13162 (N_13162,N_11298,N_11909);
nor U13163 (N_13163,N_10121,N_8697);
and U13164 (N_13164,N_8283,N_8855);
and U13165 (N_13165,N_7224,N_8896);
xnor U13166 (N_13166,N_6403,N_6689);
and U13167 (N_13167,N_10442,N_9441);
and U13168 (N_13168,N_7627,N_6721);
nand U13169 (N_13169,N_9530,N_8760);
nand U13170 (N_13170,N_7699,N_11700);
or U13171 (N_13171,N_10174,N_7819);
nand U13172 (N_13172,N_7851,N_9461);
and U13173 (N_13173,N_7758,N_10380);
or U13174 (N_13174,N_11515,N_11697);
or U13175 (N_13175,N_10643,N_10618);
or U13176 (N_13176,N_11685,N_9699);
and U13177 (N_13177,N_7465,N_9679);
xnor U13178 (N_13178,N_6558,N_8819);
and U13179 (N_13179,N_12160,N_10267);
nand U13180 (N_13180,N_8678,N_6303);
xnor U13181 (N_13181,N_10590,N_9868);
and U13182 (N_13182,N_7880,N_7294);
xor U13183 (N_13183,N_8069,N_12251);
nor U13184 (N_13184,N_10280,N_6366);
nand U13185 (N_13185,N_10252,N_10040);
xnor U13186 (N_13186,N_6718,N_11548);
and U13187 (N_13187,N_8326,N_6610);
xor U13188 (N_13188,N_10958,N_9632);
or U13189 (N_13189,N_12226,N_11114);
xnor U13190 (N_13190,N_11762,N_10402);
nor U13191 (N_13191,N_12048,N_12012);
and U13192 (N_13192,N_11157,N_12023);
xnor U13193 (N_13193,N_10201,N_7576);
or U13194 (N_13194,N_11989,N_6451);
and U13195 (N_13195,N_10672,N_9532);
nand U13196 (N_13196,N_11092,N_10913);
or U13197 (N_13197,N_6726,N_7306);
xnor U13198 (N_13198,N_11084,N_7400);
xnor U13199 (N_13199,N_10199,N_10196);
nor U13200 (N_13200,N_7823,N_9905);
and U13201 (N_13201,N_10825,N_6485);
nand U13202 (N_13202,N_12206,N_11949);
nand U13203 (N_13203,N_9986,N_9072);
xnor U13204 (N_13204,N_6561,N_12294);
and U13205 (N_13205,N_8615,N_11310);
and U13206 (N_13206,N_9672,N_11033);
and U13207 (N_13207,N_8875,N_10918);
xnor U13208 (N_13208,N_10530,N_10245);
and U13209 (N_13209,N_11221,N_12361);
xor U13210 (N_13210,N_10406,N_11444);
nand U13211 (N_13211,N_8732,N_9901);
and U13212 (N_13212,N_6947,N_9129);
xnor U13213 (N_13213,N_7373,N_9261);
and U13214 (N_13214,N_8246,N_9697);
nand U13215 (N_13215,N_10117,N_9436);
and U13216 (N_13216,N_8553,N_10456);
and U13217 (N_13217,N_9810,N_11422);
nor U13218 (N_13218,N_10805,N_6678);
xnor U13219 (N_13219,N_9278,N_8346);
nand U13220 (N_13220,N_7123,N_10683);
xor U13221 (N_13221,N_6617,N_7241);
or U13222 (N_13222,N_8131,N_12237);
nor U13223 (N_13223,N_6425,N_9071);
xnor U13224 (N_13224,N_9733,N_8318);
xor U13225 (N_13225,N_12126,N_6503);
or U13226 (N_13226,N_7771,N_9691);
or U13227 (N_13227,N_9723,N_11873);
xor U13228 (N_13228,N_11981,N_10404);
or U13229 (N_13229,N_10928,N_12387);
nor U13230 (N_13230,N_11588,N_8734);
and U13231 (N_13231,N_10328,N_8504);
and U13232 (N_13232,N_9123,N_6866);
and U13233 (N_13233,N_10526,N_10587);
xor U13234 (N_13234,N_6257,N_9351);
xnor U13235 (N_13235,N_7353,N_11790);
and U13236 (N_13236,N_10244,N_11644);
nand U13237 (N_13237,N_6742,N_6616);
and U13238 (N_13238,N_7581,N_11590);
nand U13239 (N_13239,N_9608,N_7955);
and U13240 (N_13240,N_7423,N_7963);
nor U13241 (N_13241,N_9521,N_8665);
and U13242 (N_13242,N_8378,N_9991);
xnor U13243 (N_13243,N_8144,N_10047);
or U13244 (N_13244,N_8232,N_6805);
nor U13245 (N_13245,N_11109,N_10580);
xnor U13246 (N_13246,N_9406,N_11583);
xnor U13247 (N_13247,N_10255,N_7639);
or U13248 (N_13248,N_12418,N_6565);
xnor U13249 (N_13249,N_6395,N_9427);
or U13250 (N_13250,N_9473,N_7741);
and U13251 (N_13251,N_7356,N_7264);
or U13252 (N_13252,N_10094,N_8448);
and U13253 (N_13253,N_8436,N_11691);
xor U13254 (N_13254,N_12352,N_9456);
nand U13255 (N_13255,N_11714,N_6527);
nand U13256 (N_13256,N_8158,N_6929);
and U13257 (N_13257,N_11318,N_11581);
nor U13258 (N_13258,N_11445,N_12095);
and U13259 (N_13259,N_9214,N_8124);
or U13260 (N_13260,N_10111,N_8828);
or U13261 (N_13261,N_10066,N_7489);
or U13262 (N_13262,N_11297,N_7804);
or U13263 (N_13263,N_11147,N_8183);
and U13264 (N_13264,N_6861,N_9902);
and U13265 (N_13265,N_10067,N_10570);
and U13266 (N_13266,N_12466,N_9003);
and U13267 (N_13267,N_6838,N_8288);
or U13268 (N_13268,N_7533,N_8938);
and U13269 (N_13269,N_7367,N_7173);
nand U13270 (N_13270,N_11481,N_9366);
or U13271 (N_13271,N_7678,N_8127);
or U13272 (N_13272,N_9605,N_8822);
nor U13273 (N_13273,N_9251,N_10435);
nor U13274 (N_13274,N_10696,N_10980);
xor U13275 (N_13275,N_9636,N_6990);
or U13276 (N_13276,N_7194,N_12431);
xor U13277 (N_13277,N_8189,N_11643);
and U13278 (N_13278,N_12092,N_12320);
nor U13279 (N_13279,N_11755,N_11926);
and U13280 (N_13280,N_11571,N_8498);
xnor U13281 (N_13281,N_11925,N_7534);
xnor U13282 (N_13282,N_11365,N_10528);
nand U13283 (N_13283,N_7507,N_10390);
or U13284 (N_13284,N_11847,N_9045);
nor U13285 (N_13285,N_11138,N_10419);
nand U13286 (N_13286,N_12062,N_6622);
or U13287 (N_13287,N_11108,N_8276);
nor U13288 (N_13288,N_8631,N_11267);
or U13289 (N_13289,N_7779,N_10123);
nor U13290 (N_13290,N_8294,N_10873);
or U13291 (N_13291,N_12190,N_6588);
or U13292 (N_13292,N_11503,N_9576);
or U13293 (N_13293,N_11442,N_12181);
and U13294 (N_13294,N_6723,N_10611);
xor U13295 (N_13295,N_7495,N_11622);
or U13296 (N_13296,N_11125,N_6274);
nand U13297 (N_13297,N_7505,N_10215);
nor U13298 (N_13298,N_12231,N_7301);
xnor U13299 (N_13299,N_8451,N_7897);
xnor U13300 (N_13300,N_8716,N_10710);
nor U13301 (N_13301,N_8110,N_10905);
nor U13302 (N_13302,N_11589,N_11906);
or U13303 (N_13303,N_6981,N_11200);
nand U13304 (N_13304,N_8609,N_9930);
nor U13305 (N_13305,N_6912,N_10132);
nor U13306 (N_13306,N_12347,N_11962);
xnor U13307 (N_13307,N_9259,N_11093);
and U13308 (N_13308,N_8887,N_12085);
or U13309 (N_13309,N_11288,N_10869);
nor U13310 (N_13310,N_12002,N_8044);
nand U13311 (N_13311,N_6789,N_6770);
xor U13312 (N_13312,N_10957,N_9064);
or U13313 (N_13313,N_8601,N_11461);
or U13314 (N_13314,N_12001,N_8571);
or U13315 (N_13315,N_8356,N_8642);
nand U13316 (N_13316,N_11386,N_12019);
xor U13317 (N_13317,N_12106,N_11504);
or U13318 (N_13318,N_8694,N_6259);
or U13319 (N_13319,N_11218,N_9750);
or U13320 (N_13320,N_10653,N_10865);
nor U13321 (N_13321,N_10362,N_7630);
or U13322 (N_13322,N_9146,N_8507);
and U13323 (N_13323,N_8314,N_8864);
nor U13324 (N_13324,N_6713,N_8402);
and U13325 (N_13325,N_10633,N_6301);
nor U13326 (N_13326,N_6657,N_8212);
nand U13327 (N_13327,N_8438,N_8009);
and U13328 (N_13328,N_7671,N_11499);
and U13329 (N_13329,N_11152,N_12000);
xnor U13330 (N_13330,N_12353,N_11132);
and U13331 (N_13331,N_11491,N_7836);
nand U13332 (N_13332,N_10604,N_11766);
or U13333 (N_13333,N_8628,N_7090);
xnor U13334 (N_13334,N_6349,N_7157);
or U13335 (N_13335,N_11322,N_9276);
xnor U13336 (N_13336,N_9065,N_8325);
xor U13337 (N_13337,N_12239,N_8648);
xor U13338 (N_13338,N_8570,N_12187);
and U13339 (N_13339,N_11718,N_8711);
nand U13340 (N_13340,N_12398,N_7366);
nor U13341 (N_13341,N_10606,N_7220);
nor U13342 (N_13342,N_7711,N_6361);
xor U13343 (N_13343,N_9565,N_10281);
nand U13344 (N_13344,N_8612,N_7497);
and U13345 (N_13345,N_10717,N_10102);
nor U13346 (N_13346,N_9752,N_6885);
xor U13347 (N_13347,N_9070,N_8479);
nor U13348 (N_13348,N_11551,N_10343);
nor U13349 (N_13349,N_9079,N_10859);
xnor U13350 (N_13350,N_9303,N_7372);
nor U13351 (N_13351,N_9921,N_6823);
or U13352 (N_13352,N_9654,N_12435);
nand U13353 (N_13353,N_10756,N_12309);
nor U13354 (N_13354,N_8109,N_6276);
xor U13355 (N_13355,N_8462,N_6707);
xnor U13356 (N_13356,N_11301,N_12234);
xnor U13357 (N_13357,N_8630,N_12169);
and U13358 (N_13358,N_6294,N_11453);
or U13359 (N_13359,N_9919,N_8241);
nand U13360 (N_13360,N_12139,N_6319);
nand U13361 (N_13361,N_12404,N_8091);
xor U13362 (N_13362,N_10940,N_6316);
or U13363 (N_13363,N_7290,N_9782);
or U13364 (N_13364,N_12020,N_10867);
nor U13365 (N_13365,N_11897,N_11174);
xor U13366 (N_13366,N_7885,N_8800);
xor U13367 (N_13367,N_9352,N_8000);
and U13368 (N_13368,N_8635,N_6827);
nor U13369 (N_13369,N_6841,N_10399);
nand U13370 (N_13370,N_10420,N_7203);
nor U13371 (N_13371,N_6835,N_10320);
and U13372 (N_13372,N_8753,N_7370);
xnor U13373 (N_13373,N_8386,N_7396);
xnor U13374 (N_13374,N_8412,N_9544);
and U13375 (N_13375,N_11495,N_9321);
nand U13376 (N_13376,N_11421,N_8650);
and U13377 (N_13377,N_10621,N_9175);
or U13378 (N_13378,N_6711,N_11646);
nand U13379 (N_13379,N_7139,N_9857);
nor U13380 (N_13380,N_8696,N_6358);
nand U13381 (N_13381,N_7088,N_9932);
nor U13382 (N_13382,N_9923,N_8445);
nor U13383 (N_13383,N_9874,N_10270);
nand U13384 (N_13384,N_10855,N_11019);
nor U13385 (N_13385,N_8340,N_11010);
xor U13386 (N_13386,N_7089,N_11647);
nand U13387 (N_13387,N_10473,N_11426);
and U13388 (N_13388,N_11259,N_9193);
nor U13389 (N_13389,N_10187,N_7928);
xor U13390 (N_13390,N_6673,N_10135);
xor U13391 (N_13391,N_7096,N_9145);
or U13392 (N_13392,N_10735,N_11395);
xnor U13393 (N_13393,N_12162,N_7181);
or U13394 (N_13394,N_6373,N_10272);
and U13395 (N_13395,N_8151,N_7217);
nand U13396 (N_13396,N_8173,N_11679);
or U13397 (N_13397,N_9368,N_8541);
xnor U13398 (N_13398,N_12288,N_12374);
or U13399 (N_13399,N_11514,N_10925);
nand U13400 (N_13400,N_11761,N_9973);
nor U13401 (N_13401,N_12256,N_6730);
nand U13402 (N_13402,N_7947,N_7053);
nor U13403 (N_13403,N_11014,N_6354);
nor U13404 (N_13404,N_7049,N_9591);
xor U13405 (N_13405,N_10845,N_10059);
and U13406 (N_13406,N_11466,N_8108);
nor U13407 (N_13407,N_6854,N_9536);
nand U13408 (N_13408,N_11326,N_8149);
and U13409 (N_13409,N_12067,N_7547);
or U13410 (N_13410,N_6330,N_10237);
or U13411 (N_13411,N_12099,N_8809);
nor U13412 (N_13412,N_7939,N_10617);
or U13413 (N_13413,N_8651,N_9362);
and U13414 (N_13414,N_10823,N_10130);
or U13415 (N_13415,N_6407,N_8598);
or U13416 (N_13416,N_12391,N_10513);
or U13417 (N_13417,N_6982,N_6736);
nor U13418 (N_13418,N_11465,N_7706);
xor U13419 (N_13419,N_11266,N_7929);
nor U13420 (N_13420,N_12121,N_7513);
and U13421 (N_13421,N_11111,N_8931);
nor U13422 (N_13422,N_12295,N_11530);
nor U13423 (N_13423,N_8515,N_10979);
xnor U13424 (N_13424,N_9354,N_11069);
nor U13425 (N_13425,N_7488,N_11312);
and U13426 (N_13426,N_8469,N_10950);
or U13427 (N_13427,N_11698,N_12419);
xnor U13428 (N_13428,N_9773,N_8762);
xor U13429 (N_13429,N_11314,N_10303);
xor U13430 (N_13430,N_10554,N_11850);
nand U13431 (N_13431,N_9008,N_10057);
xnor U13432 (N_13432,N_11754,N_9177);
xnor U13433 (N_13433,N_6260,N_7729);
xor U13434 (N_13434,N_6814,N_10898);
and U13435 (N_13435,N_7399,N_12350);
and U13436 (N_13436,N_8764,N_6977);
or U13437 (N_13437,N_10410,N_12238);
or U13438 (N_13438,N_6978,N_9909);
and U13439 (N_13439,N_7392,N_10605);
and U13440 (N_13440,N_6645,N_11948);
nor U13441 (N_13441,N_10157,N_6601);
xnor U13442 (N_13442,N_12259,N_6817);
nor U13443 (N_13443,N_7775,N_11277);
nand U13444 (N_13444,N_7769,N_11921);
nand U13445 (N_13445,N_8403,N_8064);
nand U13446 (N_13446,N_10891,N_11621);
or U13447 (N_13447,N_11390,N_8936);
nor U13448 (N_13448,N_12217,N_11829);
and U13449 (N_13449,N_10616,N_8980);
and U13450 (N_13450,N_9455,N_9526);
xnor U13451 (N_13451,N_7415,N_6268);
and U13452 (N_13452,N_7070,N_11334);
and U13453 (N_13453,N_8749,N_12254);
and U13454 (N_13454,N_9415,N_10931);
nand U13455 (N_13455,N_12064,N_6453);
or U13456 (N_13456,N_9088,N_6815);
or U13457 (N_13457,N_7792,N_9171);
nor U13458 (N_13458,N_10006,N_7189);
nor U13459 (N_13459,N_9794,N_8145);
and U13460 (N_13460,N_9717,N_11995);
or U13461 (N_13461,N_9563,N_11149);
and U13462 (N_13462,N_8070,N_9299);
nand U13463 (N_13463,N_12422,N_9774);
xor U13464 (N_13464,N_6900,N_6381);
xnor U13465 (N_13465,N_8567,N_10609);
nor U13466 (N_13466,N_8227,N_11494);
and U13467 (N_13467,N_11400,N_9481);
or U13468 (N_13468,N_10999,N_7943);
nand U13469 (N_13469,N_11306,N_6778);
xor U13470 (N_13470,N_12263,N_6347);
and U13471 (N_13471,N_8981,N_12289);
nand U13472 (N_13472,N_7412,N_7072);
nand U13473 (N_13473,N_8474,N_12334);
nor U13474 (N_13474,N_11278,N_6649);
or U13475 (N_13475,N_9743,N_10256);
nor U13476 (N_13476,N_10534,N_7150);
nand U13477 (N_13477,N_7592,N_8932);
and U13478 (N_13478,N_6462,N_11035);
and U13479 (N_13479,N_12384,N_6753);
and U13480 (N_13480,N_7931,N_10413);
and U13481 (N_13481,N_10056,N_6506);
xnor U13482 (N_13482,N_12433,N_11477);
and U13483 (N_13483,N_10573,N_7676);
nand U13484 (N_13484,N_10701,N_10824);
nor U13485 (N_13485,N_8892,N_8083);
xnor U13486 (N_13486,N_8526,N_8050);
nor U13487 (N_13487,N_7633,N_11025);
xnor U13488 (N_13488,N_9112,N_12495);
nand U13489 (N_13489,N_11868,N_6352);
xor U13490 (N_13490,N_11997,N_9335);
nand U13491 (N_13491,N_9485,N_10418);
nand U13492 (N_13492,N_9737,N_9104);
and U13493 (N_13493,N_6917,N_8218);
xor U13494 (N_13494,N_12488,N_9226);
nor U13495 (N_13495,N_10908,N_10355);
nand U13496 (N_13496,N_9952,N_10455);
nand U13497 (N_13497,N_8873,N_7131);
xor U13498 (N_13498,N_6435,N_11345);
nor U13499 (N_13499,N_10301,N_12299);
and U13500 (N_13500,N_7178,N_8535);
and U13501 (N_13501,N_11245,N_12297);
or U13502 (N_13502,N_8427,N_11479);
or U13503 (N_13503,N_11553,N_11520);
and U13504 (N_13504,N_6623,N_6253);
or U13505 (N_13505,N_7199,N_9945);
xor U13506 (N_13506,N_7980,N_6348);
nand U13507 (N_13507,N_6489,N_9157);
nand U13508 (N_13508,N_10798,N_11087);
nand U13509 (N_13509,N_10543,N_7020);
or U13510 (N_13510,N_10722,N_10850);
nand U13511 (N_13511,N_9785,N_12364);
or U13512 (N_13512,N_7990,N_8279);
xnor U13513 (N_13513,N_9022,N_10125);
nand U13514 (N_13514,N_7358,N_9592);
or U13515 (N_13515,N_9682,N_10105);
xnor U13516 (N_13516,N_7790,N_8959);
nand U13517 (N_13517,N_10785,N_10021);
and U13518 (N_13518,N_6792,N_12489);
or U13519 (N_13519,N_11568,N_11591);
xor U13520 (N_13520,N_10602,N_12202);
or U13521 (N_13521,N_11565,N_10361);
nand U13522 (N_13522,N_7713,N_10874);
nor U13523 (N_13523,N_8548,N_6519);
nor U13524 (N_13524,N_10385,N_9895);
and U13525 (N_13525,N_10856,N_6754);
and U13526 (N_13526,N_8181,N_8934);
xnor U13527 (N_13527,N_9616,N_8573);
and U13528 (N_13528,N_8554,N_10407);
and U13529 (N_13529,N_11523,N_12339);
nor U13530 (N_13530,N_8789,N_7109);
xor U13531 (N_13531,N_12038,N_9331);
nand U13532 (N_13532,N_8848,N_7427);
xnor U13533 (N_13533,N_9813,N_7299);
and U13534 (N_13534,N_9053,N_8861);
and U13535 (N_13535,N_7696,N_8997);
and U13536 (N_13536,N_11472,N_12113);
and U13537 (N_13537,N_8188,N_11429);
xnor U13538 (N_13538,N_12359,N_10853);
and U13539 (N_13539,N_11954,N_8019);
or U13540 (N_13540,N_11794,N_9474);
nand U13541 (N_13541,N_8437,N_9822);
and U13542 (N_13542,N_6267,N_11287);
nor U13543 (N_13543,N_9727,N_8969);
nor U13544 (N_13544,N_7434,N_6799);
nand U13545 (N_13545,N_8944,N_12428);
xor U13546 (N_13546,N_8012,N_9081);
xnor U13547 (N_13547,N_10321,N_12354);
xor U13548 (N_13548,N_8568,N_8174);
and U13549 (N_13549,N_12123,N_11451);
or U13550 (N_13550,N_7756,N_11057);
nand U13551 (N_13551,N_8228,N_10185);
nand U13552 (N_13552,N_10982,N_7824);
xor U13553 (N_13553,N_9466,N_8599);
nand U13554 (N_13554,N_7032,N_9150);
or U13555 (N_13555,N_8658,N_12197);
or U13556 (N_13556,N_8943,N_7764);
or U13557 (N_13557,N_10104,N_7114);
nand U13558 (N_13558,N_9212,N_10563);
or U13559 (N_13559,N_6356,N_6333);
xor U13560 (N_13560,N_6620,N_6948);
nand U13561 (N_13561,N_10966,N_11341);
xor U13562 (N_13562,N_6898,N_7935);
nand U13563 (N_13563,N_11399,N_11182);
xnor U13564 (N_13564,N_11036,N_7572);
or U13565 (N_13565,N_7349,N_8605);
xor U13566 (N_13566,N_6630,N_6833);
or U13567 (N_13567,N_8076,N_11768);
and U13568 (N_13568,N_6615,N_9924);
xnor U13569 (N_13569,N_10575,N_10367);
nor U13570 (N_13570,N_7649,N_12142);
nand U13571 (N_13571,N_8937,N_7517);
nand U13572 (N_13572,N_8457,N_9638);
nor U13573 (N_13573,N_11366,N_9256);
nor U13574 (N_13574,N_12159,N_10887);
nand U13575 (N_13575,N_7324,N_9589);
xnor U13576 (N_13576,N_9059,N_7918);
xor U13577 (N_13577,N_8690,N_6315);
or U13578 (N_13578,N_11211,N_10220);
xnor U13579 (N_13579,N_7431,N_7862);
and U13580 (N_13580,N_10919,N_9904);
or U13581 (N_13581,N_7761,N_6954);
nor U13582 (N_13582,N_6728,N_9110);
or U13583 (N_13583,N_6937,N_10888);
nand U13584 (N_13584,N_9228,N_7256);
nand U13585 (N_13585,N_9083,N_9194);
xnor U13586 (N_13586,N_8446,N_6559);
nor U13587 (N_13587,N_11864,N_6749);
nor U13588 (N_13588,N_6400,N_11896);
and U13589 (N_13589,N_6968,N_7483);
and U13590 (N_13590,N_10058,N_11133);
and U13591 (N_13591,N_9967,N_6295);
nor U13592 (N_13592,N_7957,N_7357);
xnor U13593 (N_13593,N_9241,N_10208);
xnor U13594 (N_13594,N_9816,N_7958);
xnor U13595 (N_13595,N_11901,N_6292);
nor U13596 (N_13596,N_9382,N_6636);
or U13597 (N_13597,N_10684,N_9404);
or U13598 (N_13598,N_7875,N_9229);
nand U13599 (N_13599,N_10497,N_7337);
and U13600 (N_13600,N_9394,N_7273);
or U13601 (N_13601,N_9855,N_6697);
nor U13602 (N_13602,N_10358,N_10042);
nand U13603 (N_13603,N_7323,N_11176);
and U13604 (N_13604,N_8415,N_7515);
nor U13605 (N_13605,N_10571,N_10053);
or U13606 (N_13606,N_11631,N_11911);
nor U13607 (N_13607,N_7691,N_11078);
or U13608 (N_13608,N_9664,N_12192);
nor U13609 (N_13609,N_11640,N_8220);
or U13610 (N_13610,N_9283,N_8426);
nor U13611 (N_13611,N_11201,N_6635);
xnor U13612 (N_13612,N_8285,N_8922);
nor U13613 (N_13613,N_9890,N_9788);
and U13614 (N_13614,N_8073,N_12054);
or U13615 (N_13615,N_11938,N_8603);
xnor U13616 (N_13616,N_11722,N_6705);
xor U13617 (N_13617,N_11971,N_12228);
xor U13618 (N_13618,N_8214,N_11615);
nand U13619 (N_13619,N_6324,N_6880);
nor U13620 (N_13620,N_9656,N_9825);
nand U13621 (N_13621,N_8234,N_10166);
xor U13622 (N_13622,N_7838,N_12144);
xor U13623 (N_13623,N_6752,N_11497);
xnor U13624 (N_13624,N_12136,N_11967);
nor U13625 (N_13625,N_10110,N_8952);
or U13626 (N_13626,N_7055,N_7705);
nand U13627 (N_13627,N_7169,N_6496);
nor U13628 (N_13628,N_10627,N_12308);
nor U13629 (N_13629,N_11203,N_10574);
or U13630 (N_13630,N_9978,N_9060);
xor U13631 (N_13631,N_7951,N_9738);
nand U13632 (N_13632,N_11773,N_9258);
and U13633 (N_13633,N_6696,N_10458);
or U13634 (N_13634,N_8721,N_7275);
or U13635 (N_13635,N_9189,N_8708);
and U13636 (N_13636,N_8377,N_8671);
and U13637 (N_13637,N_10504,N_10316);
or U13638 (N_13638,N_8001,N_10374);
nor U13639 (N_13639,N_7835,N_9620);
nand U13640 (N_13640,N_8235,N_10086);
nor U13641 (N_13641,N_8569,N_11535);
nor U13642 (N_13642,N_9484,N_8368);
nand U13643 (N_13643,N_8676,N_6712);
or U13644 (N_13644,N_10164,N_8562);
nand U13645 (N_13645,N_7308,N_11226);
nor U13646 (N_13646,N_10970,N_9683);
nand U13647 (N_13647,N_11977,N_12250);
nand U13648 (N_13648,N_11067,N_10459);
xnor U13649 (N_13649,N_8953,N_7122);
xor U13650 (N_13650,N_10638,N_6991);
nand U13651 (N_13651,N_12283,N_12120);
xnor U13652 (N_13652,N_10858,N_10516);
and U13653 (N_13653,N_6438,N_9254);
or U13654 (N_13654,N_8169,N_11032);
or U13655 (N_13655,N_6538,N_10566);
and U13656 (N_13656,N_9999,N_9706);
nor U13657 (N_13657,N_9908,N_8614);
nand U13658 (N_13658,N_10816,N_9132);
and U13659 (N_13659,N_7818,N_10376);
or U13660 (N_13660,N_11167,N_6544);
nor U13661 (N_13661,N_7609,N_9016);
nand U13662 (N_13662,N_6568,N_9821);
xnor U13663 (N_13663,N_12323,N_6740);
or U13664 (N_13664,N_8486,N_10448);
or U13665 (N_13665,N_10732,N_12168);
nand U13666 (N_13666,N_9386,N_8858);
nand U13667 (N_13667,N_9345,N_8989);
nor U13668 (N_13668,N_6768,N_11249);
or U13669 (N_13669,N_7456,N_10794);
nand U13670 (N_13670,N_11263,N_7962);
nand U13671 (N_13671,N_11828,N_6543);
or U13672 (N_13672,N_9658,N_10012);
or U13673 (N_13673,N_11086,N_10688);
xor U13674 (N_13674,N_11826,N_10558);
nor U13675 (N_13675,N_11935,N_10782);
nor U13676 (N_13676,N_9928,N_12390);
xnor U13677 (N_13677,N_12031,N_8939);
xor U13678 (N_13678,N_12033,N_11202);
nor U13679 (N_13679,N_10339,N_8674);
xor U13680 (N_13680,N_6906,N_7243);
and U13681 (N_13681,N_12110,N_9903);
or U13682 (N_13682,N_6598,N_8834);
nand U13683 (N_13683,N_9906,N_9779);
xnor U13684 (N_13684,N_8868,N_12478);
or U13685 (N_13685,N_11855,N_11215);
and U13686 (N_13686,N_7435,N_6589);
nor U13687 (N_13687,N_10932,N_7616);
nand U13688 (N_13688,N_12201,N_10603);
and U13689 (N_13689,N_8854,N_9033);
nand U13690 (N_13690,N_8534,N_9781);
or U13691 (N_13691,N_12311,N_9734);
and U13692 (N_13692,N_11813,N_6446);
nor U13693 (N_13693,N_8948,N_11602);
and U13694 (N_13694,N_10482,N_6677);
nor U13695 (N_13695,N_10962,N_11976);
and U13696 (N_13696,N_8754,N_7882);
nand U13697 (N_13697,N_7048,N_9217);
nor U13698 (N_13698,N_8543,N_10752);
or U13699 (N_13699,N_10400,N_6986);
or U13700 (N_13700,N_7809,N_6575);
xnor U13701 (N_13701,N_8844,N_11316);
xor U13702 (N_13702,N_10477,N_9117);
xor U13703 (N_13703,N_7802,N_6284);
and U13704 (N_13704,N_11183,N_7848);
xnor U13705 (N_13705,N_9783,N_10977);
nand U13706 (N_13706,N_9700,N_12018);
and U13707 (N_13707,N_10160,N_11062);
nand U13708 (N_13708,N_7227,N_10266);
nand U13709 (N_13709,N_9982,N_10242);
and U13710 (N_13710,N_12097,N_12182);
nand U13711 (N_13711,N_7643,N_8419);
xor U13712 (N_13712,N_8930,N_10801);
xnor U13713 (N_13713,N_11413,N_10424);
nand U13714 (N_13714,N_11737,N_9888);
nand U13715 (N_13715,N_6431,N_9216);
or U13716 (N_13716,N_7535,N_10276);
nand U13717 (N_13717,N_7914,N_8647);
nand U13718 (N_13718,N_6594,N_10133);
or U13719 (N_13719,N_6359,N_8252);
nor U13720 (N_13720,N_7403,N_11050);
nand U13721 (N_13721,N_6278,N_10522);
nor U13722 (N_13722,N_8138,N_8354);
and U13723 (N_13723,N_10465,N_7177);
and U13724 (N_13724,N_8964,N_8713);
or U13725 (N_13725,N_9580,N_12037);
nor U13726 (N_13726,N_9390,N_8004);
and U13727 (N_13727,N_7448,N_11524);
nor U13728 (N_13728,N_6806,N_11498);
or U13729 (N_13729,N_10545,N_9915);
nand U13730 (N_13730,N_8405,N_10797);
and U13731 (N_13731,N_11224,N_7340);
or U13732 (N_13732,N_7490,N_12013);
or U13733 (N_13733,N_8470,N_8746);
xor U13734 (N_13734,N_6600,N_8847);
xnor U13735 (N_13735,N_8418,N_7598);
xor U13736 (N_13736,N_8808,N_11117);
and U13737 (N_13737,N_9225,N_12473);
and U13738 (N_13738,N_9475,N_9980);
and U13739 (N_13739,N_10986,N_8903);
and U13740 (N_13740,N_8481,N_12274);
xnor U13741 (N_13741,N_10930,N_8529);
nand U13742 (N_13742,N_8146,N_6960);
and U13743 (N_13743,N_9953,N_7667);
and U13744 (N_13744,N_7569,N_9224);
or U13745 (N_13745,N_6942,N_11047);
or U13746 (N_13746,N_10800,N_12285);
nor U13747 (N_13747,N_6593,N_10849);
nor U13748 (N_13748,N_6872,N_10290);
and U13749 (N_13749,N_6679,N_7655);
xor U13750 (N_13750,N_8072,N_10542);
and U13751 (N_13751,N_8510,N_11907);
nor U13752 (N_13752,N_6591,N_7213);
nor U13753 (N_13753,N_9951,N_10077);
xor U13754 (N_13754,N_6533,N_7537);
nor U13755 (N_13755,N_9021,N_10572);
and U13756 (N_13756,N_10766,N_10389);
xnor U13757 (N_13757,N_12499,N_7045);
and U13758 (N_13758,N_11638,N_9911);
and U13759 (N_13759,N_9665,N_10461);
nor U13760 (N_13760,N_9615,N_11280);
nand U13761 (N_13761,N_12036,N_12386);
nor U13762 (N_13762,N_9000,N_6717);
and U13763 (N_13763,N_7499,N_6628);
and U13764 (N_13764,N_8238,N_11233);
or U13765 (N_13765,N_8455,N_9748);
nor U13766 (N_13766,N_9310,N_10436);
nor U13767 (N_13767,N_8024,N_10227);
nor U13768 (N_13768,N_8862,N_12496);
or U13769 (N_13769,N_7916,N_11975);
xor U13770 (N_13770,N_12477,N_6663);
and U13771 (N_13771,N_12049,N_12069);
nor U13772 (N_13772,N_8840,N_8941);
or U13773 (N_13773,N_9891,N_10779);
or U13774 (N_13774,N_10703,N_10239);
xnor U13775 (N_13775,N_6831,N_11474);
xnor U13776 (N_13776,N_11273,N_10562);
and U13777 (N_13777,N_7845,N_10462);
nand U13778 (N_13778,N_11468,N_6626);
and U13779 (N_13779,N_10988,N_10183);
nor U13780 (N_13780,N_9447,N_6399);
nand U13781 (N_13781,N_10758,N_11821);
and U13782 (N_13782,N_9346,N_12363);
and U13783 (N_13783,N_9492,N_7975);
or U13784 (N_13784,N_11882,N_6304);
and U13785 (N_13785,N_7033,N_7393);
nand U13786 (N_13786,N_10317,N_11705);
xnor U13787 (N_13787,N_9933,N_7041);
nand U13788 (N_13788,N_6766,N_12279);
nor U13789 (N_13789,N_6554,N_6899);
nand U13790 (N_13790,N_9359,N_7800);
and U13791 (N_13791,N_11554,N_7647);
or U13792 (N_13792,N_7681,N_12396);
xnor U13793 (N_13793,N_11876,N_11931);
xor U13794 (N_13794,N_11626,N_9710);
nand U13795 (N_13795,N_6341,N_11840);
nand U13796 (N_13796,N_7388,N_7441);
xor U13797 (N_13797,N_8132,N_10298);
xor U13798 (N_13798,N_7110,N_8079);
or U13799 (N_13799,N_11374,N_6918);
and U13800 (N_13800,N_8396,N_6501);
xor U13801 (N_13801,N_7587,N_7144);
and U13802 (N_13802,N_7010,N_7538);
or U13803 (N_13803,N_10548,N_9471);
xnor U13804 (N_13804,N_6914,N_10345);
or U13805 (N_13805,N_7811,N_11247);
nand U13806 (N_13806,N_9990,N_8248);
nand U13807 (N_13807,N_8315,N_7170);
and U13808 (N_13808,N_11090,N_8528);
nand U13809 (N_13809,N_10368,N_10091);
and U13810 (N_13810,N_11525,N_9140);
nand U13811 (N_13811,N_10679,N_7596);
and U13812 (N_13812,N_9424,N_11064);
nor U13813 (N_13813,N_12446,N_11648);
nor U13814 (N_13814,N_12349,N_10163);
nand U13815 (N_13815,N_9324,N_6690);
and U13816 (N_13816,N_10207,N_11819);
nand U13817 (N_13817,N_9808,N_6949);
nor U13818 (N_13818,N_9041,N_8395);
and U13819 (N_13819,N_7514,N_10096);
nand U13820 (N_13820,N_10128,N_10902);
nand U13821 (N_13821,N_10576,N_12039);
nor U13822 (N_13822,N_6609,N_8692);
nand U13823 (N_13823,N_6820,N_11269);
or U13824 (N_13824,N_6846,N_8488);
or U13825 (N_13825,N_7788,N_8322);
and U13826 (N_13826,N_10471,N_9454);
or U13827 (N_13827,N_12480,N_7247);
nor U13828 (N_13828,N_7197,N_7176);
nor U13829 (N_13829,N_7073,N_11541);
or U13830 (N_13830,N_11952,N_9854);
xor U13831 (N_13831,N_12479,N_6944);
nor U13832 (N_13832,N_6255,N_8394);
nor U13833 (N_13833,N_12010,N_7182);
nand U13834 (N_13834,N_7417,N_11961);
xnor U13835 (N_13835,N_12434,N_10071);
nand U13836 (N_13836,N_9548,N_10594);
and U13837 (N_13837,N_8264,N_8619);
xnor U13838 (N_13838,N_8180,N_6998);
and U13839 (N_13839,N_9247,N_9449);
nor U13840 (N_13840,N_10646,N_11789);
nand U13841 (N_13841,N_11105,N_7712);
and U13842 (N_13842,N_6971,N_10900);
xor U13843 (N_13843,N_9993,N_7381);
nand U13844 (N_13844,N_8681,N_9414);
xor U13845 (N_13845,N_11920,N_9677);
nand U13846 (N_13846,N_10369,N_8372);
nor U13847 (N_13847,N_7632,N_8874);
or U13848 (N_13848,N_8806,N_12333);
and U13849 (N_13849,N_8735,N_8748);
or U13850 (N_13850,N_9739,N_8456);
and U13851 (N_13851,N_8267,N_11998);
and U13852 (N_13852,N_7438,N_7050);
nor U13853 (N_13853,N_9105,N_8115);
and U13854 (N_13854,N_6528,N_12042);
nand U13855 (N_13855,N_9519,N_9838);
and U13856 (N_13856,N_11000,N_10490);
nor U13857 (N_13857,N_11005,N_9892);
or U13858 (N_13858,N_9204,N_7244);
xnor U13859 (N_13859,N_6443,N_11502);
or U13860 (N_13860,N_9042,N_6338);
nand U13861 (N_13861,N_11905,N_8411);
nor U13862 (N_13862,N_10536,N_11536);
or U13863 (N_13863,N_8663,N_11391);
or U13864 (N_13864,N_10363,N_8490);
nand U13865 (N_13865,N_6969,N_11169);
or U13866 (N_13866,N_9200,N_10781);
nor U13867 (N_13867,N_11531,N_9645);
or U13868 (N_13868,N_9539,N_10592);
or U13869 (N_13869,N_7798,N_7703);
or U13870 (N_13870,N_11542,N_7815);
nand U13871 (N_13871,N_12408,N_12257);
and U13872 (N_13872,N_8582,N_8424);
and U13873 (N_13873,N_11199,N_9568);
nor U13874 (N_13874,N_9446,N_9128);
nand U13875 (N_13875,N_11328,N_10388);
and U13876 (N_13876,N_12006,N_7797);
and U13877 (N_13877,N_11346,N_10650);
nand U13878 (N_13878,N_11081,N_10050);
nand U13879 (N_13879,N_8199,N_7641);
nand U13880 (N_13880,N_6418,N_8304);
nor U13881 (N_13881,N_11351,N_7269);
xnor U13882 (N_13882,N_6507,N_8122);
nor U13883 (N_13883,N_9566,N_11872);
or U13884 (N_13884,N_7205,N_7876);
or U13885 (N_13885,N_8016,N_12132);
xor U13886 (N_13886,N_10499,N_12174);
nand U13887 (N_13887,N_12065,N_7985);
xor U13888 (N_13888,N_7103,N_9800);
nor U13889 (N_13889,N_10540,N_7000);
nand U13890 (N_13890,N_7571,N_9227);
or U13891 (N_13891,N_7674,N_12215);
nand U13892 (N_13892,N_10444,N_10182);
xnor U13893 (N_13893,N_8992,N_7202);
or U13894 (N_13894,N_11459,N_10391);
and U13895 (N_13895,N_11213,N_8843);
and U13896 (N_13896,N_11289,N_6801);
and U13897 (N_13897,N_6510,N_12302);
xnor U13898 (N_13898,N_10383,N_7826);
xnor U13899 (N_13899,N_10061,N_7326);
and U13900 (N_13900,N_11060,N_9325);
and U13901 (N_13901,N_7822,N_9789);
or U13902 (N_13902,N_9764,N_8429);
xnor U13903 (N_13903,N_6973,N_10654);
or U13904 (N_13904,N_11151,N_7839);
or U13905 (N_13905,N_9383,N_11352);
and U13906 (N_13906,N_8563,N_8203);
nor U13907 (N_13907,N_6813,N_12167);
xor U13908 (N_13908,N_11576,N_6461);
and U13909 (N_13909,N_9918,N_7552);
nor U13910 (N_13910,N_6560,N_9439);
or U13911 (N_13911,N_10685,N_6322);
or U13912 (N_13912,N_11804,N_7272);
nor U13913 (N_13913,N_8006,N_8484);
or U13914 (N_13914,N_6776,N_9775);
and U13915 (N_13915,N_11972,N_8618);
or U13916 (N_13916,N_12292,N_11875);
and U13917 (N_13917,N_6308,N_8531);
xnor U13918 (N_13918,N_11599,N_8502);
nor U13919 (N_13919,N_8239,N_10582);
nand U13920 (N_13920,N_8801,N_10124);
nand U13921 (N_13921,N_8213,N_11177);
nand U13922 (N_13922,N_12225,N_11293);
xnor U13923 (N_13923,N_6708,N_7061);
nand U13924 (N_13924,N_6585,N_6727);
xnor U13925 (N_13925,N_11837,N_12457);
or U13926 (N_13926,N_10747,N_9048);
nand U13927 (N_13927,N_12140,N_9486);
xor U13928 (N_13928,N_12214,N_7152);
nor U13929 (N_13929,N_12212,N_11684);
or U13930 (N_13930,N_6313,N_9218);
xnor U13931 (N_13931,N_11378,N_7531);
nor U13932 (N_13932,N_6980,N_6921);
or U13933 (N_13933,N_9121,N_10176);
nand U13934 (N_13934,N_10879,N_10544);
xor U13935 (N_13935,N_11903,N_10481);
or U13936 (N_13936,N_12385,N_11751);
nand U13937 (N_13937,N_7146,N_8296);
and U13938 (N_13938,N_8423,N_8768);
and U13939 (N_13939,N_10377,N_7735);
or U13940 (N_13940,N_7727,N_8636);
xor U13941 (N_13941,N_10129,N_6545);
nand U13942 (N_13942,N_10069,N_6254);
xnor U13943 (N_13943,N_9419,N_10933);
xnor U13944 (N_13944,N_7158,N_7746);
and U13945 (N_13945,N_12066,N_7864);
xnor U13946 (N_13946,N_6702,N_11625);
or U13947 (N_13947,N_9111,N_9937);
and U13948 (N_13948,N_12362,N_9480);
nand U13949 (N_13949,N_10817,N_6339);
xnor U13950 (N_13950,N_10764,N_7394);
nand U13951 (N_13951,N_7494,N_11253);
nor U13952 (N_13952,N_9093,N_6513);
nor U13953 (N_13953,N_8519,N_9849);
nand U13954 (N_13954,N_10275,N_11798);
or U13955 (N_13955,N_12129,N_6759);
or U13956 (N_13956,N_7968,N_10894);
xnor U13957 (N_13957,N_9931,N_7766);
nand U13958 (N_13958,N_6704,N_9817);
or U13959 (N_13959,N_6796,N_11170);
xor U13960 (N_13960,N_11801,N_8812);
nand U13961 (N_13961,N_11435,N_9098);
nor U13962 (N_13962,N_9979,N_10230);
nand U13963 (N_13963,N_10191,N_10432);
xor U13964 (N_13964,N_9094,N_10001);
and U13965 (N_13965,N_9630,N_8955);
nand U13966 (N_13966,N_7780,N_12445);
nor U13967 (N_13967,N_7849,N_8499);
nor U13968 (N_13968,N_12004,N_10098);
nand U13969 (N_13969,N_6757,N_9757);
nand U13970 (N_13970,N_7570,N_6440);
and U13971 (N_13971,N_8467,N_10892);
nor U13972 (N_13972,N_12366,N_10938);
and U13973 (N_13973,N_6293,N_7884);
nand U13974 (N_13974,N_6271,N_6901);
or U13975 (N_13975,N_11916,N_11577);
or U13976 (N_13976,N_11377,N_6300);
xnor U13977 (N_13977,N_6746,N_8102);
and U13978 (N_13978,N_10248,N_8021);
xor U13979 (N_13979,N_7155,N_10662);
xor U13980 (N_13980,N_10716,N_9149);
xor U13981 (N_13981,N_12329,N_6950);
xnor U13982 (N_13982,N_7590,N_7398);
and U13983 (N_13983,N_9262,N_9987);
nand U13984 (N_13984,N_10247,N_7886);
nor U13985 (N_13985,N_11566,N_7714);
nand U13986 (N_13986,N_10249,N_10990);
xnor U13987 (N_13987,N_6335,N_10084);
or U13988 (N_13988,N_11963,N_9465);
xor U13989 (N_13989,N_6483,N_6367);
and U13990 (N_13990,N_6420,N_7106);
nor U13991 (N_13991,N_7915,N_7645);
or U13992 (N_13992,N_12173,N_9791);
nor U13993 (N_13993,N_9940,N_11617);
xnor U13994 (N_13994,N_8520,N_7895);
nor U13995 (N_13995,N_10386,N_8702);
nor U13996 (N_13996,N_8280,N_12372);
nand U13997 (N_13997,N_11116,N_7476);
nand U13998 (N_13998,N_8544,N_9054);
and U13999 (N_13999,N_8539,N_11791);
and U14000 (N_14000,N_11030,N_8375);
and U14001 (N_14001,N_7944,N_9845);
nand U14002 (N_14002,N_9044,N_10027);
and U14003 (N_14003,N_11835,N_7309);
nor U14004 (N_14004,N_10967,N_6436);
nand U14005 (N_14005,N_11252,N_10393);
xnor U14006 (N_14006,N_6323,N_7334);
or U14007 (N_14007,N_9130,N_11146);
xnor U14008 (N_14008,N_9718,N_7563);
nand U14009 (N_14009,N_7983,N_9043);
or U14010 (N_14010,N_10694,N_11193);
nor U14011 (N_14011,N_10158,N_6433);
nand U14012 (N_14012,N_11217,N_11376);
or U14013 (N_14013,N_6473,N_10331);
nand U14014 (N_14014,N_8097,N_11338);
and U14015 (N_14015,N_9453,N_7445);
nand U14016 (N_14016,N_10770,N_11982);
xnor U14017 (N_14017,N_11110,N_11353);
nor U14018 (N_14018,N_8114,N_7175);
nor U14019 (N_14019,N_6660,N_10214);
nand U14020 (N_14020,N_9676,N_10624);
nand U14021 (N_14021,N_7015,N_8640);
and U14022 (N_14022,N_7843,N_9747);
and U14023 (N_14023,N_10881,N_8505);
nand U14024 (N_14024,N_9056,N_8054);
nand U14025 (N_14025,N_9663,N_7744);
xor U14026 (N_14026,N_6320,N_9304);
nor U14027 (N_14027,N_12128,N_7022);
and U14028 (N_14028,N_10976,N_9440);
nor U14029 (N_14029,N_8308,N_12204);
nand U14030 (N_14030,N_12016,N_6515);
and U14031 (N_14031,N_9692,N_8305);
and U14032 (N_14032,N_9712,N_11271);
xnor U14033 (N_14033,N_10860,N_6279);
or U14034 (N_14034,N_10017,N_11385);
xor U14035 (N_14035,N_11469,N_8958);
xor U14036 (N_14036,N_10020,N_12107);
nand U14037 (N_14037,N_9167,N_9853);
and U14038 (N_14038,N_10946,N_11018);
or U14039 (N_14039,N_9848,N_10257);
xnor U14040 (N_14040,N_10070,N_6457);
or U14041 (N_14041,N_10101,N_12316);
nor U14042 (N_14042,N_10289,N_11370);
nand U14043 (N_14043,N_8833,N_8159);
xnor U14044 (N_14044,N_8865,N_10005);
nor U14045 (N_14045,N_7315,N_11205);
and U14046 (N_14046,N_10953,N_10668);
or U14047 (N_14047,N_9777,N_9378);
xor U14048 (N_14048,N_9499,N_9085);
xor U14049 (N_14049,N_12083,N_7467);
or U14050 (N_14050,N_11707,N_10054);
and U14051 (N_14051,N_8365,N_6639);
nand U14052 (N_14052,N_8673,N_10277);
xor U14053 (N_14053,N_8259,N_9553);
or U14054 (N_14054,N_10579,N_6747);
nand U14055 (N_14055,N_11808,N_12246);
xnor U14056 (N_14056,N_9515,N_9374);
xor U14057 (N_14057,N_11958,N_11180);
and U14058 (N_14058,N_11623,N_12455);
nand U14059 (N_14059,N_7120,N_12412);
and U14060 (N_14060,N_7959,N_7428);
or U14061 (N_14061,N_8233,N_11951);
and U14062 (N_14062,N_7444,N_9220);
nor U14063 (N_14063,N_7601,N_7665);
nand U14064 (N_14064,N_8163,N_8273);
and U14065 (N_14065,N_11733,N_11107);
xor U14066 (N_14066,N_10711,N_10972);
xnor U14067 (N_14067,N_8061,N_12293);
xor U14068 (N_14068,N_8794,N_7909);
nor U14069 (N_14069,N_7461,N_10365);
xnor U14070 (N_14070,N_10099,N_7362);
and U14071 (N_14071,N_7065,N_7877);
nand U14072 (N_14072,N_8336,N_6972);
and U14073 (N_14073,N_7436,N_11880);
or U14074 (N_14074,N_11029,N_7785);
nor U14075 (N_14075,N_9581,N_7879);
nor U14076 (N_14076,N_9009,N_7126);
and U14077 (N_14077,N_6959,N_8752);
xnor U14078 (N_14078,N_7683,N_7023);
nand U14079 (N_14079,N_11142,N_6286);
nor U14080 (N_14080,N_7675,N_11545);
xnor U14081 (N_14081,N_7841,N_10143);
xnor U14082 (N_14082,N_9687,N_6686);
xor U14083 (N_14083,N_8011,N_10411);
nor U14084 (N_14084,N_10833,N_7021);
nor U14085 (N_14085,N_8829,N_7056);
nor U14086 (N_14086,N_11605,N_11441);
and U14087 (N_14087,N_9829,N_11732);
nor U14088 (N_14088,N_8473,N_7937);
nand U14089 (N_14089,N_10113,N_9762);
nor U14090 (N_14090,N_7354,N_7071);
or U14091 (N_14091,N_10998,N_9879);
nand U14092 (N_14092,N_11372,N_8537);
nand U14093 (N_14093,N_7054,N_7620);
xor U14094 (N_14094,N_6688,N_12091);
nor U14095 (N_14095,N_12205,N_8954);
or U14096 (N_14096,N_11046,N_10463);
xnor U14097 (N_14097,N_12088,N_7600);
xnor U14098 (N_14098,N_7578,N_6419);
or U14099 (N_14099,N_6934,N_9574);
xor U14100 (N_14100,N_9113,N_11416);
xnor U14101 (N_14101,N_10148,N_11344);
nor U14102 (N_14102,N_8857,N_7731);
nand U14103 (N_14103,N_10114,N_6340);
nand U14104 (N_14104,N_12483,N_12461);
xnor U14105 (N_14105,N_8928,N_7164);
nor U14106 (N_14106,N_7230,N_9369);
xnor U14107 (N_14107,N_10068,N_9488);
nor U14108 (N_14108,N_9315,N_7685);
xor U14109 (N_14109,N_6536,N_7652);
nor U14110 (N_14110,N_7342,N_11870);
and U14111 (N_14111,N_12180,N_10078);
or U14112 (N_14112,N_11489,N_10695);
or U14113 (N_14113,N_11154,N_12003);
and U14114 (N_14114,N_7452,N_10519);
and U14115 (N_14115,N_11216,N_11687);
nand U14116 (N_14116,N_12022,N_9037);
and U14117 (N_14117,N_8684,N_11313);
and U14118 (N_14118,N_12209,N_8281);
nor U14119 (N_14119,N_7722,N_7532);
xor U14120 (N_14120,N_8594,N_7721);
and U14121 (N_14121,N_9402,N_11300);
nand U14122 (N_14122,N_9385,N_8971);
nand U14123 (N_14123,N_6783,N_8803);
and U14124 (N_14124,N_10478,N_8747);
xnor U14125 (N_14125,N_6500,N_11229);
and U14126 (N_14126,N_7480,N_8087);
xnor U14127 (N_14127,N_10773,N_11884);
or U14128 (N_14128,N_9336,N_8441);
nand U14129 (N_14129,N_6331,N_10635);
nand U14130 (N_14130,N_9567,N_11095);
or U14131 (N_14131,N_7698,N_10838);
xor U14132 (N_14132,N_10241,N_10080);
xnor U14133 (N_14133,N_8750,N_8645);
nor U14134 (N_14134,N_8408,N_9462);
and U14135 (N_14135,N_9073,N_8777);
or U14136 (N_14136,N_10450,N_6940);
nor U14137 (N_14137,N_11136,N_6661);
nor U14138 (N_14138,N_10553,N_9736);
and U14139 (N_14139,N_8576,N_7522);
and U14140 (N_14140,N_10921,N_7724);
and U14141 (N_14141,N_11845,N_11708);
and U14142 (N_14142,N_8883,N_8717);
or U14143 (N_14143,N_6893,N_10512);
nand U14144 (N_14144,N_9824,N_7345);
or U14145 (N_14145,N_8074,N_11927);
xnor U14146 (N_14146,N_9651,N_9028);
xnor U14147 (N_14147,N_6280,N_9897);
xor U14148 (N_14148,N_9531,N_11243);
or U14149 (N_14149,N_11928,N_6430);
xnor U14150 (N_14150,N_7673,N_12165);
nor U14151 (N_14151,N_9869,N_9380);
nor U14152 (N_14152,N_11008,N_8831);
and U14153 (N_14153,N_9894,N_6631);
or U14154 (N_14154,N_7776,N_6428);
nor U14155 (N_14155,N_7079,N_9907);
nor U14156 (N_14156,N_11163,N_7455);
nor U14157 (N_14157,N_10956,N_11261);
nor U14158 (N_14158,N_9626,N_12356);
and U14159 (N_14159,N_12325,N_11883);
nor U14160 (N_14160,N_9705,N_10354);
or U14161 (N_14161,N_11543,N_11409);
nor U14162 (N_14162,N_7902,N_12427);
or U14163 (N_14163,N_11969,N_9534);
nand U14164 (N_14164,N_6958,N_10039);
xor U14165 (N_14165,N_8194,N_11996);
xnor U14166 (N_14166,N_9255,N_7277);
nor U14167 (N_14167,N_11866,N_11802);
nor U14168 (N_14168,N_11839,N_10652);
and U14169 (N_14169,N_11701,N_8946);
nor U14170 (N_14170,N_10395,N_9389);
nand U14171 (N_14171,N_9433,N_11172);
nand U14172 (N_14172,N_9329,N_8620);
nor U14173 (N_14173,N_7556,N_6552);
nand U14174 (N_14174,N_6523,N_7287);
or U14175 (N_14175,N_9377,N_11595);
nor U14176 (N_14176,N_11219,N_11127);
nor U14177 (N_14177,N_8041,N_6857);
nor U14178 (N_14178,N_6670,N_12484);
xor U14179 (N_14179,N_10942,N_10523);
and U14180 (N_14180,N_9092,N_9689);
or U14181 (N_14181,N_7786,N_11711);
nand U14182 (N_14182,N_11570,N_6889);
xnor U14183 (N_14183,N_12024,N_11321);
xnor U14184 (N_14184,N_10649,N_10808);
and U14185 (N_14185,N_8886,N_6767);
and U14186 (N_14186,N_8085,N_12378);
nor U14187 (N_14187,N_6621,N_8565);
nor U14188 (N_14188,N_12154,N_11636);
or U14189 (N_14189,N_10929,N_7907);
and U14190 (N_14190,N_8575,N_9643);
and U14191 (N_14191,N_11734,N_8966);
nand U14192 (N_14192,N_6377,N_6848);
xor U14193 (N_14193,N_6302,N_8784);
or U14194 (N_14194,N_7657,N_6797);
nor U14195 (N_14195,N_9542,N_11329);
nand U14196 (N_14196,N_7707,N_11103);
or U14197 (N_14197,N_11681,N_11908);
nor U14198 (N_14198,N_10323,N_10334);
xnor U14199 (N_14199,N_10055,N_8918);
nor U14200 (N_14200,N_6514,N_9806);
or U14201 (N_14201,N_6572,N_8195);
nand U14202 (N_14202,N_7140,N_9403);
nand U14203 (N_14203,N_9641,N_7283);
nor U14204 (N_14204,N_10480,N_12137);
nor U14205 (N_14205,N_11490,N_8333);
or U14206 (N_14206,N_6577,N_11282);
nor U14207 (N_14207,N_9160,N_11505);
xor U14208 (N_14208,N_12269,N_11881);
xnor U14209 (N_14209,N_9069,N_12300);
and U14210 (N_14210,N_9512,N_7377);
nor U14211 (N_14211,N_12194,N_12392);
nor U14212 (N_14212,N_12486,N_10744);
nand U14213 (N_14213,N_7191,N_6640);
and U14214 (N_14214,N_12147,N_11455);
nor U14215 (N_14215,N_11788,N_6448);
or U14216 (N_14216,N_12305,N_11616);
and U14217 (N_14217,N_8123,N_7282);
nor U14218 (N_14218,N_10861,N_11516);
nand U14219 (N_14219,N_10119,N_9097);
nor U14220 (N_14220,N_11781,N_12319);
nand U14221 (N_14221,N_11240,N_11037);
nor U14222 (N_14222,N_9910,N_6553);
and U14223 (N_14223,N_9057,N_11274);
or U14224 (N_14224,N_6390,N_8282);
xnor U14225 (N_14225,N_8413,N_10072);
or U14226 (N_14226,N_8965,N_11440);
or U14227 (N_14227,N_7565,N_11726);
nand U14228 (N_14228,N_7347,N_10663);
nor U14229 (N_14229,N_6722,N_6406);
xnor U14230 (N_14230,N_10359,N_8287);
xnor U14231 (N_14231,N_9840,N_8297);
nand U14232 (N_14232,N_7313,N_9203);
and U14233 (N_14233,N_9018,N_11210);
and U14234 (N_14234,N_8047,N_9472);
nand U14235 (N_14235,N_10678,N_8116);
nand U14236 (N_14236,N_12141,N_9522);
and U14237 (N_14237,N_9047,N_11946);
and U14238 (N_14238,N_7996,N_10912);
or U14239 (N_14239,N_6845,N_6840);
xor U14240 (N_14240,N_7127,N_10127);
nor U14241 (N_14241,N_10181,N_12096);
nand U14242 (N_14242,N_7919,N_6326);
nor U14243 (N_14243,N_6825,N_9337);
nand U14244 (N_14244,N_11692,N_7679);
nand U14245 (N_14245,N_7084,N_11675);
nand U14246 (N_14246,N_8909,N_6687);
xnor U14247 (N_14247,N_8165,N_8086);
xnor U14248 (N_14248,N_10749,N_10818);
and U14249 (N_14249,N_9976,N_9917);
xor U14250 (N_14250,N_7267,N_9172);
and U14251 (N_14251,N_10830,N_7892);
or U14252 (N_14252,N_10065,N_10748);
nand U14253 (N_14253,N_8480,N_11799);
nor U14254 (N_14254,N_7551,N_9517);
xnor U14255 (N_14255,N_8596,N_12171);
xor U14256 (N_14256,N_6733,N_9770);
nand U14257 (N_14257,N_11713,N_6775);
and U14258 (N_14258,N_11598,N_8185);
and U14259 (N_14259,N_7917,N_9606);
xor U14260 (N_14260,N_12441,N_8782);
nand U14261 (N_14261,N_6895,N_10586);
xor U14262 (N_14262,N_8015,N_9703);
nand U14263 (N_14263,N_7498,N_7265);
xor U14264 (N_14264,N_9528,N_10494);
nor U14265 (N_14265,N_11295,N_8454);
and U14266 (N_14266,N_9871,N_7794);
nor U14267 (N_14267,N_9943,N_11428);
nor U14268 (N_14268,N_6569,N_9673);
nor U14269 (N_14269,N_12118,N_12143);
nor U14270 (N_14270,N_11119,N_8366);
or U14271 (N_14271,N_8926,N_10837);
nand U14272 (N_14272,N_6644,N_6903);
or U14273 (N_14273,N_10487,N_7446);
nor U14274 (N_14274,N_6675,N_8311);
or U14275 (N_14275,N_9983,N_11890);
nand U14276 (N_14276,N_8814,N_12179);
and U14277 (N_14277,N_9318,N_10786);
nand U14278 (N_14278,N_10043,N_6336);
and U14279 (N_14279,N_11727,N_9432);
xor U14280 (N_14280,N_9344,N_6282);
or U14281 (N_14281,N_11398,N_9846);
nand U14282 (N_14282,N_8089,N_11843);
and U14283 (N_14283,N_8772,N_7116);
nand U14284 (N_14284,N_8613,N_6512);
xor U14285 (N_14285,N_6824,N_11171);
or U14286 (N_14286,N_11131,N_11393);
xor U14287 (N_14287,N_8927,N_11315);
or U14288 (N_14288,N_8443,N_11418);
and U14289 (N_14289,N_10025,N_8509);
and U14290 (N_14290,N_8506,N_11511);
or U14291 (N_14291,N_6332,N_9648);
or U14292 (N_14292,N_12241,N_6522);
nor U14293 (N_14293,N_6691,N_6415);
and U14294 (N_14294,N_10821,N_7207);
xnor U14295 (N_14295,N_9195,N_10965);
nor U14296 (N_14296,N_7101,N_11194);
nand U14297 (N_14297,N_9090,N_9961);
nor U14298 (N_14298,N_11941,N_9270);
or U14299 (N_14299,N_11462,N_12443);
xor U14300 (N_14300,N_6396,N_9338);
nand U14301 (N_14301,N_9039,N_7834);
or U14302 (N_14302,N_11031,N_6682);
xnor U14303 (N_14303,N_12153,N_8224);
nor U14304 (N_14304,N_10790,N_11582);
xor U14305 (N_14305,N_7249,N_11135);
nor U14306 (N_14306,N_12035,N_7487);
or U14307 (N_14307,N_9124,N_11076);
and U14308 (N_14308,N_8982,N_10947);
and U14309 (N_14309,N_7312,N_9496);
nor U14310 (N_14310,N_11508,N_9395);
or U14311 (N_14311,N_6667,N_11634);
nand U14312 (N_14312,N_8216,N_12157);
and U14313 (N_14313,N_6265,N_9944);
nor U14314 (N_14314,N_9165,N_7930);
nand U14315 (N_14315,N_8491,N_6350);
xor U14316 (N_14316,N_8335,N_8695);
nor U14317 (N_14317,N_11383,N_12149);
and U14318 (N_14318,N_11294,N_8471);
and U14319 (N_14319,N_8170,N_9314);
xor U14320 (N_14320,N_8027,N_11102);
nand U14321 (N_14321,N_10693,N_11354);
xor U14322 (N_14322,N_10472,N_8084);
or U14323 (N_14323,N_10529,N_9509);
and U14324 (N_14324,N_10287,N_11609);
xnor U14325 (N_14325,N_8373,N_10648);
and U14326 (N_14326,N_12119,N_11533);
and U14327 (N_14327,N_10162,N_6876);
xor U14328 (N_14328,N_7635,N_8240);
or U14329 (N_14329,N_7734,N_10626);
and U14330 (N_14330,N_6619,N_11388);
or U14331 (N_14331,N_6327,N_10757);
or U14332 (N_14332,N_7450,N_7233);
or U14333 (N_14333,N_10299,N_10742);
nand U14334 (N_14334,N_9767,N_11121);
nand U14335 (N_14335,N_6964,N_7409);
xor U14336 (N_14336,N_11661,N_6452);
xor U14337 (N_14337,N_11624,N_7390);
or U14338 (N_14338,N_12348,N_11196);
nor U14339 (N_14339,N_7603,N_10292);
xor U14340 (N_14340,N_8638,N_11478);
nor U14341 (N_14341,N_12463,N_12474);
xor U14342 (N_14342,N_8728,N_9133);
xor U14343 (N_14343,N_10060,N_9995);
nor U14344 (N_14344,N_8032,N_6546);
nor U14345 (N_14345,N_10889,N_9023);
and U14346 (N_14346,N_12093,N_11325);
nor U14347 (N_14347,N_8590,N_10282);
nor U14348 (N_14348,N_7378,N_7553);
or U14349 (N_14349,N_6684,N_11449);
xor U14350 (N_14350,N_7174,N_10780);
or U14351 (N_14351,N_7085,N_7787);
xor U14352 (N_14352,N_11283,N_9839);
nor U14353 (N_14353,N_10995,N_6844);
and U14354 (N_14354,N_8901,N_8996);
and U14355 (N_14355,N_8527,N_10036);
nor U14356 (N_14356,N_8126,N_7105);
and U14357 (N_14357,N_6273,N_7024);
nand U14358 (N_14358,N_11950,N_11652);
or U14359 (N_14359,N_9108,N_11904);
and U14360 (N_14360,N_11044,N_7475);
nand U14361 (N_14361,N_7339,N_10349);
nor U14362 (N_14362,N_7622,N_10193);
and U14363 (N_14363,N_11992,N_8905);
and U14364 (N_14364,N_11320,N_10460);
and U14365 (N_14365,N_8316,N_8152);
and U14366 (N_14366,N_10763,N_7700);
nand U14367 (N_14367,N_11772,N_9010);
or U14368 (N_14368,N_6606,N_9711);
xnor U14369 (N_14369,N_7898,N_12493);
nor U14370 (N_14370,N_8291,N_7662);
xor U14371 (N_14371,N_6794,N_8693);
nor U14372 (N_14372,N_11443,N_10681);
nor U14373 (N_14373,N_12490,N_9237);
nor U14374 (N_14374,N_8103,N_8838);
xor U14375 (N_14375,N_6879,N_8987);
and U14376 (N_14376,N_9078,N_11724);
nand U14377 (N_14377,N_9731,N_9865);
nor U14378 (N_14378,N_9275,N_10578);
or U14379 (N_14379,N_12060,N_10899);
nand U14380 (N_14380,N_9912,N_7759);
or U14381 (N_14381,N_11066,N_12014);
xor U14382 (N_14382,N_8818,N_8026);
or U14383 (N_14383,N_8166,N_8644);
nand U14384 (N_14384,N_10403,N_12175);
and U14385 (N_14385,N_8897,N_7664);
xnor U14386 (N_14386,N_10559,N_6312);
xnor U14387 (N_14387,N_10623,N_8712);
nand U14388 (N_14388,N_7765,N_9392);
and U14389 (N_14389,N_10445,N_10311);
nand U14390 (N_14390,N_9579,N_7861);
nor U14391 (N_14391,N_10263,N_8243);
nand U14392 (N_14392,N_9209,N_12382);
nand U14393 (N_14393,N_7066,N_9883);
and U14394 (N_14394,N_11268,N_7457);
and U14395 (N_14395,N_10022,N_7666);
xnor U14396 (N_14396,N_9091,N_6596);
nor U14397 (N_14397,N_12073,N_12380);
nand U14398 (N_14398,N_6850,N_7058);
and U14399 (N_14399,N_6810,N_9272);
nand U14400 (N_14400,N_10414,N_10937);
nand U14401 (N_14401,N_12470,N_7866);
xor U14402 (N_14402,N_9239,N_12389);
nor U14403 (N_14403,N_12057,N_11538);
and U14404 (N_14404,N_9623,N_6380);
or U14405 (N_14405,N_9136,N_9038);
or U14406 (N_14406,N_10772,N_6869);
nor U14407 (N_14407,N_6337,N_11528);
nand U14408 (N_14408,N_8207,N_9084);
nand U14409 (N_14409,N_10760,N_12423);
and U14410 (N_14410,N_6856,N_8607);
nor U14411 (N_14411,N_6913,N_12103);
nand U14412 (N_14412,N_7768,N_9746);
or U14413 (N_14413,N_12328,N_11587);
or U14414 (N_14414,N_11106,N_10943);
and U14415 (N_14415,N_8878,N_9797);
xor U14416 (N_14416,N_8135,N_11379);
nor U14417 (N_14417,N_11143,N_12050);
and U14418 (N_14418,N_10812,N_7492);
nand U14419 (N_14419,N_10443,N_10052);
nor U14420 (N_14420,N_8555,N_9827);
xor U14421 (N_14421,N_7933,N_9320);
and U14422 (N_14422,N_10974,N_11522);
or U14423 (N_14423,N_8099,N_11686);
nor U14424 (N_14424,N_6629,N_6306);
nand U14425 (N_14425,N_10517,N_7648);
xnor U14426 (N_14426,N_11039,N_11168);
xor U14427 (N_14427,N_7896,N_8284);
or U14428 (N_14428,N_6570,N_8476);
nand U14429 (N_14429,N_7774,N_8978);
or U14430 (N_14430,N_8334,N_9678);
xnor U14431 (N_14431,N_12203,N_7260);
or U14432 (N_14432,N_9413,N_9859);
nand U14433 (N_14433,N_11242,N_9776);
nor U14434 (N_14434,N_7829,N_8669);
or U14435 (N_14435,N_9818,N_6375);
nand U14436 (N_14436,N_10154,N_6807);
nor U14437 (N_14437,N_10730,N_7288);
nand U14438 (N_14438,N_9524,N_9549);
nor U14439 (N_14439,N_9066,N_11893);
xor U14440 (N_14440,N_10826,N_8715);
nand U14441 (N_14441,N_7221,N_8428);
or U14442 (N_14442,N_6479,N_12498);
or U14443 (N_14443,N_11632,N_10496);
and U14444 (N_14444,N_9644,N_9820);
and U14445 (N_14445,N_10265,N_11089);
and U14446 (N_14446,N_7701,N_9006);
nor U14447 (N_14447,N_6731,N_11666);
or U14448 (N_14448,N_7889,N_6834);
and U14449 (N_14449,N_12376,N_9847);
and U14450 (N_14450,N_10488,N_9778);
nand U14451 (N_14451,N_8178,N_8350);
nor U14452 (N_14452,N_12275,N_7459);
nand U14453 (N_14453,N_12406,N_11427);
nor U14454 (N_14454,N_6987,N_9753);
nor U14455 (N_14455,N_7762,N_7619);
nand U14456 (N_14456,N_10951,N_8736);
nand U14457 (N_14457,N_9459,N_10634);
or U14458 (N_14458,N_9998,N_8584);
and U14459 (N_14459,N_11124,N_9833);
or U14460 (N_14460,N_10759,N_7407);
xor U14461 (N_14461,N_8447,N_8566);
xnor U14462 (N_14462,N_11797,N_7668);
and U14463 (N_14463,N_11262,N_12240);
xor U14464 (N_14464,N_7500,N_12400);
nor U14465 (N_14465,N_10217,N_7855);
nand U14466 (N_14466,N_10392,N_8052);
and U14467 (N_14467,N_8672,N_10495);
or U14468 (N_14468,N_10841,N_6437);
nor U14469 (N_14469,N_9298,N_7599);
or U14470 (N_14470,N_11639,N_8237);
or U14471 (N_14471,N_12211,N_10452);
xor U14472 (N_14472,N_11347,N_6882);
nor U14473 (N_14473,N_10877,N_8741);
nor U14474 (N_14474,N_7981,N_11191);
or U14475 (N_14475,N_11825,N_8067);
xnor U14476 (N_14476,N_9927,N_10699);
and U14477 (N_14477,N_11760,N_8577);
and U14478 (N_14478,N_11736,N_9187);
nor U14479 (N_14479,N_9877,N_7783);
nor U14480 (N_14480,N_10264,N_7229);
nand U14481 (N_14481,N_7253,N_10186);
or U14482 (N_14482,N_7237,N_11776);
xor U14483 (N_14483,N_9219,N_8698);
xnor U14484 (N_14484,N_10601,N_9661);
nand U14485 (N_14485,N_9269,N_11990);
nand U14486 (N_14486,N_12264,N_11327);
xor U14487 (N_14487,N_9399,N_9971);
or U14488 (N_14488,N_7180,N_6829);
nand U14489 (N_14489,N_7386,N_11891);
xnor U14490 (N_14490,N_9287,N_9518);
nor U14491 (N_14491,N_8776,N_8710);
or U14492 (N_14492,N_9312,N_7887);
nor U14493 (N_14493,N_9975,N_10666);
nand U14494 (N_14494,N_11402,N_9807);
and U14495 (N_14495,N_7971,N_9863);
nand U14496 (N_14496,N_10457,N_12053);
nand U14497 (N_14497,N_11406,N_10791);
nor U14498 (N_14498,N_8561,N_8434);
and U14499 (N_14499,N_11796,N_9445);
or U14500 (N_14500,N_11534,N_8053);
or U14501 (N_14501,N_9805,N_12072);
xor U14502 (N_14502,N_8774,N_11785);
or U14503 (N_14503,N_12183,N_8098);
nand U14504 (N_14504,N_10507,N_10484);
xor U14505 (N_14505,N_8493,N_10319);
or U14506 (N_14506,N_8230,N_10844);
nand U14507 (N_14507,N_7401,N_10923);
nand U14508 (N_14508,N_12074,N_6602);
nor U14509 (N_14509,N_8921,N_9600);
and U14510 (N_14510,N_8313,N_8881);
nor U14511 (N_14511,N_7091,N_9695);
and U14512 (N_14512,N_9118,N_8302);
or U14513 (N_14513,N_10008,N_6343);
and U14514 (N_14514,N_6597,N_11861);
xnor U14515 (N_14515,N_7159,N_7810);
or U14516 (N_14516,N_7238,N_6285);
nand U14517 (N_14517,N_7555,N_9080);
and U14518 (N_14518,N_7346,N_9002);
nand U14519 (N_14519,N_11811,N_7218);
or U14520 (N_14520,N_6803,N_9686);
xor U14521 (N_14521,N_10622,N_6345);
and U14522 (N_14522,N_6790,N_10229);
and U14523 (N_14523,N_9122,N_12198);
nor U14524 (N_14524,N_10993,N_9639);
nand U14525 (N_14525,N_9694,N_8299);
and U14526 (N_14526,N_10295,N_8306);
nor U14527 (N_14527,N_7095,N_8761);
or U14528 (N_14528,N_10286,N_11786);
nand U14529 (N_14529,N_8679,N_12430);
xor U14530 (N_14530,N_10503,N_10004);
nor U14531 (N_14531,N_9407,N_10409);
nand U14532 (N_14532,N_11173,N_11597);
nor U14533 (N_14533,N_9985,N_10211);
xnor U14534 (N_14534,N_6699,N_9429);
nand U14535 (N_14535,N_11651,N_10221);
and U14536 (N_14536,N_8142,N_12112);
xnor U14537 (N_14537,N_10537,N_7589);
nand U14538 (N_14538,N_11045,N_6709);
xor U14539 (N_14539,N_9527,N_9420);
xnor U14540 (N_14540,N_10862,N_8357);
nor U14541 (N_14541,N_9611,N_6378);
nor U14542 (N_14542,N_9292,N_8337);
nand U14543 (N_14543,N_7521,N_6878);
nand U14544 (N_14544,N_10216,N_11363);
xor U14545 (N_14545,N_8792,N_11683);
or U14546 (N_14546,N_7414,N_8804);
or U14547 (N_14547,N_10325,N_8341);
or U14548 (N_14548,N_8431,N_8827);
nor U14549 (N_14549,N_6870,N_10097);
and U14550 (N_14550,N_6988,N_9186);
nor U14551 (N_14551,N_10485,N_10854);
or U14552 (N_14552,N_11414,N_11239);
xnor U14553 (N_14553,N_10697,N_7355);
xnor U14554 (N_14554,N_9962,N_8095);
xor U14555 (N_14555,N_8771,N_11144);
nand U14556 (N_14556,N_6984,N_7900);
or U14557 (N_14557,N_10532,N_10509);
or U14558 (N_14558,N_8221,N_7019);
nor U14559 (N_14559,N_11915,N_11360);
and U14560 (N_14560,N_11470,N_6417);
and U14561 (N_14561,N_6516,N_7582);
xor U14562 (N_14562,N_11953,N_6884);
and U14563 (N_14563,N_6463,N_7796);
nor U14564 (N_14564,N_8500,N_10832);
xnor U14565 (N_14565,N_11251,N_11611);
xnor U14566 (N_14566,N_9941,N_9621);
nor U14567 (N_14567,N_11164,N_10525);
nor U14568 (N_14568,N_7529,N_6864);
nor U14569 (N_14569,N_6919,N_10589);
xor U14570 (N_14570,N_6764,N_11454);
or U14571 (N_14571,N_11584,N_11099);
nor U14572 (N_14572,N_7805,N_11483);
nor U14573 (N_14573,N_7222,N_9970);
xor U14574 (N_14574,N_9197,N_11290);
xor U14575 (N_14575,N_8622,N_6659);
nand U14576 (N_14576,N_11016,N_8852);
nor U14577 (N_14577,N_10483,N_11166);
xor U14578 (N_14578,N_8225,N_8920);
or U14579 (N_14579,N_6275,N_9458);
nor U14580 (N_14580,N_12009,N_10777);
nor U14581 (N_14581,N_9936,N_10806);
nand U14582 (N_14582,N_10347,N_8309);
or U14583 (N_14583,N_7577,N_8542);
nor U14584 (N_14584,N_8733,N_9745);
nor U14585 (N_14585,N_6499,N_9852);
nor U14586 (N_14586,N_11937,N_9101);
xnor U14587 (N_14587,N_8351,N_7276);
nand U14588 (N_14588,N_7847,N_12111);
and U14589 (N_14589,N_9131,N_8263);
nor U14590 (N_14590,N_10468,N_6573);
xnor U14591 (N_14591,N_6941,N_7305);
nand U14592 (N_14592,N_7588,N_8384);
xor U14593 (N_14593,N_12330,N_9450);
nor U14594 (N_14594,N_8994,N_10155);
or U14595 (N_14595,N_6478,N_10708);
nor U14596 (N_14596,N_12298,N_8999);
and U14597 (N_14597,N_10126,N_9690);
or U14598 (N_14598,N_7406,N_9755);
nor U14599 (N_14599,N_11889,N_12377);
and U14600 (N_14600,N_12417,N_6627);
and U14601 (N_14601,N_11475,N_10305);
xnor U14602 (N_14602,N_6290,N_10596);
or U14603 (N_14603,N_11658,N_10353);
nand U14604 (N_14604,N_8176,N_11254);
nand U14605 (N_14605,N_7772,N_11627);
or U14606 (N_14606,N_10541,N_11878);
and U14607 (N_14607,N_9201,N_6532);
nand U14608 (N_14608,N_6798,N_10915);
nand U14609 (N_14609,N_10776,N_11074);
xor U14610 (N_14610,N_10169,N_9635);
xnor U14611 (N_14611,N_11339,N_11965);
nand U14612 (N_14612,N_9264,N_7093);
and U14613 (N_14613,N_9634,N_12172);
nand U14614 (N_14614,N_7680,N_9913);
or U14615 (N_14615,N_6297,N_9596);
nor U14616 (N_14616,N_11923,N_10792);
and U14617 (N_14617,N_6371,N_10897);
nor U14618 (N_14618,N_10049,N_6652);
and U14619 (N_14619,N_8666,N_8798);
or U14620 (N_14620,N_8791,N_11204);
nand U14621 (N_14621,N_7484,N_11022);
xnor U14622 (N_14622,N_11671,N_11275);
and U14623 (N_14623,N_10370,N_6966);
or U14624 (N_14624,N_12080,N_10259);
nor U14625 (N_14625,N_8376,N_9642);
nand U14626 (N_14626,N_10153,N_7910);
and U14627 (N_14627,N_10651,N_10991);
xor U14628 (N_14628,N_12327,N_7035);
and U14629 (N_14629,N_9307,N_8260);
xnor U14630 (N_14630,N_11716,N_7348);
and U14631 (N_14631,N_6710,N_7694);
nand U14632 (N_14632,N_8945,N_8010);
and U14633 (N_14633,N_11403,N_12056);
and U14634 (N_14634,N_9184,N_10434);
xnor U14635 (N_14635,N_10064,N_10131);
xor U14636 (N_14636,N_7486,N_7817);
or U14637 (N_14637,N_7036,N_6943);
nor U14638 (N_14638,N_10500,N_6957);
and U14639 (N_14639,N_8492,N_9607);
nand U14640 (N_14640,N_10384,N_6531);
nand U14641 (N_14641,N_9364,N_8743);
and U14642 (N_14642,N_11480,N_12270);
nand U14643 (N_14643,N_6999,N_6975);
xnor U14644 (N_14644,N_11085,N_6365);
and U14645 (N_14645,N_9942,N_9614);
nand U14646 (N_14646,N_7121,N_6329);
or U14647 (N_14647,N_9401,N_12365);
and U14648 (N_14648,N_11974,N_11082);
nand U14649 (N_14649,N_11118,N_6491);
and U14650 (N_14650,N_9075,N_9036);
or U14651 (N_14651,N_8106,N_7335);
nor U14652 (N_14652,N_12213,N_9235);
and U14653 (N_14653,N_8078,N_10085);
nor U14654 (N_14654,N_10804,N_6962);
nand U14655 (N_14655,N_9126,N_6933);
or U14656 (N_14656,N_11806,N_11747);
or U14657 (N_14657,N_11509,N_6698);
nor U14658 (N_14658,N_10394,N_12087);
xor U14659 (N_14659,N_10062,N_10949);
nand U14660 (N_14660,N_9360,N_10667);
xor U14661 (N_14661,N_7950,N_6735);
nor U14662 (N_14662,N_10713,N_10904);
nand U14663 (N_14663,N_10288,N_10501);
or U14664 (N_14664,N_7831,N_6641);
xnor U14665 (N_14665,N_6376,N_10293);
or U14666 (N_14666,N_10774,N_10922);
and U14667 (N_14667,N_11945,N_7302);
and U14668 (N_14668,N_12343,N_8727);
and U14669 (N_14669,N_8597,N_12341);
nand U14670 (N_14670,N_10401,N_6836);
nand U14671 (N_14671,N_7137,N_7628);
nand U14672 (N_14672,N_7542,N_8031);
or U14673 (N_14673,N_8051,N_11053);
and U14674 (N_14674,N_11792,N_11284);
nor U14675 (N_14675,N_10984,N_9828);
nor U14676 (N_14676,N_10724,N_7271);
nor U14677 (N_14677,N_10871,N_6467);
nand U14678 (N_14678,N_9558,N_10076);
xor U14679 (N_14679,N_11743,N_11944);
or U14680 (N_14680,N_8763,N_10614);
or U14681 (N_14681,N_12351,N_10184);
and U14682 (N_14682,N_9125,N_11150);
nand U14683 (N_14683,N_9765,N_9106);
nor U14684 (N_14684,N_9721,N_11549);
or U14685 (N_14685,N_11112,N_12371);
or U14686 (N_14686,N_8685,N_8756);
nand U14687 (N_14687,N_8046,N_11955);
or U14688 (N_14688,N_11156,N_8327);
xnor U14689 (N_14689,N_6926,N_8392);
nor U14690 (N_14690,N_10144,N_10002);
xor U14691 (N_14691,N_10687,N_9061);
nand U14692 (N_14692,N_9729,N_10274);
xor U14693 (N_14693,N_10332,N_10689);
and U14694 (N_14694,N_11778,N_6299);
nand U14695 (N_14695,N_6384,N_12255);
nor U14696 (N_14696,N_6920,N_9426);
and U14697 (N_14697,N_6714,N_9333);
and U14698 (N_14698,N_8912,N_8802);
xor U14699 (N_14699,N_9730,N_9311);
or U14700 (N_14700,N_8361,N_9934);
nand U14701 (N_14701,N_12081,N_8317);
xor U14702 (N_14702,N_8286,N_9213);
or U14703 (N_14703,N_7506,N_7615);
nor U14704 (N_14704,N_9138,N_11567);
nor U14705 (N_14705,N_9554,N_8830);
xnor U14706 (N_14706,N_10600,N_12296);
nand U14707 (N_14707,N_11137,N_7516);
nor U14708 (N_14708,N_8068,N_8797);
or U14709 (N_14709,N_8389,N_9477);
or U14710 (N_14710,N_10702,N_6832);
or U14711 (N_14711,N_9740,N_6535);
xnor U14712 (N_14712,N_6734,N_10296);
or U14713 (N_14713,N_8593,N_9281);
nand U14714 (N_14714,N_10188,N_9886);
or U14715 (N_14715,N_10847,N_6321);
or U14716 (N_14716,N_7331,N_8643);
nand U14717 (N_14717,N_8300,N_10510);
xnor U14718 (N_14718,N_10709,N_6932);
nand U14719 (N_14719,N_7245,N_8094);
xor U14720 (N_14720,N_9332,N_7442);
nor U14721 (N_14721,N_8983,N_8821);
xor U14722 (N_14722,N_9284,N_11929);
nand U14723 (N_14723,N_9560,N_12155);
nor U14724 (N_14724,N_8268,N_12426);
or U14725 (N_14725,N_9215,N_8929);
nand U14726 (N_14726,N_7044,N_11264);
xnor U14727 (N_14727,N_8321,N_9759);
nor U14728 (N_14728,N_9355,N_10939);
and U14729 (N_14729,N_11001,N_7389);
or U14730 (N_14730,N_7482,N_8993);
and U14731 (N_14731,N_11637,N_8580);
xor U14732 (N_14732,N_10734,N_9207);
nor U14733 (N_14733,N_8759,N_11780);
nor U14734 (N_14734,N_7883,N_10479);
xor U14735 (N_14735,N_10073,N_9435);
nand U14736 (N_14736,N_10739,N_8348);
xnor U14737 (N_14737,N_11600,N_9497);
nand U14738 (N_14738,N_11065,N_9796);
nor U14739 (N_14739,N_12007,N_9698);
or U14740 (N_14740,N_10304,N_7124);
and U14741 (N_14741,N_11912,N_9823);
and U14742 (N_14742,N_7143,N_7677);
nor U14743 (N_14743,N_11723,N_8075);
and U14744 (N_14744,N_9301,N_11220);
xor U14745 (N_14745,N_12170,N_9222);
or U14746 (N_14746,N_9523,N_12332);
or U14747 (N_14747,N_9801,N_11034);
xor U14748 (N_14748,N_7078,N_12124);
nand U14749 (N_14749,N_6283,N_12011);
xor U14750 (N_14750,N_10556,N_6511);
and U14751 (N_14751,N_7059,N_11129);
xnor U14752 (N_14752,N_9334,N_11774);
or U14753 (N_14753,N_7728,N_8034);
nand U14754 (N_14754,N_7602,N_11678);
and U14755 (N_14755,N_9826,N_8730);
and U14756 (N_14756,N_8832,N_9585);
xnor U14757 (N_14757,N_8709,N_7491);
or U14758 (N_14758,N_6625,N_11933);
xor U14759 (N_14759,N_6355,N_11056);
and U14760 (N_14760,N_10552,N_7658);
and U14761 (N_14761,N_8657,N_6353);
nand U14762 (N_14762,N_10035,N_8422);
xor U14763 (N_14763,N_11728,N_7255);
nand U14764 (N_14764,N_8295,N_7007);
or U14765 (N_14765,N_8757,N_7257);
xnor U14766 (N_14766,N_6555,N_7344);
nor U14767 (N_14767,N_11507,N_12482);
and U14768 (N_14768,N_8739,N_11517);
or U14769 (N_14769,N_6927,N_7689);
nor U14770 (N_14770,N_7471,N_8120);
nand U14771 (N_14771,N_11659,N_12178);
and U14772 (N_14772,N_7236,N_10262);
or U14773 (N_14773,N_11276,N_10089);
nand U14774 (N_14774,N_10453,N_8522);
xor U14775 (N_14775,N_7663,N_8399);
nand U14776 (N_14776,N_7618,N_8860);
nor U14777 (N_14777,N_8293,N_8330);
nor U14778 (N_14778,N_7186,N_10315);
xor U14779 (N_14779,N_8036,N_7258);
or U14780 (N_14780,N_11024,N_9537);
nand U14781 (N_14781,N_8908,N_8117);
xor U14782 (N_14782,N_9593,N_9725);
nand U14783 (N_14783,N_8439,N_10381);
and U14784 (N_14784,N_8005,N_7043);
nor U14785 (N_14785,N_7873,N_10192);
or U14786 (N_14786,N_8902,N_10412);
and U14787 (N_14787,N_12086,N_11803);
nand U14788 (N_14788,N_7891,N_10147);
and U14789 (N_14789,N_6583,N_10924);
and U14790 (N_14790,N_7011,N_12467);
nor U14791 (N_14791,N_10309,N_6745);
xnor U14792 (N_14792,N_10356,N_11677);
nand U14793 (N_14793,N_11433,N_9972);
nor U14794 (N_14794,N_11160,N_8975);
nor U14795 (N_14795,N_7751,N_7856);
and U14796 (N_14796,N_6524,N_6441);
nor U14797 (N_14797,N_9013,N_11097);
and U14798 (N_14798,N_6459,N_8289);
nor U14799 (N_14799,N_11649,N_7857);
and U14800 (N_14800,N_7986,N_9408);
nand U14801 (N_14801,N_8667,N_8066);
nand U14802 (N_14802,N_10013,N_10828);
xor U14803 (N_14803,N_8579,N_7147);
xnor U14804 (N_14804,N_7736,N_12078);
nand U14805 (N_14805,N_7330,N_10387);
or U14806 (N_14806,N_10936,N_6495);
xor U14807 (N_14807,N_12196,N_6666);
nor U14808 (N_14808,N_7380,N_8610);
nor U14809 (N_14809,N_10134,N_9166);
and U14810 (N_14810,N_11188,N_9716);
and U14811 (N_14811,N_12402,N_9015);
xor U14812 (N_14812,N_8591,N_7086);
nor U14813 (N_14813,N_10351,N_12079);
nor U14814 (N_14814,N_7709,N_10116);
nor U14815 (N_14815,N_9164,N_11364);
nand U14816 (N_14816,N_11527,N_6311);
nor U14817 (N_14817,N_12265,N_7279);
and U14818 (N_14818,N_8136,N_10223);
nand U14819 (N_14819,N_12280,N_12355);
xnor U14820 (N_14820,N_8105,N_10082);
nor U14821 (N_14821,N_7702,N_10911);
nor U14822 (N_14822,N_9437,N_7539);
nor U14823 (N_14823,N_8272,N_12420);
and U14824 (N_14824,N_7321,N_12030);
and U14825 (N_14825,N_6576,N_7528);
nand U14826 (N_14826,N_11579,N_6780);
nand U14827 (N_14827,N_7424,N_6612);
xnor U14828 (N_14828,N_12284,N_9330);
nand U14829 (N_14829,N_6849,N_11775);
xnor U14830 (N_14830,N_10819,N_11704);
nor U14831 (N_14831,N_11373,N_8836);
nand U14832 (N_14832,N_12046,N_7187);
nand U14833 (N_14833,N_11750,N_11357);
xnor U14834 (N_14834,N_6793,N_11265);
xnor U14835 (N_14835,N_6816,N_7732);
nor U14836 (N_14836,N_11558,N_8177);
xnor U14837 (N_14837,N_6762,N_8904);
nand U14838 (N_14838,N_9294,N_6873);
and U14839 (N_14839,N_7359,N_11401);
or U14840 (N_14840,N_8914,N_10009);
xor U14841 (N_14841,N_12494,N_11892);
or U14842 (N_14842,N_8990,N_12045);
nand U14843 (N_14843,N_9525,N_7200);
or U14844 (N_14844,N_7799,N_11457);
nand U14845 (N_14845,N_11930,N_9297);
xnor U14846 (N_14846,N_8578,N_8559);
or U14847 (N_14847,N_11607,N_11960);
nand U14848 (N_14848,N_10736,N_11415);
xnor U14849 (N_14849,N_7154,N_10152);
and U14850 (N_14850,N_11979,N_9573);
nand U14851 (N_14851,N_10765,N_9681);
or U14852 (N_14852,N_6976,N_8383);
and U14853 (N_14853,N_9939,N_6930);
nor U14854 (N_14854,N_7773,N_10636);
or U14855 (N_14855,N_7138,N_7868);
xnor U14856 (N_14856,N_7270,N_7541);
and U14857 (N_14857,N_10271,N_6444);
nor U14858 (N_14858,N_12101,N_8275);
or U14859 (N_14859,N_11988,N_11484);
xnor U14860 (N_14860,N_7595,N_10896);
nor U14861 (N_14861,N_11888,N_9858);
nand U14862 (N_14862,N_6537,N_11042);
nor U14863 (N_14863,N_7223,N_6582);
nor U14864 (N_14864,N_11557,N_10876);
and U14865 (N_14865,N_10789,N_10665);
nand U14866 (N_14866,N_7261,N_11244);
and U14867 (N_14867,N_8223,N_7825);
or U14868 (N_14868,N_7511,N_11815);
xnor U14869 (N_14869,N_12454,N_10775);
nand U14870 (N_14870,N_7327,N_9267);
or U14871 (N_14871,N_10964,N_12158);
or U14872 (N_14872,N_10583,N_6938);
xnor U14873 (N_14873,N_7168,N_8140);
and U14874 (N_14874,N_11910,N_8342);
xor U14875 (N_14875,N_11993,N_11753);
nor U14876 (N_14876,N_6372,N_11371);
nor U14877 (N_14877,N_9535,N_6288);
xor U14878 (N_14878,N_11179,N_9358);
xor U14879 (N_14879,N_6432,N_6393);
nand U14880 (N_14880,N_8134,N_8482);
and U14881 (N_14881,N_9029,N_6442);
nand U14882 (N_14882,N_11696,N_10011);
or U14883 (N_14883,N_12260,N_9815);
nand U14884 (N_14884,N_10018,N_10941);
nand U14885 (N_14885,N_6925,N_11003);
xor U14886 (N_14886,N_12448,N_6787);
and U14887 (N_14887,N_9633,N_7708);
or U14888 (N_14888,N_6695,N_10577);
nor U14889 (N_14889,N_10212,N_7936);
or U14890 (N_14890,N_10439,N_11425);
nand U14891 (N_14891,N_6581,N_8242);
and U14892 (N_14892,N_8783,N_8162);
xor U14893 (N_14893,N_6685,N_11331);
nand U14894 (N_14894,N_8190,N_8382);
nand U14895 (N_14895,N_6360,N_8639);
nand U14896 (N_14896,N_11939,N_7607);
and U14897 (N_14897,N_6266,N_7509);
or U14898 (N_14898,N_7133,N_7001);
nand U14899 (N_14899,N_10051,N_8675);
nand U14900 (N_14900,N_8807,N_12421);
or U14901 (N_14901,N_6693,N_9087);
nand U14902 (N_14902,N_8549,N_6599);
and U14903 (N_14903,N_7162,N_6662);
and U14904 (N_14904,N_9411,N_9151);
nor U14905 (N_14905,N_8726,N_12044);
nand U14906 (N_14906,N_7594,N_6502);
nor U14907 (N_14907,N_10840,N_12210);
and U14908 (N_14908,N_10161,N_10337);
or U14909 (N_14909,N_8799,N_6963);
xnor U14910 (N_14910,N_8629,N_11769);
nor U14911 (N_14911,N_7991,N_6939);
and U14912 (N_14912,N_11874,N_7612);
or U14913 (N_14913,N_7351,N_8014);
xnor U14914 (N_14914,N_11017,N_9238);
nand U14915 (N_14915,N_10740,N_7469);
and U14916 (N_14916,N_9049,N_11744);
nand U14917 (N_14917,N_9763,N_10960);
nand U14918 (N_14918,N_7654,N_8450);
and U14919 (N_14919,N_11702,N_9938);
and U14920 (N_14920,N_7449,N_10396);
nand U14921 (N_14921,N_9169,N_7016);
nand U14922 (N_14922,N_7300,N_10754);
nor U14923 (N_14923,N_12015,N_12104);
xor U14924 (N_14924,N_12177,N_11763);
nor U14925 (N_14925,N_12135,N_9660);
nor U14926 (N_14926,N_7920,N_7111);
or U14927 (N_14927,N_9647,N_10954);
and U14928 (N_14928,N_10813,N_11041);
and U14929 (N_14929,N_9004,N_8572);
xor U14930 (N_14930,N_10048,N_7479);
nand U14931 (N_14931,N_12261,N_7193);
xor U14932 (N_14932,N_9866,N_9012);
and U14933 (N_14933,N_7869,N_9050);
nor U14934 (N_14934,N_11526,N_11002);
and U14935 (N_14935,N_8517,N_7561);
nand U14936 (N_14936,N_7793,N_10727);
nor U14937 (N_14937,N_8391,N_9100);
nand U14938 (N_14938,N_9468,N_8581);
nand U14939 (N_14939,N_12346,N_7443);
nand U14940 (N_14940,N_11260,N_7925);
xnor U14941 (N_14941,N_11198,N_6542);
and U14942 (N_14942,N_10103,N_6996);
or U14943 (N_14943,N_11770,N_9618);
and U14944 (N_14944,N_6342,N_12102);
nor U14945 (N_14945,N_10989,N_8261);
nand U14946 (N_14946,N_8038,N_7850);
or U14947 (N_14947,N_7188,N_8724);
and U14948 (N_14948,N_8432,N_7672);
xor U14949 (N_14949,N_9551,N_9158);
and U14950 (N_14950,N_10243,N_11594);
xnor U14951 (N_14951,N_7742,N_11140);
nand U14952 (N_14952,N_9520,N_9780);
or U14953 (N_14953,N_6911,N_11155);
and U14954 (N_14954,N_9464,N_11717);
and U14955 (N_14955,N_12248,N_10206);
nor U14956 (N_14956,N_10246,N_7325);
nor U14957 (N_14957,N_11343,N_6961);
xor U14958 (N_14958,N_11026,N_7807);
xor U14959 (N_14959,N_9790,N_9322);
xor U14960 (N_14960,N_11561,N_11098);
xnor U14961 (N_14961,N_11021,N_10591);
xnor U14962 (N_14962,N_6907,N_10168);
xor U14963 (N_14963,N_8312,N_10632);
nand U14964 (N_14964,N_9708,N_6455);
and U14965 (N_14965,N_9702,N_6826);
nor U14966 (N_14966,N_9657,N_9339);
xnor U14967 (N_14967,N_9819,N_8301);
and U14968 (N_14968,N_12032,N_12485);
nor U14969 (N_14969,N_7912,N_11752);
nand U14970 (N_14970,N_6383,N_7017);
nor U14971 (N_14971,N_9025,N_9575);
nor U14972 (N_14972,N_8055,N_8779);
and U14973 (N_14973,N_7737,N_6252);
nor U14974 (N_14974,N_11043,N_12040);
nor U14975 (N_14975,N_11348,N_11668);
or U14976 (N_14976,N_7808,N_9185);
and U14977 (N_14977,N_10024,N_6655);
nor U14978 (N_14978,N_6497,N_7865);
nor U14979 (N_14979,N_8976,N_11369);
nor U14980 (N_14980,N_8558,N_11943);
and U14981 (N_14981,N_9221,N_6605);
nor U14982 (N_14982,N_7391,N_8388);
nor U14983 (N_14983,N_8662,N_7303);
xnor U14984 (N_14984,N_7379,N_12152);
or U14985 (N_14985,N_7425,N_11574);
nand U14986 (N_14986,N_8813,N_8435);
nor U14987 (N_14987,N_11720,N_8258);
xnor U14988 (N_14988,N_7726,N_7753);
or U14989 (N_14989,N_11984,N_11292);
or U14990 (N_14990,N_6482,N_11879);
and U14991 (N_14991,N_6394,N_11838);
nand U14992 (N_14992,N_7034,N_11693);
nand U14993 (N_14993,N_10839,N_8463);
xor U14994 (N_14994,N_7360,N_8933);
nand U14995 (N_14995,N_12216,N_9831);
or U14996 (N_14996,N_8866,N_8077);
xor U14997 (N_14997,N_7206,N_11100);
nand U14998 (N_14998,N_9578,N_7720);
nor U14999 (N_14999,N_7504,N_11175);
and U15000 (N_15000,N_11572,N_8963);
nor U15001 (N_15001,N_9613,N_11823);
and U15002 (N_15002,N_7440,N_11187);
xnor U15003 (N_15003,N_12345,N_12272);
nor U15004 (N_15004,N_11236,N_10551);
xnor U15005 (N_15005,N_7118,N_8742);
or U15006 (N_15006,N_7212,N_10310);
nor U15007 (N_15007,N_12375,N_8689);
or U15008 (N_15008,N_12459,N_8307);
xor U15009 (N_15009,N_9313,N_8810);
and U15010 (N_15010,N_9277,N_6540);
xor U15011 (N_15011,N_8611,N_8485);
xnor U15012 (N_15012,N_11902,N_10655);
nand U15013 (N_15013,N_10620,N_12287);
nor U15014 (N_15014,N_12052,N_11130);
nand U15015 (N_15015,N_8349,N_12186);
nand U15016 (N_15016,N_7166,N_6529);
or U15017 (N_15017,N_10165,N_11335);
nand U15018 (N_15018,N_7228,N_9463);
xor U15019 (N_15019,N_9543,N_7656);
xor U15020 (N_15020,N_12465,N_9074);
nor U15021 (N_15021,N_7454,N_8236);
xnor U15022 (N_15022,N_7867,N_10903);
xnor U15023 (N_15023,N_10106,N_9963);
nand U15024 (N_15024,N_10493,N_7740);
and U15025 (N_15025,N_9493,N_7477);
or U15026 (N_15026,N_12379,N_8960);
xor U15027 (N_15027,N_6466,N_11655);
nand U15028 (N_15028,N_10203,N_11437);
or U15029 (N_15029,N_7365,N_6651);
xor U15030 (N_15030,N_10607,N_7250);
nor U15031 (N_15031,N_9206,N_8863);
nor U15032 (N_15032,N_8113,N_12252);
nor U15033 (N_15033,N_6584,N_7527);
xor U15034 (N_15034,N_7410,N_10955);
and U15035 (N_15035,N_8691,N_8101);
and U15036 (N_15036,N_8155,N_11547);
nand U15037 (N_15037,N_8585,N_6765);
xnor U15038 (N_15038,N_7292,N_12130);
nor U15039 (N_15039,N_6411,N_10793);
nor U15040 (N_15040,N_11208,N_7278);
or U15041 (N_15041,N_12357,N_6434);
nor U15042 (N_15042,N_6272,N_8028);
xnor U15043 (N_15043,N_10150,N_7611);
nor U15044 (N_15044,N_7057,N_10279);
and U15045 (N_15045,N_7038,N_10505);
nor U15046 (N_15046,N_12462,N_8775);
xnor U15047 (N_15047,N_10302,N_7266);
or U15048 (N_15048,N_11633,N_11023);
or U15049 (N_15049,N_11073,N_9317);
nor U15050 (N_15050,N_9992,N_8722);
and U15051 (N_15051,N_8182,N_8139);
nand U15052 (N_15052,N_11487,N_9541);
xnor U15053 (N_15053,N_7430,N_7585);
xor U15054 (N_15054,N_8871,N_8121);
or U15055 (N_15055,N_12344,N_10268);
nand U15056 (N_15056,N_7573,N_11667);
and U15057 (N_15057,N_10810,N_6750);
nor U15058 (N_15058,N_7995,N_6505);
or U15059 (N_15059,N_8255,N_12410);
nor U15060 (N_15060,N_9631,N_6701);
xor U15061 (N_15061,N_6281,N_12369);
or U15062 (N_15062,N_7894,N_8371);
and U15063 (N_15063,N_12230,N_6822);
and U15064 (N_15064,N_10975,N_6590);
nand U15065 (N_15065,N_9268,N_6863);
and U15066 (N_15066,N_10569,N_6910);
or U15067 (N_15067,N_9984,N_6658);
xnor U15068 (N_15068,N_9784,N_9965);
or U15069 (N_15069,N_10560,N_9850);
nand U15070 (N_15070,N_6638,N_8729);
and U15071 (N_15071,N_10100,N_7966);
nand U15072 (N_15072,N_7781,N_8731);
nand U15073 (N_15073,N_9026,N_8092);
or U15074 (N_15074,N_11257,N_11641);
and U15075 (N_15075,N_9856,N_10137);
xnor U15076 (N_15076,N_9350,N_10728);
xor U15077 (N_15077,N_11094,N_9190);
and U15078 (N_15078,N_7827,N_12161);
nand U15079 (N_15079,N_8196,N_11134);
nor U15080 (N_15080,N_10733,N_12163);
and U15081 (N_15081,N_8211,N_7481);
and U15082 (N_15082,N_8538,N_11367);
nor U15083 (N_15083,N_12068,N_7405);
or U15084 (N_15084,N_6909,N_10095);
nand U15085 (N_15085,N_12393,N_6994);
and U15086 (N_15086,N_8043,N_11853);
nand U15087 (N_15087,N_11765,N_7008);
nand U15088 (N_15088,N_9163,N_9265);
and U15089 (N_15089,N_9834,N_7536);
and U15090 (N_15090,N_6859,N_10625);
or U15091 (N_15091,N_7185,N_6851);
nor U15092 (N_15092,N_10015,N_6741);
nor U15093 (N_15093,N_9340,N_12475);
nor U15094 (N_15094,N_9704,N_8882);
nor U15095 (N_15095,N_7690,N_7361);
nor U15096 (N_15096,N_11059,N_10550);
and U15097 (N_15097,N_10416,N_12303);
or U15098 (N_15098,N_7946,N_7413);
nor U15099 (N_15099,N_8400,N_10746);
and U15100 (N_15100,N_10706,N_8489);
or U15101 (N_15101,N_7411,N_8414);
and U15102 (N_15102,N_11101,N_7812);
and U15103 (N_15103,N_8796,N_8065);
or U15104 (N_15104,N_10142,N_9882);
xnor U15105 (N_15105,N_10250,N_10567);
and U15106 (N_15106,N_11842,N_9867);
xnor U15107 (N_15107,N_8626,N_11411);
and U15108 (N_15108,N_8129,N_8037);
or U15109 (N_15109,N_9870,N_9997);
nand U15110 (N_15110,N_8888,N_7104);
or U15111 (N_15111,N_11860,N_7496);
nand U15112 (N_15112,N_11833,N_7870);
nor U15113 (N_15113,N_10322,N_11394);
nor U15114 (N_15114,N_11058,N_7755);
and U15115 (N_15115,N_8141,N_8917);
and U15116 (N_15116,N_8511,N_7710);
xor U15117 (N_15117,N_9836,N_6970);
xor U15118 (N_15118,N_7803,N_12429);
and U15119 (N_15119,N_10917,N_6890);
xor U15120 (N_15120,N_9035,N_7580);
xor U15121 (N_15121,N_10836,N_9067);
xor U15122 (N_15122,N_10297,N_9361);
or U15123 (N_15123,N_11863,N_7254);
nor U15124 (N_15124,N_9198,N_12208);
or U15125 (N_15125,N_8347,N_8907);
or U15126 (N_15126,N_7945,N_8532);
and U15127 (N_15127,N_11518,N_6860);
and U15128 (N_15128,N_11410,N_11793);
nand U15129 (N_15129,N_8998,N_7328);
xnor U15130 (N_15130,N_10884,N_6530);
nor U15131 (N_15131,N_9027,N_7201);
xor U15132 (N_15132,N_9610,N_8355);
nor U15133 (N_15133,N_6955,N_10807);
xor U15134 (N_15134,N_7421,N_10593);
nand U15135 (N_15135,N_8100,N_11712);
nor U15136 (N_15136,N_9670,N_8660);
nor U15137 (N_15137,N_6888,N_11695);
and U15138 (N_15138,N_10333,N_7148);
or U15139 (N_15139,N_9996,N_9231);
nor U15140 (N_15140,N_9423,N_12262);
xnor U15141 (N_15141,N_9652,N_8600);
or U15142 (N_15142,N_11555,N_8984);
nand U15143 (N_15143,N_9434,N_7934);
nand U15144 (N_15144,N_11189,N_6256);
and U15145 (N_15145,N_8468,N_10981);
nor U15146 (N_15146,N_11559,N_7416);
or U15147 (N_15147,N_10234,N_8641);
nor U15148 (N_15148,N_8680,N_7473);
xor U15149 (N_15149,N_6488,N_11715);
xor U15150 (N_15150,N_6563,N_8112);
nor U15151 (N_15151,N_8229,N_12222);
and U15152 (N_15152,N_11932,N_10010);
nor U15153 (N_15153,N_7211,N_9714);
or U15154 (N_15154,N_10676,N_6494);
and U15155 (N_15155,N_9017,N_7636);
and U15156 (N_15156,N_9412,N_8374);
or U15157 (N_15157,N_6786,N_10438);
xnor U15158 (N_15158,N_9768,N_7927);
nor U15159 (N_15159,N_11592,N_11434);
xor U15160 (N_15160,N_10834,N_8338);
xor U15161 (N_15161,N_8767,N_7466);
or U15162 (N_15162,N_8409,N_11319);
or U15163 (N_15163,N_7125,N_9051);
xnor U15164 (N_15164,N_11699,N_7376);
nand U15165 (N_15165,N_12326,N_12125);
nor U15166 (N_15166,N_9409,N_11424);
nor U15167 (N_15167,N_8407,N_7463);
and U15168 (N_15168,N_10761,N_9545);
and U15169 (N_15169,N_10753,N_11161);
and U15170 (N_15170,N_10408,N_9266);
nand U15171 (N_15171,N_6634,N_7828);
nor U15172 (N_15172,N_10992,N_10719);
nor U15173 (N_15173,N_9293,N_7661);
and U15174 (N_15174,N_8719,N_12221);
nor U15175 (N_15175,N_12117,N_7550);
xnor U15176 (N_15176,N_6703,N_8245);
xnor U15177 (N_15177,N_9159,N_9208);
and U15178 (N_15178,N_11304,N_7219);
and U15179 (N_15179,N_8525,N_8604);
and U15180 (N_15180,N_10210,N_6454);
nand U15181 (N_15181,N_11207,N_9144);
xor U15182 (N_15182,N_10863,N_11564);
and U15183 (N_15183,N_12338,N_7634);
nand U15184 (N_15184,N_7832,N_11942);
nand U15185 (N_15185,N_11232,N_9182);
nor U15186 (N_15186,N_7579,N_8303);
xnor U15187 (N_15187,N_9601,N_7286);
and U15188 (N_15188,N_9756,N_9196);
nand U15189 (N_15189,N_10205,N_12497);
xor U15190 (N_15190,N_8029,N_11148);
nand U15191 (N_15191,N_6989,N_11820);
nor U15192 (N_15192,N_8564,N_7129);
and U15193 (N_15193,N_6307,N_10258);
nand U15194 (N_15194,N_12414,N_10045);
and U15195 (N_15195,N_8154,N_7248);
and U15196 (N_15196,N_8850,N_12403);
nand U15197 (N_15197,N_7280,N_9959);
nor U15198 (N_15198,N_7153,N_6769);
xnor U15199 (N_15199,N_8962,N_11420);
and U15200 (N_15200,N_9726,N_9425);
xnor U15201 (N_15201,N_10660,N_6492);
or U15202 (N_15202,N_7067,N_9649);
nor U15203 (N_15203,N_12335,N_9693);
nor U15204 (N_15204,N_9583,N_12034);
xnor U15205 (N_15205,N_9153,N_6804);
xor U15206 (N_15206,N_11664,N_7291);
xor U15207 (N_15207,N_8160,N_11749);
nor U15208 (N_15208,N_11079,N_6756);
nor U15209 (N_15209,N_9946,N_8530);
nand U15210 (N_15210,N_7285,N_7748);
nor U15211 (N_15211,N_6363,N_11710);
or U15212 (N_15212,N_7821,N_11834);
nand U15213 (N_15213,N_12370,N_8870);
xor U15214 (N_15214,N_6674,N_8514);
xor U15215 (N_15215,N_6993,N_7468);
or U15216 (N_15216,N_8157,N_9572);
or U15217 (N_15217,N_8546,N_8512);
and U15218 (N_15218,N_7142,N_11206);
nand U15219 (N_15219,N_10470,N_7215);
nor U15220 (N_15220,N_9799,N_9587);
xnor U15221 (N_15221,N_11822,N_8839);
and U15222 (N_15222,N_11359,N_6800);
and U15223 (N_15223,N_7293,N_8231);
xnor U15224 (N_15224,N_11865,N_8869);
or U15225 (N_15225,N_12146,N_9505);
nand U15226 (N_15226,N_7369,N_8390);
or U15227 (N_15227,N_9668,N_7195);
xor U15228 (N_15228,N_8916,N_7608);
xor U15229 (N_15229,N_7940,N_8592);
nor U15230 (N_15230,N_6751,N_6700);
xor U15231 (N_15231,N_9842,N_9141);
nor U15232 (N_15232,N_9326,N_10893);
or U15233 (N_15233,N_7854,N_9659);
nand U15234 (N_15234,N_8360,N_10313);
nor U15235 (N_15235,N_11020,N_11324);
nand U15236 (N_15236,N_10371,N_11913);
nand U15237 (N_15237,N_7888,N_8988);
xnor U15238 (N_15238,N_8137,N_12460);
nand U15239 (N_15239,N_9211,N_11745);
xor U15240 (N_15240,N_7172,N_11052);
xor U15241 (N_15241,N_11857,N_11209);
or U15242 (N_15242,N_12134,N_8417);
and U15243 (N_15243,N_7226,N_8025);
xnor U15244 (N_15244,N_10533,N_6886);
nor U15245 (N_15245,N_8319,N_9595);
or U15246 (N_15246,N_11299,N_10561);
and U15247 (N_15247,N_9787,N_10647);
or U15248 (N_15248,N_10405,N_12290);
or U15249 (N_15249,N_10934,N_6526);
nor U15250 (N_15250,N_10118,N_7113);
nand U15251 (N_15251,N_11725,N_8503);
and U15252 (N_15252,N_11832,N_9398);
or U15253 (N_15253,N_8574,N_9062);
and U15254 (N_15254,N_11689,N_6614);
or U15255 (N_15255,N_6258,N_9922);
and U15256 (N_15256,N_11688,N_12089);
or U15257 (N_15257,N_10170,N_7760);
xnor U15258 (N_15258,N_9371,N_8842);
and U15259 (N_15259,N_9162,N_11063);
or U15260 (N_15260,N_12397,N_6729);
nand U15261 (N_15261,N_12315,N_12138);
nand U15262 (N_15262,N_7179,N_8974);
or U15263 (N_15263,N_6370,N_10705);
xor U15264 (N_15264,N_11771,N_7183);
nor U15265 (N_15265,N_11670,N_12051);
nor U15266 (N_15266,N_12070,N_10037);
nor U15267 (N_15267,N_6818,N_7997);
or U15268 (N_15268,N_11485,N_9192);
nor U15269 (N_15269,N_7374,N_9893);
nand U15270 (N_15270,N_11573,N_6672);
nor U15271 (N_15271,N_8790,N_8780);
xnor U15272 (N_15272,N_7842,N_11606);
and U15273 (N_15273,N_10671,N_8919);
xnor U15274 (N_15274,N_6891,N_7080);
nor U15275 (N_15275,N_11015,N_9356);
nor U15276 (N_15276,N_9640,N_10961);
or U15277 (N_15277,N_9900,N_12021);
xor U15278 (N_15278,N_9210,N_10260);
or U15279 (N_15279,N_11934,N_9624);
nand U15280 (N_15280,N_11120,N_8168);
nand U15281 (N_15281,N_10422,N_9504);
and U15282 (N_15282,N_6487,N_8461);
nor U15283 (N_15283,N_11214,N_10968);
xnor U15284 (N_15284,N_10506,N_7252);
nor U15285 (N_15285,N_7948,N_9328);
nand U15286 (N_15286,N_9289,N_6310);
and U15287 (N_15287,N_7081,N_11852);
or U15288 (N_15288,N_8003,N_7429);
xor U15289 (N_15289,N_11757,N_6744);
or U15290 (N_15290,N_8911,N_8049);
xor U15291 (N_15291,N_8701,N_12268);
xor U15292 (N_15292,N_9417,N_10109);
xnor U15293 (N_15293,N_7242,N_6862);
xnor U15294 (N_15294,N_8769,N_9538);
or U15295 (N_15295,N_11690,N_7316);
or U15296 (N_15296,N_7938,N_6389);
or U15297 (N_15297,N_6414,N_9650);
and U15298 (N_15298,N_11165,N_7426);
nand U15299 (N_15299,N_11071,N_11918);
nand U15300 (N_15300,N_10415,N_10446);
and U15301 (N_15301,N_8745,N_6402);
and U15302 (N_15302,N_11361,N_11192);
xor U15303 (N_15303,N_8171,N_10994);
or U15304 (N_15304,N_12100,N_7777);
xnor U15305 (N_15305,N_11620,N_7754);
and U15306 (N_15306,N_11642,N_7384);
nand U15307 (N_15307,N_8957,N_8837);
and U15308 (N_15308,N_7987,N_9675);
and U15309 (N_15309,N_11999,N_9173);
xnor U15310 (N_15310,N_6317,N_8359);
or U15311 (N_15311,N_10802,N_11450);
nand U15312 (N_15312,N_7311,N_7318);
or U15313 (N_15313,N_7371,N_12055);
nor U15314 (N_15314,N_9887,N_7747);
xnor U15315 (N_15315,N_10145,N_11886);
and U15316 (N_15316,N_12059,N_9178);
xor U15317 (N_15317,N_8466,N_7621);
nand U15318 (N_15318,N_6633,N_7978);
and U15319 (N_15319,N_7543,N_11423);
xor U15320 (N_15320,N_7965,N_11851);
or U15321 (N_15321,N_10342,N_7872);
or U15322 (N_15322,N_7644,N_12267);
and U15323 (N_15323,N_9957,N_12281);
and U15324 (N_15324,N_9724,N_8080);
xor U15325 (N_15325,N_10122,N_10093);
and U15326 (N_15326,N_6424,N_6931);
and U15327 (N_15327,N_9082,N_8071);
nor U15328 (N_15328,N_12188,N_9483);
nand U15329 (N_15329,N_8968,N_6305);
and U15330 (N_15330,N_6469,N_9977);
xnor U15331 (N_15331,N_7051,N_8949);
or U15332 (N_15332,N_9914,N_9077);
or U15333 (N_15333,N_10138,N_9291);
or U15334 (N_15334,N_7922,N_9582);
and U15335 (N_15335,N_9245,N_6611);
xnor U15336 (N_15336,N_8385,N_11827);
or U15337 (N_15337,N_11610,N_7750);
xnor U15338 (N_15338,N_11241,N_11738);
nand U15339 (N_15339,N_11895,N_11452);
nor U15340 (N_15340,N_7026,N_6388);
or U15341 (N_15341,N_11653,N_9772);
nor U15342 (N_15342,N_9516,N_12200);
xnor U15343 (N_15343,N_9958,N_10629);
nor U15344 (N_15344,N_6763,N_12307);
nor U15345 (N_15345,N_11381,N_8430);
xnor U15346 (N_15346,N_9202,N_7029);
nor U15347 (N_15347,N_11885,N_8039);
xor U15348 (N_15348,N_11396,N_9422);
or U15349 (N_15349,N_9603,N_7890);
and U15350 (N_15350,N_8148,N_6445);
xor U15351 (N_15351,N_7295,N_11195);
and U15352 (N_15352,N_11190,N_7268);
and U15353 (N_15353,N_9935,N_10926);
and U15354 (N_15354,N_8147,N_9680);
nand U15355 (N_15355,N_7806,N_6648);
and U15356 (N_15356,N_8440,N_7893);
xnor U15357 (N_15357,N_10475,N_8058);
xnor U15358 (N_15358,N_6680,N_6853);
nor U15359 (N_15359,N_11467,N_12115);
and U15360 (N_15360,N_11782,N_11519);
and U15361 (N_15361,N_6504,N_7692);
nor U15362 (N_15362,N_8107,N_9885);
nor U15363 (N_15363,N_12266,N_9491);
or U15364 (N_15364,N_9234,N_10136);
and U15365 (N_15365,N_8770,N_8420);
nand U15366 (N_15366,N_8823,N_11358);
nor U15367 (N_15367,N_7625,N_9769);
nor U15368 (N_15368,N_7813,N_12415);
and U15369 (N_15369,N_10670,N_10028);
or U15370 (N_15370,N_7697,N_8344);
xor U15371 (N_15371,N_12278,N_7653);
nor U15372 (N_15372,N_11317,N_8699);
and U15373 (N_15373,N_12491,N_10253);
xnor U15374 (N_15374,N_12306,N_9715);
xor U15375 (N_15375,N_9754,N_11340);
nand U15376 (N_15376,N_10969,N_7623);
and U15377 (N_15377,N_7989,N_12453);
or U15378 (N_15378,N_9844,N_11431);
nor U15379 (N_15379,N_8725,N_10194);
and U15380 (N_15380,N_8153,N_9040);
and U15381 (N_15381,N_11613,N_11859);
xor U15382 (N_15382,N_9442,N_10156);
or U15383 (N_15383,N_7135,N_11756);
nor U15384 (N_15384,N_10639,N_6364);
and U15385 (N_15385,N_11492,N_7640);
nor U15386 (N_15386,N_9556,N_8786);
nand U15387 (N_15387,N_6951,N_7745);
and U15388 (N_15388,N_10690,N_12447);
nor U15389 (N_15389,N_7018,N_6716);
nor U15390 (N_15390,N_8465,N_7820);
xnor U15391 (N_15391,N_8472,N_9599);
or U15392 (N_15392,N_6587,N_10430);
xor U15393 (N_15393,N_12156,N_10348);
xnor U15394 (N_15394,N_10285,N_9469);
nand U15395 (N_15395,N_12193,N_9444);
nor U15396 (N_15396,N_7899,N_8972);
nand U15397 (N_15397,N_8845,N_8656);
nand U15398 (N_15398,N_9370,N_7064);
nor U15399 (N_15399,N_6277,N_8118);
and U15400 (N_15400,N_10691,N_7145);
nand U15401 (N_15401,N_12301,N_8623);
nand U15402 (N_15402,N_12304,N_12337);
xnor U15403 (N_15403,N_11068,N_11924);
or U15404 (N_15404,N_10469,N_9561);
nand U15405 (N_15405,N_11816,N_9020);
xnor U15406 (N_15406,N_9349,N_10491);
or U15407 (N_15407,N_11660,N_9696);
or U15408 (N_15408,N_8002,N_12005);
xnor U15409 (N_15409,N_10783,N_6877);
nor U15410 (N_15410,N_10423,N_9115);
nor U15411 (N_15411,N_7650,N_6562);
xor U15412 (N_15412,N_7606,N_8290);
xnor U15413 (N_15413,N_9342,N_9792);
nor U15414 (N_15414,N_11412,N_11285);
nor U15415 (N_15415,N_8687,N_8030);
and U15416 (N_15416,N_11368,N_6896);
nor U15417 (N_15417,N_6743,N_10585);
nor U15418 (N_15418,N_10425,N_8277);
nor U15419 (N_15419,N_9898,N_6812);
xnor U15420 (N_15420,N_9546,N_8329);
or U15421 (N_15421,N_8425,N_11337);
nand U15422 (N_15422,N_11742,N_6604);
or U15423 (N_15423,N_7613,N_12245);
xnor U15424 (N_15424,N_9949,N_9669);
nand U15425 (N_15425,N_7617,N_10829);
nand U15426 (N_15426,N_8616,N_10502);
or U15427 (N_15427,N_11521,N_10112);
and U15428 (N_15428,N_9513,N_7314);
and U15429 (N_15429,N_8894,N_12166);
nand U15430 (N_15430,N_11922,N_6556);
xor U15431 (N_15431,N_7952,N_9288);
nor U15432 (N_15432,N_9134,N_7508);
and U15433 (N_15433,N_10658,N_11471);
nand U15434 (N_15434,N_6427,N_7859);
xnor U15435 (N_15435,N_8891,N_9629);
xor U15436 (N_15436,N_10538,N_6839);
nor U15437 (N_15437,N_6773,N_10901);
nand U15438 (N_15438,N_9248,N_6429);
and U15439 (N_15439,N_10014,N_8247);
xor U15440 (N_15440,N_11877,N_11680);
nor U15441 (N_15441,N_11122,N_10421);
xor U15442 (N_15442,N_7908,N_12028);
xor U15443 (N_15443,N_10088,N_11601);
or U15444 (N_15444,N_6979,N_11809);
or U15445 (N_15445,N_7132,N_8244);
xnor U15446 (N_15446,N_6668,N_10180);
or U15447 (N_15447,N_12291,N_10851);
xnor U15448 (N_15448,N_9720,N_8781);
nor U15449 (N_15449,N_9529,N_9709);
and U15450 (N_15450,N_6985,N_12340);
nor U15451 (N_15451,N_9622,N_10033);
or U15452 (N_15452,N_10397,N_6409);
nor U15453 (N_15453,N_10344,N_11145);
and U15454 (N_15454,N_10204,N_12405);
nor U15455 (N_15455,N_8652,N_10547);
nor U15456 (N_15456,N_6541,N_10219);
or U15457 (N_15457,N_10016,N_10640);
xor U15458 (N_15458,N_7322,N_7209);
nor U15459 (N_15459,N_12471,N_6858);
or U15460 (N_15460,N_10959,N_11061);
nand U15461 (N_15461,N_9467,N_7296);
nand U15462 (N_15462,N_7013,N_10715);
nand U15463 (N_15463,N_8478,N_10971);
or U15464 (N_15464,N_8893,N_8379);
nor U15465 (N_15465,N_6447,N_6534);
and U15466 (N_15466,N_9802,N_10598);
xor U15467 (N_15467,N_10762,N_12450);
or U15468 (N_15468,N_6465,N_8940);
nor U15469 (N_15469,N_7687,N_11550);
and U15470 (N_15470,N_7009,N_12189);
xnor U15471 (N_15471,N_9156,N_9604);
nand U15472 (N_15472,N_8586,N_11836);
xor U15473 (N_15473,N_11739,N_6547);
and U15474 (N_15474,N_11181,N_9955);
xor U15475 (N_15475,N_10796,N_11914);
xor U15476 (N_15476,N_7204,N_10531);
or U15477 (N_15477,N_6374,N_9758);
nand U15478 (N_15478,N_8204,N_7739);
nand U15479 (N_15479,N_11342,N_6802);
nor U15480 (N_15480,N_8217,N_12464);
nor U15481 (N_15481,N_8841,N_8755);
and U15482 (N_15482,N_10379,N_7967);
or U15483 (N_15483,N_7458,N_6477);
or U15484 (N_15484,N_10720,N_6426);
nor U15485 (N_15485,N_11831,N_9830);
nand U15486 (N_15486,N_7833,N_11645);
or U15487 (N_15487,N_9495,N_8130);
and U15488 (N_15488,N_8475,N_8040);
xnor U15489 (N_15489,N_6525,N_9479);
or U15490 (N_15490,N_12312,N_10075);
or U15491 (N_15491,N_6828,N_6264);
xor U15492 (N_15492,N_7387,N_7624);
nand U15493 (N_15493,N_10149,N_7216);
nor U15494 (N_15494,N_9102,N_8533);
or U15495 (N_15495,N_10866,N_11730);
nor U15496 (N_15496,N_7149,N_9240);
and U15497 (N_15497,N_12063,N_11841);
or U15498 (N_15498,N_8961,N_7752);
xor U15499 (N_15499,N_11614,N_8683);
and U15500 (N_15500,N_11759,N_8088);
nor U15501 (N_15501,N_12148,N_9052);
nor U15502 (N_15502,N_11539,N_8913);
xor U15503 (N_15503,N_6669,N_7117);
nor U15504 (N_15504,N_9837,N_12469);
xor U15505 (N_15505,N_7375,N_11603);
nor U15506 (N_15506,N_11619,N_7801);
or U15507 (N_15507,N_11375,N_10338);
nand U15508 (N_15508,N_11719,N_12082);
nor U15509 (N_15509,N_11476,N_9602);
nand U15510 (N_15510,N_8161,N_9489);
or U15511 (N_15511,N_10768,N_10872);
and U15512 (N_15512,N_6460,N_8627);
nor U15513 (N_15513,N_9257,N_11596);
or U15514 (N_15514,N_7259,N_9393);
xor U15515 (N_15515,N_9046,N_9751);
nand U15516 (N_15516,N_10003,N_8364);
or U15517 (N_15517,N_8625,N_7037);
and U15518 (N_15518,N_9653,N_10019);
or U15519 (N_15519,N_6974,N_9327);
nand U15520 (N_15520,N_7961,N_11721);
or U15521 (N_15521,N_11460,N_10330);
and U15522 (N_15522,N_12218,N_10907);
xnor U15523 (N_15523,N_12401,N_7161);
and U15524 (N_15524,N_7626,N_8059);
or U15525 (N_15525,N_9341,N_11510);
and U15526 (N_15526,N_6410,N_10464);
nor U15527 (N_15527,N_8766,N_7092);
and U15528 (N_15528,N_7136,N_10945);
nor U15529 (N_15529,N_8367,N_11397);
nand U15530 (N_15530,N_9766,N_8705);
nor U15531 (N_15531,N_10608,N_10584);
nor U15532 (N_15532,N_6412,N_10997);
xor U15533 (N_15533,N_6262,N_9811);
nor U15534 (N_15534,N_9376,N_9253);
xnor U15535 (N_15535,N_8119,N_11580);
nor U15536 (N_15536,N_6923,N_8900);
or U15537 (N_15537,N_6694,N_10373);
nand U15538 (N_15538,N_9482,N_7858);
nor U15539 (N_15539,N_10486,N_11562);
or U15540 (N_15540,N_6580,N_7784);
nor U15541 (N_15541,N_7548,N_7184);
nand U15542 (N_15542,N_12258,N_10341);
nand U15543 (N_15543,N_9161,N_10228);
xnor U15544 (N_15544,N_10209,N_9236);
nand U15545 (N_15545,N_7651,N_12247);
xor U15546 (N_15546,N_8703,N_7723);
xnor U15547 (N_15547,N_6905,N_9809);
or U15548 (N_15548,N_11854,N_12224);
xor U15549 (N_15549,N_9176,N_8740);
nand U15550 (N_15550,N_9555,N_9347);
nand U15551 (N_15551,N_6897,N_11848);
and U15552 (N_15552,N_11302,N_6782);
nor U15553 (N_15553,N_9063,N_10848);
xor U15554 (N_15554,N_8022,N_10090);
or U15555 (N_15555,N_8096,N_11380);
nand U15556 (N_15556,N_10546,N_6637);
nor U15557 (N_15557,N_9451,N_7871);
nor U15558 (N_15558,N_11405,N_10518);
or U15559 (N_15559,N_7878,N_9916);
xnor U15560 (N_15560,N_10799,N_9994);
nand U15561 (N_15561,N_11007,N_9430);
or U15562 (N_15562,N_8788,N_7994);
and U15563 (N_15563,N_7904,N_9609);
and U15564 (N_15564,N_6760,N_8353);
xor U15565 (N_15565,N_6566,N_11676);
nand U15566 (N_15566,N_7749,N_7568);
nor U15567 (N_15567,N_11303,N_10750);
or U15568 (N_15568,N_8271,N_9590);
or U15569 (N_15569,N_8793,N_11384);
or U15570 (N_15570,N_9438,N_8765);
and U15571 (N_15571,N_6809,N_8017);
nor U15572 (N_15572,N_11957,N_9086);
and U15573 (N_15573,N_8045,N_9713);
nand U15574 (N_15574,N_10788,N_8915);
nand U15575 (N_15575,N_10346,N_8111);
and U15576 (N_15576,N_11940,N_9309);
nand U15577 (N_15577,N_10140,N_7074);
or U15578 (N_15578,N_11665,N_10023);
or U15579 (N_15579,N_7717,N_8824);
and U15580 (N_15580,N_9250,N_12075);
or U15581 (N_15581,N_9873,N_8494);
xor U15582 (N_15582,N_9722,N_8682);
and U15583 (N_15583,N_11227,N_6946);
nor U15584 (N_15584,N_7046,N_7003);
xnor U15585 (N_15585,N_10677,N_10074);
nor U15586 (N_15586,N_7083,N_8352);
xor U15587 (N_15587,N_10741,N_6564);
xor U15588 (N_15588,N_11585,N_10437);
and U15589 (N_15589,N_8254,N_7923);
nand U15590 (N_15590,N_6517,N_6362);
xor U15591 (N_15591,N_9246,N_6344);
nor U15592 (N_15592,N_9448,N_9804);
xor U15593 (N_15593,N_12229,N_9148);
or U15594 (N_15594,N_11764,N_10139);
and U15595 (N_15595,N_9851,N_12440);
nand U15596 (N_15596,N_6852,N_8249);
or U15597 (N_15597,N_12442,N_11296);
or U15598 (N_15598,N_7307,N_11537);
and U15599 (N_15599,N_7524,N_7610);
or U15600 (N_15600,N_8560,N_6404);
or U15601 (N_15601,N_6468,N_6518);
and U15602 (N_15602,N_6607,N_10350);
nor U15603 (N_15603,N_8587,N_9242);
and U15604 (N_15604,N_12336,N_7992);
xor U15605 (N_15605,N_9707,N_10213);
nor U15606 (N_15606,N_11729,N_8677);
or U15607 (N_15607,N_7234,N_11709);
xor U15608 (N_15608,N_9191,N_10729);
xor U15609 (N_15609,N_9421,N_6784);
nand U15610 (N_15610,N_9881,N_8397);
and U15611 (N_15611,N_6458,N_11654);
nand U15612 (N_15612,N_11682,N_10745);
nor U15613 (N_15613,N_7567,N_6664);
nor U15614 (N_15614,N_6837,N_8362);
nor U15615 (N_15615,N_9154,N_6472);
nand U15616 (N_15616,N_7100,N_10641);
nand U15617 (N_15617,N_9135,N_12029);
and U15618 (N_15618,N_12223,N_6608);
xor U15619 (N_15619,N_11805,N_11305);
nand U15620 (N_15620,N_9308,N_10952);
or U15621 (N_15621,N_11552,N_9674);
xnor U15622 (N_15622,N_11703,N_10751);
and U15623 (N_15623,N_9552,N_9353);
nand U15624 (N_15624,N_8661,N_10224);
nor U15625 (N_15625,N_12028,N_8645);
or U15626 (N_15626,N_9623,N_8650);
nor U15627 (N_15627,N_9321,N_9231);
nand U15628 (N_15628,N_9826,N_6875);
and U15629 (N_15629,N_8689,N_9579);
nor U15630 (N_15630,N_10239,N_10860);
and U15631 (N_15631,N_8898,N_11332);
nor U15632 (N_15632,N_11137,N_7899);
or U15633 (N_15633,N_11790,N_10741);
or U15634 (N_15634,N_9230,N_10155);
nand U15635 (N_15635,N_10748,N_8631);
nor U15636 (N_15636,N_7223,N_11931);
nand U15637 (N_15637,N_7577,N_7960);
and U15638 (N_15638,N_7136,N_10972);
xor U15639 (N_15639,N_11342,N_10146);
xnor U15640 (N_15640,N_11827,N_8188);
xor U15641 (N_15641,N_11579,N_11648);
xor U15642 (N_15642,N_6925,N_6539);
xor U15643 (N_15643,N_10657,N_10532);
and U15644 (N_15644,N_6815,N_11474);
and U15645 (N_15645,N_11237,N_6658);
or U15646 (N_15646,N_10965,N_10761);
xnor U15647 (N_15647,N_11188,N_11263);
nand U15648 (N_15648,N_9956,N_7222);
nand U15649 (N_15649,N_9988,N_7724);
and U15650 (N_15650,N_10235,N_12203);
or U15651 (N_15651,N_10496,N_9363);
or U15652 (N_15652,N_10001,N_8806);
xor U15653 (N_15653,N_10768,N_9538);
and U15654 (N_15654,N_8279,N_8874);
or U15655 (N_15655,N_6674,N_10739);
and U15656 (N_15656,N_6567,N_7267);
or U15657 (N_15657,N_8181,N_8281);
nand U15658 (N_15658,N_7798,N_6534);
nand U15659 (N_15659,N_7832,N_8082);
xnor U15660 (N_15660,N_10103,N_10276);
and U15661 (N_15661,N_7377,N_8346);
nor U15662 (N_15662,N_10903,N_7354);
nor U15663 (N_15663,N_6750,N_6902);
nand U15664 (N_15664,N_9547,N_7351);
or U15665 (N_15665,N_8152,N_8387);
and U15666 (N_15666,N_12469,N_8322);
xor U15667 (N_15667,N_11675,N_8224);
nand U15668 (N_15668,N_12268,N_12087);
nor U15669 (N_15669,N_11475,N_8055);
and U15670 (N_15670,N_7477,N_10129);
and U15671 (N_15671,N_12086,N_7782);
or U15672 (N_15672,N_12054,N_10417);
nand U15673 (N_15673,N_6608,N_7225);
nor U15674 (N_15674,N_11871,N_10572);
nand U15675 (N_15675,N_10061,N_7424);
nor U15676 (N_15676,N_8541,N_10454);
nor U15677 (N_15677,N_9533,N_9944);
nand U15678 (N_15678,N_10500,N_7493);
nor U15679 (N_15679,N_6728,N_6682);
nor U15680 (N_15680,N_10055,N_7372);
or U15681 (N_15681,N_12459,N_9868);
and U15682 (N_15682,N_10009,N_11495);
xor U15683 (N_15683,N_9490,N_8282);
xor U15684 (N_15684,N_12359,N_12143);
and U15685 (N_15685,N_11074,N_7060);
and U15686 (N_15686,N_8576,N_11331);
nand U15687 (N_15687,N_12347,N_10880);
nand U15688 (N_15688,N_8333,N_10706);
xor U15689 (N_15689,N_10190,N_9515);
xnor U15690 (N_15690,N_12268,N_10701);
nand U15691 (N_15691,N_9144,N_7867);
or U15692 (N_15692,N_10185,N_7179);
nor U15693 (N_15693,N_8510,N_9028);
nand U15694 (N_15694,N_11431,N_9429);
and U15695 (N_15695,N_7007,N_11533);
or U15696 (N_15696,N_10956,N_8711);
xor U15697 (N_15697,N_12335,N_10661);
xor U15698 (N_15698,N_9054,N_9171);
nor U15699 (N_15699,N_7043,N_9498);
nand U15700 (N_15700,N_11273,N_8675);
and U15701 (N_15701,N_7749,N_6884);
xor U15702 (N_15702,N_11578,N_8937);
or U15703 (N_15703,N_9755,N_12359);
nor U15704 (N_15704,N_10754,N_8850);
nand U15705 (N_15705,N_10027,N_6423);
nand U15706 (N_15706,N_11293,N_9564);
xor U15707 (N_15707,N_6697,N_9135);
or U15708 (N_15708,N_12258,N_10658);
xor U15709 (N_15709,N_10405,N_9558);
nor U15710 (N_15710,N_7110,N_10915);
nand U15711 (N_15711,N_8352,N_11087);
xnor U15712 (N_15712,N_11380,N_12229);
nor U15713 (N_15713,N_8733,N_12285);
or U15714 (N_15714,N_10669,N_12490);
and U15715 (N_15715,N_8999,N_7371);
and U15716 (N_15716,N_11579,N_6896);
xor U15717 (N_15717,N_9520,N_8544);
or U15718 (N_15718,N_8311,N_11867);
nor U15719 (N_15719,N_12359,N_7689);
xnor U15720 (N_15720,N_8239,N_7436);
xor U15721 (N_15721,N_9138,N_11514);
or U15722 (N_15722,N_6424,N_7325);
and U15723 (N_15723,N_7680,N_11903);
xor U15724 (N_15724,N_9918,N_11919);
or U15725 (N_15725,N_11300,N_11719);
xnor U15726 (N_15726,N_11234,N_11850);
xnor U15727 (N_15727,N_10033,N_7631);
or U15728 (N_15728,N_7736,N_11659);
nor U15729 (N_15729,N_11934,N_11609);
nand U15730 (N_15730,N_12218,N_6790);
xor U15731 (N_15731,N_9670,N_12223);
nand U15732 (N_15732,N_7542,N_10865);
and U15733 (N_15733,N_9269,N_7149);
xor U15734 (N_15734,N_6267,N_11679);
nor U15735 (N_15735,N_11412,N_9254);
xor U15736 (N_15736,N_8724,N_7096);
and U15737 (N_15737,N_8816,N_9235);
xor U15738 (N_15738,N_9869,N_11303);
xnor U15739 (N_15739,N_7195,N_12354);
nand U15740 (N_15740,N_9350,N_8389);
and U15741 (N_15741,N_11957,N_9420);
and U15742 (N_15742,N_6809,N_6772);
xor U15743 (N_15743,N_8147,N_10006);
nor U15744 (N_15744,N_8354,N_8824);
and U15745 (N_15745,N_9426,N_6865);
and U15746 (N_15746,N_11880,N_7389);
nor U15747 (N_15747,N_6857,N_6685);
xor U15748 (N_15748,N_6862,N_6976);
or U15749 (N_15749,N_9276,N_11107);
nand U15750 (N_15750,N_10839,N_7982);
and U15751 (N_15751,N_7272,N_8213);
or U15752 (N_15752,N_8991,N_6725);
nor U15753 (N_15753,N_7217,N_11378);
nand U15754 (N_15754,N_10279,N_6580);
nor U15755 (N_15755,N_9271,N_12201);
nor U15756 (N_15756,N_7986,N_11993);
nor U15757 (N_15757,N_12405,N_12249);
nand U15758 (N_15758,N_7335,N_11391);
or U15759 (N_15759,N_7769,N_7467);
and U15760 (N_15760,N_8690,N_12000);
or U15761 (N_15761,N_11267,N_6875);
and U15762 (N_15762,N_10123,N_12032);
nor U15763 (N_15763,N_9205,N_8081);
or U15764 (N_15764,N_10983,N_11094);
or U15765 (N_15765,N_9681,N_6270);
nand U15766 (N_15766,N_11958,N_11224);
and U15767 (N_15767,N_7653,N_9494);
nand U15768 (N_15768,N_7236,N_9067);
xor U15769 (N_15769,N_6429,N_11121);
nor U15770 (N_15770,N_9822,N_10226);
xnor U15771 (N_15771,N_10393,N_10215);
xor U15772 (N_15772,N_7205,N_10982);
and U15773 (N_15773,N_9797,N_10001);
nand U15774 (N_15774,N_10189,N_7955);
nor U15775 (N_15775,N_9669,N_8145);
and U15776 (N_15776,N_11960,N_6489);
and U15777 (N_15777,N_11625,N_11862);
or U15778 (N_15778,N_11752,N_6582);
or U15779 (N_15779,N_9162,N_6737);
or U15780 (N_15780,N_7076,N_9644);
or U15781 (N_15781,N_10562,N_6290);
nor U15782 (N_15782,N_10050,N_7144);
xor U15783 (N_15783,N_10164,N_8663);
or U15784 (N_15784,N_11689,N_11875);
xnor U15785 (N_15785,N_9487,N_7219);
and U15786 (N_15786,N_11215,N_11487);
nor U15787 (N_15787,N_8175,N_9413);
nand U15788 (N_15788,N_9565,N_8832);
nor U15789 (N_15789,N_6261,N_11457);
and U15790 (N_15790,N_7361,N_11353);
xor U15791 (N_15791,N_8281,N_9667);
nor U15792 (N_15792,N_8234,N_6869);
and U15793 (N_15793,N_9847,N_10113);
nor U15794 (N_15794,N_8070,N_8193);
nand U15795 (N_15795,N_12153,N_10055);
and U15796 (N_15796,N_7712,N_11702);
nand U15797 (N_15797,N_12491,N_7683);
xnor U15798 (N_15798,N_10988,N_7747);
and U15799 (N_15799,N_9839,N_8794);
nand U15800 (N_15800,N_11035,N_7723);
or U15801 (N_15801,N_9953,N_8021);
and U15802 (N_15802,N_11762,N_6523);
xor U15803 (N_15803,N_10752,N_6781);
xor U15804 (N_15804,N_9739,N_7833);
or U15805 (N_15805,N_12423,N_8837);
nor U15806 (N_15806,N_10590,N_9127);
xnor U15807 (N_15807,N_10588,N_8129);
and U15808 (N_15808,N_10444,N_11229);
nand U15809 (N_15809,N_7058,N_7432);
or U15810 (N_15810,N_10940,N_8925);
nor U15811 (N_15811,N_10388,N_6673);
and U15812 (N_15812,N_8799,N_6603);
nand U15813 (N_15813,N_8774,N_9467);
and U15814 (N_15814,N_10651,N_11025);
and U15815 (N_15815,N_10083,N_8187);
and U15816 (N_15816,N_8723,N_11735);
nor U15817 (N_15817,N_12171,N_11755);
nand U15818 (N_15818,N_7166,N_10452);
nor U15819 (N_15819,N_7101,N_10154);
and U15820 (N_15820,N_7041,N_8323);
or U15821 (N_15821,N_7586,N_6947);
and U15822 (N_15822,N_11118,N_11694);
or U15823 (N_15823,N_10433,N_11925);
or U15824 (N_15824,N_9072,N_6991);
nor U15825 (N_15825,N_10369,N_10489);
nand U15826 (N_15826,N_9812,N_11917);
or U15827 (N_15827,N_9947,N_7772);
xor U15828 (N_15828,N_10837,N_7673);
nor U15829 (N_15829,N_7481,N_9379);
xor U15830 (N_15830,N_6990,N_11564);
nand U15831 (N_15831,N_11266,N_11543);
or U15832 (N_15832,N_7748,N_9633);
and U15833 (N_15833,N_8879,N_8105);
xor U15834 (N_15834,N_9323,N_7096);
and U15835 (N_15835,N_8496,N_11904);
or U15836 (N_15836,N_10404,N_6909);
and U15837 (N_15837,N_11255,N_10590);
and U15838 (N_15838,N_11253,N_11496);
and U15839 (N_15839,N_8222,N_12493);
and U15840 (N_15840,N_9730,N_9167);
nor U15841 (N_15841,N_12449,N_8904);
xor U15842 (N_15842,N_6542,N_7738);
nor U15843 (N_15843,N_7208,N_8319);
nand U15844 (N_15844,N_9885,N_9245);
nor U15845 (N_15845,N_11628,N_7112);
nor U15846 (N_15846,N_7624,N_7175);
or U15847 (N_15847,N_10791,N_12104);
nand U15848 (N_15848,N_9920,N_11961);
and U15849 (N_15849,N_8623,N_7804);
xor U15850 (N_15850,N_10826,N_6910);
xor U15851 (N_15851,N_12235,N_11022);
xor U15852 (N_15852,N_9237,N_10582);
xnor U15853 (N_15853,N_9233,N_10114);
and U15854 (N_15854,N_9567,N_8702);
nand U15855 (N_15855,N_7184,N_9309);
nand U15856 (N_15856,N_10630,N_9484);
nand U15857 (N_15857,N_9828,N_10599);
nand U15858 (N_15858,N_8648,N_6770);
or U15859 (N_15859,N_8608,N_7273);
nor U15860 (N_15860,N_10263,N_9477);
nor U15861 (N_15861,N_12092,N_7813);
nor U15862 (N_15862,N_12448,N_12199);
nor U15863 (N_15863,N_8088,N_12104);
or U15864 (N_15864,N_9650,N_10907);
or U15865 (N_15865,N_9075,N_10497);
xnor U15866 (N_15866,N_9599,N_9195);
xnor U15867 (N_15867,N_9286,N_10122);
nor U15868 (N_15868,N_9605,N_9639);
xor U15869 (N_15869,N_9542,N_11771);
nand U15870 (N_15870,N_6974,N_11375);
nor U15871 (N_15871,N_8492,N_7576);
nand U15872 (N_15872,N_9723,N_6915);
or U15873 (N_15873,N_7226,N_7889);
nand U15874 (N_15874,N_10370,N_10285);
xor U15875 (N_15875,N_11727,N_6440);
nand U15876 (N_15876,N_9486,N_11219);
and U15877 (N_15877,N_7717,N_9425);
and U15878 (N_15878,N_7219,N_8593);
nand U15879 (N_15879,N_9385,N_11225);
or U15880 (N_15880,N_11509,N_11803);
nand U15881 (N_15881,N_9217,N_10158);
or U15882 (N_15882,N_12366,N_9480);
or U15883 (N_15883,N_7167,N_9848);
nor U15884 (N_15884,N_9860,N_7511);
nor U15885 (N_15885,N_6706,N_8003);
xnor U15886 (N_15886,N_8090,N_8435);
nand U15887 (N_15887,N_7398,N_8394);
or U15888 (N_15888,N_10110,N_9515);
nor U15889 (N_15889,N_9737,N_10406);
nand U15890 (N_15890,N_12063,N_6889);
or U15891 (N_15891,N_6449,N_6617);
nor U15892 (N_15892,N_9130,N_9741);
xor U15893 (N_15893,N_11609,N_6297);
nor U15894 (N_15894,N_8193,N_8789);
and U15895 (N_15895,N_10041,N_7728);
nand U15896 (N_15896,N_6856,N_10946);
nor U15897 (N_15897,N_7095,N_8006);
nor U15898 (N_15898,N_8723,N_9392);
nand U15899 (N_15899,N_10798,N_6715);
nor U15900 (N_15900,N_6300,N_10800);
and U15901 (N_15901,N_9761,N_8841);
nand U15902 (N_15902,N_11416,N_11674);
xor U15903 (N_15903,N_6272,N_11540);
and U15904 (N_15904,N_12110,N_9742);
and U15905 (N_15905,N_10864,N_8853);
nor U15906 (N_15906,N_10760,N_11140);
nor U15907 (N_15907,N_7028,N_12165);
or U15908 (N_15908,N_10932,N_8743);
xnor U15909 (N_15909,N_8947,N_12478);
or U15910 (N_15910,N_8527,N_10584);
nand U15911 (N_15911,N_11531,N_10720);
and U15912 (N_15912,N_7550,N_9393);
xnor U15913 (N_15913,N_10067,N_7672);
xnor U15914 (N_15914,N_11567,N_8906);
nor U15915 (N_15915,N_9300,N_11514);
or U15916 (N_15916,N_11533,N_8275);
or U15917 (N_15917,N_7612,N_8466);
nand U15918 (N_15918,N_9382,N_6790);
or U15919 (N_15919,N_6697,N_10754);
and U15920 (N_15920,N_7007,N_11236);
or U15921 (N_15921,N_11702,N_10187);
nor U15922 (N_15922,N_8512,N_11044);
nor U15923 (N_15923,N_8229,N_12491);
or U15924 (N_15924,N_8144,N_6754);
or U15925 (N_15925,N_7303,N_7076);
or U15926 (N_15926,N_11803,N_12067);
and U15927 (N_15927,N_10311,N_9851);
nand U15928 (N_15928,N_11292,N_8442);
or U15929 (N_15929,N_6773,N_12128);
xnor U15930 (N_15930,N_12312,N_8157);
xor U15931 (N_15931,N_6710,N_9586);
xor U15932 (N_15932,N_11555,N_9941);
xnor U15933 (N_15933,N_11994,N_10275);
or U15934 (N_15934,N_9187,N_10845);
nand U15935 (N_15935,N_9277,N_6574);
nand U15936 (N_15936,N_6825,N_9532);
xnor U15937 (N_15937,N_11724,N_10227);
and U15938 (N_15938,N_8194,N_9576);
and U15939 (N_15939,N_9227,N_9720);
or U15940 (N_15940,N_8723,N_7278);
or U15941 (N_15941,N_8707,N_6372);
or U15942 (N_15942,N_9463,N_12423);
xnor U15943 (N_15943,N_11050,N_7338);
nor U15944 (N_15944,N_10667,N_10222);
xor U15945 (N_15945,N_10377,N_11122);
xnor U15946 (N_15946,N_8504,N_10954);
nand U15947 (N_15947,N_8968,N_7247);
or U15948 (N_15948,N_9001,N_10290);
and U15949 (N_15949,N_10299,N_10312);
xor U15950 (N_15950,N_9012,N_9468);
or U15951 (N_15951,N_10937,N_9576);
and U15952 (N_15952,N_11386,N_8910);
nor U15953 (N_15953,N_10974,N_9036);
xor U15954 (N_15954,N_7729,N_8497);
nor U15955 (N_15955,N_10323,N_8897);
and U15956 (N_15956,N_10545,N_11174);
xor U15957 (N_15957,N_7795,N_10233);
xnor U15958 (N_15958,N_7061,N_10026);
or U15959 (N_15959,N_6423,N_12445);
xor U15960 (N_15960,N_10270,N_7112);
and U15961 (N_15961,N_7098,N_7652);
xor U15962 (N_15962,N_11098,N_6424);
nand U15963 (N_15963,N_8153,N_11214);
nor U15964 (N_15964,N_10832,N_9913);
or U15965 (N_15965,N_8739,N_7895);
or U15966 (N_15966,N_11390,N_6840);
nand U15967 (N_15967,N_11196,N_10473);
xnor U15968 (N_15968,N_10155,N_11662);
nand U15969 (N_15969,N_10065,N_11690);
or U15970 (N_15970,N_12151,N_7045);
nand U15971 (N_15971,N_8622,N_7450);
xnor U15972 (N_15972,N_10039,N_10826);
nor U15973 (N_15973,N_7603,N_10647);
nor U15974 (N_15974,N_8144,N_8026);
xnor U15975 (N_15975,N_12244,N_7920);
nand U15976 (N_15976,N_10700,N_10415);
nor U15977 (N_15977,N_10779,N_6366);
nor U15978 (N_15978,N_12030,N_10388);
xor U15979 (N_15979,N_8806,N_12427);
nand U15980 (N_15980,N_9042,N_8036);
xnor U15981 (N_15981,N_6878,N_10115);
xnor U15982 (N_15982,N_7092,N_9741);
and U15983 (N_15983,N_10612,N_6414);
xnor U15984 (N_15984,N_10757,N_8187);
and U15985 (N_15985,N_6886,N_6844);
nand U15986 (N_15986,N_10730,N_11019);
nand U15987 (N_15987,N_9935,N_9877);
or U15988 (N_15988,N_9644,N_9146);
and U15989 (N_15989,N_9850,N_9728);
or U15990 (N_15990,N_8237,N_11481);
or U15991 (N_15991,N_9376,N_9059);
and U15992 (N_15992,N_11376,N_7887);
xor U15993 (N_15993,N_10409,N_8346);
xnor U15994 (N_15994,N_6986,N_11000);
xnor U15995 (N_15995,N_10160,N_11933);
or U15996 (N_15996,N_9468,N_12309);
or U15997 (N_15997,N_9186,N_11145);
nor U15998 (N_15998,N_8509,N_9721);
or U15999 (N_15999,N_10722,N_10159);
or U16000 (N_16000,N_11905,N_10387);
or U16001 (N_16001,N_8527,N_8971);
nand U16002 (N_16002,N_8269,N_6814);
or U16003 (N_16003,N_8347,N_7512);
xor U16004 (N_16004,N_10662,N_6872);
and U16005 (N_16005,N_8624,N_7058);
nor U16006 (N_16006,N_11712,N_7991);
xnor U16007 (N_16007,N_10174,N_8848);
nor U16008 (N_16008,N_10390,N_8643);
xnor U16009 (N_16009,N_8137,N_7890);
xnor U16010 (N_16010,N_11791,N_11069);
xnor U16011 (N_16011,N_8328,N_10757);
and U16012 (N_16012,N_6982,N_6786);
nor U16013 (N_16013,N_10251,N_8585);
nand U16014 (N_16014,N_9367,N_10669);
xnor U16015 (N_16015,N_7637,N_7025);
nand U16016 (N_16016,N_8248,N_11807);
or U16017 (N_16017,N_11762,N_9437);
or U16018 (N_16018,N_12064,N_8672);
nand U16019 (N_16019,N_9749,N_11228);
nor U16020 (N_16020,N_9808,N_8840);
and U16021 (N_16021,N_10879,N_6281);
or U16022 (N_16022,N_12139,N_12210);
and U16023 (N_16023,N_10450,N_7876);
nor U16024 (N_16024,N_9730,N_8897);
or U16025 (N_16025,N_12223,N_11710);
xor U16026 (N_16026,N_9548,N_6864);
xor U16027 (N_16027,N_6463,N_11910);
nor U16028 (N_16028,N_7521,N_11616);
xnor U16029 (N_16029,N_8782,N_10443);
xnor U16030 (N_16030,N_6853,N_11386);
and U16031 (N_16031,N_7132,N_12055);
nor U16032 (N_16032,N_10366,N_11479);
nand U16033 (N_16033,N_9620,N_11285);
nor U16034 (N_16034,N_11055,N_6501);
nand U16035 (N_16035,N_10520,N_10102);
xnor U16036 (N_16036,N_7417,N_10107);
or U16037 (N_16037,N_8258,N_11454);
xor U16038 (N_16038,N_12206,N_8414);
xnor U16039 (N_16039,N_11338,N_10542);
xor U16040 (N_16040,N_7839,N_10365);
xor U16041 (N_16041,N_8246,N_11971);
xor U16042 (N_16042,N_12025,N_6756);
or U16043 (N_16043,N_9878,N_12458);
nand U16044 (N_16044,N_8724,N_6437);
xnor U16045 (N_16045,N_6773,N_9926);
xor U16046 (N_16046,N_12008,N_9831);
nor U16047 (N_16047,N_11579,N_11970);
xor U16048 (N_16048,N_7670,N_9427);
nor U16049 (N_16049,N_8640,N_8229);
nand U16050 (N_16050,N_9438,N_10408);
xor U16051 (N_16051,N_8369,N_12119);
nand U16052 (N_16052,N_8935,N_10391);
or U16053 (N_16053,N_7663,N_7352);
nor U16054 (N_16054,N_8376,N_11959);
nand U16055 (N_16055,N_6742,N_10547);
xnor U16056 (N_16056,N_11285,N_10555);
and U16057 (N_16057,N_10596,N_10139);
and U16058 (N_16058,N_6456,N_9347);
nor U16059 (N_16059,N_7087,N_10759);
nor U16060 (N_16060,N_6981,N_8517);
and U16061 (N_16061,N_9693,N_10372);
and U16062 (N_16062,N_12468,N_10866);
nand U16063 (N_16063,N_8940,N_10868);
and U16064 (N_16064,N_9229,N_7503);
nand U16065 (N_16065,N_11937,N_10925);
or U16066 (N_16066,N_8395,N_6991);
nand U16067 (N_16067,N_10561,N_11614);
nor U16068 (N_16068,N_7616,N_9522);
xor U16069 (N_16069,N_7491,N_11791);
nand U16070 (N_16070,N_7388,N_6934);
nand U16071 (N_16071,N_7361,N_10497);
xor U16072 (N_16072,N_8504,N_8960);
nand U16073 (N_16073,N_7921,N_8781);
or U16074 (N_16074,N_6974,N_7025);
or U16075 (N_16075,N_9362,N_6331);
xor U16076 (N_16076,N_7535,N_12364);
xnor U16077 (N_16077,N_12256,N_10043);
nor U16078 (N_16078,N_9093,N_11096);
nand U16079 (N_16079,N_11335,N_8961);
nand U16080 (N_16080,N_10477,N_8946);
or U16081 (N_16081,N_7957,N_12265);
nor U16082 (N_16082,N_10532,N_8302);
or U16083 (N_16083,N_12415,N_9109);
and U16084 (N_16084,N_10576,N_8019);
or U16085 (N_16085,N_7561,N_11812);
nor U16086 (N_16086,N_10478,N_7505);
nand U16087 (N_16087,N_8963,N_7660);
or U16088 (N_16088,N_7776,N_11285);
nand U16089 (N_16089,N_7395,N_9815);
or U16090 (N_16090,N_6570,N_12447);
nand U16091 (N_16091,N_8331,N_11659);
nand U16092 (N_16092,N_7073,N_8345);
nand U16093 (N_16093,N_8638,N_7412);
nand U16094 (N_16094,N_6901,N_10699);
nor U16095 (N_16095,N_7315,N_8335);
nand U16096 (N_16096,N_12296,N_6927);
nand U16097 (N_16097,N_8328,N_8828);
nand U16098 (N_16098,N_10621,N_9168);
or U16099 (N_16099,N_8410,N_8221);
nor U16100 (N_16100,N_8866,N_8294);
or U16101 (N_16101,N_6712,N_7813);
nor U16102 (N_16102,N_11945,N_12126);
nor U16103 (N_16103,N_10651,N_10251);
nand U16104 (N_16104,N_8174,N_6292);
and U16105 (N_16105,N_6408,N_7764);
and U16106 (N_16106,N_6607,N_6466);
nor U16107 (N_16107,N_11943,N_8503);
nor U16108 (N_16108,N_10292,N_8450);
or U16109 (N_16109,N_11101,N_11945);
nand U16110 (N_16110,N_9137,N_9172);
or U16111 (N_16111,N_9390,N_11259);
and U16112 (N_16112,N_6264,N_8415);
xnor U16113 (N_16113,N_8441,N_7423);
and U16114 (N_16114,N_8837,N_11327);
nand U16115 (N_16115,N_7260,N_8690);
nand U16116 (N_16116,N_7546,N_7011);
nand U16117 (N_16117,N_6851,N_12441);
xor U16118 (N_16118,N_11429,N_7724);
nor U16119 (N_16119,N_10317,N_9415);
and U16120 (N_16120,N_8602,N_8741);
nand U16121 (N_16121,N_11101,N_10718);
nor U16122 (N_16122,N_8127,N_11377);
nand U16123 (N_16123,N_12007,N_11109);
and U16124 (N_16124,N_8634,N_7456);
xor U16125 (N_16125,N_6580,N_10061);
and U16126 (N_16126,N_11357,N_8070);
nor U16127 (N_16127,N_12107,N_11173);
nand U16128 (N_16128,N_6365,N_11501);
xor U16129 (N_16129,N_7698,N_8123);
nor U16130 (N_16130,N_6875,N_12435);
or U16131 (N_16131,N_6784,N_8777);
xor U16132 (N_16132,N_8081,N_11631);
or U16133 (N_16133,N_8343,N_9179);
nor U16134 (N_16134,N_7477,N_12030);
nor U16135 (N_16135,N_8669,N_8550);
or U16136 (N_16136,N_10051,N_9492);
nand U16137 (N_16137,N_8038,N_8011);
and U16138 (N_16138,N_7285,N_10506);
nor U16139 (N_16139,N_10621,N_8664);
nand U16140 (N_16140,N_11580,N_10726);
nor U16141 (N_16141,N_12132,N_11052);
xnor U16142 (N_16142,N_9649,N_8739);
xnor U16143 (N_16143,N_9608,N_12482);
or U16144 (N_16144,N_10593,N_9335);
or U16145 (N_16145,N_9010,N_8114);
nand U16146 (N_16146,N_9142,N_9960);
or U16147 (N_16147,N_8087,N_10891);
or U16148 (N_16148,N_10738,N_6270);
or U16149 (N_16149,N_6751,N_11696);
and U16150 (N_16150,N_9742,N_8758);
nand U16151 (N_16151,N_10696,N_10416);
nor U16152 (N_16152,N_7707,N_11936);
nand U16153 (N_16153,N_8305,N_7457);
or U16154 (N_16154,N_11545,N_8471);
xor U16155 (N_16155,N_10648,N_12424);
xor U16156 (N_16156,N_7235,N_9031);
nor U16157 (N_16157,N_8207,N_12084);
or U16158 (N_16158,N_9733,N_8072);
and U16159 (N_16159,N_7431,N_7245);
xor U16160 (N_16160,N_8979,N_8177);
xnor U16161 (N_16161,N_9184,N_10067);
and U16162 (N_16162,N_10293,N_12303);
xnor U16163 (N_16163,N_9228,N_9809);
nor U16164 (N_16164,N_6842,N_11115);
or U16165 (N_16165,N_12262,N_10405);
or U16166 (N_16166,N_9141,N_9657);
xnor U16167 (N_16167,N_6508,N_7393);
xor U16168 (N_16168,N_9191,N_9319);
nand U16169 (N_16169,N_10720,N_9987);
nor U16170 (N_16170,N_9638,N_7239);
and U16171 (N_16171,N_6323,N_11378);
and U16172 (N_16172,N_9043,N_9903);
nor U16173 (N_16173,N_11087,N_11341);
nor U16174 (N_16174,N_9860,N_6492);
nand U16175 (N_16175,N_7000,N_7889);
nand U16176 (N_16176,N_10816,N_7216);
nor U16177 (N_16177,N_9600,N_9207);
and U16178 (N_16178,N_9972,N_7432);
nor U16179 (N_16179,N_10482,N_8904);
or U16180 (N_16180,N_9201,N_8408);
xor U16181 (N_16181,N_10708,N_11978);
nor U16182 (N_16182,N_10014,N_8891);
and U16183 (N_16183,N_10975,N_8843);
nor U16184 (N_16184,N_9407,N_6489);
or U16185 (N_16185,N_6680,N_9663);
or U16186 (N_16186,N_7114,N_7353);
nand U16187 (N_16187,N_9176,N_9869);
nand U16188 (N_16188,N_10240,N_6795);
and U16189 (N_16189,N_7222,N_8930);
nand U16190 (N_16190,N_10124,N_9718);
nand U16191 (N_16191,N_12415,N_12472);
xnor U16192 (N_16192,N_11176,N_10150);
and U16193 (N_16193,N_6483,N_6868);
nand U16194 (N_16194,N_9966,N_11364);
and U16195 (N_16195,N_8651,N_8462);
xor U16196 (N_16196,N_8515,N_7398);
nor U16197 (N_16197,N_11750,N_7580);
and U16198 (N_16198,N_10900,N_6433);
nor U16199 (N_16199,N_7850,N_8879);
nor U16200 (N_16200,N_11250,N_6961);
and U16201 (N_16201,N_9067,N_12343);
nor U16202 (N_16202,N_7572,N_12163);
xor U16203 (N_16203,N_7380,N_7844);
and U16204 (N_16204,N_9000,N_11066);
and U16205 (N_16205,N_11872,N_7461);
or U16206 (N_16206,N_7608,N_11575);
xor U16207 (N_16207,N_6737,N_7021);
and U16208 (N_16208,N_9273,N_7098);
nor U16209 (N_16209,N_10790,N_11942);
nand U16210 (N_16210,N_9399,N_8632);
nand U16211 (N_16211,N_10608,N_11681);
nand U16212 (N_16212,N_11164,N_7818);
xor U16213 (N_16213,N_7939,N_11175);
or U16214 (N_16214,N_12335,N_8545);
and U16215 (N_16215,N_11928,N_7050);
nand U16216 (N_16216,N_7994,N_8290);
and U16217 (N_16217,N_10758,N_9428);
nand U16218 (N_16218,N_9565,N_11994);
xnor U16219 (N_16219,N_6434,N_8652);
xor U16220 (N_16220,N_11676,N_10095);
and U16221 (N_16221,N_12341,N_8060);
nor U16222 (N_16222,N_7582,N_8604);
or U16223 (N_16223,N_10972,N_8636);
nand U16224 (N_16224,N_12335,N_7698);
xnor U16225 (N_16225,N_9441,N_10102);
xor U16226 (N_16226,N_9253,N_10784);
nor U16227 (N_16227,N_9935,N_12262);
xor U16228 (N_16228,N_11961,N_8370);
or U16229 (N_16229,N_12338,N_6371);
or U16230 (N_16230,N_9450,N_8794);
nor U16231 (N_16231,N_10142,N_10009);
nor U16232 (N_16232,N_11375,N_8549);
xnor U16233 (N_16233,N_6889,N_10880);
nor U16234 (N_16234,N_6454,N_12267);
nand U16235 (N_16235,N_8967,N_6538);
or U16236 (N_16236,N_7597,N_8810);
or U16237 (N_16237,N_7045,N_6652);
xor U16238 (N_16238,N_8973,N_12077);
and U16239 (N_16239,N_7673,N_11468);
nor U16240 (N_16240,N_11543,N_6903);
nor U16241 (N_16241,N_7437,N_6254);
xnor U16242 (N_16242,N_9072,N_10550);
nor U16243 (N_16243,N_9689,N_9844);
xor U16244 (N_16244,N_7543,N_11197);
or U16245 (N_16245,N_7128,N_6544);
and U16246 (N_16246,N_11442,N_8031);
or U16247 (N_16247,N_12288,N_8322);
and U16248 (N_16248,N_6995,N_11338);
or U16249 (N_16249,N_11236,N_7332);
xnor U16250 (N_16250,N_12333,N_9929);
nand U16251 (N_16251,N_10634,N_11814);
and U16252 (N_16252,N_10286,N_11621);
nand U16253 (N_16253,N_11672,N_8689);
or U16254 (N_16254,N_12032,N_10183);
nand U16255 (N_16255,N_10082,N_9185);
or U16256 (N_16256,N_12213,N_8123);
xor U16257 (N_16257,N_12467,N_10375);
nand U16258 (N_16258,N_11805,N_10372);
or U16259 (N_16259,N_12172,N_8894);
nand U16260 (N_16260,N_12410,N_10284);
or U16261 (N_16261,N_9748,N_10254);
and U16262 (N_16262,N_8232,N_7174);
nand U16263 (N_16263,N_6751,N_8020);
xor U16264 (N_16264,N_11584,N_8957);
xor U16265 (N_16265,N_7971,N_10807);
xnor U16266 (N_16266,N_11381,N_11999);
nor U16267 (N_16267,N_6542,N_11614);
xor U16268 (N_16268,N_11680,N_11706);
or U16269 (N_16269,N_7071,N_7427);
and U16270 (N_16270,N_7869,N_6260);
xor U16271 (N_16271,N_9901,N_8779);
nor U16272 (N_16272,N_6280,N_8039);
or U16273 (N_16273,N_8495,N_7378);
xor U16274 (N_16274,N_10279,N_10337);
or U16275 (N_16275,N_10194,N_6679);
and U16276 (N_16276,N_6918,N_10905);
nand U16277 (N_16277,N_8783,N_10755);
nand U16278 (N_16278,N_6965,N_11102);
nand U16279 (N_16279,N_10692,N_7713);
and U16280 (N_16280,N_8083,N_7532);
nor U16281 (N_16281,N_9098,N_11022);
nor U16282 (N_16282,N_6601,N_7614);
or U16283 (N_16283,N_8675,N_9977);
nand U16284 (N_16284,N_12301,N_9124);
or U16285 (N_16285,N_10318,N_8965);
nor U16286 (N_16286,N_6376,N_12403);
nand U16287 (N_16287,N_11082,N_11107);
nand U16288 (N_16288,N_10579,N_11159);
nor U16289 (N_16289,N_12265,N_7483);
nand U16290 (N_16290,N_11084,N_9526);
xnor U16291 (N_16291,N_7464,N_12187);
and U16292 (N_16292,N_11997,N_7380);
nor U16293 (N_16293,N_6547,N_10844);
or U16294 (N_16294,N_8429,N_7609);
nor U16295 (N_16295,N_7573,N_10243);
nand U16296 (N_16296,N_8296,N_11468);
nand U16297 (N_16297,N_9918,N_10343);
and U16298 (N_16298,N_12277,N_9582);
nor U16299 (N_16299,N_7967,N_10553);
and U16300 (N_16300,N_7272,N_9608);
xnor U16301 (N_16301,N_8961,N_11100);
and U16302 (N_16302,N_11879,N_6953);
and U16303 (N_16303,N_8597,N_6474);
and U16304 (N_16304,N_8234,N_7763);
nor U16305 (N_16305,N_10471,N_11126);
nand U16306 (N_16306,N_11809,N_7094);
or U16307 (N_16307,N_9381,N_8513);
nand U16308 (N_16308,N_11493,N_11846);
and U16309 (N_16309,N_8851,N_10884);
nand U16310 (N_16310,N_9175,N_8352);
nand U16311 (N_16311,N_10150,N_8254);
nand U16312 (N_16312,N_9339,N_7042);
nor U16313 (N_16313,N_9607,N_9345);
xnor U16314 (N_16314,N_10314,N_7923);
xor U16315 (N_16315,N_8697,N_9548);
nand U16316 (N_16316,N_12497,N_8841);
xnor U16317 (N_16317,N_10941,N_8556);
nor U16318 (N_16318,N_11152,N_7158);
nor U16319 (N_16319,N_12377,N_10656);
xnor U16320 (N_16320,N_9672,N_6664);
nand U16321 (N_16321,N_8759,N_8686);
or U16322 (N_16322,N_8861,N_9258);
and U16323 (N_16323,N_8301,N_8718);
nor U16324 (N_16324,N_8982,N_12303);
xor U16325 (N_16325,N_8849,N_7249);
nand U16326 (N_16326,N_8784,N_7031);
xnor U16327 (N_16327,N_11150,N_6525);
or U16328 (N_16328,N_11895,N_8850);
and U16329 (N_16329,N_12228,N_11212);
xor U16330 (N_16330,N_11032,N_12117);
xor U16331 (N_16331,N_7270,N_7723);
nor U16332 (N_16332,N_6293,N_10994);
or U16333 (N_16333,N_11293,N_9540);
and U16334 (N_16334,N_7237,N_9074);
nor U16335 (N_16335,N_11903,N_11064);
nand U16336 (N_16336,N_7342,N_9569);
xnor U16337 (N_16337,N_7461,N_12088);
xnor U16338 (N_16338,N_11638,N_11076);
or U16339 (N_16339,N_10454,N_10693);
or U16340 (N_16340,N_8586,N_7692);
and U16341 (N_16341,N_11422,N_8243);
or U16342 (N_16342,N_6628,N_12306);
xnor U16343 (N_16343,N_11666,N_11328);
nor U16344 (N_16344,N_8270,N_9561);
and U16345 (N_16345,N_7060,N_7466);
or U16346 (N_16346,N_9066,N_9827);
nand U16347 (N_16347,N_10843,N_8394);
xnor U16348 (N_16348,N_12073,N_7545);
nand U16349 (N_16349,N_12058,N_8414);
nand U16350 (N_16350,N_10842,N_8835);
or U16351 (N_16351,N_11520,N_11249);
xor U16352 (N_16352,N_9566,N_6448);
and U16353 (N_16353,N_6402,N_11462);
nand U16354 (N_16354,N_12222,N_12103);
or U16355 (N_16355,N_9342,N_9286);
xnor U16356 (N_16356,N_7871,N_11308);
or U16357 (N_16357,N_9038,N_10360);
nor U16358 (N_16358,N_9967,N_7458);
and U16359 (N_16359,N_8430,N_7209);
xor U16360 (N_16360,N_8140,N_10267);
or U16361 (N_16361,N_8581,N_9800);
nor U16362 (N_16362,N_8518,N_9099);
or U16363 (N_16363,N_10726,N_10962);
xor U16364 (N_16364,N_8110,N_7388);
or U16365 (N_16365,N_8639,N_10552);
nor U16366 (N_16366,N_8780,N_9037);
nand U16367 (N_16367,N_8807,N_9525);
nand U16368 (N_16368,N_7183,N_8045);
xor U16369 (N_16369,N_9402,N_7081);
nor U16370 (N_16370,N_7153,N_10684);
and U16371 (N_16371,N_6851,N_11529);
nand U16372 (N_16372,N_8483,N_7742);
or U16373 (N_16373,N_10418,N_10298);
nand U16374 (N_16374,N_7907,N_9043);
xnor U16375 (N_16375,N_11610,N_10260);
and U16376 (N_16376,N_8155,N_6697);
nand U16377 (N_16377,N_11441,N_10364);
xor U16378 (N_16378,N_7506,N_12279);
nor U16379 (N_16379,N_11543,N_11620);
xor U16380 (N_16380,N_7816,N_10713);
xnor U16381 (N_16381,N_10607,N_8931);
or U16382 (N_16382,N_11073,N_10281);
nor U16383 (N_16383,N_10187,N_8017);
or U16384 (N_16384,N_8564,N_8328);
nor U16385 (N_16385,N_8278,N_11149);
or U16386 (N_16386,N_11883,N_12163);
nand U16387 (N_16387,N_7696,N_7687);
nand U16388 (N_16388,N_10263,N_10022);
nand U16389 (N_16389,N_7315,N_7194);
nor U16390 (N_16390,N_8450,N_11140);
and U16391 (N_16391,N_11699,N_8139);
xor U16392 (N_16392,N_8990,N_9789);
and U16393 (N_16393,N_11507,N_7827);
or U16394 (N_16394,N_9138,N_8914);
xor U16395 (N_16395,N_9669,N_6778);
and U16396 (N_16396,N_7217,N_8422);
nand U16397 (N_16397,N_8955,N_7397);
nor U16398 (N_16398,N_8152,N_8131);
and U16399 (N_16399,N_9277,N_8412);
nand U16400 (N_16400,N_7521,N_9921);
or U16401 (N_16401,N_8125,N_8370);
xnor U16402 (N_16402,N_11352,N_9370);
xor U16403 (N_16403,N_10115,N_10988);
xnor U16404 (N_16404,N_9702,N_12357);
and U16405 (N_16405,N_7037,N_10479);
nand U16406 (N_16406,N_11275,N_9607);
nand U16407 (N_16407,N_7769,N_10809);
nor U16408 (N_16408,N_9594,N_6756);
nand U16409 (N_16409,N_11093,N_10020);
nor U16410 (N_16410,N_12126,N_11057);
and U16411 (N_16411,N_8679,N_8835);
or U16412 (N_16412,N_11906,N_10452);
xnor U16413 (N_16413,N_8156,N_9682);
and U16414 (N_16414,N_8880,N_8134);
nor U16415 (N_16415,N_7181,N_8543);
xnor U16416 (N_16416,N_7585,N_12164);
xnor U16417 (N_16417,N_6876,N_8565);
and U16418 (N_16418,N_11823,N_12438);
xor U16419 (N_16419,N_8220,N_8649);
or U16420 (N_16420,N_11467,N_7315);
or U16421 (N_16421,N_10501,N_12101);
or U16422 (N_16422,N_7692,N_7682);
xor U16423 (N_16423,N_12139,N_7863);
nand U16424 (N_16424,N_10366,N_9082);
nor U16425 (N_16425,N_9997,N_9537);
nor U16426 (N_16426,N_11176,N_11184);
and U16427 (N_16427,N_8437,N_10430);
or U16428 (N_16428,N_12149,N_11882);
and U16429 (N_16429,N_12234,N_8814);
nor U16430 (N_16430,N_10014,N_10458);
and U16431 (N_16431,N_7199,N_12341);
nand U16432 (N_16432,N_11799,N_12383);
nor U16433 (N_16433,N_6669,N_8193);
xor U16434 (N_16434,N_9007,N_9251);
and U16435 (N_16435,N_8148,N_8524);
nand U16436 (N_16436,N_11619,N_8199);
xnor U16437 (N_16437,N_7023,N_11497);
or U16438 (N_16438,N_8011,N_9120);
xnor U16439 (N_16439,N_7665,N_12209);
or U16440 (N_16440,N_11550,N_11900);
or U16441 (N_16441,N_10637,N_12429);
or U16442 (N_16442,N_11595,N_12346);
or U16443 (N_16443,N_9253,N_6855);
nor U16444 (N_16444,N_7054,N_7604);
xnor U16445 (N_16445,N_6470,N_7023);
nor U16446 (N_16446,N_11608,N_9380);
or U16447 (N_16447,N_10926,N_12350);
and U16448 (N_16448,N_7141,N_9109);
and U16449 (N_16449,N_10954,N_6280);
or U16450 (N_16450,N_12401,N_8574);
or U16451 (N_16451,N_8586,N_6751);
nand U16452 (N_16452,N_11105,N_10198);
xor U16453 (N_16453,N_11390,N_8322);
and U16454 (N_16454,N_10352,N_8478);
or U16455 (N_16455,N_9986,N_10848);
nand U16456 (N_16456,N_9886,N_11400);
or U16457 (N_16457,N_10279,N_9770);
nor U16458 (N_16458,N_10171,N_11940);
nor U16459 (N_16459,N_9600,N_9449);
nand U16460 (N_16460,N_6644,N_8193);
or U16461 (N_16461,N_7567,N_8648);
nand U16462 (N_16462,N_7886,N_9309);
xnor U16463 (N_16463,N_7258,N_7355);
nor U16464 (N_16464,N_10346,N_9261);
nor U16465 (N_16465,N_10820,N_9023);
nor U16466 (N_16466,N_8223,N_10413);
xor U16467 (N_16467,N_6361,N_8058);
xor U16468 (N_16468,N_9112,N_6410);
nor U16469 (N_16469,N_9582,N_11350);
or U16470 (N_16470,N_7477,N_10051);
or U16471 (N_16471,N_10607,N_7206);
xor U16472 (N_16472,N_7380,N_7178);
and U16473 (N_16473,N_11104,N_8273);
nor U16474 (N_16474,N_8638,N_10652);
xor U16475 (N_16475,N_10201,N_7241);
nor U16476 (N_16476,N_11234,N_11562);
and U16477 (N_16477,N_7685,N_9849);
or U16478 (N_16478,N_11619,N_9029);
and U16479 (N_16479,N_6554,N_10932);
nor U16480 (N_16480,N_7195,N_8558);
nor U16481 (N_16481,N_11371,N_11184);
nand U16482 (N_16482,N_10960,N_10861);
or U16483 (N_16483,N_12222,N_11184);
xnor U16484 (N_16484,N_6861,N_8942);
or U16485 (N_16485,N_12208,N_11371);
and U16486 (N_16486,N_9745,N_7215);
xor U16487 (N_16487,N_11698,N_7727);
nor U16488 (N_16488,N_7478,N_8966);
and U16489 (N_16489,N_10997,N_7013);
xor U16490 (N_16490,N_7218,N_8402);
or U16491 (N_16491,N_12005,N_7520);
nor U16492 (N_16492,N_9798,N_7634);
or U16493 (N_16493,N_8868,N_9758);
and U16494 (N_16494,N_6400,N_8683);
nor U16495 (N_16495,N_9967,N_10868);
and U16496 (N_16496,N_9573,N_9670);
or U16497 (N_16497,N_10363,N_9873);
nor U16498 (N_16498,N_6303,N_9885);
and U16499 (N_16499,N_10884,N_6959);
and U16500 (N_16500,N_9929,N_8260);
xnor U16501 (N_16501,N_6576,N_6461);
and U16502 (N_16502,N_12243,N_7572);
nand U16503 (N_16503,N_11600,N_11480);
and U16504 (N_16504,N_6403,N_6412);
or U16505 (N_16505,N_11504,N_10813);
or U16506 (N_16506,N_9407,N_7943);
nor U16507 (N_16507,N_11575,N_7006);
and U16508 (N_16508,N_10436,N_8881);
nor U16509 (N_16509,N_10531,N_11455);
xor U16510 (N_16510,N_7378,N_7052);
nand U16511 (N_16511,N_8759,N_11867);
and U16512 (N_16512,N_6651,N_9418);
nor U16513 (N_16513,N_11693,N_10229);
nand U16514 (N_16514,N_12385,N_11528);
or U16515 (N_16515,N_8754,N_10360);
nand U16516 (N_16516,N_8538,N_9668);
nor U16517 (N_16517,N_10724,N_11350);
or U16518 (N_16518,N_10501,N_6950);
and U16519 (N_16519,N_7860,N_9169);
and U16520 (N_16520,N_10085,N_9954);
xnor U16521 (N_16521,N_8605,N_6413);
nand U16522 (N_16522,N_11156,N_9112);
nor U16523 (N_16523,N_8510,N_8826);
nor U16524 (N_16524,N_9746,N_10162);
nor U16525 (N_16525,N_7179,N_8566);
and U16526 (N_16526,N_9560,N_9005);
nor U16527 (N_16527,N_7491,N_9334);
nand U16528 (N_16528,N_7954,N_11188);
nor U16529 (N_16529,N_8591,N_12136);
xnor U16530 (N_16530,N_9535,N_6396);
nor U16531 (N_16531,N_9923,N_7354);
and U16532 (N_16532,N_9448,N_12119);
or U16533 (N_16533,N_11593,N_10682);
xnor U16534 (N_16534,N_9046,N_7745);
or U16535 (N_16535,N_10273,N_8610);
or U16536 (N_16536,N_8055,N_9373);
nor U16537 (N_16537,N_11662,N_9974);
and U16538 (N_16538,N_12024,N_9479);
or U16539 (N_16539,N_10037,N_12247);
or U16540 (N_16540,N_7971,N_8558);
xor U16541 (N_16541,N_7662,N_11531);
nor U16542 (N_16542,N_7595,N_7030);
nand U16543 (N_16543,N_11918,N_9110);
nor U16544 (N_16544,N_10084,N_8393);
nand U16545 (N_16545,N_7283,N_6634);
and U16546 (N_16546,N_7352,N_10183);
xor U16547 (N_16547,N_10095,N_8262);
xor U16548 (N_16548,N_10193,N_8225);
xnor U16549 (N_16549,N_6903,N_10747);
nand U16550 (N_16550,N_10958,N_8583);
or U16551 (N_16551,N_10671,N_6568);
and U16552 (N_16552,N_9529,N_6952);
xnor U16553 (N_16553,N_12411,N_9323);
and U16554 (N_16554,N_11205,N_6273);
nand U16555 (N_16555,N_11927,N_12276);
or U16556 (N_16556,N_8756,N_7659);
nand U16557 (N_16557,N_9356,N_9320);
nand U16558 (N_16558,N_8908,N_10730);
xnor U16559 (N_16559,N_12218,N_10590);
xnor U16560 (N_16560,N_10029,N_7093);
or U16561 (N_16561,N_10320,N_10637);
or U16562 (N_16562,N_7915,N_12146);
nand U16563 (N_16563,N_10575,N_10704);
nor U16564 (N_16564,N_8467,N_7271);
nor U16565 (N_16565,N_8532,N_9305);
and U16566 (N_16566,N_7187,N_11489);
nor U16567 (N_16567,N_10985,N_9945);
nor U16568 (N_16568,N_6701,N_7765);
nand U16569 (N_16569,N_10244,N_11390);
nand U16570 (N_16570,N_11138,N_8487);
nor U16571 (N_16571,N_6372,N_8830);
and U16572 (N_16572,N_9124,N_7438);
and U16573 (N_16573,N_6283,N_11719);
nand U16574 (N_16574,N_6959,N_12224);
or U16575 (N_16575,N_9411,N_11372);
or U16576 (N_16576,N_9090,N_7862);
or U16577 (N_16577,N_6811,N_11377);
nor U16578 (N_16578,N_7252,N_10316);
nand U16579 (N_16579,N_12024,N_11913);
nor U16580 (N_16580,N_10997,N_11871);
or U16581 (N_16581,N_9853,N_10886);
nor U16582 (N_16582,N_8769,N_6439);
nand U16583 (N_16583,N_11794,N_12238);
or U16584 (N_16584,N_6391,N_9881);
xnor U16585 (N_16585,N_11110,N_8404);
or U16586 (N_16586,N_10407,N_9510);
and U16587 (N_16587,N_11508,N_11700);
nor U16588 (N_16588,N_8593,N_10160);
xnor U16589 (N_16589,N_8377,N_10705);
xnor U16590 (N_16590,N_11980,N_10593);
nor U16591 (N_16591,N_9449,N_10266);
or U16592 (N_16592,N_10066,N_8268);
xnor U16593 (N_16593,N_7324,N_6907);
xor U16594 (N_16594,N_11834,N_7373);
or U16595 (N_16595,N_7265,N_11349);
xnor U16596 (N_16596,N_11678,N_10116);
xor U16597 (N_16597,N_7004,N_11756);
and U16598 (N_16598,N_7786,N_10970);
nor U16599 (N_16599,N_6588,N_10856);
nor U16600 (N_16600,N_6438,N_8372);
nand U16601 (N_16601,N_12362,N_9595);
or U16602 (N_16602,N_9598,N_8418);
nor U16603 (N_16603,N_8568,N_6931);
nor U16604 (N_16604,N_6606,N_9797);
nor U16605 (N_16605,N_9926,N_7194);
nand U16606 (N_16606,N_8982,N_7316);
nor U16607 (N_16607,N_11227,N_10276);
xnor U16608 (N_16608,N_9724,N_6482);
or U16609 (N_16609,N_9981,N_10239);
nand U16610 (N_16610,N_7050,N_12005);
or U16611 (N_16611,N_8391,N_7736);
nand U16612 (N_16612,N_6621,N_11391);
nor U16613 (N_16613,N_11442,N_7880);
and U16614 (N_16614,N_7084,N_9960);
and U16615 (N_16615,N_8705,N_7691);
or U16616 (N_16616,N_9675,N_8043);
nand U16617 (N_16617,N_8329,N_6857);
nand U16618 (N_16618,N_8187,N_8010);
or U16619 (N_16619,N_11022,N_8573);
nor U16620 (N_16620,N_12014,N_9147);
or U16621 (N_16621,N_12248,N_7978);
nand U16622 (N_16622,N_11724,N_9733);
xor U16623 (N_16623,N_10462,N_8789);
nor U16624 (N_16624,N_9881,N_10229);
nand U16625 (N_16625,N_9015,N_9101);
nand U16626 (N_16626,N_7917,N_10801);
and U16627 (N_16627,N_11364,N_6960);
nor U16628 (N_16628,N_8133,N_9216);
and U16629 (N_16629,N_8215,N_9013);
nor U16630 (N_16630,N_9412,N_9339);
or U16631 (N_16631,N_7088,N_7782);
nand U16632 (N_16632,N_10497,N_7766);
nor U16633 (N_16633,N_7144,N_9283);
nor U16634 (N_16634,N_6705,N_12181);
nand U16635 (N_16635,N_9617,N_11247);
nand U16636 (N_16636,N_11684,N_9250);
xor U16637 (N_16637,N_10667,N_6688);
or U16638 (N_16638,N_8993,N_9541);
nand U16639 (N_16639,N_11882,N_12250);
nor U16640 (N_16640,N_8755,N_6911);
xor U16641 (N_16641,N_12496,N_12353);
nand U16642 (N_16642,N_10521,N_11462);
nand U16643 (N_16643,N_8018,N_9541);
nand U16644 (N_16644,N_10207,N_11680);
nand U16645 (N_16645,N_12029,N_12196);
nand U16646 (N_16646,N_8551,N_6274);
or U16647 (N_16647,N_8329,N_11655);
xnor U16648 (N_16648,N_8303,N_7639);
nor U16649 (N_16649,N_11859,N_10478);
or U16650 (N_16650,N_7192,N_6669);
or U16651 (N_16651,N_11132,N_7912);
and U16652 (N_16652,N_10234,N_8884);
or U16653 (N_16653,N_8198,N_10587);
xor U16654 (N_16654,N_9528,N_12319);
nand U16655 (N_16655,N_6781,N_12392);
or U16656 (N_16656,N_11346,N_10811);
nor U16657 (N_16657,N_11120,N_9675);
nor U16658 (N_16658,N_7955,N_8623);
xor U16659 (N_16659,N_7480,N_6505);
and U16660 (N_16660,N_7443,N_8578);
or U16661 (N_16661,N_10780,N_7097);
xnor U16662 (N_16662,N_7533,N_7281);
nor U16663 (N_16663,N_11500,N_10304);
nand U16664 (N_16664,N_10531,N_8932);
nand U16665 (N_16665,N_11348,N_11483);
and U16666 (N_16666,N_9867,N_11541);
and U16667 (N_16667,N_10903,N_11287);
nand U16668 (N_16668,N_9970,N_10758);
nor U16669 (N_16669,N_9448,N_9753);
nor U16670 (N_16670,N_10940,N_10212);
xnor U16671 (N_16671,N_7710,N_7242);
nand U16672 (N_16672,N_10250,N_8729);
xnor U16673 (N_16673,N_8492,N_7998);
nand U16674 (N_16674,N_7758,N_11856);
nor U16675 (N_16675,N_11639,N_8121);
xor U16676 (N_16676,N_7635,N_6513);
xnor U16677 (N_16677,N_9609,N_8187);
nor U16678 (N_16678,N_11839,N_6656);
nand U16679 (N_16679,N_11824,N_7988);
nor U16680 (N_16680,N_7202,N_7272);
and U16681 (N_16681,N_10770,N_11239);
nand U16682 (N_16682,N_11600,N_9610);
or U16683 (N_16683,N_6929,N_6902);
or U16684 (N_16684,N_7023,N_11351);
nand U16685 (N_16685,N_7322,N_8288);
xor U16686 (N_16686,N_9041,N_10462);
or U16687 (N_16687,N_9198,N_8119);
or U16688 (N_16688,N_9941,N_8090);
nand U16689 (N_16689,N_11358,N_8744);
xnor U16690 (N_16690,N_8442,N_12389);
xnor U16691 (N_16691,N_9089,N_7835);
or U16692 (N_16692,N_10794,N_9797);
xor U16693 (N_16693,N_9919,N_7016);
and U16694 (N_16694,N_8858,N_10890);
nand U16695 (N_16695,N_11073,N_7688);
and U16696 (N_16696,N_7371,N_9800);
nor U16697 (N_16697,N_11841,N_12203);
nand U16698 (N_16698,N_12392,N_7945);
or U16699 (N_16699,N_12027,N_8474);
or U16700 (N_16700,N_9766,N_6781);
or U16701 (N_16701,N_6947,N_7038);
and U16702 (N_16702,N_11758,N_12174);
and U16703 (N_16703,N_10462,N_9115);
nor U16704 (N_16704,N_8507,N_12444);
and U16705 (N_16705,N_11362,N_7191);
and U16706 (N_16706,N_6511,N_12369);
and U16707 (N_16707,N_6816,N_7572);
xor U16708 (N_16708,N_10615,N_11107);
and U16709 (N_16709,N_11247,N_11777);
xor U16710 (N_16710,N_10876,N_6954);
or U16711 (N_16711,N_6819,N_9808);
and U16712 (N_16712,N_12248,N_11420);
nor U16713 (N_16713,N_6582,N_6435);
nand U16714 (N_16714,N_10289,N_12484);
nand U16715 (N_16715,N_8430,N_11286);
nand U16716 (N_16716,N_8850,N_8978);
and U16717 (N_16717,N_11717,N_8639);
nand U16718 (N_16718,N_9785,N_7431);
xnor U16719 (N_16719,N_11253,N_10416);
nor U16720 (N_16720,N_11816,N_7112);
xor U16721 (N_16721,N_7593,N_9742);
or U16722 (N_16722,N_10126,N_10786);
nand U16723 (N_16723,N_7411,N_10286);
nor U16724 (N_16724,N_8525,N_9593);
nand U16725 (N_16725,N_8884,N_12043);
xnor U16726 (N_16726,N_9148,N_10621);
nand U16727 (N_16727,N_11285,N_12092);
nor U16728 (N_16728,N_9264,N_8699);
and U16729 (N_16729,N_7364,N_9337);
or U16730 (N_16730,N_12292,N_12050);
nand U16731 (N_16731,N_9420,N_7254);
or U16732 (N_16732,N_10681,N_9242);
nand U16733 (N_16733,N_11152,N_9982);
or U16734 (N_16734,N_6884,N_7671);
nand U16735 (N_16735,N_6940,N_7799);
nor U16736 (N_16736,N_11466,N_11025);
or U16737 (N_16737,N_10047,N_10578);
xnor U16738 (N_16738,N_6596,N_11775);
nor U16739 (N_16739,N_8939,N_6661);
xor U16740 (N_16740,N_6468,N_12012);
and U16741 (N_16741,N_11095,N_8333);
and U16742 (N_16742,N_7562,N_8358);
nand U16743 (N_16743,N_10240,N_7639);
xor U16744 (N_16744,N_11950,N_10177);
and U16745 (N_16745,N_8112,N_10028);
or U16746 (N_16746,N_8069,N_10694);
nor U16747 (N_16747,N_11913,N_10472);
or U16748 (N_16748,N_11331,N_7029);
and U16749 (N_16749,N_11271,N_8633);
nand U16750 (N_16750,N_8471,N_9097);
xor U16751 (N_16751,N_12244,N_10523);
nor U16752 (N_16752,N_6851,N_11690);
nor U16753 (N_16753,N_9828,N_6587);
xor U16754 (N_16754,N_11491,N_11947);
xor U16755 (N_16755,N_7921,N_11773);
and U16756 (N_16756,N_11062,N_11315);
nand U16757 (N_16757,N_8324,N_7546);
nor U16758 (N_16758,N_8992,N_11999);
and U16759 (N_16759,N_9476,N_8196);
xor U16760 (N_16760,N_6394,N_8037);
xnor U16761 (N_16761,N_8673,N_6514);
nand U16762 (N_16762,N_12375,N_7194);
nand U16763 (N_16763,N_11054,N_6746);
nand U16764 (N_16764,N_10338,N_7576);
or U16765 (N_16765,N_9792,N_11720);
nand U16766 (N_16766,N_6962,N_10362);
or U16767 (N_16767,N_10089,N_11544);
and U16768 (N_16768,N_11368,N_11822);
or U16769 (N_16769,N_9332,N_8902);
or U16770 (N_16770,N_8986,N_7971);
nor U16771 (N_16771,N_8335,N_11758);
or U16772 (N_16772,N_7139,N_7291);
and U16773 (N_16773,N_9173,N_8022);
nand U16774 (N_16774,N_11490,N_11215);
xnor U16775 (N_16775,N_10303,N_7877);
and U16776 (N_16776,N_9972,N_9475);
and U16777 (N_16777,N_8643,N_12201);
nand U16778 (N_16778,N_6736,N_9647);
or U16779 (N_16779,N_9116,N_7827);
and U16780 (N_16780,N_9712,N_11276);
and U16781 (N_16781,N_11506,N_6854);
xor U16782 (N_16782,N_8893,N_11379);
xnor U16783 (N_16783,N_9656,N_8095);
or U16784 (N_16784,N_8808,N_12447);
nand U16785 (N_16785,N_12329,N_11734);
nand U16786 (N_16786,N_9651,N_11701);
or U16787 (N_16787,N_11162,N_6492);
nor U16788 (N_16788,N_9937,N_10066);
xnor U16789 (N_16789,N_7476,N_11861);
nor U16790 (N_16790,N_7040,N_7510);
and U16791 (N_16791,N_10005,N_11865);
and U16792 (N_16792,N_8639,N_11900);
xor U16793 (N_16793,N_7139,N_6412);
nand U16794 (N_16794,N_10051,N_6821);
xor U16795 (N_16795,N_11070,N_6334);
and U16796 (N_16796,N_10030,N_6494);
nor U16797 (N_16797,N_8141,N_9525);
and U16798 (N_16798,N_9177,N_11761);
or U16799 (N_16799,N_10660,N_6278);
xor U16800 (N_16800,N_10230,N_8348);
nand U16801 (N_16801,N_11903,N_9791);
nor U16802 (N_16802,N_7604,N_11030);
nand U16803 (N_16803,N_11501,N_9419);
or U16804 (N_16804,N_11930,N_11385);
nand U16805 (N_16805,N_6279,N_11082);
nand U16806 (N_16806,N_8284,N_8409);
nor U16807 (N_16807,N_11899,N_12478);
nand U16808 (N_16808,N_11899,N_6678);
and U16809 (N_16809,N_8802,N_11470);
nor U16810 (N_16810,N_8850,N_9490);
and U16811 (N_16811,N_10432,N_10346);
xnor U16812 (N_16812,N_10408,N_10831);
nand U16813 (N_16813,N_11853,N_8921);
and U16814 (N_16814,N_10493,N_7565);
nor U16815 (N_16815,N_9624,N_11144);
and U16816 (N_16816,N_6978,N_10474);
xor U16817 (N_16817,N_9633,N_9027);
nor U16818 (N_16818,N_9350,N_11156);
and U16819 (N_16819,N_7740,N_7507);
or U16820 (N_16820,N_10085,N_7240);
nor U16821 (N_16821,N_7030,N_10181);
or U16822 (N_16822,N_6514,N_9199);
nor U16823 (N_16823,N_8954,N_11848);
and U16824 (N_16824,N_6390,N_8456);
nand U16825 (N_16825,N_8046,N_7584);
xor U16826 (N_16826,N_9955,N_10138);
and U16827 (N_16827,N_6434,N_9907);
nor U16828 (N_16828,N_11574,N_6524);
nor U16829 (N_16829,N_10870,N_6741);
xor U16830 (N_16830,N_12234,N_8944);
xnor U16831 (N_16831,N_6251,N_8098);
and U16832 (N_16832,N_6874,N_9648);
or U16833 (N_16833,N_6724,N_8556);
and U16834 (N_16834,N_10937,N_12033);
nor U16835 (N_16835,N_10541,N_8182);
nor U16836 (N_16836,N_10747,N_8322);
or U16837 (N_16837,N_11120,N_11017);
or U16838 (N_16838,N_9981,N_12315);
nand U16839 (N_16839,N_11532,N_10752);
nand U16840 (N_16840,N_9392,N_7760);
xor U16841 (N_16841,N_6825,N_11152);
and U16842 (N_16842,N_11862,N_6786);
nor U16843 (N_16843,N_8766,N_12160);
or U16844 (N_16844,N_11067,N_12435);
xnor U16845 (N_16845,N_11689,N_11040);
and U16846 (N_16846,N_12458,N_8220);
nand U16847 (N_16847,N_7340,N_7760);
nor U16848 (N_16848,N_7255,N_8360);
nor U16849 (N_16849,N_9297,N_10935);
nand U16850 (N_16850,N_8061,N_12215);
or U16851 (N_16851,N_10539,N_6299);
and U16852 (N_16852,N_7590,N_9107);
or U16853 (N_16853,N_10770,N_8732);
nor U16854 (N_16854,N_7850,N_9849);
or U16855 (N_16855,N_7446,N_6692);
or U16856 (N_16856,N_8355,N_6358);
nand U16857 (N_16857,N_11930,N_6546);
and U16858 (N_16858,N_8750,N_6531);
and U16859 (N_16859,N_12039,N_6862);
and U16860 (N_16860,N_11784,N_11873);
nor U16861 (N_16861,N_6309,N_11452);
nand U16862 (N_16862,N_6562,N_11799);
and U16863 (N_16863,N_8122,N_10584);
and U16864 (N_16864,N_9698,N_9520);
xnor U16865 (N_16865,N_12400,N_10309);
nor U16866 (N_16866,N_7051,N_12204);
nor U16867 (N_16867,N_10615,N_9451);
xnor U16868 (N_16868,N_9167,N_10021);
or U16869 (N_16869,N_7792,N_10336);
nand U16870 (N_16870,N_8956,N_12411);
and U16871 (N_16871,N_8674,N_9548);
nand U16872 (N_16872,N_9190,N_10046);
or U16873 (N_16873,N_8641,N_10550);
nor U16874 (N_16874,N_8254,N_7777);
or U16875 (N_16875,N_11666,N_9536);
xnor U16876 (N_16876,N_8254,N_11152);
xor U16877 (N_16877,N_6978,N_11659);
and U16878 (N_16878,N_10973,N_6393);
or U16879 (N_16879,N_6615,N_7143);
and U16880 (N_16880,N_10367,N_11383);
and U16881 (N_16881,N_7765,N_7638);
and U16882 (N_16882,N_10719,N_10346);
nand U16883 (N_16883,N_8640,N_11719);
and U16884 (N_16884,N_9896,N_9403);
and U16885 (N_16885,N_11563,N_6417);
or U16886 (N_16886,N_8731,N_12430);
xnor U16887 (N_16887,N_9824,N_12135);
nand U16888 (N_16888,N_11207,N_8390);
and U16889 (N_16889,N_9064,N_7903);
nand U16890 (N_16890,N_6923,N_7407);
nor U16891 (N_16891,N_9902,N_6539);
xor U16892 (N_16892,N_6424,N_7787);
nor U16893 (N_16893,N_11469,N_8450);
or U16894 (N_16894,N_8980,N_8235);
nand U16895 (N_16895,N_8714,N_12385);
and U16896 (N_16896,N_8748,N_6912);
xor U16897 (N_16897,N_8498,N_11844);
or U16898 (N_16898,N_10569,N_10923);
xor U16899 (N_16899,N_7397,N_6957);
or U16900 (N_16900,N_7150,N_10322);
and U16901 (N_16901,N_9134,N_6922);
or U16902 (N_16902,N_8536,N_10142);
xnor U16903 (N_16903,N_10678,N_6520);
nor U16904 (N_16904,N_10847,N_10013);
or U16905 (N_16905,N_9812,N_7416);
xnor U16906 (N_16906,N_11937,N_9749);
nor U16907 (N_16907,N_8759,N_7462);
nand U16908 (N_16908,N_11178,N_7030);
nor U16909 (N_16909,N_9614,N_9983);
and U16910 (N_16910,N_9579,N_10848);
or U16911 (N_16911,N_8678,N_7977);
and U16912 (N_16912,N_10544,N_12024);
and U16913 (N_16913,N_6251,N_10233);
and U16914 (N_16914,N_12072,N_10875);
nand U16915 (N_16915,N_9642,N_7685);
and U16916 (N_16916,N_10855,N_6755);
xnor U16917 (N_16917,N_7077,N_10578);
xnor U16918 (N_16918,N_10808,N_9720);
or U16919 (N_16919,N_12153,N_12279);
and U16920 (N_16920,N_7199,N_7935);
nor U16921 (N_16921,N_11197,N_11732);
nor U16922 (N_16922,N_11935,N_10480);
nand U16923 (N_16923,N_7957,N_10741);
nand U16924 (N_16924,N_11630,N_8303);
xnor U16925 (N_16925,N_11817,N_9333);
nand U16926 (N_16926,N_7752,N_8830);
or U16927 (N_16927,N_12462,N_6990);
nand U16928 (N_16928,N_10148,N_7858);
or U16929 (N_16929,N_6865,N_7808);
nor U16930 (N_16930,N_10846,N_8523);
and U16931 (N_16931,N_11520,N_6291);
nand U16932 (N_16932,N_6826,N_9719);
nor U16933 (N_16933,N_9887,N_7873);
nand U16934 (N_16934,N_6693,N_8235);
or U16935 (N_16935,N_10819,N_10442);
xor U16936 (N_16936,N_10543,N_6363);
and U16937 (N_16937,N_6796,N_6511);
nand U16938 (N_16938,N_9323,N_9614);
nand U16939 (N_16939,N_6490,N_9698);
or U16940 (N_16940,N_10612,N_11521);
and U16941 (N_16941,N_6364,N_6904);
nand U16942 (N_16942,N_7688,N_10191);
and U16943 (N_16943,N_9753,N_11568);
and U16944 (N_16944,N_12049,N_9667);
xor U16945 (N_16945,N_10379,N_7483);
and U16946 (N_16946,N_7625,N_8003);
nand U16947 (N_16947,N_11180,N_11081);
or U16948 (N_16948,N_8687,N_11531);
nand U16949 (N_16949,N_11167,N_9631);
nand U16950 (N_16950,N_12165,N_12364);
nor U16951 (N_16951,N_8026,N_11637);
and U16952 (N_16952,N_8044,N_12112);
or U16953 (N_16953,N_7766,N_9766);
nor U16954 (N_16954,N_9227,N_7617);
nand U16955 (N_16955,N_8924,N_10574);
nand U16956 (N_16956,N_10852,N_9627);
nand U16957 (N_16957,N_8186,N_12347);
or U16958 (N_16958,N_11619,N_6866);
or U16959 (N_16959,N_9202,N_10347);
or U16960 (N_16960,N_6272,N_7547);
nand U16961 (N_16961,N_9791,N_10146);
and U16962 (N_16962,N_6365,N_12075);
nor U16963 (N_16963,N_6325,N_7532);
and U16964 (N_16964,N_7310,N_7175);
xnor U16965 (N_16965,N_8212,N_11090);
xnor U16966 (N_16966,N_8345,N_10862);
and U16967 (N_16967,N_12489,N_11526);
nor U16968 (N_16968,N_6401,N_11038);
and U16969 (N_16969,N_9799,N_12427);
nand U16970 (N_16970,N_8324,N_6957);
nand U16971 (N_16971,N_9838,N_11351);
xnor U16972 (N_16972,N_11741,N_10528);
and U16973 (N_16973,N_9490,N_8848);
nor U16974 (N_16974,N_11721,N_9335);
xor U16975 (N_16975,N_9719,N_11079);
or U16976 (N_16976,N_8546,N_9627);
nand U16977 (N_16977,N_12029,N_7863);
nand U16978 (N_16978,N_8576,N_6940);
or U16979 (N_16979,N_6840,N_7787);
or U16980 (N_16980,N_11482,N_7216);
and U16981 (N_16981,N_6443,N_7637);
nor U16982 (N_16982,N_9872,N_9754);
nor U16983 (N_16983,N_6822,N_7074);
nand U16984 (N_16984,N_9855,N_10981);
nand U16985 (N_16985,N_9579,N_7851);
xnor U16986 (N_16986,N_6381,N_7525);
xnor U16987 (N_16987,N_9095,N_9594);
or U16988 (N_16988,N_9009,N_6655);
nor U16989 (N_16989,N_10131,N_10085);
or U16990 (N_16990,N_10124,N_6574);
nor U16991 (N_16991,N_11759,N_10759);
and U16992 (N_16992,N_9225,N_6525);
or U16993 (N_16993,N_10684,N_11049);
and U16994 (N_16994,N_7402,N_6424);
nor U16995 (N_16995,N_9443,N_7333);
nor U16996 (N_16996,N_11974,N_6352);
nor U16997 (N_16997,N_9313,N_8119);
nor U16998 (N_16998,N_8164,N_10137);
nand U16999 (N_16999,N_6832,N_7412);
or U17000 (N_17000,N_7616,N_7471);
or U17001 (N_17001,N_8384,N_7252);
and U17002 (N_17002,N_10978,N_10734);
nand U17003 (N_17003,N_6434,N_9881);
or U17004 (N_17004,N_9429,N_8493);
nor U17005 (N_17005,N_8747,N_8200);
and U17006 (N_17006,N_7195,N_9876);
xnor U17007 (N_17007,N_8929,N_6891);
nor U17008 (N_17008,N_12482,N_6704);
xor U17009 (N_17009,N_8232,N_11862);
and U17010 (N_17010,N_9819,N_8390);
or U17011 (N_17011,N_6275,N_9891);
or U17012 (N_17012,N_11612,N_7892);
nand U17013 (N_17013,N_7657,N_9761);
nor U17014 (N_17014,N_8589,N_10880);
xnor U17015 (N_17015,N_8206,N_9078);
nand U17016 (N_17016,N_11294,N_10630);
nand U17017 (N_17017,N_12270,N_7365);
xnor U17018 (N_17018,N_11647,N_10728);
nand U17019 (N_17019,N_11642,N_8224);
nor U17020 (N_17020,N_11626,N_10488);
xnor U17021 (N_17021,N_6666,N_12387);
and U17022 (N_17022,N_7486,N_6796);
nand U17023 (N_17023,N_10758,N_10733);
nor U17024 (N_17024,N_9909,N_7949);
xnor U17025 (N_17025,N_12374,N_6286);
and U17026 (N_17026,N_12293,N_12035);
nor U17027 (N_17027,N_7187,N_8782);
or U17028 (N_17028,N_11038,N_7883);
and U17029 (N_17029,N_10401,N_6336);
nand U17030 (N_17030,N_11343,N_8737);
or U17031 (N_17031,N_6528,N_7484);
nor U17032 (N_17032,N_11508,N_10610);
nand U17033 (N_17033,N_7472,N_10915);
nand U17034 (N_17034,N_9477,N_10792);
and U17035 (N_17035,N_10563,N_10292);
nand U17036 (N_17036,N_10382,N_10173);
or U17037 (N_17037,N_11320,N_9552);
nor U17038 (N_17038,N_11370,N_7458);
and U17039 (N_17039,N_10275,N_6720);
or U17040 (N_17040,N_8655,N_9625);
or U17041 (N_17041,N_10036,N_11963);
nor U17042 (N_17042,N_9173,N_9558);
nand U17043 (N_17043,N_11689,N_6487);
or U17044 (N_17044,N_7355,N_9503);
and U17045 (N_17045,N_11834,N_10307);
xnor U17046 (N_17046,N_12393,N_9335);
and U17047 (N_17047,N_10406,N_9891);
or U17048 (N_17048,N_10901,N_12052);
xnor U17049 (N_17049,N_8057,N_7435);
nand U17050 (N_17050,N_10247,N_8469);
nand U17051 (N_17051,N_7984,N_7610);
xnor U17052 (N_17052,N_8591,N_10324);
and U17053 (N_17053,N_6281,N_11576);
nand U17054 (N_17054,N_11669,N_8315);
nand U17055 (N_17055,N_7988,N_6590);
and U17056 (N_17056,N_7413,N_7607);
and U17057 (N_17057,N_12414,N_7867);
nor U17058 (N_17058,N_9886,N_6747);
and U17059 (N_17059,N_10773,N_8532);
nor U17060 (N_17060,N_10013,N_8584);
xnor U17061 (N_17061,N_7424,N_11304);
xor U17062 (N_17062,N_10056,N_11998);
or U17063 (N_17063,N_9931,N_12283);
xor U17064 (N_17064,N_11005,N_7164);
nand U17065 (N_17065,N_12043,N_6772);
nor U17066 (N_17066,N_8005,N_7148);
nand U17067 (N_17067,N_10283,N_8834);
nor U17068 (N_17068,N_6632,N_9593);
nand U17069 (N_17069,N_11339,N_6345);
nand U17070 (N_17070,N_11404,N_11565);
and U17071 (N_17071,N_6274,N_7856);
nor U17072 (N_17072,N_11147,N_6290);
or U17073 (N_17073,N_7613,N_7273);
nand U17074 (N_17074,N_8727,N_9730);
nor U17075 (N_17075,N_10194,N_11556);
nand U17076 (N_17076,N_10601,N_12267);
nor U17077 (N_17077,N_12360,N_9806);
and U17078 (N_17078,N_11064,N_11361);
and U17079 (N_17079,N_8529,N_9380);
xor U17080 (N_17080,N_7983,N_9093);
xor U17081 (N_17081,N_8794,N_10697);
nor U17082 (N_17082,N_6600,N_6639);
or U17083 (N_17083,N_11973,N_8153);
nand U17084 (N_17084,N_7507,N_12240);
nor U17085 (N_17085,N_8121,N_9860);
xnor U17086 (N_17086,N_7591,N_7377);
nand U17087 (N_17087,N_6648,N_8092);
or U17088 (N_17088,N_9662,N_10329);
and U17089 (N_17089,N_6839,N_8396);
or U17090 (N_17090,N_10948,N_9683);
xnor U17091 (N_17091,N_12276,N_11001);
or U17092 (N_17092,N_9664,N_7450);
nor U17093 (N_17093,N_6351,N_9900);
xnor U17094 (N_17094,N_11822,N_8122);
nor U17095 (N_17095,N_11589,N_9109);
nand U17096 (N_17096,N_9221,N_7496);
xnor U17097 (N_17097,N_7737,N_10222);
nand U17098 (N_17098,N_11395,N_7786);
and U17099 (N_17099,N_9923,N_8531);
nand U17100 (N_17100,N_6808,N_7100);
nand U17101 (N_17101,N_7725,N_6410);
or U17102 (N_17102,N_7622,N_12222);
or U17103 (N_17103,N_11773,N_11736);
and U17104 (N_17104,N_12040,N_7801);
nor U17105 (N_17105,N_8565,N_8815);
nand U17106 (N_17106,N_8408,N_8448);
and U17107 (N_17107,N_8329,N_6477);
nor U17108 (N_17108,N_8999,N_9188);
nand U17109 (N_17109,N_7712,N_11552);
nor U17110 (N_17110,N_10378,N_11319);
and U17111 (N_17111,N_12104,N_10933);
nand U17112 (N_17112,N_7470,N_7987);
and U17113 (N_17113,N_6653,N_9618);
nand U17114 (N_17114,N_10703,N_10736);
nor U17115 (N_17115,N_8158,N_6532);
or U17116 (N_17116,N_6401,N_12249);
xnor U17117 (N_17117,N_7995,N_8554);
nand U17118 (N_17118,N_11587,N_10170);
and U17119 (N_17119,N_8242,N_11067);
nor U17120 (N_17120,N_11123,N_12036);
nand U17121 (N_17121,N_10246,N_9603);
or U17122 (N_17122,N_7856,N_12030);
nor U17123 (N_17123,N_6380,N_12087);
and U17124 (N_17124,N_6649,N_8548);
nand U17125 (N_17125,N_10659,N_6324);
or U17126 (N_17126,N_7703,N_8887);
and U17127 (N_17127,N_8975,N_9269);
and U17128 (N_17128,N_9772,N_9303);
nand U17129 (N_17129,N_11017,N_11746);
and U17130 (N_17130,N_9415,N_10490);
or U17131 (N_17131,N_7452,N_7498);
nor U17132 (N_17132,N_9398,N_10275);
or U17133 (N_17133,N_6723,N_10655);
nor U17134 (N_17134,N_8567,N_10263);
nor U17135 (N_17135,N_9718,N_10787);
or U17136 (N_17136,N_9773,N_7598);
nor U17137 (N_17137,N_7350,N_10384);
and U17138 (N_17138,N_7533,N_7393);
nand U17139 (N_17139,N_10581,N_10811);
or U17140 (N_17140,N_11306,N_7806);
xnor U17141 (N_17141,N_8959,N_11420);
or U17142 (N_17142,N_7761,N_9612);
nand U17143 (N_17143,N_11765,N_10243);
or U17144 (N_17144,N_9239,N_10071);
nor U17145 (N_17145,N_7627,N_11414);
or U17146 (N_17146,N_6344,N_10725);
nand U17147 (N_17147,N_10387,N_6923);
nand U17148 (N_17148,N_11334,N_10380);
xor U17149 (N_17149,N_8125,N_9638);
or U17150 (N_17150,N_7197,N_10245);
nand U17151 (N_17151,N_10752,N_8535);
or U17152 (N_17152,N_9701,N_6415);
nand U17153 (N_17153,N_12001,N_12481);
nand U17154 (N_17154,N_8349,N_12342);
xor U17155 (N_17155,N_12050,N_6626);
xnor U17156 (N_17156,N_8659,N_11163);
or U17157 (N_17157,N_10599,N_10318);
nand U17158 (N_17158,N_6575,N_7255);
and U17159 (N_17159,N_9740,N_12262);
xnor U17160 (N_17160,N_8996,N_6692);
and U17161 (N_17161,N_7542,N_10638);
and U17162 (N_17162,N_11743,N_12155);
nand U17163 (N_17163,N_6889,N_7425);
or U17164 (N_17164,N_7468,N_7216);
nand U17165 (N_17165,N_6817,N_8604);
or U17166 (N_17166,N_11210,N_11213);
or U17167 (N_17167,N_6485,N_7612);
nor U17168 (N_17168,N_12425,N_10688);
or U17169 (N_17169,N_7975,N_7108);
nand U17170 (N_17170,N_6388,N_6697);
nor U17171 (N_17171,N_9992,N_6314);
xnor U17172 (N_17172,N_6946,N_12326);
or U17173 (N_17173,N_8685,N_8720);
or U17174 (N_17174,N_11920,N_6476);
or U17175 (N_17175,N_10121,N_9472);
xnor U17176 (N_17176,N_6394,N_10680);
and U17177 (N_17177,N_8361,N_12160);
nor U17178 (N_17178,N_8409,N_6315);
xor U17179 (N_17179,N_10058,N_11473);
nor U17180 (N_17180,N_6991,N_8344);
xor U17181 (N_17181,N_10323,N_10137);
xnor U17182 (N_17182,N_10323,N_9842);
xnor U17183 (N_17183,N_11247,N_6327);
and U17184 (N_17184,N_6493,N_10445);
and U17185 (N_17185,N_10449,N_10941);
and U17186 (N_17186,N_12025,N_9947);
nand U17187 (N_17187,N_10771,N_11288);
nor U17188 (N_17188,N_7073,N_7516);
xnor U17189 (N_17189,N_11935,N_9613);
nor U17190 (N_17190,N_7042,N_7918);
nor U17191 (N_17191,N_7192,N_10321);
or U17192 (N_17192,N_7719,N_12288);
nand U17193 (N_17193,N_10672,N_8051);
nor U17194 (N_17194,N_9170,N_10662);
or U17195 (N_17195,N_8951,N_11480);
nor U17196 (N_17196,N_10909,N_9137);
xor U17197 (N_17197,N_11956,N_9358);
xor U17198 (N_17198,N_8642,N_6822);
nand U17199 (N_17199,N_11269,N_8903);
or U17200 (N_17200,N_7714,N_7791);
and U17201 (N_17201,N_9906,N_10529);
nand U17202 (N_17202,N_10131,N_9069);
nand U17203 (N_17203,N_8134,N_7584);
nand U17204 (N_17204,N_6535,N_12461);
nand U17205 (N_17205,N_7807,N_10438);
xnor U17206 (N_17206,N_6478,N_10176);
and U17207 (N_17207,N_12276,N_6615);
xor U17208 (N_17208,N_8464,N_9367);
nand U17209 (N_17209,N_8533,N_7454);
nor U17210 (N_17210,N_9986,N_10832);
xor U17211 (N_17211,N_6586,N_10077);
or U17212 (N_17212,N_11090,N_9824);
and U17213 (N_17213,N_9512,N_9707);
nor U17214 (N_17214,N_8966,N_9658);
xor U17215 (N_17215,N_6553,N_6744);
xor U17216 (N_17216,N_8064,N_11470);
and U17217 (N_17217,N_6818,N_10026);
nor U17218 (N_17218,N_10389,N_10256);
and U17219 (N_17219,N_10089,N_8063);
and U17220 (N_17220,N_8426,N_11316);
nor U17221 (N_17221,N_9876,N_8491);
and U17222 (N_17222,N_10432,N_10205);
and U17223 (N_17223,N_11552,N_11166);
and U17224 (N_17224,N_9700,N_8109);
nor U17225 (N_17225,N_6846,N_12264);
nor U17226 (N_17226,N_11606,N_9571);
nand U17227 (N_17227,N_7648,N_10114);
or U17228 (N_17228,N_9852,N_11635);
nand U17229 (N_17229,N_6657,N_11697);
xor U17230 (N_17230,N_7549,N_9558);
or U17231 (N_17231,N_7895,N_7683);
nor U17232 (N_17232,N_8394,N_7467);
or U17233 (N_17233,N_11151,N_11413);
xor U17234 (N_17234,N_12195,N_11868);
and U17235 (N_17235,N_8248,N_12144);
nand U17236 (N_17236,N_11076,N_8925);
and U17237 (N_17237,N_10207,N_10932);
nand U17238 (N_17238,N_8809,N_11229);
xnor U17239 (N_17239,N_10064,N_7908);
and U17240 (N_17240,N_11521,N_12451);
or U17241 (N_17241,N_6594,N_10902);
xnor U17242 (N_17242,N_8061,N_11187);
xor U17243 (N_17243,N_10913,N_9273);
nand U17244 (N_17244,N_12186,N_8948);
nor U17245 (N_17245,N_6797,N_8139);
and U17246 (N_17246,N_7157,N_7761);
xor U17247 (N_17247,N_11781,N_10906);
xnor U17248 (N_17248,N_11482,N_8792);
nand U17249 (N_17249,N_10543,N_11597);
nand U17250 (N_17250,N_8481,N_11591);
and U17251 (N_17251,N_11198,N_12132);
and U17252 (N_17252,N_11825,N_6266);
nor U17253 (N_17253,N_12468,N_6438);
xnor U17254 (N_17254,N_11653,N_12352);
xor U17255 (N_17255,N_11629,N_10768);
or U17256 (N_17256,N_10193,N_7279);
and U17257 (N_17257,N_11552,N_12396);
nor U17258 (N_17258,N_9234,N_11331);
xnor U17259 (N_17259,N_6701,N_9042);
and U17260 (N_17260,N_10747,N_7200);
xnor U17261 (N_17261,N_10965,N_6444);
and U17262 (N_17262,N_9405,N_12445);
nor U17263 (N_17263,N_6521,N_12075);
and U17264 (N_17264,N_11782,N_10617);
or U17265 (N_17265,N_7696,N_12231);
nand U17266 (N_17266,N_8284,N_10508);
nor U17267 (N_17267,N_10795,N_10433);
xnor U17268 (N_17268,N_11697,N_8025);
and U17269 (N_17269,N_8529,N_10404);
or U17270 (N_17270,N_8339,N_10643);
xnor U17271 (N_17271,N_7564,N_7238);
and U17272 (N_17272,N_9832,N_10275);
and U17273 (N_17273,N_9654,N_9148);
and U17274 (N_17274,N_6415,N_10032);
nand U17275 (N_17275,N_9495,N_9905);
xor U17276 (N_17276,N_11561,N_9765);
xor U17277 (N_17277,N_11778,N_9126);
nand U17278 (N_17278,N_9743,N_8042);
and U17279 (N_17279,N_10985,N_7323);
or U17280 (N_17280,N_6900,N_9251);
nand U17281 (N_17281,N_10195,N_11274);
nor U17282 (N_17282,N_7241,N_7578);
and U17283 (N_17283,N_11902,N_9449);
or U17284 (N_17284,N_7206,N_10317);
nand U17285 (N_17285,N_8161,N_8958);
nor U17286 (N_17286,N_11257,N_6424);
and U17287 (N_17287,N_12415,N_12216);
xor U17288 (N_17288,N_11422,N_11585);
nand U17289 (N_17289,N_10646,N_7056);
nor U17290 (N_17290,N_11858,N_7328);
nor U17291 (N_17291,N_11029,N_12004);
and U17292 (N_17292,N_11292,N_6909);
xnor U17293 (N_17293,N_6317,N_6660);
nor U17294 (N_17294,N_7253,N_6973);
and U17295 (N_17295,N_10604,N_9248);
nand U17296 (N_17296,N_10079,N_11630);
or U17297 (N_17297,N_7919,N_7054);
nor U17298 (N_17298,N_8851,N_8137);
xor U17299 (N_17299,N_11607,N_6515);
nand U17300 (N_17300,N_9819,N_9084);
nor U17301 (N_17301,N_6776,N_7474);
xor U17302 (N_17302,N_9913,N_9056);
nor U17303 (N_17303,N_12290,N_11338);
nor U17304 (N_17304,N_10877,N_10714);
and U17305 (N_17305,N_11731,N_12397);
or U17306 (N_17306,N_11643,N_9646);
nand U17307 (N_17307,N_6357,N_7821);
or U17308 (N_17308,N_10662,N_8873);
xor U17309 (N_17309,N_10938,N_8249);
nor U17310 (N_17310,N_8050,N_7357);
nor U17311 (N_17311,N_9705,N_10223);
and U17312 (N_17312,N_8241,N_7590);
nor U17313 (N_17313,N_11412,N_6524);
xnor U17314 (N_17314,N_8875,N_11229);
nand U17315 (N_17315,N_9056,N_9609);
or U17316 (N_17316,N_12339,N_7531);
nor U17317 (N_17317,N_12425,N_6798);
nand U17318 (N_17318,N_7949,N_9814);
and U17319 (N_17319,N_6517,N_7385);
nor U17320 (N_17320,N_8579,N_9489);
or U17321 (N_17321,N_10063,N_7017);
or U17322 (N_17322,N_8837,N_8293);
or U17323 (N_17323,N_11431,N_12486);
or U17324 (N_17324,N_8492,N_11890);
xnor U17325 (N_17325,N_9901,N_10959);
xor U17326 (N_17326,N_10225,N_6744);
nor U17327 (N_17327,N_12248,N_8833);
or U17328 (N_17328,N_8848,N_11722);
nor U17329 (N_17329,N_6941,N_9935);
or U17330 (N_17330,N_8783,N_12007);
and U17331 (N_17331,N_10837,N_9114);
or U17332 (N_17332,N_8846,N_8863);
xor U17333 (N_17333,N_10384,N_11315);
nand U17334 (N_17334,N_11461,N_6585);
and U17335 (N_17335,N_9444,N_10674);
nor U17336 (N_17336,N_6330,N_7962);
and U17337 (N_17337,N_6297,N_11431);
and U17338 (N_17338,N_11684,N_11130);
or U17339 (N_17339,N_10740,N_8024);
or U17340 (N_17340,N_10645,N_9937);
and U17341 (N_17341,N_8441,N_8080);
nor U17342 (N_17342,N_8262,N_8681);
or U17343 (N_17343,N_9571,N_11000);
or U17344 (N_17344,N_10711,N_8351);
nor U17345 (N_17345,N_10459,N_10746);
nand U17346 (N_17346,N_10785,N_9879);
and U17347 (N_17347,N_11377,N_11037);
nor U17348 (N_17348,N_8858,N_7424);
or U17349 (N_17349,N_9941,N_8076);
nor U17350 (N_17350,N_10176,N_7996);
nor U17351 (N_17351,N_10225,N_9339);
and U17352 (N_17352,N_7160,N_9403);
xnor U17353 (N_17353,N_8443,N_11893);
nand U17354 (N_17354,N_9626,N_8234);
nand U17355 (N_17355,N_8081,N_9889);
nor U17356 (N_17356,N_9701,N_6480);
or U17357 (N_17357,N_8166,N_7219);
and U17358 (N_17358,N_9740,N_11781);
or U17359 (N_17359,N_9423,N_10040);
or U17360 (N_17360,N_6865,N_11455);
nand U17361 (N_17361,N_7743,N_11603);
xor U17362 (N_17362,N_12422,N_7030);
xor U17363 (N_17363,N_9242,N_10967);
nand U17364 (N_17364,N_6456,N_7550);
xor U17365 (N_17365,N_9191,N_11761);
nand U17366 (N_17366,N_12177,N_8436);
xnor U17367 (N_17367,N_10557,N_7912);
xnor U17368 (N_17368,N_11107,N_8972);
nor U17369 (N_17369,N_11014,N_9764);
nor U17370 (N_17370,N_10132,N_9676);
nand U17371 (N_17371,N_11988,N_7225);
nand U17372 (N_17372,N_12178,N_10570);
and U17373 (N_17373,N_10982,N_10638);
nand U17374 (N_17374,N_11501,N_7816);
and U17375 (N_17375,N_8619,N_9465);
xnor U17376 (N_17376,N_12293,N_7221);
and U17377 (N_17377,N_11814,N_9029);
or U17378 (N_17378,N_12151,N_12055);
and U17379 (N_17379,N_11449,N_7176);
xor U17380 (N_17380,N_9774,N_8470);
nand U17381 (N_17381,N_6253,N_11151);
nor U17382 (N_17382,N_10750,N_10657);
nand U17383 (N_17383,N_10041,N_8205);
and U17384 (N_17384,N_7316,N_8005);
and U17385 (N_17385,N_10594,N_7015);
nand U17386 (N_17386,N_9979,N_9216);
and U17387 (N_17387,N_6587,N_12294);
nor U17388 (N_17388,N_10294,N_7118);
and U17389 (N_17389,N_12424,N_7701);
nand U17390 (N_17390,N_10614,N_11340);
xnor U17391 (N_17391,N_7968,N_10841);
or U17392 (N_17392,N_12376,N_12481);
and U17393 (N_17393,N_11203,N_6449);
and U17394 (N_17394,N_6562,N_11130);
and U17395 (N_17395,N_8653,N_10371);
nand U17396 (N_17396,N_6442,N_8791);
or U17397 (N_17397,N_7941,N_10209);
nand U17398 (N_17398,N_10750,N_9945);
and U17399 (N_17399,N_10878,N_10039);
xor U17400 (N_17400,N_7635,N_9133);
nor U17401 (N_17401,N_12326,N_8551);
nor U17402 (N_17402,N_8592,N_11681);
nor U17403 (N_17403,N_9162,N_11388);
nand U17404 (N_17404,N_9839,N_11959);
nand U17405 (N_17405,N_8486,N_6572);
nor U17406 (N_17406,N_10823,N_7160);
and U17407 (N_17407,N_9730,N_7085);
xnor U17408 (N_17408,N_11435,N_11232);
and U17409 (N_17409,N_8786,N_8418);
nor U17410 (N_17410,N_10470,N_10986);
and U17411 (N_17411,N_12410,N_6482);
or U17412 (N_17412,N_10997,N_11782);
nand U17413 (N_17413,N_7584,N_10884);
and U17414 (N_17414,N_8864,N_8013);
or U17415 (N_17415,N_7855,N_6970);
or U17416 (N_17416,N_9691,N_9368);
and U17417 (N_17417,N_7776,N_11071);
nor U17418 (N_17418,N_10039,N_6996);
and U17419 (N_17419,N_12352,N_9394);
and U17420 (N_17420,N_8741,N_8902);
nand U17421 (N_17421,N_7306,N_8806);
and U17422 (N_17422,N_9774,N_11166);
xor U17423 (N_17423,N_12194,N_8296);
and U17424 (N_17424,N_9249,N_11863);
xnor U17425 (N_17425,N_8707,N_10532);
nand U17426 (N_17426,N_9059,N_8451);
xor U17427 (N_17427,N_9467,N_10505);
nor U17428 (N_17428,N_11927,N_12203);
or U17429 (N_17429,N_11580,N_11016);
or U17430 (N_17430,N_8372,N_9182);
xnor U17431 (N_17431,N_8688,N_11037);
and U17432 (N_17432,N_8385,N_10154);
nand U17433 (N_17433,N_9877,N_10582);
nand U17434 (N_17434,N_7470,N_11243);
nor U17435 (N_17435,N_10010,N_10451);
nand U17436 (N_17436,N_8036,N_8002);
and U17437 (N_17437,N_10505,N_7455);
xor U17438 (N_17438,N_8998,N_10464);
xor U17439 (N_17439,N_7684,N_10480);
and U17440 (N_17440,N_11107,N_6656);
xnor U17441 (N_17441,N_7562,N_12310);
nand U17442 (N_17442,N_8257,N_9290);
and U17443 (N_17443,N_8064,N_7056);
or U17444 (N_17444,N_10004,N_7921);
or U17445 (N_17445,N_12053,N_12039);
nand U17446 (N_17446,N_9010,N_8410);
nor U17447 (N_17447,N_8899,N_7685);
nand U17448 (N_17448,N_6850,N_12466);
xnor U17449 (N_17449,N_7747,N_6349);
or U17450 (N_17450,N_6989,N_8086);
and U17451 (N_17451,N_11875,N_10602);
nand U17452 (N_17452,N_10561,N_6870);
xnor U17453 (N_17453,N_6813,N_11248);
xor U17454 (N_17454,N_6794,N_9981);
nand U17455 (N_17455,N_8033,N_9194);
nor U17456 (N_17456,N_11313,N_8137);
xnor U17457 (N_17457,N_9453,N_7894);
xor U17458 (N_17458,N_10021,N_8689);
xor U17459 (N_17459,N_11939,N_7337);
and U17460 (N_17460,N_9254,N_8177);
and U17461 (N_17461,N_11003,N_11825);
nor U17462 (N_17462,N_11035,N_10979);
or U17463 (N_17463,N_11907,N_9289);
nor U17464 (N_17464,N_11672,N_12023);
and U17465 (N_17465,N_10384,N_9805);
xnor U17466 (N_17466,N_6384,N_7454);
xor U17467 (N_17467,N_11535,N_6505);
nor U17468 (N_17468,N_9328,N_12213);
nor U17469 (N_17469,N_6827,N_11266);
nor U17470 (N_17470,N_8321,N_10453);
nor U17471 (N_17471,N_12393,N_11391);
nor U17472 (N_17472,N_7413,N_6853);
and U17473 (N_17473,N_9572,N_7029);
nand U17474 (N_17474,N_11952,N_10204);
nor U17475 (N_17475,N_6935,N_8340);
or U17476 (N_17476,N_7887,N_11561);
xnor U17477 (N_17477,N_11202,N_12396);
or U17478 (N_17478,N_6472,N_7089);
nor U17479 (N_17479,N_11950,N_10821);
xnor U17480 (N_17480,N_10473,N_10601);
xnor U17481 (N_17481,N_7044,N_9407);
or U17482 (N_17482,N_8367,N_11820);
nor U17483 (N_17483,N_6996,N_11879);
nand U17484 (N_17484,N_8315,N_8168);
nand U17485 (N_17485,N_9591,N_10306);
or U17486 (N_17486,N_6797,N_8285);
xor U17487 (N_17487,N_8843,N_11631);
nand U17488 (N_17488,N_7978,N_12195);
nor U17489 (N_17489,N_7659,N_12465);
nand U17490 (N_17490,N_6551,N_8138);
or U17491 (N_17491,N_11083,N_9155);
or U17492 (N_17492,N_8666,N_10934);
and U17493 (N_17493,N_9735,N_12167);
or U17494 (N_17494,N_12129,N_6874);
nand U17495 (N_17495,N_8223,N_12168);
nor U17496 (N_17496,N_10955,N_9015);
nor U17497 (N_17497,N_7876,N_7523);
or U17498 (N_17498,N_7021,N_8598);
nor U17499 (N_17499,N_8853,N_6937);
or U17500 (N_17500,N_8022,N_6475);
and U17501 (N_17501,N_8545,N_10586);
nand U17502 (N_17502,N_11621,N_7338);
xnor U17503 (N_17503,N_9869,N_9144);
nor U17504 (N_17504,N_6504,N_8602);
and U17505 (N_17505,N_12131,N_11775);
xor U17506 (N_17506,N_7872,N_9778);
and U17507 (N_17507,N_10873,N_9567);
nand U17508 (N_17508,N_11706,N_12053);
nor U17509 (N_17509,N_8132,N_8787);
and U17510 (N_17510,N_6376,N_12002);
or U17511 (N_17511,N_10079,N_8546);
and U17512 (N_17512,N_9119,N_11529);
and U17513 (N_17513,N_6426,N_7170);
nor U17514 (N_17514,N_8268,N_7058);
nand U17515 (N_17515,N_8431,N_10059);
nor U17516 (N_17516,N_11310,N_11510);
xnor U17517 (N_17517,N_9876,N_7492);
nor U17518 (N_17518,N_10961,N_11267);
and U17519 (N_17519,N_7059,N_6844);
nand U17520 (N_17520,N_7939,N_11676);
xnor U17521 (N_17521,N_8084,N_7253);
nor U17522 (N_17522,N_7318,N_7472);
and U17523 (N_17523,N_11525,N_7773);
nand U17524 (N_17524,N_12044,N_10537);
or U17525 (N_17525,N_7927,N_7421);
nor U17526 (N_17526,N_11536,N_6772);
nor U17527 (N_17527,N_10202,N_6838);
and U17528 (N_17528,N_12365,N_7854);
xor U17529 (N_17529,N_12267,N_10010);
nor U17530 (N_17530,N_11253,N_9641);
xnor U17531 (N_17531,N_6473,N_11759);
nor U17532 (N_17532,N_12309,N_10667);
nand U17533 (N_17533,N_10260,N_10063);
xor U17534 (N_17534,N_11883,N_10988);
and U17535 (N_17535,N_7006,N_12339);
nor U17536 (N_17536,N_9210,N_8752);
nand U17537 (N_17537,N_6790,N_7698);
nand U17538 (N_17538,N_9792,N_9625);
nand U17539 (N_17539,N_8014,N_7445);
or U17540 (N_17540,N_12012,N_8967);
xor U17541 (N_17541,N_10770,N_7074);
xor U17542 (N_17542,N_7046,N_8892);
nor U17543 (N_17543,N_11118,N_6522);
nand U17544 (N_17544,N_10052,N_7908);
xor U17545 (N_17545,N_11094,N_10266);
xor U17546 (N_17546,N_10966,N_8472);
and U17547 (N_17547,N_10229,N_7523);
nor U17548 (N_17548,N_9022,N_9845);
nand U17549 (N_17549,N_12454,N_10936);
or U17550 (N_17550,N_9976,N_11088);
and U17551 (N_17551,N_7315,N_10729);
nor U17552 (N_17552,N_12418,N_9431);
and U17553 (N_17553,N_10054,N_11267);
and U17554 (N_17554,N_7093,N_8535);
and U17555 (N_17555,N_9144,N_12156);
xnor U17556 (N_17556,N_7615,N_11230);
or U17557 (N_17557,N_7182,N_9359);
xnor U17558 (N_17558,N_9297,N_10832);
or U17559 (N_17559,N_9183,N_11651);
or U17560 (N_17560,N_11907,N_8314);
and U17561 (N_17561,N_7863,N_11672);
xor U17562 (N_17562,N_11481,N_7277);
xnor U17563 (N_17563,N_7595,N_8971);
or U17564 (N_17564,N_12334,N_9554);
and U17565 (N_17565,N_6702,N_11680);
and U17566 (N_17566,N_11324,N_6756);
and U17567 (N_17567,N_9506,N_10145);
and U17568 (N_17568,N_7109,N_11107);
nor U17569 (N_17569,N_10461,N_11109);
nand U17570 (N_17570,N_9396,N_10025);
and U17571 (N_17571,N_11789,N_8331);
nor U17572 (N_17572,N_6849,N_12054);
nand U17573 (N_17573,N_10673,N_9971);
nand U17574 (N_17574,N_11485,N_11182);
xnor U17575 (N_17575,N_8258,N_10061);
and U17576 (N_17576,N_8356,N_9315);
nand U17577 (N_17577,N_8283,N_8395);
xor U17578 (N_17578,N_10549,N_10859);
xnor U17579 (N_17579,N_11357,N_9189);
nand U17580 (N_17580,N_7152,N_12365);
xor U17581 (N_17581,N_7719,N_7517);
nand U17582 (N_17582,N_8826,N_9219);
nand U17583 (N_17583,N_6435,N_9970);
nor U17584 (N_17584,N_8679,N_9700);
and U17585 (N_17585,N_7462,N_9853);
xor U17586 (N_17586,N_11163,N_9212);
nand U17587 (N_17587,N_9884,N_6814);
or U17588 (N_17588,N_11204,N_7155);
or U17589 (N_17589,N_11371,N_11723);
or U17590 (N_17590,N_10242,N_11841);
or U17591 (N_17591,N_10158,N_11863);
nor U17592 (N_17592,N_11043,N_10174);
nor U17593 (N_17593,N_7364,N_9528);
or U17594 (N_17594,N_11789,N_7371);
and U17595 (N_17595,N_7401,N_8392);
xnor U17596 (N_17596,N_8653,N_10143);
nand U17597 (N_17597,N_9546,N_11092);
and U17598 (N_17598,N_8377,N_12048);
and U17599 (N_17599,N_9277,N_6364);
and U17600 (N_17600,N_6585,N_11194);
or U17601 (N_17601,N_7843,N_7684);
nand U17602 (N_17602,N_6562,N_11537);
nor U17603 (N_17603,N_10354,N_7133);
xor U17604 (N_17604,N_9292,N_7107);
and U17605 (N_17605,N_11096,N_8861);
nor U17606 (N_17606,N_7556,N_7793);
or U17607 (N_17607,N_9278,N_11007);
nand U17608 (N_17608,N_6518,N_6307);
or U17609 (N_17609,N_8699,N_7077);
xor U17610 (N_17610,N_9427,N_11628);
xor U17611 (N_17611,N_9710,N_6308);
nor U17612 (N_17612,N_10147,N_7059);
and U17613 (N_17613,N_9931,N_9329);
and U17614 (N_17614,N_8530,N_11332);
xnor U17615 (N_17615,N_11503,N_8607);
xor U17616 (N_17616,N_7681,N_9308);
xnor U17617 (N_17617,N_8040,N_6719);
or U17618 (N_17618,N_9416,N_8080);
nand U17619 (N_17619,N_9438,N_12180);
xor U17620 (N_17620,N_10243,N_9173);
and U17621 (N_17621,N_7926,N_8146);
nand U17622 (N_17622,N_6903,N_10839);
nand U17623 (N_17623,N_11761,N_7653);
and U17624 (N_17624,N_11058,N_7377);
xnor U17625 (N_17625,N_10925,N_12009);
nor U17626 (N_17626,N_11728,N_12138);
or U17627 (N_17627,N_12176,N_7552);
and U17628 (N_17628,N_9703,N_12094);
or U17629 (N_17629,N_9665,N_9111);
or U17630 (N_17630,N_8348,N_10687);
nor U17631 (N_17631,N_9744,N_8599);
nor U17632 (N_17632,N_10601,N_9365);
xor U17633 (N_17633,N_7541,N_9673);
and U17634 (N_17634,N_6761,N_8999);
and U17635 (N_17635,N_6798,N_11849);
or U17636 (N_17636,N_10450,N_9263);
or U17637 (N_17637,N_6445,N_10782);
or U17638 (N_17638,N_6456,N_8625);
xor U17639 (N_17639,N_12245,N_11747);
nand U17640 (N_17640,N_9502,N_9633);
nor U17641 (N_17641,N_8461,N_6706);
xnor U17642 (N_17642,N_10756,N_6683);
and U17643 (N_17643,N_12068,N_9643);
nand U17644 (N_17644,N_10118,N_9833);
xor U17645 (N_17645,N_11318,N_6317);
xor U17646 (N_17646,N_10838,N_6360);
nor U17647 (N_17647,N_11864,N_8116);
nand U17648 (N_17648,N_7227,N_8949);
nor U17649 (N_17649,N_7465,N_7358);
and U17650 (N_17650,N_7197,N_11330);
xnor U17651 (N_17651,N_8437,N_8178);
or U17652 (N_17652,N_6568,N_8345);
nor U17653 (N_17653,N_6404,N_10049);
nand U17654 (N_17654,N_10037,N_7788);
and U17655 (N_17655,N_11401,N_9617);
or U17656 (N_17656,N_6636,N_7942);
nand U17657 (N_17657,N_11633,N_12367);
or U17658 (N_17658,N_9569,N_7876);
nand U17659 (N_17659,N_9958,N_11425);
xor U17660 (N_17660,N_11608,N_9901);
or U17661 (N_17661,N_8323,N_11170);
nor U17662 (N_17662,N_9196,N_10593);
or U17663 (N_17663,N_8626,N_11251);
nor U17664 (N_17664,N_11319,N_12470);
xnor U17665 (N_17665,N_6513,N_6525);
nor U17666 (N_17666,N_7342,N_7893);
xor U17667 (N_17667,N_8078,N_11796);
or U17668 (N_17668,N_9998,N_7369);
nor U17669 (N_17669,N_10948,N_11073);
nor U17670 (N_17670,N_9277,N_10165);
or U17671 (N_17671,N_9056,N_10103);
xnor U17672 (N_17672,N_8314,N_7434);
nand U17673 (N_17673,N_7247,N_9246);
nand U17674 (N_17674,N_10230,N_9371);
or U17675 (N_17675,N_11115,N_10826);
nor U17676 (N_17676,N_11367,N_7316);
nand U17677 (N_17677,N_6264,N_10656);
nand U17678 (N_17678,N_9908,N_6454);
or U17679 (N_17679,N_10764,N_7168);
or U17680 (N_17680,N_9455,N_7061);
and U17681 (N_17681,N_6870,N_12304);
nand U17682 (N_17682,N_12003,N_8276);
and U17683 (N_17683,N_7389,N_7225);
nand U17684 (N_17684,N_8273,N_6563);
xnor U17685 (N_17685,N_7899,N_6504);
xor U17686 (N_17686,N_9469,N_9239);
or U17687 (N_17687,N_9600,N_6324);
nor U17688 (N_17688,N_7156,N_11004);
and U17689 (N_17689,N_11514,N_8814);
xor U17690 (N_17690,N_7745,N_10375);
xor U17691 (N_17691,N_8388,N_8614);
and U17692 (N_17692,N_11107,N_11763);
xor U17693 (N_17693,N_6570,N_10042);
xnor U17694 (N_17694,N_9834,N_6664);
xnor U17695 (N_17695,N_6715,N_7265);
xnor U17696 (N_17696,N_11143,N_9079);
xnor U17697 (N_17697,N_8427,N_6523);
and U17698 (N_17698,N_10019,N_9303);
nand U17699 (N_17699,N_8719,N_11736);
nor U17700 (N_17700,N_8340,N_12429);
nand U17701 (N_17701,N_9370,N_7672);
xor U17702 (N_17702,N_8060,N_8956);
and U17703 (N_17703,N_6333,N_8851);
nor U17704 (N_17704,N_11064,N_7395);
nand U17705 (N_17705,N_8290,N_10341);
and U17706 (N_17706,N_12204,N_8846);
xor U17707 (N_17707,N_11969,N_10064);
nor U17708 (N_17708,N_10406,N_8653);
nor U17709 (N_17709,N_6335,N_9685);
or U17710 (N_17710,N_6508,N_9360);
xor U17711 (N_17711,N_9982,N_8660);
or U17712 (N_17712,N_6711,N_6657);
or U17713 (N_17713,N_7158,N_11843);
and U17714 (N_17714,N_10951,N_8466);
xor U17715 (N_17715,N_7608,N_11821);
nor U17716 (N_17716,N_11120,N_7542);
nand U17717 (N_17717,N_9316,N_9014);
xor U17718 (N_17718,N_7825,N_11052);
nor U17719 (N_17719,N_7969,N_10784);
nand U17720 (N_17720,N_10033,N_10709);
xor U17721 (N_17721,N_7292,N_9994);
nand U17722 (N_17722,N_11442,N_11162);
nand U17723 (N_17723,N_6712,N_6615);
nand U17724 (N_17724,N_11718,N_9350);
nand U17725 (N_17725,N_7014,N_7643);
or U17726 (N_17726,N_8019,N_9325);
nand U17727 (N_17727,N_10914,N_7143);
and U17728 (N_17728,N_9042,N_7035);
or U17729 (N_17729,N_7396,N_7905);
nand U17730 (N_17730,N_10028,N_7037);
or U17731 (N_17731,N_9711,N_8864);
xnor U17732 (N_17732,N_10122,N_6718);
nor U17733 (N_17733,N_7103,N_8785);
nand U17734 (N_17734,N_10164,N_8227);
nor U17735 (N_17735,N_8708,N_9759);
xor U17736 (N_17736,N_6503,N_7671);
and U17737 (N_17737,N_9619,N_11596);
or U17738 (N_17738,N_12080,N_8517);
xnor U17739 (N_17739,N_8400,N_10992);
nor U17740 (N_17740,N_6915,N_10352);
nand U17741 (N_17741,N_8082,N_6560);
and U17742 (N_17742,N_11654,N_11650);
xnor U17743 (N_17743,N_10502,N_12212);
nand U17744 (N_17744,N_9732,N_9747);
nor U17745 (N_17745,N_12272,N_9340);
nor U17746 (N_17746,N_8016,N_9355);
xnor U17747 (N_17747,N_9514,N_7558);
and U17748 (N_17748,N_7501,N_10949);
or U17749 (N_17749,N_12293,N_11441);
and U17750 (N_17750,N_10281,N_7456);
or U17751 (N_17751,N_10149,N_8495);
and U17752 (N_17752,N_7582,N_8147);
nor U17753 (N_17753,N_9475,N_10818);
nor U17754 (N_17754,N_11929,N_7615);
and U17755 (N_17755,N_11528,N_6478);
nor U17756 (N_17756,N_9882,N_11766);
or U17757 (N_17757,N_10871,N_8742);
nand U17758 (N_17758,N_6402,N_10468);
nand U17759 (N_17759,N_8570,N_8013);
nand U17760 (N_17760,N_7703,N_9120);
and U17761 (N_17761,N_11281,N_12271);
nor U17762 (N_17762,N_7499,N_8109);
nand U17763 (N_17763,N_9713,N_7366);
nor U17764 (N_17764,N_12030,N_7138);
and U17765 (N_17765,N_12426,N_7779);
nand U17766 (N_17766,N_11213,N_10580);
and U17767 (N_17767,N_10769,N_11533);
and U17768 (N_17768,N_10350,N_10005);
xor U17769 (N_17769,N_9463,N_11911);
nand U17770 (N_17770,N_11693,N_9607);
nand U17771 (N_17771,N_9321,N_6612);
or U17772 (N_17772,N_7670,N_9418);
nor U17773 (N_17773,N_7625,N_6472);
or U17774 (N_17774,N_8725,N_8536);
xor U17775 (N_17775,N_6579,N_9568);
nor U17776 (N_17776,N_7933,N_8368);
nor U17777 (N_17777,N_8512,N_12449);
nor U17778 (N_17778,N_7794,N_10229);
or U17779 (N_17779,N_7419,N_10611);
nand U17780 (N_17780,N_10120,N_11972);
nor U17781 (N_17781,N_8289,N_9112);
nor U17782 (N_17782,N_12218,N_8064);
nand U17783 (N_17783,N_11223,N_11423);
and U17784 (N_17784,N_10578,N_8209);
xor U17785 (N_17785,N_10580,N_7998);
nand U17786 (N_17786,N_6670,N_10254);
xnor U17787 (N_17787,N_11090,N_10324);
and U17788 (N_17788,N_11775,N_11617);
nor U17789 (N_17789,N_11471,N_10574);
nor U17790 (N_17790,N_12131,N_11543);
xnor U17791 (N_17791,N_8464,N_10533);
nor U17792 (N_17792,N_7793,N_6532);
nor U17793 (N_17793,N_12138,N_9715);
nand U17794 (N_17794,N_7170,N_8075);
nor U17795 (N_17795,N_8480,N_10305);
nor U17796 (N_17796,N_11946,N_8623);
xnor U17797 (N_17797,N_6314,N_7074);
and U17798 (N_17798,N_7811,N_11680);
nor U17799 (N_17799,N_10474,N_7644);
nor U17800 (N_17800,N_10531,N_7517);
or U17801 (N_17801,N_6432,N_7263);
and U17802 (N_17802,N_6802,N_11869);
or U17803 (N_17803,N_11571,N_11535);
or U17804 (N_17804,N_10016,N_10139);
nand U17805 (N_17805,N_7274,N_9849);
xnor U17806 (N_17806,N_7121,N_12101);
and U17807 (N_17807,N_7807,N_10364);
or U17808 (N_17808,N_6382,N_6254);
nand U17809 (N_17809,N_10964,N_10638);
and U17810 (N_17810,N_7254,N_6830);
nor U17811 (N_17811,N_7874,N_8027);
or U17812 (N_17812,N_9225,N_8514);
nor U17813 (N_17813,N_7951,N_11764);
and U17814 (N_17814,N_9057,N_8505);
and U17815 (N_17815,N_7255,N_11543);
nand U17816 (N_17816,N_7248,N_8358);
and U17817 (N_17817,N_12398,N_10815);
and U17818 (N_17818,N_10579,N_9413);
xnor U17819 (N_17819,N_11451,N_11940);
or U17820 (N_17820,N_12224,N_8621);
nor U17821 (N_17821,N_10373,N_11451);
xnor U17822 (N_17822,N_10348,N_7345);
or U17823 (N_17823,N_11567,N_10691);
xor U17824 (N_17824,N_10198,N_7410);
nor U17825 (N_17825,N_11230,N_6866);
or U17826 (N_17826,N_8042,N_9721);
xnor U17827 (N_17827,N_8839,N_11767);
nor U17828 (N_17828,N_7510,N_11384);
and U17829 (N_17829,N_6844,N_11630);
nor U17830 (N_17830,N_10827,N_6258);
nand U17831 (N_17831,N_7179,N_8762);
nor U17832 (N_17832,N_10583,N_10244);
nand U17833 (N_17833,N_9813,N_7152);
xor U17834 (N_17834,N_10292,N_12298);
nand U17835 (N_17835,N_7317,N_12189);
and U17836 (N_17836,N_8103,N_6799);
xnor U17837 (N_17837,N_9098,N_11642);
xnor U17838 (N_17838,N_11330,N_8845);
nand U17839 (N_17839,N_8959,N_6698);
nand U17840 (N_17840,N_7406,N_8337);
nand U17841 (N_17841,N_9247,N_11745);
xnor U17842 (N_17842,N_6411,N_10324);
or U17843 (N_17843,N_6763,N_9776);
nor U17844 (N_17844,N_12105,N_7443);
and U17845 (N_17845,N_9945,N_10325);
and U17846 (N_17846,N_11595,N_10413);
or U17847 (N_17847,N_7901,N_9048);
or U17848 (N_17848,N_10543,N_10231);
nand U17849 (N_17849,N_7597,N_11326);
xor U17850 (N_17850,N_10178,N_11142);
xor U17851 (N_17851,N_11532,N_6967);
and U17852 (N_17852,N_7565,N_7110);
xor U17853 (N_17853,N_8216,N_10493);
xnor U17854 (N_17854,N_12205,N_9847);
nor U17855 (N_17855,N_12011,N_12121);
xor U17856 (N_17856,N_10762,N_8278);
nand U17857 (N_17857,N_6769,N_9764);
nor U17858 (N_17858,N_6255,N_11161);
and U17859 (N_17859,N_9269,N_11742);
and U17860 (N_17860,N_10796,N_7273);
nor U17861 (N_17861,N_7774,N_7753);
nor U17862 (N_17862,N_11872,N_7340);
and U17863 (N_17863,N_6269,N_7003);
or U17864 (N_17864,N_11084,N_7568);
nor U17865 (N_17865,N_9212,N_7518);
nor U17866 (N_17866,N_9375,N_7784);
nand U17867 (N_17867,N_10414,N_8782);
nor U17868 (N_17868,N_12383,N_8964);
nor U17869 (N_17869,N_11212,N_9710);
or U17870 (N_17870,N_6717,N_10963);
or U17871 (N_17871,N_10340,N_10576);
xnor U17872 (N_17872,N_12203,N_7276);
or U17873 (N_17873,N_11937,N_9705);
and U17874 (N_17874,N_12107,N_10351);
nand U17875 (N_17875,N_10832,N_11969);
or U17876 (N_17876,N_7201,N_10930);
nor U17877 (N_17877,N_11256,N_9613);
and U17878 (N_17878,N_10339,N_7339);
or U17879 (N_17879,N_10692,N_10208);
xnor U17880 (N_17880,N_7503,N_9336);
nor U17881 (N_17881,N_12150,N_8748);
or U17882 (N_17882,N_8592,N_8915);
nand U17883 (N_17883,N_8704,N_7329);
nand U17884 (N_17884,N_6306,N_6656);
xnor U17885 (N_17885,N_7175,N_8256);
nor U17886 (N_17886,N_12417,N_7556);
and U17887 (N_17887,N_9870,N_7184);
nor U17888 (N_17888,N_9298,N_10531);
and U17889 (N_17889,N_11556,N_10021);
xor U17890 (N_17890,N_9741,N_9351);
and U17891 (N_17891,N_7631,N_10538);
nor U17892 (N_17892,N_12442,N_7468);
xnor U17893 (N_17893,N_6619,N_7228);
nand U17894 (N_17894,N_6849,N_10862);
nand U17895 (N_17895,N_8179,N_9749);
xor U17896 (N_17896,N_9857,N_9751);
nor U17897 (N_17897,N_8763,N_10996);
xor U17898 (N_17898,N_8463,N_7160);
or U17899 (N_17899,N_12029,N_9810);
or U17900 (N_17900,N_10386,N_8543);
nand U17901 (N_17901,N_9423,N_7139);
xor U17902 (N_17902,N_8770,N_8565);
xnor U17903 (N_17903,N_11054,N_6947);
xnor U17904 (N_17904,N_10141,N_8942);
nor U17905 (N_17905,N_7009,N_7023);
xnor U17906 (N_17906,N_9853,N_8847);
and U17907 (N_17907,N_9562,N_11514);
nand U17908 (N_17908,N_7890,N_9402);
or U17909 (N_17909,N_10304,N_9079);
nand U17910 (N_17910,N_12019,N_6835);
nand U17911 (N_17911,N_10774,N_7384);
xor U17912 (N_17912,N_9130,N_11791);
and U17913 (N_17913,N_6527,N_9405);
nand U17914 (N_17914,N_7031,N_7705);
or U17915 (N_17915,N_11624,N_8476);
nor U17916 (N_17916,N_11222,N_8846);
nor U17917 (N_17917,N_8285,N_7629);
or U17918 (N_17918,N_9555,N_7890);
and U17919 (N_17919,N_9539,N_7524);
nor U17920 (N_17920,N_8127,N_8219);
nand U17921 (N_17921,N_7688,N_10212);
xor U17922 (N_17922,N_8864,N_11370);
nor U17923 (N_17923,N_8952,N_9335);
or U17924 (N_17924,N_12117,N_10727);
or U17925 (N_17925,N_8843,N_6847);
and U17926 (N_17926,N_7695,N_11181);
xnor U17927 (N_17927,N_8822,N_6988);
xor U17928 (N_17928,N_8797,N_8008);
and U17929 (N_17929,N_8484,N_8697);
or U17930 (N_17930,N_11865,N_11938);
xor U17931 (N_17931,N_8755,N_10401);
nand U17932 (N_17932,N_10999,N_8017);
nand U17933 (N_17933,N_7402,N_6526);
or U17934 (N_17934,N_8286,N_7813);
xnor U17935 (N_17935,N_10668,N_11196);
nor U17936 (N_17936,N_9015,N_9486);
and U17937 (N_17937,N_10436,N_7024);
xnor U17938 (N_17938,N_7684,N_7737);
nand U17939 (N_17939,N_11128,N_10726);
nor U17940 (N_17940,N_8840,N_7423);
nor U17941 (N_17941,N_6825,N_9390);
xnor U17942 (N_17942,N_9029,N_11776);
nand U17943 (N_17943,N_9820,N_7587);
and U17944 (N_17944,N_10702,N_11186);
nand U17945 (N_17945,N_12423,N_9062);
nor U17946 (N_17946,N_6587,N_9084);
and U17947 (N_17947,N_10453,N_8567);
and U17948 (N_17948,N_9232,N_9603);
nor U17949 (N_17949,N_7931,N_8405);
xnor U17950 (N_17950,N_10980,N_6480);
xnor U17951 (N_17951,N_10505,N_9874);
xor U17952 (N_17952,N_9937,N_11899);
or U17953 (N_17953,N_9172,N_9753);
nand U17954 (N_17954,N_10935,N_7326);
and U17955 (N_17955,N_11897,N_9457);
and U17956 (N_17956,N_9203,N_7578);
and U17957 (N_17957,N_7759,N_8069);
xnor U17958 (N_17958,N_8781,N_8003);
or U17959 (N_17959,N_7220,N_6485);
xnor U17960 (N_17960,N_6475,N_10450);
or U17961 (N_17961,N_6959,N_6402);
xnor U17962 (N_17962,N_9438,N_9580);
nand U17963 (N_17963,N_8811,N_10306);
or U17964 (N_17964,N_7645,N_6909);
and U17965 (N_17965,N_7264,N_7818);
and U17966 (N_17966,N_7728,N_12219);
and U17967 (N_17967,N_10921,N_9049);
nor U17968 (N_17968,N_6297,N_10349);
nor U17969 (N_17969,N_7179,N_6259);
xnor U17970 (N_17970,N_11954,N_7615);
xnor U17971 (N_17971,N_10306,N_11188);
or U17972 (N_17972,N_9938,N_10871);
nand U17973 (N_17973,N_7931,N_8881);
and U17974 (N_17974,N_6313,N_11784);
and U17975 (N_17975,N_10159,N_8274);
and U17976 (N_17976,N_6400,N_9936);
or U17977 (N_17977,N_6365,N_10360);
nand U17978 (N_17978,N_12241,N_12337);
nand U17979 (N_17979,N_8819,N_10630);
or U17980 (N_17980,N_10235,N_11607);
nor U17981 (N_17981,N_7574,N_8343);
nor U17982 (N_17982,N_7850,N_8622);
nand U17983 (N_17983,N_10819,N_6733);
and U17984 (N_17984,N_10879,N_9349);
nor U17985 (N_17985,N_6732,N_11063);
nor U17986 (N_17986,N_10968,N_11844);
xor U17987 (N_17987,N_8409,N_9474);
nor U17988 (N_17988,N_8357,N_11257);
xor U17989 (N_17989,N_10463,N_6888);
nand U17990 (N_17990,N_9445,N_7189);
or U17991 (N_17991,N_11980,N_11847);
or U17992 (N_17992,N_12037,N_9097);
or U17993 (N_17993,N_6707,N_10342);
or U17994 (N_17994,N_7974,N_9593);
nor U17995 (N_17995,N_6660,N_8583);
or U17996 (N_17996,N_7481,N_12414);
nand U17997 (N_17997,N_10817,N_6744);
xnor U17998 (N_17998,N_6574,N_12140);
nand U17999 (N_17999,N_11148,N_8632);
and U18000 (N_18000,N_10106,N_9230);
and U18001 (N_18001,N_6469,N_9475);
nor U18002 (N_18002,N_7897,N_12380);
nor U18003 (N_18003,N_9225,N_6631);
nand U18004 (N_18004,N_10803,N_7778);
nor U18005 (N_18005,N_9535,N_10329);
and U18006 (N_18006,N_9940,N_10425);
xor U18007 (N_18007,N_10361,N_11529);
or U18008 (N_18008,N_8451,N_7367);
or U18009 (N_18009,N_6964,N_10581);
and U18010 (N_18010,N_9178,N_6882);
nor U18011 (N_18011,N_7528,N_8352);
xor U18012 (N_18012,N_11861,N_9360);
or U18013 (N_18013,N_9940,N_11664);
or U18014 (N_18014,N_11197,N_12305);
nand U18015 (N_18015,N_7716,N_10770);
and U18016 (N_18016,N_7348,N_8717);
or U18017 (N_18017,N_10222,N_9669);
nor U18018 (N_18018,N_11798,N_10041);
nand U18019 (N_18019,N_8051,N_9485);
and U18020 (N_18020,N_7402,N_11362);
nor U18021 (N_18021,N_7435,N_6485);
xnor U18022 (N_18022,N_9508,N_11364);
nor U18023 (N_18023,N_10486,N_10960);
xor U18024 (N_18024,N_10007,N_8757);
nor U18025 (N_18025,N_11600,N_9222);
xor U18026 (N_18026,N_10164,N_9017);
nor U18027 (N_18027,N_7984,N_6805);
nor U18028 (N_18028,N_8012,N_12116);
nor U18029 (N_18029,N_10612,N_8401);
xnor U18030 (N_18030,N_7816,N_10961);
nand U18031 (N_18031,N_7246,N_11490);
nand U18032 (N_18032,N_8415,N_11917);
nand U18033 (N_18033,N_10355,N_9035);
xor U18034 (N_18034,N_8022,N_6548);
and U18035 (N_18035,N_9587,N_11732);
xor U18036 (N_18036,N_8202,N_7223);
and U18037 (N_18037,N_12240,N_6955);
nor U18038 (N_18038,N_12145,N_9806);
nor U18039 (N_18039,N_11631,N_11136);
nor U18040 (N_18040,N_10153,N_7180);
nand U18041 (N_18041,N_11451,N_9971);
nor U18042 (N_18042,N_11193,N_11769);
or U18043 (N_18043,N_9821,N_8074);
or U18044 (N_18044,N_10519,N_7955);
xor U18045 (N_18045,N_11606,N_7127);
xor U18046 (N_18046,N_6700,N_11766);
and U18047 (N_18047,N_11056,N_9996);
nand U18048 (N_18048,N_10348,N_8282);
xnor U18049 (N_18049,N_9221,N_6873);
nand U18050 (N_18050,N_9762,N_12468);
and U18051 (N_18051,N_11115,N_11977);
xnor U18052 (N_18052,N_6812,N_10534);
or U18053 (N_18053,N_8887,N_9820);
or U18054 (N_18054,N_10583,N_10350);
nor U18055 (N_18055,N_10666,N_9120);
and U18056 (N_18056,N_10021,N_12142);
or U18057 (N_18057,N_11464,N_11269);
nand U18058 (N_18058,N_9735,N_7384);
xnor U18059 (N_18059,N_8581,N_6946);
nor U18060 (N_18060,N_8475,N_10261);
nor U18061 (N_18061,N_7940,N_10157);
nor U18062 (N_18062,N_6944,N_10567);
nand U18063 (N_18063,N_8087,N_10938);
nand U18064 (N_18064,N_9924,N_10398);
and U18065 (N_18065,N_6859,N_7558);
nor U18066 (N_18066,N_7291,N_8354);
or U18067 (N_18067,N_9408,N_7632);
and U18068 (N_18068,N_12055,N_12057);
or U18069 (N_18069,N_9419,N_8959);
and U18070 (N_18070,N_8724,N_6899);
or U18071 (N_18071,N_9701,N_11946);
or U18072 (N_18072,N_8035,N_6877);
nor U18073 (N_18073,N_7670,N_11912);
xor U18074 (N_18074,N_7779,N_7604);
or U18075 (N_18075,N_11230,N_10832);
and U18076 (N_18076,N_9181,N_8313);
nor U18077 (N_18077,N_7336,N_8629);
nand U18078 (N_18078,N_8193,N_10463);
xnor U18079 (N_18079,N_11315,N_6734);
xor U18080 (N_18080,N_6536,N_7999);
xor U18081 (N_18081,N_9898,N_10889);
xnor U18082 (N_18082,N_11144,N_10285);
or U18083 (N_18083,N_8216,N_7692);
nand U18084 (N_18084,N_12081,N_7866);
nor U18085 (N_18085,N_7976,N_11950);
nor U18086 (N_18086,N_9907,N_10513);
xor U18087 (N_18087,N_11689,N_6581);
nor U18088 (N_18088,N_6546,N_7698);
xnor U18089 (N_18089,N_7400,N_8950);
or U18090 (N_18090,N_9131,N_7737);
xnor U18091 (N_18091,N_6412,N_9006);
nand U18092 (N_18092,N_11294,N_11878);
nor U18093 (N_18093,N_12233,N_6312);
xor U18094 (N_18094,N_11282,N_11106);
nand U18095 (N_18095,N_8186,N_11661);
nand U18096 (N_18096,N_9982,N_8349);
nor U18097 (N_18097,N_10524,N_9449);
or U18098 (N_18098,N_8142,N_12268);
xnor U18099 (N_18099,N_10870,N_8339);
xor U18100 (N_18100,N_11138,N_6884);
and U18101 (N_18101,N_11574,N_11495);
xnor U18102 (N_18102,N_8836,N_10845);
xor U18103 (N_18103,N_6346,N_8139);
and U18104 (N_18104,N_11110,N_10203);
nor U18105 (N_18105,N_10163,N_8667);
and U18106 (N_18106,N_11949,N_10068);
or U18107 (N_18107,N_10449,N_11435);
xnor U18108 (N_18108,N_9180,N_10981);
or U18109 (N_18109,N_7610,N_10830);
nand U18110 (N_18110,N_9885,N_8136);
nor U18111 (N_18111,N_12049,N_10230);
or U18112 (N_18112,N_6767,N_6613);
nor U18113 (N_18113,N_12328,N_7289);
xor U18114 (N_18114,N_10379,N_11074);
xor U18115 (N_18115,N_7595,N_7803);
nand U18116 (N_18116,N_9113,N_11109);
and U18117 (N_18117,N_10874,N_7567);
or U18118 (N_18118,N_9487,N_6421);
and U18119 (N_18119,N_6828,N_6391);
nor U18120 (N_18120,N_8911,N_12467);
nand U18121 (N_18121,N_10676,N_8759);
or U18122 (N_18122,N_8290,N_12340);
and U18123 (N_18123,N_9612,N_8410);
xnor U18124 (N_18124,N_8188,N_8754);
or U18125 (N_18125,N_7498,N_12244);
nand U18126 (N_18126,N_10434,N_10444);
nand U18127 (N_18127,N_12445,N_9996);
xor U18128 (N_18128,N_10092,N_7206);
xor U18129 (N_18129,N_10045,N_11033);
or U18130 (N_18130,N_11076,N_8666);
and U18131 (N_18131,N_6334,N_12081);
and U18132 (N_18132,N_7308,N_12407);
and U18133 (N_18133,N_12328,N_7143);
nand U18134 (N_18134,N_8739,N_10756);
xor U18135 (N_18135,N_10287,N_10963);
nand U18136 (N_18136,N_9652,N_9707);
and U18137 (N_18137,N_7077,N_9057);
and U18138 (N_18138,N_7863,N_9371);
and U18139 (N_18139,N_6460,N_11196);
nand U18140 (N_18140,N_12202,N_7840);
and U18141 (N_18141,N_11728,N_9497);
xnor U18142 (N_18142,N_6812,N_11890);
xor U18143 (N_18143,N_8401,N_6638);
nand U18144 (N_18144,N_6908,N_8299);
and U18145 (N_18145,N_8647,N_10958);
or U18146 (N_18146,N_8249,N_9755);
nand U18147 (N_18147,N_11726,N_9273);
nand U18148 (N_18148,N_8975,N_9678);
or U18149 (N_18149,N_11260,N_11819);
nor U18150 (N_18150,N_11943,N_12181);
xnor U18151 (N_18151,N_9315,N_10378);
nor U18152 (N_18152,N_10838,N_11023);
xor U18153 (N_18153,N_10920,N_10144);
nor U18154 (N_18154,N_9858,N_9981);
xnor U18155 (N_18155,N_10530,N_9559);
and U18156 (N_18156,N_10119,N_7104);
or U18157 (N_18157,N_11711,N_8108);
nand U18158 (N_18158,N_6357,N_10437);
or U18159 (N_18159,N_8196,N_11805);
nand U18160 (N_18160,N_9495,N_10063);
or U18161 (N_18161,N_12478,N_12110);
or U18162 (N_18162,N_10732,N_9556);
nor U18163 (N_18163,N_7534,N_11787);
or U18164 (N_18164,N_10010,N_6430);
and U18165 (N_18165,N_9853,N_11013);
and U18166 (N_18166,N_8172,N_8347);
nor U18167 (N_18167,N_12015,N_11613);
nand U18168 (N_18168,N_6570,N_7978);
xnor U18169 (N_18169,N_9029,N_6612);
and U18170 (N_18170,N_8573,N_9636);
nand U18171 (N_18171,N_6393,N_7834);
or U18172 (N_18172,N_11388,N_10450);
or U18173 (N_18173,N_10568,N_10714);
and U18174 (N_18174,N_10066,N_9289);
nand U18175 (N_18175,N_10048,N_10016);
and U18176 (N_18176,N_10694,N_7043);
nor U18177 (N_18177,N_8715,N_9537);
and U18178 (N_18178,N_9127,N_11388);
or U18179 (N_18179,N_8386,N_9591);
nor U18180 (N_18180,N_11786,N_10543);
or U18181 (N_18181,N_11246,N_7681);
xnor U18182 (N_18182,N_7417,N_12498);
nor U18183 (N_18183,N_10231,N_7304);
xor U18184 (N_18184,N_11895,N_8839);
or U18185 (N_18185,N_6497,N_9145);
nor U18186 (N_18186,N_9780,N_9686);
nand U18187 (N_18187,N_6852,N_8465);
nor U18188 (N_18188,N_6781,N_12359);
xor U18189 (N_18189,N_9568,N_9501);
xor U18190 (N_18190,N_7177,N_9769);
nor U18191 (N_18191,N_7237,N_12245);
nor U18192 (N_18192,N_11812,N_7441);
or U18193 (N_18193,N_9642,N_10463);
or U18194 (N_18194,N_11117,N_6956);
and U18195 (N_18195,N_9931,N_11314);
or U18196 (N_18196,N_9519,N_7675);
xnor U18197 (N_18197,N_8218,N_11516);
nor U18198 (N_18198,N_8997,N_7046);
or U18199 (N_18199,N_8811,N_12474);
nand U18200 (N_18200,N_9128,N_6722);
or U18201 (N_18201,N_10991,N_8912);
or U18202 (N_18202,N_9474,N_9215);
nor U18203 (N_18203,N_8741,N_12449);
or U18204 (N_18204,N_9519,N_11829);
nand U18205 (N_18205,N_9583,N_12375);
xnor U18206 (N_18206,N_11846,N_10834);
xor U18207 (N_18207,N_8332,N_10684);
and U18208 (N_18208,N_9922,N_11187);
nor U18209 (N_18209,N_8521,N_7101);
nand U18210 (N_18210,N_10130,N_11726);
or U18211 (N_18211,N_8099,N_9125);
nor U18212 (N_18212,N_10037,N_7654);
xor U18213 (N_18213,N_10136,N_6410);
xnor U18214 (N_18214,N_10697,N_7012);
or U18215 (N_18215,N_10195,N_6936);
nand U18216 (N_18216,N_10028,N_11746);
nand U18217 (N_18217,N_10908,N_8982);
or U18218 (N_18218,N_6963,N_7781);
nand U18219 (N_18219,N_6430,N_6928);
nand U18220 (N_18220,N_12320,N_12392);
nand U18221 (N_18221,N_7442,N_12019);
nand U18222 (N_18222,N_6391,N_11518);
and U18223 (N_18223,N_6467,N_7764);
nor U18224 (N_18224,N_7323,N_7487);
and U18225 (N_18225,N_11992,N_8979);
or U18226 (N_18226,N_6364,N_11368);
nand U18227 (N_18227,N_9504,N_6749);
nor U18228 (N_18228,N_8654,N_10428);
nand U18229 (N_18229,N_8468,N_8680);
nand U18230 (N_18230,N_10175,N_11701);
and U18231 (N_18231,N_8722,N_10034);
and U18232 (N_18232,N_11472,N_7230);
nor U18233 (N_18233,N_6251,N_6305);
and U18234 (N_18234,N_8481,N_8580);
and U18235 (N_18235,N_7718,N_6787);
and U18236 (N_18236,N_7226,N_11646);
xnor U18237 (N_18237,N_8069,N_8916);
or U18238 (N_18238,N_10429,N_8616);
or U18239 (N_18239,N_9045,N_7265);
nand U18240 (N_18240,N_10864,N_6504);
nor U18241 (N_18241,N_8982,N_8356);
and U18242 (N_18242,N_8665,N_6591);
xor U18243 (N_18243,N_6522,N_7981);
or U18244 (N_18244,N_8208,N_8668);
nor U18245 (N_18245,N_12130,N_10974);
xor U18246 (N_18246,N_7812,N_6552);
or U18247 (N_18247,N_9631,N_9603);
xnor U18248 (N_18248,N_9731,N_9783);
nand U18249 (N_18249,N_9582,N_10544);
nor U18250 (N_18250,N_6559,N_12281);
or U18251 (N_18251,N_8428,N_7926);
and U18252 (N_18252,N_8324,N_8897);
nor U18253 (N_18253,N_9364,N_8873);
nand U18254 (N_18254,N_10538,N_9857);
xor U18255 (N_18255,N_10804,N_6965);
nand U18256 (N_18256,N_9728,N_11015);
nor U18257 (N_18257,N_8055,N_12481);
or U18258 (N_18258,N_10569,N_7634);
xnor U18259 (N_18259,N_11673,N_6416);
nand U18260 (N_18260,N_8709,N_6569);
or U18261 (N_18261,N_10688,N_12074);
nor U18262 (N_18262,N_8524,N_10110);
and U18263 (N_18263,N_10635,N_10878);
xnor U18264 (N_18264,N_12447,N_12376);
nand U18265 (N_18265,N_9240,N_8910);
or U18266 (N_18266,N_10235,N_6359);
and U18267 (N_18267,N_10404,N_12451);
nand U18268 (N_18268,N_6577,N_12077);
nand U18269 (N_18269,N_9231,N_10162);
nor U18270 (N_18270,N_8885,N_12354);
nor U18271 (N_18271,N_10599,N_6811);
or U18272 (N_18272,N_8171,N_12010);
nor U18273 (N_18273,N_8613,N_11968);
xor U18274 (N_18274,N_6332,N_7433);
or U18275 (N_18275,N_8758,N_11362);
nand U18276 (N_18276,N_10713,N_12152);
xnor U18277 (N_18277,N_7456,N_10670);
nand U18278 (N_18278,N_11592,N_12449);
or U18279 (N_18279,N_7634,N_7249);
nand U18280 (N_18280,N_9420,N_10953);
nand U18281 (N_18281,N_6637,N_10402);
nand U18282 (N_18282,N_8345,N_10663);
nand U18283 (N_18283,N_12115,N_10429);
xor U18284 (N_18284,N_10822,N_8128);
nor U18285 (N_18285,N_8866,N_7441);
xor U18286 (N_18286,N_6963,N_8194);
xor U18287 (N_18287,N_7177,N_11131);
xor U18288 (N_18288,N_12189,N_7181);
nand U18289 (N_18289,N_6849,N_10967);
or U18290 (N_18290,N_9271,N_10620);
or U18291 (N_18291,N_11107,N_7964);
or U18292 (N_18292,N_11978,N_11975);
xnor U18293 (N_18293,N_7953,N_10458);
and U18294 (N_18294,N_10473,N_7725);
nand U18295 (N_18295,N_10299,N_6746);
xor U18296 (N_18296,N_8004,N_6568);
and U18297 (N_18297,N_6326,N_9222);
and U18298 (N_18298,N_10350,N_6843);
nand U18299 (N_18299,N_8087,N_12469);
or U18300 (N_18300,N_9037,N_6719);
nand U18301 (N_18301,N_7819,N_11851);
nand U18302 (N_18302,N_6261,N_10926);
nand U18303 (N_18303,N_11347,N_9672);
or U18304 (N_18304,N_6592,N_10220);
nor U18305 (N_18305,N_10300,N_6355);
nand U18306 (N_18306,N_6652,N_7062);
xor U18307 (N_18307,N_7351,N_7643);
xor U18308 (N_18308,N_12433,N_7754);
xnor U18309 (N_18309,N_6625,N_8116);
nor U18310 (N_18310,N_10790,N_6787);
nand U18311 (N_18311,N_6732,N_7136);
nand U18312 (N_18312,N_8919,N_8751);
nor U18313 (N_18313,N_10393,N_8436);
and U18314 (N_18314,N_7614,N_7835);
xnor U18315 (N_18315,N_8918,N_8396);
or U18316 (N_18316,N_8511,N_11358);
nand U18317 (N_18317,N_11457,N_9802);
or U18318 (N_18318,N_6473,N_9106);
nor U18319 (N_18319,N_7245,N_7788);
nor U18320 (N_18320,N_9045,N_6628);
and U18321 (N_18321,N_10598,N_11064);
nor U18322 (N_18322,N_11964,N_8971);
xor U18323 (N_18323,N_6833,N_11645);
nand U18324 (N_18324,N_9818,N_7893);
nor U18325 (N_18325,N_7853,N_10154);
nand U18326 (N_18326,N_6412,N_11179);
nor U18327 (N_18327,N_9138,N_6470);
or U18328 (N_18328,N_7233,N_10205);
xnor U18329 (N_18329,N_8912,N_8422);
and U18330 (N_18330,N_6474,N_10382);
or U18331 (N_18331,N_7540,N_11143);
or U18332 (N_18332,N_11759,N_10788);
and U18333 (N_18333,N_12366,N_10548);
and U18334 (N_18334,N_6260,N_7206);
and U18335 (N_18335,N_8656,N_10847);
nor U18336 (N_18336,N_11122,N_8269);
or U18337 (N_18337,N_9390,N_9486);
and U18338 (N_18338,N_6352,N_8010);
xnor U18339 (N_18339,N_9081,N_11024);
xor U18340 (N_18340,N_8681,N_6805);
nor U18341 (N_18341,N_9856,N_10700);
xor U18342 (N_18342,N_11604,N_8442);
and U18343 (N_18343,N_9350,N_11447);
nand U18344 (N_18344,N_8517,N_7583);
nand U18345 (N_18345,N_11396,N_10971);
or U18346 (N_18346,N_8773,N_12098);
nor U18347 (N_18347,N_9311,N_6565);
or U18348 (N_18348,N_11052,N_10245);
and U18349 (N_18349,N_9531,N_10624);
nand U18350 (N_18350,N_9063,N_10732);
xnor U18351 (N_18351,N_12293,N_7294);
or U18352 (N_18352,N_8126,N_10464);
xnor U18353 (N_18353,N_11602,N_8099);
nor U18354 (N_18354,N_8018,N_11098);
xor U18355 (N_18355,N_6330,N_10090);
nand U18356 (N_18356,N_10225,N_9077);
nor U18357 (N_18357,N_9613,N_9914);
nor U18358 (N_18358,N_7854,N_9129);
or U18359 (N_18359,N_8797,N_9330);
nand U18360 (N_18360,N_8595,N_11429);
or U18361 (N_18361,N_6923,N_10751);
and U18362 (N_18362,N_7907,N_8958);
xnor U18363 (N_18363,N_10298,N_8935);
nand U18364 (N_18364,N_7176,N_9369);
xor U18365 (N_18365,N_6775,N_11529);
nand U18366 (N_18366,N_9616,N_11972);
xor U18367 (N_18367,N_8254,N_7291);
xnor U18368 (N_18368,N_10464,N_7266);
nor U18369 (N_18369,N_11133,N_11598);
or U18370 (N_18370,N_11377,N_10377);
or U18371 (N_18371,N_8271,N_8923);
nor U18372 (N_18372,N_12175,N_8499);
or U18373 (N_18373,N_7012,N_8377);
and U18374 (N_18374,N_8871,N_12322);
xor U18375 (N_18375,N_6496,N_8290);
xor U18376 (N_18376,N_10787,N_10799);
and U18377 (N_18377,N_11766,N_6513);
and U18378 (N_18378,N_9439,N_7534);
or U18379 (N_18379,N_6384,N_8301);
nor U18380 (N_18380,N_10915,N_6486);
xor U18381 (N_18381,N_10205,N_7805);
or U18382 (N_18382,N_10007,N_11674);
nor U18383 (N_18383,N_11205,N_8156);
xnor U18384 (N_18384,N_7771,N_7722);
or U18385 (N_18385,N_11788,N_10499);
nor U18386 (N_18386,N_7140,N_11364);
xnor U18387 (N_18387,N_7131,N_10646);
nand U18388 (N_18388,N_9920,N_9978);
xnor U18389 (N_18389,N_10689,N_7211);
and U18390 (N_18390,N_10440,N_9661);
xnor U18391 (N_18391,N_9416,N_12021);
xor U18392 (N_18392,N_7530,N_7159);
nor U18393 (N_18393,N_8375,N_9841);
nand U18394 (N_18394,N_12184,N_7587);
and U18395 (N_18395,N_12030,N_11214);
xnor U18396 (N_18396,N_6763,N_6502);
nor U18397 (N_18397,N_9697,N_11200);
xnor U18398 (N_18398,N_12005,N_9166);
or U18399 (N_18399,N_7549,N_12297);
nor U18400 (N_18400,N_7304,N_7627);
and U18401 (N_18401,N_8521,N_8287);
or U18402 (N_18402,N_11810,N_6906);
xnor U18403 (N_18403,N_7551,N_10074);
or U18404 (N_18404,N_12151,N_9463);
nand U18405 (N_18405,N_8911,N_7810);
or U18406 (N_18406,N_6401,N_11343);
nand U18407 (N_18407,N_9310,N_12377);
and U18408 (N_18408,N_10288,N_11502);
and U18409 (N_18409,N_9838,N_11372);
and U18410 (N_18410,N_11511,N_9831);
and U18411 (N_18411,N_11248,N_6466);
or U18412 (N_18412,N_7343,N_7773);
or U18413 (N_18413,N_12497,N_12110);
nor U18414 (N_18414,N_10922,N_9623);
xnor U18415 (N_18415,N_7665,N_6601);
or U18416 (N_18416,N_7741,N_10888);
or U18417 (N_18417,N_8648,N_7117);
xor U18418 (N_18418,N_6683,N_12187);
nand U18419 (N_18419,N_11129,N_7124);
and U18420 (N_18420,N_6871,N_6941);
nor U18421 (N_18421,N_6568,N_6454);
xor U18422 (N_18422,N_10656,N_8789);
and U18423 (N_18423,N_7198,N_7151);
or U18424 (N_18424,N_10402,N_10966);
nor U18425 (N_18425,N_9179,N_8680);
or U18426 (N_18426,N_6783,N_8636);
xnor U18427 (N_18427,N_9029,N_7630);
xnor U18428 (N_18428,N_10885,N_7901);
or U18429 (N_18429,N_9908,N_10622);
nor U18430 (N_18430,N_11856,N_8141);
nand U18431 (N_18431,N_7762,N_9301);
or U18432 (N_18432,N_7709,N_6787);
nand U18433 (N_18433,N_11334,N_7338);
or U18434 (N_18434,N_8930,N_11249);
nand U18435 (N_18435,N_7043,N_8759);
nor U18436 (N_18436,N_11276,N_6907);
xor U18437 (N_18437,N_9506,N_7818);
nand U18438 (N_18438,N_11254,N_8251);
xnor U18439 (N_18439,N_9440,N_6990);
nor U18440 (N_18440,N_8833,N_9190);
or U18441 (N_18441,N_6664,N_11885);
xor U18442 (N_18442,N_8799,N_9907);
or U18443 (N_18443,N_7585,N_11517);
or U18444 (N_18444,N_11731,N_7800);
xnor U18445 (N_18445,N_12460,N_9760);
nand U18446 (N_18446,N_7899,N_11102);
nor U18447 (N_18447,N_9296,N_12376);
and U18448 (N_18448,N_9685,N_9008);
nor U18449 (N_18449,N_7322,N_8065);
or U18450 (N_18450,N_9946,N_7818);
nand U18451 (N_18451,N_10572,N_7233);
nor U18452 (N_18452,N_8984,N_7232);
or U18453 (N_18453,N_11456,N_8020);
nand U18454 (N_18454,N_10648,N_8392);
nor U18455 (N_18455,N_6643,N_6280);
or U18456 (N_18456,N_8429,N_8830);
xor U18457 (N_18457,N_7590,N_11927);
and U18458 (N_18458,N_11169,N_12144);
and U18459 (N_18459,N_11578,N_9135);
and U18460 (N_18460,N_9386,N_8100);
nand U18461 (N_18461,N_7812,N_9011);
nor U18462 (N_18462,N_12222,N_11212);
nor U18463 (N_18463,N_9305,N_9261);
or U18464 (N_18464,N_9768,N_9751);
or U18465 (N_18465,N_7906,N_7892);
and U18466 (N_18466,N_11835,N_8467);
or U18467 (N_18467,N_7376,N_9640);
and U18468 (N_18468,N_9159,N_10128);
xnor U18469 (N_18469,N_8450,N_8533);
nor U18470 (N_18470,N_11599,N_8279);
nand U18471 (N_18471,N_12368,N_7764);
nor U18472 (N_18472,N_11876,N_7847);
and U18473 (N_18473,N_10793,N_9808);
xnor U18474 (N_18474,N_9439,N_11782);
xor U18475 (N_18475,N_10502,N_10618);
and U18476 (N_18476,N_10155,N_7314);
xor U18477 (N_18477,N_10580,N_11607);
and U18478 (N_18478,N_10186,N_6262);
nor U18479 (N_18479,N_7806,N_7152);
and U18480 (N_18480,N_12314,N_9193);
nor U18481 (N_18481,N_6691,N_9671);
nor U18482 (N_18482,N_7579,N_8945);
nand U18483 (N_18483,N_9303,N_10398);
xnor U18484 (N_18484,N_8893,N_9773);
nor U18485 (N_18485,N_10901,N_6276);
xor U18486 (N_18486,N_7250,N_8922);
nand U18487 (N_18487,N_8083,N_11263);
or U18488 (N_18488,N_6346,N_7435);
nor U18489 (N_18489,N_8743,N_11516);
or U18490 (N_18490,N_12453,N_10686);
or U18491 (N_18491,N_9324,N_7171);
xnor U18492 (N_18492,N_7969,N_6836);
nand U18493 (N_18493,N_11271,N_7930);
nor U18494 (N_18494,N_7765,N_11277);
nand U18495 (N_18495,N_12079,N_9362);
nand U18496 (N_18496,N_11992,N_9052);
or U18497 (N_18497,N_11870,N_6736);
and U18498 (N_18498,N_6924,N_8152);
xnor U18499 (N_18499,N_7592,N_11364);
and U18500 (N_18500,N_6898,N_6610);
nor U18501 (N_18501,N_10951,N_8364);
nand U18502 (N_18502,N_9565,N_7735);
and U18503 (N_18503,N_12406,N_6653);
nor U18504 (N_18504,N_12168,N_11949);
and U18505 (N_18505,N_7293,N_9669);
nor U18506 (N_18506,N_7387,N_9381);
nor U18507 (N_18507,N_8212,N_9160);
nand U18508 (N_18508,N_10827,N_6673);
or U18509 (N_18509,N_7996,N_11507);
xor U18510 (N_18510,N_6879,N_10141);
nand U18511 (N_18511,N_8316,N_8239);
xnor U18512 (N_18512,N_11136,N_7936);
nor U18513 (N_18513,N_9001,N_7071);
and U18514 (N_18514,N_6281,N_11408);
nor U18515 (N_18515,N_12047,N_7294);
nor U18516 (N_18516,N_7525,N_12056);
and U18517 (N_18517,N_12386,N_12042);
nand U18518 (N_18518,N_10077,N_8366);
nand U18519 (N_18519,N_6483,N_6519);
nand U18520 (N_18520,N_8425,N_9015);
nand U18521 (N_18521,N_8890,N_6966);
nand U18522 (N_18522,N_12006,N_6315);
nor U18523 (N_18523,N_9978,N_8332);
and U18524 (N_18524,N_7877,N_8238);
or U18525 (N_18525,N_7411,N_11783);
xnor U18526 (N_18526,N_7897,N_7136);
xor U18527 (N_18527,N_9297,N_10783);
nor U18528 (N_18528,N_8239,N_9163);
and U18529 (N_18529,N_9197,N_11071);
nand U18530 (N_18530,N_10375,N_10009);
and U18531 (N_18531,N_9597,N_10283);
and U18532 (N_18532,N_10227,N_11450);
nand U18533 (N_18533,N_7315,N_6648);
or U18534 (N_18534,N_10840,N_9613);
nand U18535 (N_18535,N_11305,N_10594);
or U18536 (N_18536,N_6554,N_6834);
nor U18537 (N_18537,N_9834,N_8180);
xor U18538 (N_18538,N_7048,N_11028);
or U18539 (N_18539,N_8822,N_10172);
nand U18540 (N_18540,N_7335,N_12100);
nor U18541 (N_18541,N_6594,N_7600);
or U18542 (N_18542,N_6317,N_10212);
or U18543 (N_18543,N_7060,N_11928);
nand U18544 (N_18544,N_12264,N_9430);
and U18545 (N_18545,N_10759,N_10262);
xnor U18546 (N_18546,N_10412,N_7348);
nor U18547 (N_18547,N_9309,N_7541);
xnor U18548 (N_18548,N_7882,N_8905);
nor U18549 (N_18549,N_12114,N_8012);
xor U18550 (N_18550,N_11223,N_6935);
xnor U18551 (N_18551,N_10035,N_11533);
or U18552 (N_18552,N_6889,N_9170);
nand U18553 (N_18553,N_11556,N_7097);
and U18554 (N_18554,N_9463,N_9702);
nor U18555 (N_18555,N_10374,N_11143);
nor U18556 (N_18556,N_6604,N_10639);
nor U18557 (N_18557,N_8217,N_7603);
nand U18558 (N_18558,N_7480,N_9593);
or U18559 (N_18559,N_12498,N_8525);
nor U18560 (N_18560,N_8435,N_8429);
xor U18561 (N_18561,N_10754,N_10261);
and U18562 (N_18562,N_8349,N_8826);
or U18563 (N_18563,N_9892,N_7447);
or U18564 (N_18564,N_10200,N_11611);
and U18565 (N_18565,N_11915,N_10130);
nor U18566 (N_18566,N_8421,N_12339);
nor U18567 (N_18567,N_9172,N_7889);
nand U18568 (N_18568,N_8699,N_9206);
and U18569 (N_18569,N_11285,N_10318);
xnor U18570 (N_18570,N_10596,N_11364);
and U18571 (N_18571,N_7841,N_6645);
nand U18572 (N_18572,N_10465,N_11695);
and U18573 (N_18573,N_12264,N_12249);
xor U18574 (N_18574,N_8487,N_11364);
xor U18575 (N_18575,N_12234,N_11977);
nor U18576 (N_18576,N_7941,N_7602);
nand U18577 (N_18577,N_6907,N_8144);
and U18578 (N_18578,N_11163,N_10675);
or U18579 (N_18579,N_9729,N_6305);
and U18580 (N_18580,N_11454,N_8461);
xnor U18581 (N_18581,N_8179,N_10385);
nand U18582 (N_18582,N_10615,N_9643);
xor U18583 (N_18583,N_8630,N_11690);
nand U18584 (N_18584,N_9085,N_9465);
and U18585 (N_18585,N_6738,N_11657);
xnor U18586 (N_18586,N_10554,N_11446);
xnor U18587 (N_18587,N_9969,N_7109);
or U18588 (N_18588,N_10766,N_11424);
or U18589 (N_18589,N_7827,N_9466);
or U18590 (N_18590,N_9135,N_7823);
or U18591 (N_18591,N_9713,N_7534);
nor U18592 (N_18592,N_10983,N_10481);
and U18593 (N_18593,N_8556,N_7518);
nand U18594 (N_18594,N_11245,N_10263);
and U18595 (N_18595,N_6772,N_8107);
and U18596 (N_18596,N_7814,N_7414);
or U18597 (N_18597,N_10225,N_6264);
xnor U18598 (N_18598,N_9377,N_6560);
or U18599 (N_18599,N_10995,N_7982);
nor U18600 (N_18600,N_9904,N_11977);
nor U18601 (N_18601,N_11550,N_8729);
xor U18602 (N_18602,N_12226,N_10495);
nand U18603 (N_18603,N_11824,N_6251);
and U18604 (N_18604,N_8922,N_6470);
nand U18605 (N_18605,N_8932,N_9070);
nor U18606 (N_18606,N_8768,N_7278);
xor U18607 (N_18607,N_12384,N_9909);
or U18608 (N_18608,N_9053,N_7401);
nand U18609 (N_18609,N_7694,N_10635);
or U18610 (N_18610,N_6511,N_11215);
xor U18611 (N_18611,N_8791,N_11423);
nand U18612 (N_18612,N_8641,N_9717);
and U18613 (N_18613,N_10556,N_10991);
and U18614 (N_18614,N_11887,N_10895);
nand U18615 (N_18615,N_8920,N_6517);
and U18616 (N_18616,N_8736,N_9049);
nand U18617 (N_18617,N_8329,N_10407);
nor U18618 (N_18618,N_12160,N_10533);
xnor U18619 (N_18619,N_6661,N_6891);
or U18620 (N_18620,N_10558,N_11286);
or U18621 (N_18621,N_8808,N_6776);
or U18622 (N_18622,N_11745,N_10184);
or U18623 (N_18623,N_10571,N_9107);
and U18624 (N_18624,N_7360,N_8957);
nand U18625 (N_18625,N_6380,N_6442);
nor U18626 (N_18626,N_9114,N_12062);
nand U18627 (N_18627,N_6281,N_7735);
and U18628 (N_18628,N_11398,N_8419);
and U18629 (N_18629,N_9074,N_7703);
and U18630 (N_18630,N_11137,N_10262);
xor U18631 (N_18631,N_12443,N_6862);
xnor U18632 (N_18632,N_11569,N_10794);
or U18633 (N_18633,N_8770,N_9541);
nor U18634 (N_18634,N_6849,N_9684);
nand U18635 (N_18635,N_11078,N_9363);
nor U18636 (N_18636,N_11926,N_10560);
xnor U18637 (N_18637,N_6608,N_11723);
xor U18638 (N_18638,N_10151,N_8883);
nor U18639 (N_18639,N_9228,N_9879);
nand U18640 (N_18640,N_11923,N_7058);
xor U18641 (N_18641,N_6603,N_8456);
nand U18642 (N_18642,N_10239,N_10558);
nand U18643 (N_18643,N_11492,N_12083);
or U18644 (N_18644,N_9540,N_10541);
and U18645 (N_18645,N_11678,N_12056);
or U18646 (N_18646,N_11114,N_11952);
nand U18647 (N_18647,N_6429,N_8152);
and U18648 (N_18648,N_6432,N_9461);
nand U18649 (N_18649,N_7414,N_10768);
xnor U18650 (N_18650,N_10850,N_8446);
xor U18651 (N_18651,N_10563,N_7344);
or U18652 (N_18652,N_12055,N_11021);
or U18653 (N_18653,N_6671,N_9722);
nand U18654 (N_18654,N_6613,N_12079);
nor U18655 (N_18655,N_8599,N_6705);
or U18656 (N_18656,N_8221,N_8935);
or U18657 (N_18657,N_9273,N_8089);
or U18658 (N_18658,N_7481,N_9932);
or U18659 (N_18659,N_7346,N_9660);
or U18660 (N_18660,N_6317,N_10133);
nor U18661 (N_18661,N_9151,N_7759);
nor U18662 (N_18662,N_12231,N_10337);
and U18663 (N_18663,N_7694,N_12188);
or U18664 (N_18664,N_10735,N_8698);
and U18665 (N_18665,N_9157,N_11652);
nand U18666 (N_18666,N_6776,N_7659);
nand U18667 (N_18667,N_8542,N_11488);
nor U18668 (N_18668,N_7049,N_11652);
nand U18669 (N_18669,N_8946,N_10429);
or U18670 (N_18670,N_7267,N_7590);
nand U18671 (N_18671,N_7148,N_6973);
and U18672 (N_18672,N_9203,N_8130);
and U18673 (N_18673,N_7994,N_11011);
nor U18674 (N_18674,N_11625,N_10412);
nand U18675 (N_18675,N_11537,N_7252);
and U18676 (N_18676,N_6908,N_11313);
nand U18677 (N_18677,N_7450,N_11529);
nor U18678 (N_18678,N_11270,N_7837);
nand U18679 (N_18679,N_8344,N_10111);
nor U18680 (N_18680,N_9030,N_10023);
and U18681 (N_18681,N_9212,N_8297);
xnor U18682 (N_18682,N_7884,N_11813);
nand U18683 (N_18683,N_6792,N_9175);
nand U18684 (N_18684,N_7175,N_12268);
and U18685 (N_18685,N_8731,N_11457);
nor U18686 (N_18686,N_9693,N_11300);
nor U18687 (N_18687,N_11821,N_6696);
nand U18688 (N_18688,N_9996,N_11266);
nand U18689 (N_18689,N_9276,N_6662);
xnor U18690 (N_18690,N_11136,N_6343);
or U18691 (N_18691,N_8833,N_10750);
or U18692 (N_18692,N_12011,N_8461);
xor U18693 (N_18693,N_7746,N_11465);
xor U18694 (N_18694,N_12029,N_9884);
or U18695 (N_18695,N_10632,N_8589);
xnor U18696 (N_18696,N_7866,N_7983);
nand U18697 (N_18697,N_9653,N_11427);
and U18698 (N_18698,N_11082,N_10127);
xor U18699 (N_18699,N_8919,N_9149);
nor U18700 (N_18700,N_9777,N_7227);
and U18701 (N_18701,N_9623,N_11219);
and U18702 (N_18702,N_8425,N_10995);
xnor U18703 (N_18703,N_11107,N_8403);
and U18704 (N_18704,N_9846,N_12128);
xor U18705 (N_18705,N_10834,N_12075);
or U18706 (N_18706,N_12402,N_9684);
nand U18707 (N_18707,N_10111,N_7952);
nand U18708 (N_18708,N_7510,N_11141);
nor U18709 (N_18709,N_12407,N_8467);
nand U18710 (N_18710,N_7733,N_12164);
xor U18711 (N_18711,N_8834,N_7831);
xor U18712 (N_18712,N_7985,N_9523);
or U18713 (N_18713,N_10056,N_6806);
and U18714 (N_18714,N_7762,N_11633);
or U18715 (N_18715,N_6656,N_10237);
xor U18716 (N_18716,N_11215,N_9870);
or U18717 (N_18717,N_7640,N_10951);
nor U18718 (N_18718,N_9831,N_11888);
and U18719 (N_18719,N_6449,N_7370);
and U18720 (N_18720,N_7522,N_12135);
xor U18721 (N_18721,N_9289,N_10696);
nand U18722 (N_18722,N_11709,N_12488);
and U18723 (N_18723,N_11243,N_11203);
nand U18724 (N_18724,N_12186,N_10526);
nand U18725 (N_18725,N_11981,N_9749);
xor U18726 (N_18726,N_9050,N_7494);
and U18727 (N_18727,N_10167,N_11879);
or U18728 (N_18728,N_11992,N_11301);
and U18729 (N_18729,N_6423,N_12006);
nor U18730 (N_18730,N_12393,N_9177);
xor U18731 (N_18731,N_8483,N_9878);
nand U18732 (N_18732,N_6813,N_12479);
and U18733 (N_18733,N_11751,N_8755);
nand U18734 (N_18734,N_10790,N_8471);
nand U18735 (N_18735,N_9100,N_8780);
or U18736 (N_18736,N_11324,N_8626);
nor U18737 (N_18737,N_7588,N_7508);
or U18738 (N_18738,N_11777,N_9073);
nand U18739 (N_18739,N_8906,N_10556);
xnor U18740 (N_18740,N_7670,N_8459);
and U18741 (N_18741,N_6465,N_11588);
nor U18742 (N_18742,N_11714,N_8988);
and U18743 (N_18743,N_6637,N_6391);
or U18744 (N_18744,N_6836,N_12194);
nand U18745 (N_18745,N_7800,N_6471);
or U18746 (N_18746,N_6279,N_7390);
and U18747 (N_18747,N_12072,N_8068);
xor U18748 (N_18748,N_9077,N_7916);
nand U18749 (N_18749,N_9613,N_8378);
and U18750 (N_18750,N_15840,N_17786);
and U18751 (N_18751,N_17093,N_17319);
or U18752 (N_18752,N_14424,N_18182);
nand U18753 (N_18753,N_16838,N_17777);
and U18754 (N_18754,N_17069,N_14060);
nand U18755 (N_18755,N_15751,N_16654);
and U18756 (N_18756,N_14553,N_17809);
nand U18757 (N_18757,N_16632,N_14879);
xnor U18758 (N_18758,N_16096,N_16079);
and U18759 (N_18759,N_16401,N_13141);
or U18760 (N_18760,N_18520,N_12668);
and U18761 (N_18761,N_17680,N_17966);
and U18762 (N_18762,N_18496,N_18329);
or U18763 (N_18763,N_14741,N_15848);
nor U18764 (N_18764,N_18076,N_12836);
and U18765 (N_18765,N_13105,N_14167);
xnor U18766 (N_18766,N_14863,N_13727);
nand U18767 (N_18767,N_13953,N_12998);
xnor U18768 (N_18768,N_17372,N_13991);
nand U18769 (N_18769,N_12666,N_16695);
nand U18770 (N_18770,N_13114,N_16009);
or U18771 (N_18771,N_16068,N_18024);
or U18772 (N_18772,N_13169,N_17818);
nand U18773 (N_18773,N_12734,N_17737);
xnor U18774 (N_18774,N_18469,N_17018);
or U18775 (N_18775,N_18016,N_13485);
or U18776 (N_18776,N_15235,N_16550);
xor U18777 (N_18777,N_16679,N_13276);
nand U18778 (N_18778,N_14570,N_17105);
nand U18779 (N_18779,N_15243,N_15043);
or U18780 (N_18780,N_15306,N_15687);
or U18781 (N_18781,N_13340,N_13873);
or U18782 (N_18782,N_17104,N_15232);
xor U18783 (N_18783,N_18624,N_17147);
or U18784 (N_18784,N_14201,N_13206);
xnor U18785 (N_18785,N_17635,N_18162);
xor U18786 (N_18786,N_13997,N_17548);
nand U18787 (N_18787,N_16479,N_13531);
or U18788 (N_18788,N_18585,N_17206);
nor U18789 (N_18789,N_18159,N_16565);
xor U18790 (N_18790,N_14023,N_17977);
xor U18791 (N_18791,N_16081,N_15433);
nor U18792 (N_18792,N_13263,N_14439);
nand U18793 (N_18793,N_17914,N_15230);
or U18794 (N_18794,N_16849,N_15518);
nand U18795 (N_18795,N_15729,N_18261);
xor U18796 (N_18796,N_15620,N_18243);
or U18797 (N_18797,N_15271,N_12800);
or U18798 (N_18798,N_17456,N_18006);
nor U18799 (N_18799,N_15111,N_14667);
nor U18800 (N_18800,N_13603,N_16604);
and U18801 (N_18801,N_17858,N_13788);
and U18802 (N_18802,N_14003,N_16258);
nand U18803 (N_18803,N_16242,N_15185);
and U18804 (N_18804,N_16366,N_14441);
xnor U18805 (N_18805,N_16237,N_18687);
nor U18806 (N_18806,N_13190,N_18035);
nand U18807 (N_18807,N_17621,N_15430);
nor U18808 (N_18808,N_15570,N_16141);
xor U18809 (N_18809,N_14123,N_16508);
and U18810 (N_18810,N_14071,N_16014);
and U18811 (N_18811,N_17895,N_13745);
or U18812 (N_18812,N_14541,N_12948);
nor U18813 (N_18813,N_14674,N_14375);
or U18814 (N_18814,N_17435,N_12761);
nor U18815 (N_18815,N_17851,N_14015);
and U18816 (N_18816,N_18644,N_16888);
nor U18817 (N_18817,N_15238,N_13399);
nand U18818 (N_18818,N_15484,N_13082);
and U18819 (N_18819,N_14236,N_16767);
xor U18820 (N_18820,N_13125,N_17926);
nand U18821 (N_18821,N_16215,N_13995);
nor U18822 (N_18822,N_17587,N_12944);
and U18823 (N_18823,N_17763,N_15097);
and U18824 (N_18824,N_16563,N_12736);
or U18825 (N_18825,N_13471,N_14226);
nand U18826 (N_18826,N_15046,N_15593);
and U18827 (N_18827,N_14505,N_16688);
nor U18828 (N_18828,N_13884,N_14809);
and U18829 (N_18829,N_14630,N_14457);
nand U18830 (N_18830,N_18150,N_12595);
nand U18831 (N_18831,N_15019,N_12895);
nor U18832 (N_18832,N_17005,N_16245);
or U18833 (N_18833,N_16217,N_13560);
and U18834 (N_18834,N_12546,N_14550);
or U18835 (N_18835,N_15821,N_18032);
and U18836 (N_18836,N_15812,N_13961);
or U18837 (N_18837,N_15356,N_15252);
nor U18838 (N_18838,N_17611,N_16906);
nor U18839 (N_18839,N_13306,N_17986);
nor U18840 (N_18840,N_15437,N_13433);
nand U18841 (N_18841,N_14820,N_15837);
xor U18842 (N_18842,N_12722,N_17046);
nand U18843 (N_18843,N_14361,N_13047);
nand U18844 (N_18844,N_18555,N_12986);
nor U18845 (N_18845,N_17051,N_15688);
xnor U18846 (N_18846,N_15073,N_16641);
nand U18847 (N_18847,N_17111,N_15917);
and U18848 (N_18848,N_18093,N_13470);
nor U18849 (N_18849,N_17664,N_15063);
or U18850 (N_18850,N_15968,N_16647);
xor U18851 (N_18851,N_16620,N_17097);
or U18852 (N_18852,N_14240,N_15706);
xor U18853 (N_18853,N_15815,N_13481);
nor U18854 (N_18854,N_17506,N_13432);
and U18855 (N_18855,N_14971,N_14476);
nor U18856 (N_18856,N_16470,N_13930);
xor U18857 (N_18857,N_15052,N_15517);
xor U18858 (N_18858,N_15148,N_14908);
and U18859 (N_18859,N_14503,N_15014);
or U18860 (N_18860,N_13073,N_12773);
nand U18861 (N_18861,N_13784,N_14716);
nand U18862 (N_18862,N_14680,N_13015);
and U18863 (N_18863,N_17126,N_15739);
nand U18864 (N_18864,N_18417,N_16896);
xor U18865 (N_18865,N_14887,N_15948);
xor U18866 (N_18866,N_16182,N_17006);
nand U18867 (N_18867,N_18322,N_16640);
xnor U18868 (N_18868,N_16117,N_13006);
nand U18869 (N_18869,N_13680,N_14185);
or U18870 (N_18870,N_14335,N_16509);
and U18871 (N_18871,N_12712,N_18548);
and U18872 (N_18872,N_13748,N_17103);
and U18873 (N_18873,N_13061,N_15728);
xnor U18874 (N_18874,N_12762,N_17296);
nand U18875 (N_18875,N_15344,N_18107);
nor U18876 (N_18876,N_16843,N_13504);
xnor U18877 (N_18877,N_13024,N_15126);
and U18878 (N_18878,N_15548,N_13708);
xor U18879 (N_18879,N_18245,N_14431);
xor U18880 (N_18880,N_13529,N_17203);
xnor U18881 (N_18881,N_17642,N_16124);
nor U18882 (N_18882,N_16286,N_13809);
nor U18883 (N_18883,N_12933,N_14601);
xnor U18884 (N_18884,N_13076,N_16898);
and U18885 (N_18885,N_17637,N_12534);
or U18886 (N_18886,N_17640,N_15464);
xor U18887 (N_18887,N_17466,N_14992);
xnor U18888 (N_18888,N_14493,N_14684);
or U18889 (N_18889,N_14610,N_13608);
nand U18890 (N_18890,N_14398,N_16073);
and U18891 (N_18891,N_12821,N_17188);
nand U18892 (N_18892,N_14477,N_15256);
nand U18893 (N_18893,N_13167,N_18034);
xnor U18894 (N_18894,N_18257,N_18675);
nand U18895 (N_18895,N_15236,N_15583);
nor U18896 (N_18896,N_16492,N_18022);
or U18897 (N_18897,N_18726,N_17474);
nor U18898 (N_18898,N_18229,N_16092);
and U18899 (N_18899,N_13418,N_16530);
nand U18900 (N_18900,N_15267,N_13746);
xnor U18901 (N_18901,N_14462,N_12618);
nand U18902 (N_18902,N_16965,N_15684);
and U18903 (N_18903,N_12807,N_13844);
nor U18904 (N_18904,N_17359,N_16078);
nor U18905 (N_18905,N_17565,N_15847);
or U18906 (N_18906,N_15836,N_14665);
nand U18907 (N_18907,N_16744,N_15530);
nand U18908 (N_18908,N_16210,N_15114);
or U18909 (N_18909,N_14107,N_13028);
xnor U18910 (N_18910,N_15979,N_18449);
or U18911 (N_18911,N_16507,N_14738);
or U18912 (N_18912,N_14347,N_15928);
or U18913 (N_18913,N_16814,N_16760);
nor U18914 (N_18914,N_16300,N_16815);
or U18915 (N_18915,N_17911,N_14872);
nor U18916 (N_18916,N_18226,N_13630);
or U18917 (N_18917,N_13092,N_13403);
nand U18918 (N_18918,N_13508,N_18693);
or U18919 (N_18919,N_14289,N_17865);
and U18920 (N_18920,N_15598,N_12901);
xor U18921 (N_18921,N_14877,N_16728);
nor U18922 (N_18922,N_17861,N_17526);
nand U18923 (N_18923,N_15206,N_15782);
and U18924 (N_18924,N_13657,N_13696);
or U18925 (N_18925,N_17318,N_15479);
and U18926 (N_18926,N_16047,N_14425);
and U18927 (N_18927,N_12662,N_17017);
and U18928 (N_18928,N_13888,N_15218);
nand U18929 (N_18929,N_17461,N_16336);
or U18930 (N_18930,N_14899,N_15402);
xor U18931 (N_18931,N_12567,N_16209);
and U18932 (N_18932,N_12679,N_16428);
nor U18933 (N_18933,N_15958,N_12760);
and U18934 (N_18934,N_12920,N_16069);
or U18935 (N_18935,N_17504,N_15446);
nor U18936 (N_18936,N_18542,N_14752);
nor U18937 (N_18937,N_16091,N_16072);
and U18938 (N_18938,N_17146,N_17703);
nor U18939 (N_18939,N_13863,N_13720);
or U18940 (N_18940,N_13257,N_18321);
nand U18941 (N_18941,N_17509,N_13450);
nand U18942 (N_18942,N_14718,N_12506);
and U18943 (N_18943,N_12687,N_16955);
nor U18944 (N_18944,N_14765,N_13240);
xor U18945 (N_18945,N_15285,N_12932);
nor U18946 (N_18946,N_15577,N_15042);
and U18947 (N_18947,N_15559,N_15784);
or U18948 (N_18948,N_16880,N_14987);
or U18949 (N_18949,N_14701,N_18036);
nor U18950 (N_18950,N_14170,N_17169);
or U18951 (N_18951,N_14244,N_17328);
xnor U18952 (N_18952,N_17238,N_15299);
xor U18953 (N_18953,N_13520,N_13402);
or U18954 (N_18954,N_17756,N_14896);
or U18955 (N_18955,N_16846,N_14266);
or U18956 (N_18956,N_16134,N_16518);
xnor U18957 (N_18957,N_15427,N_12768);
nor U18958 (N_18958,N_15108,N_14836);
nand U18959 (N_18959,N_13145,N_16235);
xnor U18960 (N_18960,N_16425,N_16155);
and U18961 (N_18961,N_15936,N_14782);
nand U18962 (N_18962,N_12779,N_16720);
and U18963 (N_18963,N_16189,N_15867);
or U18964 (N_18964,N_16875,N_16927);
nand U18965 (N_18965,N_13133,N_17262);
or U18966 (N_18966,N_14970,N_18495);
xnor U18967 (N_18967,N_13049,N_14504);
nand U18968 (N_18968,N_16146,N_17837);
and U18969 (N_18969,N_17876,N_14543);
xnor U18970 (N_18970,N_14581,N_15735);
xnor U18971 (N_18971,N_13713,N_16510);
and U18972 (N_18972,N_17370,N_14306);
nand U18973 (N_18973,N_14233,N_16032);
nor U18974 (N_18974,N_14161,N_16414);
nor U18975 (N_18975,N_16471,N_16982);
xor U18976 (N_18976,N_18552,N_17915);
xor U18977 (N_18977,N_12623,N_13463);
nand U18978 (N_18978,N_17698,N_14039);
nor U18979 (N_18979,N_16163,N_13139);
and U18980 (N_18980,N_15254,N_16973);
nor U18981 (N_18981,N_15322,N_13147);
nand U18982 (N_18982,N_16388,N_14898);
nor U18983 (N_18983,N_14303,N_13187);
xnor U18984 (N_18984,N_14006,N_15803);
or U18985 (N_18985,N_18130,N_14978);
nor U18986 (N_18986,N_18152,N_15138);
and U18987 (N_18987,N_15745,N_17313);
nor U18988 (N_18988,N_14077,N_15002);
or U18989 (N_18989,N_14612,N_13093);
or U18990 (N_18990,N_15279,N_14824);
nor U18991 (N_18991,N_14184,N_15830);
xor U18992 (N_18992,N_18031,N_17622);
nor U18993 (N_18993,N_13118,N_15793);
or U18994 (N_18994,N_16709,N_13699);
xor U18995 (N_18995,N_14400,N_14745);
nand U18996 (N_18996,N_18330,N_12995);
or U18997 (N_18997,N_13044,N_18201);
xor U18998 (N_18998,N_15513,N_14996);
nor U18999 (N_18999,N_14090,N_13786);
nand U19000 (N_19000,N_15631,N_12811);
and U19001 (N_19001,N_14265,N_18060);
nor U19002 (N_19002,N_18025,N_15152);
xnor U19003 (N_19003,N_16132,N_13434);
or U19004 (N_19004,N_15970,N_14203);
nand U19005 (N_19005,N_17508,N_15511);
xor U19006 (N_19006,N_16944,N_15333);
nand U19007 (N_19007,N_12574,N_15417);
or U19008 (N_19008,N_12974,N_15089);
and U19009 (N_19009,N_15361,N_17213);
nand U19010 (N_19010,N_13327,N_14239);
nand U19011 (N_19011,N_13641,N_13212);
nor U19012 (N_19012,N_12796,N_14685);
and U19013 (N_19013,N_15656,N_13950);
or U19014 (N_19014,N_16299,N_17128);
and U19015 (N_19015,N_12825,N_17862);
or U19016 (N_19016,N_12514,N_18611);
and U19017 (N_19017,N_16349,N_15181);
xor U19018 (N_19018,N_16523,N_14479);
nor U19019 (N_19019,N_16756,N_17430);
nor U19020 (N_19020,N_13666,N_15457);
nor U19021 (N_19021,N_13328,N_16658);
and U19022 (N_19022,N_18214,N_14276);
xnor U19023 (N_19023,N_17360,N_15671);
nor U19024 (N_19024,N_18559,N_13527);
xnor U19025 (N_19025,N_14731,N_16522);
nor U19026 (N_19026,N_15494,N_16588);
xnor U19027 (N_19027,N_13298,N_16030);
and U19028 (N_19028,N_12544,N_13495);
nand U19029 (N_19029,N_16517,N_14029);
or U19030 (N_19030,N_15365,N_13837);
or U19031 (N_19031,N_14713,N_13106);
xnor U19032 (N_19032,N_18311,N_16467);
nor U19033 (N_19033,N_13894,N_13429);
and U19034 (N_19034,N_16040,N_12660);
nor U19035 (N_19035,N_14911,N_17157);
xor U19036 (N_19036,N_13038,N_18317);
or U19037 (N_19037,N_18018,N_17588);
nand U19038 (N_19038,N_13782,N_12577);
nor U19039 (N_19039,N_12717,N_18085);
nor U19040 (N_19040,N_14960,N_14366);
and U19041 (N_19041,N_12648,N_14677);
xnor U19042 (N_19042,N_16437,N_17249);
xor U19043 (N_19043,N_17714,N_17473);
nand U19044 (N_19044,N_13494,N_17905);
nor U19045 (N_19045,N_17218,N_17530);
xnor U19046 (N_19046,N_16084,N_15297);
nand U19047 (N_19047,N_14914,N_14257);
nor U19048 (N_19048,N_16120,N_14604);
and U19049 (N_19049,N_12581,N_15696);
nand U19050 (N_19050,N_14147,N_15032);
or U19051 (N_19051,N_13408,N_16034);
and U19052 (N_19052,N_16956,N_17729);
and U19053 (N_19053,N_15217,N_15080);
nor U19054 (N_19054,N_15198,N_15748);
and U19055 (N_19055,N_16244,N_15959);
xor U19056 (N_19056,N_16177,N_16703);
nand U19057 (N_19057,N_15887,N_13893);
and U19058 (N_19058,N_16558,N_15145);
and U19059 (N_19059,N_14654,N_16232);
nand U19060 (N_19060,N_15119,N_18683);
or U19061 (N_19061,N_14949,N_13668);
and U19062 (N_19062,N_17358,N_18728);
and U19063 (N_19063,N_15594,N_13763);
xor U19064 (N_19064,N_17779,N_16998);
nand U19065 (N_19065,N_18220,N_16332);
nor U19066 (N_19066,N_18462,N_14330);
and U19067 (N_19067,N_16308,N_12670);
xor U19068 (N_19068,N_14251,N_12904);
and U19069 (N_19069,N_16468,N_15225);
xnor U19070 (N_19070,N_16741,N_17919);
and U19071 (N_19071,N_12755,N_13659);
xor U19072 (N_19072,N_15208,N_14825);
nor U19073 (N_19073,N_15421,N_18471);
nor U19074 (N_19074,N_15794,N_16478);
and U19075 (N_19075,N_13921,N_18425);
xnor U19076 (N_19076,N_13820,N_14946);
or U19077 (N_19077,N_17833,N_17750);
nand U19078 (N_19078,N_13663,N_15955);
or U19079 (N_19079,N_18474,N_16983);
or U19080 (N_19080,N_15618,N_12624);
or U19081 (N_19081,N_15930,N_18454);
and U19082 (N_19082,N_18702,N_15429);
nand U19083 (N_19083,N_15122,N_13737);
or U19084 (N_19084,N_16905,N_12777);
xnor U19085 (N_19085,N_13008,N_13739);
xor U19086 (N_19086,N_14297,N_15658);
or U19087 (N_19087,N_12798,N_18446);
nand U19088 (N_19088,N_14332,N_14501);
and U19089 (N_19089,N_15186,N_18593);
nand U19090 (N_19090,N_14806,N_15143);
nand U19091 (N_19091,N_13021,N_15645);
or U19092 (N_19092,N_16891,N_14428);
and U19093 (N_19093,N_16823,N_14129);
nand U19094 (N_19094,N_12806,N_18394);
nand U19095 (N_19095,N_13319,N_13389);
nand U19096 (N_19096,N_18731,N_16502);
nand U19097 (N_19097,N_15015,N_14430);
and U19098 (N_19098,N_15331,N_14865);
nand U19099 (N_19099,N_17037,N_18406);
xor U19100 (N_19100,N_17382,N_16455);
xor U19101 (N_19101,N_14611,N_16036);
nor U19102 (N_19102,N_16088,N_13036);
nand U19103 (N_19103,N_17364,N_12885);
xor U19104 (N_19104,N_14108,N_16037);
or U19105 (N_19105,N_16020,N_15025);
xnor U19106 (N_19106,N_14281,N_16580);
nand U19107 (N_19107,N_12523,N_16740);
nand U19108 (N_19108,N_13261,N_13564);
or U19109 (N_19109,N_17476,N_17271);
or U19110 (N_19110,N_13152,N_13312);
xnor U19111 (N_19111,N_17971,N_15180);
or U19112 (N_19112,N_18529,N_15519);
and U19113 (N_19113,N_18364,N_16923);
or U19114 (N_19114,N_12831,N_12621);
or U19115 (N_19115,N_14407,N_15506);
or U19116 (N_19116,N_14418,N_13417);
or U19117 (N_19117,N_18197,N_14056);
and U19118 (N_19118,N_16249,N_16024);
nand U19119 (N_19119,N_13381,N_13906);
nand U19120 (N_19120,N_17056,N_15453);
xor U19121 (N_19121,N_12820,N_16175);
nand U19122 (N_19122,N_18275,N_15661);
xor U19123 (N_19123,N_15280,N_15632);
nor U19124 (N_19124,N_13168,N_12958);
nor U19125 (N_19125,N_13524,N_16298);
nand U19126 (N_19126,N_16243,N_17590);
or U19127 (N_19127,N_17736,N_13670);
nand U19128 (N_19128,N_17492,N_17990);
nand U19129 (N_19129,N_18480,N_13774);
nor U19130 (N_19130,N_14054,N_16190);
and U19131 (N_19131,N_17502,N_16592);
xor U19132 (N_19132,N_17092,N_16737);
xor U19133 (N_19133,N_18013,N_17802);
and U19134 (N_19134,N_17404,N_18352);
nand U19135 (N_19135,N_13819,N_15284);
or U19136 (N_19136,N_16352,N_13395);
xor U19137 (N_19137,N_15375,N_12969);
nor U19138 (N_19138,N_14443,N_14302);
nor U19139 (N_19139,N_16745,N_16748);
and U19140 (N_19140,N_17280,N_16197);
xor U19141 (N_19141,N_16104,N_16464);
nor U19142 (N_19142,N_16960,N_17518);
and U19143 (N_19143,N_16600,N_12602);
or U19144 (N_19144,N_15991,N_16852);
and U19145 (N_19145,N_16871,N_16701);
and U19146 (N_19146,N_14294,N_13215);
nand U19147 (N_19147,N_12586,N_15949);
nand U19148 (N_19148,N_14962,N_12803);
nand U19149 (N_19149,N_15229,N_16606);
nand U19150 (N_19150,N_13081,N_15068);
nor U19151 (N_19151,N_17609,N_18384);
xor U19152 (N_19152,N_14316,N_15578);
nor U19153 (N_19153,N_14647,N_14127);
or U19154 (N_19154,N_17302,N_14177);
nor U19155 (N_19155,N_16975,N_15714);
and U19156 (N_19156,N_15588,N_14285);
nor U19157 (N_19157,N_17574,N_13729);
and U19158 (N_19158,N_16279,N_13932);
and U19159 (N_19159,N_13363,N_14109);
xor U19160 (N_19160,N_16089,N_18716);
xnor U19161 (N_19161,N_12971,N_17131);
xor U19162 (N_19162,N_18273,N_16904);
and U19163 (N_19163,N_18569,N_14691);
xor U19164 (N_19164,N_13196,N_12559);
or U19165 (N_19165,N_17836,N_16706);
or U19166 (N_19166,N_13738,N_18522);
nor U19167 (N_19167,N_15546,N_17731);
or U19168 (N_19168,N_12810,N_17045);
nand U19169 (N_19169,N_17931,N_17434);
nand U19170 (N_19170,N_13959,N_16276);
xnor U19171 (N_19171,N_12614,N_14644);
xor U19172 (N_19172,N_13568,N_17568);
and U19173 (N_19173,N_14307,N_18099);
nand U19174 (N_19174,N_14811,N_13525);
and U19175 (N_19175,N_14900,N_13791);
xnor U19176 (N_19176,N_17171,N_13839);
xor U19177 (N_19177,N_14846,N_17482);
xnor U19178 (N_19178,N_14510,N_17228);
or U19179 (N_19179,N_18707,N_12645);
and U19180 (N_19180,N_18416,N_18077);
or U19181 (N_19181,N_13929,N_16553);
xnor U19182 (N_19182,N_15873,N_16556);
nor U19183 (N_19183,N_13996,N_17490);
or U19184 (N_19184,N_13326,N_15493);
xnor U19185 (N_19185,N_18238,N_14508);
nor U19186 (N_19186,N_16650,N_15312);
nand U19187 (N_19187,N_15483,N_13732);
xor U19188 (N_19188,N_15157,N_13980);
or U19189 (N_19189,N_15293,N_13194);
xnor U19190 (N_19190,N_14867,N_15844);
xnor U19191 (N_19191,N_13755,N_16685);
xnor U19192 (N_19192,N_16666,N_14044);
nand U19193 (N_19193,N_17689,N_14920);
and U19194 (N_19194,N_15387,N_18249);
xnor U19195 (N_19195,N_12770,N_18211);
xor U19196 (N_19196,N_15458,N_16793);
nand U19197 (N_19197,N_16689,N_14246);
nor U19198 (N_19198,N_13886,N_17969);
xor U19199 (N_19199,N_16821,N_13679);
or U19200 (N_19200,N_15298,N_15366);
or U19201 (N_19201,N_15767,N_15600);
nand U19202 (N_19202,N_13468,N_16221);
nand U19203 (N_19203,N_17438,N_16946);
nand U19204 (N_19204,N_12695,N_18266);
nor U19205 (N_19205,N_12612,N_17282);
nand U19206 (N_19206,N_13626,N_15807);
or U19207 (N_19207,N_13437,N_13370);
and U19208 (N_19208,N_18524,N_12700);
and U19209 (N_19209,N_18540,N_16489);
xor U19210 (N_19210,N_18483,N_17278);
xnor U19211 (N_19211,N_13658,N_16344);
xor U19212 (N_19212,N_14173,N_14864);
nand U19213 (N_19213,N_14277,N_16067);
and U19214 (N_19214,N_16594,N_13155);
nor U19215 (N_19215,N_16044,N_15159);
nor U19216 (N_19216,N_14641,N_16306);
and U19217 (N_19217,N_15395,N_17335);
and U19218 (N_19218,N_15286,N_17952);
nor U19219 (N_19219,N_16534,N_15726);
xor U19220 (N_19220,N_15731,N_18344);
nor U19221 (N_19221,N_13225,N_14059);
xnor U19222 (N_19222,N_16951,N_13834);
nand U19223 (N_19223,N_17344,N_17399);
or U19224 (N_19224,N_15529,N_16984);
nand U19225 (N_19225,N_17844,N_18127);
nor U19226 (N_19226,N_12951,N_12788);
xor U19227 (N_19227,N_14858,N_18043);
nor U19228 (N_19228,N_13349,N_15076);
and U19229 (N_19229,N_15248,N_16870);
nand U19230 (N_19230,N_13831,N_17657);
nor U19231 (N_19231,N_17822,N_14165);
or U19232 (N_19232,N_17804,N_16377);
nand U19233 (N_19233,N_12869,N_14926);
xnor U19234 (N_19234,N_18608,N_14102);
nor U19235 (N_19235,N_18456,N_16704);
xnor U19236 (N_19236,N_13054,N_17405);
xnor U19237 (N_19237,N_17726,N_16656);
xor U19238 (N_19238,N_15859,N_13271);
xor U19239 (N_19239,N_17770,N_13661);
xor U19240 (N_19240,N_18413,N_17260);
nand U19241 (N_19241,N_18375,N_17783);
and U19242 (N_19242,N_17348,N_17088);
xnor U19243 (N_19243,N_16811,N_15537);
or U19244 (N_19244,N_13273,N_18461);
and U19245 (N_19245,N_14878,N_18408);
and U19246 (N_19246,N_14582,N_13002);
nor U19247 (N_19247,N_16976,N_14989);
xnor U19248 (N_19248,N_16813,N_17628);
nand U19249 (N_19249,N_16928,N_14256);
nand U19250 (N_19250,N_16648,N_18388);
and U19251 (N_19251,N_15674,N_18641);
and U19252 (N_19252,N_14781,N_15700);
and U19253 (N_19253,N_17057,N_18662);
xor U19254 (N_19254,N_15151,N_13416);
and U19255 (N_19255,N_16261,N_14817);
and U19256 (N_19256,N_18534,N_16251);
xnor U19257 (N_19257,N_12947,N_17441);
or U19258 (N_19258,N_17384,N_17566);
nor U19259 (N_19259,N_14459,N_16736);
nor U19260 (N_19260,N_14725,N_13704);
nor U19261 (N_19261,N_17699,N_14859);
nand U19262 (N_19262,N_17553,N_16433);
and U19263 (N_19263,N_15353,N_15061);
and U19264 (N_19264,N_14934,N_12686);
and U19265 (N_19265,N_18195,N_17350);
or U19266 (N_19266,N_18103,N_16697);
nor U19267 (N_19267,N_18360,N_18105);
and U19268 (N_19268,N_18227,N_17402);
nor U19269 (N_19269,N_16103,N_16564);
and U19270 (N_19270,N_14771,N_15103);
xnor U19271 (N_19271,N_14755,N_17541);
or U19272 (N_19272,N_12654,N_13643);
or U19273 (N_19273,N_18224,N_15792);
nor U19274 (N_19274,N_17042,N_12929);
nor U19275 (N_19275,N_13011,N_14881);
xnor U19276 (N_19276,N_17788,N_13892);
and U19277 (N_19277,N_13549,N_12797);
nor U19278 (N_19278,N_17572,N_14097);
nor U19279 (N_19279,N_17082,N_15553);
nand U19280 (N_19280,N_16605,N_18289);
or U19281 (N_19281,N_14670,N_14942);
xnor U19282 (N_19282,N_13461,N_17838);
or U19283 (N_19283,N_15326,N_13052);
nor U19284 (N_19284,N_14888,N_12889);
and U19285 (N_19285,N_13935,N_14464);
xor U19286 (N_19286,N_16790,N_13513);
xor U19287 (N_19287,N_12804,N_12667);
xnor U19288 (N_19288,N_13390,N_15200);
nor U19289 (N_19289,N_14822,N_13369);
or U19290 (N_19290,N_13760,N_15099);
or U19291 (N_19291,N_18636,N_13224);
nand U19292 (N_19292,N_14134,N_14437);
nand U19293 (N_19293,N_16143,N_17667);
and U19294 (N_19294,N_18473,N_13592);
and U19295 (N_19295,N_14954,N_13401);
and U19296 (N_19296,N_15443,N_14828);
nor U19297 (N_19297,N_14195,N_15734);
nor U19298 (N_19298,N_16419,N_15644);
nand U19299 (N_19299,N_13157,N_17101);
nor U19300 (N_19300,N_18096,N_14319);
xor U19301 (N_19301,N_12517,N_15370);
and U19302 (N_19302,N_15343,N_16486);
nor U19303 (N_19303,N_14043,N_15263);
or U19304 (N_19304,N_14795,N_12740);
nand U19305 (N_19305,N_17728,N_15819);
and U19306 (N_19306,N_18027,N_17314);
nand U19307 (N_19307,N_16841,N_16183);
nor U19308 (N_19308,N_18572,N_16561);
or U19309 (N_19309,N_15635,N_13664);
and U19310 (N_19310,N_16546,N_14968);
nand U19311 (N_19311,N_13104,N_15999);
or U19312 (N_19312,N_14176,N_15246);
and U19313 (N_19313,N_13778,N_12794);
nand U19314 (N_19314,N_16739,N_17850);
nand U19315 (N_19315,N_15095,N_16885);
or U19316 (N_19316,N_15678,N_15045);
or U19317 (N_19317,N_12547,N_12500);
or U19318 (N_19318,N_16797,N_13158);
and U19319 (N_19319,N_18650,N_14166);
nor U19320 (N_19320,N_17383,N_14948);
nor U19321 (N_19321,N_18686,N_17880);
nor U19322 (N_19322,N_17646,N_17484);
and U19323 (N_19323,N_15934,N_13936);
nand U19324 (N_19324,N_13260,N_12742);
and U19325 (N_19325,N_17874,N_12688);
nor U19326 (N_19326,N_17415,N_13796);
or U19327 (N_19327,N_16268,N_17178);
xnor U19328 (N_19328,N_18042,N_16466);
or U19329 (N_19329,N_17711,N_15222);
and U19330 (N_19330,N_13986,N_13459);
or U19331 (N_19331,N_13631,N_15829);
xor U19332 (N_19332,N_14310,N_17747);
nand U19333 (N_19333,N_18690,N_16528);
and U19334 (N_19334,N_17007,N_17825);
nor U19335 (N_19335,N_16651,N_18114);
or U19336 (N_19336,N_15897,N_14341);
and U19337 (N_19337,N_17197,N_16917);
or U19338 (N_19338,N_15691,N_15137);
nand U19339 (N_19339,N_16262,N_13719);
xor U19340 (N_19340,N_18165,N_17960);
and U19341 (N_19341,N_15923,N_16584);
nor U19342 (N_19342,N_13323,N_16363);
nor U19343 (N_19343,N_14120,N_13540);
and U19344 (N_19344,N_18251,N_12950);
or U19345 (N_19345,N_15879,N_17710);
and U19346 (N_19346,N_14579,N_16614);
and U19347 (N_19347,N_13101,N_18260);
nand U19348 (N_19348,N_13779,N_12968);
nand U19349 (N_19349,N_18685,N_18326);
xnor U19350 (N_19350,N_15313,N_18663);
xnor U19351 (N_19351,N_17613,N_18654);
xnor U19352 (N_19352,N_15701,N_15462);
nor U19353 (N_19353,N_17935,N_14144);
or U19354 (N_19354,N_13602,N_12721);
and U19355 (N_19355,N_17240,N_12630);
or U19356 (N_19356,N_14608,N_13069);
nor U19357 (N_19357,N_18286,N_17424);
or U19358 (N_19358,N_16005,N_14370);
or U19359 (N_19359,N_14305,N_16342);
xnor U19360 (N_19360,N_16293,N_18597);
and U19361 (N_19361,N_17653,N_13171);
xor U19362 (N_19362,N_16461,N_18270);
nand U19363 (N_19363,N_12819,N_12626);
nand U19364 (N_19364,N_17661,N_18639);
or U19365 (N_19365,N_13348,N_17062);
or U19366 (N_19366,N_14769,N_15787);
and U19367 (N_19367,N_16660,N_13456);
and U19368 (N_19368,N_13136,N_13574);
and U19369 (N_19369,N_16201,N_14522);
and U19370 (N_19370,N_17472,N_14729);
and U19371 (N_19371,N_12542,N_13415);
and U19372 (N_19372,N_14849,N_18359);
or U19373 (N_19373,N_15178,N_17380);
and U19374 (N_19374,N_12940,N_14288);
and U19375 (N_19375,N_13955,N_14287);
or U19376 (N_19376,N_15692,N_14599);
nor U19377 (N_19377,N_15708,N_17894);
nor U19378 (N_19378,N_17321,N_16400);
xnor U19379 (N_19379,N_13304,N_13046);
nand U19380 (N_19380,N_17170,N_12661);
nand U19381 (N_19381,N_13259,N_13222);
and U19382 (N_19382,N_17885,N_16150);
nor U19383 (N_19383,N_15841,N_18598);
or U19384 (N_19384,N_14221,N_13770);
nand U19385 (N_19385,N_17365,N_14512);
or U19386 (N_19386,N_15287,N_18711);
xor U19387 (N_19387,N_14636,N_16351);
and U19388 (N_19388,N_14453,N_13575);
or U19389 (N_19389,N_15386,N_18297);
nand U19390 (N_19390,N_15850,N_17958);
and U19391 (N_19391,N_18710,N_13130);
or U19392 (N_19392,N_18614,N_13301);
nor U19393 (N_19393,N_14214,N_13938);
nand U19394 (N_19394,N_13126,N_14063);
and U19395 (N_19395,N_14497,N_16252);
nand U19396 (N_19396,N_13102,N_12750);
or U19397 (N_19397,N_13464,N_14249);
or U19398 (N_19398,N_16586,N_17735);
nor U19399 (N_19399,N_14818,N_14035);
nor U19400 (N_19400,N_14019,N_15098);
nor U19401 (N_19401,N_16469,N_13411);
nand U19402 (N_19402,N_14548,N_14928);
and U19403 (N_19403,N_13963,N_15191);
xnor U19404 (N_19404,N_14136,N_13164);
xor U19405 (N_19405,N_13579,N_16149);
xor U19406 (N_19406,N_17215,N_18506);
nor U19407 (N_19407,N_15391,N_13973);
and U19408 (N_19408,N_15962,N_13705);
or U19409 (N_19409,N_13067,N_17079);
nand U19410 (N_19410,N_17470,N_17923);
or U19411 (N_19411,N_16220,N_15189);
xnor U19412 (N_19412,N_12844,N_16882);
nor U19413 (N_19413,N_14478,N_17495);
xnor U19414 (N_19414,N_14363,N_15209);
and U19415 (N_19415,N_12813,N_15890);
and U19416 (N_19416,N_18622,N_13903);
nand U19417 (N_19417,N_16013,N_16002);
and U19418 (N_19418,N_15475,N_15115);
nor U19419 (N_19419,N_17925,N_16585);
nor U19420 (N_19420,N_17872,N_13230);
xor U19421 (N_19421,N_16962,N_15637);
or U19422 (N_19422,N_14135,N_14314);
nor U19423 (N_19423,N_13914,N_15935);
nor U19424 (N_19424,N_15907,N_17224);
nand U19425 (N_19425,N_12724,N_14979);
xor U19426 (N_19426,N_14835,N_14267);
xor U19427 (N_19427,N_14458,N_18267);
or U19428 (N_19428,N_12598,N_15590);
nor U19429 (N_19429,N_17841,N_16285);
and U19430 (N_19430,N_12997,N_13282);
xnor U19431 (N_19431,N_13889,N_12557);
or U19432 (N_19432,N_14923,N_16596);
and U19433 (N_19433,N_14767,N_13397);
nand U19434 (N_19434,N_14523,N_15822);
or U19435 (N_19435,N_17299,N_17853);
xor U19436 (N_19436,N_15039,N_13683);
nor U19437 (N_19437,N_15495,N_17189);
xor U19438 (N_19438,N_14432,N_18213);
nand U19439 (N_19439,N_17847,N_15811);
nor U19440 (N_19440,N_14391,N_16968);
nor U19441 (N_19441,N_17346,N_17706);
and U19442 (N_19442,N_16557,N_18280);
nand U19443 (N_19443,N_14095,N_18179);
and U19444 (N_19444,N_14245,N_13635);
nand U19445 (N_19445,N_15649,N_15900);
nand U19446 (N_19446,N_16116,N_14311);
nand U19447 (N_19447,N_12552,N_18349);
nor U19448 (N_19448,N_17368,N_14254);
nand U19449 (N_19449,N_16850,N_18504);
xor U19450 (N_19450,N_14619,N_12867);
nor U19451 (N_19451,N_15174,N_17610);
xnor U19452 (N_19452,N_15946,N_18479);
xnor U19453 (N_19453,N_13992,N_17546);
or U19454 (N_19454,N_18741,N_16909);
nand U19455 (N_19455,N_12701,N_14140);
nand U19456 (N_19456,N_12891,N_13232);
and U19457 (N_19457,N_15893,N_15166);
xor U19458 (N_19458,N_14365,N_15587);
and U19459 (N_19459,N_15489,N_14707);
or U19460 (N_19460,N_16953,N_17601);
xor U19461 (N_19461,N_15766,N_15033);
xor U19462 (N_19462,N_18231,N_16726);
nand U19463 (N_19463,N_15662,N_14931);
nand U19464 (N_19464,N_15158,N_13897);
nor U19465 (N_19465,N_16187,N_15888);
or U19466 (N_19466,N_13591,N_13290);
and U19467 (N_19467,N_14372,N_12886);
xnor U19468 (N_19468,N_14403,N_13785);
xor U19469 (N_19469,N_13129,N_13233);
nand U19470 (N_19470,N_17556,N_12590);
xnor U19471 (N_19471,N_16374,N_14852);
xnor U19472 (N_19472,N_16314,N_16538);
xnor U19473 (N_19473,N_12582,N_14350);
nor U19474 (N_19474,N_13536,N_17389);
nor U19475 (N_19475,N_14087,N_13887);
nand U19476 (N_19476,N_14150,N_14646);
and U19477 (N_19477,N_15008,N_12878);
xnor U19478 (N_19478,N_18205,N_16385);
nand U19479 (N_19479,N_15093,N_14255);
or U19480 (N_19480,N_14791,N_16246);
and U19481 (N_19481,N_13428,N_17050);
nor U19482 (N_19482,N_12587,N_18560);
or U19483 (N_19483,N_16458,N_17995);
and U19484 (N_19484,N_15663,N_17086);
nand U19485 (N_19485,N_12593,N_16499);
and U19486 (N_19486,N_18217,N_18183);
nor U19487 (N_19487,N_18334,N_14894);
nand U19488 (N_19488,N_18448,N_17676);
nand U19489 (N_19489,N_12890,N_17307);
xor U19490 (N_19490,N_14317,N_13469);
nand U19491 (N_19491,N_16749,N_13108);
or U19492 (N_19492,N_16435,N_16731);
nand U19493 (N_19493,N_18719,N_15013);
nor U19494 (N_19494,N_14761,N_13874);
or U19495 (N_19495,N_14146,N_17968);
xnor U19496 (N_19496,N_15965,N_12876);
nand U19497 (N_19497,N_13638,N_18578);
nand U19498 (N_19498,N_13615,N_14719);
and U19499 (N_19499,N_15491,N_14093);
xnor U19500 (N_19500,N_15736,N_16317);
and U19501 (N_19501,N_15278,N_13297);
xnor U19502 (N_19502,N_17581,N_17666);
xor U19503 (N_19503,N_16997,N_18324);
nand U19504 (N_19504,N_13858,N_16506);
or U19505 (N_19505,N_13341,N_13740);
nor U19506 (N_19506,N_18588,N_13912);
xnor U19507 (N_19507,N_12877,N_16178);
nor U19508 (N_19508,N_12503,N_16125);
nor U19509 (N_19509,N_18605,N_16274);
nor U19510 (N_19510,N_12650,N_16567);
nand U19511 (N_19511,N_13458,N_15981);
nor U19512 (N_19512,N_13879,N_13070);
nor U19513 (N_19513,N_15057,N_13681);
nor U19514 (N_19514,N_18065,N_14151);
or U19515 (N_19515,N_18119,N_15768);
nor U19516 (N_19516,N_13535,N_12738);
nor U19517 (N_19517,N_14525,N_14569);
xnor U19518 (N_19518,N_13596,N_14614);
xor U19519 (N_19519,N_14618,N_13042);
nand U19520 (N_19520,N_15969,N_18402);
nor U19521 (N_19521,N_17311,N_14890);
and U19522 (N_19522,N_14560,N_16828);
nand U19523 (N_19523,N_17882,N_17907);
and U19524 (N_19524,N_16281,N_13940);
and U19525 (N_19525,N_17266,N_18175);
xnor U19526 (N_19526,N_13115,N_15295);
nand U19527 (N_19527,N_16832,N_17252);
nand U19528 (N_19528,N_13578,N_17924);
xor U19529 (N_19529,N_13810,N_17810);
nand U19530 (N_19530,N_18430,N_16105);
nor U19531 (N_19531,N_14004,N_17532);
nor U19532 (N_19532,N_16136,N_17113);
and U19533 (N_19533,N_15857,N_17281);
and U19534 (N_19534,N_13515,N_15738);
and U19535 (N_19535,N_18445,N_16755);
nor U19536 (N_19536,N_18580,N_17663);
nand U19537 (N_19537,N_14377,N_13559);
or U19538 (N_19538,N_13751,N_13933);
and U19539 (N_19539,N_14955,N_16057);
nand U19540 (N_19540,N_18110,N_17643);
nor U19541 (N_19541,N_15608,N_15876);
nor U19542 (N_19542,N_15772,N_14066);
nor U19543 (N_19543,N_14111,N_18033);
nor U19544 (N_19544,N_15290,N_17649);
and U19545 (N_19545,N_13359,N_15301);
and U19546 (N_19546,N_15616,N_16196);
or U19547 (N_19547,N_12972,N_16788);
nor U19548 (N_19548,N_14356,N_14386);
and U19549 (N_19549,N_14325,N_12710);
or U19550 (N_19550,N_16061,N_18681);
and U19551 (N_19551,N_13012,N_16834);
and U19552 (N_19552,N_13045,N_17648);
nor U19553 (N_19553,N_14704,N_12791);
and U19554 (N_19554,N_17976,N_18295);
nor U19555 (N_19555,N_14784,N_17781);
or U19556 (N_19556,N_18594,N_18431);
and U19557 (N_19557,N_16277,N_16925);
nand U19558 (N_19558,N_16633,N_15694);
xor U19559 (N_19559,N_15504,N_17323);
nand U19560 (N_19560,N_13925,N_18678);
nor U19561 (N_19561,N_14532,N_18255);
nor U19562 (N_19562,N_14449,N_14779);
or U19563 (N_19563,N_15617,N_17595);
or U19564 (N_19564,N_14785,N_14104);
or U19565 (N_19565,N_13007,N_12729);
xor U19566 (N_19566,N_17469,N_13388);
nand U19567 (N_19567,N_13928,N_14149);
and U19568 (N_19568,N_18527,N_16354);
and U19569 (N_19569,N_17032,N_16610);
nor U19570 (N_19570,N_18166,N_18163);
nor U19571 (N_19571,N_12859,N_12528);
nor U19572 (N_19572,N_13112,N_17903);
or U19573 (N_19573,N_18237,N_14450);
nand U19574 (N_19574,N_17413,N_17496);
nor U19575 (N_19575,N_18008,N_15827);
or U19576 (N_19576,N_18482,N_17498);
nand U19577 (N_19577,N_17417,N_14735);
nor U19578 (N_19578,N_18230,N_17896);
or U19579 (N_19579,N_13019,N_13336);
or U19580 (N_19580,N_12509,N_15994);
xor U19581 (N_19581,N_12706,N_17927);
and U19582 (N_19582,N_15425,N_14230);
or U19583 (N_19583,N_18399,N_13414);
or U19584 (N_19584,N_15374,N_14540);
and U19585 (N_19585,N_15054,N_14326);
xnor U19586 (N_19586,N_13993,N_13354);
or U19587 (N_19587,N_13474,N_13802);
or U19588 (N_19588,N_16664,N_15780);
nor U19589 (N_19589,N_18320,N_16514);
xnor U19590 (N_19590,N_15078,N_15394);
nand U19591 (N_19591,N_14885,N_15455);
nand U19592 (N_19592,N_17343,N_13448);
or U19593 (N_19593,N_15021,N_18185);
or U19594 (N_19594,N_14295,N_18368);
and U19595 (N_19595,N_15802,N_17125);
nor U19596 (N_19596,N_13072,N_13211);
xnor U19597 (N_19597,N_18634,N_17257);
xor U19598 (N_19598,N_15535,N_18523);
and U19599 (N_19599,N_13677,N_15652);
xor U19600 (N_19600,N_17899,N_17038);
nor U19601 (N_19601,N_12815,N_14848);
or U19602 (N_19602,N_18673,N_18133);
nand U19603 (N_19603,N_14435,N_15693);
or U19604 (N_19604,N_15665,N_13371);
or U19605 (N_19605,N_17164,N_13454);
nor U19606 (N_19606,N_12651,N_15340);
or U19607 (N_19607,N_14966,N_16853);
nor U19608 (N_19608,N_12862,N_15964);
or U19609 (N_19609,N_15851,N_13913);
xor U19610 (N_19610,N_17583,N_15749);
nand U19611 (N_19611,N_17563,N_17080);
and U19612 (N_19612,N_14855,N_14279);
xnor U19613 (N_19613,N_15001,N_16240);
and U19614 (N_19614,N_17870,N_17087);
xnor U19615 (N_19615,N_16520,N_13573);
and U19616 (N_19616,N_18549,N_13812);
nor U19617 (N_19617,N_18064,N_13446);
nand U19618 (N_19618,N_17599,N_18351);
xnor U19619 (N_19619,N_16874,N_13096);
xnor U19620 (N_19620,N_16952,N_17377);
nor U19621 (N_19621,N_18184,N_16348);
or U19622 (N_19622,N_18298,N_17964);
and U19623 (N_19623,N_16153,N_15654);
xnor U19624 (N_19624,N_12603,N_17805);
or U19625 (N_19625,N_17690,N_17668);
nand U19626 (N_19626,N_16250,N_16899);
or U19627 (N_19627,N_13207,N_13922);
or U19628 (N_19628,N_13647,N_14841);
nor U19629 (N_19629,N_13043,N_17725);
xor U19630 (N_19630,N_16082,N_15554);
nor U19631 (N_19631,N_15711,N_12771);
xor U19632 (N_19632,N_16436,N_13697);
or U19633 (N_19633,N_18629,N_18571);
nor U19634 (N_19634,N_12580,N_17800);
and U19635 (N_19635,N_13835,N_16933);
and U19636 (N_19636,N_13709,N_18432);
or U19637 (N_19637,N_15788,N_16599);
or U19638 (N_19638,N_17855,N_14892);
or U19639 (N_19639,N_15630,N_15846);
nand U19640 (N_19640,N_15354,N_12718);
or U19641 (N_19641,N_12531,N_13733);
and U19642 (N_19642,N_15419,N_15234);
nand U19643 (N_19643,N_15627,N_14645);
xnor U19644 (N_19644,N_14024,N_17945);
nand U19645 (N_19645,N_14264,N_14426);
xor U19646 (N_19646,N_16048,N_18029);
and U19647 (N_19647,N_12977,N_16533);
nand U19648 (N_19648,N_16996,N_18308);
nand U19649 (N_19649,N_14470,N_13182);
and U19650 (N_19650,N_16087,N_18403);
and U19651 (N_19651,N_13173,N_18228);
nand U19652 (N_19652,N_18082,N_14814);
nor U19653 (N_19653,N_16859,N_17427);
nand U19654 (N_19654,N_14536,N_16759);
nor U19655 (N_19655,N_18513,N_16423);
or U19656 (N_19656,N_14652,N_13789);
nor U19657 (N_19657,N_15149,N_18073);
and U19658 (N_19658,N_17798,N_18037);
and U19659 (N_19659,N_15562,N_15120);
nand U19660 (N_19660,N_17806,N_15384);
nor U19661 (N_19661,N_16413,N_15607);
nand U19662 (N_19662,N_13055,N_15539);
xor U19663 (N_19663,N_13688,N_12516);
nand U19664 (N_19664,N_18083,N_12824);
and U19665 (N_19665,N_17273,N_15336);
and U19666 (N_19666,N_15373,N_17808);
nand U19667 (N_19667,N_16802,N_15385);
nand U19668 (N_19668,N_17759,N_17001);
xor U19669 (N_19669,N_15170,N_14686);
or U19670 (N_19670,N_15150,N_15393);
xnor U19671 (N_19671,N_13964,N_13116);
and U19672 (N_19672,N_13761,N_12591);
or U19673 (N_19673,N_15109,N_16929);
xor U19674 (N_19674,N_17720,N_13945);
and U19675 (N_19675,N_15129,N_15592);
and U19676 (N_19676,N_18465,N_16108);
and U19677 (N_19677,N_15797,N_15398);
xor U19678 (N_19678,N_12837,N_13752);
or U19679 (N_19679,N_12583,N_14743);
or U19680 (N_19680,N_18007,N_15029);
nand U19681 (N_19681,N_16054,N_14062);
nor U19682 (N_19682,N_15785,N_14554);
nand U19683 (N_19683,N_13840,N_15503);
nor U19684 (N_19684,N_16411,N_16683);
and U19685 (N_19685,N_14301,N_17602);
nor U19686 (N_19686,N_17204,N_16806);
nor U19687 (N_19687,N_17608,N_18003);
or U19688 (N_19688,N_13821,N_14629);
nor U19689 (N_19689,N_18747,N_17366);
xnor U19690 (N_19690,N_16851,N_18058);
nor U19691 (N_19691,N_17701,N_12953);
nand U19692 (N_19692,N_16026,N_16548);
xor U19693 (N_19693,N_12606,N_13287);
or U19694 (N_19694,N_17109,N_17791);
or U19695 (N_19695,N_17332,N_18434);
or U19696 (N_19696,N_15016,N_18088);
xor U19697 (N_19697,N_15709,N_14296);
and U19698 (N_19698,N_18285,N_13451);
and U19699 (N_19699,N_17219,N_16330);
nor U19700 (N_19700,N_17451,N_13965);
and U19701 (N_19701,N_16058,N_16675);
and U19702 (N_19702,N_17177,N_15144);
and U19703 (N_19703,N_15899,N_12549);
and U19704 (N_19704,N_15834,N_15622);
nand U19705 (N_19705,N_16051,N_12505);
nand U19706 (N_19706,N_17558,N_16776);
xor U19707 (N_19707,N_16617,N_12954);
or U19708 (N_19708,N_18709,N_16707);
xnor U19709 (N_19709,N_16635,N_13501);
or U19710 (N_19710,N_13804,N_13662);
nand U19711 (N_19711,N_18044,N_15752);
xnor U19712 (N_19712,N_13510,N_15156);
xnor U19713 (N_19713,N_16979,N_14880);
nor U19714 (N_19714,N_15468,N_17091);
nand U19715 (N_19715,N_13216,N_13714);
nand U19716 (N_19716,N_15947,N_17235);
nand U19717 (N_19717,N_18137,N_14770);
or U19718 (N_19718,N_15030,N_17349);
nor U19719 (N_19719,N_17153,N_17898);
or U19720 (N_19720,N_13877,N_18011);
nor U19721 (N_19721,N_13756,N_16004);
or U19722 (N_19722,N_14596,N_17181);
xnor U19723 (N_19723,N_16536,N_16901);
or U19724 (N_19724,N_13780,N_12880);
or U19725 (N_19725,N_14530,N_13057);
and U19726 (N_19726,N_14145,N_13178);
or U19727 (N_19727,N_13907,N_14857);
and U19728 (N_19728,N_16970,N_12960);
or U19729 (N_19729,N_16000,N_13827);
nand U19730 (N_19730,N_13333,N_13503);
nand U19731 (N_19731,N_12748,N_12672);
xnor U19732 (N_19732,N_14475,N_14633);
nand U19733 (N_19733,N_17021,N_12918);
or U19734 (N_19734,N_18341,N_12521);
nand U19735 (N_19735,N_18092,N_18475);
nor U19736 (N_19736,N_14001,N_14247);
xor U19737 (N_19737,N_15912,N_14988);
nor U19738 (N_19738,N_18147,N_15308);
xnor U19739 (N_19739,N_14706,N_12747);
nand U19740 (N_19740,N_13000,N_16271);
nor U19741 (N_19741,N_13084,N_18596);
nor U19742 (N_19742,N_16050,N_16169);
nor U19743 (N_19743,N_12839,N_17993);
or U19744 (N_19744,N_13871,N_15585);
and U19745 (N_19745,N_14205,N_14694);
and U19746 (N_19746,N_14498,N_17782);
nand U19747 (N_19747,N_15038,N_12931);
and U19748 (N_19748,N_14383,N_18271);
or U19749 (N_19749,N_13201,N_16621);
nand U19750 (N_19750,N_13356,N_16023);
nor U19751 (N_19751,N_17537,N_13452);
or U19752 (N_19752,N_13975,N_18531);
or U19753 (N_19753,N_12539,N_18049);
or U19754 (N_19754,N_13883,N_13644);
nor U19755 (N_19755,N_18697,N_14360);
and U19756 (N_19756,N_17963,N_16031);
xor U19757 (N_19757,N_15853,N_13423);
nand U19758 (N_19758,N_14008,N_15172);
nand U19759 (N_19759,N_15224,N_13478);
or U19760 (N_19760,N_12983,N_12555);
nand U19761 (N_19761,N_15515,N_14940);
and U19762 (N_19762,N_13176,N_13383);
and U19763 (N_19763,N_17799,N_18242);
or U19764 (N_19764,N_17277,N_17084);
xnor U19765 (N_19765,N_15882,N_13947);
or U19766 (N_19766,N_18481,N_13911);
nor U19767 (N_19767,N_15698,N_16902);
nand U19768 (N_19768,N_18292,N_13283);
or U19769 (N_19769,N_15404,N_15214);
or U19770 (N_19770,N_15480,N_13843);
nor U19771 (N_19771,N_17849,N_15940);
nand U19772 (N_19772,N_16937,N_13278);
xnor U19773 (N_19773,N_18115,N_15118);
xnor U19774 (N_19774,N_15753,N_16302);
and U19775 (N_19775,N_16770,N_18219);
xnor U19776 (N_19776,N_16637,N_14597);
and U19777 (N_19777,N_14119,N_17677);
nor U19778 (N_19778,N_14943,N_14549);
xnor U19779 (N_19779,N_17584,N_15081);
xor U19780 (N_19780,N_14414,N_16642);
and U19781 (N_19781,N_18209,N_16303);
and U19782 (N_19782,N_18583,N_18030);
nor U19783 (N_19783,N_18498,N_18095);
xor U19784 (N_19784,N_15000,N_16636);
xor U19785 (N_19785,N_16121,N_15604);
and U19786 (N_19786,N_13537,N_13583);
nand U19787 (N_19787,N_18356,N_16265);
and U19788 (N_19788,N_18187,N_17843);
nand U19789 (N_19789,N_16042,N_12941);
or U19790 (N_19790,N_15091,N_18447);
or U19791 (N_19791,N_14483,N_16964);
nor U19792 (N_19792,N_14681,N_17909);
xor U19793 (N_19793,N_13248,N_17269);
nand U19794 (N_19794,N_12763,N_13200);
and U19795 (N_19795,N_13226,N_13509);
nor U19796 (N_19796,N_16109,N_16495);
xor U19797 (N_19797,N_17336,N_15872);
and U19798 (N_19798,N_14639,N_16474);
or U19799 (N_19799,N_18252,N_15465);
nand U19800 (N_19800,N_16778,N_18294);
xnor U19801 (N_19801,N_15956,N_16990);
nor U19802 (N_19802,N_15621,N_15490);
nand U19803 (N_19803,N_12634,N_14950);
and U19804 (N_19804,N_15360,N_17073);
nand U19805 (N_19805,N_16692,N_13962);
or U19806 (N_19806,N_18325,N_18010);
nor U19807 (N_19807,N_14137,N_15545);
and U19808 (N_19808,N_18511,N_13978);
nand U19809 (N_19809,N_13421,N_16626);
or U19810 (N_19810,N_15251,N_13144);
nor U19811 (N_19811,N_13308,N_16646);
nand U19812 (N_19812,N_16684,N_16691);
nor U19813 (N_19813,N_18499,N_15237);
nor U19814 (N_19814,N_16180,N_14659);
or U19815 (N_19815,N_17829,N_17665);
and U19816 (N_19816,N_13186,N_15750);
xnor U19817 (N_19817,N_17724,N_16628);
xnor U19818 (N_19818,N_12584,N_15624);
and U19819 (N_19819,N_17761,N_18508);
nor U19820 (N_19820,N_15995,N_13694);
or U19821 (N_19821,N_12720,N_12605);
nor U19822 (N_19822,N_14697,N_15265);
and U19823 (N_19823,N_16012,N_14045);
or U19824 (N_19824,N_18316,N_18056);
nand U19825 (N_19825,N_13482,N_16629);
nand U19826 (N_19826,N_12887,N_17234);
or U19827 (N_19827,N_14293,N_18331);
nand U19828 (N_19828,N_14939,N_15774);
or U19829 (N_19829,N_13543,N_12871);
xor U19830 (N_19830,N_18459,N_16269);
and U19831 (N_19831,N_17554,N_13256);
or U19832 (N_19832,N_13797,N_16021);
and U19833 (N_19833,N_15342,N_15710);
nor U19834 (N_19834,N_14546,N_12674);
nor U19835 (N_19835,N_16310,N_14671);
xor U19836 (N_19836,N_15805,N_12578);
nand U19837 (N_19837,N_14405,N_17460);
and U19838 (N_19838,N_13498,N_16321);
or U19839 (N_19839,N_13967,N_12942);
xor U19840 (N_19840,N_13299,N_14169);
xor U19841 (N_19841,N_18199,N_16402);
or U19842 (N_19842,N_18743,N_16820);
and U19843 (N_19843,N_16607,N_12934);
nand U19844 (N_19844,N_12732,N_13375);
nor U19845 (N_19845,N_18725,N_17422);
xnor U19846 (N_19846,N_16341,N_12646);
xnor U19847 (N_19847,N_16543,N_17732);
nand U19848 (N_19848,N_12658,N_16959);
xnor U19849 (N_19849,N_17651,N_17166);
xnor U19850 (N_19850,N_17738,N_14193);
or U19851 (N_19851,N_14313,N_17216);
xnor U19852 (N_19852,N_18268,N_13590);
or U19853 (N_19853,N_17937,N_16372);
nand U19854 (N_19854,N_17652,N_17888);
nor U19855 (N_19855,N_15565,N_16516);
xnor U19856 (N_19856,N_18601,N_17414);
xnor U19857 (N_19857,N_16708,N_16062);
and U19858 (N_19858,N_15798,N_17752);
nand U19859 (N_19859,N_17276,N_18602);
nor U19860 (N_19860,N_16529,N_17974);
nor U19861 (N_19861,N_15641,N_14026);
nand U19862 (N_19862,N_15183,N_17551);
nand U19863 (N_19863,N_14075,N_16110);
xnor U19864 (N_19864,N_13237,N_16743);
nor U19865 (N_19865,N_14234,N_17467);
and U19866 (N_19866,N_12980,N_16066);
xnor U19867 (N_19867,N_18422,N_16074);
nand U19868 (N_19868,N_13747,N_16705);
or U19869 (N_19869,N_15127,N_16872);
or U19870 (N_19870,N_18015,N_15258);
nand U19871 (N_19871,N_16077,N_17934);
xnor U19872 (N_19872,N_14756,N_17156);
nor U19873 (N_19873,N_12719,N_17119);
or U19874 (N_19874,N_14562,N_13566);
or U19875 (N_19875,N_18642,N_15132);
xnor U19876 (N_19876,N_16319,N_18592);
xnor U19877 (N_19877,N_18733,N_15094);
or U19878 (N_19878,N_15070,N_12639);
and U19879 (N_19879,N_14328,N_12530);
xnor U19880 (N_19880,N_14571,N_13236);
or U19881 (N_19881,N_14708,N_14447);
nand U19882 (N_19882,N_16817,N_14613);
and U19883 (N_19883,N_16856,N_16950);
nor U19884 (N_19884,N_14064,N_13621);
or U19885 (N_19885,N_15771,N_13565);
and U19886 (N_19886,N_15004,N_16729);
or U19887 (N_19887,N_15770,N_13035);
nor U19888 (N_19888,N_14223,N_12576);
nor U19889 (N_19889,N_12592,N_13701);
nor U19890 (N_19890,N_18712,N_12640);
nor U19891 (N_19891,N_13499,N_17272);
nor U19892 (N_19892,N_13649,N_13184);
xor U19893 (N_19893,N_17394,N_12894);
nand U19894 (N_19894,N_15826,N_14786);
or U19895 (N_19895,N_12924,N_13466);
or U19896 (N_19896,N_16329,N_13322);
or U19897 (N_19897,N_12769,N_12697);
or U19898 (N_19898,N_13551,N_16029);
nor U19899 (N_19899,N_13483,N_16106);
nand U19900 (N_19900,N_14874,N_18713);
nor U19901 (N_19901,N_13998,N_15675);
nor U19902 (N_19902,N_15463,N_13958);
nor U19903 (N_19903,N_16680,N_16830);
or U19904 (N_19904,N_18390,N_16218);
nor U19905 (N_19905,N_16315,N_14870);
nand U19906 (N_19906,N_17773,N_15059);
nor U19907 (N_19907,N_17352,N_13005);
nand U19908 (N_19908,N_16173,N_17024);
nor U19909 (N_19909,N_15806,N_16475);
nand U19910 (N_19910,N_16095,N_17174);
or U19911 (N_19911,N_15531,N_13205);
xor U19912 (N_19912,N_13633,N_13792);
xnor U19913 (N_19913,N_13300,N_17542);
nor U19914 (N_19914,N_13742,N_15884);
and U19915 (N_19915,N_14722,N_17790);
nand U19916 (N_19916,N_15161,N_15201);
or U19917 (N_19917,N_15576,N_14714);
and U19918 (N_19918,N_13134,N_15866);
nand U19919 (N_19919,N_13413,N_14788);
nand U19920 (N_19920,N_18094,N_12527);
or U19921 (N_19921,N_15507,N_17134);
nand U19922 (N_19922,N_13899,N_17449);
and U19923 (N_19923,N_15134,N_16792);
nand U19924 (N_19924,N_14873,N_15006);
nor U19925 (N_19925,N_17639,N_17973);
or U19926 (N_19926,N_14259,N_14032);
and U19927 (N_19927,N_14951,N_13969);
or U19928 (N_19928,N_17893,N_16335);
or U19929 (N_19929,N_18490,N_14566);
or U19930 (N_19930,N_17812,N_18066);
or U19931 (N_19931,N_13179,N_14773);
xor U19932 (N_19932,N_17524,N_17334);
nor U19933 (N_19933,N_17774,N_12928);
and U19934 (N_19934,N_14695,N_15196);
xnor U19935 (N_19935,N_17475,N_18272);
or U19936 (N_19936,N_13511,N_14105);
xor U19937 (N_19937,N_13624,N_15591);
nand U19938 (N_19938,N_18665,N_14212);
nand U19939 (N_19939,N_14929,N_14138);
xnor U19940 (N_19940,N_14511,N_18189);
xnor U19941 (N_19941,N_18589,N_17398);
nand U19942 (N_19942,N_16481,N_17796);
nand U19943 (N_19943,N_18054,N_13926);
xor U19944 (N_19944,N_14994,N_12816);
and U19945 (N_19945,N_18149,N_13850);
nor U19946 (N_19946,N_16541,N_16501);
or U19947 (N_19947,N_18055,N_16378);
or U19948 (N_19948,N_13801,N_18235);
nand U19949 (N_19949,N_12822,N_14442);
nand U19950 (N_19950,N_15371,N_13870);
or U19951 (N_19951,N_14844,N_15997);
and U19952 (N_19952,N_15540,N_15699);
or U19953 (N_19953,N_17939,N_13762);
nand U19954 (N_19954,N_16139,N_18570);
and U19955 (N_19955,N_15773,N_17933);
or U19956 (N_19956,N_16426,N_13872);
nand U19957 (N_19957,N_14340,N_12938);
and U19958 (N_19958,N_18440,N_17429);
nand U19959 (N_19959,N_13859,N_12657);
and U19960 (N_19960,N_18414,N_18132);
nor U19961 (N_19961,N_16723,N_13514);
xnor U19962 (N_19962,N_13919,N_12772);
xnor U19963 (N_19963,N_13868,N_18486);
xor U19964 (N_19964,N_12752,N_13063);
nor U19965 (N_19965,N_17824,N_17387);
xor U19966 (N_19966,N_13502,N_17658);
nor U19967 (N_19967,N_16202,N_18424);
and U19968 (N_19968,N_12962,N_12848);
xor U19969 (N_19969,N_14235,N_15307);
and U19970 (N_19970,N_17765,N_17199);
xor U19971 (N_19971,N_15219,N_18134);
nor U19972 (N_19972,N_13695,N_16371);
and U19973 (N_19973,N_13616,N_14758);
nand U19974 (N_19974,N_17463,N_14976);
xnor U19975 (N_19975,N_14723,N_15204);
or U19976 (N_19976,N_12616,N_15833);
and U19977 (N_19977,N_12562,N_16491);
and U19978 (N_19978,N_15758,N_16296);
and U19979 (N_19979,N_14164,N_14038);
xnor U19980 (N_19980,N_15349,N_15300);
nand U19981 (N_19981,N_17586,N_12541);
xnor U19982 (N_19982,N_15603,N_18263);
or U19983 (N_19983,N_17688,N_16071);
and U19984 (N_19984,N_14110,N_14698);
nand U19985 (N_19985,N_16450,N_16662);
nor U19986 (N_19986,N_13170,N_16144);
or U19987 (N_19987,N_13522,N_17625);
nor U19988 (N_19988,N_15415,N_14789);
or U19989 (N_19989,N_15226,N_13976);
nand U19990 (N_19990,N_18279,N_16119);
nor U19991 (N_19991,N_15823,N_15071);
nor U19992 (N_19992,N_16916,N_13878);
nor U19993 (N_19993,N_13339,N_18372);
xnor U19994 (N_19994,N_13385,N_18223);
xnor U19995 (N_19995,N_13487,N_17454);
nor U19996 (N_19996,N_17705,N_14101);
xor U19997 (N_19997,N_13703,N_14993);
nand U19998 (N_19998,N_17254,N_12766);
xnor U19999 (N_19999,N_14742,N_12601);
or U20000 (N_20000,N_17612,N_14634);
xor U20001 (N_20001,N_15740,N_17355);
or U20002 (N_20002,N_15613,N_15497);
nor U20003 (N_20003,N_15352,N_16889);
and U20004 (N_20004,N_15403,N_15611);
xnor U20005 (N_20005,N_14353,N_18509);
xor U20006 (N_20006,N_16272,N_13771);
or U20007 (N_20007,N_14871,N_14514);
xor U20008 (N_20008,N_17529,N_15664);
nand U20009 (N_20009,N_12919,N_14565);
and U20010 (N_20010,N_16460,N_15672);
xor U20011 (N_20011,N_16289,N_18014);
and U20012 (N_20012,N_15399,N_12847);
or U20013 (N_20013,N_16195,N_16255);
nand U20014 (N_20014,N_13479,N_12993);
xor U20015 (N_20015,N_17265,N_16867);
xnor U20016 (N_20016,N_16799,N_18264);
xor U20017 (N_20017,N_18108,N_17397);
nand U20018 (N_20018,N_18748,N_18613);
and U20019 (N_20019,N_18505,N_17624);
nand U20020 (N_20020,N_15801,N_13849);
xnor U20021 (N_20021,N_12959,N_16540);
nand U20022 (N_20022,N_14126,N_17450);
xor U20023 (N_20023,N_14191,N_13954);
and U20024 (N_20024,N_15937,N_15983);
or U20025 (N_20025,N_16613,N_17168);
nand U20026 (N_20026,N_15442,N_17700);
xor U20027 (N_20027,N_17285,N_16663);
or U20028 (N_20028,N_13086,N_18180);
or U20029 (N_20029,N_18561,N_15355);
and U20030 (N_20030,N_13163,N_12817);
nor U20031 (N_20031,N_14132,N_16900);
nor U20032 (N_20032,N_14772,N_13905);
or U20033 (N_20033,N_17815,N_17194);
nand U20034 (N_20034,N_16359,N_15273);
nor U20035 (N_20035,N_17210,N_13966);
or U20036 (N_20036,N_16231,N_18477);
xnor U20037 (N_20037,N_15582,N_13146);
and U20038 (N_20038,N_16225,N_16128);
nand U20039 (N_20039,N_14381,N_13431);
and U20040 (N_20040,N_18218,N_14709);
nor U20041 (N_20041,N_16667,N_16016);
xor U20042 (N_20042,N_15669,N_16715);
nor U20043 (N_20043,N_14598,N_14378);
and U20044 (N_20044,N_12787,N_12911);
nor U20045 (N_20045,N_17848,N_16831);
nand U20046 (N_20046,N_14808,N_13174);
nand U20047 (N_20047,N_17386,N_17196);
nand U20048 (N_20048,N_12622,N_16844);
nand U20049 (N_20049,N_17478,N_14945);
and U20050 (N_20050,N_12597,N_14415);
nand U20051 (N_20051,N_13109,N_13866);
and U20052 (N_20052,N_14975,N_13646);
or U20053 (N_20053,N_14640,N_16893);
and U20054 (N_20054,N_15789,N_16404);
or U20055 (N_20055,N_18069,N_17339);
and U20056 (N_20056,N_12838,N_13288);
nand U20057 (N_20057,N_15828,N_18525);
or U20058 (N_20058,N_18172,N_13107);
xor U20059 (N_20059,N_15104,N_13331);
or U20060 (N_20060,N_13284,N_18736);
nor U20061 (N_20061,N_13422,N_15023);
nand U20062 (N_20062,N_16949,N_15963);
xor U20063 (N_20063,N_16170,N_14524);
nor U20064 (N_20064,N_18104,N_18336);
nand U20065 (N_20065,N_16734,N_18101);
nand U20066 (N_20066,N_18457,N_18615);
and U20067 (N_20067,N_17745,N_15175);
xor U20068 (N_20068,N_15347,N_13384);
or U20069 (N_20069,N_15260,N_13692);
nor U20070 (N_20070,N_17785,N_14260);
nor U20071 (N_20071,N_17695,N_15467);
xnor U20072 (N_20072,N_17220,N_14211);
or U20073 (N_20073,N_14000,N_15220);
nor U20074 (N_20074,N_15049,N_16212);
or U20075 (N_20075,N_15534,N_17523);
nand U20076 (N_20076,N_14679,N_16764);
nand U20077 (N_20077,N_15012,N_18026);
nor U20078 (N_20078,N_17173,N_13294);
nand U20079 (N_20079,N_12702,N_15532);
nor U20080 (N_20080,N_17444,N_16611);
or U20081 (N_20081,N_14446,N_18493);
xor U20082 (N_20082,N_16732,N_15274);
nor U20083 (N_20083,N_17373,N_18314);
and U20084 (N_20084,N_13314,N_13269);
or U20085 (N_20085,N_14617,N_15843);
nor U20086 (N_20086,N_12585,N_17944);
xor U20087 (N_20087,N_17410,N_12912);
xnor U20088 (N_20088,N_15133,N_15107);
nor U20089 (N_20089,N_16772,N_16757);
nor U20090 (N_20090,N_18274,N_14275);
or U20091 (N_20091,N_15414,N_14997);
or U20092 (N_20092,N_15925,N_17244);
and U20093 (N_20093,N_16930,N_17327);
nor U20094 (N_20094,N_18074,N_17538);
nand U20095 (N_20095,N_17721,N_13255);
nand U20096 (N_20096,N_17712,N_17807);
nand U20097 (N_20097,N_13317,N_14304);
nand U20098 (N_20098,N_14278,N_13253);
nor U20099 (N_20099,N_15009,N_14944);
xor U20100 (N_20100,N_12545,N_13223);
or U20101 (N_20101,N_18575,N_12522);
xor U20102 (N_20102,N_16181,N_13293);
or U20103 (N_20103,N_14762,N_15242);
nand U20104 (N_20104,N_17525,N_18518);
nor U20105 (N_20105,N_18420,N_14157);
or U20106 (N_20106,N_16822,N_14396);
nand U20107 (N_20107,N_15597,N_15296);
nand U20108 (N_20108,N_16229,N_16601);
nor U20109 (N_20109,N_15377,N_18657);
nor U20110 (N_20110,N_13175,N_12636);
nor U20111 (N_20111,N_17412,N_14346);
nor U20112 (N_20112,N_15952,N_16472);
and U20113 (N_20113,N_18667,N_16525);
nor U20114 (N_20114,N_13062,N_12780);
nand U20115 (N_20115,N_16198,N_18453);
xnor U20116 (N_20116,N_16049,N_15845);
nor U20117 (N_20117,N_18173,N_18401);
nand U20118 (N_20118,N_15160,N_15020);
nand U20119 (N_20119,N_17008,N_15908);
or U20120 (N_20120,N_12902,N_18086);
or U20121 (N_20121,N_12745,N_12827);
nor U20122 (N_20122,N_13542,N_15896);
or U20123 (N_20123,N_13764,N_17004);
nor U20124 (N_20124,N_16159,N_13009);
and U20125 (N_20125,N_12520,N_13489);
or U20126 (N_20126,N_17287,N_17052);
and U20127 (N_20127,N_13855,N_12799);
nor U20128 (N_20128,N_17432,N_18288);
nor U20129 (N_20129,N_17819,N_16549);
nor U20130 (N_20130,N_16320,N_14017);
or U20131 (N_20131,N_15659,N_18045);
nand U20132 (N_20132,N_13484,N_17407);
nor U20133 (N_20133,N_16358,N_18221);
or U20134 (N_20134,N_16111,N_18738);
xor U20135 (N_20135,N_15241,N_13861);
and U20136 (N_20136,N_16248,N_17392);
and U20137 (N_20137,N_15376,N_13117);
nor U20138 (N_20138,N_14812,N_15339);
nor U20139 (N_20139,N_18299,N_14322);
xor U20140 (N_20140,N_13392,N_17716);
and U20141 (N_20141,N_14991,N_17820);
xor U20142 (N_20142,N_15202,N_15584);
and U20143 (N_20143,N_18398,N_15476);
or U20144 (N_20144,N_13252,N_14682);
xnor U20145 (N_20145,N_18749,N_17261);
nand U20146 (N_20146,N_15210,N_14648);
and U20147 (N_20147,N_15707,N_13931);
or U20148 (N_20148,N_13650,N_16297);
and U20149 (N_20149,N_18487,N_17110);
nand U20150 (N_20150,N_18470,N_16992);
or U20151 (N_20151,N_14033,N_14436);
nand U20152 (N_20152,N_16630,N_17867);
or U20153 (N_20153,N_15760,N_14444);
xor U20154 (N_20154,N_13094,N_13974);
and U20155 (N_20155,N_16236,N_14687);
or U20156 (N_20156,N_12625,N_17251);
and U20157 (N_20157,N_17253,N_15130);
and U20158 (N_20158,N_16700,N_17544);
nor U20159 (N_20159,N_15596,N_16941);
and U20160 (N_20160,N_13480,N_15413);
xnor U20161 (N_20161,N_18502,N_17719);
nand U20162 (N_20162,N_16652,N_13120);
or U20163 (N_20163,N_15456,N_17946);
or U20164 (N_20164,N_12725,N_12535);
nor U20165 (N_20165,N_18186,N_15272);
xor U20166 (N_20166,N_13406,N_17440);
nor U20167 (N_20167,N_13013,N_13245);
or U20168 (N_20168,N_13360,N_17683);
or U20169 (N_20169,N_13665,N_17922);
and U20170 (N_20170,N_14854,N_15589);
xnor U20171 (N_20171,N_16443,N_14124);
nand U20172 (N_20172,N_12989,N_14049);
or U20173 (N_20173,N_17292,N_13191);
or U20174 (N_20174,N_16151,N_14076);
or U20175 (N_20175,N_17019,N_16135);
or U20176 (N_20176,N_13229,N_17338);
or U20177 (N_20177,N_17230,N_14843);
nor U20178 (N_20178,N_18118,N_14465);
and U20179 (N_20179,N_14672,N_18004);
nand U20180 (N_20180,N_15216,N_16389);
xor U20181 (N_20181,N_14580,N_18362);
or U20182 (N_20182,N_15646,N_15581);
or U20183 (N_20183,N_15825,N_12696);
nor U20184 (N_20184,N_14632,N_16603);
xor U20185 (N_20185,N_15187,N_16207);
and U20186 (N_20186,N_17263,N_13412);
and U20187 (N_20187,N_17201,N_17615);
nor U20188 (N_20188,N_15615,N_18418);
nand U20189 (N_20189,N_18072,N_13845);
xnor U20190 (N_20190,N_18048,N_13281);
nand U20191 (N_20191,N_13188,N_15875);
xnor U20192 (N_20192,N_15498,N_14710);
nand U20193 (N_20193,N_16920,N_18019);
or U20194 (N_20194,N_17419,N_14816);
and U20195 (N_20195,N_15407,N_12842);
nand U20196 (N_20196,N_12502,N_18718);
and U20197 (N_20197,N_18648,N_14631);
or U20198 (N_20198,N_17912,N_14010);
and U20199 (N_20199,N_14832,N_13442);
and U20200 (N_20200,N_14448,N_13453);
nor U20201 (N_20201,N_16459,N_15682);
xor U20202 (N_20202,N_14609,N_17957);
or U20203 (N_20203,N_18684,N_16978);
nor U20204 (N_20204,N_13266,N_17310);
and U20205 (N_20205,N_18140,N_14084);
nand U20206 (N_20206,N_18706,N_16162);
nor U20207 (N_20207,N_15369,N_17378);
nand U20208 (N_20208,N_13342,N_14935);
and U20209 (N_20209,N_14218,N_17112);
nor U20210 (N_20210,N_13832,N_16527);
or U20211 (N_20211,N_13655,N_15110);
or U20212 (N_20212,N_16713,N_18631);
xnor U20213 (N_20213,N_17436,N_14517);
nor U20214 (N_20214,N_14154,N_13335);
or U20215 (N_20215,N_15390,N_17956);
nand U20216 (N_20216,N_17459,N_17951);
xor U20217 (N_20217,N_16986,N_15759);
nor U20218 (N_20218,N_14777,N_14783);
and U20219 (N_20219,N_12939,N_12507);
and U20220 (N_20220,N_13419,N_16768);
and U20221 (N_20221,N_13346,N_18234);
nor U20222 (N_20222,N_13856,N_14011);
nand U20223 (N_20223,N_13089,N_17687);
or U20224 (N_20224,N_18722,N_14367);
and U20225 (N_20225,N_17772,N_18645);
or U20226 (N_20226,N_17433,N_18519);
or U20227 (N_20227,N_15264,N_14956);
nand U20228 (N_20228,N_15556,N_14925);
nand U20229 (N_20229,N_12713,N_13445);
nand U20230 (N_20230,N_15880,N_14172);
or U20231 (N_20231,N_14889,N_18124);
xor U20232 (N_20232,N_16370,N_15988);
and U20233 (N_20233,N_15520,N_15139);
and U20234 (N_20234,N_18225,N_13165);
or U20235 (N_20235,N_13439,N_17873);
nand U20236 (N_20236,N_16803,N_13585);
or U20237 (N_20237,N_14683,N_13275);
nor U20238 (N_20238,N_15190,N_14790);
nor U20239 (N_20239,N_14041,N_17997);
xnor U20240 (N_20240,N_13841,N_13860);
xor U20241 (N_20241,N_16158,N_12610);
and U20242 (N_20242,N_17797,N_15657);
nor U20243 (N_20243,N_16206,N_17751);
nand U20244 (N_20244,N_15207,N_18562);
xor U20245 (N_20245,N_13267,N_13885);
nor U20246 (N_20246,N_18192,N_18246);
nand U20247 (N_20247,N_16356,N_15112);
nand U20248 (N_20248,N_16631,N_13927);
xnor U20249 (N_20249,N_14397,N_14220);
nor U20250 (N_20250,N_14181,N_15318);
xnor U20251 (N_20251,N_15055,N_17520);
nand U20252 (N_20252,N_15942,N_16786);
nor U20253 (N_20253,N_16041,N_16113);
and U20254 (N_20254,N_15211,N_18627);
xnor U20255 (N_20255,N_13238,N_14180);
and U20256 (N_20256,N_12537,N_18000);
nor U20257 (N_20257,N_13833,N_15341);
xnor U20258 (N_20258,N_17304,N_17764);
nand U20259 (N_20259,N_16526,N_14027);
nand U20260 (N_20260,N_13074,N_14337);
xor U20261 (N_20261,N_18366,N_17167);
nor U20262 (N_20262,N_18595,N_14379);
xnor U20263 (N_20263,N_17144,N_15919);
nor U20264 (N_20264,N_16373,N_14197);
or U20265 (N_20265,N_13048,N_14484);
xor U20266 (N_20266,N_16290,N_18156);
or U20267 (N_20267,N_18421,N_12548);
nor U20268 (N_20268,N_14196,N_17857);
xnor U20269 (N_20269,N_13496,N_15011);
and U20270 (N_20270,N_18746,N_14081);
or U20271 (N_20271,N_18135,N_13744);
nand U20272 (N_20272,N_18579,N_18637);
nor U20273 (N_20273,N_14567,N_15487);
or U20274 (N_20274,N_17727,N_17041);
or U20275 (N_20275,N_16687,N_14085);
xnor U20276 (N_20276,N_13066,N_16780);
nor U20277 (N_20277,N_13078,N_13715);
xor U20278 (N_20278,N_17638,N_16328);
and U20279 (N_20279,N_15449,N_17317);
xnor U20280 (N_20280,N_13824,N_17312);
and U20281 (N_20281,N_13209,N_16609);
and U20282 (N_20282,N_16393,N_18696);
nor U20283 (N_20283,N_18680,N_16288);
nor U20284 (N_20284,N_18563,N_13706);
nand U20285 (N_20285,N_18660,N_13235);
nand U20286 (N_20286,N_17258,N_12510);
xor U20287 (N_20287,N_15878,N_14474);
nand U20288 (N_20288,N_16076,N_12784);
nand U20289 (N_20289,N_13068,N_15901);
and U20290 (N_20290,N_14273,N_13517);
or U20291 (N_20291,N_17341,N_16204);
nand U20292 (N_20292,N_14607,N_15892);
nor U20293 (N_20293,N_14733,N_15852);
nand U20294 (N_20294,N_16619,N_17290);
or U20295 (N_20295,N_18131,N_17375);
xnor U20296 (N_20296,N_12619,N_17055);
or U20297 (N_20297,N_16256,N_17161);
xnor U20298 (N_20298,N_12566,N_12861);
xor U20299 (N_20299,N_13758,N_14274);
nand U20300 (N_20300,N_17030,N_14286);
or U20301 (N_20301,N_16848,N_13307);
nand U20302 (N_20302,N_15660,N_17259);
nand U20303 (N_20303,N_16138,N_16919);
and U20304 (N_20304,N_18444,N_15199);
xnor U20305 (N_20305,N_17604,N_14036);
nor U20306 (N_20306,N_18122,N_15918);
nand U20307 (N_20307,N_15136,N_18158);
xnor U20308 (N_20308,N_18567,N_17605);
or U20309 (N_20309,N_14489,N_16194);
nand U20310 (N_20310,N_16539,N_17540);
or U20311 (N_20311,N_16939,N_15676);
nor U20312 (N_20312,N_15502,N_15281);
xnor U20313 (N_20313,N_17160,N_15528);
nor U20314 (N_20314,N_13823,N_14897);
or U20315 (N_20315,N_14651,N_16769);
and U20316 (N_20316,N_14916,N_14990);
nor U20317 (N_20317,N_13247,N_16824);
nor U20318 (N_20318,N_15612,N_13753);
and U20319 (N_20319,N_14242,N_12882);
nand U20320 (N_20320,N_14981,N_17275);
nor U20321 (N_20321,N_13987,N_14393);
nand U20322 (N_20322,N_12782,N_14801);
nor U20323 (N_20323,N_18415,N_15860);
nand U20324 (N_20324,N_15856,N_16322);
or U20325 (N_20325,N_12515,N_17767);
xor U20326 (N_20326,N_18692,N_18371);
nand U20327 (N_20327,N_13599,N_14933);
or U20328 (N_20328,N_12519,N_17138);
nand U20329 (N_20329,N_13795,N_15088);
and U20330 (N_20330,N_17231,N_13059);
and U20331 (N_20331,N_15717,N_15477);
or U20332 (N_20332,N_13982,N_15069);
or U20333 (N_20333,N_17522,N_17182);
or U20334 (N_20334,N_18239,N_12802);
and U20335 (N_20335,N_16361,N_13132);
nor U20336 (N_20336,N_14411,N_18668);
nand U20337 (N_20337,N_14973,N_12965);
nor U20338 (N_20338,N_17293,N_14179);
xor U20339 (N_20339,N_12828,N_15140);
nand U20340 (N_20340,N_15324,N_18515);
or U20341 (N_20341,N_15165,N_16283);
nor U20342 (N_20342,N_18666,N_16241);
and U20343 (N_20343,N_13981,N_16678);
and U20344 (N_20344,N_17846,N_14385);
nand U20345 (N_20345,N_14394,N_14065);
and U20346 (N_20346,N_13904,N_14373);
or U20347 (N_20347,N_17647,N_15311);
and U20348 (N_20348,N_12978,N_13805);
nand U20349 (N_20349,N_13541,N_18537);
nand U20350 (N_20350,N_17757,N_15067);
nor U20351 (N_20351,N_14615,N_18584);
nor U20352 (N_20352,N_15550,N_12900);
or U20353 (N_20353,N_17155,N_16018);
and U20354 (N_20354,N_16161,N_17010);
xnor U20355 (N_20355,N_18625,N_12937);
nand U20356 (N_20356,N_14206,N_16434);
and U20357 (N_20357,N_16383,N_17545);
nor U20358 (N_20358,N_15182,N_18409);
xnor U20359 (N_20359,N_15245,N_18365);
nand U20360 (N_20360,N_17579,N_16783);
nor U20361 (N_20361,N_14413,N_15712);
nand U20362 (N_20362,N_14526,N_13777);
xnor U20363 (N_20363,N_18142,N_16711);
xor U20364 (N_20364,N_16987,N_14965);
nand U20365 (N_20365,N_17061,N_13582);
nand U20366 (N_20366,N_14850,N_18672);
nor U20367 (N_20367,N_18541,N_12809);
nand U20368 (N_20368,N_13318,N_13943);
nor U20369 (N_20369,N_13195,N_18052);
xor U20370 (N_20370,N_14545,N_14884);
xor U20371 (N_20371,N_16800,N_18116);
xor U20372 (N_20372,N_18640,N_15388);
and U20373 (N_20373,N_16551,N_17468);
nand U20374 (N_20374,N_16869,N_13258);
nor U20375 (N_20375,N_17979,N_15179);
xor U20376 (N_20376,N_15775,N_13660);
xnor U20377 (N_20377,N_12757,N_18161);
nand U20378 (N_20378,N_14182,N_15075);
xnor U20379 (N_20379,N_14106,N_16164);
nor U20380 (N_20380,N_14938,N_12571);
or U20381 (N_20381,N_15982,N_18171);
nor U20382 (N_20382,N_18405,N_17243);
and U20383 (N_20383,N_12863,N_15650);
nor U20384 (N_20384,N_16673,N_18553);
nand U20385 (N_20385,N_13077,N_14650);
nand U20386 (N_20386,N_14868,N_14091);
xor U20387 (N_20387,N_14794,N_17437);
nor U20388 (N_20388,N_16943,N_14320);
or U20389 (N_20389,N_15084,N_18328);
and U20390 (N_20390,N_12881,N_13135);
xnor U20391 (N_20391,N_16910,N_12538);
or U20392 (N_20392,N_18494,N_16494);
xor U20393 (N_20393,N_14657,N_14122);
nand U20394 (N_20394,N_18177,N_14371);
or U20395 (N_20395,N_16052,N_12872);
nor U20396 (N_20396,N_18253,N_16521);
nand U20397 (N_20397,N_16657,N_13321);
nor U20398 (N_20398,N_13507,N_14628);
nor U20399 (N_20399,N_18193,N_14963);
nor U20400 (N_20400,N_18112,N_16477);
and U20401 (N_20401,N_16337,N_16796);
nor U20402 (N_20402,N_12996,N_13398);
and U20403 (N_20403,N_15525,N_15381);
or U20404 (N_20404,N_17068,N_15197);
and U20405 (N_20405,N_14803,N_16773);
xor U20406 (N_20406,N_14901,N_15903);
xor U20407 (N_20407,N_13736,N_13058);
or U20408 (N_20408,N_14600,N_13915);
or U20409 (N_20409,N_15783,N_18100);
nor U20410 (N_20410,N_14283,N_13923);
and U20411 (N_20411,N_15469,N_17116);
nand U20412 (N_20412,N_17988,N_17121);
nor U20413 (N_20413,N_13669,N_15485);
or U20414 (N_20414,N_17060,N_16829);
xor U20415 (N_20415,N_16738,N_14018);
nor U20416 (N_20416,N_18507,N_13405);
nor U20417 (N_20417,N_12767,N_14445);
and U20418 (N_20418,N_13337,N_14021);
and U20419 (N_20419,N_13472,N_12865);
and U20420 (N_20420,N_15721,N_15579);
nand U20421 (N_20421,N_15987,N_15854);
xor U20422 (N_20422,N_15633,N_18464);
and U20423 (N_20423,N_14563,N_13040);
or U20424 (N_20424,N_14088,N_15954);
nand U20425 (N_20425,N_16313,N_17403);
xnor U20426 (N_20426,N_13846,N_12764);
and U20427 (N_20427,N_14507,N_16676);
and U20428 (N_20428,N_14797,N_18126);
nand U20429 (N_20429,N_15213,N_17681);
nand U20430 (N_20430,N_16230,N_18353);
xor U20431 (N_20431,N_17744,N_15523);
or U20432 (N_20432,N_16376,N_14155);
nand U20433 (N_20433,N_16227,N_18210);
or U20434 (N_20434,N_17053,N_16166);
or U20435 (N_20435,N_16624,N_14280);
and U20436 (N_20436,N_15886,N_15765);
nor U20437 (N_20437,N_15889,N_15704);
and U20438 (N_20438,N_14057,N_17445);
and U20439 (N_20439,N_17095,N_18370);
or U20440 (N_20440,N_13382,N_15764);
nand U20441 (N_20441,N_13743,N_17892);
nand U20442 (N_20442,N_12945,N_17531);
or U20443 (N_20443,N_12818,N_15253);
or U20444 (N_20444,N_16350,N_17616);
or U20445 (N_20445,N_14653,N_18606);
nor U20446 (N_20446,N_18730,N_15062);
xnor U20447 (N_20447,N_16948,N_17078);
nand U20448 (N_20448,N_12759,N_17143);
nand U20449 (N_20449,N_14556,N_13814);
and U20450 (N_20450,N_15329,N_17162);
or U20451 (N_20451,N_15976,N_17570);
or U20452 (N_20452,N_14591,N_15392);
nor U20453 (N_20453,N_14190,N_16440);
nor U20454 (N_20454,N_13601,N_18699);
nand U20455 (N_20455,N_15677,N_18658);
nand U20456 (N_20456,N_17515,N_16223);
or U20457 (N_20457,N_13984,N_14469);
nor U20458 (N_20458,N_15106,N_15746);
xor U20459 (N_20459,N_13426,N_13822);
and U20460 (N_20460,N_15642,N_14482);
xnor U20461 (N_20461,N_15317,N_18377);
and U20462 (N_20462,N_14186,N_16094);
or U20463 (N_20463,N_16090,N_17527);
xor U20464 (N_20464,N_12753,N_13368);
and U20465 (N_20465,N_16991,N_18097);
nand U20466 (N_20466,N_16781,N_16722);
and U20467 (N_20467,N_18001,N_16010);
xor U20468 (N_20468,N_13613,N_14416);
nor U20469 (N_20469,N_15639,N_15951);
nand U20470 (N_20470,N_18284,N_16887);
or U20471 (N_20471,N_18050,N_16945);
xnor U20472 (N_20472,N_13900,N_17868);
and U20473 (N_20473,N_14116,N_13587);
nor U20474 (N_20474,N_15212,N_13407);
or U20475 (N_20475,N_12781,N_18089);
and U20476 (N_20476,N_16926,N_12504);
xnor U20477 (N_20477,N_12649,N_17447);
xor U20478 (N_20478,N_12834,N_14388);
or U20479 (N_20479,N_17620,N_18355);
nand U20480 (N_20480,N_16721,N_14717);
and U20481 (N_20481,N_12905,N_18040);
or U20482 (N_20482,N_17297,N_13722);
xnor U20483 (N_20483,N_13217,N_12899);
nand U20484 (N_20484,N_12665,N_13023);
nand U20485 (N_20485,N_17575,N_18510);
xnor U20486 (N_20486,N_16392,N_16672);
nor U20487 (N_20487,N_15382,N_12792);
nor U20488 (N_20488,N_12984,N_13438);
or U20489 (N_20489,N_14673,N_16362);
or U20490 (N_20490,N_16989,N_18410);
and U20491 (N_20491,N_14799,N_14917);
or U20492 (N_20492,N_16903,N_14070);
nand U20493 (N_20493,N_16659,N_13305);
and U20494 (N_20494,N_17662,N_17998);
and U20495 (N_20495,N_15813,N_14547);
and U20496 (N_20496,N_16934,N_15640);
and U20497 (N_20497,N_12921,N_17324);
nand U20498 (N_20498,N_18727,N_17330);
nor U20499 (N_20499,N_17067,N_13121);
nor U20500 (N_20500,N_16410,N_14837);
xor U20501 (N_20501,N_15724,N_16441);
nand U20502 (N_20502,N_16511,N_15302);
and U20503 (N_20503,N_16129,N_18516);
nor U20504 (N_20504,N_14417,N_17536);
xor U20505 (N_20505,N_14421,N_14074);
and U20506 (N_20506,N_14380,N_16038);
or U20507 (N_20507,N_17889,N_12990);
xnor U20508 (N_20508,N_17827,N_15551);
and U20509 (N_20509,N_15436,N_17854);
nor U20510 (N_20510,N_15761,N_15609);
or U20511 (N_20511,N_15966,N_12917);
nor U20512 (N_20512,N_16323,N_18168);
and U20513 (N_20513,N_18369,N_15044);
or U20514 (N_20514,N_17811,N_16544);
xnor U20515 (N_20515,N_17950,N_16653);
or U20516 (N_20516,N_13244,N_14712);
nand U20517 (N_20517,N_12875,N_14485);
nand U20518 (N_20518,N_16699,N_18621);
nand U20519 (N_20519,N_16774,N_14354);
nor U20520 (N_20520,N_17185,N_17674);
and U20521 (N_20521,N_15816,N_17048);
or U20522 (N_20522,N_18148,N_17965);
and U20523 (N_20523,N_14114,N_12735);
xnor U20524 (N_20524,N_17600,N_15432);
nor U20525 (N_20525,N_16122,N_13724);
xnor U20526 (N_20526,N_15064,N_18389);
and U20527 (N_20527,N_13547,N_15719);
nand U20528 (N_20528,N_12641,N_14702);
xor U20529 (N_20529,N_16993,N_15066);
nor U20530 (N_20530,N_18204,N_14643);
nor U20531 (N_20531,N_14339,N_15162);
and U20532 (N_20532,N_12600,N_13548);
nand U20533 (N_20533,N_15722,N_18489);
nand U20534 (N_20534,N_17054,N_14986);
and U20535 (N_20535,N_16827,N_13443);
nor U20536 (N_20536,N_15538,N_17906);
nand U20537 (N_20537,N_13865,N_18215);
nand U20538 (N_20538,N_15113,N_15756);
nor U20539 (N_20539,N_17284,N_14666);
nand U20540 (N_20540,N_14572,N_13562);
nand U20541 (N_20541,N_17630,N_14472);
or U20542 (N_20542,N_15409,N_17264);
or U20543 (N_20543,N_14839,N_16011);
or U20544 (N_20544,N_13497,N_18038);
nand U20545 (N_20545,N_16883,N_16914);
nor U20546 (N_20546,N_14224,N_17499);
nand U20547 (N_20547,N_13667,N_16775);
xor U20548 (N_20548,N_15090,N_13600);
nor U20549 (N_20549,N_17878,N_13909);
and U20550 (N_20550,N_17333,N_14807);
xor U20551 (N_20551,N_13033,N_17491);
xor U20552 (N_20552,N_15625,N_18435);
nand U20553 (N_20553,N_17457,N_18591);
nor U20554 (N_20554,N_13598,N_14083);
nand U20555 (N_20555,N_13544,N_16762);
and U20556 (N_20556,N_13289,N_16463);
xnor U20557 (N_20557,N_17739,N_16338);
or U20558 (N_20558,N_17748,N_12678);
or U20559 (N_20559,N_13609,N_14290);
xnor U20560 (N_20560,N_13037,N_14334);
or U20561 (N_20561,N_14559,N_18476);
xor U20562 (N_20562,N_13526,N_14488);
nand U20563 (N_20563,N_17320,N_18607);
and U20564 (N_20564,N_16307,N_13122);
and U20565 (N_20565,N_14390,N_17357);
nor U20566 (N_20566,N_14906,N_15400);
nor U20567 (N_20567,N_17142,N_17081);
or U20568 (N_20568,N_14327,N_16644);
or U20569 (N_20569,N_14148,N_18576);
nand U20570 (N_20570,N_12676,N_18632);
or U20571 (N_20571,N_17596,N_18265);
nor U20572 (N_20572,N_17573,N_12728);
xor U20573 (N_20573,N_18138,N_15448);
xnor U20574 (N_20574,N_12943,N_18412);
nor U20575 (N_20575,N_14739,N_14936);
xor U20576 (N_20576,N_14705,N_17221);
xnor U20577 (N_20577,N_15294,N_14152);
xor U20578 (N_20578,N_17301,N_16750);
nand U20579 (N_20579,N_15048,N_17465);
nand U20580 (N_20580,N_13404,N_17733);
xor U20581 (N_20581,N_15911,N_13242);
or U20582 (N_20582,N_16789,N_18307);
xor U20583 (N_20583,N_13942,N_16295);
nor U20584 (N_20584,N_18539,N_15800);
nand U20585 (N_20585,N_14433,N_16572);
nor U20586 (N_20586,N_16879,N_14040);
xnor U20587 (N_20587,N_17023,N_18327);
xnor U20588 (N_20588,N_13546,N_14977);
and U20589 (N_20589,N_14315,N_17452);
xor U20590 (N_20590,N_14774,N_18558);
and U20591 (N_20591,N_12858,N_17223);
and U20592 (N_20592,N_13614,N_16545);
nor U20593 (N_20593,N_17014,N_12511);
xnor U20594 (N_20594,N_16583,N_16432);
xor U20595 (N_20595,N_17418,N_18545);
xor U20596 (N_20596,N_14014,N_13948);
or U20597 (N_20597,N_13787,N_17477);
nand U20598 (N_20598,N_16291,N_14125);
nor U20599 (N_20599,N_17871,N_16938);
nor U20600 (N_20600,N_13320,N_14387);
or U20601 (N_20601,N_17983,N_16725);
xnor U20602 (N_20602,N_18492,N_14576);
nor U20603 (N_20603,N_16309,N_16498);
xnor U20604 (N_20604,N_14830,N_17326);
nor U20605 (N_20605,N_17122,N_17741);
xor U20606 (N_20606,N_17256,N_15804);
xor U20607 (N_20607,N_16531,N_14238);
xor U20608 (N_20608,N_18550,N_13315);
nor U20609 (N_20609,N_14467,N_18247);
xnor U20610 (N_20610,N_17154,N_14207);
and U20611 (N_20611,N_13532,N_13853);
nand U20612 (N_20612,N_13561,N_16247);
xnor U20613 (N_20613,N_16669,N_14401);
xor U20614 (N_20614,N_13095,N_15877);
and U20615 (N_20615,N_16453,N_15894);
nand U20616 (N_20616,N_18109,N_14649);
xnor U20617 (N_20617,N_14568,N_18437);
nand U20618 (N_20618,N_15777,N_13772);
nor U20619 (N_20619,N_15117,N_13119);
nand U20620 (N_20620,N_17948,N_18244);
nor U20621 (N_20621,N_16184,N_14958);
or U20622 (N_20622,N_17817,N_15303);
nor U20623 (N_20623,N_17300,N_12615);
and U20624 (N_20624,N_17209,N_17233);
nor U20625 (N_20625,N_15474,N_12685);
and U20626 (N_20626,N_14168,N_14969);
nor U20627 (N_20627,N_14736,N_17685);
or U20628 (N_20628,N_15411,N_14595);
xnor U20629 (N_20629,N_14284,N_15441);
and U20630 (N_20630,N_17396,N_18203);
nand U20631 (N_20631,N_17840,N_16616);
nor U20632 (N_20632,N_17930,N_15440);
nor U20633 (N_20633,N_13097,N_16211);
xnor U20634 (N_20634,N_17618,N_17559);
xor U20635 (N_20635,N_17222,N_15941);
or U20636 (N_20636,N_15338,N_13316);
and U20637 (N_20637,N_13516,N_18535);
nor U20638 (N_20638,N_16396,N_18315);
nand U20639 (N_20639,N_14983,N_18191);
and U20640 (N_20640,N_12501,N_14079);
or U20641 (N_20641,N_18113,N_12656);
nor U20642 (N_20642,N_13123,N_15305);
xor U20643 (N_20643,N_16429,N_13376);
and U20644 (N_20644,N_17766,N_17793);
xor U20645 (N_20645,N_17176,N_17673);
xnor U20646 (N_20646,N_16947,N_13193);
nor U20647 (N_20647,N_12910,N_16156);
nand U20648 (N_20648,N_13512,N_14904);
nand U20649 (N_20649,N_17306,N_13475);
and U20650 (N_20650,N_16131,N_13029);
and U20651 (N_20651,N_17283,N_13571);
nand U20652 (N_20652,N_15037,N_16615);
nor U20653 (N_20653,N_18478,N_14776);
nor U20654 (N_20654,N_13651,N_15679);
nor U20655 (N_20655,N_18128,N_17401);
nor U20656 (N_20656,N_15683,N_18310);
xor U20657 (N_20657,N_12833,N_12808);
nor U20658 (N_20658,N_15895,N_13400);
nand U20659 (N_20659,N_18120,N_18216);
nor U20660 (N_20660,N_12893,N_18626);
and U20661 (N_20661,N_15244,N_18423);
or U20662 (N_20662,N_14535,N_18222);
nor U20663 (N_20663,N_13391,N_15561);
nor U20664 (N_20664,N_13597,N_14312);
xor U20665 (N_20665,N_17369,N_14225);
or U20666 (N_20666,N_14527,N_12607);
and U20667 (N_20667,N_15077,N_18300);
and U20668 (N_20668,N_13607,N_13968);
nand U20669 (N_20669,N_13010,N_14359);
nand U20670 (N_20670,N_16147,N_18651);
nand U20671 (N_20671,N_16418,N_13357);
and U20672 (N_20672,N_16482,N_14638);
nand U20673 (N_20673,N_15288,N_17028);
nand U20674 (N_20674,N_12575,N_13563);
nand U20675 (N_20675,N_17000,N_17821);
xnor U20676 (N_20676,N_14732,N_15171);
xnor U20677 (N_20677,N_15795,N_16595);
or U20678 (N_20678,N_14210,N_13890);
nand U20679 (N_20679,N_18190,N_13113);
and U20680 (N_20680,N_13818,N_14198);
nor U20681 (N_20681,N_14531,N_13457);
or U20682 (N_20682,N_16127,N_12892);
nand U20683 (N_20683,N_15193,N_12746);
nor U20684 (N_20684,N_18682,N_14903);
or U20685 (N_20685,N_14231,N_14492);
nor U20686 (N_20686,N_15496,N_12955);
or U20687 (N_20687,N_16086,N_15927);
nand U20688 (N_20688,N_14821,N_13775);
nor U20689 (N_20689,N_16913,N_16591);
and U20690 (N_20690,N_13350,N_18463);
xnor U20691 (N_20691,N_14031,N_16114);
and U20692 (N_20692,N_13440,N_15634);
nand U20693 (N_20693,N_12703,N_15397);
xor U20694 (N_20694,N_13003,N_17489);
or U20695 (N_20695,N_17149,N_17165);
nand U20696 (N_20696,N_12683,N_16334);
and U20697 (N_20697,N_16199,N_17869);
and U20698 (N_20698,N_12991,N_15454);
nor U20699 (N_20699,N_16967,N_13741);
nand U20700 (N_20700,N_17416,N_17636);
and U20701 (N_20701,N_13355,N_16093);
xor U20702 (N_20702,N_16397,N_18233);
and U20703 (N_20703,N_17845,N_17190);
or U20704 (N_20704,N_13917,N_16981);
and U20705 (N_20705,N_13161,N_12853);
nand U20706 (N_20706,N_18340,N_13239);
and U20707 (N_20707,N_17044,N_14834);
and U20708 (N_20708,N_17132,N_15362);
and U20709 (N_20709,N_13534,N_15695);
nand U20710 (N_20710,N_15486,N_13816);
or U20711 (N_20711,N_14583,N_13065);
and U20712 (N_20712,N_16571,N_13569);
nor U20713 (N_20713,N_15434,N_12840);
nand U20714 (N_20714,N_15898,N_13781);
or U20715 (N_20715,N_12795,N_12830);
xor U20716 (N_20716,N_17345,N_16969);
and U20717 (N_20717,N_15350,N_12652);
and U20718 (N_20718,N_14804,N_12564);
nor U20719 (N_20719,N_12952,N_16075);
or U20720 (N_20720,N_18121,N_18373);
nor U20721 (N_20721,N_18262,N_13589);
or U20722 (N_20722,N_14909,N_13292);
xor U20723 (N_20723,N_13435,N_16008);
nor U20724 (N_20724,N_16278,N_15905);
nand U20725 (N_20725,N_15791,N_16346);
or U20726 (N_20726,N_17379,N_14200);
or U20727 (N_20727,N_16980,N_13410);
nor U20728 (N_20728,N_17431,N_15259);
and U20729 (N_20729,N_17560,N_18715);
and U20730 (N_20730,N_16794,N_18703);
and U20731 (N_20731,N_14593,N_16515);
nand U20732 (N_20732,N_16456,N_14964);
xor U20733 (N_20733,N_13862,N_13447);
and U20734 (N_20734,N_18620,N_16115);
or U20735 (N_20735,N_18655,N_16167);
nor U20736 (N_20736,N_16837,N_14972);
or U20737 (N_20737,N_17395,N_17458);
or U20738 (N_20738,N_14740,N_13150);
nor U20739 (N_20739,N_17329,N_17981);
or U20740 (N_20740,N_13956,N_12994);
and U20741 (N_20741,N_16007,N_14592);
nand U20742 (N_20742,N_15292,N_17856);
xnor U20743 (N_20743,N_16100,N_15488);
or U20744 (N_20744,N_16327,N_14660);
nor U20745 (N_20745,N_16677,N_13344);
nor U20746 (N_20746,N_14715,N_15638);
xnor U20747 (N_20747,N_15079,N_17775);
nand U20748 (N_20748,N_18155,N_18343);
or U20749 (N_20749,N_16779,N_12572);
or U20750 (N_20750,N_13181,N_17696);
nor U20751 (N_20751,N_17309,N_17686);
or U20752 (N_20752,N_16379,N_17034);
xnor U20753 (N_20753,N_17943,N_16275);
nand U20754 (N_20754,N_13723,N_16364);
and U20755 (N_20755,N_14819,N_18053);
or U20756 (N_20756,N_18443,N_13783);
and U20757 (N_20757,N_15779,N_18671);
or U20758 (N_20758,N_13875,N_18491);
and U20759 (N_20759,N_15215,N_16884);
xnor U20760 (N_20760,N_15626,N_16107);
and U20761 (N_20761,N_14486,N_18698);
or U20762 (N_20762,N_15871,N_16524);
xnor U20763 (N_20763,N_18304,N_16408);
or U20764 (N_20764,N_13711,N_18590);
and U20765 (N_20765,N_13538,N_18737);
nor U20766 (N_20766,N_17207,N_14851);
xor U20767 (N_20767,N_13262,N_15147);
and U20768 (N_20768,N_16503,N_18102);
and U20769 (N_20769,N_13465,N_15060);
nand U20770 (N_20770,N_15431,N_18256);
or U20771 (N_20771,N_18538,N_14800);
and U20772 (N_20772,N_17671,N_17255);
and U20773 (N_20773,N_14423,N_15072);
nor U20774 (N_20774,N_16420,N_15192);
nand U20775 (N_20775,N_15891,N_18452);
and U20776 (N_20776,N_16301,N_18305);
nor U20777 (N_20777,N_16025,N_15334);
or U20778 (N_20778,N_16442,N_12935);
nor U20779 (N_20779,N_17723,N_15524);
nor U20780 (N_20780,N_14675,N_12967);
nor U20781 (N_20781,N_17985,N_16260);
and U20782 (N_20782,N_14344,N_12982);
or U20783 (N_20783,N_14912,N_15558);
and U20784 (N_20784,N_14506,N_16547);
nand U20785 (N_20785,N_13924,N_12681);
nand U20786 (N_20786,N_14429,N_13882);
nand U20787 (N_20787,N_14389,N_12906);
nand U20788 (N_20788,N_16380,N_17205);
or U20789 (N_20789,N_13896,N_17577);
nand U20790 (N_20790,N_13629,N_12551);
or U20791 (N_20791,N_15602,N_12611);
nor U20792 (N_20792,N_18198,N_17571);
or U20793 (N_20793,N_14959,N_17768);
or U20794 (N_20794,N_16639,N_13099);
nor U20795 (N_20795,N_17367,N_17607);
nand U20796 (N_20796,N_15989,N_15123);
or U20797 (N_20797,N_12854,N_14308);
nand U20798 (N_20798,N_18385,N_17684);
xor U20799 (N_20799,N_16326,N_16399);
xor U20800 (N_20800,N_16083,N_16590);
xnor U20801 (N_20801,N_17202,N_16771);
and U20802 (N_20802,N_14324,N_13022);
and U20803 (N_20803,N_17555,N_14012);
nand U20804 (N_20804,N_15231,N_17955);
nor U20805 (N_20805,N_13916,N_16568);
and U20806 (N_20806,N_16907,N_15568);
xor U20807 (N_20807,N_15885,N_13811);
and U20808 (N_20808,N_16487,N_13154);
nand U20809 (N_20809,N_18472,N_18143);
nor U20810 (N_20810,N_14542,N_15653);
xnor U20811 (N_20811,N_18543,N_13672);
xnor U20812 (N_20812,N_16931,N_16855);
and U20813 (N_20813,N_16598,N_13759);
or U20814 (N_20814,N_16267,N_14915);
xor U20815 (N_20815,N_14258,N_13971);
or U20816 (N_20816,N_14588,N_18574);
xor U20817 (N_20817,N_13270,N_15842);
nand U20818 (N_20818,N_14460,N_12663);
xnor U20819 (N_20819,N_13702,N_16039);
nor U20820 (N_20820,N_16608,N_14602);
nor U20821 (N_20821,N_15314,N_12554);
nor U20822 (N_20822,N_17713,N_15345);
nand U20823 (N_20823,N_14537,N_13864);
and U20824 (N_20824,N_14833,N_13228);
and U20825 (N_20825,N_13303,N_15990);
nand U20826 (N_20826,N_17246,N_17391);
xor U20827 (N_20827,N_12638,N_17598);
and U20828 (N_20828,N_13420,N_14237);
and U20829 (N_20829,N_14384,N_15086);
nor U20830 (N_20830,N_18376,N_17140);
and U20831 (N_20831,N_16908,N_15808);
xnor U20832 (N_20832,N_14455,N_12850);
nor U20833 (N_20833,N_15980,N_14720);
xnor U20834 (N_20834,N_12914,N_14408);
or U20835 (N_20835,N_16504,N_16576);
nand U20836 (N_20836,N_13825,N_16259);
xor U20837 (N_20837,N_13654,N_15450);
nor U20838 (N_20838,N_17913,N_17374);
nor U20839 (N_20839,N_18646,N_13567);
xor U20840 (N_20840,N_15105,N_13477);
nor U20841 (N_20841,N_15327,N_16085);
or U20842 (N_20842,N_17517,N_17982);
nand U20843 (N_20843,N_12569,N_12961);
xnor U20844 (N_20844,N_17002,N_18339);
or U20845 (N_20845,N_18411,N_15092);
xor U20846 (N_20846,N_14924,N_16457);
nor U20847 (N_20847,N_15359,N_16448);
or U20848 (N_20848,N_14626,N_13908);
nand U20849 (N_20849,N_17094,N_15571);
nor U20850 (N_20850,N_15420,N_15372);
or U20851 (N_20851,N_14792,N_17114);
nor U20852 (N_20852,N_15547,N_17929);
or U20853 (N_20853,N_15406,N_16602);
nor U20854 (N_20854,N_14128,N_13347);
xor U20855 (N_20855,N_18466,N_14869);
nand U20856 (N_20856,N_18386,N_16496);
nand U20857 (N_20857,N_14072,N_18565);
nor U20858 (N_20858,N_13750,N_12897);
nand U20859 (N_20859,N_16055,N_17881);
xor U20860 (N_20860,N_14728,N_17117);
xor U20861 (N_20861,N_16473,N_17886);
or U20862 (N_20862,N_13642,N_17708);
or U20863 (N_20863,N_14624,N_13552);
nor U20864 (N_20864,N_13218,N_16382);
nand U20865 (N_20865,N_14451,N_17623);
xnor U20866 (N_20866,N_13734,N_12694);
and U20867 (N_20867,N_16160,N_18071);
and U20868 (N_20868,N_13060,N_15291);
or U20869 (N_20869,N_18512,N_18674);
xnor U20870 (N_20870,N_17771,N_15953);
or U20871 (N_20871,N_16316,N_17158);
xor U20872 (N_20872,N_15741,N_13577);
or U20873 (N_20873,N_13800,N_14764);
and U20874 (N_20874,N_14661,N_17884);
and U20875 (N_20875,N_18670,N_17183);
and U20876 (N_20876,N_13768,N_17141);
nand U20877 (N_20877,N_14333,N_18129);
or U20878 (N_20878,N_14974,N_14555);
xnor U20879 (N_20879,N_17179,N_16569);
and U20880 (N_20880,N_15505,N_12949);
nor U20881 (N_20881,N_18379,N_16421);
or U20882 (N_20882,N_16046,N_12988);
nor U20883 (N_20883,N_17730,N_16911);
nor U20884 (N_20884,N_14875,N_17828);
nand U20885 (N_20885,N_17245,N_13296);
nand U20886 (N_20886,N_16842,N_17232);
and U20887 (N_20887,N_15323,N_14616);
nor U20888 (N_20888,N_13090,N_13486);
nor U20889 (N_20889,N_18450,N_14292);
nand U20890 (N_20890,N_13234,N_15461);
and U20891 (N_20891,N_16742,N_13131);
xor U20892 (N_20892,N_15723,N_16191);
nor U20893 (N_20893,N_13648,N_15552);
and U20894 (N_20894,N_13757,N_15614);
xnor U20895 (N_20895,N_14253,N_13625);
and U20896 (N_20896,N_13324,N_17064);
nor U20897 (N_20897,N_16570,N_12512);
xnor U20898 (N_20898,N_15435,N_14961);
xnor U20899 (N_20899,N_17816,N_17830);
or U20900 (N_20900,N_13880,N_17237);
or U20901 (N_20901,N_17875,N_16579);
or U20902 (N_20902,N_13386,N_14985);
or U20903 (N_20903,N_16782,N_18287);
nor U20904 (N_20904,N_15481,N_16484);
xnor U20905 (N_20905,N_14355,N_16578);
and U20906 (N_20906,N_15855,N_13377);
and U20907 (N_20907,N_18146,N_16465);
nor U20908 (N_20908,N_17552,N_13185);
nor U20909 (N_20909,N_17286,N_13550);
nand U20910 (N_20910,N_16761,N_14921);
nor U20911 (N_20911,N_14187,N_12758);
or U20912 (N_20912,N_15810,N_13295);
xnor U20913 (N_20913,N_13127,N_16219);
nor U20914 (N_20914,N_17959,N_17778);
nor U20915 (N_20915,N_14509,N_13836);
nand U20916 (N_20916,N_15378,N_12689);
nor U20917 (N_20917,N_15164,N_13393);
xor U20918 (N_20918,N_17085,N_13606);
and U20919 (N_20919,N_16395,N_16216);
xnor U20920 (N_20920,N_17633,N_18669);
or U20921 (N_20921,N_18439,N_14349);
nand U20922 (N_20922,N_13881,N_16733);
xnor U20923 (N_20923,N_18649,N_17163);
nand U20924 (N_20924,N_16403,N_14473);
or U20925 (N_20925,N_14727,N_14902);
or U20926 (N_20926,N_15154,N_18612);
nor U20927 (N_20927,N_18057,N_17136);
nand U20928 (N_20928,N_18503,N_16325);
xor U20929 (N_20929,N_16873,N_17755);
nor U20930 (N_20930,N_13586,N_14061);
xnor U20931 (N_20931,N_16718,N_15416);
xor U20932 (N_20932,N_12633,N_18174);
nor U20933 (N_20933,N_18200,N_17917);
nand U20934 (N_20934,N_14845,N_13177);
xor U20935 (N_20935,N_13091,N_15628);
and U20936 (N_20936,N_17099,N_14192);
nand U20937 (N_20937,N_15040,N_15058);
or U20938 (N_20938,N_18676,N_16581);
or U20939 (N_20939,N_13949,N_13367);
or U20940 (N_20940,N_14578,N_18397);
nand U20941 (N_20941,N_15367,N_16895);
or U20942 (N_20942,N_14269,N_14299);
nand U20943 (N_20943,N_12801,N_13343);
xor U20944 (N_20944,N_17992,N_14189);
and U20945 (N_20945,N_18258,N_13210);
or U20946 (N_20946,N_14768,N_12936);
nor U20947 (N_20947,N_13521,N_14544);
and U20948 (N_20948,N_17059,N_13619);
nor U20949 (N_20949,N_14957,N_17511);
or U20950 (N_20950,N_13286,N_15926);
or U20951 (N_20951,N_16142,N_16347);
nor U20952 (N_20952,N_14539,N_16188);
and U20953 (N_20953,N_18041,N_16535);
xnor U20954 (N_20954,N_17949,N_17029);
and U20955 (N_20955,N_18358,N_17792);
and U20956 (N_20956,N_18573,N_18167);
and U20957 (N_20957,N_14261,N_14827);
nand U20958 (N_20958,N_15648,N_15379);
nand U20959 (N_20959,N_17617,N_14272);
or U20960 (N_20960,N_16735,N_14734);
or U20961 (N_20961,N_17591,N_16942);
xnor U20962 (N_20962,N_17991,N_16668);
nand U20963 (N_20963,N_12596,N_17107);
nor U20964 (N_20964,N_15423,N_17016);
nor U20965 (N_20965,N_13506,N_13192);
or U20966 (N_20966,N_16043,N_12829);
nor U20967 (N_20967,N_15010,N_16263);
xnor U20968 (N_20968,N_15250,N_14907);
or U20969 (N_20969,N_17031,N_12751);
or U20970 (N_20970,N_13166,N_14813);
nor U20971 (N_20971,N_18123,N_13110);
or U20972 (N_20972,N_15543,N_13910);
or U20973 (N_20973,N_12835,N_15730);
or U20974 (N_20974,N_17065,N_15439);
xor U20975 (N_20975,N_16368,N_16200);
xnor U20976 (N_20976,N_14069,N_13213);
or U20977 (N_20977,N_15986,N_18616);
nor U20978 (N_20978,N_14013,N_16645);
xnor U20979 (N_20979,N_15915,N_17606);
and U20980 (N_20980,N_15320,N_17562);
nand U20981 (N_20981,N_13572,N_15839);
or U20982 (N_20982,N_13793,N_12913);
or U20983 (N_20983,N_17362,N_13999);
nor U20984 (N_20984,N_17803,N_17547);
nand U20985 (N_20985,N_13584,N_12841);
and U20986 (N_20986,N_17193,N_13854);
nor U20987 (N_20987,N_13353,N_12711);
nand U20988 (N_20988,N_18254,N_14747);
xor U20989 (N_20989,N_13251,N_18603);
nand U20990 (N_20990,N_15668,N_17298);
nor U20991 (N_20991,N_15869,N_18248);
or U20992 (N_20992,N_14905,N_18346);
and U20993 (N_20993,N_14689,N_16812);
nand U20994 (N_20994,N_14112,N_13274);
nor U20995 (N_20995,N_12927,N_18623);
nand U20996 (N_20996,N_14886,N_17100);
and U20997 (N_20997,N_13372,N_16140);
nand U20998 (N_20998,N_18664,N_16940);
or U20999 (N_20999,N_18051,N_17058);
nor U21000 (N_21000,N_17497,N_18293);
nor U21001 (N_21001,N_13250,N_13610);
or U21002 (N_21002,N_17942,N_16710);
nand U21003 (N_21003,N_16339,N_15337);
xnor U21004 (N_21004,N_16682,N_15018);
nand U21005 (N_21005,N_17071,N_18391);
and U21006 (N_21006,N_15762,N_14103);
xor U21007 (N_21007,N_12874,N_17961);
and U21008 (N_21008,N_16698,N_13826);
xor U21009 (N_21009,N_13148,N_17102);
nor U21010 (N_21010,N_14348,N_17656);
nand U21011 (N_21011,N_16059,N_13640);
xnor U21012 (N_21012,N_17936,N_15276);
nand U21013 (N_21013,N_14621,N_16053);
xor U21014 (N_21014,N_14860,N_18153);
nor U21015 (N_21015,N_13111,N_14726);
or U21016 (N_21016,N_18723,N_15838);
nand U21017 (N_21017,N_15383,N_14853);
nand U21018 (N_21018,N_14664,N_14209);
nor U21019 (N_21019,N_15459,N_12870);
or U21020 (N_21020,N_18488,N_13765);
nor U21021 (N_21021,N_18740,N_17120);
and U21022 (N_21022,N_15858,N_13989);
or U21023 (N_21023,N_13988,N_14456);
nand U21024 (N_21024,N_14984,N_14953);
xor U21025 (N_21025,N_12903,N_12536);
nor U21026 (N_21026,N_17813,N_17692);
nand U21027 (N_21027,N_13698,N_14268);
and U21028 (N_21028,N_17740,N_17443);
and U21029 (N_21029,N_14392,N_16921);
nor U21030 (N_21030,N_17354,N_17659);
nor U21031 (N_21031,N_16203,N_14374);
nand U21032 (N_21032,N_14564,N_13243);
xnor U21033 (N_21033,N_13852,N_18313);
or U21034 (N_21034,N_14658,N_18354);
or U21035 (N_21035,N_15472,N_12677);
and U21036 (N_21036,N_15544,N_13128);
nor U21037 (N_21037,N_16148,N_16690);
nand U21038 (N_21038,N_15321,N_12987);
nand U21039 (N_21039,N_14427,N_16625);
or U21040 (N_21040,N_15228,N_13689);
and U21041 (N_21041,N_16826,N_15720);
nand U21042 (N_21042,N_16439,N_13137);
or U21043 (N_21043,N_13798,N_13684);
nand U21044 (N_21044,N_14053,N_15309);
nor U21045 (N_21045,N_12533,N_13268);
nor U21046 (N_21046,N_15998,N_18396);
or U21047 (N_21047,N_17702,N_14481);
nor U21048 (N_21048,N_16355,N_15051);
xor U21049 (N_21049,N_13467,N_15121);
and U21050 (N_21050,N_12992,N_13265);
xnor U21051 (N_21051,N_18067,N_17115);
and U21052 (N_21052,N_15778,N_14228);
and U21053 (N_21053,N_18618,N_13533);
or U21054 (N_21054,N_14529,N_14055);
xnor U21055 (N_21055,N_13430,N_18154);
nand U21056 (N_21056,N_16758,N_13580);
xnor U21057 (N_21057,N_13876,N_14603);
nor U21058 (N_21058,N_16412,N_14409);
and U21059 (N_21059,N_18241,N_18196);
or U21060 (N_21060,N_13627,N_13153);
and U21061 (N_21061,N_16763,N_13990);
and U21062 (N_21062,N_15188,N_18318);
nand U21063 (N_21063,N_15233,N_14323);
nand U21064 (N_21064,N_15522,N_18206);
nor U21065 (N_21065,N_14141,N_18691);
nand U21066 (N_21066,N_13473,N_16222);
and U21067 (N_21067,N_15422,N_13556);
and U21068 (N_21068,N_12868,N_14919);
nand U21069 (N_21069,N_18387,N_17212);
nand U21070 (N_21070,N_17996,N_14241);
or U21071 (N_21071,N_14440,N_12785);
and U21072 (N_21072,N_12754,N_16712);
or U21073 (N_21073,N_16957,N_17916);
nor U21074 (N_21074,N_17208,N_16415);
and U21075 (N_21075,N_14829,N_17866);
xor U21076 (N_21076,N_17442,N_13103);
nand U21077 (N_21077,N_16681,N_16234);
nand U21078 (N_21078,N_17187,N_12518);
xor U21079 (N_21079,N_14656,N_18337);
and U21080 (N_21080,N_15725,N_14051);
and U21081 (N_21081,N_13254,N_15031);
nand U21082 (N_21082,N_18404,N_12852);
or U21083 (N_21083,N_13491,N_15028);
nand U21084 (N_21084,N_18361,N_15047);
xnor U21085 (N_21085,N_15027,N_12898);
and U21086 (N_21086,N_15595,N_15277);
and U21087 (N_21087,N_14118,N_16671);
or U21088 (N_21088,N_18581,N_16807);
nand U21089 (N_21089,N_14815,N_12556);
nor U21090 (N_21090,N_16006,N_13424);
and U21091 (N_21091,N_15655,N_12704);
nor U21092 (N_21092,N_13676,N_15261);
nor U21093 (N_21093,N_16798,N_17503);
nor U21094 (N_21094,N_16719,N_12692);
xnor U21095 (N_21095,N_13151,N_16454);
and U21096 (N_21096,N_13088,N_15358);
nor U21097 (N_21097,N_17342,N_15647);
and U21098 (N_21098,N_15101,N_14050);
xor U21099 (N_21099,N_18348,N_14998);
nor U21100 (N_21100,N_17879,N_15572);
nand U21101 (N_21101,N_18181,N_18012);
nand U21102 (N_21102,N_18441,N_17954);
nand U21103 (N_21103,N_18332,N_13493);
and U21104 (N_21104,N_18433,N_13634);
or U21105 (N_21105,N_16932,N_16292);
nor U21106 (N_21106,N_16449,N_14746);
or U21107 (N_21107,N_17691,N_12730);
nor U21108 (N_21108,N_15163,N_18170);
nand U21109 (N_21109,N_16566,N_14910);
and U21110 (N_21110,N_15697,N_18630);
nand U21111 (N_21111,N_16280,N_18701);
nand U21112 (N_21112,N_16532,N_15514);
nor U21113 (N_21113,N_16126,N_16022);
xnor U21114 (N_21114,N_13142,N_18139);
xor U21115 (N_21115,N_17512,N_17239);
nand U21116 (N_21116,N_17013,N_13554);
or U21117 (N_21117,N_14174,N_14422);
nand U21118 (N_21118,N_15904,N_17567);
xnor U21119 (N_21119,N_17920,N_18136);
xor U21120 (N_21120,N_13362,N_17172);
xnor U21121 (N_21121,N_15195,N_14793);
and U21122 (N_21122,N_15961,N_17137);
xor U21123 (N_21123,N_16560,N_14480);
nor U21124 (N_21124,N_18301,N_13018);
xnor U21125 (N_21125,N_13983,N_15862);
or U21126 (N_21126,N_16112,N_12532);
or U21127 (N_21127,N_16638,N_18458);
xor U21128 (N_21128,N_14162,N_16390);
and U21129 (N_21129,N_17479,N_12957);
and U21130 (N_21130,N_15549,N_18028);
nand U21131 (N_21131,N_14861,N_14183);
and U21132 (N_21132,N_15863,N_14655);
nor U21133 (N_21133,N_14862,N_15247);
nand U21134 (N_21134,N_18556,N_15270);
xor U21135 (N_21135,N_14046,N_17890);
and U21136 (N_21136,N_18383,N_16804);
nand U21137 (N_21137,N_15346,N_14020);
xnor U21138 (N_21138,N_13249,N_15573);
nor U21139 (N_21139,N_17557,N_18380);
nand U21140 (N_21140,N_15575,N_14495);
nand U21141 (N_21141,N_15606,N_13159);
nand U21142 (N_21142,N_14751,N_16157);
xnor U21143 (N_21143,N_14419,N_16935);
xnor U21144 (N_21144,N_17787,N_14252);
nor U21145 (N_21145,N_15824,N_18021);
nor U21146 (N_21146,N_13313,N_15065);
nand U21147 (N_21147,N_15396,N_18061);
nor U21148 (N_21148,N_13449,N_14528);
and U21149 (N_21149,N_14078,N_14842);
nand U21150 (N_21150,N_13031,N_15924);
nor U21151 (N_21151,N_15992,N_18661);
xor U21152 (N_21152,N_17980,N_15737);
nor U21153 (N_21153,N_13639,N_15289);
nor U21154 (N_21154,N_12925,N_16238);
or U21155 (N_21155,N_17083,N_14099);
nand U21156 (N_21156,N_16480,N_14194);
xor U21157 (N_21157,N_16661,N_18566);
or U21158 (N_21158,N_13588,N_15146);
and U21159 (N_21159,N_17776,N_18278);
xor U21160 (N_21160,N_14534,N_16854);
and U21161 (N_21161,N_16101,N_16333);
nor U21162 (N_21162,N_15939,N_13231);
xor U21163 (N_21163,N_13396,N_16833);
and U21164 (N_21164,N_17521,N_14016);
xor U21165 (N_21165,N_13162,N_13241);
or U21166 (N_21166,N_17152,N_12845);
or U21167 (N_21167,N_18717,N_12908);
or U21168 (N_21168,N_13149,N_12741);
and U21169 (N_21169,N_17025,N_17742);
xor U21170 (N_21170,N_16582,N_17904);
xnor U21171 (N_21171,N_18544,N_14922);
and U21172 (N_21172,N_16282,N_12923);
nor U21173 (N_21173,N_14175,N_14663);
xor U21174 (N_21174,N_18652,N_15389);
xor U21175 (N_21175,N_13124,N_14780);
or U21176 (N_21176,N_16118,N_12778);
nor U21177 (N_21177,N_14787,N_14587);
and U21178 (N_21178,N_13539,N_17315);
or U21179 (N_21179,N_18342,N_18744);
and U21180 (N_21180,N_17535,N_14291);
xnor U21181 (N_21181,N_15831,N_17096);
or U21182 (N_21182,N_18694,N_14487);
nand U21183 (N_21183,N_14468,N_12765);
xor U21184 (N_21184,N_17127,N_18708);
nor U21185 (N_21185,N_16233,N_14763);
or U21186 (N_21186,N_15053,N_14321);
xor U21187 (N_21187,N_17075,N_13080);
and U21188 (N_21188,N_12594,N_17795);
xnor U21189 (N_21189,N_13518,N_18426);
and U21190 (N_21190,N_14094,N_13728);
or U21191 (N_21191,N_17576,N_18428);
nand U21192 (N_21192,N_18604,N_18532);
or U21193 (N_21193,N_14096,N_15007);
and U21194 (N_21194,N_17353,N_15977);
or U21195 (N_21195,N_15176,N_15984);
nand U21196 (N_21196,N_13202,N_17762);
xor U21197 (N_21197,N_14622,N_15586);
nand U21198 (N_21198,N_14757,N_14980);
nor U21199 (N_21199,N_14404,N_12793);
and U21200 (N_21200,N_13352,N_16977);
and U21201 (N_21201,N_12981,N_14693);
xor U21202 (N_21202,N_16513,N_12737);
and U21203 (N_21203,N_17455,N_17303);
and U21204 (N_21204,N_15282,N_16176);
and U21205 (N_21205,N_16985,N_15960);
xnor U21206 (N_21206,N_15082,N_13361);
or U21207 (N_21207,N_15666,N_14737);
xor U21208 (N_21208,N_18005,N_16027);
nand U21209 (N_21209,N_15315,N_15050);
and U21210 (N_21210,N_14067,N_13334);
xor U21211 (N_21211,N_13557,N_14047);
nor U21212 (N_21212,N_17421,N_16391);
or U21213 (N_21213,N_18164,N_14042);
nand U21214 (N_21214,N_13605,N_13280);
nand U21215 (N_21215,N_13409,N_12637);
nor U21216 (N_21216,N_17483,N_14082);
nor U21217 (N_21217,N_18282,N_17928);
or U21218 (N_21218,N_15727,N_16445);
nand U21219 (N_21219,N_14499,N_16462);
xnor U21220 (N_21220,N_16253,N_17133);
or U21221 (N_21221,N_15364,N_12570);
nor U21222 (N_21222,N_16593,N_17697);
and U21223 (N_21223,N_13425,N_12620);
xor U21224 (N_21224,N_14941,N_14627);
and U21225 (N_21225,N_15357,N_15835);
and U21226 (N_21226,N_16890,N_18635);
and U21227 (N_21227,N_17655,N_17801);
xor U21228 (N_21228,N_14156,N_14009);
or U21229 (N_21229,N_17718,N_15527);
or U21230 (N_21230,N_17106,N_17462);
or U21231 (N_21231,N_14376,N_15820);
or U21232 (N_21232,N_18157,N_14490);
xnor U21233 (N_21233,N_18111,N_14318);
nand U21234 (N_21234,N_14692,N_15619);
nor U21235 (N_21235,N_14005,N_15881);
xnor U21236 (N_21236,N_16791,N_15380);
nand U21237 (N_21237,N_15957,N_16999);
nand U21238 (N_21238,N_17900,N_15124);
or U21239 (N_21239,N_16213,N_18078);
and U21240 (N_21240,N_17288,N_17186);
nor U21241 (N_21241,N_17371,N_14402);
nor U21242 (N_21242,N_14520,N_17746);
nor U21243 (N_21243,N_15471,N_17641);
xor U21244 (N_21244,N_18070,N_15169);
and U21245 (N_21245,N_14882,N_13204);
or U21246 (N_21246,N_14199,N_18345);
nor U21247 (N_21247,N_12786,N_17863);
nor U21248 (N_21248,N_18419,N_16493);
xor U21249 (N_21249,N_14721,N_13808);
or U21250 (N_21250,N_13098,N_18514);
and U21251 (N_21251,N_15221,N_17972);
or U21252 (N_21252,N_13842,N_16001);
and U21253 (N_21253,N_14577,N_16324);
nand U21254 (N_21254,N_16205,N_14805);
nand U21255 (N_21255,N_18679,N_12973);
nor U21256 (N_21256,N_15541,N_14575);
xnor U21257 (N_21257,N_12930,N_15203);
xnor U21258 (N_21258,N_14471,N_17514);
or U21259 (N_21259,N_17578,N_15861);
and U21260 (N_21260,N_16438,N_15950);
and U21261 (N_21261,N_17226,N_17011);
xor U21262 (N_21262,N_13285,N_14967);
or U21263 (N_21263,N_15368,N_17831);
xnor U21264 (N_21264,N_16424,N_14700);
and U21265 (N_21265,N_15470,N_12966);
nor U21266 (N_21266,N_17274,N_13617);
nand U21267 (N_21267,N_17749,N_18587);
or U21268 (N_21268,N_14369,N_18068);
and U21269 (N_21269,N_16444,N_15533);
xnor U21270 (N_21270,N_14282,N_15024);
nand U21271 (N_21271,N_12714,N_18063);
and U21272 (N_21272,N_13030,N_13920);
nor U21273 (N_21273,N_17994,N_16099);
or U21274 (N_21274,N_13977,N_15167);
nand U21275 (N_21275,N_14153,N_17543);
and U21276 (N_21276,N_13806,N_17063);
nand U21277 (N_21277,N_17519,N_16431);
xnor U21278 (N_21278,N_12560,N_14412);
nand U21279 (N_21279,N_16294,N_13979);
xor U21280 (N_21280,N_13172,N_17200);
nor U21281 (N_21281,N_14213,N_17242);
and U21282 (N_21282,N_18568,N_17564);
nor U21283 (N_21283,N_14952,N_16353);
xnor U21284 (N_21284,N_17887,N_17709);
and U21285 (N_21285,N_17012,N_15451);
and U21286 (N_21286,N_15269,N_15223);
or U21287 (N_21287,N_14142,N_16752);
nand U21288 (N_21288,N_13330,N_13016);
and U21289 (N_21289,N_14037,N_17385);
nand U21290 (N_21290,N_15623,N_14937);
xor U21291 (N_21291,N_17932,N_12669);
nor U21292 (N_21292,N_18208,N_13140);
xor U21293 (N_21293,N_14159,N_18046);
nand U21294 (N_21294,N_15026,N_17393);
xor U21295 (N_21295,N_16994,N_14590);
xor U21296 (N_21296,N_14080,N_14668);
and U21297 (N_21297,N_17337,N_13766);
nor U21298 (N_21298,N_12956,N_18599);
and U21299 (N_21299,N_16618,N_17629);
nor U21300 (N_21300,N_13056,N_15566);
and U21301 (N_21301,N_18536,N_16070);
nor U21302 (N_21302,N_13620,N_16224);
and U21303 (N_21303,N_14678,N_12553);
and U21304 (N_21304,N_14676,N_14802);
nor U21305 (N_21305,N_18742,N_17860);
and U21306 (N_21306,N_16386,N_12540);
xor U21307 (N_21307,N_12716,N_17022);
or U21308 (N_21308,N_13790,N_15335);
xnor U21309 (N_21309,N_12682,N_17978);
and U21310 (N_21310,N_14133,N_16694);
nor U21311 (N_21311,N_13272,N_17340);
nor U21312 (N_21312,N_16519,N_14766);
nand U21313 (N_21313,N_13700,N_16787);
xnor U21314 (N_21314,N_13682,N_15703);
nand U21315 (N_21315,N_15348,N_15564);
nor U21316 (N_21316,N_17139,N_15452);
and U21317 (N_21317,N_16963,N_15428);
xor U21318 (N_21318,N_17897,N_13302);
nand U21319 (N_21319,N_12508,N_17734);
and U21320 (N_21320,N_16714,N_17076);
nand U21321 (N_21321,N_18395,N_14810);
xnor U21322 (N_21322,N_16098,N_13951);
or U21323 (N_21323,N_16483,N_17090);
and U21324 (N_21324,N_16696,N_16490);
nor U21325 (N_21325,N_16154,N_15883);
and U21326 (N_21326,N_14753,N_15141);
nor U21327 (N_21327,N_18357,N_16340);
and U21328 (N_21328,N_15445,N_17411);
and U21329 (N_21329,N_12860,N_18600);
or U21330 (N_21330,N_14999,N_14215);
xor U21331 (N_21331,N_15473,N_12653);
xor U21332 (N_21332,N_14798,N_17089);
and U21333 (N_21333,N_14724,N_15447);
nand U21334 (N_21334,N_15460,N_16060);
or U21335 (N_21335,N_18240,N_15567);
or U21336 (N_21336,N_14759,N_17967);
xnor U21337 (N_21337,N_14711,N_17704);
or U21338 (N_21338,N_15799,N_14163);
xnor U21339 (N_21339,N_14115,N_13199);
nand U21340 (N_21340,N_18084,N_16512);
and U21341 (N_21341,N_14331,N_14930);
nor U21342 (N_21342,N_14100,N_13345);
xnor U21343 (N_21343,N_13767,N_16972);
nand U21344 (N_21344,N_14030,N_18023);
or U21345 (N_21345,N_12744,N_16387);
or U21346 (N_21346,N_15283,N_18350);
and U21347 (N_21347,N_15003,N_12789);
or U21348 (N_21348,N_18438,N_14760);
xnor U21349 (N_21349,N_12873,N_13749);
nand U21350 (N_21350,N_16612,N_16369);
and U21351 (N_21351,N_13027,N_14068);
and U21352 (N_21352,N_16747,N_17682);
and U21353 (N_21353,N_18455,N_17679);
xnor U21354 (N_21354,N_12849,N_17331);
nor U21355 (N_21355,N_15266,N_14662);
and U21356 (N_21356,N_13957,N_12579);
and U21357 (N_21357,N_16730,N_13830);
nand U21358 (N_21358,N_14130,N_13686);
or U21359 (N_21359,N_17145,N_15536);
nand U21360 (N_21360,N_12826,N_15832);
xnor U21361 (N_21361,N_15681,N_13553);
xor U21362 (N_21362,N_15747,N_15085);
nor U21363 (N_21363,N_13636,N_17481);
nand U21364 (N_21364,N_17439,N_15557);
nor U21365 (N_21365,N_17561,N_13530);
and U21366 (N_21366,N_16562,N_17036);
or U21367 (N_21367,N_13570,N_12749);
nand U21368 (N_21368,N_13380,N_12573);
or U21369 (N_21369,N_17488,N_12926);
or U21370 (N_21370,N_15931,N_14229);
xor U21371 (N_21371,N_13100,N_17124);
and U21372 (N_21372,N_12659,N_13898);
and U21373 (N_21373,N_17501,N_18610);
or U21374 (N_21374,N_18381,N_14461);
nor U21375 (N_21375,N_14271,N_14840);
and U21376 (N_21376,N_14594,N_17118);
nor U21377 (N_21377,N_16430,N_17409);
and U21378 (N_21378,N_17769,N_15685);
nand U21379 (N_21379,N_13735,N_16264);
or U21380 (N_21380,N_16174,N_16825);
nand U21381 (N_21381,N_15102,N_17580);
nor U21382 (N_21382,N_13365,N_15809);
or U21383 (N_21383,N_13611,N_17159);
or U21384 (N_21384,N_13064,N_17420);
xor U21385 (N_21385,N_15521,N_17074);
or U21386 (N_21386,N_13279,N_14558);
nand U21387 (N_21387,N_16622,N_14113);
nor U21388 (N_21388,N_14552,N_18695);
or U21389 (N_21389,N_12726,N_14222);
and U21390 (N_21390,N_16312,N_16367);
or U21391 (N_21391,N_16171,N_14362);
xnor U21392 (N_21392,N_16753,N_12529);
nor U21393 (N_21393,N_17150,N_18306);
nor U21394 (N_21394,N_16257,N_15316);
or U21395 (N_21395,N_13246,N_17644);
xor U21396 (N_21396,N_15743,N_18141);
and U21397 (N_21397,N_13754,N_18577);
nor U21398 (N_21398,N_17316,N_17486);
or U21399 (N_21399,N_18323,N_15776);
and U21400 (N_21400,N_17534,N_17987);
xor U21401 (N_21401,N_14342,N_14913);
or U21402 (N_21402,N_13026,N_12922);
nand U21403 (N_21403,N_15310,N_15563);
nor U21404 (N_21404,N_18633,N_16015);
xnor U21405 (N_21405,N_18429,N_13829);
xnor U21406 (N_21406,N_14551,N_15205);
and U21407 (N_21407,N_12775,N_17191);
nor U21408 (N_21408,N_18714,N_18125);
nand U21409 (N_21409,N_18169,N_12909);
xor U21410 (N_21410,N_17098,N_15128);
and U21411 (N_21411,N_13460,N_14519);
xnor U21412 (N_21412,N_13220,N_18151);
nor U21413 (N_21413,N_15705,N_13197);
nand U21414 (N_21414,N_14635,N_16304);
xor U21415 (N_21415,N_16886,N_12558);
nor U21416 (N_21416,N_12814,N_17015);
and U21417 (N_21417,N_12846,N_16597);
nand U21418 (N_21418,N_16405,N_17009);
xor U21419 (N_21419,N_16407,N_16555);
and U21420 (N_21420,N_12563,N_12884);
nor U21421 (N_21421,N_13656,N_16270);
and U21422 (N_21422,N_16836,N_13807);
xnor U21423 (N_21423,N_15715,N_17493);
nand U21424 (N_21424,N_14382,N_16500);
xor U21425 (N_21425,N_14538,N_15786);
nand U21426 (N_21426,N_16452,N_13939);
and U21427 (N_21427,N_17594,N_16019);
or U21428 (N_21428,N_16554,N_16193);
or U21429 (N_21429,N_18586,N_14744);
nand U21430 (N_21430,N_13379,N_13085);
xor U21431 (N_21431,N_15651,N_16587);
xnor U21432 (N_21432,N_13594,N_17852);
nand U21433 (N_21433,N_15732,N_17027);
xor U21434 (N_21434,N_17516,N_12916);
nand U21435 (N_21435,N_16878,N_16627);
and U21436 (N_21436,N_14357,N_15932);
or U21437 (N_21437,N_16894,N_13221);
or U21438 (N_21438,N_16868,N_14158);
nand U21439 (N_21439,N_15438,N_13622);
xnor U21440 (N_21440,N_18517,N_18547);
and U21441 (N_21441,N_12698,N_13492);
nor U21442 (N_21442,N_13505,N_12756);
nand U21443 (N_21443,N_18617,N_17582);
nand U21444 (N_21444,N_17020,N_17135);
nor U21445 (N_21445,N_14927,N_16003);
nand U21446 (N_21446,N_16384,N_15702);
xor U21447 (N_21447,N_18232,N_15239);
or U21448 (N_21448,N_15227,N_13488);
nor U21449 (N_21449,N_17549,N_12851);
xor U21450 (N_21450,N_14847,N_14932);
xnor U21451 (N_21451,N_15035,N_16961);
nor U21452 (N_21452,N_18338,N_12565);
nor U21453 (N_21453,N_17669,N_15405);
or U21454 (N_21454,N_12629,N_18467);
nand U21455 (N_21455,N_18451,N_13050);
nor U21456 (N_21456,N_18407,N_14589);
nor U21457 (N_21457,N_15249,N_13079);
or U21458 (N_21458,N_15444,N_18659);
xnor U21459 (N_21459,N_12743,N_13901);
and U21460 (N_21460,N_13671,N_14336);
xnor U21461 (N_21461,N_17908,N_13087);
xnor U21462 (N_21462,N_17539,N_13528);
xnor U21463 (N_21463,N_12647,N_13311);
nor U21464 (N_21464,N_17593,N_12568);
or U21465 (N_21465,N_18688,N_14625);
nand U21466 (N_21466,N_17989,N_13576);
nand U21467 (N_21467,N_18501,N_17631);
or U21468 (N_21468,N_18628,N_17236);
or U21469 (N_21469,N_15083,N_16045);
nor U21470 (N_21470,N_17129,N_14345);
xor U21471 (N_21471,N_16505,N_17351);
nand U21472 (N_21472,N_16056,N_16394);
nor U21473 (N_21473,N_15636,N_12664);
or U21474 (N_21474,N_17250,N_15177);
xnor U21475 (N_21475,N_15041,N_18442);
nor U21476 (N_21476,N_18202,N_12964);
xnor U21477 (N_21477,N_13455,N_14748);
xor U21478 (N_21478,N_15945,N_17789);
and U21479 (N_21479,N_17072,N_17494);
nand U21480 (N_21480,N_18363,N_17589);
nand U21481 (N_21481,N_17123,N_14533);
or U21482 (N_21482,N_16835,N_16845);
and U21483 (N_21483,N_12857,N_16365);
nor U21484 (N_21484,N_12774,N_15555);
and U21485 (N_21485,N_14358,N_17043);
or U21486 (N_21486,N_15686,N_13208);
or U21487 (N_21487,N_16574,N_13071);
nor U21488 (N_21488,N_13558,N_17480);
or U21489 (N_21489,N_15319,N_18734);
nor U21490 (N_21490,N_16033,N_12999);
nand U21491 (N_21491,N_15909,N_15922);
and U21492 (N_21492,N_16670,N_15974);
xnor U21493 (N_21493,N_17291,N_17984);
and U21494 (N_21494,N_12684,N_14574);
or U21495 (N_21495,N_16398,N_12675);
nor U21496 (N_21496,N_14364,N_13937);
nand U21497 (N_21497,N_18564,N_15944);
nor U21498 (N_21498,N_15870,N_13053);
nand U21499 (N_21499,N_16409,N_13075);
or U21500 (N_21500,N_17627,N_13691);
or U21501 (N_21501,N_14034,N_16974);
and U21502 (N_21502,N_13794,N_12699);
xor U21503 (N_21503,N_16577,N_12642);
and U21504 (N_21504,N_17047,N_16318);
or U21505 (N_21505,N_12705,N_15629);
nor U21506 (N_21506,N_12609,N_18484);
nand U21507 (N_21507,N_14300,N_14516);
and U21508 (N_21508,N_17428,N_17241);
and U21509 (N_21509,N_15713,N_13918);
nand U21510 (N_21510,N_16228,N_17834);
xor U21511 (N_21511,N_13799,N_14775);
nor U21512 (N_21512,N_17550,N_14463);
xor U21513 (N_21513,N_14343,N_12631);
nand U21514 (N_21514,N_17654,N_17279);
nand U21515 (N_21515,N_13017,N_16693);
nand U21516 (N_21516,N_17227,N_13712);
nand U21517 (N_21517,N_12680,N_17603);
nand U21518 (N_21518,N_12970,N_14086);
or U21519 (N_21519,N_14585,N_17794);
or U21520 (N_21520,N_13946,N_13366);
xnor U21521 (N_21521,N_15542,N_16028);
or U21522 (N_21522,N_14826,N_17678);
xnor U21523 (N_21523,N_17528,N_12805);
nand U21524 (N_21524,N_18009,N_15424);
nand U21525 (N_21525,N_15689,N_14351);
xor U21526 (N_21526,N_16918,N_16922);
xnor U21527 (N_21527,N_17195,N_14143);
xnor U21528 (N_21528,N_17918,N_12864);
or U21529 (N_21529,N_13325,N_14227);
and U21530 (N_21530,N_15131,N_14454);
and U21531 (N_21531,N_14121,N_12513);
xnor U21532 (N_21532,N_14586,N_18106);
nor U21533 (N_21533,N_18497,N_16777);
and U21534 (N_21534,N_17585,N_14117);
nor U21535 (N_21535,N_18319,N_16311);
nand U21536 (N_21536,N_14893,N_17891);
and U21537 (N_21537,N_17175,N_15996);
xnor U21538 (N_21538,N_16958,N_18277);
nor U21539 (N_21539,N_16080,N_17938);
and U21540 (N_21540,N_15754,N_15967);
nor U21541 (N_21541,N_17826,N_16537);
nor U21542 (N_21542,N_12707,N_13847);
xor U21543 (N_21543,N_15920,N_18117);
xor U21544 (N_21544,N_16847,N_16476);
xnor U21545 (N_21545,N_15142,N_16876);
nor U21546 (N_21546,N_17151,N_15412);
xor U21547 (N_21547,N_13769,N_13623);
and U21548 (N_21548,N_15478,N_12628);
and U21549 (N_21549,N_13083,N_13813);
xor U21550 (N_21550,N_14699,N_16488);
xnor U21551 (N_21551,N_17381,N_16097);
and U21552 (N_21552,N_14188,N_15418);
and U21553 (N_21553,N_15074,N_13970);
nor U21554 (N_21554,N_13462,N_15332);
nand U21555 (N_21555,N_16254,N_14584);
and U21556 (N_21556,N_18382,N_15125);
nor U21557 (N_21557,N_13687,N_17513);
or U21558 (N_21558,N_13693,N_18392);
nor U21559 (N_21559,N_14502,N_13373);
xor U21560 (N_21560,N_18460,N_15516);
and U21561 (N_21561,N_12915,N_17295);
nand U21562 (N_21562,N_18062,N_16643);
xnor U21563 (N_21563,N_14028,N_17214);
and U21564 (N_21564,N_13014,N_17634);
or U21565 (N_21565,N_15173,N_13653);
xor U21566 (N_21566,N_14139,N_16168);
nor U21567 (N_21567,N_18427,N_13838);
nor U21568 (N_21568,N_14178,N_16406);
nand U21569 (N_21569,N_17902,N_16381);
xor U21570 (N_21570,N_15943,N_13051);
nand U21571 (N_21571,N_16746,N_17632);
nor U21572 (N_21572,N_18647,N_13960);
or U21573 (N_21573,N_12627,N_14491);
xnor U21574 (N_21574,N_17270,N_12635);
nor U21575 (N_21575,N_18485,N_16766);
and U21576 (N_21576,N_17760,N_15194);
nor U21577 (N_21577,N_14515,N_15755);
xnor U21578 (N_21578,N_18020,N_13490);
or U21579 (N_21579,N_14947,N_17672);
xnor U21580 (N_21580,N_15865,N_13329);
or U21581 (N_21581,N_18039,N_14007);
and U21582 (N_21582,N_18526,N_13645);
or U21583 (N_21583,N_13675,N_15482);
xor U21584 (N_21584,N_16422,N_12979);
nand U21585 (N_21585,N_16860,N_13374);
nand U21586 (N_21586,N_13189,N_12708);
or U21587 (N_21587,N_15744,N_16924);
or U21588 (N_21588,N_17715,N_13994);
xnor U21589 (N_21589,N_15508,N_15100);
xnor U21590 (N_21590,N_13674,N_13725);
nor U21591 (N_21591,N_15670,N_16754);
and U21592 (N_21592,N_17753,N_14496);
nor U21593 (N_21593,N_17184,N_18378);
nand U21594 (N_21594,N_17626,N_17423);
and U21595 (N_21595,N_16017,N_18468);
or U21596 (N_21596,N_17040,N_15168);
or U21597 (N_21597,N_17505,N_18546);
or U21598 (N_21598,N_17670,N_13555);
or U21599 (N_21599,N_14831,N_18721);
nand U21600 (N_21600,N_12907,N_16239);
nor U21601 (N_21601,N_15466,N_15512);
nand U21602 (N_21602,N_18367,N_17294);
xor U21603 (N_21603,N_14248,N_12525);
or U21604 (N_21604,N_17842,N_17962);
xnor U21605 (N_21605,N_17305,N_16724);
xnor U21606 (N_21606,N_13351,N_13593);
nand U21607 (N_21607,N_14232,N_17487);
xor U21608 (N_21608,N_14982,N_12739);
or U21609 (N_21609,N_14270,N_16172);
xnor U21610 (N_21610,N_14002,N_16063);
nand U21611 (N_21611,N_17425,N_13545);
nor U21612 (N_21612,N_14171,N_17448);
xnor U21613 (N_21613,N_15929,N_16864);
or U21614 (N_21614,N_18309,N_14866);
nor U21615 (N_21615,N_16634,N_13934);
nand U21616 (N_21616,N_17035,N_14406);
nor U21617 (N_21617,N_16877,N_16192);
nand U21618 (N_21618,N_16208,N_15938);
nor U21619 (N_21619,N_16915,N_15056);
nand U21620 (N_21620,N_13143,N_15933);
and U21621 (N_21621,N_16936,N_15408);
and U21622 (N_21622,N_15818,N_13364);
or U21623 (N_21623,N_15921,N_14995);
or U21624 (N_21624,N_14466,N_15817);
nor U21625 (N_21625,N_16866,N_18145);
xnor U21626 (N_21626,N_16954,N_15716);
nand U21627 (N_21627,N_16559,N_17859);
nor U21628 (N_21628,N_14730,N_16226);
xor U21629 (N_21629,N_18269,N_17108);
nor U21630 (N_21630,N_14434,N_15742);
or U21631 (N_21631,N_15601,N_16727);
or U21632 (N_21632,N_15275,N_16360);
nor U21633 (N_21633,N_13710,N_16179);
and U21634 (N_21634,N_12783,N_12715);
or U21635 (N_21635,N_15985,N_13441);
or U21636 (N_21636,N_12655,N_18207);
and U21637 (N_21637,N_12855,N_17308);
or U21638 (N_21638,N_16416,N_16751);
nand U21639 (N_21639,N_14637,N_16819);
and U21640 (N_21640,N_17953,N_12733);
nor U21641 (N_21641,N_17743,N_13444);
or U21642 (N_21642,N_15363,N_17592);
and U21643 (N_21643,N_14219,N_14329);
nor U21644 (N_21644,N_18347,N_12723);
or U21645 (N_21645,N_12526,N_15910);
nor U21646 (N_21646,N_16686,N_15680);
or U21647 (N_21647,N_16784,N_14518);
xnor U21648 (N_21648,N_12843,N_16674);
xnor U21649 (N_21649,N_18290,N_14243);
or U21650 (N_21650,N_18530,N_18250);
and U21651 (N_21651,N_12896,N_15914);
nand U21652 (N_21652,N_18002,N_18656);
xnor U21653 (N_21653,N_15184,N_13025);
and U21654 (N_21654,N_17347,N_13891);
nor U21655 (N_21655,N_15569,N_14025);
or U21656 (N_21656,N_16064,N_16808);
nand U21657 (N_21657,N_18689,N_16702);
nor U21658 (N_21658,N_13717,N_14089);
nand U21659 (N_21659,N_15005,N_17693);
and U21660 (N_21660,N_17645,N_17675);
xnor U21661 (N_21661,N_12643,N_16839);
or U21662 (N_21662,N_13004,N_16065);
nand U21663 (N_21663,N_13138,N_13160);
nand U21664 (N_21664,N_14058,N_16862);
xnor U21665 (N_21665,N_13219,N_13678);
or U21666 (N_21666,N_14620,N_17614);
nor U21667 (N_21667,N_12883,N_15796);
and U21668 (N_21668,N_15769,N_15330);
nand U21669 (N_21669,N_17864,N_15580);
nor U21670 (N_21670,N_14399,N_12823);
or U21671 (N_21671,N_12524,N_14891);
nor U21672 (N_21672,N_14557,N_17033);
nor U21673 (N_21673,N_18554,N_16623);
or U21674 (N_21674,N_18557,N_15510);
nor U21675 (N_21675,N_13034,N_16451);
nand U21676 (N_21676,N_13581,N_15978);
and U21677 (N_21677,N_14048,N_15034);
or U21678 (N_21678,N_12790,N_18144);
and U21679 (N_21679,N_18729,N_15971);
or U21680 (N_21680,N_14131,N_14208);
and U21681 (N_21681,N_16130,N_17694);
nand U21682 (N_21682,N_17970,N_18091);
or U21683 (N_21683,N_15153,N_13685);
xnor U21684 (N_21684,N_17510,N_18188);
or U21685 (N_21685,N_17229,N_13944);
and U21686 (N_21686,N_14298,N_17940);
nand U21687 (N_21687,N_14688,N_17148);
xnor U21688 (N_21688,N_13731,N_16417);
nand U21689 (N_21689,N_13378,N_14823);
nor U21690 (N_21690,N_18080,N_15426);
nand U21691 (N_21691,N_14895,N_15790);
nor U21692 (N_21692,N_12690,N_16305);
or U21693 (N_21693,N_18178,N_17619);
or U21694 (N_21694,N_18098,N_14410);
or U21695 (N_21695,N_13203,N_15814);
nand U21696 (N_21696,N_15022,N_13523);
nor U21697 (N_21697,N_13020,N_13427);
xnor U21698 (N_21698,N_14368,N_15916);
nand U21699 (N_21699,N_15906,N_17211);
nand U21700 (N_21700,N_13436,N_14669);
or U21701 (N_21701,N_16765,N_18677);
nor U21702 (N_21702,N_13632,N_18276);
nand U21703 (N_21703,N_17376,N_17289);
nor U21704 (N_21704,N_16343,N_15913);
and U21705 (N_21705,N_18704,N_18081);
or U21706 (N_21706,N_13637,N_16649);
or U21707 (N_21707,N_17569,N_13895);
nand U21708 (N_21708,N_16345,N_17832);
nor U21709 (N_21709,N_14642,N_18259);
nand U21710 (N_21710,N_14796,N_14309);
nand U21711 (N_21711,N_18528,N_17784);
or U21712 (N_21712,N_18079,N_18735);
nand U21713 (N_21713,N_16446,N_15509);
xnor U21714 (N_21714,N_14160,N_16785);
nand U21715 (N_21715,N_17003,N_17901);
xor U21716 (N_21716,N_18638,N_15325);
and U21717 (N_21717,N_17361,N_16801);
nor U21718 (N_21718,N_12617,N_13264);
or U21719 (N_21719,N_15605,N_14052);
or U21720 (N_21720,N_15328,N_15401);
nand U21721 (N_21721,N_16497,N_12812);
nand U21722 (N_21722,N_13332,N_14749);
or U21723 (N_21723,N_18500,N_17247);
nand U21724 (N_21724,N_17722,N_18619);
and U21725 (N_21725,N_12550,N_16865);
xor U21726 (N_21726,N_17248,N_17325);
xnor U21727 (N_21727,N_15610,N_16881);
and U21728 (N_21728,N_17975,N_16858);
or U21729 (N_21729,N_17198,N_12888);
and U21730 (N_21730,N_14883,N_17408);
and U21731 (N_21731,N_14606,N_16805);
and U21732 (N_21732,N_15116,N_18521);
and U21733 (N_21733,N_15096,N_16357);
or U21734 (N_21734,N_16284,N_17533);
xnor U21735 (N_21735,N_17225,N_17941);
nand U21736 (N_21736,N_13726,N_15526);
nor U21737 (N_21737,N_14217,N_15036);
nor U21738 (N_21738,N_17597,N_16861);
nor U21739 (N_21739,N_16152,N_13828);
nand U21740 (N_21740,N_18176,N_18075);
and U21741 (N_21741,N_13985,N_13039);
and U21742 (N_21742,N_17049,N_16816);
or U21743 (N_21743,N_14500,N_12976);
xnor U21744 (N_21744,N_14561,N_13773);
xnor U21745 (N_21745,N_15733,N_16287);
and U21746 (N_21746,N_18333,N_16892);
nor U21747 (N_21747,N_17823,N_16716);
or U21748 (N_21748,N_17717,N_17400);
nor U21749 (N_21749,N_16818,N_15499);
and U21750 (N_21750,N_15864,N_13227);
or U21751 (N_21751,N_16186,N_13277);
and U21752 (N_21752,N_17426,N_13815);
nor U21753 (N_21753,N_17446,N_12608);
and U21754 (N_21754,N_15690,N_18312);
nand U21755 (N_21755,N_18582,N_18643);
xnor U21756 (N_21756,N_14690,N_16795);
nand U21757 (N_21757,N_15902,N_14754);
and U21758 (N_21758,N_14098,N_15868);
nor U21759 (N_21759,N_13690,N_18533);
and U21760 (N_21760,N_15087,N_18087);
or U21761 (N_21761,N_12589,N_18291);
nand U21762 (N_21762,N_12561,N_17707);
xnor U21763 (N_21763,N_13032,N_15757);
or U21764 (N_21764,N_14438,N_17883);
nand U21765 (N_21765,N_13358,N_13776);
or U21766 (N_21766,N_18653,N_15135);
nor U21767 (N_21767,N_14395,N_15560);
xnor U21768 (N_21768,N_13519,N_17066);
or U21769 (N_21769,N_15351,N_15781);
xor U21770 (N_21770,N_16542,N_16966);
nor U21771 (N_21771,N_18732,N_16035);
or U21772 (N_21772,N_17471,N_18059);
nor U21773 (N_21773,N_14605,N_18739);
xor U21774 (N_21774,N_12644,N_16123);
nand U21775 (N_21775,N_16185,N_12588);
or U21776 (N_21776,N_18303,N_18745);
or U21777 (N_21777,N_17077,N_17835);
nand U21778 (N_21778,N_15874,N_12599);
and U21779 (N_21779,N_12693,N_13952);
xor U21780 (N_21780,N_15667,N_18705);
nand U21781 (N_21781,N_12856,N_17130);
nor U21782 (N_21782,N_12709,N_14022);
xor U21783 (N_21783,N_17999,N_18236);
xor U21784 (N_21784,N_16810,N_15849);
nor U21785 (N_21785,N_16133,N_17947);
nand U21786 (N_21786,N_12963,N_17390);
nor U21787 (N_21787,N_12985,N_15240);
nand U21788 (N_21788,N_17500,N_17839);
and U21789 (N_21789,N_18281,N_16273);
and U21790 (N_21790,N_13612,N_18609);
or U21791 (N_21791,N_17877,N_18296);
nand U21792 (N_21792,N_17267,N_16552);
and U21793 (N_21793,N_16863,N_12613);
and U21794 (N_21794,N_18017,N_14352);
nand U21795 (N_21795,N_18551,N_15643);
xnor U21796 (N_21796,N_14876,N_17507);
or U21797 (N_21797,N_16589,N_14216);
nor U21798 (N_21798,N_13001,N_14838);
xor U21799 (N_21799,N_16655,N_16912);
nand U21800 (N_21800,N_13972,N_12832);
or U21801 (N_21801,N_14262,N_16857);
or U21802 (N_21802,N_13595,N_13338);
or U21803 (N_21803,N_15975,N_14202);
nand U21804 (N_21804,N_14263,N_12866);
nand U21805 (N_21805,N_16266,N_18090);
nand U21806 (N_21806,N_13707,N_13730);
or U21807 (N_21807,N_13716,N_14452);
nor U21808 (N_21808,N_17406,N_17814);
and U21809 (N_21809,N_18724,N_12975);
or U21810 (N_21810,N_15268,N_15500);
nor U21811 (N_21811,N_16971,N_18436);
nand U21812 (N_21812,N_13183,N_18400);
or U21813 (N_21813,N_14696,N_17070);
and U21814 (N_21814,N_16717,N_17388);
xnor U21815 (N_21815,N_15155,N_18194);
nand U21816 (N_21816,N_13848,N_16897);
and U21817 (N_21817,N_14073,N_12604);
or U21818 (N_21818,N_13387,N_17660);
nand U21819 (N_21819,N_13291,N_13180);
xor U21820 (N_21820,N_14856,N_18212);
and U21821 (N_21821,N_16102,N_18283);
and U21822 (N_21822,N_16447,N_17322);
or U21823 (N_21823,N_18720,N_15599);
or U21824 (N_21824,N_14521,N_16995);
or U21825 (N_21825,N_16575,N_17453);
nor U21826 (N_21826,N_13867,N_16214);
nand U21827 (N_21827,N_13721,N_13156);
xnor U21828 (N_21828,N_14750,N_18335);
nand U21829 (N_21829,N_13869,N_18374);
or U21830 (N_21830,N_12879,N_17464);
nor U21831 (N_21831,N_17180,N_16427);
nor U21832 (N_21832,N_13628,N_18700);
nand U21833 (N_21833,N_12671,N_18047);
nor U21834 (N_21834,N_17921,N_16840);
or U21835 (N_21835,N_14573,N_12543);
and U21836 (N_21836,N_15973,N_17026);
xor U21837 (N_21837,N_17363,N_13718);
xnor U21838 (N_21838,N_13214,N_16573);
or U21839 (N_21839,N_14778,N_16145);
nor U21840 (N_21840,N_14513,N_13673);
nand U21841 (N_21841,N_14092,N_12691);
or U21842 (N_21842,N_17268,N_17356);
or U21843 (N_21843,N_13817,N_16988);
or U21844 (N_21844,N_16485,N_13476);
or U21845 (N_21845,N_18302,N_13310);
nand U21846 (N_21846,N_18393,N_14918);
or U21847 (N_21847,N_17650,N_17780);
nor U21848 (N_21848,N_16665,N_14338);
or U21849 (N_21849,N_13618,N_16809);
nand U21850 (N_21850,N_15993,N_15501);
nor U21851 (N_21851,N_15972,N_15763);
or U21852 (N_21852,N_15017,N_17754);
xnor U21853 (N_21853,N_12727,N_17910);
xnor U21854 (N_21854,N_15718,N_17485);
nand U21855 (N_21855,N_13198,N_15262);
or U21856 (N_21856,N_13851,N_13500);
and U21857 (N_21857,N_14204,N_13857);
and U21858 (N_21858,N_15255,N_12673);
or U21859 (N_21859,N_13803,N_15257);
nor U21860 (N_21860,N_12731,N_15673);
xor U21861 (N_21861,N_14494,N_17039);
xor U21862 (N_21862,N_14623,N_16375);
nand U21863 (N_21863,N_16165,N_15410);
nor U21864 (N_21864,N_13041,N_17192);
and U21865 (N_21865,N_13604,N_14420);
xnor U21866 (N_21866,N_14250,N_14703);
nand U21867 (N_21867,N_16331,N_16137);
and U21868 (N_21868,N_12946,N_12632);
nor U21869 (N_21869,N_12776,N_13941);
nand U21870 (N_21870,N_17217,N_15492);
nor U21871 (N_21871,N_15574,N_13394);
xor U21872 (N_21872,N_13652,N_18160);
or U21873 (N_21873,N_15304,N_17758);
or U21874 (N_21874,N_13902,N_13309);
nor U21875 (N_21875,N_17512,N_17696);
nand U21876 (N_21876,N_16225,N_13971);
nand U21877 (N_21877,N_17124,N_13279);
and U21878 (N_21878,N_15145,N_13783);
or U21879 (N_21879,N_18014,N_12752);
and U21880 (N_21880,N_17219,N_13850);
nand U21881 (N_21881,N_13888,N_13800);
nor U21882 (N_21882,N_14304,N_17609);
nand U21883 (N_21883,N_12876,N_18399);
or U21884 (N_21884,N_14827,N_13180);
nor U21885 (N_21885,N_18376,N_17589);
nor U21886 (N_21886,N_16326,N_15932);
xnor U21887 (N_21887,N_18564,N_16312);
or U21888 (N_21888,N_17544,N_17484);
and U21889 (N_21889,N_14296,N_15321);
xor U21890 (N_21890,N_14439,N_17009);
nand U21891 (N_21891,N_16917,N_15403);
or U21892 (N_21892,N_13261,N_16291);
xor U21893 (N_21893,N_14624,N_16454);
and U21894 (N_21894,N_13718,N_17555);
or U21895 (N_21895,N_13313,N_16092);
or U21896 (N_21896,N_16310,N_17091);
nor U21897 (N_21897,N_15481,N_14162);
xnor U21898 (N_21898,N_13615,N_14721);
xor U21899 (N_21899,N_14173,N_14216);
nand U21900 (N_21900,N_16170,N_12852);
nand U21901 (N_21901,N_13571,N_16812);
xor U21902 (N_21902,N_16740,N_17933);
xnor U21903 (N_21903,N_15883,N_16975);
nor U21904 (N_21904,N_17714,N_17555);
nor U21905 (N_21905,N_14337,N_14825);
or U21906 (N_21906,N_12647,N_13822);
and U21907 (N_21907,N_17430,N_17157);
nor U21908 (N_21908,N_16695,N_13099);
and U21909 (N_21909,N_14261,N_13943);
or U21910 (N_21910,N_12965,N_13373);
nor U21911 (N_21911,N_16419,N_14679);
and U21912 (N_21912,N_18689,N_15943);
and U21913 (N_21913,N_13551,N_15549);
nand U21914 (N_21914,N_15224,N_15562);
and U21915 (N_21915,N_17813,N_15565);
nor U21916 (N_21916,N_17641,N_16835);
and U21917 (N_21917,N_17354,N_14542);
or U21918 (N_21918,N_13750,N_13567);
nor U21919 (N_21919,N_14434,N_18408);
and U21920 (N_21920,N_13941,N_15210);
and U21921 (N_21921,N_16871,N_12521);
nand U21922 (N_21922,N_15234,N_17970);
or U21923 (N_21923,N_15266,N_13306);
xor U21924 (N_21924,N_13159,N_14374);
or U21925 (N_21925,N_16932,N_13088);
and U21926 (N_21926,N_17000,N_12911);
and U21927 (N_21927,N_18539,N_12580);
xnor U21928 (N_21928,N_16167,N_16274);
nand U21929 (N_21929,N_15166,N_18538);
xor U21930 (N_21930,N_16992,N_12797);
xnor U21931 (N_21931,N_17180,N_18243);
nor U21932 (N_21932,N_15792,N_17539);
nor U21933 (N_21933,N_13154,N_16438);
or U21934 (N_21934,N_12943,N_17891);
xor U21935 (N_21935,N_14146,N_16076);
nor U21936 (N_21936,N_17198,N_17071);
nand U21937 (N_21937,N_15669,N_12670);
nor U21938 (N_21938,N_15375,N_17179);
nor U21939 (N_21939,N_17840,N_15792);
xnor U21940 (N_21940,N_15635,N_12849);
or U21941 (N_21941,N_13659,N_12651);
and U21942 (N_21942,N_14710,N_12801);
or U21943 (N_21943,N_15967,N_15073);
nand U21944 (N_21944,N_15077,N_13223);
xor U21945 (N_21945,N_15831,N_18535);
or U21946 (N_21946,N_17495,N_13990);
nor U21947 (N_21947,N_18313,N_15489);
or U21948 (N_21948,N_14708,N_14377);
and U21949 (N_21949,N_17014,N_14182);
and U21950 (N_21950,N_14880,N_18083);
or U21951 (N_21951,N_12721,N_14714);
nor U21952 (N_21952,N_13287,N_16419);
nor U21953 (N_21953,N_17925,N_16463);
nor U21954 (N_21954,N_16236,N_15261);
and U21955 (N_21955,N_12566,N_12848);
and U21956 (N_21956,N_14580,N_18522);
and U21957 (N_21957,N_15841,N_16225);
nor U21958 (N_21958,N_18473,N_12928);
nand U21959 (N_21959,N_12805,N_17899);
xor U21960 (N_21960,N_13809,N_16962);
nor U21961 (N_21961,N_15179,N_15467);
nand U21962 (N_21962,N_13314,N_17631);
or U21963 (N_21963,N_16228,N_17060);
or U21964 (N_21964,N_18486,N_14608);
xnor U21965 (N_21965,N_17519,N_17620);
xnor U21966 (N_21966,N_16954,N_15959);
or U21967 (N_21967,N_16136,N_15556);
and U21968 (N_21968,N_17905,N_17076);
and U21969 (N_21969,N_15352,N_17991);
nor U21970 (N_21970,N_13762,N_16567);
or U21971 (N_21971,N_17006,N_16388);
nor U21972 (N_21972,N_16893,N_18298);
xnor U21973 (N_21973,N_13128,N_12819);
or U21974 (N_21974,N_18053,N_18170);
or U21975 (N_21975,N_13131,N_17516);
and U21976 (N_21976,N_18413,N_17900);
and U21977 (N_21977,N_17621,N_17961);
nor U21978 (N_21978,N_15880,N_13241);
nor U21979 (N_21979,N_16983,N_18650);
and U21980 (N_21980,N_14915,N_13400);
and U21981 (N_21981,N_17319,N_15494);
nand U21982 (N_21982,N_18283,N_17526);
or U21983 (N_21983,N_13466,N_18356);
nand U21984 (N_21984,N_15451,N_17881);
and U21985 (N_21985,N_16324,N_17868);
xnor U21986 (N_21986,N_15245,N_18560);
xor U21987 (N_21987,N_12663,N_14813);
nand U21988 (N_21988,N_13453,N_16152);
and U21989 (N_21989,N_13507,N_18322);
xnor U21990 (N_21990,N_14416,N_16377);
nand U21991 (N_21991,N_16785,N_15159);
or U21992 (N_21992,N_17032,N_16195);
and U21993 (N_21993,N_13872,N_17689);
nand U21994 (N_21994,N_15536,N_14535);
nand U21995 (N_21995,N_16621,N_15776);
nor U21996 (N_21996,N_12518,N_17528);
nor U21997 (N_21997,N_18231,N_15374);
and U21998 (N_21998,N_13644,N_13328);
xor U21999 (N_21999,N_12833,N_16618);
and U22000 (N_22000,N_17451,N_16262);
or U22001 (N_22001,N_17545,N_14718);
or U22002 (N_22002,N_17655,N_15751);
xnor U22003 (N_22003,N_14719,N_14506);
or U22004 (N_22004,N_12846,N_17673);
nor U22005 (N_22005,N_13498,N_13641);
nor U22006 (N_22006,N_18681,N_17835);
xnor U22007 (N_22007,N_14750,N_14327);
and U22008 (N_22008,N_12639,N_16699);
nor U22009 (N_22009,N_13375,N_17392);
or U22010 (N_22010,N_12683,N_16791);
or U22011 (N_22011,N_13509,N_18346);
xnor U22012 (N_22012,N_16752,N_16960);
or U22013 (N_22013,N_14860,N_16416);
and U22014 (N_22014,N_18282,N_13731);
nand U22015 (N_22015,N_15598,N_14079);
nor U22016 (N_22016,N_18541,N_17569);
xnor U22017 (N_22017,N_13445,N_16441);
or U22018 (N_22018,N_14951,N_15757);
nand U22019 (N_22019,N_15472,N_13656);
xnor U22020 (N_22020,N_17755,N_12777);
nand U22021 (N_22021,N_13231,N_12604);
nand U22022 (N_22022,N_15354,N_15330);
or U22023 (N_22023,N_14208,N_16104);
nor U22024 (N_22024,N_18211,N_14361);
nand U22025 (N_22025,N_15191,N_15212);
nor U22026 (N_22026,N_16605,N_13534);
nor U22027 (N_22027,N_16117,N_14035);
nand U22028 (N_22028,N_16446,N_14858);
or U22029 (N_22029,N_12759,N_17202);
xnor U22030 (N_22030,N_15729,N_15404);
nand U22031 (N_22031,N_13421,N_13202);
nand U22032 (N_22032,N_18542,N_13151);
or U22033 (N_22033,N_16332,N_14503);
nor U22034 (N_22034,N_12738,N_14224);
or U22035 (N_22035,N_14421,N_13854);
or U22036 (N_22036,N_17795,N_15781);
xnor U22037 (N_22037,N_14142,N_13363);
or U22038 (N_22038,N_12917,N_13266);
xor U22039 (N_22039,N_17997,N_16841);
or U22040 (N_22040,N_14049,N_17810);
and U22041 (N_22041,N_14372,N_16127);
or U22042 (N_22042,N_16829,N_13464);
and U22043 (N_22043,N_16369,N_18204);
nand U22044 (N_22044,N_12739,N_14620);
and U22045 (N_22045,N_16110,N_13030);
and U22046 (N_22046,N_14745,N_16849);
xnor U22047 (N_22047,N_17498,N_13249);
nand U22048 (N_22048,N_18369,N_16618);
nor U22049 (N_22049,N_15173,N_16472);
or U22050 (N_22050,N_14187,N_16054);
nor U22051 (N_22051,N_18257,N_14939);
or U22052 (N_22052,N_12632,N_16653);
and U22053 (N_22053,N_17012,N_18386);
nor U22054 (N_22054,N_12590,N_13914);
nor U22055 (N_22055,N_13148,N_18184);
nand U22056 (N_22056,N_13946,N_16887);
and U22057 (N_22057,N_17847,N_12870);
nor U22058 (N_22058,N_17555,N_16148);
and U22059 (N_22059,N_14107,N_17148);
xnor U22060 (N_22060,N_18365,N_16607);
nor U22061 (N_22061,N_15449,N_12854);
and U22062 (N_22062,N_18627,N_15613);
xnor U22063 (N_22063,N_15411,N_15094);
nand U22064 (N_22064,N_17039,N_15608);
nor U22065 (N_22065,N_13384,N_15512);
nor U22066 (N_22066,N_13322,N_13107);
xnor U22067 (N_22067,N_16746,N_15580);
nor U22068 (N_22068,N_15572,N_14341);
and U22069 (N_22069,N_13819,N_16067);
and U22070 (N_22070,N_13991,N_15115);
and U22071 (N_22071,N_18436,N_17100);
or U22072 (N_22072,N_16483,N_17252);
nor U22073 (N_22073,N_14946,N_13264);
and U22074 (N_22074,N_18670,N_13832);
nand U22075 (N_22075,N_13893,N_15099);
nand U22076 (N_22076,N_15908,N_14941);
or U22077 (N_22077,N_13987,N_16924);
and U22078 (N_22078,N_14371,N_12582);
xor U22079 (N_22079,N_15805,N_13915);
and U22080 (N_22080,N_17732,N_13648);
xor U22081 (N_22081,N_15396,N_16697);
nand U22082 (N_22082,N_17231,N_17607);
or U22083 (N_22083,N_12776,N_18501);
or U22084 (N_22084,N_13030,N_14749);
nand U22085 (N_22085,N_17391,N_16533);
nor U22086 (N_22086,N_17248,N_17778);
or U22087 (N_22087,N_14771,N_13498);
xor U22088 (N_22088,N_14428,N_14036);
nand U22089 (N_22089,N_17346,N_14659);
nor U22090 (N_22090,N_16447,N_14544);
and U22091 (N_22091,N_15693,N_12845);
or U22092 (N_22092,N_15929,N_14481);
nor U22093 (N_22093,N_15604,N_17264);
nand U22094 (N_22094,N_16988,N_13654);
and U22095 (N_22095,N_16149,N_16329);
nand U22096 (N_22096,N_18536,N_17047);
nand U22097 (N_22097,N_14476,N_17116);
nand U22098 (N_22098,N_15277,N_16402);
or U22099 (N_22099,N_15176,N_18272);
nor U22100 (N_22100,N_13114,N_17771);
or U22101 (N_22101,N_18561,N_18551);
nand U22102 (N_22102,N_14230,N_14411);
xnor U22103 (N_22103,N_16747,N_18149);
nor U22104 (N_22104,N_16359,N_17962);
or U22105 (N_22105,N_18076,N_17221);
xnor U22106 (N_22106,N_15867,N_18262);
xor U22107 (N_22107,N_15836,N_14205);
and U22108 (N_22108,N_13980,N_15539);
or U22109 (N_22109,N_13984,N_17822);
nor U22110 (N_22110,N_16138,N_17004);
nand U22111 (N_22111,N_17002,N_14213);
or U22112 (N_22112,N_14846,N_18471);
xnor U22113 (N_22113,N_13229,N_17273);
and U22114 (N_22114,N_14740,N_16271);
nand U22115 (N_22115,N_18475,N_13116);
or U22116 (N_22116,N_16697,N_13573);
nor U22117 (N_22117,N_16540,N_14495);
and U22118 (N_22118,N_13363,N_15404);
and U22119 (N_22119,N_12866,N_15816);
nand U22120 (N_22120,N_18063,N_18051);
nand U22121 (N_22121,N_13335,N_13856);
and U22122 (N_22122,N_12961,N_17150);
nor U22123 (N_22123,N_12515,N_12627);
xnor U22124 (N_22124,N_18149,N_17120);
xnor U22125 (N_22125,N_17641,N_12502);
nand U22126 (N_22126,N_15424,N_17620);
nor U22127 (N_22127,N_17826,N_14548);
or U22128 (N_22128,N_16599,N_15293);
nor U22129 (N_22129,N_18746,N_16909);
nand U22130 (N_22130,N_16498,N_14541);
xnor U22131 (N_22131,N_18087,N_15771);
xnor U22132 (N_22132,N_17865,N_15105);
and U22133 (N_22133,N_12761,N_14740);
nor U22134 (N_22134,N_13871,N_14380);
xnor U22135 (N_22135,N_12671,N_13097);
and U22136 (N_22136,N_17606,N_12964);
or U22137 (N_22137,N_16257,N_13619);
and U22138 (N_22138,N_13597,N_14028);
xor U22139 (N_22139,N_13858,N_15960);
and U22140 (N_22140,N_14948,N_15993);
nand U22141 (N_22141,N_17115,N_16246);
xnor U22142 (N_22142,N_12557,N_14515);
xor U22143 (N_22143,N_18337,N_12561);
or U22144 (N_22144,N_15451,N_18080);
xor U22145 (N_22145,N_16862,N_13903);
or U22146 (N_22146,N_14813,N_13861);
nor U22147 (N_22147,N_17716,N_16369);
nor U22148 (N_22148,N_13713,N_15208);
and U22149 (N_22149,N_16879,N_13205);
and U22150 (N_22150,N_18311,N_16011);
or U22151 (N_22151,N_17503,N_13305);
nor U22152 (N_22152,N_18678,N_13418);
and U22153 (N_22153,N_13050,N_13782);
nor U22154 (N_22154,N_15992,N_15279);
nand U22155 (N_22155,N_17042,N_14037);
xnor U22156 (N_22156,N_15289,N_17693);
or U22157 (N_22157,N_15854,N_18084);
or U22158 (N_22158,N_17605,N_13585);
and U22159 (N_22159,N_18132,N_14423);
nor U22160 (N_22160,N_13115,N_17497);
or U22161 (N_22161,N_18263,N_14336);
nand U22162 (N_22162,N_16950,N_15208);
nor U22163 (N_22163,N_16867,N_12533);
xor U22164 (N_22164,N_16329,N_13576);
nand U22165 (N_22165,N_16852,N_18015);
or U22166 (N_22166,N_14032,N_18080);
xnor U22167 (N_22167,N_18142,N_18133);
nor U22168 (N_22168,N_17796,N_15842);
xor U22169 (N_22169,N_18309,N_17745);
xnor U22170 (N_22170,N_15528,N_13201);
xnor U22171 (N_22171,N_15062,N_15055);
nor U22172 (N_22172,N_16621,N_18198);
or U22173 (N_22173,N_13147,N_14650);
xnor U22174 (N_22174,N_17285,N_16088);
nand U22175 (N_22175,N_15444,N_12531);
nand U22176 (N_22176,N_16058,N_16212);
xor U22177 (N_22177,N_14898,N_18473);
xor U22178 (N_22178,N_17743,N_16520);
or U22179 (N_22179,N_15457,N_17169);
or U22180 (N_22180,N_12863,N_18356);
and U22181 (N_22181,N_17819,N_17997);
nand U22182 (N_22182,N_13974,N_14386);
or U22183 (N_22183,N_16410,N_12656);
or U22184 (N_22184,N_15968,N_16630);
and U22185 (N_22185,N_12594,N_17329);
xor U22186 (N_22186,N_12574,N_12872);
xor U22187 (N_22187,N_16338,N_16828);
and U22188 (N_22188,N_13588,N_14504);
nand U22189 (N_22189,N_18058,N_13451);
nand U22190 (N_22190,N_18625,N_17033);
nor U22191 (N_22191,N_17490,N_16691);
nand U22192 (N_22192,N_14978,N_17659);
nand U22193 (N_22193,N_13396,N_17004);
nor U22194 (N_22194,N_12518,N_17192);
and U22195 (N_22195,N_12540,N_17865);
nor U22196 (N_22196,N_14716,N_16169);
nor U22197 (N_22197,N_18543,N_16540);
xnor U22198 (N_22198,N_14417,N_17994);
nand U22199 (N_22199,N_15501,N_12868);
nor U22200 (N_22200,N_13237,N_12913);
and U22201 (N_22201,N_17295,N_13230);
xor U22202 (N_22202,N_13396,N_14119);
nand U22203 (N_22203,N_18502,N_16220);
or U22204 (N_22204,N_17199,N_17642);
xnor U22205 (N_22205,N_13684,N_12529);
or U22206 (N_22206,N_18399,N_16883);
and U22207 (N_22207,N_16015,N_16291);
or U22208 (N_22208,N_15388,N_15108);
nor U22209 (N_22209,N_16541,N_16105);
xor U22210 (N_22210,N_13358,N_17440);
nor U22211 (N_22211,N_13247,N_13527);
xnor U22212 (N_22212,N_14905,N_13301);
xnor U22213 (N_22213,N_13188,N_18618);
nor U22214 (N_22214,N_16223,N_13138);
nand U22215 (N_22215,N_18334,N_16324);
and U22216 (N_22216,N_14044,N_16610);
nand U22217 (N_22217,N_13894,N_14687);
nand U22218 (N_22218,N_13959,N_14027);
nand U22219 (N_22219,N_12993,N_13764);
xor U22220 (N_22220,N_15672,N_17179);
xnor U22221 (N_22221,N_13631,N_15405);
and U22222 (N_22222,N_15973,N_17871);
and U22223 (N_22223,N_16106,N_18179);
nor U22224 (N_22224,N_16602,N_16177);
and U22225 (N_22225,N_17192,N_17100);
xnor U22226 (N_22226,N_13084,N_17825);
and U22227 (N_22227,N_15433,N_13463);
nand U22228 (N_22228,N_17007,N_14586);
nor U22229 (N_22229,N_12895,N_16057);
nand U22230 (N_22230,N_17256,N_15305);
and U22231 (N_22231,N_13343,N_17686);
or U22232 (N_22232,N_16508,N_14409);
nor U22233 (N_22233,N_14928,N_17423);
or U22234 (N_22234,N_14203,N_14730);
or U22235 (N_22235,N_17426,N_18644);
nand U22236 (N_22236,N_13054,N_14039);
nand U22237 (N_22237,N_14186,N_12991);
and U22238 (N_22238,N_14190,N_14074);
nand U22239 (N_22239,N_13867,N_13749);
or U22240 (N_22240,N_12508,N_15446);
xor U22241 (N_22241,N_12842,N_13308);
and U22242 (N_22242,N_14154,N_18071);
nand U22243 (N_22243,N_13072,N_17731);
nand U22244 (N_22244,N_14631,N_15904);
nand U22245 (N_22245,N_17904,N_15512);
xor U22246 (N_22246,N_12764,N_16153);
xnor U22247 (N_22247,N_12926,N_15338);
and U22248 (N_22248,N_17406,N_13706);
and U22249 (N_22249,N_13800,N_14641);
or U22250 (N_22250,N_14801,N_17207);
and U22251 (N_22251,N_17622,N_12607);
nor U22252 (N_22252,N_15151,N_18040);
nor U22253 (N_22253,N_14145,N_16062);
and U22254 (N_22254,N_18706,N_17351);
xnor U22255 (N_22255,N_12939,N_13522);
nor U22256 (N_22256,N_15106,N_18485);
nand U22257 (N_22257,N_13636,N_14758);
or U22258 (N_22258,N_15172,N_12860);
nand U22259 (N_22259,N_14783,N_13632);
or U22260 (N_22260,N_15650,N_13520);
and U22261 (N_22261,N_13953,N_13299);
and U22262 (N_22262,N_13812,N_17934);
xor U22263 (N_22263,N_13212,N_14274);
or U22264 (N_22264,N_17070,N_15484);
nand U22265 (N_22265,N_13732,N_15860);
nor U22266 (N_22266,N_15983,N_15378);
and U22267 (N_22267,N_16889,N_13947);
xnor U22268 (N_22268,N_18488,N_15028);
and U22269 (N_22269,N_12912,N_16411);
nand U22270 (N_22270,N_18441,N_17257);
xnor U22271 (N_22271,N_14194,N_18478);
or U22272 (N_22272,N_15285,N_14050);
nor U22273 (N_22273,N_12967,N_14620);
nand U22274 (N_22274,N_15787,N_12886);
or U22275 (N_22275,N_18701,N_12763);
or U22276 (N_22276,N_13813,N_14176);
nor U22277 (N_22277,N_17744,N_15722);
nor U22278 (N_22278,N_17609,N_13252);
or U22279 (N_22279,N_13827,N_16436);
nand U22280 (N_22280,N_16499,N_14041);
nor U22281 (N_22281,N_16685,N_17246);
nand U22282 (N_22282,N_18663,N_17281);
xnor U22283 (N_22283,N_14322,N_13790);
xor U22284 (N_22284,N_17085,N_18100);
or U22285 (N_22285,N_15537,N_17404);
nor U22286 (N_22286,N_16661,N_17148);
and U22287 (N_22287,N_17501,N_15607);
and U22288 (N_22288,N_16814,N_17052);
nand U22289 (N_22289,N_15789,N_12826);
xor U22290 (N_22290,N_14253,N_15784);
nand U22291 (N_22291,N_17784,N_12953);
nand U22292 (N_22292,N_15662,N_18473);
xnor U22293 (N_22293,N_16425,N_16006);
or U22294 (N_22294,N_13260,N_17894);
nand U22295 (N_22295,N_14728,N_13439);
nor U22296 (N_22296,N_16733,N_15138);
nand U22297 (N_22297,N_13231,N_14487);
nor U22298 (N_22298,N_15422,N_17679);
or U22299 (N_22299,N_13670,N_15708);
nand U22300 (N_22300,N_15964,N_16819);
nand U22301 (N_22301,N_16632,N_16368);
or U22302 (N_22302,N_15285,N_17173);
nor U22303 (N_22303,N_14970,N_14493);
or U22304 (N_22304,N_16947,N_12864);
nand U22305 (N_22305,N_14628,N_12699);
nand U22306 (N_22306,N_15998,N_13579);
and U22307 (N_22307,N_15682,N_17163);
and U22308 (N_22308,N_16345,N_13302);
nor U22309 (N_22309,N_16105,N_15286);
xnor U22310 (N_22310,N_13102,N_14895);
xnor U22311 (N_22311,N_17897,N_18160);
or U22312 (N_22312,N_12769,N_17198);
xnor U22313 (N_22313,N_15566,N_15447);
or U22314 (N_22314,N_15343,N_14109);
and U22315 (N_22315,N_13829,N_14157);
nand U22316 (N_22316,N_16484,N_14712);
and U22317 (N_22317,N_17858,N_15834);
xnor U22318 (N_22318,N_12549,N_15548);
and U22319 (N_22319,N_14999,N_13194);
nor U22320 (N_22320,N_17717,N_12630);
nor U22321 (N_22321,N_17595,N_12635);
nand U22322 (N_22322,N_14528,N_17935);
nor U22323 (N_22323,N_13688,N_17308);
xor U22324 (N_22324,N_13718,N_14903);
nor U22325 (N_22325,N_16160,N_18591);
xnor U22326 (N_22326,N_14057,N_15376);
xor U22327 (N_22327,N_17439,N_13839);
or U22328 (N_22328,N_14005,N_18148);
or U22329 (N_22329,N_13084,N_17332);
and U22330 (N_22330,N_17043,N_17216);
xor U22331 (N_22331,N_13236,N_13592);
and U22332 (N_22332,N_13358,N_15407);
xnor U22333 (N_22333,N_13661,N_14148);
and U22334 (N_22334,N_14215,N_15375);
and U22335 (N_22335,N_12942,N_16246);
and U22336 (N_22336,N_13611,N_17012);
or U22337 (N_22337,N_17565,N_18011);
nor U22338 (N_22338,N_15605,N_14128);
and U22339 (N_22339,N_16638,N_16981);
or U22340 (N_22340,N_16821,N_12587);
or U22341 (N_22341,N_14344,N_18576);
xnor U22342 (N_22342,N_15634,N_18656);
nor U22343 (N_22343,N_17741,N_13502);
nor U22344 (N_22344,N_15943,N_15160);
xnor U22345 (N_22345,N_16895,N_16532);
or U22346 (N_22346,N_18248,N_17699);
and U22347 (N_22347,N_12689,N_16676);
nor U22348 (N_22348,N_14351,N_13648);
xnor U22349 (N_22349,N_16482,N_17745);
nor U22350 (N_22350,N_16456,N_15468);
or U22351 (N_22351,N_14059,N_15362);
nor U22352 (N_22352,N_18273,N_17459);
nor U22353 (N_22353,N_14628,N_16141);
xor U22354 (N_22354,N_15570,N_18056);
and U22355 (N_22355,N_15089,N_14054);
nand U22356 (N_22356,N_17094,N_15837);
nand U22357 (N_22357,N_15444,N_18262);
and U22358 (N_22358,N_13433,N_13921);
xnor U22359 (N_22359,N_17960,N_13257);
and U22360 (N_22360,N_16503,N_18342);
nand U22361 (N_22361,N_12969,N_17979);
nand U22362 (N_22362,N_13848,N_13096);
nor U22363 (N_22363,N_14994,N_14783);
nand U22364 (N_22364,N_15102,N_12655);
xnor U22365 (N_22365,N_18281,N_15103);
xnor U22366 (N_22366,N_15841,N_14357);
and U22367 (N_22367,N_15422,N_15691);
nor U22368 (N_22368,N_16328,N_15170);
xnor U22369 (N_22369,N_14666,N_16158);
xor U22370 (N_22370,N_14266,N_14423);
nand U22371 (N_22371,N_16568,N_18495);
or U22372 (N_22372,N_17528,N_13455);
nand U22373 (N_22373,N_18526,N_15826);
nor U22374 (N_22374,N_14811,N_13427);
nor U22375 (N_22375,N_18726,N_15706);
nand U22376 (N_22376,N_16386,N_17046);
and U22377 (N_22377,N_17383,N_17277);
nand U22378 (N_22378,N_16910,N_14291);
nand U22379 (N_22379,N_16135,N_18190);
xnor U22380 (N_22380,N_18516,N_16421);
xor U22381 (N_22381,N_12885,N_17069);
nor U22382 (N_22382,N_16499,N_17263);
nand U22383 (N_22383,N_17747,N_15883);
nand U22384 (N_22384,N_12637,N_12629);
nand U22385 (N_22385,N_17658,N_16296);
or U22386 (N_22386,N_15034,N_13911);
nand U22387 (N_22387,N_14693,N_13282);
nand U22388 (N_22388,N_12848,N_17344);
nand U22389 (N_22389,N_15268,N_13140);
or U22390 (N_22390,N_16231,N_15071);
and U22391 (N_22391,N_13767,N_16218);
xnor U22392 (N_22392,N_13307,N_12534);
nor U22393 (N_22393,N_18730,N_17218);
and U22394 (N_22394,N_16646,N_13888);
and U22395 (N_22395,N_16630,N_14075);
nor U22396 (N_22396,N_14113,N_14834);
or U22397 (N_22397,N_15620,N_18329);
nor U22398 (N_22398,N_18018,N_18504);
nand U22399 (N_22399,N_12912,N_18368);
nand U22400 (N_22400,N_15687,N_14049);
and U22401 (N_22401,N_17360,N_14936);
and U22402 (N_22402,N_13946,N_17836);
xor U22403 (N_22403,N_16105,N_15057);
or U22404 (N_22404,N_13176,N_13758);
or U22405 (N_22405,N_17106,N_16996);
xor U22406 (N_22406,N_16856,N_14850);
xnor U22407 (N_22407,N_12766,N_17312);
xnor U22408 (N_22408,N_13620,N_18440);
and U22409 (N_22409,N_15019,N_15098);
nor U22410 (N_22410,N_18279,N_17892);
nand U22411 (N_22411,N_18446,N_12661);
and U22412 (N_22412,N_14088,N_16632);
nor U22413 (N_22413,N_15491,N_12744);
and U22414 (N_22414,N_12782,N_17588);
nor U22415 (N_22415,N_12633,N_14565);
nand U22416 (N_22416,N_13923,N_17915);
nand U22417 (N_22417,N_16386,N_17300);
nand U22418 (N_22418,N_13971,N_17875);
nor U22419 (N_22419,N_16945,N_18394);
and U22420 (N_22420,N_16665,N_18491);
nor U22421 (N_22421,N_13894,N_14422);
or U22422 (N_22422,N_16699,N_18422);
and U22423 (N_22423,N_18374,N_18430);
and U22424 (N_22424,N_16149,N_15516);
nor U22425 (N_22425,N_14894,N_17921);
and U22426 (N_22426,N_14670,N_17207);
or U22427 (N_22427,N_14097,N_14145);
or U22428 (N_22428,N_13123,N_18374);
or U22429 (N_22429,N_15082,N_12693);
nor U22430 (N_22430,N_14128,N_18206);
xnor U22431 (N_22431,N_17316,N_15633);
nand U22432 (N_22432,N_13490,N_18184);
or U22433 (N_22433,N_16975,N_17320);
and U22434 (N_22434,N_17279,N_16856);
xnor U22435 (N_22435,N_13859,N_13087);
xor U22436 (N_22436,N_17525,N_16227);
or U22437 (N_22437,N_14574,N_17269);
nand U22438 (N_22438,N_16206,N_15897);
xor U22439 (N_22439,N_18162,N_16102);
and U22440 (N_22440,N_15835,N_16250);
or U22441 (N_22441,N_18236,N_16787);
and U22442 (N_22442,N_15930,N_17663);
nand U22443 (N_22443,N_16240,N_17165);
nor U22444 (N_22444,N_17470,N_17035);
and U22445 (N_22445,N_16632,N_15728);
nor U22446 (N_22446,N_16466,N_12724);
or U22447 (N_22447,N_12770,N_17221);
xnor U22448 (N_22448,N_17790,N_16945);
nand U22449 (N_22449,N_16787,N_15908);
nand U22450 (N_22450,N_16306,N_14476);
nor U22451 (N_22451,N_15360,N_12678);
or U22452 (N_22452,N_15936,N_12674);
and U22453 (N_22453,N_16512,N_16294);
and U22454 (N_22454,N_16004,N_18473);
or U22455 (N_22455,N_14401,N_18438);
or U22456 (N_22456,N_18209,N_17979);
or U22457 (N_22457,N_17665,N_16534);
or U22458 (N_22458,N_16542,N_15877);
nand U22459 (N_22459,N_14363,N_18692);
xor U22460 (N_22460,N_13865,N_16978);
or U22461 (N_22461,N_13991,N_14313);
nor U22462 (N_22462,N_18682,N_12908);
or U22463 (N_22463,N_17855,N_16126);
nand U22464 (N_22464,N_17157,N_14591);
nor U22465 (N_22465,N_13781,N_13970);
nor U22466 (N_22466,N_12858,N_14632);
xor U22467 (N_22467,N_15131,N_16578);
or U22468 (N_22468,N_12966,N_16095);
or U22469 (N_22469,N_15894,N_13356);
nand U22470 (N_22470,N_14998,N_12585);
nor U22471 (N_22471,N_12947,N_14619);
and U22472 (N_22472,N_16549,N_14763);
or U22473 (N_22473,N_13477,N_14557);
nor U22474 (N_22474,N_18192,N_16003);
or U22475 (N_22475,N_15680,N_18322);
or U22476 (N_22476,N_16516,N_17838);
or U22477 (N_22477,N_18420,N_18555);
or U22478 (N_22478,N_15444,N_15646);
or U22479 (N_22479,N_18447,N_17540);
and U22480 (N_22480,N_12558,N_14889);
nand U22481 (N_22481,N_17054,N_14695);
nor U22482 (N_22482,N_16436,N_18023);
nor U22483 (N_22483,N_15166,N_13378);
and U22484 (N_22484,N_12823,N_12906);
nor U22485 (N_22485,N_13299,N_17187);
xnor U22486 (N_22486,N_13161,N_16399);
nand U22487 (N_22487,N_17127,N_13487);
nor U22488 (N_22488,N_13142,N_14654);
nand U22489 (N_22489,N_14621,N_13086);
and U22490 (N_22490,N_15013,N_18396);
or U22491 (N_22491,N_12608,N_16289);
xnor U22492 (N_22492,N_17781,N_15874);
nand U22493 (N_22493,N_12535,N_17902);
nor U22494 (N_22494,N_14227,N_15603);
xor U22495 (N_22495,N_17632,N_17604);
nor U22496 (N_22496,N_15063,N_13649);
or U22497 (N_22497,N_17884,N_17321);
and U22498 (N_22498,N_12878,N_12730);
or U22499 (N_22499,N_16782,N_15777);
nor U22500 (N_22500,N_14746,N_14047);
nor U22501 (N_22501,N_14458,N_14815);
nand U22502 (N_22502,N_13874,N_17056);
or U22503 (N_22503,N_13737,N_15352);
nand U22504 (N_22504,N_14693,N_12763);
nand U22505 (N_22505,N_13510,N_18401);
or U22506 (N_22506,N_14948,N_18516);
or U22507 (N_22507,N_13471,N_14290);
nor U22508 (N_22508,N_18104,N_16317);
and U22509 (N_22509,N_17902,N_13904);
xnor U22510 (N_22510,N_13229,N_17087);
xor U22511 (N_22511,N_15371,N_14431);
and U22512 (N_22512,N_14676,N_12865);
nand U22513 (N_22513,N_13516,N_16308);
nor U22514 (N_22514,N_18408,N_15053);
nand U22515 (N_22515,N_14597,N_18485);
nor U22516 (N_22516,N_12690,N_17062);
or U22517 (N_22517,N_17783,N_13679);
and U22518 (N_22518,N_14251,N_14107);
and U22519 (N_22519,N_14555,N_17139);
nand U22520 (N_22520,N_17860,N_18006);
nor U22521 (N_22521,N_13115,N_13440);
nand U22522 (N_22522,N_18326,N_16660);
and U22523 (N_22523,N_16875,N_17711);
xnor U22524 (N_22524,N_17500,N_14232);
nand U22525 (N_22525,N_14382,N_15689);
or U22526 (N_22526,N_14737,N_15101);
xor U22527 (N_22527,N_13623,N_13921);
xor U22528 (N_22528,N_17151,N_17808);
xnor U22529 (N_22529,N_16561,N_14914);
nor U22530 (N_22530,N_16019,N_17743);
xnor U22531 (N_22531,N_17121,N_15232);
xnor U22532 (N_22532,N_16046,N_16126);
and U22533 (N_22533,N_13147,N_18338);
or U22534 (N_22534,N_18457,N_17508);
xnor U22535 (N_22535,N_15027,N_18287);
nand U22536 (N_22536,N_15991,N_16504);
nor U22537 (N_22537,N_14983,N_16820);
xnor U22538 (N_22538,N_13100,N_16625);
xnor U22539 (N_22539,N_18390,N_16234);
and U22540 (N_22540,N_18723,N_16790);
or U22541 (N_22541,N_16574,N_13641);
nor U22542 (N_22542,N_14798,N_18091);
and U22543 (N_22543,N_14594,N_13243);
and U22544 (N_22544,N_15638,N_13883);
nor U22545 (N_22545,N_17757,N_14401);
nand U22546 (N_22546,N_14218,N_16439);
xnor U22547 (N_22547,N_15719,N_17861);
nor U22548 (N_22548,N_16836,N_17380);
and U22549 (N_22549,N_13980,N_14463);
nor U22550 (N_22550,N_13349,N_14557);
xnor U22551 (N_22551,N_17985,N_15913);
xor U22552 (N_22552,N_16833,N_15112);
and U22553 (N_22553,N_15264,N_14803);
nor U22554 (N_22554,N_17215,N_16843);
or U22555 (N_22555,N_17455,N_15451);
xnor U22556 (N_22556,N_15927,N_16508);
or U22557 (N_22557,N_15742,N_15151);
xor U22558 (N_22558,N_15061,N_17281);
nor U22559 (N_22559,N_13026,N_16099);
nand U22560 (N_22560,N_12723,N_16878);
nand U22561 (N_22561,N_18694,N_13428);
nand U22562 (N_22562,N_14832,N_18530);
nor U22563 (N_22563,N_13271,N_16679);
nor U22564 (N_22564,N_13770,N_15787);
or U22565 (N_22565,N_16405,N_15640);
nor U22566 (N_22566,N_16810,N_17060);
nand U22567 (N_22567,N_12668,N_14373);
and U22568 (N_22568,N_12803,N_15594);
or U22569 (N_22569,N_15570,N_13560);
xnor U22570 (N_22570,N_16735,N_12962);
xnor U22571 (N_22571,N_13477,N_17417);
nor U22572 (N_22572,N_18086,N_15132);
or U22573 (N_22573,N_15092,N_14617);
and U22574 (N_22574,N_17441,N_16695);
xnor U22575 (N_22575,N_14903,N_13839);
xnor U22576 (N_22576,N_17919,N_14014);
xor U22577 (N_22577,N_15602,N_13851);
and U22578 (N_22578,N_16730,N_15256);
and U22579 (N_22579,N_14408,N_14854);
nand U22580 (N_22580,N_14311,N_18713);
nor U22581 (N_22581,N_14863,N_14160);
nor U22582 (N_22582,N_13891,N_17992);
nand U22583 (N_22583,N_13997,N_15883);
xor U22584 (N_22584,N_16228,N_16521);
and U22585 (N_22585,N_16738,N_13177);
and U22586 (N_22586,N_15877,N_14659);
nor U22587 (N_22587,N_15787,N_16156);
nor U22588 (N_22588,N_15908,N_14942);
or U22589 (N_22589,N_17996,N_18690);
xor U22590 (N_22590,N_15660,N_17662);
nor U22591 (N_22591,N_16232,N_16291);
xor U22592 (N_22592,N_15490,N_13918);
nor U22593 (N_22593,N_13158,N_12954);
nor U22594 (N_22594,N_13939,N_14180);
and U22595 (N_22595,N_13681,N_12958);
and U22596 (N_22596,N_17624,N_12666);
xor U22597 (N_22597,N_13683,N_18304);
nand U22598 (N_22598,N_17914,N_15849);
or U22599 (N_22599,N_13432,N_18226);
or U22600 (N_22600,N_16487,N_12541);
xnor U22601 (N_22601,N_13822,N_14819);
nor U22602 (N_22602,N_13201,N_12681);
and U22603 (N_22603,N_14214,N_16142);
or U22604 (N_22604,N_18274,N_15064);
or U22605 (N_22605,N_14240,N_18042);
or U22606 (N_22606,N_15846,N_13769);
or U22607 (N_22607,N_16840,N_14902);
and U22608 (N_22608,N_12826,N_15103);
and U22609 (N_22609,N_18250,N_14670);
nand U22610 (N_22610,N_12840,N_13943);
or U22611 (N_22611,N_17026,N_15106);
nor U22612 (N_22612,N_16912,N_18694);
nand U22613 (N_22613,N_17924,N_13422);
nor U22614 (N_22614,N_15723,N_18260);
or U22615 (N_22615,N_12852,N_17270);
xor U22616 (N_22616,N_14396,N_16733);
or U22617 (N_22617,N_17898,N_14653);
nand U22618 (N_22618,N_16249,N_17933);
or U22619 (N_22619,N_14311,N_17149);
nor U22620 (N_22620,N_16097,N_15265);
xor U22621 (N_22621,N_16531,N_14806);
or U22622 (N_22622,N_17767,N_17554);
or U22623 (N_22623,N_12715,N_12890);
or U22624 (N_22624,N_15838,N_16352);
or U22625 (N_22625,N_14334,N_15975);
xnor U22626 (N_22626,N_17191,N_15416);
or U22627 (N_22627,N_13350,N_14344);
or U22628 (N_22628,N_15550,N_18691);
xnor U22629 (N_22629,N_15474,N_18333);
nor U22630 (N_22630,N_17427,N_14753);
nand U22631 (N_22631,N_13627,N_15565);
nand U22632 (N_22632,N_16952,N_16687);
nor U22633 (N_22633,N_18304,N_12648);
or U22634 (N_22634,N_14939,N_14285);
nand U22635 (N_22635,N_13249,N_12856);
xor U22636 (N_22636,N_13252,N_12643);
nor U22637 (N_22637,N_14475,N_17241);
or U22638 (N_22638,N_13818,N_14602);
nor U22639 (N_22639,N_12957,N_13607);
xnor U22640 (N_22640,N_13132,N_14664);
xnor U22641 (N_22641,N_13478,N_15923);
or U22642 (N_22642,N_15321,N_17583);
nor U22643 (N_22643,N_16024,N_16589);
nor U22644 (N_22644,N_17490,N_15366);
nand U22645 (N_22645,N_17269,N_15568);
nor U22646 (N_22646,N_17481,N_17841);
xnor U22647 (N_22647,N_17832,N_17533);
xor U22648 (N_22648,N_15308,N_12669);
or U22649 (N_22649,N_18313,N_13548);
or U22650 (N_22650,N_17885,N_17837);
xnor U22651 (N_22651,N_18227,N_16217);
nand U22652 (N_22652,N_15432,N_13921);
nand U22653 (N_22653,N_16433,N_13402);
or U22654 (N_22654,N_16696,N_12868);
and U22655 (N_22655,N_12875,N_18234);
or U22656 (N_22656,N_15933,N_17681);
nor U22657 (N_22657,N_12754,N_18247);
and U22658 (N_22658,N_15651,N_17780);
xnor U22659 (N_22659,N_15677,N_14772);
and U22660 (N_22660,N_13595,N_18326);
or U22661 (N_22661,N_17510,N_13095);
nand U22662 (N_22662,N_18465,N_17281);
and U22663 (N_22663,N_14598,N_15657);
and U22664 (N_22664,N_16840,N_14627);
or U22665 (N_22665,N_14367,N_17693);
nand U22666 (N_22666,N_16231,N_17637);
and U22667 (N_22667,N_15980,N_18465);
nor U22668 (N_22668,N_12683,N_16057);
xor U22669 (N_22669,N_13256,N_18027);
xor U22670 (N_22670,N_15146,N_14980);
nand U22671 (N_22671,N_13582,N_18499);
nor U22672 (N_22672,N_17249,N_15754);
nor U22673 (N_22673,N_13361,N_15009);
xnor U22674 (N_22674,N_15595,N_16260);
nor U22675 (N_22675,N_18739,N_18294);
nor U22676 (N_22676,N_16081,N_17474);
nor U22677 (N_22677,N_17414,N_14024);
xor U22678 (N_22678,N_17900,N_18429);
nor U22679 (N_22679,N_12550,N_14049);
nand U22680 (N_22680,N_14563,N_16609);
nor U22681 (N_22681,N_12801,N_14313);
and U22682 (N_22682,N_13346,N_16308);
and U22683 (N_22683,N_15747,N_16855);
or U22684 (N_22684,N_15159,N_15348);
nand U22685 (N_22685,N_12526,N_13830);
nand U22686 (N_22686,N_13509,N_16527);
nor U22687 (N_22687,N_18123,N_18332);
xnor U22688 (N_22688,N_14910,N_14931);
and U22689 (N_22689,N_12659,N_13713);
xnor U22690 (N_22690,N_16912,N_16064);
or U22691 (N_22691,N_15569,N_13839);
or U22692 (N_22692,N_17054,N_16884);
or U22693 (N_22693,N_14314,N_13999);
xor U22694 (N_22694,N_18374,N_15585);
or U22695 (N_22695,N_17764,N_14260);
and U22696 (N_22696,N_13565,N_14996);
and U22697 (N_22697,N_15379,N_14458);
or U22698 (N_22698,N_15624,N_14982);
nand U22699 (N_22699,N_14135,N_17782);
nand U22700 (N_22700,N_16535,N_15321);
nand U22701 (N_22701,N_13552,N_12586);
xnor U22702 (N_22702,N_15052,N_18601);
nand U22703 (N_22703,N_13546,N_16218);
nand U22704 (N_22704,N_16623,N_18661);
xnor U22705 (N_22705,N_17401,N_16240);
xnor U22706 (N_22706,N_17623,N_16668);
and U22707 (N_22707,N_12621,N_17428);
nor U22708 (N_22708,N_16742,N_14119);
and U22709 (N_22709,N_17484,N_14201);
nor U22710 (N_22710,N_18144,N_18625);
and U22711 (N_22711,N_14142,N_17144);
nand U22712 (N_22712,N_14007,N_17727);
xnor U22713 (N_22713,N_12973,N_15951);
xnor U22714 (N_22714,N_17142,N_12952);
nand U22715 (N_22715,N_15561,N_15262);
and U22716 (N_22716,N_15267,N_14348);
and U22717 (N_22717,N_12822,N_16902);
and U22718 (N_22718,N_16362,N_13948);
and U22719 (N_22719,N_18381,N_15204);
and U22720 (N_22720,N_18706,N_16466);
or U22721 (N_22721,N_14251,N_18017);
nand U22722 (N_22722,N_15362,N_16348);
or U22723 (N_22723,N_12781,N_14521);
nor U22724 (N_22724,N_12997,N_18640);
xor U22725 (N_22725,N_16577,N_15260);
and U22726 (N_22726,N_17479,N_13238);
nand U22727 (N_22727,N_14948,N_16221);
nor U22728 (N_22728,N_15910,N_18521);
xnor U22729 (N_22729,N_15175,N_13390);
or U22730 (N_22730,N_16269,N_12674);
nor U22731 (N_22731,N_14123,N_18325);
xnor U22732 (N_22732,N_16156,N_16081);
and U22733 (N_22733,N_17424,N_16968);
nor U22734 (N_22734,N_16838,N_16120);
and U22735 (N_22735,N_15742,N_17791);
nand U22736 (N_22736,N_14182,N_14503);
nor U22737 (N_22737,N_16621,N_16996);
and U22738 (N_22738,N_16716,N_15534);
or U22739 (N_22739,N_13250,N_17340);
or U22740 (N_22740,N_15432,N_16022);
xnor U22741 (N_22741,N_16854,N_16298);
nor U22742 (N_22742,N_17939,N_13690);
xor U22743 (N_22743,N_14785,N_13572);
or U22744 (N_22744,N_16097,N_14181);
nand U22745 (N_22745,N_16039,N_16201);
xor U22746 (N_22746,N_14333,N_17440);
or U22747 (N_22747,N_17441,N_18243);
or U22748 (N_22748,N_14414,N_12986);
and U22749 (N_22749,N_18657,N_13681);
and U22750 (N_22750,N_17157,N_12996);
or U22751 (N_22751,N_18628,N_13094);
nand U22752 (N_22752,N_12954,N_14167);
xnor U22753 (N_22753,N_14315,N_17887);
xor U22754 (N_22754,N_16395,N_14821);
or U22755 (N_22755,N_14774,N_14666);
or U22756 (N_22756,N_13789,N_16199);
or U22757 (N_22757,N_15779,N_14669);
and U22758 (N_22758,N_17753,N_17998);
nor U22759 (N_22759,N_18479,N_13363);
nor U22760 (N_22760,N_12662,N_14948);
xor U22761 (N_22761,N_13305,N_17716);
xnor U22762 (N_22762,N_15883,N_13568);
nor U22763 (N_22763,N_18719,N_15632);
nor U22764 (N_22764,N_15553,N_15830);
and U22765 (N_22765,N_16248,N_12655);
xor U22766 (N_22766,N_14673,N_16070);
and U22767 (N_22767,N_13619,N_16261);
and U22768 (N_22768,N_18490,N_13061);
xnor U22769 (N_22769,N_13794,N_13772);
nand U22770 (N_22770,N_15245,N_18019);
nor U22771 (N_22771,N_18699,N_16409);
nand U22772 (N_22772,N_13308,N_18437);
nor U22773 (N_22773,N_14434,N_15954);
or U22774 (N_22774,N_13605,N_18003);
nand U22775 (N_22775,N_16620,N_16653);
nand U22776 (N_22776,N_16970,N_16800);
nand U22777 (N_22777,N_15311,N_18263);
nor U22778 (N_22778,N_17013,N_13721);
nor U22779 (N_22779,N_14637,N_17775);
nand U22780 (N_22780,N_15732,N_12563);
or U22781 (N_22781,N_12829,N_14301);
nand U22782 (N_22782,N_14332,N_13195);
nor U22783 (N_22783,N_13508,N_16052);
xor U22784 (N_22784,N_13689,N_17795);
xor U22785 (N_22785,N_12522,N_14374);
nor U22786 (N_22786,N_17422,N_15205);
nor U22787 (N_22787,N_15767,N_16969);
nand U22788 (N_22788,N_15487,N_16530);
or U22789 (N_22789,N_15555,N_15225);
and U22790 (N_22790,N_14428,N_14243);
and U22791 (N_22791,N_14443,N_13812);
nand U22792 (N_22792,N_13316,N_15936);
nand U22793 (N_22793,N_15268,N_17241);
or U22794 (N_22794,N_15755,N_15925);
or U22795 (N_22795,N_17922,N_14572);
nor U22796 (N_22796,N_12995,N_13098);
and U22797 (N_22797,N_14738,N_18248);
nand U22798 (N_22798,N_18655,N_14449);
and U22799 (N_22799,N_17758,N_18420);
or U22800 (N_22800,N_12857,N_17453);
nand U22801 (N_22801,N_17514,N_13228);
or U22802 (N_22802,N_17883,N_17639);
or U22803 (N_22803,N_15737,N_17120);
and U22804 (N_22804,N_14006,N_17199);
and U22805 (N_22805,N_15160,N_16863);
xor U22806 (N_22806,N_12767,N_17755);
nor U22807 (N_22807,N_18235,N_17012);
or U22808 (N_22808,N_15690,N_17427);
xor U22809 (N_22809,N_12816,N_17926);
nand U22810 (N_22810,N_15581,N_16385);
or U22811 (N_22811,N_17841,N_13349);
nor U22812 (N_22812,N_15186,N_16226);
nand U22813 (N_22813,N_14130,N_13720);
and U22814 (N_22814,N_18075,N_16518);
and U22815 (N_22815,N_14532,N_12790);
nand U22816 (N_22816,N_16853,N_15376);
nor U22817 (N_22817,N_17281,N_18496);
nor U22818 (N_22818,N_14627,N_18263);
xnor U22819 (N_22819,N_15268,N_12852);
nand U22820 (N_22820,N_17014,N_18160);
or U22821 (N_22821,N_16075,N_18492);
nor U22822 (N_22822,N_12704,N_16022);
xor U22823 (N_22823,N_12727,N_14699);
xnor U22824 (N_22824,N_13251,N_17493);
and U22825 (N_22825,N_12913,N_18179);
xor U22826 (N_22826,N_16940,N_17111);
nor U22827 (N_22827,N_16911,N_16143);
and U22828 (N_22828,N_13181,N_13429);
or U22829 (N_22829,N_16143,N_17192);
or U22830 (N_22830,N_17952,N_15612);
nand U22831 (N_22831,N_17515,N_17378);
xnor U22832 (N_22832,N_12514,N_18045);
nor U22833 (N_22833,N_13997,N_15682);
nor U22834 (N_22834,N_15560,N_17415);
nand U22835 (N_22835,N_16919,N_12762);
or U22836 (N_22836,N_12850,N_18117);
and U22837 (N_22837,N_18488,N_17528);
nor U22838 (N_22838,N_16845,N_14812);
or U22839 (N_22839,N_18433,N_14267);
or U22840 (N_22840,N_16572,N_15364);
or U22841 (N_22841,N_14194,N_12952);
xor U22842 (N_22842,N_16123,N_18259);
or U22843 (N_22843,N_16806,N_15970);
nand U22844 (N_22844,N_15963,N_12836);
xnor U22845 (N_22845,N_14163,N_16060);
nand U22846 (N_22846,N_13836,N_14858);
nand U22847 (N_22847,N_13089,N_14593);
xnor U22848 (N_22848,N_17569,N_18159);
nor U22849 (N_22849,N_12856,N_18342);
or U22850 (N_22850,N_15382,N_13544);
xnor U22851 (N_22851,N_12753,N_17066);
nand U22852 (N_22852,N_12856,N_17917);
or U22853 (N_22853,N_12691,N_15714);
xor U22854 (N_22854,N_16814,N_18225);
nor U22855 (N_22855,N_13034,N_14961);
xor U22856 (N_22856,N_13477,N_14200);
and U22857 (N_22857,N_14547,N_17890);
xor U22858 (N_22858,N_14429,N_14181);
or U22859 (N_22859,N_13532,N_17732);
nand U22860 (N_22860,N_13595,N_17655);
nor U22861 (N_22861,N_13918,N_15338);
and U22862 (N_22862,N_13785,N_17262);
nor U22863 (N_22863,N_17871,N_13309);
nand U22864 (N_22864,N_13613,N_17141);
xor U22865 (N_22865,N_17894,N_18366);
nor U22866 (N_22866,N_15373,N_16146);
or U22867 (N_22867,N_13047,N_17896);
nand U22868 (N_22868,N_18729,N_13614);
xnor U22869 (N_22869,N_17017,N_16761);
or U22870 (N_22870,N_14449,N_13067);
nand U22871 (N_22871,N_15690,N_14739);
nor U22872 (N_22872,N_14680,N_13702);
or U22873 (N_22873,N_15444,N_13452);
nor U22874 (N_22874,N_13023,N_13331);
xnor U22875 (N_22875,N_13629,N_16312);
and U22876 (N_22876,N_17468,N_17652);
nand U22877 (N_22877,N_15859,N_15891);
nand U22878 (N_22878,N_14306,N_14831);
and U22879 (N_22879,N_14278,N_15946);
or U22880 (N_22880,N_12740,N_15648);
xnor U22881 (N_22881,N_16973,N_17501);
or U22882 (N_22882,N_15188,N_17402);
or U22883 (N_22883,N_18382,N_17110);
nor U22884 (N_22884,N_13293,N_16248);
xor U22885 (N_22885,N_18167,N_17555);
and U22886 (N_22886,N_16477,N_14365);
xor U22887 (N_22887,N_13373,N_14891);
or U22888 (N_22888,N_18407,N_13279);
nor U22889 (N_22889,N_18077,N_12712);
or U22890 (N_22890,N_17094,N_17978);
or U22891 (N_22891,N_15785,N_14527);
or U22892 (N_22892,N_17699,N_13959);
nor U22893 (N_22893,N_16495,N_18623);
xnor U22894 (N_22894,N_14289,N_16376);
or U22895 (N_22895,N_16851,N_15124);
nand U22896 (N_22896,N_14386,N_17613);
or U22897 (N_22897,N_12905,N_17831);
and U22898 (N_22898,N_16754,N_13443);
xnor U22899 (N_22899,N_14029,N_17394);
or U22900 (N_22900,N_18511,N_18630);
nor U22901 (N_22901,N_12539,N_13705);
nand U22902 (N_22902,N_13323,N_12965);
and U22903 (N_22903,N_16873,N_14075);
xor U22904 (N_22904,N_13590,N_17016);
xnor U22905 (N_22905,N_18525,N_14014);
and U22906 (N_22906,N_12763,N_16441);
and U22907 (N_22907,N_13710,N_14998);
or U22908 (N_22908,N_14473,N_12754);
or U22909 (N_22909,N_14329,N_17037);
nand U22910 (N_22910,N_17770,N_14325);
or U22911 (N_22911,N_16978,N_16761);
or U22912 (N_22912,N_18406,N_15420);
nand U22913 (N_22913,N_15910,N_15097);
or U22914 (N_22914,N_13974,N_17136);
nor U22915 (N_22915,N_17088,N_12879);
xnor U22916 (N_22916,N_13298,N_15856);
nand U22917 (N_22917,N_14355,N_14999);
nand U22918 (N_22918,N_12532,N_13832);
or U22919 (N_22919,N_18006,N_14185);
xnor U22920 (N_22920,N_17053,N_18014);
nand U22921 (N_22921,N_15634,N_17311);
nand U22922 (N_22922,N_17030,N_16976);
nand U22923 (N_22923,N_16581,N_12963);
or U22924 (N_22924,N_13094,N_17714);
and U22925 (N_22925,N_13735,N_14359);
nand U22926 (N_22926,N_13398,N_17618);
xor U22927 (N_22927,N_13577,N_16259);
nand U22928 (N_22928,N_13952,N_15622);
or U22929 (N_22929,N_16060,N_14584);
xnor U22930 (N_22930,N_15740,N_14895);
nor U22931 (N_22931,N_17413,N_17150);
and U22932 (N_22932,N_14168,N_16973);
nor U22933 (N_22933,N_16946,N_16515);
nand U22934 (N_22934,N_17238,N_16712);
nand U22935 (N_22935,N_17866,N_14851);
nor U22936 (N_22936,N_16250,N_13335);
and U22937 (N_22937,N_15384,N_15192);
xor U22938 (N_22938,N_16780,N_17402);
xnor U22939 (N_22939,N_15353,N_17854);
xnor U22940 (N_22940,N_12569,N_15003);
xnor U22941 (N_22941,N_15557,N_13460);
nand U22942 (N_22942,N_13035,N_13609);
nand U22943 (N_22943,N_13717,N_13902);
nand U22944 (N_22944,N_16903,N_15975);
and U22945 (N_22945,N_17547,N_12659);
nor U22946 (N_22946,N_15665,N_15544);
xor U22947 (N_22947,N_13102,N_15478);
nor U22948 (N_22948,N_16861,N_15187);
and U22949 (N_22949,N_18377,N_15076);
or U22950 (N_22950,N_13590,N_18209);
xnor U22951 (N_22951,N_12553,N_17236);
or U22952 (N_22952,N_18746,N_14361);
nor U22953 (N_22953,N_18028,N_18355);
xor U22954 (N_22954,N_14162,N_17192);
xnor U22955 (N_22955,N_17717,N_13646);
nand U22956 (N_22956,N_14253,N_12558);
xnor U22957 (N_22957,N_15714,N_18218);
nand U22958 (N_22958,N_12529,N_14239);
nor U22959 (N_22959,N_17275,N_17829);
or U22960 (N_22960,N_16414,N_14439);
or U22961 (N_22961,N_15006,N_14476);
and U22962 (N_22962,N_15896,N_16096);
nor U22963 (N_22963,N_15420,N_13429);
nor U22964 (N_22964,N_15717,N_17091);
and U22965 (N_22965,N_16240,N_17853);
xor U22966 (N_22966,N_12587,N_15231);
xor U22967 (N_22967,N_17639,N_18553);
xor U22968 (N_22968,N_16475,N_14336);
and U22969 (N_22969,N_18088,N_15872);
and U22970 (N_22970,N_15326,N_13057);
xnor U22971 (N_22971,N_14401,N_15492);
xor U22972 (N_22972,N_15827,N_18354);
and U22973 (N_22973,N_15733,N_13977);
or U22974 (N_22974,N_15393,N_13294);
and U22975 (N_22975,N_17978,N_17939);
nor U22976 (N_22976,N_14995,N_17633);
xnor U22977 (N_22977,N_16055,N_16025);
nand U22978 (N_22978,N_16187,N_12934);
or U22979 (N_22979,N_14023,N_15225);
nand U22980 (N_22980,N_15204,N_12961);
xnor U22981 (N_22981,N_14981,N_16667);
and U22982 (N_22982,N_17197,N_12964);
and U22983 (N_22983,N_15084,N_16171);
nor U22984 (N_22984,N_17102,N_13541);
nor U22985 (N_22985,N_12757,N_15655);
nand U22986 (N_22986,N_15048,N_18560);
xnor U22987 (N_22987,N_13975,N_13123);
nor U22988 (N_22988,N_18707,N_15971);
or U22989 (N_22989,N_18300,N_15731);
nor U22990 (N_22990,N_15382,N_18266);
or U22991 (N_22991,N_14503,N_13902);
nand U22992 (N_22992,N_16166,N_15228);
or U22993 (N_22993,N_14959,N_12676);
or U22994 (N_22994,N_16775,N_14169);
nor U22995 (N_22995,N_15245,N_13971);
or U22996 (N_22996,N_16262,N_13821);
xor U22997 (N_22997,N_17700,N_18428);
and U22998 (N_22998,N_13494,N_18231);
nor U22999 (N_22999,N_15239,N_18405);
and U23000 (N_23000,N_16381,N_15200);
xnor U23001 (N_23001,N_17476,N_16501);
nor U23002 (N_23002,N_17405,N_12687);
or U23003 (N_23003,N_13892,N_14375);
xnor U23004 (N_23004,N_15663,N_18699);
nand U23005 (N_23005,N_17102,N_13215);
nor U23006 (N_23006,N_15157,N_15139);
xnor U23007 (N_23007,N_15419,N_17780);
nor U23008 (N_23008,N_15289,N_15941);
or U23009 (N_23009,N_18105,N_16649);
xnor U23010 (N_23010,N_15305,N_16377);
and U23011 (N_23011,N_14692,N_17355);
and U23012 (N_23012,N_18698,N_17243);
xnor U23013 (N_23013,N_15527,N_12632);
nor U23014 (N_23014,N_18480,N_14933);
and U23015 (N_23015,N_12947,N_17162);
or U23016 (N_23016,N_17543,N_14277);
nand U23017 (N_23017,N_18307,N_16869);
and U23018 (N_23018,N_12933,N_17522);
nor U23019 (N_23019,N_15501,N_17722);
or U23020 (N_23020,N_14235,N_16638);
and U23021 (N_23021,N_15752,N_16522);
or U23022 (N_23022,N_17809,N_17530);
xnor U23023 (N_23023,N_15042,N_13028);
nand U23024 (N_23024,N_18652,N_15158);
and U23025 (N_23025,N_14596,N_14816);
or U23026 (N_23026,N_12597,N_17484);
and U23027 (N_23027,N_16006,N_16250);
nand U23028 (N_23028,N_16211,N_15707);
nor U23029 (N_23029,N_16065,N_14965);
nand U23030 (N_23030,N_18469,N_14789);
nor U23031 (N_23031,N_16826,N_16074);
and U23032 (N_23032,N_15021,N_16252);
or U23033 (N_23033,N_17224,N_17402);
nor U23034 (N_23034,N_12807,N_17031);
nand U23035 (N_23035,N_14524,N_12699);
and U23036 (N_23036,N_16725,N_15651);
or U23037 (N_23037,N_13136,N_14721);
and U23038 (N_23038,N_14832,N_17990);
nor U23039 (N_23039,N_18274,N_18675);
nand U23040 (N_23040,N_17511,N_18100);
or U23041 (N_23041,N_15973,N_16298);
or U23042 (N_23042,N_16087,N_16542);
xor U23043 (N_23043,N_15902,N_15839);
xor U23044 (N_23044,N_14016,N_16345);
nor U23045 (N_23045,N_13805,N_14427);
xnor U23046 (N_23046,N_13044,N_18710);
and U23047 (N_23047,N_13350,N_15361);
or U23048 (N_23048,N_15749,N_13429);
nand U23049 (N_23049,N_13344,N_16321);
xnor U23050 (N_23050,N_14323,N_15421);
or U23051 (N_23051,N_18250,N_16921);
and U23052 (N_23052,N_13140,N_13564);
xnor U23053 (N_23053,N_17926,N_13717);
and U23054 (N_23054,N_14989,N_13609);
and U23055 (N_23055,N_17946,N_16672);
and U23056 (N_23056,N_18294,N_13467);
nor U23057 (N_23057,N_15137,N_17099);
nand U23058 (N_23058,N_14182,N_12541);
nand U23059 (N_23059,N_14156,N_18275);
nor U23060 (N_23060,N_18336,N_18245);
xnor U23061 (N_23061,N_15983,N_17185);
nor U23062 (N_23062,N_14511,N_16640);
or U23063 (N_23063,N_17874,N_13735);
nand U23064 (N_23064,N_14117,N_14931);
and U23065 (N_23065,N_14534,N_16252);
and U23066 (N_23066,N_18200,N_17502);
and U23067 (N_23067,N_14663,N_13062);
xor U23068 (N_23068,N_12795,N_14276);
and U23069 (N_23069,N_14538,N_14321);
xnor U23070 (N_23070,N_14419,N_15864);
nor U23071 (N_23071,N_18471,N_16546);
or U23072 (N_23072,N_15682,N_15753);
nand U23073 (N_23073,N_17593,N_18461);
and U23074 (N_23074,N_12864,N_18164);
xnor U23075 (N_23075,N_17769,N_16450);
and U23076 (N_23076,N_18141,N_14440);
nand U23077 (N_23077,N_16648,N_17861);
and U23078 (N_23078,N_14009,N_13020);
or U23079 (N_23079,N_14746,N_18509);
nand U23080 (N_23080,N_14035,N_13788);
or U23081 (N_23081,N_12893,N_13600);
nand U23082 (N_23082,N_15716,N_17759);
nor U23083 (N_23083,N_16640,N_16795);
or U23084 (N_23084,N_18430,N_16636);
nor U23085 (N_23085,N_17921,N_14912);
nand U23086 (N_23086,N_16786,N_18331);
xor U23087 (N_23087,N_14871,N_12864);
and U23088 (N_23088,N_18008,N_15503);
nor U23089 (N_23089,N_15569,N_16153);
nor U23090 (N_23090,N_15343,N_13837);
or U23091 (N_23091,N_14027,N_16196);
nand U23092 (N_23092,N_13164,N_17036);
or U23093 (N_23093,N_18096,N_14186);
nor U23094 (N_23094,N_16546,N_13079);
or U23095 (N_23095,N_15605,N_17499);
xnor U23096 (N_23096,N_17418,N_15318);
xnor U23097 (N_23097,N_13678,N_18210);
xor U23098 (N_23098,N_12964,N_12972);
nor U23099 (N_23099,N_18402,N_14246);
nand U23100 (N_23100,N_17863,N_18060);
or U23101 (N_23101,N_15514,N_15001);
xor U23102 (N_23102,N_15873,N_16138);
and U23103 (N_23103,N_14621,N_18585);
xnor U23104 (N_23104,N_17596,N_17201);
xor U23105 (N_23105,N_18369,N_14739);
and U23106 (N_23106,N_18670,N_14835);
or U23107 (N_23107,N_18483,N_16900);
and U23108 (N_23108,N_17829,N_12969);
or U23109 (N_23109,N_13367,N_17278);
nor U23110 (N_23110,N_13503,N_17542);
and U23111 (N_23111,N_17707,N_18346);
or U23112 (N_23112,N_16952,N_12754);
nand U23113 (N_23113,N_14689,N_16274);
or U23114 (N_23114,N_14901,N_17397);
and U23115 (N_23115,N_17133,N_13989);
and U23116 (N_23116,N_16332,N_15686);
nor U23117 (N_23117,N_15079,N_15821);
xor U23118 (N_23118,N_13475,N_15514);
nor U23119 (N_23119,N_17602,N_15450);
and U23120 (N_23120,N_18051,N_13907);
and U23121 (N_23121,N_17892,N_15718);
or U23122 (N_23122,N_13500,N_14559);
and U23123 (N_23123,N_13205,N_15176);
nand U23124 (N_23124,N_17975,N_14584);
nor U23125 (N_23125,N_16838,N_17843);
or U23126 (N_23126,N_18471,N_15551);
xnor U23127 (N_23127,N_13634,N_14905);
xor U23128 (N_23128,N_14793,N_16555);
nor U23129 (N_23129,N_17005,N_18476);
or U23130 (N_23130,N_14894,N_12780);
or U23131 (N_23131,N_16201,N_14842);
nor U23132 (N_23132,N_17884,N_12691);
nor U23133 (N_23133,N_14555,N_16112);
xor U23134 (N_23134,N_16009,N_18270);
or U23135 (N_23135,N_17380,N_18349);
nor U23136 (N_23136,N_17342,N_18077);
xnor U23137 (N_23137,N_14571,N_15794);
and U23138 (N_23138,N_17270,N_14553);
xor U23139 (N_23139,N_16733,N_17844);
and U23140 (N_23140,N_16747,N_13044);
or U23141 (N_23141,N_14360,N_14715);
xor U23142 (N_23142,N_14940,N_13385);
and U23143 (N_23143,N_15225,N_14781);
xnor U23144 (N_23144,N_13097,N_12997);
xor U23145 (N_23145,N_16855,N_14707);
nor U23146 (N_23146,N_17981,N_14593);
nand U23147 (N_23147,N_14379,N_17396);
nand U23148 (N_23148,N_15973,N_16284);
or U23149 (N_23149,N_14407,N_16309);
nand U23150 (N_23150,N_18738,N_14992);
or U23151 (N_23151,N_13367,N_18245);
xor U23152 (N_23152,N_18357,N_17502);
xnor U23153 (N_23153,N_15154,N_17332);
or U23154 (N_23154,N_18283,N_17525);
nor U23155 (N_23155,N_12588,N_18553);
and U23156 (N_23156,N_13790,N_16630);
xnor U23157 (N_23157,N_16226,N_17408);
and U23158 (N_23158,N_17794,N_15832);
nand U23159 (N_23159,N_13177,N_14671);
or U23160 (N_23160,N_17348,N_16946);
or U23161 (N_23161,N_18478,N_17228);
nand U23162 (N_23162,N_17048,N_13423);
or U23163 (N_23163,N_14984,N_16593);
nand U23164 (N_23164,N_17378,N_14550);
and U23165 (N_23165,N_13548,N_15100);
or U23166 (N_23166,N_14292,N_15075);
nor U23167 (N_23167,N_15051,N_12868);
xor U23168 (N_23168,N_18146,N_15002);
or U23169 (N_23169,N_14550,N_15766);
xnor U23170 (N_23170,N_18475,N_17529);
and U23171 (N_23171,N_16761,N_18145);
xor U23172 (N_23172,N_18716,N_15560);
xor U23173 (N_23173,N_16982,N_17423);
and U23174 (N_23174,N_13361,N_13686);
nor U23175 (N_23175,N_16714,N_15035);
nand U23176 (N_23176,N_16364,N_15362);
nand U23177 (N_23177,N_12852,N_14264);
or U23178 (N_23178,N_12772,N_16201);
xor U23179 (N_23179,N_18181,N_15834);
nor U23180 (N_23180,N_18156,N_17880);
or U23181 (N_23181,N_14292,N_17621);
nor U23182 (N_23182,N_13066,N_17396);
nor U23183 (N_23183,N_13979,N_13923);
xnor U23184 (N_23184,N_13374,N_17467);
and U23185 (N_23185,N_15545,N_15518);
and U23186 (N_23186,N_15316,N_16696);
nor U23187 (N_23187,N_13375,N_16275);
xnor U23188 (N_23188,N_18062,N_17145);
nor U23189 (N_23189,N_18388,N_12708);
xor U23190 (N_23190,N_15628,N_14101);
or U23191 (N_23191,N_18645,N_18609);
and U23192 (N_23192,N_17254,N_16974);
or U23193 (N_23193,N_18663,N_17839);
or U23194 (N_23194,N_18276,N_14576);
nor U23195 (N_23195,N_13227,N_18300);
nand U23196 (N_23196,N_18619,N_15401);
or U23197 (N_23197,N_15791,N_15121);
or U23198 (N_23198,N_17102,N_15860);
and U23199 (N_23199,N_18542,N_17777);
and U23200 (N_23200,N_15369,N_17364);
nor U23201 (N_23201,N_15140,N_18608);
and U23202 (N_23202,N_14022,N_13795);
xnor U23203 (N_23203,N_13253,N_15537);
nand U23204 (N_23204,N_14476,N_12517);
nor U23205 (N_23205,N_13501,N_14302);
xnor U23206 (N_23206,N_14977,N_16870);
or U23207 (N_23207,N_13668,N_14357);
nand U23208 (N_23208,N_12784,N_12820);
nand U23209 (N_23209,N_15632,N_15137);
xor U23210 (N_23210,N_16102,N_12572);
xor U23211 (N_23211,N_17363,N_12542);
nor U23212 (N_23212,N_16793,N_15391);
xnor U23213 (N_23213,N_15918,N_17333);
nand U23214 (N_23214,N_14043,N_14798);
and U23215 (N_23215,N_13868,N_17759);
nand U23216 (N_23216,N_14396,N_18301);
nand U23217 (N_23217,N_14507,N_15170);
nand U23218 (N_23218,N_13453,N_16955);
xor U23219 (N_23219,N_16373,N_13909);
nand U23220 (N_23220,N_15312,N_17333);
nor U23221 (N_23221,N_12912,N_13614);
nand U23222 (N_23222,N_15550,N_15657);
and U23223 (N_23223,N_15505,N_18428);
and U23224 (N_23224,N_15905,N_13561);
xnor U23225 (N_23225,N_13990,N_14839);
and U23226 (N_23226,N_15256,N_16697);
and U23227 (N_23227,N_17609,N_18041);
xor U23228 (N_23228,N_15644,N_18619);
nor U23229 (N_23229,N_15643,N_16495);
nand U23230 (N_23230,N_14224,N_17125);
nand U23231 (N_23231,N_15622,N_17857);
or U23232 (N_23232,N_14849,N_12731);
xnor U23233 (N_23233,N_13281,N_14086);
or U23234 (N_23234,N_17984,N_13789);
nand U23235 (N_23235,N_14694,N_14369);
and U23236 (N_23236,N_16506,N_13558);
xnor U23237 (N_23237,N_18023,N_17564);
xnor U23238 (N_23238,N_14273,N_16464);
nand U23239 (N_23239,N_16150,N_16407);
and U23240 (N_23240,N_16679,N_14605);
and U23241 (N_23241,N_17144,N_18138);
or U23242 (N_23242,N_14299,N_13737);
and U23243 (N_23243,N_16137,N_15216);
nor U23244 (N_23244,N_17985,N_17525);
xnor U23245 (N_23245,N_13135,N_13674);
and U23246 (N_23246,N_18606,N_16284);
xor U23247 (N_23247,N_13502,N_17495);
or U23248 (N_23248,N_13255,N_16939);
xor U23249 (N_23249,N_17629,N_13676);
or U23250 (N_23250,N_14695,N_15950);
nand U23251 (N_23251,N_13800,N_18239);
xnor U23252 (N_23252,N_15780,N_18602);
nor U23253 (N_23253,N_18599,N_17848);
nor U23254 (N_23254,N_17417,N_15239);
xor U23255 (N_23255,N_16156,N_17648);
xnor U23256 (N_23256,N_13270,N_15488);
and U23257 (N_23257,N_14277,N_16870);
nand U23258 (N_23258,N_13651,N_14902);
or U23259 (N_23259,N_15612,N_15613);
xnor U23260 (N_23260,N_12830,N_15795);
xor U23261 (N_23261,N_15758,N_12973);
nor U23262 (N_23262,N_14228,N_13017);
and U23263 (N_23263,N_16049,N_14272);
xnor U23264 (N_23264,N_14100,N_17384);
or U23265 (N_23265,N_18392,N_17145);
and U23266 (N_23266,N_14968,N_15220);
nor U23267 (N_23267,N_13773,N_17096);
xnor U23268 (N_23268,N_13271,N_16159);
or U23269 (N_23269,N_12985,N_15156);
nand U23270 (N_23270,N_16935,N_16235);
xor U23271 (N_23271,N_16648,N_17051);
nor U23272 (N_23272,N_18418,N_16654);
xor U23273 (N_23273,N_17062,N_14879);
xor U23274 (N_23274,N_18567,N_16118);
or U23275 (N_23275,N_17122,N_15787);
xnor U23276 (N_23276,N_16166,N_12859);
and U23277 (N_23277,N_14120,N_13759);
and U23278 (N_23278,N_15686,N_17061);
nand U23279 (N_23279,N_14214,N_13513);
nand U23280 (N_23280,N_14602,N_14574);
or U23281 (N_23281,N_15917,N_15192);
and U23282 (N_23282,N_18522,N_15889);
nor U23283 (N_23283,N_17001,N_15860);
xnor U23284 (N_23284,N_14394,N_13953);
nand U23285 (N_23285,N_18068,N_17858);
nor U23286 (N_23286,N_13009,N_14473);
or U23287 (N_23287,N_15098,N_16044);
nor U23288 (N_23288,N_13466,N_15610);
nor U23289 (N_23289,N_17284,N_13486);
xnor U23290 (N_23290,N_17052,N_15089);
and U23291 (N_23291,N_13876,N_12887);
or U23292 (N_23292,N_12963,N_17817);
xnor U23293 (N_23293,N_18217,N_14363);
nand U23294 (N_23294,N_17540,N_18125);
xor U23295 (N_23295,N_14322,N_17198);
nor U23296 (N_23296,N_14274,N_13761);
or U23297 (N_23297,N_12843,N_18105);
nand U23298 (N_23298,N_14874,N_15006);
nand U23299 (N_23299,N_17518,N_15947);
and U23300 (N_23300,N_14439,N_18384);
and U23301 (N_23301,N_15692,N_17666);
nor U23302 (N_23302,N_17618,N_17903);
or U23303 (N_23303,N_13809,N_16125);
nor U23304 (N_23304,N_17076,N_18040);
nand U23305 (N_23305,N_16505,N_14535);
nand U23306 (N_23306,N_13787,N_15566);
nor U23307 (N_23307,N_14972,N_16230);
nand U23308 (N_23308,N_18493,N_15535);
nand U23309 (N_23309,N_16953,N_15357);
or U23310 (N_23310,N_12559,N_17091);
nor U23311 (N_23311,N_14349,N_15335);
xnor U23312 (N_23312,N_12816,N_16465);
and U23313 (N_23313,N_16284,N_14702);
xor U23314 (N_23314,N_15678,N_17806);
and U23315 (N_23315,N_14128,N_13030);
nor U23316 (N_23316,N_14819,N_17304);
nor U23317 (N_23317,N_18715,N_15729);
and U23318 (N_23318,N_14009,N_15028);
nand U23319 (N_23319,N_14957,N_18573);
nor U23320 (N_23320,N_17696,N_18682);
nor U23321 (N_23321,N_17652,N_16023);
xor U23322 (N_23322,N_17047,N_16590);
or U23323 (N_23323,N_18637,N_16757);
xor U23324 (N_23324,N_16779,N_18468);
and U23325 (N_23325,N_18576,N_16322);
and U23326 (N_23326,N_14155,N_15566);
xor U23327 (N_23327,N_16242,N_16571);
or U23328 (N_23328,N_16887,N_15767);
xnor U23329 (N_23329,N_15836,N_17858);
or U23330 (N_23330,N_17882,N_12862);
xor U23331 (N_23331,N_16037,N_15925);
nand U23332 (N_23332,N_14470,N_16856);
xor U23333 (N_23333,N_18601,N_18074);
and U23334 (N_23334,N_14741,N_15002);
nor U23335 (N_23335,N_12606,N_14894);
and U23336 (N_23336,N_15328,N_14733);
xnor U23337 (N_23337,N_16889,N_14444);
xnor U23338 (N_23338,N_18408,N_16165);
and U23339 (N_23339,N_17034,N_17788);
or U23340 (N_23340,N_16526,N_15758);
nor U23341 (N_23341,N_15786,N_14485);
nand U23342 (N_23342,N_16061,N_18245);
nand U23343 (N_23343,N_14247,N_16527);
nand U23344 (N_23344,N_15957,N_17459);
or U23345 (N_23345,N_13697,N_15384);
and U23346 (N_23346,N_16804,N_16801);
or U23347 (N_23347,N_13813,N_15276);
nor U23348 (N_23348,N_18127,N_15703);
and U23349 (N_23349,N_15261,N_14006);
xnor U23350 (N_23350,N_17909,N_13406);
or U23351 (N_23351,N_17596,N_13815);
nor U23352 (N_23352,N_15406,N_18623);
nand U23353 (N_23353,N_14855,N_15905);
and U23354 (N_23354,N_17137,N_15725);
nor U23355 (N_23355,N_13211,N_16314);
or U23356 (N_23356,N_18432,N_13409);
and U23357 (N_23357,N_17318,N_17233);
xnor U23358 (N_23358,N_13058,N_18153);
or U23359 (N_23359,N_17802,N_16451);
and U23360 (N_23360,N_15782,N_16825);
xnor U23361 (N_23361,N_16812,N_18733);
nand U23362 (N_23362,N_12797,N_18501);
nand U23363 (N_23363,N_14458,N_13277);
xor U23364 (N_23364,N_15223,N_15963);
nand U23365 (N_23365,N_16099,N_15230);
nand U23366 (N_23366,N_14983,N_14265);
or U23367 (N_23367,N_16947,N_17136);
nor U23368 (N_23368,N_18398,N_14954);
and U23369 (N_23369,N_17727,N_13655);
nor U23370 (N_23370,N_18604,N_17147);
nand U23371 (N_23371,N_14177,N_15844);
or U23372 (N_23372,N_18748,N_18644);
nor U23373 (N_23373,N_14066,N_18398);
and U23374 (N_23374,N_16456,N_17756);
nor U23375 (N_23375,N_16840,N_13611);
and U23376 (N_23376,N_17574,N_14898);
nand U23377 (N_23377,N_16194,N_14088);
nor U23378 (N_23378,N_13172,N_15857);
nor U23379 (N_23379,N_14591,N_18100);
or U23380 (N_23380,N_17542,N_13216);
or U23381 (N_23381,N_13105,N_13923);
and U23382 (N_23382,N_16102,N_12834);
nand U23383 (N_23383,N_14838,N_13406);
nand U23384 (N_23384,N_17486,N_17069);
and U23385 (N_23385,N_13869,N_16164);
xor U23386 (N_23386,N_15772,N_15341);
or U23387 (N_23387,N_17887,N_12519);
nor U23388 (N_23388,N_16448,N_15774);
nor U23389 (N_23389,N_18593,N_16458);
and U23390 (N_23390,N_13799,N_14832);
and U23391 (N_23391,N_12870,N_14308);
and U23392 (N_23392,N_18478,N_13904);
or U23393 (N_23393,N_13802,N_14189);
nor U23394 (N_23394,N_18387,N_16960);
nand U23395 (N_23395,N_13010,N_17935);
nand U23396 (N_23396,N_14915,N_17091);
nor U23397 (N_23397,N_16917,N_14789);
and U23398 (N_23398,N_15675,N_17200);
nand U23399 (N_23399,N_14356,N_16498);
nand U23400 (N_23400,N_15153,N_17500);
nor U23401 (N_23401,N_16116,N_16589);
and U23402 (N_23402,N_12849,N_13557);
nand U23403 (N_23403,N_18615,N_14495);
or U23404 (N_23404,N_17208,N_17519);
xor U23405 (N_23405,N_15755,N_15556);
and U23406 (N_23406,N_17712,N_15482);
nor U23407 (N_23407,N_18013,N_13036);
nor U23408 (N_23408,N_15353,N_12520);
xor U23409 (N_23409,N_16662,N_14897);
and U23410 (N_23410,N_15080,N_15878);
nand U23411 (N_23411,N_18643,N_15390);
nor U23412 (N_23412,N_17711,N_18280);
xnor U23413 (N_23413,N_13385,N_16514);
xnor U23414 (N_23414,N_13447,N_14457);
or U23415 (N_23415,N_16378,N_14353);
or U23416 (N_23416,N_18193,N_17572);
and U23417 (N_23417,N_15243,N_12731);
or U23418 (N_23418,N_12596,N_13429);
or U23419 (N_23419,N_13162,N_15720);
or U23420 (N_23420,N_18624,N_14017);
xor U23421 (N_23421,N_15773,N_13289);
nor U23422 (N_23422,N_18499,N_17923);
xor U23423 (N_23423,N_18581,N_15418);
xor U23424 (N_23424,N_13041,N_17884);
and U23425 (N_23425,N_13920,N_17332);
nor U23426 (N_23426,N_18126,N_12904);
nand U23427 (N_23427,N_15557,N_12751);
nor U23428 (N_23428,N_13991,N_16719);
nand U23429 (N_23429,N_12788,N_13586);
and U23430 (N_23430,N_17078,N_15607);
and U23431 (N_23431,N_16300,N_16098);
or U23432 (N_23432,N_14290,N_16623);
nand U23433 (N_23433,N_12639,N_16287);
nand U23434 (N_23434,N_13848,N_18041);
or U23435 (N_23435,N_17502,N_15744);
nand U23436 (N_23436,N_16656,N_13958);
nand U23437 (N_23437,N_17509,N_14708);
or U23438 (N_23438,N_17534,N_15918);
nand U23439 (N_23439,N_14501,N_15943);
and U23440 (N_23440,N_14265,N_17719);
and U23441 (N_23441,N_17334,N_16845);
nor U23442 (N_23442,N_13030,N_12827);
xnor U23443 (N_23443,N_13937,N_16343);
and U23444 (N_23444,N_13083,N_17828);
nand U23445 (N_23445,N_18533,N_15457);
nand U23446 (N_23446,N_15323,N_13842);
nand U23447 (N_23447,N_16762,N_13620);
and U23448 (N_23448,N_14251,N_15513);
xor U23449 (N_23449,N_15511,N_14468);
xor U23450 (N_23450,N_16809,N_16401);
nand U23451 (N_23451,N_18013,N_13894);
or U23452 (N_23452,N_14058,N_18247);
and U23453 (N_23453,N_13648,N_15174);
or U23454 (N_23454,N_15604,N_15959);
xnor U23455 (N_23455,N_14143,N_13362);
or U23456 (N_23456,N_13955,N_13746);
nand U23457 (N_23457,N_15912,N_15256);
or U23458 (N_23458,N_16746,N_13572);
or U23459 (N_23459,N_13987,N_17786);
or U23460 (N_23460,N_17038,N_14616);
and U23461 (N_23461,N_18654,N_17115);
xnor U23462 (N_23462,N_18237,N_12777);
nand U23463 (N_23463,N_13083,N_16660);
nand U23464 (N_23464,N_16340,N_17522);
and U23465 (N_23465,N_15652,N_18490);
or U23466 (N_23466,N_14558,N_14221);
and U23467 (N_23467,N_14825,N_17850);
nand U23468 (N_23468,N_16376,N_18474);
and U23469 (N_23469,N_13646,N_12698);
xnor U23470 (N_23470,N_18648,N_13408);
and U23471 (N_23471,N_18308,N_17533);
nor U23472 (N_23472,N_12964,N_18693);
and U23473 (N_23473,N_12727,N_16234);
and U23474 (N_23474,N_15251,N_16142);
nand U23475 (N_23475,N_13456,N_13912);
and U23476 (N_23476,N_14225,N_12605);
nor U23477 (N_23477,N_13292,N_16407);
and U23478 (N_23478,N_13288,N_15676);
and U23479 (N_23479,N_17299,N_12823);
or U23480 (N_23480,N_14760,N_14024);
nand U23481 (N_23481,N_13532,N_16603);
nor U23482 (N_23482,N_16469,N_14660);
nand U23483 (N_23483,N_17127,N_15062);
or U23484 (N_23484,N_17664,N_16655);
and U23485 (N_23485,N_16836,N_17005);
and U23486 (N_23486,N_12912,N_16784);
xor U23487 (N_23487,N_14063,N_12735);
xor U23488 (N_23488,N_13016,N_14496);
and U23489 (N_23489,N_13199,N_15029);
nand U23490 (N_23490,N_16111,N_17759);
nand U23491 (N_23491,N_15854,N_17115);
nand U23492 (N_23492,N_16930,N_16580);
and U23493 (N_23493,N_16897,N_15351);
nor U23494 (N_23494,N_12996,N_18341);
xnor U23495 (N_23495,N_14122,N_15913);
nand U23496 (N_23496,N_17462,N_18537);
nand U23497 (N_23497,N_14647,N_16250);
xor U23498 (N_23498,N_14550,N_14632);
and U23499 (N_23499,N_17149,N_14023);
nand U23500 (N_23500,N_14384,N_12696);
nor U23501 (N_23501,N_17578,N_12816);
nor U23502 (N_23502,N_14960,N_17016);
or U23503 (N_23503,N_18299,N_14397);
nand U23504 (N_23504,N_12993,N_17971);
xnor U23505 (N_23505,N_13887,N_16957);
xor U23506 (N_23506,N_17288,N_14034);
nor U23507 (N_23507,N_12884,N_14843);
nand U23508 (N_23508,N_15965,N_14537);
xor U23509 (N_23509,N_13436,N_13003);
nand U23510 (N_23510,N_15074,N_17863);
xnor U23511 (N_23511,N_17217,N_15050);
xnor U23512 (N_23512,N_14586,N_15856);
and U23513 (N_23513,N_15632,N_18265);
nor U23514 (N_23514,N_13390,N_14648);
xnor U23515 (N_23515,N_16074,N_13899);
nor U23516 (N_23516,N_17354,N_15445);
or U23517 (N_23517,N_17036,N_18017);
and U23518 (N_23518,N_15557,N_15588);
xnor U23519 (N_23519,N_18358,N_16973);
xnor U23520 (N_23520,N_15071,N_15162);
xor U23521 (N_23521,N_15352,N_14424);
and U23522 (N_23522,N_14323,N_16029);
nor U23523 (N_23523,N_18446,N_16933);
or U23524 (N_23524,N_17065,N_14789);
nand U23525 (N_23525,N_14185,N_12754);
or U23526 (N_23526,N_15860,N_12605);
and U23527 (N_23527,N_17889,N_15724);
xnor U23528 (N_23528,N_13799,N_18172);
nor U23529 (N_23529,N_14815,N_15406);
and U23530 (N_23530,N_16489,N_14123);
xor U23531 (N_23531,N_14792,N_15211);
nand U23532 (N_23532,N_17296,N_18409);
nor U23533 (N_23533,N_15062,N_18665);
nand U23534 (N_23534,N_13364,N_16229);
or U23535 (N_23535,N_15687,N_15024);
xor U23536 (N_23536,N_15066,N_12920);
or U23537 (N_23537,N_12548,N_12805);
or U23538 (N_23538,N_18118,N_18635);
nor U23539 (N_23539,N_13140,N_17385);
and U23540 (N_23540,N_12925,N_13474);
xor U23541 (N_23541,N_13887,N_13371);
or U23542 (N_23542,N_13724,N_15107);
nand U23543 (N_23543,N_15500,N_16474);
nor U23544 (N_23544,N_16330,N_14321);
nor U23545 (N_23545,N_17238,N_17958);
nor U23546 (N_23546,N_14199,N_13487);
and U23547 (N_23547,N_17630,N_13964);
and U23548 (N_23548,N_15543,N_16891);
or U23549 (N_23549,N_14921,N_16089);
xor U23550 (N_23550,N_17193,N_14061);
nor U23551 (N_23551,N_14052,N_17139);
nor U23552 (N_23552,N_17577,N_16208);
xor U23553 (N_23553,N_18178,N_16972);
nor U23554 (N_23554,N_13075,N_17383);
and U23555 (N_23555,N_15340,N_16560);
xor U23556 (N_23556,N_16199,N_13714);
or U23557 (N_23557,N_17802,N_12720);
nand U23558 (N_23558,N_17590,N_17470);
nand U23559 (N_23559,N_14750,N_16547);
nand U23560 (N_23560,N_16514,N_14563);
xnor U23561 (N_23561,N_13340,N_18678);
xor U23562 (N_23562,N_13438,N_15406);
nand U23563 (N_23563,N_18145,N_14974);
and U23564 (N_23564,N_18222,N_18619);
nor U23565 (N_23565,N_15601,N_14339);
or U23566 (N_23566,N_12760,N_14174);
nand U23567 (N_23567,N_16540,N_13891);
and U23568 (N_23568,N_16092,N_17759);
and U23569 (N_23569,N_14427,N_12790);
nand U23570 (N_23570,N_13647,N_15125);
nor U23571 (N_23571,N_15590,N_17275);
or U23572 (N_23572,N_15733,N_16987);
nor U23573 (N_23573,N_14411,N_18250);
or U23574 (N_23574,N_15670,N_16061);
nand U23575 (N_23575,N_14204,N_16378);
or U23576 (N_23576,N_13778,N_13445);
and U23577 (N_23577,N_13379,N_13491);
nand U23578 (N_23578,N_12963,N_15665);
nor U23579 (N_23579,N_12628,N_18371);
and U23580 (N_23580,N_15976,N_18113);
and U23581 (N_23581,N_16100,N_18328);
or U23582 (N_23582,N_15611,N_13605);
xnor U23583 (N_23583,N_16879,N_18006);
or U23584 (N_23584,N_13703,N_17462);
nor U23585 (N_23585,N_16279,N_17369);
and U23586 (N_23586,N_12812,N_16223);
or U23587 (N_23587,N_17809,N_15167);
or U23588 (N_23588,N_12500,N_18412);
nor U23589 (N_23589,N_17311,N_13452);
and U23590 (N_23590,N_13049,N_16051);
and U23591 (N_23591,N_18453,N_17649);
nand U23592 (N_23592,N_13619,N_15703);
nand U23593 (N_23593,N_16859,N_17841);
xnor U23594 (N_23594,N_13436,N_18362);
and U23595 (N_23595,N_13546,N_16718);
xnor U23596 (N_23596,N_16672,N_14769);
or U23597 (N_23597,N_16427,N_18161);
and U23598 (N_23598,N_13794,N_14255);
or U23599 (N_23599,N_13102,N_16211);
nand U23600 (N_23600,N_13747,N_17095);
or U23601 (N_23601,N_15099,N_18108);
or U23602 (N_23602,N_15174,N_16132);
and U23603 (N_23603,N_18619,N_16099);
nand U23604 (N_23604,N_18149,N_16067);
or U23605 (N_23605,N_14605,N_15604);
or U23606 (N_23606,N_17350,N_18152);
and U23607 (N_23607,N_16062,N_18138);
and U23608 (N_23608,N_18359,N_12661);
nand U23609 (N_23609,N_13818,N_16125);
nand U23610 (N_23610,N_18532,N_18502);
or U23611 (N_23611,N_17651,N_16960);
or U23612 (N_23612,N_14665,N_16323);
nand U23613 (N_23613,N_15872,N_17943);
or U23614 (N_23614,N_16788,N_15907);
and U23615 (N_23615,N_14871,N_15334);
and U23616 (N_23616,N_13147,N_17460);
or U23617 (N_23617,N_14469,N_15624);
nor U23618 (N_23618,N_18632,N_15139);
nand U23619 (N_23619,N_18198,N_13399);
xor U23620 (N_23620,N_17610,N_13801);
or U23621 (N_23621,N_13657,N_13876);
nand U23622 (N_23622,N_16055,N_13328);
or U23623 (N_23623,N_17185,N_12767);
nor U23624 (N_23624,N_13088,N_14352);
or U23625 (N_23625,N_14308,N_14685);
xnor U23626 (N_23626,N_15397,N_16160);
and U23627 (N_23627,N_18594,N_13898);
xnor U23628 (N_23628,N_15648,N_17914);
xnor U23629 (N_23629,N_18227,N_17600);
nor U23630 (N_23630,N_18372,N_15830);
xor U23631 (N_23631,N_15720,N_17612);
or U23632 (N_23632,N_13955,N_12958);
nand U23633 (N_23633,N_14705,N_16279);
or U23634 (N_23634,N_15898,N_14687);
or U23635 (N_23635,N_12605,N_17437);
or U23636 (N_23636,N_15545,N_15295);
and U23637 (N_23637,N_14310,N_15107);
and U23638 (N_23638,N_12540,N_15704);
and U23639 (N_23639,N_13673,N_17224);
nand U23640 (N_23640,N_13595,N_17165);
or U23641 (N_23641,N_13738,N_12526);
nor U23642 (N_23642,N_15898,N_13951);
nor U23643 (N_23643,N_12724,N_14901);
nand U23644 (N_23644,N_17638,N_13229);
and U23645 (N_23645,N_12965,N_18115);
nor U23646 (N_23646,N_17945,N_17049);
or U23647 (N_23647,N_16011,N_16888);
xnor U23648 (N_23648,N_12605,N_15310);
nor U23649 (N_23649,N_14548,N_13203);
nand U23650 (N_23650,N_16248,N_17200);
nor U23651 (N_23651,N_13043,N_14510);
and U23652 (N_23652,N_15989,N_13253);
nand U23653 (N_23653,N_14605,N_14138);
and U23654 (N_23654,N_16420,N_14889);
xor U23655 (N_23655,N_15453,N_14726);
nand U23656 (N_23656,N_17228,N_13467);
nand U23657 (N_23657,N_15337,N_17412);
nand U23658 (N_23658,N_15892,N_17180);
or U23659 (N_23659,N_18742,N_14296);
and U23660 (N_23660,N_16301,N_17230);
nand U23661 (N_23661,N_16576,N_16662);
xnor U23662 (N_23662,N_12583,N_15736);
or U23663 (N_23663,N_17351,N_14616);
or U23664 (N_23664,N_15570,N_13374);
nor U23665 (N_23665,N_14540,N_15700);
and U23666 (N_23666,N_15560,N_13951);
xor U23667 (N_23667,N_18556,N_13810);
and U23668 (N_23668,N_18289,N_17995);
nand U23669 (N_23669,N_17081,N_15938);
nand U23670 (N_23670,N_16456,N_13228);
or U23671 (N_23671,N_15176,N_14266);
xor U23672 (N_23672,N_14996,N_13920);
nor U23673 (N_23673,N_17311,N_12503);
nand U23674 (N_23674,N_17302,N_16045);
or U23675 (N_23675,N_14174,N_15745);
or U23676 (N_23676,N_14169,N_18334);
or U23677 (N_23677,N_13758,N_15326);
xnor U23678 (N_23678,N_14143,N_16497);
or U23679 (N_23679,N_12935,N_13709);
xor U23680 (N_23680,N_18202,N_13807);
nand U23681 (N_23681,N_16412,N_15313);
or U23682 (N_23682,N_16896,N_13932);
and U23683 (N_23683,N_15484,N_12768);
or U23684 (N_23684,N_13503,N_16295);
nor U23685 (N_23685,N_16667,N_13279);
and U23686 (N_23686,N_17264,N_13929);
or U23687 (N_23687,N_17309,N_17148);
xor U23688 (N_23688,N_15386,N_17529);
nand U23689 (N_23689,N_14396,N_15334);
nor U23690 (N_23690,N_14593,N_16812);
nor U23691 (N_23691,N_14048,N_14617);
nand U23692 (N_23692,N_13355,N_16622);
nand U23693 (N_23693,N_18013,N_12686);
nor U23694 (N_23694,N_13577,N_13984);
nor U23695 (N_23695,N_13387,N_17018);
and U23696 (N_23696,N_16256,N_17572);
xor U23697 (N_23697,N_12920,N_17649);
or U23698 (N_23698,N_12884,N_14315);
xnor U23699 (N_23699,N_17791,N_14422);
nor U23700 (N_23700,N_13959,N_14417);
or U23701 (N_23701,N_15387,N_17211);
xnor U23702 (N_23702,N_16381,N_15479);
and U23703 (N_23703,N_14249,N_12914);
nand U23704 (N_23704,N_13518,N_18624);
nor U23705 (N_23705,N_18438,N_17687);
and U23706 (N_23706,N_15203,N_14923);
nand U23707 (N_23707,N_17373,N_12835);
or U23708 (N_23708,N_18001,N_17293);
xor U23709 (N_23709,N_18280,N_13108);
or U23710 (N_23710,N_12712,N_17654);
and U23711 (N_23711,N_13513,N_18341);
xnor U23712 (N_23712,N_17210,N_15014);
xor U23713 (N_23713,N_15602,N_14989);
or U23714 (N_23714,N_12794,N_15091);
nor U23715 (N_23715,N_17395,N_12812);
and U23716 (N_23716,N_18140,N_18413);
nand U23717 (N_23717,N_14838,N_16770);
or U23718 (N_23718,N_18147,N_15578);
nand U23719 (N_23719,N_16602,N_14069);
nor U23720 (N_23720,N_13594,N_14477);
nand U23721 (N_23721,N_17555,N_14501);
nor U23722 (N_23722,N_17914,N_14276);
nand U23723 (N_23723,N_12539,N_15700);
and U23724 (N_23724,N_17106,N_16196);
nor U23725 (N_23725,N_18494,N_18357);
nand U23726 (N_23726,N_14566,N_12885);
xor U23727 (N_23727,N_16365,N_16277);
nor U23728 (N_23728,N_13084,N_16306);
and U23729 (N_23729,N_16254,N_12997);
nand U23730 (N_23730,N_15367,N_18603);
and U23731 (N_23731,N_12822,N_18656);
or U23732 (N_23732,N_13693,N_13406);
and U23733 (N_23733,N_12561,N_13264);
or U23734 (N_23734,N_18395,N_14209);
and U23735 (N_23735,N_13897,N_18206);
and U23736 (N_23736,N_18647,N_18749);
and U23737 (N_23737,N_15680,N_17305);
nor U23738 (N_23738,N_16082,N_14163);
nand U23739 (N_23739,N_18496,N_15513);
nand U23740 (N_23740,N_13685,N_18704);
xor U23741 (N_23741,N_14842,N_13450);
or U23742 (N_23742,N_16132,N_13746);
xnor U23743 (N_23743,N_13100,N_17688);
nand U23744 (N_23744,N_18162,N_13613);
or U23745 (N_23745,N_12894,N_18689);
and U23746 (N_23746,N_13232,N_13606);
or U23747 (N_23747,N_17807,N_16490);
nor U23748 (N_23748,N_15739,N_18202);
nor U23749 (N_23749,N_18142,N_17743);
or U23750 (N_23750,N_17282,N_14467);
and U23751 (N_23751,N_14276,N_12755);
or U23752 (N_23752,N_18227,N_18232);
nor U23753 (N_23753,N_16075,N_17715);
or U23754 (N_23754,N_13640,N_17946);
or U23755 (N_23755,N_12928,N_12548);
nor U23756 (N_23756,N_14009,N_15179);
xor U23757 (N_23757,N_17595,N_18451);
nor U23758 (N_23758,N_17914,N_16951);
and U23759 (N_23759,N_14920,N_16563);
or U23760 (N_23760,N_14146,N_18062);
xnor U23761 (N_23761,N_16309,N_17765);
nor U23762 (N_23762,N_18553,N_17192);
nor U23763 (N_23763,N_12645,N_18433);
nand U23764 (N_23764,N_12651,N_17406);
and U23765 (N_23765,N_17636,N_16914);
or U23766 (N_23766,N_14442,N_16097);
nor U23767 (N_23767,N_17179,N_15735);
and U23768 (N_23768,N_15079,N_14976);
nand U23769 (N_23769,N_16076,N_17747);
nand U23770 (N_23770,N_13978,N_17034);
xnor U23771 (N_23771,N_13337,N_17820);
nand U23772 (N_23772,N_12918,N_16032);
and U23773 (N_23773,N_13085,N_15173);
nand U23774 (N_23774,N_14804,N_18664);
xnor U23775 (N_23775,N_17288,N_16907);
and U23776 (N_23776,N_14051,N_17883);
xor U23777 (N_23777,N_18705,N_16134);
or U23778 (N_23778,N_15553,N_18446);
nand U23779 (N_23779,N_15457,N_14049);
nand U23780 (N_23780,N_16693,N_16162);
and U23781 (N_23781,N_17955,N_17474);
nand U23782 (N_23782,N_17107,N_15591);
xor U23783 (N_23783,N_15729,N_12643);
or U23784 (N_23784,N_13602,N_16034);
or U23785 (N_23785,N_16168,N_13416);
nand U23786 (N_23786,N_15758,N_12725);
xor U23787 (N_23787,N_14680,N_14879);
or U23788 (N_23788,N_14469,N_16241);
nor U23789 (N_23789,N_17566,N_18407);
nand U23790 (N_23790,N_14922,N_17837);
nand U23791 (N_23791,N_17740,N_18074);
or U23792 (N_23792,N_17853,N_13521);
xor U23793 (N_23793,N_17198,N_15997);
xnor U23794 (N_23794,N_13813,N_15767);
or U23795 (N_23795,N_15947,N_13423);
nor U23796 (N_23796,N_15436,N_13693);
nor U23797 (N_23797,N_17430,N_14947);
and U23798 (N_23798,N_15214,N_18060);
xor U23799 (N_23799,N_14362,N_18128);
or U23800 (N_23800,N_13893,N_14278);
or U23801 (N_23801,N_12816,N_18486);
nor U23802 (N_23802,N_13996,N_18259);
nor U23803 (N_23803,N_12579,N_14926);
and U23804 (N_23804,N_16940,N_15492);
xor U23805 (N_23805,N_18660,N_13706);
nand U23806 (N_23806,N_14223,N_14097);
nor U23807 (N_23807,N_13992,N_13171);
xor U23808 (N_23808,N_14293,N_12745);
or U23809 (N_23809,N_18158,N_15658);
or U23810 (N_23810,N_13089,N_18337);
xor U23811 (N_23811,N_18480,N_14553);
nor U23812 (N_23812,N_13479,N_14313);
and U23813 (N_23813,N_15275,N_15234);
xor U23814 (N_23814,N_14366,N_15428);
and U23815 (N_23815,N_14655,N_13506);
and U23816 (N_23816,N_12762,N_15795);
nor U23817 (N_23817,N_16362,N_13911);
nand U23818 (N_23818,N_16176,N_16199);
xnor U23819 (N_23819,N_13923,N_16652);
or U23820 (N_23820,N_14955,N_16840);
nor U23821 (N_23821,N_15171,N_14391);
nor U23822 (N_23822,N_18535,N_17127);
xor U23823 (N_23823,N_17479,N_13918);
or U23824 (N_23824,N_14021,N_16412);
xnor U23825 (N_23825,N_15463,N_13190);
or U23826 (N_23826,N_15955,N_14333);
or U23827 (N_23827,N_18245,N_17332);
or U23828 (N_23828,N_17993,N_17004);
xor U23829 (N_23829,N_14182,N_16697);
and U23830 (N_23830,N_16885,N_14508);
nor U23831 (N_23831,N_16534,N_16372);
and U23832 (N_23832,N_17130,N_13903);
and U23833 (N_23833,N_13106,N_13213);
nand U23834 (N_23834,N_13348,N_12904);
xnor U23835 (N_23835,N_17088,N_17186);
nand U23836 (N_23836,N_13122,N_15855);
xnor U23837 (N_23837,N_15430,N_14456);
and U23838 (N_23838,N_12897,N_13681);
nor U23839 (N_23839,N_16632,N_14083);
xnor U23840 (N_23840,N_15750,N_18042);
or U23841 (N_23841,N_15020,N_18684);
or U23842 (N_23842,N_14226,N_12666);
xor U23843 (N_23843,N_12586,N_13489);
nand U23844 (N_23844,N_17835,N_15652);
nand U23845 (N_23845,N_15474,N_14710);
nand U23846 (N_23846,N_18732,N_13216);
and U23847 (N_23847,N_16699,N_15617);
and U23848 (N_23848,N_16328,N_12748);
and U23849 (N_23849,N_18678,N_15053);
xnor U23850 (N_23850,N_14395,N_12643);
nand U23851 (N_23851,N_15470,N_15091);
nand U23852 (N_23852,N_13461,N_18645);
and U23853 (N_23853,N_16024,N_12615);
or U23854 (N_23854,N_13176,N_14683);
or U23855 (N_23855,N_17557,N_15668);
xor U23856 (N_23856,N_13398,N_18457);
or U23857 (N_23857,N_14412,N_13237);
nor U23858 (N_23858,N_15257,N_17439);
xor U23859 (N_23859,N_18690,N_18331);
or U23860 (N_23860,N_15606,N_14705);
nand U23861 (N_23861,N_17127,N_13310);
nor U23862 (N_23862,N_13061,N_16579);
nand U23863 (N_23863,N_18658,N_13723);
and U23864 (N_23864,N_14359,N_14249);
or U23865 (N_23865,N_15604,N_15095);
nand U23866 (N_23866,N_14811,N_14204);
or U23867 (N_23867,N_17420,N_12751);
and U23868 (N_23868,N_13015,N_14067);
xor U23869 (N_23869,N_15971,N_15041);
or U23870 (N_23870,N_16174,N_12797);
and U23871 (N_23871,N_18183,N_18097);
xor U23872 (N_23872,N_18317,N_14655);
nand U23873 (N_23873,N_17546,N_17355);
or U23874 (N_23874,N_18143,N_13401);
nor U23875 (N_23875,N_17063,N_14628);
nor U23876 (N_23876,N_14800,N_18166);
or U23877 (N_23877,N_17221,N_13085);
nand U23878 (N_23878,N_14363,N_18274);
or U23879 (N_23879,N_14493,N_18191);
nand U23880 (N_23880,N_13620,N_12642);
nand U23881 (N_23881,N_17543,N_15686);
nor U23882 (N_23882,N_14765,N_14120);
and U23883 (N_23883,N_12884,N_16176);
nand U23884 (N_23884,N_13357,N_14766);
or U23885 (N_23885,N_14531,N_14753);
xor U23886 (N_23886,N_13635,N_13738);
xnor U23887 (N_23887,N_18447,N_15877);
nand U23888 (N_23888,N_15138,N_16195);
or U23889 (N_23889,N_15392,N_12957);
xor U23890 (N_23890,N_16451,N_13683);
nor U23891 (N_23891,N_14056,N_18678);
or U23892 (N_23892,N_18458,N_18260);
nor U23893 (N_23893,N_16346,N_13406);
or U23894 (N_23894,N_13823,N_15479);
and U23895 (N_23895,N_17904,N_13775);
nand U23896 (N_23896,N_17615,N_13112);
xnor U23897 (N_23897,N_16416,N_16881);
and U23898 (N_23898,N_16059,N_13598);
nor U23899 (N_23899,N_15516,N_16297);
and U23900 (N_23900,N_12842,N_14260);
and U23901 (N_23901,N_13118,N_18404);
nand U23902 (N_23902,N_13884,N_14118);
xnor U23903 (N_23903,N_14820,N_17298);
and U23904 (N_23904,N_12577,N_18171);
and U23905 (N_23905,N_12938,N_13133);
or U23906 (N_23906,N_17539,N_14382);
or U23907 (N_23907,N_17825,N_18449);
and U23908 (N_23908,N_14983,N_16824);
nand U23909 (N_23909,N_16015,N_13961);
and U23910 (N_23910,N_12844,N_13699);
nand U23911 (N_23911,N_17439,N_14291);
or U23912 (N_23912,N_13039,N_14802);
and U23913 (N_23913,N_18159,N_15458);
or U23914 (N_23914,N_18193,N_13956);
and U23915 (N_23915,N_12963,N_17876);
or U23916 (N_23916,N_14245,N_15024);
or U23917 (N_23917,N_12593,N_14752);
or U23918 (N_23918,N_16382,N_15899);
nand U23919 (N_23919,N_13510,N_15319);
and U23920 (N_23920,N_18407,N_16837);
nor U23921 (N_23921,N_16781,N_15159);
and U23922 (N_23922,N_15837,N_16667);
or U23923 (N_23923,N_15355,N_12651);
xor U23924 (N_23924,N_15993,N_17164);
nor U23925 (N_23925,N_16284,N_15085);
and U23926 (N_23926,N_16502,N_13529);
or U23927 (N_23927,N_17097,N_15311);
nand U23928 (N_23928,N_14596,N_18296);
or U23929 (N_23929,N_13457,N_17909);
and U23930 (N_23930,N_16722,N_13987);
and U23931 (N_23931,N_17145,N_18550);
nand U23932 (N_23932,N_14531,N_14721);
nor U23933 (N_23933,N_13229,N_13465);
nor U23934 (N_23934,N_17980,N_14444);
or U23935 (N_23935,N_17882,N_17635);
or U23936 (N_23936,N_14741,N_13382);
and U23937 (N_23937,N_13573,N_13677);
and U23938 (N_23938,N_16154,N_16854);
nor U23939 (N_23939,N_16147,N_13107);
or U23940 (N_23940,N_16399,N_14959);
xor U23941 (N_23941,N_14161,N_14749);
or U23942 (N_23942,N_12684,N_18399);
or U23943 (N_23943,N_18609,N_16930);
and U23944 (N_23944,N_17833,N_15761);
nand U23945 (N_23945,N_13812,N_13117);
xor U23946 (N_23946,N_12649,N_18498);
nor U23947 (N_23947,N_17233,N_12722);
or U23948 (N_23948,N_17101,N_17958);
xor U23949 (N_23949,N_13166,N_14986);
nand U23950 (N_23950,N_13389,N_16565);
xor U23951 (N_23951,N_17913,N_15544);
xor U23952 (N_23952,N_15888,N_17765);
or U23953 (N_23953,N_17057,N_17568);
nor U23954 (N_23954,N_16239,N_15416);
nand U23955 (N_23955,N_14522,N_13403);
xor U23956 (N_23956,N_13317,N_12631);
nand U23957 (N_23957,N_15141,N_14410);
and U23958 (N_23958,N_15659,N_14243);
and U23959 (N_23959,N_17612,N_16018);
and U23960 (N_23960,N_13289,N_12673);
nand U23961 (N_23961,N_13955,N_18342);
or U23962 (N_23962,N_15312,N_17821);
nor U23963 (N_23963,N_17046,N_18302);
and U23964 (N_23964,N_16169,N_14426);
nor U23965 (N_23965,N_18249,N_13557);
xnor U23966 (N_23966,N_16206,N_12959);
and U23967 (N_23967,N_16699,N_14001);
nand U23968 (N_23968,N_18472,N_14662);
nor U23969 (N_23969,N_17335,N_13434);
or U23970 (N_23970,N_17976,N_16862);
xnor U23971 (N_23971,N_15209,N_15627);
or U23972 (N_23972,N_16187,N_15949);
xnor U23973 (N_23973,N_12702,N_16996);
and U23974 (N_23974,N_15071,N_18440);
nand U23975 (N_23975,N_17063,N_13673);
nor U23976 (N_23976,N_15748,N_17392);
nor U23977 (N_23977,N_14578,N_14369);
nor U23978 (N_23978,N_12931,N_14930);
xnor U23979 (N_23979,N_16339,N_14766);
or U23980 (N_23980,N_18274,N_16822);
nand U23981 (N_23981,N_15280,N_17362);
or U23982 (N_23982,N_15291,N_15060);
nor U23983 (N_23983,N_16482,N_15102);
or U23984 (N_23984,N_12670,N_17874);
xor U23985 (N_23985,N_12660,N_17745);
and U23986 (N_23986,N_13042,N_14115);
nor U23987 (N_23987,N_17868,N_14686);
xnor U23988 (N_23988,N_17917,N_15421);
or U23989 (N_23989,N_14980,N_15132);
nand U23990 (N_23990,N_12851,N_12512);
or U23991 (N_23991,N_17987,N_12971);
nand U23992 (N_23992,N_12846,N_13605);
nor U23993 (N_23993,N_18458,N_15295);
nor U23994 (N_23994,N_18684,N_12692);
nand U23995 (N_23995,N_17631,N_13441);
nand U23996 (N_23996,N_12710,N_16284);
xnor U23997 (N_23997,N_18083,N_12781);
and U23998 (N_23998,N_16448,N_13655);
nand U23999 (N_23999,N_17802,N_15349);
or U24000 (N_24000,N_18483,N_13586);
or U24001 (N_24001,N_12960,N_15441);
and U24002 (N_24002,N_17325,N_16023);
xnor U24003 (N_24003,N_14968,N_15778);
or U24004 (N_24004,N_13107,N_13261);
nand U24005 (N_24005,N_16687,N_17072);
nand U24006 (N_24006,N_14336,N_15588);
and U24007 (N_24007,N_13304,N_18096);
and U24008 (N_24008,N_14365,N_13872);
xnor U24009 (N_24009,N_17665,N_13721);
nor U24010 (N_24010,N_13285,N_18022);
nand U24011 (N_24011,N_14559,N_17096);
or U24012 (N_24012,N_16834,N_16305);
or U24013 (N_24013,N_18389,N_18078);
and U24014 (N_24014,N_17634,N_16328);
nand U24015 (N_24015,N_16459,N_17210);
xor U24016 (N_24016,N_17977,N_15319);
nand U24017 (N_24017,N_18084,N_13565);
nor U24018 (N_24018,N_16501,N_16927);
nand U24019 (N_24019,N_17074,N_14236);
xnor U24020 (N_24020,N_17528,N_12872);
or U24021 (N_24021,N_14208,N_18426);
nand U24022 (N_24022,N_15049,N_15161);
nor U24023 (N_24023,N_13087,N_15884);
xnor U24024 (N_24024,N_17631,N_17475);
or U24025 (N_24025,N_13081,N_18068);
and U24026 (N_24026,N_13126,N_15782);
nor U24027 (N_24027,N_16619,N_13808);
or U24028 (N_24028,N_15375,N_13916);
xnor U24029 (N_24029,N_14983,N_14785);
nor U24030 (N_24030,N_15870,N_13478);
and U24031 (N_24031,N_16936,N_12758);
nand U24032 (N_24032,N_16492,N_18701);
or U24033 (N_24033,N_16498,N_14074);
nor U24034 (N_24034,N_14996,N_14917);
or U24035 (N_24035,N_15725,N_17970);
nand U24036 (N_24036,N_13767,N_17464);
nor U24037 (N_24037,N_16587,N_14646);
or U24038 (N_24038,N_14304,N_18533);
nor U24039 (N_24039,N_13811,N_15149);
nand U24040 (N_24040,N_18413,N_17807);
and U24041 (N_24041,N_16867,N_15578);
xnor U24042 (N_24042,N_18054,N_14134);
and U24043 (N_24043,N_17161,N_18283);
xnor U24044 (N_24044,N_17240,N_15385);
nor U24045 (N_24045,N_17902,N_14572);
xor U24046 (N_24046,N_15102,N_15242);
or U24047 (N_24047,N_15830,N_16825);
xnor U24048 (N_24048,N_13659,N_12897);
nor U24049 (N_24049,N_13017,N_18616);
xor U24050 (N_24050,N_16894,N_16210);
and U24051 (N_24051,N_16783,N_15617);
or U24052 (N_24052,N_18279,N_18669);
nor U24053 (N_24053,N_14990,N_15756);
or U24054 (N_24054,N_13118,N_14516);
nor U24055 (N_24055,N_18289,N_16908);
xor U24056 (N_24056,N_12745,N_15013);
and U24057 (N_24057,N_15538,N_13321);
nor U24058 (N_24058,N_16831,N_14659);
or U24059 (N_24059,N_14708,N_13379);
or U24060 (N_24060,N_12679,N_17625);
and U24061 (N_24061,N_18257,N_18049);
nand U24062 (N_24062,N_13597,N_15491);
or U24063 (N_24063,N_18195,N_12936);
or U24064 (N_24064,N_16266,N_14305);
and U24065 (N_24065,N_15217,N_17410);
xnor U24066 (N_24066,N_13127,N_17154);
xnor U24067 (N_24067,N_14337,N_12513);
nand U24068 (N_24068,N_13061,N_14730);
nor U24069 (N_24069,N_12958,N_15473);
xor U24070 (N_24070,N_14558,N_14156);
xor U24071 (N_24071,N_17150,N_16259);
xor U24072 (N_24072,N_17484,N_13369);
and U24073 (N_24073,N_15746,N_17018);
or U24074 (N_24074,N_16890,N_17528);
and U24075 (N_24075,N_13378,N_18389);
xnor U24076 (N_24076,N_12976,N_16021);
nand U24077 (N_24077,N_14028,N_17110);
or U24078 (N_24078,N_14657,N_16698);
xnor U24079 (N_24079,N_17730,N_18488);
nand U24080 (N_24080,N_12930,N_13014);
or U24081 (N_24081,N_14115,N_15225);
and U24082 (N_24082,N_17595,N_13762);
nand U24083 (N_24083,N_16089,N_13941);
xor U24084 (N_24084,N_16007,N_15511);
xor U24085 (N_24085,N_12677,N_13963);
xor U24086 (N_24086,N_16480,N_15819);
xor U24087 (N_24087,N_13994,N_13057);
nor U24088 (N_24088,N_14894,N_13594);
xor U24089 (N_24089,N_12900,N_17801);
xor U24090 (N_24090,N_17243,N_13472);
nor U24091 (N_24091,N_17363,N_18478);
or U24092 (N_24092,N_13539,N_14358);
and U24093 (N_24093,N_12608,N_15702);
nor U24094 (N_24094,N_16703,N_14006);
nor U24095 (N_24095,N_18345,N_12662);
and U24096 (N_24096,N_18708,N_13821);
nand U24097 (N_24097,N_18554,N_16215);
xnor U24098 (N_24098,N_18229,N_15800);
xor U24099 (N_24099,N_13312,N_18171);
nand U24100 (N_24100,N_12573,N_16956);
nor U24101 (N_24101,N_14852,N_17394);
xor U24102 (N_24102,N_15621,N_17266);
nor U24103 (N_24103,N_17920,N_12667);
or U24104 (N_24104,N_15079,N_14836);
nor U24105 (N_24105,N_14353,N_13689);
nand U24106 (N_24106,N_16491,N_17441);
or U24107 (N_24107,N_15048,N_18698);
nor U24108 (N_24108,N_17436,N_18098);
xor U24109 (N_24109,N_18647,N_14190);
and U24110 (N_24110,N_13115,N_15888);
nand U24111 (N_24111,N_14847,N_17234);
xnor U24112 (N_24112,N_18404,N_13174);
nor U24113 (N_24113,N_14911,N_16134);
nand U24114 (N_24114,N_17297,N_13151);
nor U24115 (N_24115,N_13546,N_16418);
and U24116 (N_24116,N_14817,N_14803);
and U24117 (N_24117,N_14922,N_13270);
xnor U24118 (N_24118,N_12972,N_15145);
nor U24119 (N_24119,N_13187,N_18005);
nand U24120 (N_24120,N_15753,N_15849);
nor U24121 (N_24121,N_13275,N_13085);
and U24122 (N_24122,N_13775,N_14178);
nor U24123 (N_24123,N_15932,N_14125);
xnor U24124 (N_24124,N_16105,N_16062);
or U24125 (N_24125,N_15265,N_15781);
or U24126 (N_24126,N_18625,N_17453);
xor U24127 (N_24127,N_15296,N_17409);
xor U24128 (N_24128,N_15541,N_14192);
and U24129 (N_24129,N_13340,N_17669);
nand U24130 (N_24130,N_18300,N_13784);
nor U24131 (N_24131,N_18728,N_15140);
xnor U24132 (N_24132,N_14431,N_12658);
and U24133 (N_24133,N_13667,N_18013);
xor U24134 (N_24134,N_14249,N_15222);
or U24135 (N_24135,N_18278,N_18685);
xor U24136 (N_24136,N_13858,N_12751);
or U24137 (N_24137,N_16670,N_15222);
nand U24138 (N_24138,N_13154,N_12643);
xor U24139 (N_24139,N_18638,N_13095);
nand U24140 (N_24140,N_16892,N_12694);
xnor U24141 (N_24141,N_13277,N_18198);
or U24142 (N_24142,N_13808,N_14962);
xor U24143 (N_24143,N_18498,N_16873);
and U24144 (N_24144,N_18080,N_14147);
and U24145 (N_24145,N_16037,N_16057);
nor U24146 (N_24146,N_15648,N_13242);
nand U24147 (N_24147,N_12647,N_15123);
or U24148 (N_24148,N_16163,N_13822);
xnor U24149 (N_24149,N_15397,N_12734);
nand U24150 (N_24150,N_12987,N_18066);
xnor U24151 (N_24151,N_16937,N_17822);
nand U24152 (N_24152,N_18170,N_15013);
nand U24153 (N_24153,N_13856,N_17524);
and U24154 (N_24154,N_16109,N_16135);
or U24155 (N_24155,N_14698,N_14715);
xnor U24156 (N_24156,N_17850,N_16085);
or U24157 (N_24157,N_14408,N_14568);
xor U24158 (N_24158,N_14083,N_14794);
and U24159 (N_24159,N_17971,N_18485);
or U24160 (N_24160,N_15329,N_12770);
xor U24161 (N_24161,N_13595,N_18375);
nor U24162 (N_24162,N_16047,N_12931);
xnor U24163 (N_24163,N_15459,N_16352);
or U24164 (N_24164,N_15684,N_16129);
xor U24165 (N_24165,N_13293,N_15199);
and U24166 (N_24166,N_13749,N_17098);
or U24167 (N_24167,N_17095,N_13923);
nor U24168 (N_24168,N_17981,N_18132);
nand U24169 (N_24169,N_15685,N_13204);
nor U24170 (N_24170,N_14089,N_17226);
nor U24171 (N_24171,N_13950,N_16029);
nand U24172 (N_24172,N_14997,N_18141);
and U24173 (N_24173,N_18011,N_15330);
or U24174 (N_24174,N_17851,N_12785);
nand U24175 (N_24175,N_13532,N_16474);
and U24176 (N_24176,N_17613,N_14701);
xor U24177 (N_24177,N_17619,N_13412);
xor U24178 (N_24178,N_14081,N_17109);
nand U24179 (N_24179,N_15930,N_17083);
and U24180 (N_24180,N_16529,N_15450);
nand U24181 (N_24181,N_18620,N_16241);
nand U24182 (N_24182,N_12651,N_14894);
or U24183 (N_24183,N_14114,N_17857);
nand U24184 (N_24184,N_17016,N_12847);
nand U24185 (N_24185,N_13518,N_14063);
nor U24186 (N_24186,N_17605,N_13551);
or U24187 (N_24187,N_16302,N_14198);
nor U24188 (N_24188,N_17717,N_13175);
nor U24189 (N_24189,N_17378,N_15550);
nor U24190 (N_24190,N_13295,N_15072);
or U24191 (N_24191,N_16942,N_14421);
or U24192 (N_24192,N_15575,N_12947);
nand U24193 (N_24193,N_15729,N_16541);
nand U24194 (N_24194,N_12980,N_15044);
or U24195 (N_24195,N_17081,N_18168);
nor U24196 (N_24196,N_14647,N_18623);
or U24197 (N_24197,N_14298,N_18646);
nand U24198 (N_24198,N_15201,N_12981);
and U24199 (N_24199,N_15535,N_16517);
nor U24200 (N_24200,N_17115,N_15982);
or U24201 (N_24201,N_14289,N_15825);
nand U24202 (N_24202,N_15542,N_16608);
nand U24203 (N_24203,N_13425,N_15098);
and U24204 (N_24204,N_14052,N_14627);
xor U24205 (N_24205,N_15965,N_12802);
xor U24206 (N_24206,N_16406,N_16326);
or U24207 (N_24207,N_15533,N_15355);
nand U24208 (N_24208,N_17492,N_15359);
nor U24209 (N_24209,N_15884,N_16632);
and U24210 (N_24210,N_12538,N_17881);
nand U24211 (N_24211,N_17824,N_13307);
and U24212 (N_24212,N_15393,N_15866);
and U24213 (N_24213,N_15402,N_13922);
xnor U24214 (N_24214,N_15099,N_17169);
nor U24215 (N_24215,N_14677,N_16637);
or U24216 (N_24216,N_16040,N_14268);
or U24217 (N_24217,N_12587,N_13102);
xnor U24218 (N_24218,N_16486,N_15067);
and U24219 (N_24219,N_18069,N_13250);
nor U24220 (N_24220,N_16995,N_13066);
or U24221 (N_24221,N_14892,N_18644);
and U24222 (N_24222,N_14177,N_17909);
nor U24223 (N_24223,N_17874,N_17556);
nor U24224 (N_24224,N_17729,N_17890);
xnor U24225 (N_24225,N_14921,N_15905);
or U24226 (N_24226,N_17156,N_13588);
nand U24227 (N_24227,N_16809,N_16162);
and U24228 (N_24228,N_14984,N_18647);
nor U24229 (N_24229,N_16358,N_14858);
nor U24230 (N_24230,N_15209,N_15108);
nand U24231 (N_24231,N_17628,N_17704);
xor U24232 (N_24232,N_14141,N_18358);
or U24233 (N_24233,N_13335,N_18159);
xor U24234 (N_24234,N_14470,N_14711);
nor U24235 (N_24235,N_15605,N_14906);
xor U24236 (N_24236,N_13495,N_13087);
and U24237 (N_24237,N_14935,N_13332);
nor U24238 (N_24238,N_18571,N_16650);
nor U24239 (N_24239,N_16884,N_18096);
xor U24240 (N_24240,N_18292,N_16091);
or U24241 (N_24241,N_14859,N_15141);
nor U24242 (N_24242,N_14445,N_13529);
xnor U24243 (N_24243,N_14412,N_18109);
nand U24244 (N_24244,N_13064,N_14421);
nor U24245 (N_24245,N_14422,N_15601);
and U24246 (N_24246,N_16223,N_13309);
and U24247 (N_24247,N_13482,N_16888);
nand U24248 (N_24248,N_18412,N_13104);
nand U24249 (N_24249,N_13704,N_14412);
xor U24250 (N_24250,N_15345,N_12654);
nor U24251 (N_24251,N_16139,N_15702);
nor U24252 (N_24252,N_12600,N_16816);
nand U24253 (N_24253,N_18365,N_15735);
xnor U24254 (N_24254,N_13426,N_13863);
and U24255 (N_24255,N_17144,N_13450);
nor U24256 (N_24256,N_18660,N_12553);
nor U24257 (N_24257,N_12813,N_14947);
nor U24258 (N_24258,N_15403,N_13982);
nor U24259 (N_24259,N_15392,N_16022);
or U24260 (N_24260,N_13892,N_16983);
xor U24261 (N_24261,N_17692,N_15774);
xor U24262 (N_24262,N_16146,N_14461);
and U24263 (N_24263,N_13827,N_15177);
xor U24264 (N_24264,N_13793,N_13734);
or U24265 (N_24265,N_13630,N_17494);
or U24266 (N_24266,N_12775,N_18457);
xnor U24267 (N_24267,N_16480,N_16722);
xnor U24268 (N_24268,N_13419,N_12724);
or U24269 (N_24269,N_16959,N_14399);
xnor U24270 (N_24270,N_15192,N_13969);
and U24271 (N_24271,N_14832,N_18423);
and U24272 (N_24272,N_17298,N_17559);
nand U24273 (N_24273,N_12529,N_18653);
nor U24274 (N_24274,N_15618,N_17949);
nand U24275 (N_24275,N_17599,N_14899);
nand U24276 (N_24276,N_17519,N_14697);
nor U24277 (N_24277,N_12632,N_17129);
xor U24278 (N_24278,N_13122,N_14801);
nor U24279 (N_24279,N_17181,N_15388);
or U24280 (N_24280,N_13861,N_13303);
nor U24281 (N_24281,N_18599,N_17475);
nand U24282 (N_24282,N_16990,N_13933);
xor U24283 (N_24283,N_13721,N_16720);
xor U24284 (N_24284,N_15690,N_15691);
xnor U24285 (N_24285,N_15096,N_16148);
nand U24286 (N_24286,N_17879,N_16002);
xnor U24287 (N_24287,N_16470,N_16622);
xor U24288 (N_24288,N_15349,N_17813);
xnor U24289 (N_24289,N_15369,N_12827);
and U24290 (N_24290,N_12505,N_15973);
nand U24291 (N_24291,N_16626,N_15700);
xnor U24292 (N_24292,N_15427,N_16537);
and U24293 (N_24293,N_17953,N_17120);
nor U24294 (N_24294,N_13639,N_14628);
nand U24295 (N_24295,N_15361,N_18370);
or U24296 (N_24296,N_14258,N_18315);
and U24297 (N_24297,N_13316,N_12870);
and U24298 (N_24298,N_17340,N_15542);
xnor U24299 (N_24299,N_18563,N_15223);
and U24300 (N_24300,N_17941,N_16260);
nor U24301 (N_24301,N_14406,N_13092);
nand U24302 (N_24302,N_14435,N_18275);
or U24303 (N_24303,N_16803,N_16542);
nand U24304 (N_24304,N_17296,N_14529);
or U24305 (N_24305,N_12691,N_14611);
or U24306 (N_24306,N_17995,N_18384);
nor U24307 (N_24307,N_14189,N_16157);
or U24308 (N_24308,N_15481,N_18359);
or U24309 (N_24309,N_15653,N_13945);
nor U24310 (N_24310,N_13541,N_15288);
or U24311 (N_24311,N_16942,N_16387);
and U24312 (N_24312,N_18034,N_18313);
or U24313 (N_24313,N_16925,N_14568);
xnor U24314 (N_24314,N_18364,N_17512);
nand U24315 (N_24315,N_18682,N_13507);
or U24316 (N_24316,N_14029,N_18150);
nand U24317 (N_24317,N_13255,N_13349);
nand U24318 (N_24318,N_18174,N_14069);
nand U24319 (N_24319,N_15517,N_15409);
nor U24320 (N_24320,N_14562,N_16624);
or U24321 (N_24321,N_12960,N_13096);
nor U24322 (N_24322,N_16246,N_13836);
and U24323 (N_24323,N_13727,N_12580);
and U24324 (N_24324,N_16634,N_16211);
nand U24325 (N_24325,N_17165,N_15250);
or U24326 (N_24326,N_14151,N_18256);
xnor U24327 (N_24327,N_12685,N_14888);
xnor U24328 (N_24328,N_12558,N_17056);
nor U24329 (N_24329,N_14295,N_14928);
or U24330 (N_24330,N_14717,N_14634);
nand U24331 (N_24331,N_14071,N_13143);
xnor U24332 (N_24332,N_12504,N_18415);
nand U24333 (N_24333,N_16430,N_16148);
nand U24334 (N_24334,N_15250,N_16962);
or U24335 (N_24335,N_16665,N_15310);
xor U24336 (N_24336,N_17992,N_12996);
or U24337 (N_24337,N_16558,N_17754);
or U24338 (N_24338,N_15755,N_12669);
or U24339 (N_24339,N_16207,N_15440);
nand U24340 (N_24340,N_16841,N_15906);
or U24341 (N_24341,N_15130,N_13419);
or U24342 (N_24342,N_17400,N_13822);
or U24343 (N_24343,N_13377,N_13565);
xnor U24344 (N_24344,N_14595,N_16698);
nand U24345 (N_24345,N_12968,N_13337);
xor U24346 (N_24346,N_16485,N_12882);
nor U24347 (N_24347,N_14340,N_15105);
nand U24348 (N_24348,N_15981,N_15741);
and U24349 (N_24349,N_16503,N_13695);
nand U24350 (N_24350,N_13609,N_14614);
or U24351 (N_24351,N_17978,N_15044);
and U24352 (N_24352,N_15965,N_16789);
and U24353 (N_24353,N_17390,N_15085);
xnor U24354 (N_24354,N_17872,N_17991);
nand U24355 (N_24355,N_15449,N_15062);
xor U24356 (N_24356,N_17775,N_13397);
xor U24357 (N_24357,N_13933,N_17280);
xor U24358 (N_24358,N_15069,N_13388);
and U24359 (N_24359,N_16813,N_14806);
nor U24360 (N_24360,N_16080,N_14749);
nor U24361 (N_24361,N_15651,N_17323);
xnor U24362 (N_24362,N_12645,N_12710);
xnor U24363 (N_24363,N_14077,N_17400);
and U24364 (N_24364,N_14897,N_16434);
xor U24365 (N_24365,N_13963,N_17231);
nor U24366 (N_24366,N_15217,N_13344);
nor U24367 (N_24367,N_13344,N_14712);
and U24368 (N_24368,N_17315,N_17730);
or U24369 (N_24369,N_16270,N_13821);
nor U24370 (N_24370,N_12899,N_13124);
and U24371 (N_24371,N_14950,N_18463);
and U24372 (N_24372,N_14603,N_14656);
nand U24373 (N_24373,N_16457,N_18263);
nand U24374 (N_24374,N_17541,N_14650);
nor U24375 (N_24375,N_15306,N_13480);
xnor U24376 (N_24376,N_18542,N_15397);
or U24377 (N_24377,N_12960,N_15288);
or U24378 (N_24378,N_16674,N_14577);
or U24379 (N_24379,N_14364,N_16537);
xor U24380 (N_24380,N_18042,N_13164);
and U24381 (N_24381,N_15833,N_17228);
and U24382 (N_24382,N_13293,N_17860);
and U24383 (N_24383,N_12590,N_17777);
nand U24384 (N_24384,N_18515,N_17293);
nor U24385 (N_24385,N_17865,N_17496);
or U24386 (N_24386,N_17858,N_16507);
and U24387 (N_24387,N_13201,N_16450);
nand U24388 (N_24388,N_17591,N_12644);
xor U24389 (N_24389,N_13365,N_17062);
xnor U24390 (N_24390,N_17637,N_13622);
xnor U24391 (N_24391,N_17777,N_12744);
xor U24392 (N_24392,N_18231,N_15939);
nor U24393 (N_24393,N_12995,N_16132);
nand U24394 (N_24394,N_18548,N_15996);
or U24395 (N_24395,N_13715,N_18107);
xnor U24396 (N_24396,N_14607,N_13809);
nor U24397 (N_24397,N_17652,N_18070);
and U24398 (N_24398,N_18210,N_18059);
or U24399 (N_24399,N_13054,N_13381);
xnor U24400 (N_24400,N_12657,N_18562);
nand U24401 (N_24401,N_13415,N_17431);
and U24402 (N_24402,N_16765,N_17122);
and U24403 (N_24403,N_17101,N_14887);
nor U24404 (N_24404,N_16003,N_18179);
xor U24405 (N_24405,N_14463,N_18035);
or U24406 (N_24406,N_13564,N_17514);
or U24407 (N_24407,N_18706,N_18711);
or U24408 (N_24408,N_17238,N_16723);
nand U24409 (N_24409,N_16109,N_16040);
xor U24410 (N_24410,N_17472,N_16239);
xnor U24411 (N_24411,N_15548,N_16628);
or U24412 (N_24412,N_15857,N_12885);
and U24413 (N_24413,N_17023,N_17779);
nand U24414 (N_24414,N_15315,N_17585);
and U24415 (N_24415,N_17093,N_13287);
or U24416 (N_24416,N_17631,N_14681);
or U24417 (N_24417,N_14825,N_18645);
or U24418 (N_24418,N_15762,N_17943);
xnor U24419 (N_24419,N_14397,N_16383);
nand U24420 (N_24420,N_14537,N_13855);
and U24421 (N_24421,N_18678,N_13064);
or U24422 (N_24422,N_16880,N_13826);
and U24423 (N_24423,N_13638,N_13724);
and U24424 (N_24424,N_14187,N_13554);
or U24425 (N_24425,N_18235,N_13690);
and U24426 (N_24426,N_15338,N_15698);
nor U24427 (N_24427,N_13373,N_16811);
xor U24428 (N_24428,N_12704,N_16481);
or U24429 (N_24429,N_17157,N_12771);
nor U24430 (N_24430,N_17731,N_13458);
or U24431 (N_24431,N_13695,N_17119);
or U24432 (N_24432,N_18746,N_16495);
nand U24433 (N_24433,N_12789,N_15569);
nand U24434 (N_24434,N_13365,N_16871);
nor U24435 (N_24435,N_17080,N_12564);
or U24436 (N_24436,N_17014,N_14113);
xnor U24437 (N_24437,N_18602,N_13633);
nor U24438 (N_24438,N_18705,N_13669);
and U24439 (N_24439,N_13370,N_15091);
xor U24440 (N_24440,N_16128,N_13957);
xor U24441 (N_24441,N_16888,N_14879);
and U24442 (N_24442,N_16068,N_18490);
xnor U24443 (N_24443,N_16322,N_16332);
xor U24444 (N_24444,N_17183,N_17168);
nand U24445 (N_24445,N_14289,N_17493);
xnor U24446 (N_24446,N_18198,N_17564);
nand U24447 (N_24447,N_18739,N_12760);
nor U24448 (N_24448,N_15835,N_12855);
nor U24449 (N_24449,N_16002,N_14053);
nor U24450 (N_24450,N_17005,N_12758);
nand U24451 (N_24451,N_13857,N_13855);
xor U24452 (N_24452,N_18624,N_12541);
nor U24453 (N_24453,N_13730,N_18648);
xor U24454 (N_24454,N_17784,N_17306);
nand U24455 (N_24455,N_14304,N_17014);
xnor U24456 (N_24456,N_12891,N_14131);
or U24457 (N_24457,N_17585,N_17281);
and U24458 (N_24458,N_13074,N_17978);
nand U24459 (N_24459,N_13417,N_15385);
or U24460 (N_24460,N_18563,N_17494);
nor U24461 (N_24461,N_17608,N_17843);
and U24462 (N_24462,N_15124,N_17000);
or U24463 (N_24463,N_15885,N_16002);
xor U24464 (N_24464,N_15311,N_16088);
xnor U24465 (N_24465,N_13394,N_12851);
xor U24466 (N_24466,N_16468,N_15184);
nor U24467 (N_24467,N_16066,N_14349);
xor U24468 (N_24468,N_17859,N_15492);
nand U24469 (N_24469,N_16963,N_13589);
xnor U24470 (N_24470,N_12909,N_13026);
and U24471 (N_24471,N_18603,N_13281);
nor U24472 (N_24472,N_14284,N_15509);
nand U24473 (N_24473,N_13868,N_16756);
or U24474 (N_24474,N_12587,N_14443);
nor U24475 (N_24475,N_13296,N_15297);
xnor U24476 (N_24476,N_14947,N_13303);
and U24477 (N_24477,N_13866,N_12771);
nor U24478 (N_24478,N_16343,N_13321);
xor U24479 (N_24479,N_14237,N_16384);
or U24480 (N_24480,N_16704,N_14433);
xor U24481 (N_24481,N_16371,N_17294);
xor U24482 (N_24482,N_15546,N_17433);
and U24483 (N_24483,N_15745,N_14533);
xor U24484 (N_24484,N_15873,N_13832);
nand U24485 (N_24485,N_15022,N_14551);
xor U24486 (N_24486,N_13681,N_14650);
xnor U24487 (N_24487,N_15288,N_13192);
nor U24488 (N_24488,N_17889,N_15719);
xor U24489 (N_24489,N_18627,N_16936);
or U24490 (N_24490,N_14374,N_15522);
nand U24491 (N_24491,N_15333,N_14498);
xor U24492 (N_24492,N_15456,N_16675);
nor U24493 (N_24493,N_18444,N_13313);
and U24494 (N_24494,N_18320,N_17008);
xor U24495 (N_24495,N_13806,N_18647);
nor U24496 (N_24496,N_14420,N_17319);
or U24497 (N_24497,N_13202,N_13601);
and U24498 (N_24498,N_13334,N_13775);
nand U24499 (N_24499,N_15322,N_17796);
or U24500 (N_24500,N_16059,N_18060);
nor U24501 (N_24501,N_17785,N_15454);
nand U24502 (N_24502,N_14913,N_13661);
or U24503 (N_24503,N_15775,N_12939);
xnor U24504 (N_24504,N_15932,N_17260);
nand U24505 (N_24505,N_16269,N_13731);
and U24506 (N_24506,N_17073,N_13197);
nand U24507 (N_24507,N_15091,N_14250);
nor U24508 (N_24508,N_15179,N_14944);
and U24509 (N_24509,N_18600,N_13948);
nor U24510 (N_24510,N_12706,N_15551);
nand U24511 (N_24511,N_14053,N_16879);
and U24512 (N_24512,N_18713,N_12857);
xor U24513 (N_24513,N_16966,N_12747);
xor U24514 (N_24514,N_13181,N_14291);
and U24515 (N_24515,N_12970,N_14930);
xor U24516 (N_24516,N_16843,N_16238);
nor U24517 (N_24517,N_15151,N_14460);
and U24518 (N_24518,N_18029,N_12745);
nand U24519 (N_24519,N_17891,N_16765);
nand U24520 (N_24520,N_15114,N_16237);
nor U24521 (N_24521,N_14325,N_17290);
and U24522 (N_24522,N_12681,N_12590);
nand U24523 (N_24523,N_14283,N_12621);
nand U24524 (N_24524,N_14095,N_16290);
nor U24525 (N_24525,N_18035,N_15447);
nand U24526 (N_24526,N_15250,N_16688);
nor U24527 (N_24527,N_14261,N_13571);
nand U24528 (N_24528,N_14341,N_18542);
and U24529 (N_24529,N_17556,N_15165);
or U24530 (N_24530,N_13683,N_17184);
nand U24531 (N_24531,N_16061,N_12563);
nor U24532 (N_24532,N_14486,N_13580);
nor U24533 (N_24533,N_17240,N_14023);
and U24534 (N_24534,N_17673,N_16333);
nor U24535 (N_24535,N_18322,N_16862);
nand U24536 (N_24536,N_15452,N_16811);
and U24537 (N_24537,N_15843,N_14772);
nand U24538 (N_24538,N_15322,N_17481);
or U24539 (N_24539,N_18371,N_12775);
or U24540 (N_24540,N_14078,N_16754);
or U24541 (N_24541,N_13023,N_13851);
nor U24542 (N_24542,N_16465,N_16088);
nand U24543 (N_24543,N_12938,N_17584);
xnor U24544 (N_24544,N_13989,N_17867);
and U24545 (N_24545,N_14444,N_14189);
or U24546 (N_24546,N_14209,N_16226);
and U24547 (N_24547,N_15054,N_13494);
nand U24548 (N_24548,N_17985,N_15872);
xor U24549 (N_24549,N_14686,N_18482);
nor U24550 (N_24550,N_17543,N_14666);
and U24551 (N_24551,N_18675,N_15393);
nand U24552 (N_24552,N_12524,N_13975);
xnor U24553 (N_24553,N_14776,N_16294);
xor U24554 (N_24554,N_12839,N_13039);
or U24555 (N_24555,N_16000,N_13615);
and U24556 (N_24556,N_16422,N_15606);
nor U24557 (N_24557,N_13581,N_14069);
nand U24558 (N_24558,N_12962,N_17289);
nor U24559 (N_24559,N_14357,N_17321);
nor U24560 (N_24560,N_18070,N_15475);
or U24561 (N_24561,N_16061,N_16915);
nor U24562 (N_24562,N_12657,N_18600);
nor U24563 (N_24563,N_17826,N_17496);
nor U24564 (N_24564,N_14649,N_15462);
xor U24565 (N_24565,N_17577,N_17347);
nand U24566 (N_24566,N_13090,N_18577);
nand U24567 (N_24567,N_16985,N_14407);
nand U24568 (N_24568,N_14773,N_16573);
nand U24569 (N_24569,N_16971,N_17269);
or U24570 (N_24570,N_18152,N_14160);
and U24571 (N_24571,N_15448,N_14602);
xnor U24572 (N_24572,N_16808,N_16275);
nand U24573 (N_24573,N_13913,N_16177);
and U24574 (N_24574,N_16295,N_16770);
nand U24575 (N_24575,N_13452,N_15664);
or U24576 (N_24576,N_15845,N_13534);
and U24577 (N_24577,N_14672,N_12725);
nor U24578 (N_24578,N_14674,N_14476);
nor U24579 (N_24579,N_17959,N_13344);
and U24580 (N_24580,N_13915,N_12832);
xor U24581 (N_24581,N_14292,N_14840);
or U24582 (N_24582,N_16835,N_17849);
or U24583 (N_24583,N_13838,N_13019);
nand U24584 (N_24584,N_12860,N_14758);
nand U24585 (N_24585,N_13171,N_18723);
nor U24586 (N_24586,N_14060,N_17736);
nor U24587 (N_24587,N_18484,N_15039);
and U24588 (N_24588,N_16446,N_14107);
nand U24589 (N_24589,N_16459,N_17587);
nor U24590 (N_24590,N_17993,N_14572);
nand U24591 (N_24591,N_13116,N_15354);
nor U24592 (N_24592,N_14559,N_16591);
or U24593 (N_24593,N_18166,N_18450);
or U24594 (N_24594,N_14449,N_17560);
and U24595 (N_24595,N_16414,N_17592);
nand U24596 (N_24596,N_18641,N_16108);
nor U24597 (N_24597,N_13034,N_13845);
nor U24598 (N_24598,N_13257,N_17901);
nand U24599 (N_24599,N_12575,N_18186);
and U24600 (N_24600,N_12994,N_13317);
or U24601 (N_24601,N_14697,N_18445);
and U24602 (N_24602,N_14416,N_18696);
or U24603 (N_24603,N_18683,N_16628);
and U24604 (N_24604,N_18378,N_13345);
xor U24605 (N_24605,N_15467,N_12569);
and U24606 (N_24606,N_15639,N_17904);
or U24607 (N_24607,N_15930,N_17263);
nand U24608 (N_24608,N_14824,N_12621);
and U24609 (N_24609,N_12839,N_17032);
or U24610 (N_24610,N_18253,N_18128);
and U24611 (N_24611,N_15263,N_18485);
xnor U24612 (N_24612,N_13771,N_15988);
or U24613 (N_24613,N_16129,N_18346);
and U24614 (N_24614,N_14701,N_15117);
or U24615 (N_24615,N_14072,N_13463);
xnor U24616 (N_24616,N_17049,N_17721);
xnor U24617 (N_24617,N_16942,N_13771);
xnor U24618 (N_24618,N_14369,N_15561);
nor U24619 (N_24619,N_13326,N_14980);
and U24620 (N_24620,N_12718,N_16706);
and U24621 (N_24621,N_18715,N_12849);
nor U24622 (N_24622,N_12827,N_14851);
and U24623 (N_24623,N_15698,N_14353);
and U24624 (N_24624,N_16331,N_18696);
nor U24625 (N_24625,N_14311,N_13028);
nand U24626 (N_24626,N_14820,N_15711);
or U24627 (N_24627,N_15232,N_17778);
and U24628 (N_24628,N_17830,N_16529);
nand U24629 (N_24629,N_17197,N_14101);
nor U24630 (N_24630,N_17061,N_15692);
and U24631 (N_24631,N_12754,N_14298);
nor U24632 (N_24632,N_13058,N_14031);
xor U24633 (N_24633,N_18473,N_12601);
xor U24634 (N_24634,N_14686,N_16965);
nand U24635 (N_24635,N_13885,N_14407);
nand U24636 (N_24636,N_15297,N_14185);
nor U24637 (N_24637,N_16604,N_16423);
nand U24638 (N_24638,N_17956,N_17766);
nor U24639 (N_24639,N_17281,N_12653);
or U24640 (N_24640,N_13309,N_15604);
nor U24641 (N_24641,N_14582,N_18003);
xor U24642 (N_24642,N_16735,N_13583);
and U24643 (N_24643,N_14476,N_13143);
nand U24644 (N_24644,N_16780,N_14544);
xnor U24645 (N_24645,N_14122,N_14783);
nor U24646 (N_24646,N_18185,N_17023);
nand U24647 (N_24647,N_16261,N_18520);
and U24648 (N_24648,N_14740,N_12548);
nor U24649 (N_24649,N_15853,N_13952);
nand U24650 (N_24650,N_14267,N_16825);
nand U24651 (N_24651,N_15582,N_15141);
xnor U24652 (N_24652,N_13042,N_17256);
nand U24653 (N_24653,N_13572,N_15057);
or U24654 (N_24654,N_13323,N_17175);
or U24655 (N_24655,N_13197,N_16399);
or U24656 (N_24656,N_12678,N_12526);
or U24657 (N_24657,N_16829,N_15120);
and U24658 (N_24658,N_17202,N_15066);
or U24659 (N_24659,N_15974,N_13706);
nor U24660 (N_24660,N_12860,N_12522);
nand U24661 (N_24661,N_14516,N_18641);
nand U24662 (N_24662,N_15308,N_15409);
nand U24663 (N_24663,N_14832,N_17343);
xnor U24664 (N_24664,N_15895,N_14126);
xor U24665 (N_24665,N_18666,N_17611);
or U24666 (N_24666,N_13328,N_12969);
and U24667 (N_24667,N_15993,N_17616);
and U24668 (N_24668,N_14490,N_18320);
or U24669 (N_24669,N_15314,N_13980);
nor U24670 (N_24670,N_12698,N_17631);
and U24671 (N_24671,N_14249,N_16527);
nor U24672 (N_24672,N_14912,N_13897);
or U24673 (N_24673,N_14367,N_14963);
nand U24674 (N_24674,N_15497,N_18164);
and U24675 (N_24675,N_13301,N_14895);
and U24676 (N_24676,N_18538,N_12659);
xnor U24677 (N_24677,N_16651,N_13824);
or U24678 (N_24678,N_16158,N_13023);
nor U24679 (N_24679,N_17521,N_12509);
or U24680 (N_24680,N_15156,N_16906);
nand U24681 (N_24681,N_15493,N_17296);
nand U24682 (N_24682,N_15472,N_18745);
nor U24683 (N_24683,N_13933,N_16607);
nand U24684 (N_24684,N_18306,N_13315);
nor U24685 (N_24685,N_13191,N_15285);
xor U24686 (N_24686,N_17196,N_18524);
nand U24687 (N_24687,N_18699,N_16251);
nor U24688 (N_24688,N_14472,N_14991);
or U24689 (N_24689,N_13836,N_17186);
and U24690 (N_24690,N_15399,N_16674);
and U24691 (N_24691,N_18699,N_16263);
nor U24692 (N_24692,N_16805,N_13555);
or U24693 (N_24693,N_18576,N_17567);
or U24694 (N_24694,N_18748,N_12750);
and U24695 (N_24695,N_13921,N_18448);
nand U24696 (N_24696,N_12644,N_18280);
nand U24697 (N_24697,N_14127,N_15274);
and U24698 (N_24698,N_13687,N_13030);
or U24699 (N_24699,N_17962,N_14285);
or U24700 (N_24700,N_16781,N_13616);
or U24701 (N_24701,N_18088,N_13700);
nand U24702 (N_24702,N_16044,N_12519);
or U24703 (N_24703,N_12604,N_13504);
nor U24704 (N_24704,N_12891,N_16763);
nand U24705 (N_24705,N_15873,N_13948);
or U24706 (N_24706,N_14829,N_15176);
or U24707 (N_24707,N_17904,N_14326);
xnor U24708 (N_24708,N_17679,N_13596);
or U24709 (N_24709,N_14566,N_17524);
and U24710 (N_24710,N_18701,N_13118);
nand U24711 (N_24711,N_16643,N_14692);
nor U24712 (N_24712,N_16724,N_15914);
nand U24713 (N_24713,N_15367,N_14365);
nor U24714 (N_24714,N_17469,N_18491);
nor U24715 (N_24715,N_17438,N_14070);
xnor U24716 (N_24716,N_18402,N_13270);
nand U24717 (N_24717,N_14350,N_16673);
xor U24718 (N_24718,N_17477,N_14261);
or U24719 (N_24719,N_17356,N_13593);
or U24720 (N_24720,N_18357,N_18323);
and U24721 (N_24721,N_13907,N_17016);
xor U24722 (N_24722,N_13519,N_14751);
xnor U24723 (N_24723,N_18488,N_15322);
or U24724 (N_24724,N_16983,N_15423);
nand U24725 (N_24725,N_13400,N_12988);
nand U24726 (N_24726,N_13899,N_16001);
nand U24727 (N_24727,N_15655,N_15182);
xor U24728 (N_24728,N_15302,N_14279);
nand U24729 (N_24729,N_15590,N_12599);
xnor U24730 (N_24730,N_16861,N_13014);
or U24731 (N_24731,N_17717,N_12689);
nand U24732 (N_24732,N_14453,N_12586);
xnor U24733 (N_24733,N_14531,N_17687);
xnor U24734 (N_24734,N_17984,N_16860);
or U24735 (N_24735,N_16509,N_16955);
nand U24736 (N_24736,N_14025,N_14374);
nor U24737 (N_24737,N_16613,N_13520);
nand U24738 (N_24738,N_15939,N_13998);
nand U24739 (N_24739,N_14626,N_13289);
xnor U24740 (N_24740,N_15882,N_17034);
nor U24741 (N_24741,N_13112,N_18046);
nor U24742 (N_24742,N_15055,N_15264);
xnor U24743 (N_24743,N_15579,N_14535);
or U24744 (N_24744,N_14602,N_18529);
or U24745 (N_24745,N_15142,N_16346);
xnor U24746 (N_24746,N_12605,N_15488);
and U24747 (N_24747,N_16987,N_17276);
nand U24748 (N_24748,N_15527,N_16296);
xor U24749 (N_24749,N_14228,N_14663);
and U24750 (N_24750,N_18244,N_18604);
or U24751 (N_24751,N_17848,N_18596);
nor U24752 (N_24752,N_14575,N_13220);
xnor U24753 (N_24753,N_16734,N_18457);
and U24754 (N_24754,N_14228,N_18676);
or U24755 (N_24755,N_16598,N_15387);
and U24756 (N_24756,N_16053,N_18733);
nor U24757 (N_24757,N_13150,N_16527);
nand U24758 (N_24758,N_16090,N_12829);
xnor U24759 (N_24759,N_17309,N_15726);
xnor U24760 (N_24760,N_17154,N_13991);
xor U24761 (N_24761,N_17567,N_17940);
nand U24762 (N_24762,N_16300,N_18675);
and U24763 (N_24763,N_14951,N_18327);
nor U24764 (N_24764,N_17457,N_18612);
or U24765 (N_24765,N_17542,N_14795);
xnor U24766 (N_24766,N_17238,N_15182);
nor U24767 (N_24767,N_18477,N_15833);
and U24768 (N_24768,N_15185,N_12703);
or U24769 (N_24769,N_18543,N_17144);
or U24770 (N_24770,N_17507,N_17246);
or U24771 (N_24771,N_18102,N_16569);
or U24772 (N_24772,N_17123,N_14657);
or U24773 (N_24773,N_13557,N_15381);
or U24774 (N_24774,N_15112,N_14895);
or U24775 (N_24775,N_15139,N_13275);
nand U24776 (N_24776,N_18209,N_13441);
nand U24777 (N_24777,N_15714,N_15848);
nand U24778 (N_24778,N_13338,N_18253);
nand U24779 (N_24779,N_13289,N_15825);
or U24780 (N_24780,N_16682,N_14717);
nand U24781 (N_24781,N_13397,N_12644);
nand U24782 (N_24782,N_14601,N_12858);
and U24783 (N_24783,N_18546,N_15289);
nand U24784 (N_24784,N_16170,N_16514);
nor U24785 (N_24785,N_13506,N_17953);
xnor U24786 (N_24786,N_13831,N_14971);
nor U24787 (N_24787,N_14906,N_12549);
or U24788 (N_24788,N_17608,N_17949);
or U24789 (N_24789,N_16159,N_16567);
xnor U24790 (N_24790,N_15368,N_18653);
nor U24791 (N_24791,N_12718,N_13025);
nand U24792 (N_24792,N_15786,N_13836);
nor U24793 (N_24793,N_17972,N_12562);
and U24794 (N_24794,N_12725,N_16556);
or U24795 (N_24795,N_17986,N_17930);
xnor U24796 (N_24796,N_18279,N_12702);
and U24797 (N_24797,N_16546,N_18426);
nor U24798 (N_24798,N_14140,N_13011);
or U24799 (N_24799,N_18524,N_16306);
nand U24800 (N_24800,N_17418,N_13418);
nor U24801 (N_24801,N_14375,N_13885);
and U24802 (N_24802,N_16809,N_18700);
nor U24803 (N_24803,N_15162,N_13879);
nand U24804 (N_24804,N_17163,N_13118);
nor U24805 (N_24805,N_18414,N_16165);
or U24806 (N_24806,N_15489,N_17628);
nor U24807 (N_24807,N_13791,N_17532);
and U24808 (N_24808,N_13542,N_17045);
or U24809 (N_24809,N_15983,N_13335);
xnor U24810 (N_24810,N_18521,N_17235);
xnor U24811 (N_24811,N_17629,N_12666);
nor U24812 (N_24812,N_17516,N_13419);
or U24813 (N_24813,N_17695,N_13693);
nand U24814 (N_24814,N_16361,N_18122);
nor U24815 (N_24815,N_15966,N_13285);
nand U24816 (N_24816,N_18349,N_17385);
nor U24817 (N_24817,N_14453,N_15248);
nor U24818 (N_24818,N_15491,N_15034);
nand U24819 (N_24819,N_17988,N_13658);
or U24820 (N_24820,N_12677,N_13684);
xnor U24821 (N_24821,N_18185,N_13530);
nand U24822 (N_24822,N_16024,N_17266);
and U24823 (N_24823,N_16233,N_17467);
nand U24824 (N_24824,N_17722,N_13135);
and U24825 (N_24825,N_18373,N_15967);
or U24826 (N_24826,N_13572,N_17699);
nand U24827 (N_24827,N_18225,N_13125);
xnor U24828 (N_24828,N_13318,N_17174);
nor U24829 (N_24829,N_13664,N_14033);
or U24830 (N_24830,N_18136,N_13920);
nand U24831 (N_24831,N_17467,N_18538);
xnor U24832 (N_24832,N_13842,N_14630);
or U24833 (N_24833,N_18193,N_12872);
nand U24834 (N_24834,N_17242,N_17023);
nand U24835 (N_24835,N_15109,N_18490);
or U24836 (N_24836,N_18484,N_15118);
or U24837 (N_24837,N_13034,N_14304);
or U24838 (N_24838,N_16886,N_17540);
and U24839 (N_24839,N_15660,N_13556);
nand U24840 (N_24840,N_18130,N_16923);
and U24841 (N_24841,N_14905,N_15475);
or U24842 (N_24842,N_16939,N_18331);
nand U24843 (N_24843,N_17944,N_17266);
nor U24844 (N_24844,N_14050,N_14734);
nor U24845 (N_24845,N_13935,N_14957);
nor U24846 (N_24846,N_13025,N_17811);
or U24847 (N_24847,N_15533,N_12902);
nor U24848 (N_24848,N_15984,N_17148);
nand U24849 (N_24849,N_12774,N_14669);
and U24850 (N_24850,N_15891,N_17663);
nand U24851 (N_24851,N_16832,N_18704);
xor U24852 (N_24852,N_16456,N_17871);
nor U24853 (N_24853,N_13724,N_15271);
xor U24854 (N_24854,N_16604,N_16258);
nand U24855 (N_24855,N_17648,N_17500);
or U24856 (N_24856,N_17033,N_14877);
or U24857 (N_24857,N_15848,N_16558);
xor U24858 (N_24858,N_14921,N_18156);
xnor U24859 (N_24859,N_16073,N_13053);
nand U24860 (N_24860,N_16007,N_15925);
nor U24861 (N_24861,N_13498,N_13658);
and U24862 (N_24862,N_16392,N_17201);
xnor U24863 (N_24863,N_15543,N_14826);
xnor U24864 (N_24864,N_17743,N_16278);
xnor U24865 (N_24865,N_12522,N_15853);
xor U24866 (N_24866,N_16091,N_13522);
and U24867 (N_24867,N_18020,N_13857);
nor U24868 (N_24868,N_18336,N_14537);
and U24869 (N_24869,N_16314,N_13141);
nand U24870 (N_24870,N_16712,N_13510);
and U24871 (N_24871,N_13278,N_18405);
xor U24872 (N_24872,N_17724,N_16503);
or U24873 (N_24873,N_18613,N_13023);
nand U24874 (N_24874,N_15813,N_14793);
or U24875 (N_24875,N_16497,N_15263);
nor U24876 (N_24876,N_15034,N_15690);
nor U24877 (N_24877,N_14196,N_16298);
nand U24878 (N_24878,N_17308,N_12912);
or U24879 (N_24879,N_13829,N_14193);
nor U24880 (N_24880,N_14178,N_18161);
xor U24881 (N_24881,N_13667,N_18412);
or U24882 (N_24882,N_17407,N_18074);
or U24883 (N_24883,N_17576,N_17311);
xor U24884 (N_24884,N_17170,N_12689);
xnor U24885 (N_24885,N_17598,N_14169);
and U24886 (N_24886,N_13579,N_18398);
nand U24887 (N_24887,N_13200,N_18026);
nor U24888 (N_24888,N_17593,N_14350);
and U24889 (N_24889,N_12854,N_13781);
nor U24890 (N_24890,N_17248,N_16879);
and U24891 (N_24891,N_13419,N_13921);
and U24892 (N_24892,N_14822,N_16004);
and U24893 (N_24893,N_18257,N_14226);
nor U24894 (N_24894,N_16824,N_15213);
nor U24895 (N_24895,N_14015,N_18652);
nor U24896 (N_24896,N_15413,N_16393);
and U24897 (N_24897,N_14412,N_14788);
xnor U24898 (N_24898,N_15288,N_15921);
xor U24899 (N_24899,N_15128,N_13673);
nor U24900 (N_24900,N_14709,N_17590);
xor U24901 (N_24901,N_16659,N_12550);
nand U24902 (N_24902,N_14237,N_12894);
or U24903 (N_24903,N_18042,N_16911);
nor U24904 (N_24904,N_17398,N_17493);
and U24905 (N_24905,N_16739,N_14592);
or U24906 (N_24906,N_16848,N_16700);
xnor U24907 (N_24907,N_17197,N_13588);
nor U24908 (N_24908,N_14668,N_15064);
nand U24909 (N_24909,N_13122,N_14481);
and U24910 (N_24910,N_12636,N_16025);
nand U24911 (N_24911,N_13592,N_14784);
nor U24912 (N_24912,N_18688,N_14334);
nand U24913 (N_24913,N_17312,N_12675);
and U24914 (N_24914,N_14371,N_14470);
or U24915 (N_24915,N_15110,N_12636);
or U24916 (N_24916,N_13381,N_12596);
xor U24917 (N_24917,N_17595,N_14734);
or U24918 (N_24918,N_17143,N_14138);
nor U24919 (N_24919,N_15008,N_17097);
and U24920 (N_24920,N_13551,N_14430);
nand U24921 (N_24921,N_16309,N_17797);
or U24922 (N_24922,N_13895,N_16406);
xor U24923 (N_24923,N_14905,N_17602);
xor U24924 (N_24924,N_12672,N_15379);
or U24925 (N_24925,N_13830,N_13136);
or U24926 (N_24926,N_18713,N_13185);
or U24927 (N_24927,N_15488,N_16556);
and U24928 (N_24928,N_13382,N_15101);
nand U24929 (N_24929,N_14393,N_17515);
nor U24930 (N_24930,N_17208,N_16309);
xor U24931 (N_24931,N_16019,N_14774);
or U24932 (N_24932,N_16762,N_16091);
nand U24933 (N_24933,N_14357,N_15808);
or U24934 (N_24934,N_17651,N_15660);
nor U24935 (N_24935,N_14515,N_13583);
xor U24936 (N_24936,N_13600,N_14997);
nand U24937 (N_24937,N_15172,N_13340);
nor U24938 (N_24938,N_13266,N_14398);
or U24939 (N_24939,N_12691,N_13316);
and U24940 (N_24940,N_13213,N_12626);
and U24941 (N_24941,N_13176,N_13374);
xnor U24942 (N_24942,N_17532,N_15048);
xnor U24943 (N_24943,N_14814,N_13873);
xor U24944 (N_24944,N_13865,N_14029);
or U24945 (N_24945,N_17126,N_13414);
or U24946 (N_24946,N_17139,N_17191);
and U24947 (N_24947,N_14595,N_12656);
nand U24948 (N_24948,N_15297,N_17105);
xnor U24949 (N_24949,N_15098,N_13609);
and U24950 (N_24950,N_13879,N_17033);
or U24951 (N_24951,N_14030,N_13034);
or U24952 (N_24952,N_16386,N_14106);
xnor U24953 (N_24953,N_17236,N_15622);
or U24954 (N_24954,N_14475,N_16264);
and U24955 (N_24955,N_12619,N_17015);
nand U24956 (N_24956,N_13920,N_14370);
and U24957 (N_24957,N_13810,N_16926);
or U24958 (N_24958,N_16562,N_18338);
or U24959 (N_24959,N_14222,N_13062);
xnor U24960 (N_24960,N_14305,N_13755);
and U24961 (N_24961,N_16743,N_15366);
nor U24962 (N_24962,N_15074,N_15850);
nor U24963 (N_24963,N_12504,N_14119);
and U24964 (N_24964,N_16179,N_15191);
nor U24965 (N_24965,N_15727,N_16763);
xor U24966 (N_24966,N_14762,N_15793);
xor U24967 (N_24967,N_17431,N_17225);
nor U24968 (N_24968,N_17729,N_13744);
xnor U24969 (N_24969,N_17217,N_17062);
and U24970 (N_24970,N_13823,N_15507);
nand U24971 (N_24971,N_13125,N_13338);
nand U24972 (N_24972,N_14919,N_12875);
nor U24973 (N_24973,N_17837,N_17122);
nand U24974 (N_24974,N_16996,N_15428);
nand U24975 (N_24975,N_15212,N_18243);
nand U24976 (N_24976,N_17087,N_15475);
and U24977 (N_24977,N_18084,N_13421);
nor U24978 (N_24978,N_18733,N_14515);
and U24979 (N_24979,N_18557,N_17260);
nor U24980 (N_24980,N_12840,N_17956);
nor U24981 (N_24981,N_13628,N_18104);
or U24982 (N_24982,N_14819,N_13833);
xnor U24983 (N_24983,N_17146,N_12890);
xnor U24984 (N_24984,N_13109,N_16339);
nor U24985 (N_24985,N_16705,N_15059);
or U24986 (N_24986,N_14428,N_16729);
nand U24987 (N_24987,N_14917,N_14457);
and U24988 (N_24988,N_13382,N_15089);
and U24989 (N_24989,N_14515,N_17918);
xor U24990 (N_24990,N_15434,N_13603);
nand U24991 (N_24991,N_13478,N_16022);
or U24992 (N_24992,N_14870,N_16656);
xor U24993 (N_24993,N_14891,N_16171);
xnor U24994 (N_24994,N_13365,N_13078);
and U24995 (N_24995,N_18425,N_12682);
or U24996 (N_24996,N_12740,N_14754);
nand U24997 (N_24997,N_12916,N_16759);
and U24998 (N_24998,N_13768,N_12671);
nand U24999 (N_24999,N_18206,N_18448);
and UO_0 (O_0,N_19453,N_22345);
xor UO_1 (O_1,N_20337,N_23903);
xnor UO_2 (O_2,N_18798,N_22996);
or UO_3 (O_3,N_22767,N_24563);
nand UO_4 (O_4,N_19491,N_19270);
xnor UO_5 (O_5,N_19442,N_21769);
and UO_6 (O_6,N_19633,N_24557);
xor UO_7 (O_7,N_24853,N_23235);
xor UO_8 (O_8,N_22230,N_22620);
nand UO_9 (O_9,N_20547,N_20861);
and UO_10 (O_10,N_24531,N_22253);
and UO_11 (O_11,N_23265,N_24220);
and UO_12 (O_12,N_21866,N_21756);
xnor UO_13 (O_13,N_19001,N_24455);
nor UO_14 (O_14,N_24325,N_18855);
nor UO_15 (O_15,N_24822,N_23727);
nor UO_16 (O_16,N_19920,N_24834);
nand UO_17 (O_17,N_24634,N_19333);
nor UO_18 (O_18,N_24584,N_20251);
and UO_19 (O_19,N_23674,N_22537);
and UO_20 (O_20,N_24875,N_21146);
and UO_21 (O_21,N_19496,N_19718);
nand UO_22 (O_22,N_24988,N_23454);
and UO_23 (O_23,N_21301,N_24336);
xor UO_24 (O_24,N_22735,N_20959);
and UO_25 (O_25,N_22210,N_24337);
xnor UO_26 (O_26,N_20850,N_24075);
nand UO_27 (O_27,N_24049,N_24029);
nand UO_28 (O_28,N_22698,N_23046);
xor UO_29 (O_29,N_23192,N_19824);
xnor UO_30 (O_30,N_22671,N_22830);
xnor UO_31 (O_31,N_24045,N_19924);
nand UO_32 (O_32,N_24639,N_22902);
xor UO_33 (O_33,N_24258,N_21595);
nor UO_34 (O_34,N_19710,N_21912);
and UO_35 (O_35,N_21350,N_21247);
or UO_36 (O_36,N_18895,N_21919);
nor UO_37 (O_37,N_24462,N_19766);
and UO_38 (O_38,N_21670,N_19683);
nor UO_39 (O_39,N_21940,N_18818);
xor UO_40 (O_40,N_22485,N_20461);
nor UO_41 (O_41,N_19880,N_19087);
xnor UO_42 (O_42,N_18755,N_19897);
nor UO_43 (O_43,N_22019,N_19437);
nor UO_44 (O_44,N_22314,N_18817);
nor UO_45 (O_45,N_21251,N_21693);
xor UO_46 (O_46,N_24957,N_20854);
xor UO_47 (O_47,N_19157,N_20667);
and UO_48 (O_48,N_19999,N_22927);
nand UO_49 (O_49,N_24934,N_19988);
or UO_50 (O_50,N_20605,N_21227);
nand UO_51 (O_51,N_22301,N_18925);
and UO_52 (O_52,N_20834,N_20971);
nor UO_53 (O_53,N_23677,N_20774);
nand UO_54 (O_54,N_20589,N_24637);
and UO_55 (O_55,N_21926,N_20713);
or UO_56 (O_56,N_24299,N_23226);
nand UO_57 (O_57,N_23323,N_22038);
and UO_58 (O_58,N_20211,N_23260);
and UO_59 (O_59,N_22388,N_22484);
nand UO_60 (O_60,N_23813,N_22398);
nor UO_61 (O_61,N_24737,N_24546);
nor UO_62 (O_62,N_21763,N_22150);
and UO_63 (O_63,N_20816,N_18885);
nor UO_64 (O_64,N_22521,N_20577);
xor UO_65 (O_65,N_24688,N_22156);
xnor UO_66 (O_66,N_23380,N_24483);
and UO_67 (O_67,N_21674,N_22960);
nor UO_68 (O_68,N_22407,N_24063);
nor UO_69 (O_69,N_20779,N_20644);
nand UO_70 (O_70,N_21373,N_20927);
xor UO_71 (O_71,N_23304,N_19393);
xnor UO_72 (O_72,N_23015,N_22157);
or UO_73 (O_73,N_20883,N_19737);
nand UO_74 (O_74,N_23305,N_21521);
and UO_75 (O_75,N_21203,N_23966);
xnor UO_76 (O_76,N_20218,N_24799);
or UO_77 (O_77,N_22041,N_21111);
nor UO_78 (O_78,N_19484,N_24361);
and UO_79 (O_79,N_24689,N_18921);
and UO_80 (O_80,N_21526,N_23453);
nand UO_81 (O_81,N_22612,N_20091);
nor UO_82 (O_82,N_23723,N_20098);
nand UO_83 (O_83,N_21596,N_19726);
nor UO_84 (O_84,N_19755,N_20486);
or UO_85 (O_85,N_20729,N_23361);
nor UO_86 (O_86,N_23514,N_21974);
and UO_87 (O_87,N_21436,N_23427);
nor UO_88 (O_88,N_23846,N_22410);
nand UO_89 (O_89,N_20210,N_20941);
nor UO_90 (O_90,N_21392,N_22775);
nand UO_91 (O_91,N_22602,N_24198);
nand UO_92 (O_92,N_19457,N_24260);
xnor UO_93 (O_93,N_20873,N_20466);
and UO_94 (O_94,N_23633,N_19613);
or UO_95 (O_95,N_18830,N_24190);
or UO_96 (O_96,N_21677,N_22932);
xor UO_97 (O_97,N_22514,N_19774);
or UO_98 (O_98,N_23045,N_22616);
and UO_99 (O_99,N_20471,N_22886);
nand UO_100 (O_100,N_24903,N_24250);
nand UO_101 (O_101,N_24982,N_23063);
nor UO_102 (O_102,N_22419,N_22549);
nand UO_103 (O_103,N_20954,N_24293);
nor UO_104 (O_104,N_20165,N_22013);
nor UO_105 (O_105,N_20428,N_19231);
xnor UO_106 (O_106,N_20167,N_19587);
xnor UO_107 (O_107,N_22931,N_22974);
and UO_108 (O_108,N_22732,N_21744);
xor UO_109 (O_109,N_19528,N_18974);
nor UO_110 (O_110,N_23199,N_24393);
nand UO_111 (O_111,N_23049,N_20092);
and UO_112 (O_112,N_21664,N_21802);
nand UO_113 (O_113,N_21405,N_21776);
or UO_114 (O_114,N_23696,N_22141);
nand UO_115 (O_115,N_21126,N_24964);
nor UO_116 (O_116,N_24669,N_24797);
nor UO_117 (O_117,N_20268,N_21532);
and UO_118 (O_118,N_23073,N_22009);
or UO_119 (O_119,N_20451,N_18916);
and UO_120 (O_120,N_20651,N_24241);
nor UO_121 (O_121,N_18757,N_21856);
xnor UO_122 (O_122,N_19301,N_23294);
nor UO_123 (O_123,N_21904,N_21394);
nor UO_124 (O_124,N_22145,N_18891);
xor UO_125 (O_125,N_19638,N_23208);
xnor UO_126 (O_126,N_24864,N_21982);
or UO_127 (O_127,N_20204,N_19636);
nor UO_128 (O_128,N_24774,N_22244);
and UO_129 (O_129,N_24969,N_20159);
xor UO_130 (O_130,N_20701,N_21407);
nor UO_131 (O_131,N_20258,N_22010);
and UO_132 (O_132,N_21470,N_18811);
xnor UO_133 (O_133,N_21001,N_20117);
and UO_134 (O_134,N_19791,N_19062);
or UO_135 (O_135,N_21662,N_21055);
nor UO_136 (O_136,N_19074,N_19730);
nand UO_137 (O_137,N_19521,N_19435);
xor UO_138 (O_138,N_21345,N_23911);
and UO_139 (O_139,N_24363,N_19721);
or UO_140 (O_140,N_21360,N_23409);
and UO_141 (O_141,N_21232,N_24611);
nor UO_142 (O_142,N_21419,N_23341);
or UO_143 (O_143,N_21398,N_24503);
and UO_144 (O_144,N_22466,N_21032);
or UO_145 (O_145,N_22395,N_19973);
or UO_146 (O_146,N_20002,N_24240);
and UO_147 (O_147,N_22770,N_24953);
and UO_148 (O_148,N_19494,N_24463);
nand UO_149 (O_149,N_21481,N_22779);
xnor UO_150 (O_150,N_19653,N_19674);
or UO_151 (O_151,N_24370,N_21796);
nand UO_152 (O_152,N_22976,N_22734);
nor UO_153 (O_153,N_20707,N_22346);
nor UO_154 (O_154,N_21509,N_19332);
nor UO_155 (O_155,N_20588,N_20592);
and UO_156 (O_156,N_21009,N_20988);
nand UO_157 (O_157,N_24847,N_21827);
xnor UO_158 (O_158,N_24811,N_19339);
xnor UO_159 (O_159,N_23850,N_21936);
and UO_160 (O_160,N_20473,N_20570);
xnor UO_161 (O_161,N_24161,N_21819);
nor UO_162 (O_162,N_23624,N_23164);
and UO_163 (O_163,N_23489,N_24769);
and UO_164 (O_164,N_22335,N_24050);
or UO_165 (O_165,N_24789,N_23246);
xnor UO_166 (O_166,N_20297,N_24861);
nand UO_167 (O_167,N_19566,N_23152);
xor UO_168 (O_168,N_19035,N_19517);
or UO_169 (O_169,N_19776,N_24873);
nor UO_170 (O_170,N_22804,N_22105);
nand UO_171 (O_171,N_22656,N_22309);
or UO_172 (O_172,N_20662,N_23729);
xnor UO_173 (O_173,N_24651,N_23993);
and UO_174 (O_174,N_21946,N_21703);
and UO_175 (O_175,N_22796,N_21489);
nand UO_176 (O_176,N_24713,N_20256);
nand UO_177 (O_177,N_19198,N_21543);
or UO_178 (O_178,N_20699,N_19141);
and UO_179 (O_179,N_19129,N_19458);
xnor UO_180 (O_180,N_18982,N_24907);
xor UO_181 (O_181,N_23457,N_23515);
nand UO_182 (O_182,N_23755,N_24730);
nand UO_183 (O_183,N_20311,N_22838);
or UO_184 (O_184,N_20418,N_23103);
nor UO_185 (O_185,N_24910,N_22468);
xor UO_186 (O_186,N_20213,N_24901);
and UO_187 (O_187,N_22972,N_20758);
nand UO_188 (O_188,N_19402,N_23722);
and UO_189 (O_189,N_22686,N_20705);
xor UO_190 (O_190,N_21401,N_20366);
or UO_191 (O_191,N_22845,N_24263);
nor UO_192 (O_192,N_23784,N_22965);
or UO_193 (O_193,N_23408,N_24012);
nand UO_194 (O_194,N_22206,N_20770);
or UO_195 (O_195,N_19773,N_19156);
nor UO_196 (O_196,N_21014,N_19903);
and UO_197 (O_197,N_21655,N_20431);
nor UO_198 (O_198,N_20754,N_22531);
and UO_199 (O_199,N_22077,N_20782);
nand UO_200 (O_200,N_19133,N_19095);
or UO_201 (O_201,N_20944,N_23744);
nand UO_202 (O_202,N_24835,N_24465);
or UO_203 (O_203,N_21039,N_22042);
and UO_204 (O_204,N_22294,N_24351);
or UO_205 (O_205,N_20304,N_24586);
nand UO_206 (O_206,N_22945,N_24279);
nand UO_207 (O_207,N_20090,N_19618);
nand UO_208 (O_208,N_19276,N_24504);
nor UO_209 (O_209,N_20613,N_20684);
nand UO_210 (O_210,N_21808,N_19930);
and UO_211 (O_211,N_21892,N_23626);
and UO_212 (O_212,N_22115,N_20374);
nand UO_213 (O_213,N_22577,N_23259);
nand UO_214 (O_214,N_24272,N_23228);
and UO_215 (O_215,N_19452,N_24083);
xor UO_216 (O_216,N_24410,N_19214);
or UO_217 (O_217,N_21459,N_20261);
nor UO_218 (O_218,N_23950,N_20745);
and UO_219 (O_219,N_24522,N_19306);
or UO_220 (O_220,N_20125,N_18843);
and UO_221 (O_221,N_22919,N_22982);
nor UO_222 (O_222,N_22975,N_21088);
nand UO_223 (O_223,N_20511,N_22034);
nor UO_224 (O_224,N_23030,N_22282);
xor UO_225 (O_225,N_24484,N_21909);
nor UO_226 (O_226,N_23517,N_19697);
or UO_227 (O_227,N_20700,N_20848);
or UO_228 (O_228,N_19530,N_23666);
xor UO_229 (O_229,N_24793,N_23516);
nor UO_230 (O_230,N_21824,N_22625);
and UO_231 (O_231,N_21850,N_24328);
xor UO_232 (O_232,N_24018,N_20717);
or UO_233 (O_233,N_23367,N_19682);
nand UO_234 (O_234,N_21252,N_19196);
and UO_235 (O_235,N_20922,N_20271);
or UO_236 (O_236,N_21905,N_23610);
xor UO_237 (O_237,N_24666,N_19463);
or UO_238 (O_238,N_20783,N_23472);
xor UO_239 (O_239,N_23375,N_20238);
and UO_240 (O_240,N_20171,N_21463);
or UO_241 (O_241,N_23252,N_21632);
xor UO_242 (O_242,N_24461,N_22343);
and UO_243 (O_243,N_22328,N_21991);
nor UO_244 (O_244,N_22432,N_23614);
nand UO_245 (O_245,N_20500,N_22634);
nor UO_246 (O_246,N_20518,N_23686);
xnor UO_247 (O_247,N_23175,N_19298);
or UO_248 (O_248,N_24618,N_22439);
xnor UO_249 (O_249,N_21434,N_19844);
and UO_250 (O_250,N_23845,N_24765);
xnor UO_251 (O_251,N_18950,N_21404);
and UO_252 (O_252,N_24828,N_23940);
nor UO_253 (O_253,N_22883,N_20727);
and UO_254 (O_254,N_20043,N_21626);
xnor UO_255 (O_255,N_19789,N_23658);
nand UO_256 (O_256,N_24001,N_21049);
or UO_257 (O_257,N_19693,N_18874);
nor UO_258 (O_258,N_20763,N_20544);
or UO_259 (O_259,N_21480,N_20893);
nand UO_260 (O_260,N_19412,N_24340);
nand UO_261 (O_261,N_24905,N_20969);
and UO_262 (O_262,N_23053,N_24432);
and UO_263 (O_263,N_20599,N_23358);
xnor UO_264 (O_264,N_19644,N_22578);
nor UO_265 (O_265,N_24918,N_22112);
or UO_266 (O_266,N_23431,N_23593);
xnor UO_267 (O_267,N_19659,N_24549);
and UO_268 (O_268,N_23001,N_19676);
nand UO_269 (O_269,N_19628,N_22292);
nand UO_270 (O_270,N_21250,N_23261);
xor UO_271 (O_271,N_24997,N_23806);
xor UO_272 (O_272,N_21058,N_21229);
and UO_273 (O_273,N_19394,N_19936);
nor UO_274 (O_274,N_21402,N_19868);
xor UO_275 (O_275,N_23012,N_19797);
nor UO_276 (O_276,N_18881,N_23715);
nand UO_277 (O_277,N_24353,N_23079);
or UO_278 (O_278,N_24927,N_24207);
and UO_279 (O_279,N_18839,N_21957);
nor UO_280 (O_280,N_18954,N_21200);
nor UO_281 (O_281,N_21233,N_24124);
nor UO_282 (O_282,N_19976,N_24216);
xor UO_283 (O_283,N_23708,N_21018);
or UO_284 (O_284,N_22757,N_18952);
nand UO_285 (O_285,N_20665,N_22237);
xnor UO_286 (O_286,N_24696,N_19863);
nand UO_287 (O_287,N_22753,N_22682);
xnor UO_288 (O_288,N_23823,N_20572);
or UO_289 (O_289,N_22662,N_18825);
nor UO_290 (O_290,N_23041,N_20409);
and UO_291 (O_291,N_23299,N_20618);
nand UO_292 (O_292,N_21895,N_22074);
and UO_293 (O_293,N_20842,N_22582);
nand UO_294 (O_294,N_18847,N_22628);
and UO_295 (O_295,N_20637,N_24543);
or UO_296 (O_296,N_19342,N_20643);
and UO_297 (O_297,N_21450,N_20427);
xnor UO_298 (O_298,N_19071,N_20269);
xor UO_299 (O_299,N_20414,N_23527);
nor UO_300 (O_300,N_20382,N_23444);
nor UO_301 (O_301,N_23975,N_24379);
nor UO_302 (O_302,N_21334,N_22385);
xor UO_303 (O_303,N_23086,N_24172);
nor UO_304 (O_304,N_23925,N_22096);
nor UO_305 (O_305,N_21184,N_23748);
nand UO_306 (O_306,N_23440,N_20504);
or UO_307 (O_307,N_24373,N_22502);
nor UO_308 (O_308,N_23741,N_21134);
and UO_309 (O_309,N_19706,N_21370);
and UO_310 (O_310,N_21965,N_19830);
xnor UO_311 (O_311,N_23313,N_21574);
xnor UO_312 (O_312,N_21682,N_21217);
and UO_313 (O_313,N_18775,N_19550);
and UO_314 (O_314,N_22386,N_22673);
or UO_315 (O_315,N_20812,N_20935);
nand UO_316 (O_316,N_23652,N_19963);
and UO_317 (O_317,N_19687,N_18863);
xor UO_318 (O_318,N_20747,N_21514);
and UO_319 (O_319,N_21613,N_23526);
and UO_320 (O_320,N_22725,N_20048);
and UO_321 (O_321,N_23097,N_23205);
and UO_322 (O_322,N_20458,N_22261);
nand UO_323 (O_323,N_20849,N_21412);
nand UO_324 (O_324,N_22259,N_19689);
nand UO_325 (O_325,N_24398,N_23118);
or UO_326 (O_326,N_22833,N_23819);
nor UO_327 (O_327,N_24675,N_22469);
or UO_328 (O_328,N_23155,N_19312);
and UO_329 (O_329,N_20233,N_21133);
nand UO_330 (O_330,N_19227,N_22006);
and UO_331 (O_331,N_20005,N_22704);
and UO_332 (O_332,N_22088,N_22037);
and UO_333 (O_333,N_20021,N_19281);
nand UO_334 (O_334,N_21860,N_22888);
or UO_335 (O_335,N_24523,N_23370);
nand UO_336 (O_336,N_24805,N_22128);
or UO_337 (O_337,N_22851,N_19349);
or UO_338 (O_338,N_21903,N_22797);
nand UO_339 (O_339,N_20336,N_18983);
xnor UO_340 (O_340,N_24273,N_21935);
xnor UO_341 (O_341,N_23301,N_19405);
nand UO_342 (O_342,N_20906,N_21520);
or UO_343 (O_343,N_23709,N_19049);
and UO_344 (O_344,N_20319,N_22822);
nor UO_345 (O_345,N_23270,N_21578);
nor UO_346 (O_346,N_22563,N_23583);
and UO_347 (O_347,N_19749,N_24959);
nand UO_348 (O_348,N_21076,N_19401);
or UO_349 (O_349,N_19732,N_23297);
nand UO_350 (O_350,N_19576,N_20680);
nor UO_351 (O_351,N_23679,N_19099);
xor UO_352 (O_352,N_22646,N_18927);
xor UO_353 (O_353,N_22046,N_21708);
nor UO_354 (O_354,N_24092,N_24958);
or UO_355 (O_355,N_22270,N_24709);
nand UO_356 (O_356,N_24388,N_19395);
nor UO_357 (O_357,N_24854,N_23601);
nor UO_358 (O_358,N_24107,N_20843);
and UO_359 (O_359,N_24986,N_24101);
xor UO_360 (O_360,N_24118,N_19900);
and UO_361 (O_361,N_22754,N_23498);
nor UO_362 (O_362,N_24719,N_18848);
nand UO_363 (O_363,N_21259,N_18842);
and UO_364 (O_364,N_19450,N_22979);
nor UO_365 (O_365,N_20846,N_19769);
or UO_366 (O_366,N_24609,N_18866);
nand UO_367 (O_367,N_24387,N_18896);
and UO_368 (O_368,N_21159,N_19883);
nor UO_369 (O_369,N_20001,N_18918);
or UO_370 (O_370,N_19712,N_20346);
nor UO_371 (O_371,N_20892,N_20659);
xor UO_372 (O_372,N_23417,N_23974);
xor UO_373 (O_373,N_23833,N_23128);
xor UO_374 (O_374,N_21706,N_22773);
nor UO_375 (O_375,N_23182,N_18899);
nand UO_376 (O_376,N_22835,N_23555);
or UO_377 (O_377,N_23345,N_23736);
xnor UO_378 (O_378,N_24419,N_20732);
xnor UO_379 (O_379,N_19629,N_24322);
nor UO_380 (O_380,N_22266,N_24048);
nand UO_381 (O_381,N_21652,N_19722);
and UO_382 (O_382,N_23485,N_20786);
and UO_383 (O_383,N_20611,N_19839);
and UO_384 (O_384,N_24515,N_20503);
nor UO_385 (O_385,N_24800,N_20265);
xor UO_386 (O_386,N_21971,N_19390);
or UO_387 (O_387,N_23185,N_22813);
and UO_388 (O_388,N_21410,N_19723);
nor UO_389 (O_389,N_21135,N_20405);
or UO_390 (O_390,N_21472,N_22921);
and UO_391 (O_391,N_21336,N_23861);
nor UO_392 (O_392,N_21363,N_23076);
nand UO_393 (O_393,N_22944,N_23754);
nor UO_394 (O_394,N_23216,N_23766);
xnor UO_395 (O_395,N_20756,N_20270);
nor UO_396 (O_396,N_21060,N_23546);
and UO_397 (O_397,N_20314,N_24960);
xor UO_398 (O_398,N_18912,N_23363);
xnor UO_399 (O_399,N_21641,N_23145);
nor UO_400 (O_400,N_23924,N_21539);
or UO_401 (O_401,N_23376,N_24436);
and UO_402 (O_402,N_22941,N_20447);
and UO_403 (O_403,N_20004,N_21791);
nand UO_404 (O_404,N_21953,N_21603);
or UO_405 (O_405,N_24290,N_19564);
or UO_406 (O_406,N_19321,N_21792);
nand UO_407 (O_407,N_20197,N_23539);
and UO_408 (O_408,N_24017,N_23504);
nor UO_409 (O_409,N_23604,N_22110);
and UO_410 (O_410,N_20811,N_21725);
or UO_411 (O_411,N_21242,N_23600);
xor UO_412 (O_412,N_19831,N_20813);
nor UO_413 (O_413,N_23282,N_20138);
xor UO_414 (O_414,N_20194,N_24303);
or UO_415 (O_415,N_24281,N_22431);
nor UO_416 (O_416,N_23738,N_19965);
or UO_417 (O_417,N_19640,N_23797);
nand UO_418 (O_418,N_18980,N_19508);
nor UO_419 (O_419,N_22289,N_21396);
or UO_420 (O_420,N_20826,N_19376);
nand UO_421 (O_421,N_22418,N_22052);
nor UO_422 (O_422,N_20416,N_22087);
nor UO_423 (O_423,N_22561,N_22790);
nor UO_424 (O_424,N_23424,N_20633);
or UO_425 (O_425,N_20120,N_19030);
or UO_426 (O_426,N_19854,N_18849);
or UO_427 (O_427,N_23929,N_21296);
nor UO_428 (O_428,N_23963,N_19359);
nand UO_429 (O_429,N_22321,N_21276);
and UO_430 (O_430,N_23979,N_19247);
nand UO_431 (O_431,N_24844,N_21799);
xnor UO_432 (O_432,N_24791,N_22890);
nor UO_433 (O_433,N_23855,N_23069);
or UO_434 (O_434,N_21676,N_23255);
and UO_435 (O_435,N_19004,N_22905);
nand UO_436 (O_436,N_21506,N_20371);
nand UO_437 (O_437,N_23354,N_23133);
and UO_438 (O_438,N_20679,N_20086);
or UO_439 (O_439,N_20057,N_21701);
nand UO_440 (O_440,N_24255,N_20554);
nor UO_441 (O_441,N_20844,N_20760);
xnor UO_442 (O_442,N_21959,N_24291);
nand UO_443 (O_443,N_19507,N_20836);
xor UO_444 (O_444,N_20660,N_22535);
and UO_445 (O_445,N_24715,N_21305);
and UO_446 (O_446,N_23811,N_22879);
nor UO_447 (O_447,N_23072,N_24980);
nand UO_448 (O_448,N_21540,N_19186);
or UO_449 (O_449,N_22303,N_23163);
nor UO_450 (O_450,N_19382,N_22774);
and UO_451 (O_451,N_18877,N_19264);
nor UO_452 (O_452,N_24418,N_23992);
or UO_453 (O_453,N_23753,N_20578);
and UO_454 (O_454,N_22316,N_23894);
or UO_455 (O_455,N_18766,N_19998);
or UO_456 (O_456,N_24058,N_21601);
and UO_457 (O_457,N_20406,N_23656);
nand UO_458 (O_458,N_21562,N_23768);
and UO_459 (O_459,N_22049,N_23106);
nor UO_460 (O_460,N_19083,N_24139);
or UO_461 (O_461,N_24610,N_22044);
nor UO_462 (O_462,N_19245,N_23335);
and UO_463 (O_463,N_20038,N_22766);
xnor UO_464 (O_464,N_23720,N_18997);
nor UO_465 (O_465,N_21314,N_18765);
and UO_466 (O_466,N_21341,N_24098);
xnor UO_467 (O_467,N_19703,N_20403);
or UO_468 (O_468,N_24282,N_20074);
and UO_469 (O_469,N_19972,N_24184);
nand UO_470 (O_470,N_21798,N_19066);
and UO_471 (O_471,N_20991,N_20272);
nor UO_472 (O_472,N_20997,N_24526);
nor UO_473 (O_473,N_19250,N_21057);
or UO_474 (O_474,N_21650,N_23085);
and UO_475 (O_475,N_18944,N_24838);
and UO_476 (O_476,N_19279,N_21635);
or UO_477 (O_477,N_19919,N_19090);
and UO_478 (O_478,N_23225,N_23126);
nand UO_479 (O_479,N_24081,N_24602);
xnor UO_480 (O_480,N_19315,N_21493);
nor UO_481 (O_481,N_24194,N_20909);
or UO_482 (O_482,N_23207,N_20648);
and UO_483 (O_483,N_24946,N_20533);
nand UO_484 (O_484,N_23897,N_21445);
nand UO_485 (O_485,N_23714,N_24074);
nand UO_486 (O_486,N_24159,N_21839);
xnor UO_487 (O_487,N_20041,N_22403);
and UO_488 (O_488,N_20006,N_22939);
or UO_489 (O_489,N_23698,N_23764);
xor UO_490 (O_490,N_20962,N_19785);
nand UO_491 (O_491,N_24792,N_24377);
and UO_492 (O_492,N_23143,N_19775);
nor UO_493 (O_493,N_23038,N_22660);
and UO_494 (O_494,N_24879,N_23557);
or UO_495 (O_495,N_24620,N_18812);
and UO_496 (O_496,N_19310,N_21313);
or UO_497 (O_497,N_22866,N_21986);
xor UO_498 (O_498,N_20438,N_23661);
nor UO_499 (O_499,N_24530,N_19150);
and UO_500 (O_500,N_22228,N_19858);
xnor UO_501 (O_501,N_23272,N_20115);
and UO_502 (O_502,N_21879,N_19064);
nand UO_503 (O_503,N_23662,N_23864);
and UO_504 (O_504,N_19421,N_23473);
and UO_505 (O_505,N_20444,N_24928);
or UO_506 (O_506,N_21930,N_24038);
or UO_507 (O_507,N_21256,N_23247);
xnor UO_508 (O_508,N_20231,N_23311);
nand UO_509 (O_509,N_22842,N_21980);
nand UO_510 (O_510,N_21928,N_22839);
nand UO_511 (O_511,N_19163,N_19161);
nand UO_512 (O_512,N_22478,N_24421);
nor UO_513 (O_513,N_22436,N_24703);
xor UO_514 (O_514,N_21177,N_21157);
nor UO_515 (O_515,N_20837,N_21462);
nand UO_516 (O_516,N_19172,N_22613);
xnor UO_517 (O_517,N_20858,N_22165);
xnor UO_518 (O_518,N_19182,N_24488);
xnor UO_519 (O_519,N_24940,N_23730);
and UO_520 (O_520,N_22777,N_18774);
nand UO_521 (O_521,N_23102,N_21780);
nor UO_522 (O_522,N_24011,N_19274);
nor UO_523 (O_523,N_21033,N_24306);
xnor UO_524 (O_524,N_19877,N_23248);
and UO_525 (O_525,N_20830,N_20472);
or UO_526 (O_526,N_21634,N_19311);
xnor UO_527 (O_527,N_23937,N_21028);
nand UO_528 (O_528,N_20178,N_22329);
nand UO_529 (O_529,N_19180,N_24545);
and UO_530 (O_530,N_21510,N_20051);
xnor UO_531 (O_531,N_20827,N_20122);
or UO_532 (O_532,N_24084,N_19093);
nand UO_533 (O_533,N_22323,N_24444);
or UO_534 (O_534,N_20093,N_19975);
and UO_535 (O_535,N_21628,N_21533);
nor UO_536 (O_536,N_21346,N_22274);
nor UO_537 (O_537,N_20439,N_19403);
xnor UO_538 (O_538,N_23962,N_24016);
nand UO_539 (O_539,N_24391,N_19962);
nand UO_540 (O_540,N_23694,N_22812);
xnor UO_541 (O_541,N_20252,N_20030);
nor UO_542 (O_542,N_22901,N_19146);
nor UO_543 (O_543,N_24493,N_24020);
nor UO_544 (O_544,N_24528,N_23016);
and UO_545 (O_545,N_23108,N_24383);
nor UO_546 (O_546,N_22718,N_24392);
nand UO_547 (O_547,N_24454,N_21093);
and UO_548 (O_548,N_24815,N_23826);
nor UO_549 (O_549,N_24131,N_22405);
xor UO_550 (O_550,N_20334,N_19286);
and UO_551 (O_551,N_20666,N_21762);
or UO_552 (O_552,N_23487,N_21581);
nand UO_553 (O_553,N_24191,N_18893);
nand UO_554 (O_554,N_21888,N_22364);
nand UO_555 (O_555,N_23997,N_18962);
nand UO_556 (O_556,N_21209,N_21732);
or UO_557 (O_557,N_24096,N_19343);
nor UO_558 (O_558,N_23074,N_24591);
nor UO_559 (O_559,N_23415,N_21213);
nor UO_560 (O_560,N_19347,N_24922);
or UO_561 (O_561,N_23476,N_24888);
xor UO_562 (O_562,N_21335,N_24949);
nor UO_563 (O_563,N_20510,N_24725);
and UO_564 (O_564,N_20731,N_21245);
nor UO_565 (O_565,N_21501,N_24640);
nor UO_566 (O_566,N_21783,N_21061);
nand UO_567 (O_567,N_20388,N_22816);
and UO_568 (O_568,N_19119,N_23988);
xnor UO_569 (O_569,N_19094,N_22684);
or UO_570 (O_570,N_23776,N_22477);
and UO_571 (O_571,N_19360,N_23202);
nor UO_572 (O_572,N_21052,N_21270);
nand UO_573 (O_573,N_22277,N_23721);
xor UO_574 (O_574,N_20343,N_22848);
nor UO_575 (O_575,N_24453,N_22127);
nor UO_576 (O_576,N_22570,N_22164);
nand UO_577 (O_577,N_23553,N_21359);
or UO_578 (O_578,N_21967,N_20046);
nor UO_579 (O_579,N_21185,N_20212);
nor UO_580 (O_580,N_24156,N_20623);
or UO_581 (O_581,N_18946,N_22852);
and UO_582 (O_582,N_23757,N_20410);
nor UO_583 (O_583,N_22786,N_20255);
nand UO_584 (O_584,N_24775,N_22709);
and UO_585 (O_585,N_19750,N_20965);
and UO_586 (O_586,N_18876,N_24372);
nor UO_587 (O_587,N_23122,N_19847);
or UO_588 (O_588,N_19251,N_24819);
xor UO_589 (O_589,N_21559,N_22663);
nor UO_590 (O_590,N_24056,N_20301);
nor UO_591 (O_591,N_23702,N_23818);
nor UO_592 (O_592,N_20321,N_18751);
or UO_593 (O_593,N_23176,N_19980);
and UO_594 (O_594,N_19006,N_21711);
nor UO_595 (O_595,N_23004,N_20294);
xor UO_596 (O_596,N_21849,N_20126);
nand UO_597 (O_597,N_24825,N_19023);
or UO_598 (O_598,N_23276,N_24238);
and UO_599 (O_599,N_20323,N_21546);
or UO_600 (O_600,N_21830,N_23190);
and UO_601 (O_601,N_24520,N_24019);
nor UO_602 (O_602,N_19731,N_19707);
nor UO_603 (O_603,N_18789,N_21374);
and UO_604 (O_604,N_23127,N_23807);
and UO_605 (O_605,N_24938,N_24365);
nor UO_606 (O_606,N_21931,N_21890);
nor UO_607 (O_607,N_22648,N_21611);
nand UO_608 (O_608,N_20945,N_21475);
nor UO_609 (O_609,N_20363,N_22999);
or UO_610 (O_610,N_21145,N_20445);
nor UO_611 (O_611,N_24064,N_21500);
or UO_612 (O_612,N_21303,N_21016);
nor UO_613 (O_613,N_24105,N_21364);
and UO_614 (O_614,N_22676,N_22552);
and UO_615 (O_615,N_22212,N_23373);
or UO_616 (O_616,N_19211,N_20446);
xor UO_617 (O_617,N_20996,N_24909);
or UO_618 (O_618,N_22809,N_19248);
xnor UO_619 (O_619,N_22614,N_23439);
or UO_620 (O_620,N_22463,N_19373);
and UO_621 (O_621,N_23901,N_19079);
xor UO_622 (O_622,N_20530,N_19979);
nor UO_623 (O_623,N_21787,N_23809);
xor UO_624 (O_624,N_20529,N_23550);
nor UO_625 (O_625,N_21181,N_20436);
xnor UO_626 (O_626,N_24644,N_23078);
nand UO_627 (O_627,N_19896,N_19433);
or UO_628 (O_628,N_21343,N_23343);
xnor UO_629 (O_629,N_22860,N_23663);
nand UO_630 (O_630,N_22401,N_22085);
nand UO_631 (O_631,N_23179,N_19594);
and UO_632 (O_632,N_22685,N_20113);
xnor UO_633 (O_633,N_19529,N_21512);
or UO_634 (O_634,N_18941,N_23328);
nand UO_635 (O_635,N_22065,N_24254);
nand UO_636 (O_636,N_20757,N_19226);
xnor UO_637 (O_637,N_21182,N_22173);
nor UO_638 (O_638,N_21822,N_22420);
nand UO_639 (O_639,N_21355,N_21240);
and UO_640 (O_640,N_24417,N_19968);
xor UO_641 (O_641,N_20963,N_18926);
xor UO_642 (O_642,N_20037,N_23058);
nor UO_643 (O_643,N_24598,N_22119);
or UO_644 (O_644,N_24551,N_21901);
nor UO_645 (O_645,N_19801,N_20200);
xnor UO_646 (O_646,N_19626,N_23693);
and UO_647 (O_647,N_20034,N_21767);
xor UO_648 (O_648,N_21588,N_20895);
or UO_649 (O_649,N_22155,N_24846);
xor UO_650 (O_650,N_22397,N_21140);
nor UO_651 (O_651,N_20356,N_24331);
xnor UO_652 (O_652,N_23563,N_19649);
nor UO_653 (O_653,N_24646,N_22365);
xor UO_654 (O_654,N_20320,N_19852);
and UO_655 (O_655,N_19153,N_24966);
nand UO_656 (O_656,N_23595,N_18786);
xor UO_657 (O_657,N_22440,N_20557);
xnor UO_658 (O_658,N_22557,N_20062);
xor UO_659 (O_659,N_23355,N_21439);
nand UO_660 (O_660,N_24518,N_19867);
and UO_661 (O_661,N_22130,N_21285);
and UO_662 (O_662,N_24758,N_24532);
nand UO_663 (O_663,N_23796,N_22211);
nor UO_664 (O_664,N_19840,N_24314);
and UO_665 (O_665,N_20661,N_23853);
and UO_666 (O_666,N_22904,N_24262);
nor UO_667 (O_667,N_20627,N_19320);
nand UO_668 (O_668,N_24876,N_22413);
nand UO_669 (O_669,N_22863,N_21716);
or UO_670 (O_670,N_24079,N_22491);
and UO_671 (O_671,N_24776,N_20259);
and UO_672 (O_672,N_21691,N_21196);
xnor UO_673 (O_673,N_20743,N_20071);
nor UO_674 (O_674,N_20109,N_24567);
nor UO_675 (O_675,N_20548,N_19881);
nand UO_676 (O_676,N_21768,N_22146);
nor UO_677 (O_677,N_20766,N_24227);
and UO_678 (O_678,N_20603,N_24158);
nand UO_679 (O_679,N_20278,N_19503);
and UO_680 (O_680,N_21083,N_24978);
or UO_681 (O_681,N_24193,N_24936);
and UO_682 (O_682,N_21294,N_19355);
xor UO_683 (O_683,N_23456,N_18851);
nor UO_684 (O_684,N_19236,N_21805);
nand UO_685 (O_685,N_20710,N_24228);
and UO_686 (O_686,N_21646,N_19469);
and UO_687 (O_687,N_23574,N_18988);
or UO_688 (O_688,N_18934,N_22588);
or UO_689 (O_689,N_23759,N_20976);
nor UO_690 (O_690,N_22964,N_20101);
nor UO_691 (O_691,N_20741,N_23432);
xnor UO_692 (O_692,N_19967,N_23168);
xor UO_693 (O_693,N_19178,N_20240);
or UO_694 (O_694,N_22174,N_21672);
or UO_695 (O_695,N_20938,N_21536);
and UO_696 (O_696,N_23920,N_23281);
nor UO_697 (O_697,N_24065,N_19542);
or UO_698 (O_698,N_23407,N_19451);
xnor UO_699 (O_699,N_23681,N_22826);
or UO_700 (O_700,N_22740,N_23752);
and UO_701 (O_701,N_20274,N_21411);
and UO_702 (O_702,N_24313,N_20576);
or UO_703 (O_703,N_21007,N_23441);
nand UO_704 (O_704,N_21637,N_24559);
xor UO_705 (O_705,N_19837,N_24347);
xor UO_706 (O_706,N_19436,N_21087);
nor UO_707 (O_707,N_24973,N_23874);
and UO_708 (O_708,N_23318,N_22649);
xnor UO_709 (O_709,N_24356,N_20100);
and UO_710 (O_710,N_19598,N_21630);
xnor UO_711 (O_711,N_23147,N_22254);
nand UO_712 (O_712,N_24604,N_19991);
and UO_713 (O_713,N_23482,N_22186);
xor UO_714 (O_714,N_21128,N_24037);
and UO_715 (O_715,N_19971,N_22352);
or UO_716 (O_716,N_20003,N_22586);
or UO_717 (O_717,N_20966,N_20296);
and UO_718 (O_718,N_19384,N_22639);
nor UO_719 (O_719,N_24008,N_20007);
and UO_720 (O_720,N_22655,N_21257);
nor UO_721 (O_721,N_19614,N_22400);
nor UO_722 (O_722,N_22720,N_21243);
xnor UO_723 (O_723,N_24459,N_21114);
xor UO_724 (O_724,N_19921,N_24548);
and UO_725 (O_725,N_20485,N_23314);
nand UO_726 (O_726,N_20375,N_21253);
and UO_727 (O_727,N_20580,N_18984);
nor UO_728 (O_728,N_22810,N_19523);
xnor UO_729 (O_729,N_19265,N_19029);
and UO_730 (O_730,N_20910,N_23840);
and UO_731 (O_731,N_24734,N_24007);
and UO_732 (O_732,N_21899,N_21752);
and UO_733 (O_733,N_23243,N_20325);
nand UO_734 (O_734,N_23223,N_21961);
or UO_735 (O_735,N_18756,N_21354);
nor UO_736 (O_736,N_18875,N_20395);
nor UO_737 (O_737,N_20546,N_21705);
nand UO_738 (O_738,N_21979,N_23560);
nand UO_739 (O_739,N_20566,N_20876);
xnor UO_740 (O_740,N_22559,N_23336);
nand UO_741 (O_741,N_20106,N_20629);
xnor UO_742 (O_742,N_24416,N_19558);
nand UO_743 (O_743,N_21453,N_24731);
nor UO_744 (O_744,N_21862,N_21604);
nor UO_745 (O_745,N_24899,N_21851);
xnor UO_746 (O_746,N_21143,N_24832);
nor UO_747 (O_747,N_20016,N_19228);
and UO_748 (O_748,N_22233,N_20284);
nor UO_749 (O_749,N_24619,N_21013);
nor UO_750 (O_750,N_18867,N_22638);
nor UO_751 (O_751,N_20082,N_23391);
nor UO_752 (O_752,N_21668,N_21137);
or UO_753 (O_753,N_21102,N_19970);
nand UO_754 (O_754,N_22801,N_19651);
and UO_755 (O_755,N_20772,N_22035);
nand UO_756 (O_756,N_18958,N_21272);
and UO_757 (O_757,N_22370,N_24534);
or UO_758 (O_758,N_20008,N_23493);
nand UO_759 (O_759,N_23201,N_21062);
and UO_760 (O_760,N_23778,N_22417);
xor UO_761 (O_761,N_24685,N_21881);
nor UO_762 (O_762,N_21273,N_22969);
nand UO_763 (O_763,N_22688,N_22635);
and UO_764 (O_764,N_19116,N_22415);
and UO_765 (O_765,N_23598,N_22229);
and UO_766 (O_766,N_19535,N_22971);
or UO_767 (O_767,N_20359,N_21187);
or UO_768 (O_768,N_23219,N_19798);
nor UO_769 (O_769,N_20450,N_19708);
xor UO_770 (O_770,N_23726,N_19978);
or UO_771 (O_771,N_23771,N_21599);
or UO_772 (O_772,N_23203,N_19850);
and UO_773 (O_773,N_22126,N_19813);
or UO_774 (O_774,N_24711,N_21577);
nor UO_775 (O_775,N_22427,N_19428);
or UO_776 (O_776,N_22028,N_20985);
and UO_777 (O_777,N_19539,N_20047);
xnor UO_778 (O_778,N_19670,N_22297);
xor UO_779 (O_779,N_21022,N_21910);
or UO_780 (O_780,N_22093,N_24470);
or UO_781 (O_781,N_23635,N_18806);
or UO_782 (O_782,N_19643,N_23668);
or UO_783 (O_783,N_19037,N_20131);
xor UO_784 (O_784,N_22550,N_19055);
nor UO_785 (O_785,N_22481,N_24732);
and UO_786 (O_786,N_21105,N_21863);
xor UO_787 (O_787,N_22219,N_21954);
nor UO_788 (O_788,N_21331,N_19190);
and UO_789 (O_789,N_24592,N_23397);
or UO_790 (O_790,N_22554,N_23359);
nand UO_791 (O_791,N_23009,N_24886);
xnor UO_792 (O_792,N_21781,N_21810);
nor UO_793 (O_793,N_21999,N_24097);
xnor UO_794 (O_794,N_24175,N_21081);
or UO_795 (O_795,N_24450,N_20733);
nor UO_796 (O_796,N_24893,N_23385);
or UO_797 (O_797,N_24593,N_22027);
and UO_798 (O_798,N_22967,N_21560);
or UO_799 (O_799,N_19325,N_22922);
or UO_800 (O_800,N_20313,N_21978);
or UO_801 (O_801,N_19429,N_24167);
nor UO_802 (O_802,N_22234,N_24256);
nand UO_803 (O_803,N_21987,N_21047);
or UO_804 (O_804,N_22269,N_21449);
and UO_805 (O_805,N_19176,N_23703);
or UO_806 (O_806,N_20610,N_24067);
and UO_807 (O_807,N_22392,N_22565);
nor UO_808 (O_808,N_23938,N_20350);
nand UO_809 (O_809,N_22092,N_20787);
and UO_810 (O_810,N_22151,N_19427);
nor UO_811 (O_811,N_18971,N_21997);
and UO_812 (O_812,N_21947,N_21558);
nor UO_813 (O_813,N_23339,N_22576);
or UO_814 (O_814,N_22925,N_19516);
nand UO_815 (O_815,N_22933,N_24108);
xnor UO_816 (O_816,N_20208,N_18992);
nor UO_817 (O_817,N_22763,N_21920);
xnor UO_818 (O_818,N_24452,N_20358);
xor UO_819 (O_819,N_22344,N_19611);
nor UO_820 (O_820,N_23450,N_20386);
or UO_821 (O_821,N_24752,N_23887);
nor UO_822 (O_822,N_21921,N_19140);
and UO_823 (O_823,N_20879,N_23973);
xor UO_824 (O_824,N_21094,N_21323);
or UO_825 (O_825,N_19765,N_20614);
nor UO_826 (O_826,N_22963,N_24041);
and UO_827 (O_827,N_23524,N_19799);
nand UO_828 (O_828,N_21169,N_20917);
nor UO_829 (O_829,N_21186,N_24892);
nor UO_830 (O_830,N_20688,N_20293);
nand UO_831 (O_831,N_24872,N_21089);
nor UO_832 (O_832,N_20118,N_24334);
nand UO_833 (O_833,N_21609,N_23309);
xnor UO_834 (O_834,N_19461,N_21733);
nor UO_835 (O_835,N_21258,N_20513);
nand UO_836 (O_836,N_18801,N_22859);
or UO_837 (O_837,N_18796,N_24259);
xor UO_838 (O_838,N_19271,N_22681);
nand UO_839 (O_839,N_19167,N_23116);
nand UO_840 (O_840,N_19448,N_19745);
xnor UO_841 (O_841,N_19297,N_18762);
nor UO_842 (O_842,N_23372,N_19162);
or UO_843 (O_843,N_21108,N_22171);
and UO_844 (O_844,N_19024,N_19354);
and UO_845 (O_845,N_23561,N_20537);
and UO_846 (O_846,N_20726,N_18813);
xor UO_847 (O_847,N_20042,N_23791);
nand UO_848 (O_848,N_20437,N_24535);
xor UO_849 (O_849,N_20460,N_20506);
nand UO_850 (O_850,N_24102,N_23562);
xor UO_851 (O_851,N_21050,N_21138);
or UO_852 (O_852,N_21889,N_24676);
or UO_853 (O_853,N_22122,N_21748);
nor UO_854 (O_854,N_20574,N_23984);
xnor UO_855 (O_855,N_19028,N_23888);
nor UO_856 (O_856,N_19296,N_19929);
nand UO_857 (O_857,N_23334,N_19009);
nand UO_858 (O_858,N_21996,N_19341);
nor UO_859 (O_859,N_23572,N_19958);
xnor UO_860 (O_860,N_20425,N_19111);
or UO_861 (O_861,N_19475,N_20764);
or UO_862 (O_862,N_21970,N_21778);
xor UO_863 (O_863,N_20998,N_24968);
xor UO_864 (O_864,N_24271,N_19788);
and UO_865 (O_865,N_21198,N_21421);
nor UO_866 (O_866,N_23530,N_21441);
or UO_867 (O_867,N_20124,N_24767);
or UO_868 (O_868,N_19181,N_22759);
and UO_869 (O_869,N_22355,N_21096);
or UO_870 (O_870,N_22194,N_24507);
nand UO_871 (O_871,N_20536,N_23559);
and UO_872 (O_872,N_24179,N_19002);
xnor UO_873 (O_873,N_23695,N_22260);
and UO_874 (O_874,N_22538,N_23765);
or UO_875 (O_875,N_23365,N_23346);
xnor UO_876 (O_876,N_23065,N_22772);
nand UO_877 (O_877,N_22079,N_23253);
xor UO_878 (O_878,N_21984,N_19016);
or UO_879 (O_879,N_24430,N_19950);
nor UO_880 (O_880,N_20957,N_24916);
or UO_881 (O_881,N_23718,N_19100);
nand UO_882 (O_882,N_19607,N_22885);
xor UO_883 (O_883,N_21823,N_19070);
or UO_884 (O_884,N_23616,N_20932);
nand UO_885 (O_885,N_18948,N_22652);
nand UO_886 (O_886,N_23511,N_22665);
nor UO_887 (O_887,N_24176,N_20318);
nor UO_888 (O_888,N_19893,N_24381);
or UO_889 (O_889,N_22235,N_22849);
xnor UO_890 (O_890,N_22643,N_23865);
xor UO_891 (O_891,N_21833,N_20845);
or UO_892 (O_892,N_21255,N_23465);
nor UO_893 (O_893,N_20788,N_23783);
nor UO_894 (O_894,N_24569,N_23262);
xnor UO_895 (O_895,N_21095,N_23613);
xnor UO_896 (O_896,N_24168,N_20686);
and UO_897 (O_897,N_22784,N_20540);
nand UO_898 (O_898,N_20397,N_19901);
nor UO_899 (O_899,N_21395,N_21908);
nand UO_900 (O_900,N_23958,N_19187);
and UO_901 (O_901,N_19862,N_18816);
or UO_902 (O_902,N_21854,N_24439);
or UO_903 (O_903,N_24482,N_24962);
or UO_904 (O_904,N_20058,N_24330);
or UO_905 (O_905,N_21365,N_20582);
xor UO_906 (O_906,N_19305,N_24197);
nor UO_907 (O_907,N_22920,N_20137);
and UO_908 (O_908,N_24577,N_20602);
xor UO_909 (O_909,N_24568,N_24160);
and UO_910 (O_910,N_21681,N_20778);
nor UO_911 (O_911,N_20166,N_24140);
nor UO_912 (O_912,N_21720,N_24210);
nand UO_913 (O_913,N_19524,N_21275);
nor UO_914 (O_914,N_21107,N_24320);
nand UO_915 (O_915,N_23566,N_20153);
nand UO_916 (O_916,N_22680,N_23538);
and UO_917 (O_917,N_20309,N_23490);
and UO_918 (O_918,N_19459,N_24062);
or UO_919 (O_919,N_22728,N_23399);
nor UO_920 (O_920,N_24656,N_20805);
xor UO_921 (O_921,N_24277,N_19698);
nand UO_922 (O_922,N_21254,N_19147);
or UO_923 (O_923,N_20527,N_19956);
and UO_924 (O_924,N_23433,N_20604);
and UO_925 (O_925,N_23543,N_21597);
xor UO_926 (O_926,N_22412,N_19548);
and UO_927 (O_927,N_23519,N_21148);
or UO_928 (O_928,N_21753,N_21503);
and UO_929 (O_929,N_24150,N_20097);
nor UO_930 (O_930,N_21821,N_23934);
or UO_931 (O_931,N_24580,N_22111);
nand UO_932 (O_932,N_19702,N_24460);
or UO_933 (O_933,N_23327,N_22387);
nand UO_934 (O_934,N_24824,N_22528);
xnor UO_935 (O_935,N_22597,N_24466);
or UO_936 (O_936,N_21511,N_20480);
nand UO_937 (O_937,N_24687,N_19168);
or UO_938 (O_938,N_20517,N_24708);
or UO_939 (O_939,N_20183,N_23447);
xor UO_940 (O_940,N_20257,N_20292);
nor UO_941 (O_941,N_23580,N_22506);
nor UO_942 (O_942,N_24898,N_24665);
nand UO_943 (O_943,N_20432,N_22125);
or UO_944 (O_944,N_19113,N_23954);
or UO_945 (O_945,N_24200,N_21100);
nor UO_946 (O_946,N_22970,N_21557);
xnor UO_947 (O_947,N_24638,N_20443);
nand UO_948 (O_948,N_19038,N_20865);
nand UO_949 (O_949,N_20925,N_22714);
xnor UO_950 (O_950,N_23576,N_23837);
and UO_951 (O_951,N_22072,N_21125);
nor UO_952 (O_952,N_19632,N_19927);
or UO_953 (O_953,N_24148,N_23957);
and UO_954 (O_954,N_21633,N_24692);
or UO_955 (O_955,N_24573,N_23077);
nand UO_956 (O_956,N_21587,N_23540);
nor UO_957 (O_957,N_21078,N_24120);
nor UO_958 (O_958,N_20463,N_19589);
nand UO_959 (O_959,N_19821,N_24858);
nand UO_960 (O_960,N_20647,N_23382);
nand UO_961 (O_961,N_24442,N_22324);
nor UO_962 (O_962,N_24028,N_20641);
xor UO_963 (O_963,N_23919,N_18810);
and UO_964 (O_964,N_23849,N_24113);
and UO_965 (O_965,N_20023,N_22823);
or UO_966 (O_966,N_20874,N_24981);
xor UO_967 (O_967,N_19907,N_24471);
xnor UO_968 (O_968,N_23536,N_22911);
and UO_969 (O_969,N_21570,N_20593);
xnor UO_970 (O_970,N_24304,N_24855);
nor UO_971 (O_971,N_20434,N_20672);
nand UO_972 (O_972,N_22179,N_23620);
nand UO_973 (O_973,N_24857,N_24681);
xnor UO_974 (O_974,N_19866,N_21621);
and UO_975 (O_975,N_22936,N_24914);
and UO_976 (O_976,N_21988,N_21841);
nor UO_977 (O_977,N_21333,N_19400);
or UO_978 (O_978,N_20682,N_20793);
or UO_979 (O_979,N_19817,N_23129);
nand UO_980 (O_980,N_19114,N_24270);
and UO_981 (O_981,N_21413,N_19326);
xor UO_982 (O_982,N_19527,N_21846);
nor UO_983 (O_983,N_20054,N_21368);
xor UO_984 (O_984,N_19822,N_24206);
or UO_985 (O_985,N_20878,N_22683);
and UO_986 (O_986,N_22340,N_19838);
and UO_987 (O_987,N_21523,N_22043);
or UO_988 (O_988,N_20498,N_22441);
xor UO_989 (O_989,N_20401,N_24761);
or UO_990 (O_990,N_20930,N_22099);
xor UO_991 (O_991,N_20851,N_24581);
or UO_992 (O_992,N_23584,N_20979);
xor UO_993 (O_993,N_21973,N_23209);
nand UO_994 (O_994,N_23429,N_22878);
xnor UO_995 (O_995,N_22836,N_23998);
and UO_996 (O_996,N_22262,N_23050);
xor UO_997 (O_997,N_18904,N_22915);
xnor UO_998 (O_998,N_22283,N_22479);
or UO_999 (O_999,N_24143,N_19282);
nor UO_1000 (O_1000,N_19101,N_22086);
nand UO_1001 (O_1001,N_22433,N_23256);
and UO_1002 (O_1002,N_19859,N_24833);
nor UO_1003 (O_1003,N_19219,N_21485);
nor UO_1004 (O_1004,N_24491,N_23389);
or UO_1005 (O_1005,N_24297,N_22906);
nand UO_1006 (O_1006,N_21654,N_19572);
and UO_1007 (O_1007,N_23854,N_22462);
xor UO_1008 (O_1008,N_22311,N_24153);
or UO_1009 (O_1009,N_23939,N_22811);
nand UO_1010 (O_1010,N_23542,N_18955);
xor UO_1011 (O_1011,N_22980,N_21167);
xnor UO_1012 (O_1012,N_22372,N_23032);
or UO_1013 (O_1013,N_23333,N_19369);
xor UO_1014 (O_1014,N_23627,N_20799);
or UO_1015 (O_1015,N_24448,N_24287);
or UO_1016 (O_1016,N_21316,N_20217);
nand UO_1017 (O_1017,N_21906,N_21147);
nand UO_1018 (O_1018,N_18782,N_19345);
and UO_1019 (O_1019,N_21328,N_19627);
nor UO_1020 (O_1020,N_24795,N_19631);
nor UO_1021 (O_1021,N_20921,N_22207);
nand UO_1022 (O_1022,N_19717,N_22990);
nor UO_1023 (O_1023,N_19806,N_21161);
nor UO_1024 (O_1024,N_22242,N_22090);
or UO_1025 (O_1025,N_24601,N_19191);
xor UO_1026 (O_1026,N_23657,N_21831);
nand UO_1027 (O_1027,N_24989,N_23716);
nor UO_1028 (O_1028,N_21829,N_19869);
nor UO_1029 (O_1029,N_18938,N_20449);
and UO_1030 (O_1030,N_20612,N_19879);
nand UO_1031 (O_1031,N_19569,N_19138);
nand UO_1032 (O_1032,N_23590,N_19084);
nor UO_1033 (O_1033,N_18836,N_24913);
xnor UO_1034 (O_1034,N_24987,N_20150);
and UO_1035 (O_1035,N_20649,N_21636);
nor UO_1036 (O_1036,N_23578,N_18973);
nor UO_1037 (O_1037,N_24746,N_19193);
and UO_1038 (O_1038,N_21929,N_18903);
nand UO_1039 (O_1039,N_19225,N_23374);
xnor UO_1040 (O_1040,N_24562,N_23435);
and UO_1041 (O_1041,N_21068,N_22286);
and UO_1042 (O_1042,N_21788,N_24995);
nor UO_1043 (O_1043,N_21614,N_20833);
or UO_1044 (O_1044,N_23608,N_18873);
and UO_1045 (O_1045,N_21963,N_20229);
or UO_1046 (O_1046,N_23951,N_24183);
or UO_1047 (O_1047,N_19054,N_19356);
nand UO_1048 (O_1048,N_20396,N_19201);
nand UO_1049 (O_1049,N_21315,N_20136);
and UO_1050 (O_1050,N_24807,N_20453);
and UO_1051 (O_1051,N_22762,N_23649);
and UO_1052 (O_1052,N_19665,N_24856);
and UO_1053 (O_1053,N_21339,N_23788);
and UO_1054 (O_1054,N_19909,N_21150);
and UO_1055 (O_1055,N_21223,N_19679);
and UO_1056 (O_1056,N_22654,N_21492);
nand UO_1057 (O_1057,N_24527,N_24426);
xnor UO_1058 (O_1058,N_22589,N_21238);
nand UO_1059 (O_1059,N_24225,N_22781);
nand UO_1060 (O_1060,N_24015,N_21040);
nor UO_1061 (O_1061,N_24326,N_19424);
nand UO_1062 (O_1062,N_24623,N_22568);
or UO_1063 (O_1063,N_21131,N_19912);
nand UO_1064 (O_1064,N_24477,N_23160);
or UO_1065 (O_1065,N_21448,N_23056);
and UO_1066 (O_1066,N_21813,N_24046);
or UO_1067 (O_1067,N_21127,N_21782);
nand UO_1068 (O_1068,N_24757,N_23183);
and UO_1069 (O_1069,N_24726,N_24820);
nor UO_1070 (O_1070,N_23956,N_19994);
xor UO_1071 (O_1071,N_21380,N_22987);
xnor UO_1072 (O_1072,N_23655,N_23105);
and UO_1073 (O_1073,N_22788,N_22703);
nand UO_1074 (O_1074,N_24103,N_24921);
and UO_1075 (O_1075,N_22956,N_21535);
nor UO_1076 (O_1076,N_21443,N_24605);
nor UO_1077 (O_1077,N_20952,N_19443);
xnor UO_1078 (O_1078,N_23648,N_19175);
and UO_1079 (O_1079,N_19386,N_23969);
xnor UO_1080 (O_1080,N_20095,N_23296);
nor UO_1081 (O_1081,N_19704,N_19338);
nor UO_1082 (O_1082,N_24871,N_24394);
and UO_1083 (O_1083,N_20140,N_20978);
nor UO_1084 (O_1084,N_23994,N_21865);
or UO_1085 (O_1085,N_20228,N_20354);
and UO_1086 (O_1086,N_21119,N_23673);
or UO_1087 (O_1087,N_24412,N_21897);
nand UO_1088 (O_1088,N_21771,N_24839);
or UO_1089 (O_1089,N_20994,N_23856);
and UO_1090 (O_1090,N_19284,N_22778);
or UO_1091 (O_1091,N_19738,N_20856);
or UO_1092 (O_1092,N_18821,N_20653);
xor UO_1093 (O_1093,N_21617,N_19447);
or UO_1094 (O_1094,N_20066,N_20180);
or UO_1095 (O_1095,N_22153,N_20831);
nor UO_1096 (O_1096,N_23039,N_19701);
and UO_1097 (O_1097,N_20056,N_23055);
or UO_1098 (O_1098,N_24380,N_19918);
nor UO_1099 (O_1099,N_22825,N_22307);
nor UO_1100 (O_1100,N_20722,N_23104);
or UO_1101 (O_1101,N_19551,N_24185);
xnor UO_1102 (O_1102,N_19892,N_22161);
nand UO_1103 (O_1103,N_18845,N_19039);
nor UO_1104 (O_1104,N_24908,N_19604);
nand UO_1105 (O_1105,N_23245,N_23719);
and UO_1106 (O_1106,N_22426,N_22545);
or UO_1107 (O_1107,N_24040,N_19580);
nand UO_1108 (O_1108,N_22383,N_19229);
nor UO_1109 (O_1109,N_22390,N_20276);
nor UO_1110 (O_1110,N_21917,N_21552);
nand UO_1111 (O_1111,N_19164,N_22599);
or UO_1112 (O_1112,N_24246,N_20759);
or UO_1113 (O_1113,N_23496,N_18853);
nand UO_1114 (O_1114,N_19777,N_22896);
nand UO_1115 (O_1115,N_20829,N_18834);
nand UO_1116 (O_1116,N_22706,N_21966);
xor UO_1117 (O_1117,N_19522,N_23640);
xnor UO_1118 (O_1118,N_23960,N_20541);
nor UO_1119 (O_1119,N_21199,N_19559);
nor UO_1120 (O_1120,N_22624,N_22872);
nor UO_1121 (O_1121,N_18769,N_24119);
and UO_1122 (O_1122,N_23689,N_19602);
and UO_1123 (O_1123,N_19000,N_19058);
xnor UO_1124 (O_1124,N_24991,N_19374);
xnor UO_1125 (O_1125,N_22674,N_19645);
or UO_1126 (O_1126,N_24486,N_22166);
nand UO_1127 (O_1127,N_20575,N_21564);
nor UO_1128 (O_1128,N_19675,N_18778);
and UO_1129 (O_1129,N_19300,N_23603);
and UO_1130 (O_1130,N_20803,N_20622);
and UO_1131 (O_1131,N_24047,N_23642);
or UO_1132 (O_1132,N_23132,N_21714);
and UO_1133 (O_1133,N_22071,N_23112);
and UO_1134 (O_1134,N_21054,N_22923);
xnor UO_1135 (O_1135,N_22302,N_21300);
xor UO_1136 (O_1136,N_20785,N_18869);
nor UO_1137 (O_1137,N_22951,N_21261);
xnor UO_1138 (O_1138,N_22189,N_24253);
or UO_1139 (O_1139,N_21853,N_19582);
or UO_1140 (O_1140,N_19855,N_22255);
nor UO_1141 (O_1141,N_22650,N_23193);
and UO_1142 (O_1142,N_24121,N_23117);
nand UO_1143 (O_1143,N_22679,N_20119);
and UO_1144 (O_1144,N_21101,N_20315);
and UO_1145 (O_1145,N_21576,N_20762);
nor UO_1146 (O_1146,N_24782,N_21554);
nor UO_1147 (O_1147,N_23273,N_20198);
nand UO_1148 (O_1148,N_24274,N_21219);
nand UO_1149 (O_1149,N_21764,N_23413);
nand UO_1150 (O_1150,N_23451,N_18986);
and UO_1151 (O_1151,N_24906,N_20995);
xor UO_1152 (O_1152,N_20088,N_22382);
or UO_1153 (O_1153,N_24424,N_22985);
and UO_1154 (O_1154,N_20499,N_24305);
nand UO_1155 (O_1155,N_20636,N_23761);
and UO_1156 (O_1156,N_18939,N_24641);
nand UO_1157 (O_1157,N_22000,N_20528);
nor UO_1158 (O_1158,N_19327,N_24214);
and UO_1159 (O_1159,N_21795,N_21490);
nor UO_1160 (O_1160,N_24723,N_20694);
nor UO_1161 (O_1161,N_21298,N_20908);
xnor UO_1162 (O_1162,N_24975,N_23144);
or UO_1163 (O_1163,N_22490,N_22930);
and UO_1164 (O_1164,N_24174,N_20108);
and UO_1165 (O_1165,N_23428,N_22226);
nor UO_1166 (O_1166,N_19188,N_20796);
nor UO_1167 (O_1167,N_20163,N_19025);
or UO_1168 (O_1168,N_22464,N_18907);
xnor UO_1169 (O_1169,N_20841,N_20027);
and UO_1170 (O_1170,N_23599,N_24743);
nor UO_1171 (O_1171,N_24467,N_20081);
nand UO_1172 (O_1172,N_18781,N_18923);
nand UO_1173 (O_1173,N_19984,N_19414);
nor UO_1174 (O_1174,N_23071,N_23321);
nor UO_1175 (O_1175,N_18758,N_24192);
nor UO_1176 (O_1176,N_24896,N_24289);
nor UO_1177 (O_1177,N_24123,N_22584);
nor UO_1178 (O_1178,N_18943,N_24180);
or UO_1179 (O_1179,N_24492,N_20288);
or UO_1180 (O_1180,N_21431,N_19720);
xor UO_1181 (O_1181,N_24446,N_24375);
or UO_1182 (O_1182,N_21804,N_22236);
and UO_1183 (O_1183,N_24597,N_23872);
and UO_1184 (O_1184,N_19672,N_21585);
nor UO_1185 (O_1185,N_18793,N_22575);
xor UO_1186 (O_1186,N_19195,N_21666);
nand UO_1187 (O_1187,N_22834,N_19536);
nand UO_1188 (O_1188,N_24312,N_19540);
or UO_1189 (O_1189,N_19205,N_22583);
nor UO_1190 (O_1190,N_20172,N_23461);
nand UO_1191 (O_1191,N_21180,N_24574);
nor UO_1192 (O_1192,N_19782,N_18965);
nor UO_1193 (O_1193,N_23772,N_19505);
nand UO_1194 (O_1194,N_23468,N_19068);
nor UO_1195 (O_1195,N_20236,N_20595);
or UO_1196 (O_1196,N_21221,N_18906);
nand UO_1197 (O_1197,N_18856,N_21012);
xnor UO_1198 (O_1198,N_19865,N_24413);
or UO_1199 (O_1199,N_22224,N_19959);
nor UO_1200 (O_1200,N_21583,N_23204);
xor UO_1201 (O_1201,N_23234,N_22172);
xnor UO_1202 (O_1202,N_21132,N_20377);
xor UO_1203 (O_1203,N_23706,N_22997);
nand UO_1204 (O_1204,N_18979,N_18976);
nand UO_1205 (O_1205,N_23965,N_19277);
xor UO_1206 (O_1206,N_21228,N_23257);
or UO_1207 (O_1207,N_22733,N_18833);
nand UO_1208 (O_1208,N_19783,N_20266);
or UO_1209 (O_1209,N_23737,N_23292);
nor UO_1210 (O_1210,N_21994,N_19700);
xor UO_1211 (O_1211,N_19473,N_20009);
nand UO_1212 (O_1212,N_22348,N_23062);
and UO_1213 (O_1213,N_23981,N_24702);
and UO_1214 (O_1214,N_21623,N_21918);
xor UO_1215 (O_1215,N_23615,N_22421);
nand UO_1216 (O_1216,N_23596,N_24804);
or UO_1217 (O_1217,N_20133,N_23089);
nand UO_1218 (O_1218,N_23426,N_21842);
nor UO_1219 (O_1219,N_24630,N_20479);
nor UO_1220 (O_1220,N_24948,N_21727);
and UO_1221 (O_1221,N_23851,N_22494);
nor UO_1222 (O_1222,N_22670,N_23114);
nand UO_1223 (O_1223,N_24624,N_21488);
nand UO_1224 (O_1224,N_19579,N_24177);
and UO_1225 (O_1225,N_23885,N_20675);
or UO_1226 (O_1226,N_22334,N_19466);
nand UO_1227 (O_1227,N_23494,N_22899);
and UO_1228 (O_1228,N_24733,N_23844);
nor UO_1229 (O_1229,N_23229,N_23534);
and UO_1230 (O_1230,N_21403,N_19685);
xor UO_1231 (O_1231,N_22942,N_20657);
nor UO_1232 (O_1232,N_22339,N_23535);
nand UO_1233 (O_1233,N_19096,N_21673);
nand UO_1234 (O_1234,N_22573,N_21484);
xor UO_1235 (O_1235,N_23134,N_21289);
and UO_1236 (O_1236,N_22450,N_23421);
nor UO_1237 (O_1237,N_18990,N_24475);
nor UO_1238 (O_1238,N_21801,N_23269);
and UO_1239 (O_1239,N_23839,N_22605);
nand UO_1240 (O_1240,N_21642,N_21482);
nor UO_1241 (O_1241,N_22148,N_22752);
nor UO_1242 (O_1242,N_24558,N_23827);
nand UO_1243 (O_1243,N_24234,N_19547);
and UO_1244 (O_1244,N_20053,N_21835);
or UO_1245 (O_1245,N_22116,N_22791);
xnor UO_1246 (O_1246,N_20695,N_19861);
nor UO_1247 (O_1247,N_19455,N_24126);
nor UO_1248 (O_1248,N_22995,N_24677);
nand UO_1249 (O_1249,N_19391,N_21505);
and UO_1250 (O_1250,N_24877,N_21498);
nor UO_1251 (O_1251,N_23337,N_19234);
and UO_1252 (O_1252,N_21579,N_20509);
and UO_1253 (O_1253,N_21415,N_24728);
or UO_1254 (O_1254,N_24750,N_21277);
and UO_1255 (O_1255,N_24237,N_22331);
and UO_1256 (O_1256,N_22299,N_23692);
and UO_1257 (O_1257,N_21896,N_24881);
nand UO_1258 (O_1258,N_19050,N_24547);
and UO_1259 (O_1259,N_19379,N_23701);
and UO_1260 (O_1260,N_22667,N_23678);
nand UO_1261 (O_1261,N_20435,N_23602);
nor UO_1262 (O_1262,N_22630,N_23775);
nor UO_1263 (O_1263,N_21423,N_24883);
nand UO_1264 (O_1264,N_23889,N_20721);
nor UO_1265 (O_1265,N_22222,N_21989);
and UO_1266 (O_1266,N_23139,N_23430);
or UO_1267 (O_1267,N_23059,N_24556);
nor UO_1268 (O_1268,N_22699,N_20207);
nor UO_1269 (O_1269,N_23876,N_21019);
nor UO_1270 (O_1270,N_23617,N_23713);
and UO_1271 (O_1271,N_24359,N_19439);
xor UO_1272 (O_1272,N_20968,N_19983);
nand UO_1273 (O_1273,N_20492,N_23914);
or UO_1274 (O_1274,N_19608,N_19511);
or UO_1275 (O_1275,N_21483,N_19914);
xor UO_1276 (O_1276,N_24435,N_24283);
xor UO_1277 (O_1277,N_20940,N_23005);
xnor UO_1278 (O_1278,N_23332,N_21884);
or UO_1279 (O_1279,N_20380,N_20399);
nor UO_1280 (O_1280,N_20103,N_22059);
nand UO_1281 (O_1281,N_24408,N_22051);
xor UO_1282 (O_1282,N_20600,N_19260);
xnor UO_1283 (O_1283,N_19170,N_21955);
nand UO_1284 (O_1284,N_24233,N_22084);
xnor UO_1285 (O_1285,N_23933,N_23968);
xnor UO_1286 (O_1286,N_24533,N_21786);
nand UO_1287 (O_1287,N_19895,N_18981);
nand UO_1288 (O_1288,N_21809,N_22591);
xor UO_1289 (O_1289,N_21249,N_24114);
or UO_1290 (O_1290,N_24705,N_21207);
and UO_1291 (O_1291,N_22363,N_19993);
xor UO_1292 (O_1292,N_21442,N_23750);
nor UO_1293 (O_1293,N_23395,N_20075);
nor UO_1294 (O_1294,N_22522,N_24992);
and UO_1295 (O_1295,N_20160,N_21834);
and UO_1296 (O_1296,N_21379,N_22341);
or UO_1297 (O_1297,N_24053,N_21629);
nor UO_1298 (O_1298,N_21729,N_24397);
nand UO_1299 (O_1299,N_21063,N_19173);
nand UO_1300 (O_1300,N_22454,N_22447);
or UO_1301 (O_1301,N_21042,N_23787);
xnor UO_1302 (O_1302,N_24891,N_19076);
nand UO_1303 (O_1303,N_24162,N_22140);
and UO_1304 (O_1304,N_18951,N_20568);
and UO_1305 (O_1305,N_19294,N_23785);
nor UO_1306 (O_1306,N_21774,N_18947);
nor UO_1307 (O_1307,N_24489,N_24812);
nor UO_1308 (O_1308,N_24133,N_23130);
nand UO_1309 (O_1309,N_21538,N_23758);
and UO_1310 (O_1310,N_22123,N_18991);
xor UO_1311 (O_1311,N_24541,N_21724);
and UO_1312 (O_1312,N_20981,N_24817);
or UO_1313 (O_1313,N_21618,N_23817);
and UO_1314 (O_1314,N_20621,N_20379);
nand UO_1315 (O_1315,N_23350,N_22103);
xor UO_1316 (O_1316,N_21175,N_22004);
nand UO_1317 (O_1317,N_22701,N_19544);
nand UO_1318 (O_1318,N_24382,N_22225);
or UO_1319 (O_1319,N_22892,N_23137);
nor UO_1320 (O_1320,N_19888,N_24112);
or UO_1321 (O_1321,N_24690,N_19660);
nor UO_1322 (O_1322,N_19696,N_22633);
nor UO_1323 (O_1323,N_22846,N_22169);
nor UO_1324 (O_1324,N_24550,N_21218);
and UO_1325 (O_1325,N_24571,N_20299);
nor UO_1326 (O_1326,N_19605,N_23735);
nor UO_1327 (O_1327,N_22075,N_20141);
nand UO_1328 (O_1328,N_20168,N_24748);
xnor UO_1329 (O_1329,N_20352,N_20389);
and UO_1330 (O_1330,N_21964,N_20077);
or UO_1331 (O_1331,N_23906,N_21469);
nand UO_1332 (O_1332,N_22327,N_19894);
nor UO_1333 (O_1333,N_21287,N_20224);
nor UO_1334 (O_1334,N_20860,N_23609);
xor UO_1335 (O_1335,N_24511,N_19954);
nand UO_1336 (O_1336,N_19493,N_20055);
nand UO_1337 (O_1337,N_23042,N_21353);
or UO_1338 (O_1338,N_22642,N_19951);
nor UO_1339 (O_1339,N_21598,N_19987);
or UO_1340 (O_1340,N_24235,N_22461);
nor UO_1341 (O_1341,N_22107,N_20491);
or UO_1342 (O_1342,N_19011,N_23500);
xnor UO_1343 (O_1343,N_19681,N_22789);
and UO_1344 (O_1344,N_23860,N_19746);
and UO_1345 (O_1345,N_19378,N_22814);
or UO_1346 (O_1346,N_24066,N_22358);
xor UO_1347 (O_1347,N_20761,N_22739);
nand UO_1348 (O_1348,N_21487,N_24880);
nor UO_1349 (O_1349,N_22098,N_20128);
nor UO_1350 (O_1350,N_21266,N_24134);
nor UO_1351 (O_1351,N_22175,N_24691);
and UO_1352 (O_1352,N_23022,N_24521);
xor UO_1353 (O_1353,N_22608,N_20226);
nor UO_1354 (O_1354,N_18911,N_22332);
and UO_1355 (O_1355,N_19288,N_22296);
and UO_1356 (O_1356,N_23098,N_23606);
or UO_1357 (O_1357,N_24933,N_23023);
xnor UO_1358 (O_1358,N_22512,N_23942);
xnor UO_1359 (O_1359,N_21660,N_20697);
and UO_1360 (O_1360,N_19555,N_19018);
nor UO_1361 (O_1361,N_21004,N_22272);
or UO_1362 (O_1362,N_18905,N_22245);
and UO_1363 (O_1363,N_20279,N_20671);
nor UO_1364 (O_1364,N_19468,N_24582);
nor UO_1365 (O_1365,N_21438,N_23518);
and UO_1366 (O_1366,N_21985,N_19584);
nand UO_1367 (O_1367,N_24784,N_23033);
nand UO_1368 (O_1368,N_21679,N_22744);
and UO_1369 (O_1369,N_22805,N_19960);
xor UO_1370 (O_1370,N_22138,N_23991);
nor UO_1371 (O_1371,N_22200,N_21222);
nand UO_1372 (O_1372,N_22442,N_23859);
nor UO_1373 (O_1373,N_19570,N_21074);
and UO_1374 (O_1374,N_23362,N_19389);
nand UO_1375 (O_1375,N_24645,N_19878);
or UO_1376 (O_1376,N_21284,N_23213);
xor UO_1377 (O_1377,N_22330,N_21452);
xor UO_1378 (O_1378,N_21923,N_19948);
or UO_1379 (O_1379,N_22267,N_22756);
or UO_1380 (O_1380,N_20061,N_21356);
nor UO_1381 (O_1381,N_22668,N_22176);
nand UO_1382 (O_1382,N_20332,N_24085);
nand UO_1383 (O_1383,N_18932,N_20052);
nand UO_1384 (O_1384,N_24636,N_23774);
nand UO_1385 (O_1385,N_24249,N_22677);
xnor UO_1386 (O_1386,N_22727,N_21109);
nor UO_1387 (O_1387,N_22089,N_21568);
nor UO_1388 (O_1388,N_22039,N_24600);
nor UO_1389 (O_1389,N_20896,N_21206);
xor UO_1390 (O_1390,N_24680,N_24395);
nor UO_1391 (O_1391,N_19757,N_19454);
xnor UO_1392 (O_1392,N_22247,N_22184);
nand UO_1393 (O_1393,N_20316,N_19152);
xor UO_1394 (O_1394,N_22868,N_23918);
and UO_1395 (O_1395,N_23623,N_22167);
and UO_1396 (O_1396,N_20348,N_18935);
and UO_1397 (O_1397,N_19753,N_24699);
nand UO_1398 (O_1398,N_23371,N_23575);
or UO_1399 (O_1399,N_20740,N_24631);
or UO_1400 (O_1400,N_20809,N_22950);
nor UO_1401 (O_1401,N_22142,N_21925);
and UO_1402 (O_1402,N_19768,N_23688);
nor UO_1403 (O_1403,N_23125,N_19073);
nand UO_1404 (O_1404,N_24106,N_22113);
nand UO_1405 (O_1405,N_24524,N_23277);
or UO_1406 (O_1406,N_21855,N_21507);
nand UO_1407 (O_1407,N_21942,N_20044);
nand UO_1408 (O_1408,N_22081,N_20933);
nand UO_1409 (O_1409,N_24327,N_21730);
and UO_1410 (O_1410,N_21308,N_20182);
xnor UO_1411 (O_1411,N_21066,N_21458);
nand UO_1412 (O_1412,N_21807,N_23438);
xnor UO_1413 (O_1413,N_22188,N_23976);
nand UO_1414 (O_1414,N_21607,N_21428);
and UO_1415 (O_1415,N_20475,N_20989);
xor UO_1416 (O_1416,N_19751,N_19184);
nor UO_1417 (O_1417,N_24787,N_23419);
nor UO_1418 (O_1418,N_23241,N_22029);
nor UO_1419 (O_1419,N_23986,N_22882);
nand UO_1420 (O_1420,N_22747,N_23641);
and UO_1421 (O_1421,N_21418,N_21914);
nor UO_1422 (O_1422,N_24268,N_22264);
nor UO_1423 (O_1423,N_22404,N_20646);
and UO_1424 (O_1424,N_19445,N_20369);
and UO_1425 (O_1425,N_20949,N_19552);
or UO_1426 (O_1426,N_18924,N_20579);
and UO_1427 (O_1427,N_21123,N_22889);
or UO_1428 (O_1428,N_24087,N_22136);
and UO_1429 (O_1429,N_19481,N_24510);
xnor UO_1430 (O_1430,N_20105,N_19692);
nand UO_1431 (O_1431,N_19922,N_24710);
or UO_1432 (O_1432,N_21165,N_23070);
xor UO_1433 (O_1433,N_20489,N_24366);
or UO_1434 (O_1434,N_20804,N_20049);
or UO_1435 (O_1435,N_18760,N_22487);
nand UO_1436 (O_1436,N_22697,N_24924);
nor UO_1437 (O_1437,N_22149,N_22564);
or UO_1438 (O_1438,N_23732,N_22185);
nor UO_1439 (O_1439,N_20096,N_20495);
and UO_1440 (O_1440,N_21847,N_24943);
and UO_1441 (O_1441,N_22864,N_18960);
nor UO_1442 (O_1442,N_24744,N_20070);
and UO_1443 (O_1443,N_24201,N_21624);
nor UO_1444 (O_1444,N_22218,N_18823);
xor UO_1445 (O_1445,N_22083,N_20505);
nor UO_1446 (O_1446,N_19860,N_20345);
and UO_1447 (O_1447,N_20645,N_20690);
and UO_1448 (O_1448,N_22106,N_24315);
or UO_1449 (O_1449,N_24513,N_21606);
or UO_1450 (O_1450,N_19261,N_19889);
or UO_1451 (O_1451,N_22422,N_24818);
nor UO_1452 (O_1452,N_18878,N_21065);
nand UO_1453 (O_1453,N_20322,N_23947);
and UO_1454 (O_1454,N_23731,N_19397);
xnor UO_1455 (O_1455,N_18794,N_20420);
and UO_1456 (O_1456,N_20640,N_22929);
or UO_1457 (O_1457,N_19853,N_23815);
nand UO_1458 (O_1458,N_22631,N_24998);
nand UO_1459 (O_1459,N_20277,N_22008);
nand UO_1460 (O_1460,N_20626,N_24578);
xnor UO_1461 (O_1461,N_22032,N_21178);
nand UO_1462 (O_1462,N_19514,N_20426);
nand UO_1463 (O_1463,N_20891,N_21789);
nor UO_1464 (O_1464,N_23685,N_23922);
nand UO_1465 (O_1465,N_20022,N_23782);
and UO_1466 (O_1466,N_22986,N_18945);
nor UO_1467 (O_1467,N_21858,N_21112);
and UO_1468 (O_1468,N_22907,N_22288);
nor UO_1469 (O_1469,N_19122,N_22509);
and UO_1470 (O_1470,N_23064,N_22066);
xnor UO_1471 (O_1471,N_23944,N_21286);
xor UO_1472 (O_1472,N_22857,N_24944);
nor UO_1473 (O_1473,N_19033,N_20185);
nor UO_1474 (O_1474,N_24501,N_22300);
nor UO_1475 (O_1475,N_24840,N_21992);
and UO_1476 (O_1476,N_23324,N_19331);
nand UO_1477 (O_1477,N_21757,N_24343);
xor UO_1478 (O_1478,N_19210,N_22276);
xor UO_1479 (O_1479,N_19744,N_20984);
nor UO_1480 (O_1480,N_19615,N_22319);
xor UO_1481 (O_1481,N_18880,N_22705);
or UO_1482 (O_1482,N_23835,N_20807);
xor UO_1483 (O_1483,N_22821,N_24704);
nor UO_1484 (O_1484,N_18972,N_19470);
xor UO_1485 (O_1485,N_18959,N_22546);
nor UO_1486 (O_1486,N_20367,N_20913);
xor UO_1487 (O_1487,N_19127,N_21735);
nand UO_1488 (O_1488,N_24786,N_18995);
and UO_1489 (O_1489,N_19224,N_23099);
nor UO_1490 (O_1490,N_19873,N_24332);
nand UO_1491 (O_1491,N_20591,N_19885);
nand UO_1492 (O_1492,N_22180,N_19192);
nand UO_1493 (O_1493,N_19736,N_22120);
xor UO_1494 (O_1494,N_22021,N_23892);
and UO_1495 (O_1495,N_21097,N_22501);
or UO_1496 (O_1496,N_23165,N_18800);
and UO_1497 (O_1497,N_23414,N_19489);
nand UO_1498 (O_1498,N_20730,N_21545);
nand UO_1499 (O_1499,N_23832,N_21811);
nand UO_1500 (O_1500,N_19828,N_24814);
or UO_1501 (O_1501,N_21943,N_20539);
nand UO_1502 (O_1502,N_24154,N_19926);
and UO_1503 (O_1503,N_21017,N_19664);
xor UO_1504 (O_1504,N_24607,N_19086);
xor UO_1505 (O_1505,N_20454,N_20866);
and UO_1506 (O_1506,N_23479,N_23597);
nand UO_1507 (O_1507,N_23239,N_21685);
nor UO_1508 (O_1508,N_19764,N_24051);
nand UO_1509 (O_1509,N_24870,N_24054);
nand UO_1510 (O_1510,N_20441,N_23366);
nand UO_1511 (O_1511,N_21425,N_23186);
nand UO_1512 (O_1512,N_23675,N_23329);
nand UO_1513 (O_1513,N_23319,N_21179);
or UO_1514 (O_1514,N_21902,N_24362);
or UO_1515 (O_1515,N_20983,N_18937);
or UO_1516 (O_1516,N_23364,N_19065);
nor UO_1517 (O_1517,N_22369,N_24199);
nor UO_1518 (O_1518,N_24346,N_22070);
nand UO_1519 (O_1519,N_21657,N_24494);
nand UO_1520 (O_1520,N_20907,N_19290);
nand UO_1521 (O_1521,N_24842,N_21590);
nand UO_1522 (O_1522,N_24643,N_22928);
or UO_1523 (O_1523,N_24663,N_20448);
nor UO_1524 (O_1524,N_21473,N_20711);
or UO_1525 (O_1525,N_19293,N_22063);
xor UO_1526 (O_1526,N_24229,N_22867);
or UO_1527 (O_1527,N_23862,N_22456);
nor UO_1528 (O_1528,N_19253,N_21383);
nor UO_1529 (O_1529,N_20429,N_19677);
xnor UO_1530 (O_1530,N_20817,N_20169);
and UO_1531 (O_1531,N_23214,N_21556);
or UO_1532 (O_1532,N_23420,N_19008);
nor UO_1533 (O_1533,N_24759,N_23943);
xor UO_1534 (O_1534,N_22360,N_21754);
nand UO_1535 (O_1535,N_22831,N_24307);
and UO_1536 (O_1536,N_19603,N_23900);
and UO_1537 (O_1537,N_24165,N_22627);
nor UO_1538 (O_1538,N_22617,N_24937);
and UO_1539 (O_1539,N_22776,N_23838);
and UO_1540 (O_1540,N_19771,N_20868);
nor UO_1541 (O_1541,N_21188,N_21348);
or UO_1542 (O_1542,N_19808,N_24658);
xnor UO_1543 (O_1543,N_19313,N_22312);
nand UO_1544 (O_1544,N_20442,N_19989);
nor UO_1545 (O_1545,N_20302,N_19059);
and UO_1546 (O_1546,N_24755,N_23215);
or UO_1547 (O_1547,N_21319,N_22702);
nand UO_1548 (O_1548,N_19786,N_21352);
and UO_1549 (O_1549,N_20583,N_22601);
and UO_1550 (O_1550,N_23970,N_18787);
xnor UO_1551 (O_1551,N_23174,N_24802);
nor UO_1552 (O_1552,N_24963,N_18828);
xor UO_1553 (O_1553,N_19363,N_21457);
nor UO_1554 (O_1554,N_24243,N_24400);
and UO_1555 (O_1555,N_23638,N_21944);
and UO_1556 (O_1556,N_24753,N_22910);
nor UO_1557 (O_1557,N_22492,N_20673);
nor UO_1558 (O_1558,N_23258,N_22134);
xor UO_1559 (O_1559,N_21194,N_22829);
or UO_1560 (O_1560,N_19158,N_19620);
and UO_1561 (O_1561,N_24724,N_21265);
and UO_1562 (O_1562,N_23443,N_20347);
nor UO_1563 (O_1563,N_19304,N_20750);
or UO_1564 (O_1564,N_24443,N_20289);
nor UO_1565 (O_1565,N_19479,N_21911);
or UO_1566 (O_1566,N_18783,N_23266);
xnor UO_1567 (O_1567,N_23508,N_20929);
and UO_1568 (O_1568,N_22516,N_21653);
nor UO_1569 (O_1569,N_21739,N_21872);
and UO_1570 (O_1570,N_20508,N_23031);
nor UO_1571 (O_1571,N_19169,N_21766);
and UO_1572 (O_1572,N_20156,N_21197);
xor UO_1573 (O_1573,N_19787,N_22689);
xor UO_1574 (O_1574,N_21837,N_23416);
nor UO_1575 (O_1575,N_24095,N_21154);
xnor UO_1576 (O_1576,N_22840,N_19513);
or UO_1577 (O_1577,N_23977,N_22057);
or UO_1578 (O_1578,N_20476,N_21171);
xnor UO_1579 (O_1579,N_20456,N_22472);
and UO_1580 (O_1580,N_20617,N_20215);
or UO_1581 (O_1581,N_20114,N_22722);
xor UO_1582 (O_1582,N_19289,N_24170);
and UO_1583 (O_1583,N_19825,N_20863);
or UO_1584 (O_1584,N_21734,N_23710);
and UO_1585 (O_1585,N_19032,N_22874);
or UO_1586 (O_1586,N_22017,N_24714);
nand UO_1587 (O_1587,N_22742,N_23463);
or UO_1588 (O_1588,N_21938,N_23905);
nor UO_1589 (O_1589,N_23263,N_22659);
nand UO_1590 (O_1590,N_22855,N_22056);
or UO_1591 (O_1591,N_21378,N_24740);
nand UO_1592 (O_1592,N_20084,N_19478);
xnor UO_1593 (O_1593,N_22750,N_21045);
and UO_1594 (O_1594,N_19361,N_22787);
xnor UO_1595 (O_1595,N_24441,N_19056);
xnor UO_1596 (O_1596,N_22637,N_21627);
and UO_1597 (O_1597,N_20852,N_19565);
nor UO_1598 (O_1598,N_19942,N_22871);
and UO_1599 (O_1599,N_23841,N_22238);
xor UO_1600 (O_1600,N_24930,N_23857);
nand UO_1601 (O_1601,N_22124,N_23935);
or UO_1602 (O_1602,N_18763,N_19399);
xnor UO_1603 (O_1603,N_21293,N_20970);
and UO_1604 (O_1604,N_22610,N_22908);
nand UO_1605 (O_1605,N_19882,N_20918);
nor UO_1606 (O_1606,N_21281,N_21046);
xor UO_1607 (O_1607,N_23060,N_20597);
and UO_1608 (O_1608,N_21357,N_20328);
nand UO_1609 (O_1609,N_20835,N_24751);
xor UO_1610 (O_1610,N_24635,N_24099);
xnor UO_1611 (O_1611,N_22661,N_24707);
and UO_1612 (O_1612,N_19415,N_24429);
or UO_1613 (O_1613,N_20638,N_24002);
nor UO_1614 (O_1614,N_24564,N_24345);
or UO_1615 (O_1615,N_21387,N_19654);
and UO_1616 (O_1616,N_23331,N_22532);
and UO_1617 (O_1617,N_22062,N_19624);
nor UO_1618 (O_1618,N_22209,N_20975);
nand UO_1619 (O_1619,N_23288,N_23184);
or UO_1620 (O_1620,N_22870,N_19467);
nand UO_1621 (O_1621,N_23491,N_23303);
nor UO_1622 (O_1622,N_22938,N_24542);
and UO_1623 (O_1623,N_20784,N_24440);
xnor UO_1624 (O_1624,N_20862,N_24252);
xor UO_1625 (O_1625,N_23338,N_19588);
nand UO_1626 (O_1626,N_19418,N_19934);
xnor UO_1627 (O_1627,N_24912,N_24369);
xor UO_1628 (O_1628,N_23221,N_20871);
xnor UO_1629 (O_1629,N_20515,N_21377);
xnor UO_1630 (O_1630,N_20561,N_20263);
xnor UO_1631 (O_1631,N_20024,N_21941);
nand UO_1632 (O_1632,N_23167,N_22018);
xor UO_1633 (O_1633,N_19725,N_23111);
and UO_1634 (O_1634,N_19387,N_24585);
or UO_1635 (O_1635,N_19254,N_19137);
xnor UO_1636 (O_1636,N_20936,N_21785);
or UO_1637 (O_1637,N_22240,N_19742);
nor UO_1638 (O_1638,N_19952,N_24771);
nand UO_1639 (O_1639,N_22580,N_22903);
xor UO_1640 (O_1640,N_21351,N_22025);
nor UO_1641 (O_1641,N_22060,N_21342);
or UO_1642 (O_1642,N_21740,N_23880);
or UO_1643 (O_1643,N_23805,N_22541);
nand UO_1644 (O_1644,N_19218,N_22480);
or UO_1645 (O_1645,N_22875,N_23670);
nand UO_1646 (O_1646,N_20488,N_24529);
or UO_1647 (O_1647,N_23789,N_23672);
xnor UO_1648 (O_1648,N_22239,N_18928);
nand UO_1649 (O_1649,N_19635,N_19206);
and UO_1650 (O_1650,N_22423,N_23581);
nand UO_1651 (O_1651,N_23622,N_20394);
and UO_1652 (O_1652,N_24803,N_20497);
xnor UO_1653 (O_1653,N_21429,N_19818);
xnor UO_1654 (O_1654,N_18799,N_23025);
or UO_1655 (O_1655,N_22445,N_22444);
nand UO_1656 (O_1656,N_19273,N_22806);
nand UO_1657 (O_1657,N_23667,N_23330);
nand UO_1658 (O_1658,N_19933,N_21779);
nand UO_1659 (O_1659,N_19504,N_24027);
xnor UO_1660 (O_1660,N_21385,N_20407);
nor UO_1661 (O_1661,N_20735,N_19501);
or UO_1662 (O_1662,N_24718,N_24579);
or UO_1663 (O_1663,N_23196,N_22590);
nand UO_1664 (O_1664,N_24476,N_23882);
and UO_1665 (O_1665,N_22946,N_19586);
xnor UO_1666 (O_1666,N_20678,N_18859);
or UO_1667 (O_1667,N_23244,N_24479);
xnor UO_1668 (O_1668,N_22317,N_20164);
nor UO_1669 (O_1669,N_20619,N_20650);
and UO_1670 (O_1670,N_20771,N_21871);
nand UO_1671 (O_1671,N_19690,N_22373);
nor UO_1672 (O_1672,N_19969,N_20928);
nor UO_1673 (O_1673,N_20905,N_23291);
or UO_1674 (O_1674,N_23792,N_20391);
nand UO_1675 (O_1675,N_20050,N_20065);
and UO_1676 (O_1676,N_22991,N_24984);
and UO_1677 (O_1677,N_21710,N_19941);
nor UO_1678 (O_1678,N_22508,N_20739);
and UO_1679 (O_1679,N_23019,N_20305);
and UO_1680 (O_1680,N_23153,N_21115);
nand UO_1681 (O_1681,N_19678,N_22203);
nor UO_1682 (O_1682,N_22014,N_24664);
and UO_1683 (O_1683,N_23728,N_18784);
or UO_1684 (O_1684,N_20550,N_24821);
xnor UO_1685 (O_1685,N_19044,N_21843);
nand UO_1686 (O_1686,N_19072,N_22475);
and UO_1687 (O_1687,N_19434,N_19060);
and UO_1688 (O_1688,N_23497,N_21683);
nand UO_1689 (O_1689,N_22160,N_24248);
nand UO_1690 (O_1690,N_19724,N_24932);
xor UO_1691 (O_1691,N_22271,N_19502);
and UO_1692 (O_1692,N_24205,N_20368);
nand UO_1693 (O_1693,N_21857,N_22359);
and UO_1694 (O_1694,N_21868,N_22696);
nor UO_1695 (O_1695,N_19886,N_20381);
or UO_1696 (O_1696,N_22281,N_20039);
nor UO_1697 (O_1697,N_18978,N_19790);
nor UO_1698 (O_1698,N_19319,N_18805);
and UO_1699 (O_1699,N_22322,N_19812);
nand UO_1700 (O_1700,N_21644,N_20064);
or UO_1701 (O_1701,N_19334,N_21332);
and UO_1702 (O_1702,N_23211,N_21124);
and UO_1703 (O_1703,N_21214,N_22769);
nand UO_1704 (O_1704,N_21440,N_19739);
nand UO_1705 (O_1705,N_18889,N_24845);
nor UO_1706 (O_1706,N_22505,N_23987);
nor UO_1707 (O_1707,N_20398,N_20246);
and UO_1708 (O_1708,N_24244,N_22877);
or UO_1709 (O_1709,N_22992,N_23631);
nand UO_1710 (O_1710,N_24135,N_19573);
nor UO_1711 (O_1711,N_23238,N_19243);
nor UO_1712 (O_1712,N_20598,N_23286);
nor UO_1713 (O_1713,N_23149,N_22959);
xor UO_1714 (O_1714,N_22163,N_24232);
xnor UO_1715 (O_1715,N_21023,N_24736);
xor UO_1716 (O_1716,N_21268,N_20080);
xnor UO_1717 (O_1717,N_18809,N_20559);
and UO_1718 (O_1718,N_20980,N_24324);
and UO_1719 (O_1719,N_23513,N_22252);
xnor UO_1720 (O_1720,N_20033,N_24032);
or UO_1721 (O_1721,N_20630,N_18753);
and UO_1722 (O_1722,N_19606,N_19761);
or UO_1723 (O_1723,N_24505,N_22749);
nor UO_1724 (O_1724,N_19842,N_19365);
or UO_1725 (O_1725,N_24647,N_19045);
or UO_1726 (O_1726,N_21612,N_21697);
and UO_1727 (O_1727,N_23000,N_21318);
and UO_1728 (O_1728,N_23173,N_24781);
and UO_1729 (O_1729,N_20587,N_22651);
or UO_1730 (O_1730,N_20887,N_23971);
xnor UO_1731 (O_1731,N_23150,N_20362);
and UO_1732 (O_1732,N_19966,N_22737);
xor UO_1733 (O_1733,N_20201,N_20029);
or UO_1734 (O_1734,N_19302,N_24284);
nand UO_1735 (O_1735,N_19728,N_24868);
or UO_1736 (O_1736,N_21950,N_22325);
nor UO_1737 (O_1737,N_19490,N_21665);
and UO_1738 (O_1738,N_19237,N_24667);
and UO_1739 (O_1739,N_22220,N_23843);
nand UO_1740 (O_1740,N_21005,N_24866);
and UO_1741 (O_1741,N_23043,N_19027);
and UO_1742 (O_1742,N_22596,N_20249);
or UO_1743 (O_1743,N_18894,N_22579);
nor UO_1744 (O_1744,N_19735,N_18792);
nand UO_1745 (O_1745,N_22379,N_24762);
xnor UO_1746 (O_1746,N_18892,N_20719);
nor UO_1747 (O_1747,N_21376,N_20078);
and UO_1748 (O_1748,N_24560,N_18879);
and UO_1749 (O_1749,N_20552,N_19832);
or UO_1750 (O_1750,N_22820,N_19241);
xor UO_1751 (O_1751,N_19007,N_23250);
and UO_1752 (O_1752,N_23895,N_20094);
xor UO_1753 (O_1753,N_21362,N_19848);
xor UO_1754 (O_1754,N_22504,N_24716);
or UO_1755 (O_1755,N_21084,N_21565);
nand UO_1756 (O_1756,N_20977,N_22556);
nand UO_1757 (O_1757,N_18989,N_23492);
nor UO_1758 (O_1758,N_21329,N_22310);
nor UO_1759 (O_1759,N_20129,N_18858);
or UO_1760 (O_1760,N_20028,N_22320);
nor UO_1761 (O_1761,N_24445,N_22989);
and UO_1762 (O_1762,N_20281,N_19174);
or UO_1763 (O_1763,N_18942,N_23644);
xnor UO_1764 (O_1764,N_20718,N_22182);
and UO_1765 (O_1765,N_21934,N_19425);
xor UO_1766 (O_1766,N_24301,N_19142);
nor UO_1767 (O_1767,N_22530,N_20317);
nand UO_1768 (O_1768,N_21409,N_19335);
xor UO_1769 (O_1769,N_20596,N_21494);
nand UO_1770 (O_1770,N_21317,N_23786);
and UO_1771 (O_1771,N_19585,N_22869);
nor UO_1772 (O_1772,N_19426,N_23501);
xnor UO_1773 (O_1773,N_22465,N_20958);
and UO_1774 (O_1774,N_20819,N_19884);
and UO_1775 (O_1775,N_23875,N_19639);
or UO_1776 (O_1776,N_24137,N_19574);
nor UO_1777 (O_1777,N_20417,N_23878);
or UO_1778 (O_1778,N_24091,N_21993);
nand UO_1779 (O_1779,N_20112,N_20828);
or UO_1780 (O_1780,N_24077,N_22144);
and UO_1781 (O_1781,N_21790,N_20147);
nand UO_1782 (O_1782,N_24384,N_19985);
xor UO_1783 (O_1783,N_22937,N_24890);
and UO_1784 (O_1784,N_22690,N_19021);
nor UO_1785 (O_1785,N_24747,N_21968);
or UO_1786 (O_1786,N_23825,N_19995);
xor UO_1787 (O_1787,N_24204,N_19741);
or UO_1788 (O_1788,N_23119,N_20972);
or UO_1789 (O_1789,N_21471,N_22298);
xor UO_1790 (O_1790,N_24447,N_23308);
nor UO_1791 (O_1791,N_21010,N_24311);
xor UO_1792 (O_1792,N_23587,N_23948);
and UO_1793 (O_1793,N_20872,N_20520);
or UO_1794 (O_1794,N_20832,N_19352);
or UO_1795 (O_1795,N_22473,N_20810);
xnor UO_1796 (O_1796,N_19557,N_23240);
and UO_1797 (O_1797,N_22187,N_23967);
nor UO_1798 (O_1798,N_23037,N_19846);
xor UO_1799 (O_1799,N_19910,N_23344);
or UO_1800 (O_1800,N_21122,N_20481);
or UO_1801 (O_1801,N_22603,N_20408);
nand UO_1802 (O_1802,N_19449,N_22694);
nor UO_1803 (O_1803,N_19946,N_18956);
or UO_1804 (O_1804,N_21059,N_20716);
and UO_1805 (O_1805,N_22800,N_18772);
and UO_1806 (O_1806,N_18901,N_24076);
and UO_1807 (O_1807,N_21566,N_21529);
or UO_1808 (O_1808,N_23899,N_19684);
nand UO_1809 (O_1809,N_23044,N_19543);
nand UO_1810 (O_1810,N_24497,N_23829);
xor UO_1811 (O_1811,N_23393,N_22204);
and UO_1812 (O_1812,N_24219,N_22351);
nand UO_1813 (O_1813,N_20815,N_19317);
xor UO_1814 (O_1814,N_21283,N_24187);
nand UO_1815 (O_1815,N_24514,N_19440);
and UO_1816 (O_1816,N_19396,N_22227);
or UO_1817 (O_1817,N_20877,N_21104);
nor UO_1818 (O_1818,N_19267,N_20870);
or UO_1819 (O_1819,N_19430,N_21814);
xnor UO_1820 (O_1820,N_23551,N_22957);
nand UO_1821 (O_1821,N_24480,N_23820);
or UO_1822 (O_1822,N_21960,N_23368);
nand UO_1823 (O_1823,N_19183,N_22482);
or UO_1824 (O_1824,N_23093,N_21031);
nor UO_1825 (O_1825,N_22983,N_22657);
and UO_1826 (O_1826,N_24144,N_22799);
xnor UO_1827 (O_1827,N_20285,N_19040);
nor UO_1828 (O_1828,N_24693,N_24403);
or UO_1829 (O_1829,N_24386,N_24660);
or UO_1830 (O_1830,N_21386,N_19416);
nor UO_1831 (O_1831,N_22916,N_20746);
nand UO_1832 (O_1832,N_22824,N_24626);
and UO_1833 (O_1833,N_23684,N_18804);
and UO_1834 (O_1834,N_24764,N_23177);
and UO_1835 (O_1835,N_22782,N_24039);
and UO_1836 (O_1836,N_21537,N_19199);
nor UO_1837 (O_1837,N_23315,N_24276);
nand UO_1838 (O_1838,N_24695,N_19792);
or UO_1839 (O_1839,N_21278,N_24086);
or UO_1840 (O_1840,N_24034,N_22217);
or UO_1841 (O_1841,N_24088,N_19977);
xor UO_1842 (O_1842,N_24659,N_19562);
xnor UO_1843 (O_1843,N_23469,N_22876);
nor UO_1844 (O_1844,N_23466,N_21225);
nand UO_1845 (O_1845,N_19003,N_24976);
xnor UO_1846 (O_1846,N_21044,N_19733);
and UO_1847 (O_1847,N_23705,N_21172);
nor UO_1848 (O_1848,N_19747,N_24189);
xor UO_1849 (O_1849,N_22536,N_23659);
and UO_1850 (O_1850,N_24349,N_21322);
nand UO_1851 (O_1851,N_23448,N_21176);
and UO_1852 (O_1852,N_24145,N_20947);
and UO_1853 (O_1853,N_22794,N_20015);
nand UO_1854 (O_1854,N_23083,N_22198);
xor UO_1855 (O_1855,N_24849,N_20806);
nand UO_1856 (O_1856,N_22873,N_22912);
and UO_1857 (O_1857,N_21572,N_19408);
nor UO_1858 (O_1858,N_22162,N_21113);
and UO_1859 (O_1859,N_21291,N_20656);
xnor UO_1860 (O_1860,N_20987,N_23777);
or UO_1861 (O_1861,N_23528,N_21794);
xnor UO_1862 (O_1862,N_20931,N_20676);
nand UO_1863 (O_1863,N_24221,N_19108);
nor UO_1864 (O_1864,N_24625,N_24195);
xnor UO_1865 (O_1865,N_19136,N_18994);
or UO_1866 (O_1866,N_22808,N_22526);
nor UO_1867 (O_1867,N_18963,N_23101);
or UO_1868 (O_1868,N_21534,N_22048);
or UO_1869 (O_1869,N_23351,N_19875);
and UO_1870 (O_1870,N_19655,N_20795);
nor UO_1871 (O_1871,N_22055,N_23437);
xor UO_1872 (O_1872,N_19625,N_23509);
nand UO_1873 (O_1873,N_23628,N_19308);
nor UO_1874 (O_1874,N_23654,N_21041);
or UO_1875 (O_1875,N_20487,N_24670);
and UO_1876 (O_1876,N_23464,N_21721);
and UO_1877 (O_1877,N_19476,N_24796);
nand UO_1878 (O_1878,N_22147,N_21192);
xnor UO_1879 (O_1879,N_22745,N_24005);
or UO_1880 (O_1880,N_19990,N_21825);
and UO_1881 (O_1881,N_19263,N_21694);
nor UO_1882 (O_1882,N_19103,N_22534);
nor UO_1883 (O_1883,N_21620,N_21349);
nor UO_1884 (O_1884,N_21237,N_22819);
and UO_1885 (O_1885,N_19553,N_21215);
or UO_1886 (O_1886,N_22016,N_21927);
nor UO_1887 (O_1887,N_22349,N_21667);
and UO_1888 (O_1888,N_19283,N_23236);
xnor UO_1889 (O_1889,N_23394,N_19619);
and UO_1890 (O_1890,N_19110,N_20413);
xor UO_1891 (O_1891,N_24230,N_19752);
and UO_1892 (O_1892,N_22926,N_19829);
and UO_1893 (O_1893,N_24952,N_19657);
or UO_1894 (O_1894,N_22555,N_21139);
nand UO_1895 (O_1895,N_21508,N_20523);
and UO_1896 (O_1896,N_19992,N_24935);
and UO_1897 (O_1897,N_19204,N_24756);
nor UO_1898 (O_1898,N_21324,N_23651);
nor UO_1899 (O_1899,N_20219,N_23293);
nand UO_1900 (O_1900,N_23054,N_21183);
nor UO_1901 (O_1901,N_24862,N_24779);
nor UO_1902 (O_1902,N_22137,N_22347);
nor UO_1903 (O_1903,N_19080,N_20242);
nor UO_1904 (O_1904,N_20250,N_24269);
xnor UO_1905 (O_1905,N_23446,N_19996);
and UO_1906 (O_1906,N_19671,N_23110);
xnor UO_1907 (O_1907,N_24859,N_24411);
nand UO_1908 (O_1908,N_22452,N_21591);
nand UO_1909 (O_1909,N_20031,N_21420);
xor UO_1910 (O_1910,N_24006,N_19358);
and UO_1911 (O_1911,N_18910,N_21338);
and UO_1912 (O_1912,N_21034,N_21212);
and UO_1913 (O_1913,N_21738,N_20189);
and UO_1914 (O_1914,N_19711,N_22058);
xnor UO_1915 (O_1915,N_24884,N_20749);
or UO_1916 (O_1916,N_24813,N_19131);
and UO_1917 (O_1917,N_23360,N_22497);
xnor UO_1918 (O_1918,N_24401,N_19328);
nand UO_1919 (O_1919,N_19217,N_21304);
or UO_1920 (O_1920,N_23084,N_20079);
or UO_1921 (O_1921,N_19974,N_22847);
or UO_1922 (O_1922,N_22891,N_22214);
or UO_1923 (O_1923,N_24848,N_24317);
and UO_1924 (O_1924,N_21962,N_21717);
or UO_1925 (O_1925,N_23388,N_22827);
nor UO_1926 (O_1926,N_20331,N_19537);
xnor UO_1927 (O_1927,N_24517,N_24052);
nand UO_1928 (O_1928,N_21886,N_22213);
or UO_1929 (O_1929,N_23579,N_22966);
nand UO_1930 (O_1930,N_21079,N_22792);
xor UO_1931 (O_1931,N_21474,N_23477);
xnor UO_1932 (O_1932,N_24157,N_24122);
nor UO_1933 (O_1933,N_22053,N_19596);
xor UO_1934 (O_1934,N_22622,N_19285);
xor UO_1935 (O_1935,N_19781,N_22333);
or UO_1936 (O_1936,N_24371,N_20130);
or UO_1937 (O_1937,N_24251,N_20484);
and UO_1938 (O_1938,N_19348,N_20326);
and UO_1939 (O_1939,N_24788,N_18871);
and UO_1940 (O_1940,N_20776,N_19077);
and UO_1941 (O_1941,N_20516,N_21638);
or UO_1942 (O_1942,N_24512,N_22947);
xnor UO_1943 (O_1943,N_21103,N_24422);
nand UO_1944 (O_1944,N_20538,N_19075);
and UO_1945 (O_1945,N_24310,N_22731);
nand UO_1946 (O_1946,N_21168,N_21800);
nand UO_1947 (O_1947,N_24576,N_19532);
and UO_1948 (O_1948,N_20748,N_24994);
nand UO_1949 (O_1949,N_23996,N_20157);
or UO_1950 (O_1950,N_23348,N_20915);
nor UO_1951 (O_1951,N_22636,N_21226);
and UO_1952 (O_1952,N_22844,N_23556);
nand UO_1953 (O_1953,N_24561,N_22640);
or UO_1954 (O_1954,N_21594,N_20355);
nand UO_1955 (O_1955,N_20869,N_23224);
nand UO_1956 (O_1956,N_20652,N_24983);
and UO_1957 (O_1957,N_19997,N_23952);
or UO_1958 (O_1958,N_21551,N_21056);
nor UO_1959 (O_1959,N_19052,N_19597);
nand UO_1960 (O_1960,N_22707,N_21035);
and UO_1961 (O_1961,N_23024,N_19051);
nor UO_1962 (O_1962,N_24544,N_21467);
xnor UO_1963 (O_1963,N_23452,N_21937);
and UO_1964 (O_1964,N_18822,N_19851);
nand UO_1965 (O_1965,N_24552,N_19291);
nor UO_1966 (O_1966,N_22114,N_23697);
and UO_1967 (O_1967,N_21048,N_22513);
and UO_1968 (O_1968,N_19482,N_19509);
and UO_1969 (O_1969,N_19662,N_24882);
nand UO_1970 (O_1970,N_20658,N_22389);
and UO_1971 (O_1971,N_24894,N_18768);
nor UO_1972 (O_1972,N_19160,N_22195);
xor UO_1973 (O_1973,N_23283,N_18754);
and UO_1974 (O_1974,N_21647,N_21086);
xnor UO_1975 (O_1975,N_22817,N_19836);
or UO_1976 (O_1976,N_22458,N_24117);
or UO_1977 (O_1977,N_19364,N_20339);
nor UO_1978 (O_1978,N_20525,N_23591);
xor UO_1979 (O_1979,N_23711,N_23502);
and UO_1980 (O_1980,N_21430,N_20139);
and UO_1981 (O_1981,N_22023,N_18993);
nand UO_1982 (O_1982,N_20781,N_23621);
nand UO_1983 (O_1983,N_19371,N_19257);
nand UO_1984 (O_1984,N_20901,N_23802);
or UO_1985 (O_1985,N_24655,N_19577);
xor UO_1986 (O_1986,N_23161,N_21164);
nor UO_1987 (O_1987,N_22399,N_21136);
nand UO_1988 (O_1988,N_21142,N_23131);
nor UO_1989 (O_1989,N_19043,N_24406);
nand UO_1990 (O_1990,N_21476,N_19610);
nand UO_1991 (O_1991,N_18785,N_23852);
xnor UO_1992 (O_1992,N_24414,N_20040);
xnor UO_1993 (O_1993,N_24596,N_21584);
or UO_1994 (O_1994,N_22366,N_22152);
or UO_1995 (O_1995,N_24374,N_18870);
xor UO_1996 (O_1996,N_24485,N_23930);
and UO_1997 (O_1997,N_22700,N_19203);
xnor UO_1998 (O_1998,N_19067,N_20507);
and UO_1999 (O_1999,N_24142,N_20132);
nand UO_2000 (O_2000,N_19132,N_19423);
xnor UO_2001 (O_2001,N_19612,N_23449);
nand UO_2002 (O_2002,N_24823,N_21758);
and UO_2003 (O_2003,N_23267,N_24954);
and UO_2004 (O_2004,N_20889,N_20820);
or UO_2005 (O_2005,N_19171,N_21692);
nor UO_2006 (O_2006,N_22743,N_24745);
xor UO_2007 (O_2007,N_20223,N_22350);
nand UO_2008 (O_2008,N_20248,N_21723);
or UO_2009 (O_2009,N_20999,N_19019);
nand UO_2010 (O_2010,N_21347,N_18864);
nand UO_2011 (O_2011,N_19650,N_19760);
or UO_2012 (O_2012,N_22223,N_21689);
or UO_2013 (O_2013,N_23745,N_23830);
xnor UO_2014 (O_2014,N_22507,N_23512);
and UO_2015 (O_2015,N_20608,N_21477);
and UO_2016 (O_2016,N_21092,N_23520);
and UO_2017 (O_2017,N_19392,N_21515);
nor UO_2018 (O_2018,N_23251,N_22687);
xnor UO_2019 (O_2019,N_21311,N_24972);
and UO_2020 (O_2020,N_23195,N_21887);
nor UO_2021 (O_2021,N_20360,N_20469);
nor UO_2022 (O_2022,N_23588,N_21116);
nor UO_2023 (O_2023,N_22523,N_23798);
and UO_2024 (O_2024,N_24261,N_23912);
nand UO_2025 (O_2025,N_22726,N_22843);
or UO_2026 (O_2026,N_23769,N_24203);
or UO_2027 (O_2027,N_22158,N_22132);
and UO_2028 (O_2028,N_21290,N_18929);
or UO_2029 (O_2029,N_23770,N_24321);
and UO_2030 (O_2030,N_23867,N_19525);
xnor UO_2031 (O_2031,N_21478,N_21325);
or UO_2032 (O_2032,N_21759,N_21575);
xor UO_2033 (O_2033,N_19767,N_20423);
nand UO_2034 (O_2034,N_24164,N_22558);
xnor UO_2035 (O_2035,N_24539,N_22437);
nor UO_2036 (O_2036,N_20654,N_22002);
and UO_2037 (O_2037,N_22672,N_21210);
nand UO_2038 (O_2038,N_20919,N_23916);
xnor UO_2039 (O_2039,N_23035,N_20534);
or UO_2040 (O_2040,N_23347,N_23381);
xnor UO_2041 (O_2041,N_22221,N_24538);
nand UO_2042 (O_2042,N_19500,N_24629);
and UO_2043 (O_2043,N_19246,N_21454);
xnor UO_2044 (O_2044,N_22940,N_22898);
nor UO_2045 (O_2045,N_20468,N_21726);
nor UO_2046 (O_2046,N_20253,N_24236);
xor UO_2047 (O_2047,N_21675,N_22438);
or UO_2048 (O_2048,N_18915,N_22593);
or UO_2049 (O_2049,N_23166,N_22368);
or UO_2050 (O_2050,N_21163,N_24583);
xnor UO_2051 (O_2051,N_24035,N_21461);
nor UO_2052 (O_2052,N_24587,N_19533);
and UO_2053 (O_2053,N_20737,N_24295);
or UO_2054 (O_2054,N_20365,N_19124);
nor UO_2055 (O_2055,N_21728,N_19727);
or UO_2056 (O_2056,N_19346,N_23404);
nor UO_2057 (O_2057,N_24810,N_18771);
xnor UO_2058 (O_2058,N_19647,N_20245);
nor UO_2059 (O_2059,N_20857,N_20286);
and UO_2060 (O_2060,N_23831,N_20298);
or UO_2061 (O_2061,N_20310,N_22313);
or UO_2062 (O_2062,N_19020,N_19656);
nor UO_2063 (O_2063,N_23569,N_22647);
nor UO_2064 (O_2064,N_23507,N_19902);
xnor UO_2065 (O_2065,N_21307,N_24127);
nand UO_2066 (O_2066,N_19567,N_19510);
nor UO_2067 (O_2067,N_22338,N_21155);
or UO_2068 (O_2068,N_23980,N_19870);
nand UO_2069 (O_2069,N_23403,N_19549);
nand UO_2070 (O_2070,N_20225,N_22443);
and UO_2071 (O_2071,N_23972,N_22736);
or UO_2072 (O_2072,N_24537,N_19931);
nand UO_2073 (O_2073,N_22476,N_22357);
and UO_2074 (O_2074,N_23733,N_20017);
nor UO_2075 (O_2075,N_23326,N_24627);
xor UO_2076 (O_2076,N_21026,N_22414);
nor UO_2077 (O_2077,N_18967,N_21861);
and UO_2078 (O_2078,N_23717,N_21173);
or UO_2079 (O_2079,N_21282,N_23704);
nand UO_2080 (O_2080,N_20549,N_20349);
xor UO_2081 (O_2081,N_21141,N_20220);
or UO_2082 (O_2082,N_18779,N_22765);
xnor UO_2083 (O_2083,N_19404,N_21263);
or UO_2084 (O_2084,N_20177,N_23289);
xnor UO_2085 (O_2085,N_21358,N_19249);
and UO_2086 (O_2086,N_19209,N_20121);
xor UO_2087 (O_2087,N_20904,N_24712);
or UO_2088 (O_2088,N_19012,N_21391);
nor UO_2089 (O_2089,N_20669,N_21812);
and UO_2090 (O_2090,N_19729,N_23423);
xnor UO_2091 (O_2091,N_24171,N_20780);
nand UO_2092 (O_2092,N_22196,N_20308);
nand UO_2093 (O_2093,N_22362,N_23896);
or UO_2094 (O_2094,N_21876,N_19340);
xor UO_2095 (O_2095,N_23699,N_21417);
xnor UO_2096 (O_2096,N_21156,N_23923);
xor UO_2097 (O_2097,N_19194,N_20601);
xor UO_2098 (O_2098,N_24806,N_20341);
nand UO_2099 (O_2099,N_24481,N_18999);
nor UO_2100 (O_2100,N_22371,N_21121);
and UO_2101 (O_2101,N_22955,N_21110);
and UO_2102 (O_2102,N_22828,N_21486);
or UO_2103 (O_2103,N_18872,N_21956);
nor UO_2104 (O_2104,N_24904,N_24727);
or UO_2105 (O_2105,N_19105,N_19556);
and UO_2106 (O_2106,N_20144,N_22073);
xnor UO_2107 (O_2107,N_22500,N_22273);
nand UO_2108 (O_2108,N_20011,N_22961);
xnor UO_2109 (O_2109,N_24717,N_21773);
and UO_2110 (O_2110,N_18808,N_21414);
or UO_2111 (O_2111,N_18807,N_20411);
and UO_2112 (O_2112,N_20151,N_19233);
nand UO_2113 (O_2113,N_19819,N_22935);
and UO_2114 (O_2114,N_20155,N_19816);
nand UO_2115 (O_2115,N_24057,N_18913);
nand UO_2116 (O_2116,N_23306,N_20801);
xor UO_2117 (O_2117,N_24130,N_19215);
xnor UO_2118 (O_2118,N_22336,N_23274);
or UO_2119 (O_2119,N_22658,N_23396);
or UO_2120 (O_2120,N_24729,N_22448);
or UO_2121 (O_2121,N_19474,N_20424);
and UO_2122 (O_2122,N_21661,N_22315);
or UO_2123 (O_2123,N_20742,N_19135);
nand UO_2124 (O_2124,N_19575,N_23170);
xor UO_2125 (O_2125,N_23510,N_24895);
or UO_2126 (O_2126,N_20283,N_21772);
or UO_2127 (O_2127,N_18824,N_23172);
nand UO_2128 (O_2128,N_22862,N_23884);
nor UO_2129 (O_2129,N_21527,N_23544);
or UO_2130 (O_2130,N_20663,N_19109);
or UO_2131 (O_2131,N_22047,N_20111);
nor UO_2132 (O_2132,N_20775,N_21891);
xnor UO_2133 (O_2133,N_24223,N_18819);
or UO_2134 (O_2134,N_21687,N_22897);
nand UO_2135 (O_2135,N_19961,N_20190);
nand UO_2136 (O_2136,N_20586,N_20744);
nor UO_2137 (O_2137,N_22738,N_23322);
or UO_2138 (O_2138,N_22170,N_22375);
nor UO_2139 (O_2139,N_21051,N_20902);
and UO_2140 (O_2140,N_23138,N_23178);
nand UO_2141 (O_2141,N_24525,N_23548);
nand UO_2142 (O_2142,N_19916,N_23505);
nand UO_2143 (O_2143,N_20227,N_23171);
and UO_2144 (O_2144,N_20898,N_19519);
and UO_2145 (O_2145,N_23198,N_22716);
xor UO_2146 (O_2146,N_20357,N_18902);
or UO_2147 (O_2147,N_24302,N_19890);
xor UO_2148 (O_2148,N_24368,N_19843);
nor UO_2149 (O_2149,N_22361,N_19928);
nand UO_2150 (O_2150,N_20961,N_24000);
and UO_2151 (O_2151,N_23470,N_19123);
and UO_2152 (O_2152,N_23521,N_24070);
or UO_2153 (O_2153,N_23455,N_20738);
or UO_2154 (O_2154,N_19179,N_20765);
nand UO_2155 (O_2155,N_20421,N_20703);
nor UO_2156 (O_2156,N_23525,N_24683);
and UO_2157 (O_2157,N_22715,N_20383);
xnor UO_2158 (O_2158,N_20553,N_22012);
nor UO_2159 (O_2159,N_20696,N_21976);
and UO_2160 (O_2160,N_23650,N_24970);
xnor UO_2161 (O_2161,N_23091,N_21153);
xor UO_2162 (O_2162,N_20152,N_21704);
nand UO_2163 (O_2163,N_21312,N_19541);
nand UO_2164 (O_2164,N_22251,N_22425);
nand UO_2165 (O_2165,N_23002,N_19600);
xnor UO_2166 (O_2166,N_24915,N_22215);
xnor UO_2167 (O_2167,N_24536,N_24285);
nor UO_2168 (O_2168,N_21639,N_23803);
nor UO_2169 (O_2169,N_22295,N_23931);
nand UO_2170 (O_2170,N_23904,N_22293);
nand UO_2171 (O_2171,N_23445,N_23237);
xor UO_2172 (O_2172,N_23645,N_21880);
or UO_2173 (O_2173,N_23891,N_23349);
and UO_2174 (O_2174,N_22653,N_21826);
and UO_2175 (O_2175,N_22856,N_20330);
xnor UO_2176 (O_2176,N_19337,N_19802);
and UO_2177 (O_2177,N_20199,N_20312);
and UO_2178 (O_2178,N_23353,N_22434);
nand UO_2179 (O_2179,N_22900,N_21549);
nor UO_2180 (O_2180,N_23568,N_24653);
nor UO_2181 (O_2181,N_22880,N_22695);
nor UO_2182 (O_2182,N_20173,N_23082);
nor UO_2183 (O_2183,N_23180,N_21949);
or UO_2184 (O_2184,N_24633,N_23011);
xor UO_2185 (O_2185,N_21874,N_22510);
nor UO_2186 (O_2186,N_21071,N_24778);
xor UO_2187 (O_2187,N_23793,N_24617);
xnor UO_2188 (O_2188,N_22569,N_18920);
nand UO_2189 (O_2189,N_20720,N_24785);
or UO_2190 (O_2190,N_19571,N_19053);
and UO_2191 (O_2191,N_22710,N_20875);
xnor UO_2192 (O_2192,N_22760,N_23873);
or UO_2193 (O_2193,N_22003,N_20116);
nand UO_2194 (O_2194,N_24682,N_24590);
xnor UO_2195 (O_2195,N_19388,N_21569);
xnor UO_2196 (O_2196,N_22430,N_22914);
nand UO_2197 (O_2197,N_24042,N_24111);
nor UO_2198 (O_2198,N_19259,N_21983);
nor UO_2199 (O_2199,N_21736,N_23162);
and UO_2200 (O_2200,N_21969,N_19106);
or UO_2201 (O_2201,N_19026,N_21437);
nand UO_2202 (O_2202,N_23227,N_20753);
nand UO_2203 (O_2203,N_24355,N_23136);
or UO_2204 (O_2204,N_23158,N_21731);
or UO_2205 (O_2205,N_23690,N_21859);
or UO_2206 (O_2206,N_24885,N_18764);
and UO_2207 (O_2207,N_18933,N_21815);
nor UO_2208 (O_2208,N_24068,N_24979);
or UO_2209 (O_2209,N_18820,N_19595);
nor UO_2210 (O_2210,N_22798,N_21516);
nor UO_2211 (O_2211,N_21743,N_18780);
or UO_2212 (O_2212,N_22881,N_24950);
or UO_2213 (O_2213,N_20882,N_24971);
and UO_2214 (O_2214,N_23573,N_20419);
or UO_2215 (O_2215,N_20026,N_22973);
and UO_2216 (O_2216,N_20264,N_20206);
nand UO_2217 (O_2217,N_21747,N_19705);
nor UO_2218 (O_2218,N_20191,N_19069);
or UO_2219 (O_2219,N_23545,N_19486);
or UO_2220 (O_2220,N_23917,N_23401);
nor UO_2221 (O_2221,N_20254,N_21649);
nor UO_2222 (O_2222,N_19208,N_21326);
nor UO_2223 (O_2223,N_20899,N_21381);
nor UO_2224 (O_2224,N_24929,N_20216);
or UO_2225 (O_2225,N_24431,N_19222);
xnor UO_2226 (O_2226,N_20110,N_24508);
nand UO_2227 (O_2227,N_19581,N_20241);
nand UO_2228 (O_2228,N_24025,N_22861);
or UO_2229 (O_2229,N_21260,N_23400);
and UO_2230 (O_2230,N_21616,N_24338);
nand UO_2231 (O_2231,N_20545,N_22393);
or UO_2232 (O_2232,N_20825,N_20295);
nor UO_2233 (O_2233,N_20668,N_23036);
xnor UO_2234 (O_2234,N_21836,N_21699);
xor UO_2235 (O_2235,N_21948,N_23639);
and UO_2236 (O_2236,N_23549,N_22353);
xnor UO_2237 (O_2237,N_19795,N_18846);
nand UO_2238 (O_2238,N_20333,N_19089);
or UO_2239 (O_2239,N_20821,N_21170);
or UO_2240 (O_2240,N_19939,N_20338);
nand UO_2241 (O_2241,N_19081,N_22326);
and UO_2242 (O_2242,N_21230,N_23634);
nor UO_2243 (O_2243,N_18919,N_21369);
and UO_2244 (O_2244,N_21236,N_24358);
and UO_2245 (O_2245,N_19368,N_18840);
xnor UO_2246 (O_2246,N_20457,N_24500);
xor UO_2247 (O_2247,N_21707,N_24468);
nand UO_2248 (O_2248,N_22783,N_21806);
or UO_2249 (O_2249,N_19688,N_21793);
nor UO_2250 (O_2250,N_21977,N_21513);
xor UO_2251 (O_2251,N_21975,N_24215);
nor UO_2252 (O_2252,N_24553,N_21499);
nor UO_2253 (O_2253,N_19512,N_19125);
or UO_2254 (O_2254,N_24902,N_21021);
or UO_2255 (O_2255,N_24956,N_23902);
nand UO_2256 (O_2256,N_21497,N_22751);
or UO_2257 (O_2257,N_21306,N_20202);
nor UO_2258 (O_2258,N_22572,N_19316);
and UO_2259 (O_2259,N_23157,N_19309);
or UO_2260 (O_2260,N_23646,N_24749);
nor UO_2261 (O_2261,N_20205,N_19793);
or UO_2262 (O_2262,N_21528,N_20792);
nand UO_2263 (O_2263,N_22064,N_20894);
nand UO_2264 (O_2264,N_19014,N_24469);
nand UO_2265 (O_2265,N_21592,N_19144);
nor UO_2266 (O_2266,N_23148,N_24735);
nor UO_2267 (O_2267,N_22978,N_23848);
nand UO_2268 (O_2268,N_24125,N_21877);
xor UO_2269 (O_2269,N_20076,N_19464);
xor UO_2270 (O_2270,N_20452,N_19329);
and UO_2271 (O_2271,N_24044,N_18883);
nor UO_2272 (O_2272,N_22396,N_22280);
xnor UO_2273 (O_2273,N_21820,N_24023);
or UO_2274 (O_2274,N_22376,N_21267);
and UO_2275 (O_2275,N_22977,N_22449);
xor UO_2276 (O_2276,N_24615,N_21321);
nand UO_2277 (O_2277,N_20923,N_23379);
xnor UO_2278 (O_2278,N_20459,N_19609);
nand UO_2279 (O_2279,N_24354,N_21375);
xor UO_2280 (O_2280,N_23386,N_22455);
nor UO_2281 (O_2281,N_20728,N_23822);
nor UO_2282 (O_2282,N_19554,N_19362);
xnor UO_2283 (O_2283,N_19212,N_19213);
xnor UO_2284 (O_2284,N_21400,N_23010);
nand UO_2285 (O_2285,N_23499,N_19949);
and UO_2286 (O_2286,N_22489,N_20376);
nor UO_2287 (O_2287,N_20524,N_20127);
nand UO_2288 (O_2288,N_23863,N_22078);
or UO_2289 (O_2289,N_20247,N_19117);
xnor UO_2290 (O_2290,N_23881,N_19756);
xor UO_2291 (O_2291,N_21803,N_21205);
or UO_2292 (O_2292,N_21713,N_21274);
or UO_2293 (O_2293,N_21320,N_24721);
xor UO_2294 (O_2294,N_20179,N_20543);
nand UO_2295 (O_2295,N_23094,N_21894);
nor UO_2296 (O_2296,N_22571,N_23081);
nor UO_2297 (O_2297,N_20402,N_19734);
nand UO_2298 (O_2298,N_23961,N_19041);
and UO_2299 (O_2299,N_20493,N_20692);
and UO_2300 (O_2300,N_20674,N_21496);
xor UO_2301 (O_2301,N_20823,N_24495);
and UO_2302 (O_2302,N_21422,N_23558);
or UO_2303 (O_2303,N_22641,N_22248);
xor UO_2304 (O_2304,N_20324,N_22470);
xor UO_2305 (O_2305,N_22374,N_20467);
xnor UO_2306 (O_2306,N_21561,N_20085);
nor UO_2307 (O_2307,N_20951,N_21659);
xnor UO_2308 (O_2308,N_19252,N_22268);
and UO_2309 (O_2309,N_22865,N_21160);
nand UO_2310 (O_2310,N_19149,N_22257);
nor UO_2311 (O_2311,N_21224,N_22533);
xor UO_2312 (O_2312,N_21435,N_20960);
nor UO_2313 (O_2313,N_22594,N_24648);
nand UO_2314 (O_2314,N_24264,N_24265);
nor UO_2315 (O_2315,N_19088,N_18917);
nor UO_2316 (O_2316,N_23921,N_20502);
or UO_2317 (O_2317,N_23637,N_19268);
nor UO_2318 (O_2318,N_21563,N_24947);
nand UO_2319 (O_2319,N_20072,N_21742);
nand UO_2320 (O_2320,N_24673,N_24830);
nor UO_2321 (O_2321,N_19487,N_24869);
and UO_2322 (O_2322,N_19385,N_19800);
nand UO_2323 (O_2323,N_19145,N_20364);
and UO_2324 (O_2324,N_20287,N_19078);
nand UO_2325 (O_2325,N_22755,N_22542);
xnor UO_2326 (O_2326,N_23057,N_21000);
or UO_2327 (O_2327,N_21995,N_23484);
or UO_2328 (O_2328,N_21070,N_20161);
xor UO_2329 (O_2329,N_23115,N_21690);
or UO_2330 (O_2330,N_21939,N_22496);
and UO_2331 (O_2331,N_20239,N_20020);
and UO_2332 (O_2332,N_19472,N_19709);
xor UO_2333 (O_2333,N_21680,N_22474);
and UO_2334 (O_2334,N_18777,N_23724);
xnor UO_2335 (O_2335,N_23027,N_19370);
xnor UO_2336 (O_2336,N_20221,N_21002);
nor UO_2337 (O_2337,N_21777,N_20808);
nor UO_2338 (O_2338,N_20142,N_24004);
or UO_2339 (O_2339,N_19515,N_20154);
and UO_2340 (O_2340,N_21898,N_19834);
xnor UO_2341 (O_2341,N_22540,N_22011);
nand UO_2342 (O_2342,N_21432,N_20412);
xnor UO_2343 (O_2343,N_19013,N_21544);
or UO_2344 (O_2344,N_20087,N_21433);
xnor UO_2345 (O_2345,N_22459,N_19857);
nand UO_2346 (O_2346,N_19772,N_19155);
nor UO_2347 (O_2347,N_23739,N_22104);
nand UO_2348 (O_2348,N_23222,N_21719);
xor UO_2349 (O_2349,N_23109,N_18922);
or UO_2350 (O_2350,N_20470,N_23671);
xor UO_2351 (O_2351,N_23669,N_19372);
nor UO_2352 (O_2352,N_23567,N_22381);
or UO_2353 (O_2353,N_22416,N_23312);
xor UO_2354 (O_2354,N_19357,N_21090);
xnor UO_2355 (O_2355,N_22118,N_21737);
or UO_2356 (O_2356,N_24608,N_24955);
nor UO_2357 (O_2357,N_24116,N_20924);
and UO_2358 (O_2358,N_22717,N_24152);
nor UO_2359 (O_2359,N_21053,N_24589);
nand UO_2360 (O_2360,N_22803,N_19578);
xor UO_2361 (O_2361,N_23800,N_23123);
or UO_2362 (O_2362,N_18914,N_20032);
or UO_2363 (O_2363,N_20725,N_19322);
nand UO_2364 (O_2364,N_20010,N_19130);
and UO_2365 (O_2365,N_21718,N_19630);
and UO_2366 (O_2366,N_22669,N_19462);
nor UO_2367 (O_2367,N_23218,N_24739);
or UO_2368 (O_2368,N_22354,N_22287);
nand UO_2369 (O_2369,N_21567,N_24760);
xnor UO_2370 (O_2370,N_23794,N_19483);
and UO_2371 (O_2371,N_20393,N_24033);
or UO_2372 (O_2372,N_24202,N_19258);
and UO_2373 (O_2373,N_19809,N_23481);
and UO_2374 (O_2374,N_20797,N_21446);
nor UO_2375 (O_2375,N_18759,N_24420);
and UO_2376 (O_2376,N_20677,N_20490);
xnor UO_2377 (O_2377,N_23316,N_21688);
and UO_2378 (O_2378,N_19048,N_23824);
nand UO_2379 (O_2379,N_23869,N_22199);
and UO_2380 (O_2380,N_22457,N_24013);
nor UO_2381 (O_2381,N_23964,N_19456);
or UO_2382 (O_2382,N_24754,N_22832);
xor UO_2383 (O_2383,N_19833,N_20912);
xnor UO_2384 (O_2384,N_20724,N_19235);
xnor UO_2385 (O_2385,N_24329,N_19669);
or UO_2386 (O_2386,N_21600,N_19098);
xnor UO_2387 (O_2387,N_21750,N_22741);
xnor UO_2388 (O_2388,N_21548,N_24376);
nor UO_2389 (O_2389,N_22948,N_22177);
xnor UO_2390 (O_2390,N_21038,N_19891);
and UO_2391 (O_2391,N_20158,N_19871);
nand UO_2392 (O_2392,N_24090,N_21913);
nor UO_2393 (O_2393,N_21195,N_23398);
nor UO_2394 (O_2394,N_23458,N_24961);
xor UO_2395 (O_2395,N_20262,N_22258);
and UO_2396 (O_2396,N_22551,N_19652);
xor UO_2397 (O_2397,N_22033,N_23087);
xor UO_2398 (O_2398,N_21455,N_23506);
nand UO_2399 (O_2399,N_23008,N_18790);
or UO_2400 (O_2400,N_21174,N_22519);
or UO_2401 (O_2401,N_21408,N_20143);
nand UO_2402 (O_2402,N_24309,N_22101);
and UO_2403 (O_2403,N_23653,N_24865);
xnor UO_2404 (O_2404,N_23300,N_21292);
and UO_2405 (O_2405,N_23552,N_19957);
xor UO_2406 (O_2406,N_23406,N_24649);
nand UO_2407 (O_2407,N_23529,N_20400);
nand UO_2408 (O_2408,N_21008,N_22918);
and UO_2409 (O_2409,N_20590,N_20404);
and UO_2410 (O_2410,N_24925,N_20687);
nand UO_2411 (O_2411,N_20193,N_21696);
or UO_2412 (O_2412,N_24794,N_24977);
nand UO_2413 (O_2413,N_21722,N_20946);
or UO_2414 (O_2414,N_19444,N_20609);
nor UO_2415 (O_2415,N_19216,N_18996);
and UO_2416 (O_2416,N_20885,N_24650);
or UO_2417 (O_2417,N_19139,N_19905);
nor UO_2418 (O_2418,N_21241,N_23564);
nand UO_2419 (O_2419,N_19299,N_20237);
and UO_2420 (O_2420,N_21530,N_19590);
xor UO_2421 (O_2421,N_21262,N_19599);
and UO_2422 (O_2422,N_19112,N_19307);
nand UO_2423 (O_2423,N_24110,N_23378);
or UO_2424 (O_2424,N_20494,N_20565);
or UO_2425 (O_2425,N_20542,N_24060);
xnor UO_2426 (O_2426,N_18953,N_24575);
nor UO_2427 (O_2427,N_24129,N_24128);
or UO_2428 (O_2428,N_23307,N_20477);
and UO_2429 (O_2429,N_24109,N_19292);
or UO_2430 (O_2430,N_24827,N_20709);
or UO_2431 (O_2431,N_21915,N_23647);
xnor UO_2432 (O_2432,N_24222,N_19118);
or UO_2433 (O_2433,N_19805,N_22256);
and UO_2434 (O_2434,N_24456,N_19906);
or UO_2435 (O_2435,N_19324,N_20615);
or UO_2436 (O_2436,N_19872,N_22424);
and UO_2437 (O_2437,N_24209,N_23475);
nor UO_2438 (O_2438,N_20964,N_21883);
nor UO_2439 (O_2439,N_24024,N_22318);
and UO_2440 (O_2440,N_19022,N_24911);
nand UO_2441 (O_2441,N_23749,N_20522);
xnor UO_2442 (O_2442,N_22208,N_19538);
and UO_2443 (O_2443,N_22402,N_18829);
nor UO_2444 (O_2444,N_24720,N_23422);
and UO_2445 (O_2445,N_19981,N_23926);
xnor UO_2446 (O_2446,N_24926,N_22621);
nor UO_2447 (O_2447,N_21640,N_21479);
xor UO_2448 (O_2448,N_23537,N_24671);
nand UO_2449 (O_2449,N_23197,N_24996);
xnor UO_2450 (O_2450,N_21755,N_23866);
and UO_2451 (O_2451,N_19623,N_18931);
xnor UO_2452 (O_2452,N_19695,N_21030);
xor UO_2453 (O_2453,N_24808,N_23523);
nand UO_2454 (O_2454,N_21189,N_24499);
nand UO_2455 (O_2455,N_24498,N_21518);
or UO_2456 (O_2456,N_19438,N_23369);
and UO_2457 (O_2457,N_20594,N_23021);
or UO_2458 (O_2458,N_24694,N_22435);
nand UO_2459 (O_2459,N_24662,N_24874);
nor UO_2460 (O_2460,N_18860,N_24178);
nand UO_2461 (O_2461,N_22486,N_22909);
xor UO_2462 (O_2462,N_23936,N_21502);
nand UO_2463 (O_2463,N_23040,N_22618);
xor UO_2464 (O_2464,N_20934,N_24115);
xor UO_2465 (O_2465,N_23995,N_22953);
xor UO_2466 (O_2466,N_24186,N_22592);
xnor UO_2467 (O_2467,N_19899,N_22562);
nand UO_2468 (O_2468,N_23121,N_18977);
or UO_2469 (O_2469,N_20993,N_19953);
or UO_2470 (O_2470,N_24094,N_19887);
or UO_2471 (O_2471,N_23858,N_24166);
nand UO_2472 (O_2472,N_21397,N_19754);
or UO_2473 (O_2473,N_21234,N_23531);
xor UO_2474 (O_2474,N_19488,N_21271);
and UO_2475 (O_2475,N_23217,N_24438);
and UO_2476 (O_2476,N_18844,N_19410);
and UO_2477 (O_2477,N_24031,N_21295);
or UO_2478 (O_2478,N_24679,N_23188);
nor UO_2479 (O_2479,N_24554,N_23928);
xor UO_2480 (O_2480,N_23909,N_23990);
xor UO_2481 (O_2481,N_21211,N_20838);
and UO_2482 (O_2482,N_19010,N_21120);
and UO_2483 (O_2483,N_23442,N_21297);
nor UO_2484 (O_2484,N_23285,N_19864);
or UO_2485 (O_2485,N_20275,N_22998);
and UO_2486 (O_2486,N_24078,N_20069);
or UO_2487 (O_2487,N_23034,N_20532);
nor UO_2488 (O_2488,N_23088,N_23411);
nand UO_2489 (O_2489,N_20769,N_21998);
xor UO_2490 (O_2490,N_18964,N_19220);
xor UO_2491 (O_2491,N_23636,N_23605);
nor UO_2492 (O_2492,N_22954,N_21922);
and UO_2493 (O_2493,N_24809,N_20884);
xor UO_2494 (O_2494,N_23612,N_19005);
nand UO_2495 (O_2495,N_22666,N_21447);
xnor UO_2496 (O_2496,N_23541,N_24149);
nand UO_2497 (O_2497,N_24674,N_23870);
xor UO_2498 (O_2498,N_24742,N_20014);
or UO_2499 (O_2499,N_19823,N_21550);
nor UO_2500 (O_2500,N_21981,N_24009);
and UO_2501 (O_2501,N_22837,N_20606);
xnor UO_2502 (O_2502,N_21663,N_18998);
xor UO_2503 (O_2503,N_23383,N_19422);
xnor UO_2504 (O_2504,N_21149,N_22232);
xor UO_2505 (O_2505,N_20462,N_22895);
or UO_2506 (O_2506,N_19200,N_18841);
nor UO_2507 (O_2507,N_22858,N_24415);
and UO_2508 (O_2508,N_20018,N_18852);
nor UO_2509 (O_2509,N_23425,N_22453);
xnor UO_2510 (O_2510,N_24226,N_20840);
and UO_2511 (O_2511,N_21648,N_22305);
or UO_2512 (O_2512,N_20068,N_20888);
xor UO_2513 (O_2513,N_23585,N_19350);
xnor UO_2514 (O_2514,N_20573,N_21302);
xnor UO_2515 (O_2515,N_20881,N_23756);
xor UO_2516 (O_2516,N_21602,N_24684);
nor UO_2517 (O_2517,N_19561,N_22560);
or UO_2518 (O_2518,N_24628,N_23280);
xor UO_2519 (O_2519,N_22178,N_21924);
nand UO_2520 (O_2520,N_24298,N_19256);
nor UO_2521 (O_2521,N_22604,N_21525);
and UO_2522 (O_2522,N_20025,N_22664);
and UO_2523 (O_2523,N_22181,N_20392);
or UO_2524 (O_2524,N_23532,N_19637);
xnor UO_2525 (O_2525,N_22645,N_18767);
nand UO_2526 (O_2526,N_23949,N_21117);
xor UO_2527 (O_2527,N_19151,N_19431);
nand UO_2528 (O_2528,N_23985,N_20385);
nand UO_2529 (O_2529,N_22761,N_18900);
or UO_2530 (O_2530,N_19778,N_22304);
and UO_2531 (O_2531,N_22378,N_23436);
and UO_2532 (O_2532,N_24738,N_24409);
or UO_2533 (O_2533,N_23999,N_23007);
xnor UO_2534 (O_2534,N_20723,N_21784);
nand UO_2535 (O_2535,N_24348,N_23522);
or UO_2536 (O_2536,N_22391,N_20581);
xnor UO_2537 (O_2537,N_23018,N_21761);
nand UO_2538 (O_2538,N_23268,N_23712);
nand UO_2539 (O_2539,N_23142,N_22143);
and UO_2540 (O_2540,N_19545,N_24266);
nand UO_2541 (O_2541,N_19713,N_23676);
or UO_2542 (O_2542,N_23459,N_24777);
xnor UO_2543 (O_2543,N_24080,N_24763);
nand UO_2544 (O_2544,N_24887,N_24212);
nand UO_2545 (O_2545,N_24247,N_24965);
and UO_2546 (O_2546,N_22924,N_20755);
xnor UO_2547 (O_2547,N_24487,N_23357);
or UO_2548 (O_2548,N_20698,N_24093);
xnor UO_2549 (O_2549,N_22764,N_20063);
or UO_2550 (O_2550,N_20482,N_21130);
xor UO_2551 (O_2551,N_21631,N_23804);
xor UO_2552 (O_2552,N_18838,N_19419);
xnor UO_2553 (O_2553,N_20967,N_19794);
and UO_2554 (O_2554,N_19856,N_23682);
and UO_2555 (O_2555,N_18857,N_20789);
xnor UO_2556 (O_2556,N_24173,N_21344);
xnor UO_2557 (O_2557,N_21248,N_20478);
or UO_2558 (O_2558,N_23983,N_24026);
nand UO_2559 (O_2559,N_22993,N_21399);
nor UO_2560 (O_2560,N_19938,N_22515);
and UO_2561 (O_2561,N_18750,N_24917);
or UO_2562 (O_2562,N_23589,N_19518);
and UO_2563 (O_2563,N_23959,N_22201);
or UO_2564 (O_2564,N_22581,N_23392);
xnor UO_2565 (O_2565,N_24389,N_23740);
nand UO_2566 (O_2566,N_19380,N_21460);
nor UO_2567 (O_2567,N_20802,N_20982);
or UO_2568 (O_2568,N_23342,N_19097);
xnor UO_2569 (O_2569,N_20824,N_24570);
xor UO_2570 (O_2570,N_21427,N_21091);
nand UO_2571 (O_2571,N_19694,N_19534);
nor UO_2572 (O_2572,N_22962,N_23799);
nand UO_2573 (O_2573,N_21069,N_23151);
nor UO_2574 (O_2574,N_19159,N_20635);
nor UO_2575 (O_2575,N_23052,N_21309);
and UO_2576 (O_2576,N_20099,N_21547);
xor UO_2577 (O_2577,N_19262,N_22815);
nor UO_2578 (O_2578,N_20535,N_22587);
xor UO_2579 (O_2579,N_19057,N_22713);
nor UO_2580 (O_2580,N_21099,N_19381);
or UO_2581 (O_2581,N_19185,N_20329);
or UO_2582 (O_2582,N_20624,N_20628);
and UO_2583 (O_2583,N_23763,N_22493);
or UO_2584 (O_2584,N_19202,N_24945);
nand UO_2585 (O_2585,N_23801,N_22619);
or UO_2586 (O_2586,N_21698,N_19485);
and UO_2587 (O_2587,N_24701,N_19943);
nor UO_2588 (O_2588,N_22135,N_20814);
xnor UO_2589 (O_2589,N_24836,N_21077);
and UO_2590 (O_2590,N_20187,N_20897);
or UO_2591 (O_2591,N_21468,N_21541);
nor UO_2592 (O_2592,N_20560,N_24661);
and UO_2593 (O_2593,N_19432,N_20045);
nand UO_2594 (O_2594,N_22567,N_23594);
nand UO_2595 (O_2595,N_20736,N_21867);
nand UO_2596 (O_2596,N_19668,N_21495);
and UO_2597 (O_2597,N_21684,N_21416);
nand UO_2598 (O_2598,N_19465,N_21231);
nand UO_2599 (O_2599,N_23978,N_18837);
and UO_2600 (O_2600,N_24843,N_20900);
or UO_2601 (O_2601,N_21106,N_18802);
xnor UO_2602 (O_2602,N_21118,N_24851);
xor UO_2603 (O_2603,N_19269,N_24072);
or UO_2604 (O_2604,N_20616,N_20214);
or UO_2605 (O_2605,N_24657,N_21907);
nor UO_2606 (O_2606,N_18897,N_24621);
nor UO_2607 (O_2607,N_24985,N_22216);
and UO_2608 (O_2608,N_23945,N_19498);
nor UO_2609 (O_2609,N_24831,N_22994);
nor UO_2610 (O_2610,N_23061,N_23140);
xor UO_2611 (O_2611,N_22040,N_20013);
xnor UO_2612 (O_2612,N_24224,N_23462);
xnor UO_2613 (O_2613,N_20800,N_24308);
and UO_2614 (O_2614,N_23169,N_22384);
nor UO_2615 (O_2615,N_24036,N_22600);
nor UO_2616 (O_2616,N_19287,N_21869);
and UO_2617 (O_2617,N_19661,N_23582);
nor UO_2618 (O_2618,N_24423,N_23210);
nand UO_2619 (O_2619,N_23547,N_20422);
or UO_2620 (O_2620,N_22197,N_18936);
or UO_2621 (O_2621,N_21390,N_21715);
and UO_2622 (O_2622,N_22595,N_22102);
nor UO_2623 (O_2623,N_21216,N_24852);
or UO_2624 (O_2624,N_22076,N_24698);
nor UO_2625 (O_2625,N_23868,N_21589);
xor UO_2626 (O_2626,N_21852,N_21073);
nor UO_2627 (O_2627,N_20102,N_20950);
and UO_2628 (O_2628,N_21166,N_20571);
or UO_2629 (O_2629,N_20195,N_24147);
or UO_2630 (O_2630,N_23680,N_23687);
xor UO_2631 (O_2631,N_23029,N_23233);
nor UO_2632 (O_2632,N_20689,N_19925);
nor UO_2633 (O_2633,N_23707,N_19964);
xnor UO_2634 (O_2634,N_22050,N_19715);
xnor UO_2635 (O_2635,N_19223,N_24316);
nor UO_2636 (O_2636,N_23135,N_19407);
nor UO_2637 (O_2637,N_23271,N_20558);
nor UO_2638 (O_2638,N_21571,N_22884);
nor UO_2639 (O_2639,N_24428,N_23982);
nor UO_2640 (O_2640,N_24816,N_19166);
and UO_2641 (O_2641,N_20440,N_21818);
and UO_2642 (O_2642,N_24211,N_19420);
and UO_2643 (O_2643,N_24242,N_19898);
nand UO_2644 (O_2644,N_20465,N_23828);
nor UO_2645 (O_2645,N_19740,N_22131);
nor UO_2646 (O_2646,N_23488,N_18975);
nand UO_2647 (O_2647,N_23842,N_22409);
nand UO_2648 (O_2648,N_19814,N_22574);
nor UO_2649 (O_2649,N_20890,N_24335);
nand UO_2650 (O_2650,N_21193,N_18835);
and UO_2651 (O_2651,N_23377,N_21817);
xnor UO_2652 (O_2652,N_20914,N_23028);
nand UO_2653 (O_2653,N_21695,N_24850);
or UO_2654 (O_2654,N_22054,N_18761);
xnor UO_2655 (O_2655,N_22377,N_23068);
and UO_2656 (O_2656,N_19827,N_21848);
or UO_2657 (O_2657,N_23467,N_24073);
nand UO_2658 (O_2658,N_22746,N_23107);
xor UO_2659 (O_2659,N_20464,N_23665);
xnor UO_2660 (O_2660,N_22607,N_21745);
or UO_2661 (O_2661,N_21337,N_21816);
or UO_2662 (O_2662,N_19622,N_21129);
nor UO_2663 (O_2663,N_20073,N_20563);
or UO_2664 (O_2664,N_22793,N_23156);
nor UO_2665 (O_2665,N_23014,N_22693);
nand UO_2666 (O_2666,N_19409,N_20992);
nor UO_2667 (O_2667,N_23570,N_24700);
nand UO_2668 (O_2668,N_19255,N_24245);
or UO_2669 (O_2669,N_24801,N_23302);
nor UO_2670 (O_2670,N_23814,N_19015);
xor UO_2671 (O_2671,N_22278,N_23200);
and UO_2672 (O_2672,N_23220,N_24612);
and UO_2673 (O_2673,N_19017,N_22193);
xor UO_2674 (O_2674,N_21760,N_19344);
and UO_2675 (O_2675,N_21190,N_20986);
nor UO_2676 (O_2676,N_21519,N_22850);
or UO_2677 (O_2677,N_20715,N_24296);
nand UO_2678 (O_2678,N_23390,N_18752);
nand UO_2679 (O_2679,N_20953,N_23910);
xor UO_2680 (O_2680,N_19758,N_23746);
and UO_2681 (O_2681,N_18827,N_20378);
and UO_2682 (O_2682,N_21201,N_24333);
or UO_2683 (O_2683,N_19841,N_20244);
nand UO_2684 (O_2684,N_22748,N_19673);
nor UO_2685 (O_2685,N_23989,N_19849);
nor UO_2686 (O_2686,N_23908,N_21746);
or UO_2687 (O_2687,N_22981,N_18985);
nor UO_2688 (O_2688,N_22615,N_21709);
and UO_2689 (O_2689,N_23790,N_22768);
and UO_2690 (O_2690,N_24069,N_19207);
or UO_2691 (O_2691,N_21916,N_20012);
nand UO_2692 (O_2692,N_24055,N_18908);
nand UO_2693 (O_2693,N_24286,N_19593);
nand UO_2694 (O_2694,N_18987,N_21288);
xor UO_2695 (O_2695,N_24138,N_20655);
or UO_2696 (O_2696,N_23886,N_21645);
nand UO_2697 (O_2697,N_20134,N_23883);
nor UO_2698 (O_2698,N_24043,N_19874);
nor UO_2699 (O_2699,N_20585,N_24021);
nand UO_2700 (O_2700,N_24427,N_23495);
or UO_2701 (O_2701,N_19495,N_24433);
or UO_2702 (O_2702,N_21027,N_20714);
nor UO_2703 (O_2703,N_24188,N_19908);
or UO_2704 (O_2704,N_21878,N_20886);
or UO_2705 (O_2705,N_22943,N_23287);
or UO_2706 (O_2706,N_19280,N_20685);
and UO_2707 (O_2707,N_21244,N_21553);
xor UO_2708 (O_2708,N_23295,N_21011);
and UO_2709 (O_2709,N_24790,N_19716);
or UO_2710 (O_2710,N_24257,N_21686);
nor UO_2711 (O_2711,N_22291,N_23310);
and UO_2712 (O_2712,N_21064,N_22279);
and UO_2713 (O_2713,N_19042,N_19563);
or UO_2714 (O_2714,N_23020,N_20584);
xnor UO_2715 (O_2715,N_24449,N_19913);
and UO_2716 (O_2716,N_18791,N_24155);
nand UO_2717 (O_2717,N_23298,N_19616);
nand UO_2718 (O_2718,N_24473,N_23751);
nor UO_2719 (O_2719,N_19804,N_20555);
or UO_2720 (O_2720,N_23095,N_24999);
nor UO_2721 (O_2721,N_24104,N_19398);
nor UO_2722 (O_2722,N_22894,N_23890);
or UO_2723 (O_2723,N_24010,N_19601);
or UO_2724 (O_2724,N_22026,N_23317);
nor UO_2725 (O_2725,N_19667,N_21932);
or UO_2726 (O_2726,N_24502,N_20232);
xor UO_2727 (O_2727,N_22539,N_22460);
or UO_2728 (O_2728,N_24974,N_23080);
nand UO_2729 (O_2729,N_18861,N_18957);
and UO_2730 (O_2730,N_22853,N_21464);
and UO_2731 (O_2731,N_23017,N_19314);
nor UO_2732 (O_2732,N_24434,N_24319);
and UO_2733 (O_2733,N_22795,N_24474);
and UO_2734 (O_2734,N_21990,N_20433);
and UO_2735 (O_2735,N_24780,N_20519);
nand UO_2736 (O_2736,N_23480,N_22190);
nand UO_2737 (O_2737,N_23586,N_19221);
xor UO_2738 (O_2738,N_19242,N_22082);
nor UO_2739 (O_2739,N_24614,N_19583);
xnor UO_2740 (O_2740,N_21037,N_20060);
xnor UO_2741 (O_2741,N_21393,N_23629);
nor UO_2742 (O_2742,N_24506,N_22020);
or UO_2743 (O_2743,N_20664,N_21389);
or UO_2744 (O_2744,N_20569,N_19762);
and UO_2745 (O_2745,N_23290,N_21067);
or UO_2746 (O_2746,N_21098,N_22544);
nor UO_2747 (O_2747,N_24278,N_21015);
or UO_2748 (O_2748,N_23141,N_24478);
and UO_2749 (O_2749,N_23742,N_23254);
xor UO_2750 (O_2750,N_24196,N_23503);
or UO_2751 (O_2751,N_19061,N_23836);
xnor UO_2752 (O_2752,N_22467,N_23434);
xnor UO_2753 (O_2753,N_24181,N_19499);
nor UO_2754 (O_2754,N_23249,N_18773);
nand UO_2755 (O_2755,N_21384,N_22629);
xor UO_2756 (O_2756,N_21840,N_24829);
nand UO_2757 (O_2757,N_19318,N_21085);
nor UO_2758 (O_2758,N_21702,N_20867);
or UO_2759 (O_2759,N_19743,N_23013);
and UO_2760 (O_2760,N_23278,N_23212);
or UO_2761 (O_2761,N_23618,N_22408);
nand UO_2762 (O_2762,N_22024,N_22644);
or UO_2763 (O_2763,N_21191,N_24889);
nor UO_2764 (O_2764,N_23194,N_20794);
nand UO_2765 (O_2765,N_22202,N_19165);
or UO_2766 (O_2766,N_21605,N_21582);
or UO_2767 (O_2767,N_24231,N_24773);
xnor UO_2768 (O_2768,N_22566,N_22117);
xnor UO_2769 (O_2769,N_22771,N_18850);
xnor UO_2770 (O_2770,N_24878,N_18961);
xor UO_2771 (O_2771,N_19780,N_19531);
or UO_2772 (O_2772,N_21310,N_19336);
or UO_2773 (O_2773,N_18966,N_20752);
nand UO_2774 (O_2774,N_19353,N_24941);
nand UO_2775 (O_2775,N_22129,N_21643);
and UO_2776 (O_2776,N_22724,N_21864);
or UO_2777 (O_2777,N_22758,N_23565);
and UO_2778 (O_2778,N_22243,N_24672);
nand UO_2779 (O_2779,N_24280,N_23953);
or UO_2780 (O_2780,N_21451,N_22022);
and UO_2781 (O_2781,N_19520,N_24288);
nor UO_2782 (O_2782,N_23352,N_21144);
or UO_2783 (O_2783,N_20839,N_22265);
and UO_2784 (O_2784,N_22080,N_19923);
nand UO_2785 (O_2785,N_18770,N_20943);
nor UO_2786 (O_2786,N_23100,N_24239);
or UO_2787 (O_2787,N_18854,N_20415);
or UO_2788 (O_2788,N_20384,N_23747);
or UO_2789 (O_2789,N_18862,N_21299);
nand UO_2790 (O_2790,N_18890,N_22183);
nor UO_2791 (O_2791,N_22917,N_20335);
and UO_2792 (O_2792,N_19642,N_23264);
and UO_2793 (O_2793,N_24003,N_19811);
nor UO_2794 (O_2794,N_19634,N_24367);
and UO_2795 (O_2795,N_20148,N_20642);
xnor UO_2796 (O_2796,N_22394,N_24867);
nor UO_2797 (O_2797,N_21656,N_23816);
nor UO_2798 (O_2798,N_20327,N_20708);
nor UO_2799 (O_2799,N_18814,N_24594);
xnor UO_2800 (O_2800,N_24919,N_24318);
and UO_2801 (O_2801,N_23320,N_19460);
nor UO_2802 (O_2802,N_19641,N_21367);
or UO_2803 (O_2803,N_24509,N_21424);
xor UO_2804 (O_2804,N_22308,N_19189);
and UO_2805 (O_2805,N_20083,N_22529);
and UO_2806 (O_2806,N_24516,N_23356);
or UO_2807 (O_2807,N_22031,N_19763);
nand UO_2808 (O_2808,N_21712,N_21933);
nand UO_2809 (O_2809,N_20196,N_21371);
xor UO_2810 (O_2810,N_19784,N_23893);
nor UO_2811 (O_2811,N_20853,N_22949);
nor UO_2812 (O_2812,N_18803,N_23325);
xor UO_2813 (O_2813,N_24722,N_21608);
nor UO_2814 (O_2814,N_22609,N_20526);
xnor UO_2815 (O_2815,N_19810,N_20631);
nand UO_2816 (O_2816,N_23927,N_22692);
nand UO_2817 (O_2817,N_24942,N_19621);
nor UO_2818 (O_2818,N_20818,N_20145);
and UO_2819 (O_2819,N_20734,N_23643);
xnor UO_2820 (O_2820,N_24613,N_23113);
nor UO_2821 (O_2821,N_19876,N_19278);
and UO_2822 (O_2822,N_19351,N_19917);
xnor UO_2823 (O_2823,N_21491,N_20222);
nor UO_2824 (O_2824,N_23760,N_23191);
and UO_2825 (O_2825,N_23146,N_23154);
and UO_2826 (O_2826,N_22543,N_21873);
nor UO_2827 (O_2827,N_20192,N_23159);
and UO_2828 (O_2828,N_23231,N_22121);
nor UO_2829 (O_2829,N_22045,N_19295);
nor UO_2830 (O_2830,N_20521,N_22168);
or UO_2831 (O_2831,N_23405,N_19560);
and UO_2832 (O_2832,N_20948,N_22097);
or UO_2833 (O_2833,N_21610,N_23048);
xor UO_2834 (O_2834,N_18940,N_21388);
xor UO_2835 (O_2835,N_18865,N_19303);
and UO_2836 (O_2836,N_23124,N_22451);
xor UO_2837 (O_2837,N_22192,N_24405);
xnor UO_2838 (O_2838,N_22471,N_24595);
nor UO_2839 (O_2839,N_21006,N_20089);
or UO_2840 (O_2840,N_20562,N_24540);
and UO_2841 (O_2841,N_24360,N_18795);
nand UO_2842 (O_2842,N_20273,N_22446);
or UO_2843 (O_2843,N_22356,N_24136);
and UO_2844 (O_2844,N_18776,N_19417);
xor UO_2845 (O_2845,N_19143,N_24352);
or UO_2846 (O_2846,N_24826,N_22585);
nor UO_2847 (O_2847,N_19748,N_23189);
nand UO_2848 (O_2848,N_22719,N_20186);
xnor UO_2849 (O_2849,N_19686,N_19082);
xnor UO_2850 (O_2850,N_21361,N_20123);
and UO_2851 (O_2851,N_19272,N_20260);
xor UO_2852 (O_2852,N_21043,N_20135);
nor UO_2853 (O_2853,N_22108,N_21875);
and UO_2854 (O_2854,N_24407,N_20181);
xnor UO_2855 (O_2855,N_24208,N_20920);
xor UO_2856 (O_2856,N_20855,N_24275);
and UO_2857 (O_2857,N_20300,N_22780);
and UO_2858 (O_2858,N_23003,N_19658);
nor UO_2859 (O_2859,N_19377,N_23554);
nand UO_2860 (O_2860,N_23577,N_21264);
xor UO_2861 (O_2861,N_22290,N_21080);
and UO_2862 (O_2862,N_18898,N_20203);
nor UO_2863 (O_2863,N_23767,N_20019);
and UO_2864 (O_2864,N_22001,N_22488);
or UO_2865 (O_2865,N_18815,N_20501);
nor UO_2866 (O_2866,N_22495,N_23387);
nand UO_2867 (O_2867,N_22527,N_18868);
and UO_2868 (O_2868,N_23275,N_19441);
nand UO_2869 (O_2869,N_23340,N_19091);
nand UO_2870 (O_2870,N_23946,N_24390);
xor UO_2871 (O_2871,N_21622,N_22675);
xnor UO_2872 (O_2872,N_22094,N_19121);
nand UO_2873 (O_2873,N_19154,N_20773);
or UO_2874 (O_2874,N_20956,N_20567);
and UO_2875 (O_2875,N_19835,N_23700);
nor UO_2876 (O_2876,N_22095,N_18949);
or UO_2877 (O_2877,N_19238,N_21555);
nor UO_2878 (O_2878,N_23187,N_19904);
nor UO_2879 (O_2879,N_23242,N_24642);
and UO_2880 (O_2880,N_19036,N_21580);
or UO_2881 (O_2881,N_22988,N_21615);
nor UO_2882 (O_2882,N_23471,N_24616);
or UO_2883 (O_2883,N_24344,N_20564);
nand UO_2884 (O_2884,N_20632,N_24863);
or UO_2885 (O_2885,N_23611,N_24678);
nand UO_2886 (O_2886,N_20822,N_20768);
or UO_2887 (O_2887,N_19330,N_19134);
or UO_2888 (O_2888,N_19120,N_24741);
xor UO_2889 (O_2889,N_24385,N_24770);
xor UO_2890 (O_2890,N_22711,N_20767);
or UO_2891 (O_2891,N_19128,N_20916);
xnor UO_2892 (O_2892,N_24768,N_21075);
nand UO_2893 (O_2893,N_20706,N_20175);
or UO_2894 (O_2894,N_22807,N_23206);
nand UO_2895 (O_2895,N_24565,N_24967);
nor UO_2896 (O_2896,N_21972,N_23660);
and UO_2897 (O_2897,N_21945,N_21327);
nor UO_2898 (O_2898,N_21444,N_21204);
nand UO_2899 (O_2899,N_20209,N_21669);
xnor UO_2900 (O_2900,N_22632,N_23460);
nor UO_2901 (O_2901,N_19719,N_22275);
xor UO_2902 (O_2902,N_24163,N_19383);
nor UO_2903 (O_2903,N_19648,N_23781);
nand UO_2904 (O_2904,N_20702,N_24300);
nor UO_2905 (O_2905,N_21020,N_23571);
xor UO_2906 (O_2906,N_24458,N_19546);
nor UO_2907 (O_2907,N_22005,N_23533);
nand UO_2908 (O_2908,N_22231,N_22284);
nand UO_2909 (O_2909,N_23691,N_24652);
and UO_2910 (O_2910,N_19796,N_20683);
nand UO_2911 (O_2911,N_23075,N_21456);
or UO_2912 (O_2912,N_20230,N_19232);
xor UO_2913 (O_2913,N_20174,N_22518);
nand UO_2914 (O_2914,N_19691,N_23847);
xor UO_2915 (O_2915,N_20344,N_21838);
nand UO_2916 (O_2916,N_20864,N_18968);
nand UO_2917 (O_2917,N_24014,N_22428);
and UO_2918 (O_2918,N_24841,N_21531);
nand UO_2919 (O_2919,N_24146,N_22721);
nand UO_2920 (O_2920,N_24082,N_22547);
and UO_2921 (O_2921,N_24606,N_24399);
nor UO_2922 (O_2922,N_20607,N_21426);
and UO_2923 (O_2923,N_24860,N_23780);
nand UO_2924 (O_2924,N_20990,N_20184);
xor UO_2925 (O_2925,N_23834,N_24897);
xnor UO_2926 (O_2926,N_22524,N_22498);
nand UO_2927 (O_2927,N_19092,N_24993);
or UO_2928 (O_2928,N_20942,N_23066);
or UO_2929 (O_2929,N_19986,N_21280);
xor UO_2930 (O_2930,N_20903,N_21072);
xor UO_2931 (O_2931,N_19945,N_22691);
nor UO_2932 (O_2932,N_21029,N_24071);
nand UO_2933 (O_2933,N_20777,N_19826);
or UO_2934 (O_2934,N_23181,N_21751);
or UO_2935 (O_2935,N_22708,N_24357);
nor UO_2936 (O_2936,N_19779,N_23725);
or UO_2937 (O_2937,N_21082,N_23619);
and UO_2938 (O_2938,N_23915,N_23955);
nor UO_2939 (O_2939,N_18884,N_21797);
nand UO_2940 (O_2940,N_19955,N_23592);
nand UO_2941 (O_2941,N_20390,N_20035);
and UO_2942 (O_2942,N_19932,N_19820);
nand UO_2943 (O_2943,N_22626,N_20059);
or UO_2944 (O_2944,N_19411,N_24182);
or UO_2945 (O_2945,N_23879,N_24772);
and UO_2946 (O_2946,N_18826,N_19663);
nand UO_2947 (O_2947,N_24555,N_22191);
or UO_2948 (O_2948,N_20790,N_19666);
or UO_2949 (O_2949,N_22499,N_21952);
or UO_2950 (O_2950,N_22598,N_21524);
nand UO_2951 (O_2951,N_22785,N_24697);
nor UO_2952 (O_2952,N_21885,N_19126);
xor UO_2953 (O_2953,N_24350,N_21832);
xnor UO_2954 (O_2954,N_24341,N_23932);
or UO_2955 (O_2955,N_21586,N_24061);
nor UO_2956 (O_2956,N_22205,N_18797);
nor UO_2957 (O_2957,N_23096,N_22249);
nor UO_2958 (O_2958,N_22036,N_24323);
nor UO_2959 (O_2959,N_20474,N_22015);
nor UO_2960 (O_2960,N_20625,N_23779);
and UO_2961 (O_2961,N_24900,N_22337);
or UO_2962 (O_2962,N_23486,N_19375);
or UO_2963 (O_2963,N_21025,N_20791);
xnor UO_2964 (O_2964,N_21235,N_21522);
xor UO_2965 (O_2965,N_23810,N_18887);
xor UO_2966 (O_2966,N_23279,N_19239);
nand UO_2967 (O_2967,N_18930,N_24920);
xor UO_2968 (O_2968,N_22285,N_20880);
nand UO_2969 (O_2969,N_21741,N_21651);
or UO_2970 (O_2970,N_21465,N_19759);
xor UO_2971 (O_2971,N_23410,N_19323);
nor UO_2972 (O_2972,N_22611,N_22154);
and UO_2973 (O_2973,N_24100,N_20859);
and UO_2974 (O_2974,N_23092,N_21828);
nor UO_2975 (O_2975,N_20551,N_22503);
xnor UO_2976 (O_2976,N_21882,N_19807);
xor UO_2977 (O_2977,N_22893,N_19115);
nand UO_2978 (O_2978,N_23284,N_23808);
xnor UO_2979 (O_2979,N_19982,N_20176);
xor UO_2980 (O_2980,N_22818,N_22061);
nor UO_2981 (O_2981,N_19406,N_20704);
xor UO_2982 (O_2982,N_23898,N_20000);
and UO_2983 (O_2983,N_23230,N_20162);
nor UO_2984 (O_2984,N_20955,N_21900);
or UO_2985 (O_2985,N_23743,N_24030);
and UO_2986 (O_2986,N_21765,N_20514);
or UO_2987 (O_2987,N_23664,N_22712);
nor UO_2988 (O_2988,N_22406,N_24622);
or UO_2989 (O_2989,N_20496,N_19592);
nor UO_2990 (O_2990,N_22934,N_19845);
xor UO_2991 (O_2991,N_23762,N_20531);
nand UO_2992 (O_2992,N_23625,N_21406);
and UO_2993 (O_2993,N_21749,N_20170);
and UO_2994 (O_2994,N_23026,N_24169);
or UO_2995 (O_2995,N_20267,N_21330);
and UO_2996 (O_2996,N_23478,N_23067);
nor UO_2997 (O_2997,N_24218,N_24686);
or UO_2998 (O_2998,N_20290,N_18886);
or UO_2999 (O_2999,N_24668,N_22241);
endmodule