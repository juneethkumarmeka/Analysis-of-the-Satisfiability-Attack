module basic_2500_25000_3000_100_levels_1xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
nor U0 (N_0,In_1444,In_1892);
nand U1 (N_1,In_1685,In_729);
and U2 (N_2,In_679,In_2083);
nor U3 (N_3,In_1753,In_718);
nor U4 (N_4,In_1814,In_1445);
xor U5 (N_5,In_728,In_471);
nand U6 (N_6,In_1370,In_983);
nor U7 (N_7,In_882,In_670);
or U8 (N_8,In_1772,In_991);
nor U9 (N_9,In_2323,In_2229);
nor U10 (N_10,In_1475,In_154);
nand U11 (N_11,In_1851,In_1338);
nor U12 (N_12,In_2458,In_227);
nor U13 (N_13,In_9,In_1426);
or U14 (N_14,In_2173,In_74);
and U15 (N_15,In_862,In_1835);
and U16 (N_16,In_1183,In_594);
and U17 (N_17,In_1353,In_985);
nor U18 (N_18,In_1960,In_2187);
nor U19 (N_19,In_2484,In_1480);
nand U20 (N_20,In_1442,In_2223);
xor U21 (N_21,In_1800,In_1491);
nand U22 (N_22,In_1005,In_2071);
and U23 (N_23,In_1100,In_1189);
nor U24 (N_24,In_1429,In_2281);
nand U25 (N_25,In_2077,In_1257);
nor U26 (N_26,In_1381,In_977);
and U27 (N_27,In_2389,In_1948);
and U28 (N_28,In_1586,In_229);
nor U29 (N_29,In_327,In_158);
and U30 (N_30,In_2248,In_2125);
nand U31 (N_31,In_1090,In_2112);
nor U32 (N_32,In_1541,In_1282);
or U33 (N_33,In_1049,In_606);
or U34 (N_34,In_2217,In_2340);
nor U35 (N_35,In_222,In_736);
or U36 (N_36,In_1664,In_63);
nand U37 (N_37,In_156,In_1523);
nor U38 (N_38,In_1618,In_529);
nor U39 (N_39,In_1749,In_805);
nand U40 (N_40,In_799,In_909);
and U41 (N_41,In_896,In_1173);
nor U42 (N_42,In_2039,In_742);
nor U43 (N_43,In_1879,In_2275);
or U44 (N_44,In_972,In_331);
and U45 (N_45,In_1963,In_1050);
or U46 (N_46,In_1982,In_307);
nor U47 (N_47,In_1401,In_5);
nor U48 (N_48,In_548,In_1387);
or U49 (N_49,In_1743,In_635);
or U50 (N_50,In_1497,In_569);
nand U51 (N_51,In_1018,In_175);
nor U52 (N_52,In_145,In_276);
or U53 (N_53,In_2170,In_7);
or U54 (N_54,In_1791,In_1327);
and U55 (N_55,In_657,In_199);
nor U56 (N_56,In_2437,In_660);
or U57 (N_57,In_255,In_2249);
and U58 (N_58,In_2232,In_2407);
nor U59 (N_59,In_1680,In_1634);
or U60 (N_60,In_1230,In_1094);
nor U61 (N_61,In_565,In_1572);
nand U62 (N_62,In_1437,In_386);
or U63 (N_63,In_608,In_147);
nor U64 (N_64,In_1591,In_539);
nand U65 (N_65,In_1410,In_1767);
or U66 (N_66,In_2344,In_609);
and U67 (N_67,In_1862,In_837);
nand U68 (N_68,In_1638,In_2036);
or U69 (N_69,In_2098,In_2157);
or U70 (N_70,In_2369,In_1330);
nor U71 (N_71,In_686,In_2162);
or U72 (N_72,In_1253,In_1540);
and U73 (N_73,In_208,In_823);
and U74 (N_74,In_642,In_1885);
nand U75 (N_75,In_137,In_586);
nand U76 (N_76,In_500,In_1737);
nor U77 (N_77,In_1468,In_900);
and U78 (N_78,In_2226,In_1020);
nor U79 (N_79,In_727,In_1300);
and U80 (N_80,In_2104,In_1299);
nand U81 (N_81,In_211,In_1996);
nor U82 (N_82,In_563,In_814);
and U83 (N_83,In_2148,In_2424);
and U84 (N_84,In_1489,In_648);
and U85 (N_85,In_2449,In_2411);
or U86 (N_86,In_2183,In_1956);
or U87 (N_87,In_323,In_1110);
nor U88 (N_88,In_1361,In_1169);
or U89 (N_89,In_1708,In_2314);
nand U90 (N_90,In_730,In_1527);
nand U91 (N_91,In_2433,In_1555);
and U92 (N_92,In_1343,In_1718);
nor U93 (N_93,In_1348,In_2312);
nand U94 (N_94,In_38,In_1896);
and U95 (N_95,In_1212,In_152);
nor U96 (N_96,In_404,In_816);
or U97 (N_97,In_16,In_1735);
nor U98 (N_98,In_1726,In_481);
or U99 (N_99,In_1435,In_1219);
xnor U100 (N_100,In_2175,In_853);
nand U101 (N_101,In_1953,In_1817);
nor U102 (N_102,In_62,In_1380);
and U103 (N_103,In_334,In_891);
nor U104 (N_104,In_2485,In_1820);
nand U105 (N_105,In_1265,In_1962);
or U106 (N_106,In_680,In_975);
nor U107 (N_107,In_1287,In_895);
and U108 (N_108,In_1935,In_1310);
or U109 (N_109,In_644,In_1660);
nand U110 (N_110,In_1754,In_758);
and U111 (N_111,In_2499,In_993);
nand U112 (N_112,In_1436,In_2054);
or U113 (N_113,In_2295,In_960);
or U114 (N_114,In_583,In_631);
or U115 (N_115,In_782,In_478);
nor U116 (N_116,In_1509,In_982);
and U117 (N_117,In_913,In_1030);
nor U118 (N_118,In_1231,In_677);
nand U119 (N_119,In_1066,In_1121);
and U120 (N_120,In_501,In_1407);
nand U121 (N_121,In_2415,In_984);
nand U122 (N_122,In_1865,In_505);
and U123 (N_123,In_2368,In_626);
and U124 (N_124,In_1467,In_2438);
nor U125 (N_125,In_113,In_146);
nand U126 (N_126,In_2258,In_1195);
or U127 (N_127,In_1164,In_536);
or U128 (N_128,In_804,In_1929);
nand U129 (N_129,In_207,In_2075);
nand U130 (N_130,In_650,In_462);
nand U131 (N_131,In_1710,In_1432);
nor U132 (N_132,In_1829,In_1345);
nor U133 (N_133,In_952,In_301);
and U134 (N_134,In_2359,In_434);
or U135 (N_135,In_1803,In_1793);
nor U136 (N_136,In_885,In_2285);
or U137 (N_137,In_1071,In_160);
or U138 (N_138,In_1106,In_1796);
and U139 (N_139,In_1416,In_1887);
and U140 (N_140,In_1097,In_220);
and U141 (N_141,In_2302,In_2355);
or U142 (N_142,In_1010,In_224);
nor U143 (N_143,In_1850,In_511);
nor U144 (N_144,In_2114,In_1667);
nor U145 (N_145,In_1473,In_791);
nor U146 (N_146,In_1993,In_1304);
and U147 (N_147,In_1639,In_14);
nand U148 (N_148,In_1420,In_1730);
or U149 (N_149,In_1342,In_414);
or U150 (N_150,In_1611,In_912);
or U151 (N_151,In_1825,In_1021);
nor U152 (N_152,In_1248,In_1070);
and U153 (N_153,In_1715,In_636);
nand U154 (N_154,In_260,In_387);
nand U155 (N_155,In_504,In_369);
nand U156 (N_156,In_1549,In_1596);
nand U157 (N_157,In_56,In_1924);
or U158 (N_158,In_1252,In_1792);
nand U159 (N_159,In_2044,In_174);
nor U160 (N_160,In_2130,In_2284);
nand U161 (N_161,In_2043,In_1458);
and U162 (N_162,In_1209,In_70);
and U163 (N_163,In_325,In_614);
nor U164 (N_164,In_585,In_2230);
and U165 (N_165,In_1334,In_2047);
or U166 (N_166,In_920,In_690);
or U167 (N_167,In_1367,In_1014);
or U168 (N_168,In_1119,In_465);
nor U169 (N_169,In_272,In_1619);
or U170 (N_170,In_21,In_1606);
nor U171 (N_171,In_974,In_2108);
nor U172 (N_172,In_1970,In_1303);
or U173 (N_173,In_1315,In_946);
xnor U174 (N_174,In_218,In_2321);
nand U175 (N_175,In_1839,In_1723);
nand U176 (N_176,In_2236,In_820);
and U177 (N_177,In_477,In_1925);
nand U178 (N_178,In_1544,In_48);
nor U179 (N_179,In_1724,In_1980);
and U180 (N_180,In_305,In_710);
and U181 (N_181,In_2289,In_2427);
and U182 (N_182,In_1609,In_2416);
or U183 (N_183,In_1229,In_487);
and U184 (N_184,In_1856,In_130);
or U185 (N_185,In_405,In_1968);
nand U186 (N_186,In_1588,In_835);
nor U187 (N_187,In_1194,In_1125);
xnor U188 (N_188,In_2069,In_904);
or U189 (N_189,In_2028,In_676);
and U190 (N_190,In_696,In_1272);
nor U191 (N_191,In_148,In_1044);
and U192 (N_192,In_2,In_774);
nand U193 (N_193,In_338,In_163);
or U194 (N_194,In_1777,In_732);
nor U195 (N_195,In_1889,In_817);
or U196 (N_196,In_1156,In_185);
nor U197 (N_197,In_2124,In_776);
nor U198 (N_198,In_1823,In_1656);
nor U199 (N_199,In_202,In_2293);
and U200 (N_200,In_1494,In_197);
nor U201 (N_201,In_1613,In_1827);
and U202 (N_202,In_1919,In_2351);
nand U203 (N_203,In_294,In_470);
nand U204 (N_204,In_750,In_2441);
or U205 (N_205,In_2127,In_2270);
or U206 (N_206,In_859,In_1185);
nor U207 (N_207,In_528,In_808);
xor U208 (N_208,In_372,In_2430);
nand U209 (N_209,In_721,In_905);
nand U210 (N_210,In_298,In_926);
nor U211 (N_211,In_1648,In_1760);
nand U212 (N_212,In_1386,In_2345);
and U213 (N_213,In_671,In_1339);
nand U214 (N_214,In_664,In_1105);
or U215 (N_215,In_2330,In_2346);
nand U216 (N_216,In_884,In_2448);
or U217 (N_217,In_495,In_215);
nor U218 (N_218,In_362,In_1612);
nor U219 (N_219,In_1113,In_1716);
or U220 (N_220,In_140,In_928);
nor U221 (N_221,In_1075,In_577);
nand U222 (N_222,In_532,In_329);
or U223 (N_223,In_1412,In_99);
nand U224 (N_224,In_136,In_2471);
nor U225 (N_225,In_2360,In_1061);
nor U226 (N_226,In_2107,In_1806);
nor U227 (N_227,In_2474,In_2265);
or U228 (N_228,In_590,In_1936);
or U229 (N_229,In_393,In_770);
or U230 (N_230,In_291,In_1971);
and U231 (N_231,In_1251,In_385);
nor U232 (N_232,In_1199,In_360);
or U233 (N_233,In_392,In_625);
or U234 (N_234,In_1759,In_2166);
and U235 (N_235,In_1493,In_483);
nand U236 (N_236,In_903,In_653);
nand U237 (N_237,In_1439,In_964);
or U238 (N_238,In_1268,In_124);
nor U239 (N_239,In_411,In_430);
nor U240 (N_240,In_701,In_1693);
nor U241 (N_241,In_1376,In_2213);
and U242 (N_242,In_942,In_17);
nand U243 (N_243,In_2269,In_1262);
xnor U244 (N_244,In_2453,In_513);
nand U245 (N_245,In_872,In_1139);
or U246 (N_246,In_1686,In_2182);
and U247 (N_247,In_426,In_1898);
and U248 (N_248,In_1597,In_1720);
or U249 (N_249,In_2037,In_1765);
xor U250 (N_250,In_1868,In_269);
or U251 (N_251,In_1625,In_682);
or U252 (N_252,In_219,In_1312);
and U253 (N_253,In_76,N_98);
nand U254 (N_254,In_605,In_2201);
or U255 (N_255,In_1883,In_1488);
nand U256 (N_256,In_1949,N_135);
and U257 (N_257,N_247,In_268);
and U258 (N_258,In_901,In_877);
nor U259 (N_259,In_182,In_852);
or U260 (N_260,In_2451,In_2056);
nand U261 (N_261,In_1474,In_2325);
and U262 (N_262,N_111,In_2109);
nor U263 (N_263,In_2079,In_2397);
nor U264 (N_264,N_93,In_368);
nand U265 (N_265,In_1396,In_81);
xor U266 (N_266,In_2348,In_1564);
or U267 (N_267,In_2337,In_1688);
nand U268 (N_268,In_1174,In_166);
nor U269 (N_269,In_123,In_1039);
xnor U270 (N_270,In_951,In_1967);
and U271 (N_271,In_878,In_2385);
nor U272 (N_272,In_2349,In_345);
and U273 (N_273,In_1178,In_785);
or U274 (N_274,In_2417,In_15);
nand U275 (N_275,N_61,N_170);
or U276 (N_276,In_1787,In_1040);
nor U277 (N_277,In_812,In_1154);
nor U278 (N_278,In_1331,In_1866);
nor U279 (N_279,In_865,In_1502);
and U280 (N_280,In_748,In_2216);
nor U281 (N_281,In_560,In_422);
nand U282 (N_282,In_827,N_119);
and U283 (N_283,In_1166,In_969);
or U284 (N_284,In_973,In_1291);
nand U285 (N_285,N_57,In_1975);
and U286 (N_286,In_637,In_2381);
nor U287 (N_287,In_2222,In_86);
or U288 (N_288,N_183,In_64);
nand U289 (N_289,In_1114,In_1104);
nor U290 (N_290,In_856,N_68);
nand U291 (N_291,In_1908,In_2147);
nand U292 (N_292,In_1159,In_380);
and U293 (N_293,In_1500,In_1266);
nand U294 (N_294,In_1563,In_383);
or U295 (N_295,In_310,In_1860);
or U296 (N_296,In_285,In_1152);
nor U297 (N_297,N_226,In_674);
and U298 (N_298,In_1786,In_2080);
or U299 (N_299,In_1578,In_935);
and U300 (N_300,In_1292,In_1043);
or U301 (N_301,In_2167,In_1109);
and U302 (N_302,In_2008,In_1130);
or U303 (N_303,In_2200,In_2257);
nand U304 (N_304,N_21,In_2482);
or U305 (N_305,In_834,In_443);
or U306 (N_306,In_1200,In_1160);
nor U307 (N_307,In_1990,N_187);
and U308 (N_308,In_1031,In_1542);
or U309 (N_309,In_1550,In_464);
nand U310 (N_310,In_18,In_407);
or U311 (N_311,In_2189,In_436);
nor U312 (N_312,In_712,In_1214);
or U313 (N_313,In_1072,In_1873);
or U314 (N_314,In_297,In_641);
nand U315 (N_315,In_250,N_106);
nor U316 (N_316,In_1988,In_1831);
xnor U317 (N_317,In_1641,N_156);
or U318 (N_318,In_1546,In_668);
nor U319 (N_319,N_153,In_97);
nor U320 (N_320,In_1187,N_168);
and U321 (N_321,In_514,In_1145);
and U322 (N_322,In_2221,In_863);
and U323 (N_323,In_2252,In_1890);
nor U324 (N_324,In_745,In_1459);
nand U325 (N_325,In_1408,In_1208);
nor U326 (N_326,In_704,In_1559);
and U327 (N_327,In_246,In_1450);
nand U328 (N_328,In_328,In_122);
nor U329 (N_329,In_2101,In_1972);
nand U330 (N_330,In_1142,In_384);
nand U331 (N_331,N_129,N_193);
or U332 (N_332,In_1736,In_2191);
and U333 (N_333,In_1614,In_1143);
nor U334 (N_334,In_716,In_2146);
or U335 (N_335,In_242,In_2475);
or U336 (N_336,In_2404,In_1930);
or U337 (N_337,In_1966,In_1379);
nor U338 (N_338,In_181,In_2260);
nand U339 (N_339,In_601,In_2264);
nor U340 (N_340,N_17,In_1496);
nor U341 (N_341,In_225,In_2145);
nor U342 (N_342,N_120,In_1317);
and U343 (N_343,In_1676,In_1309);
and U344 (N_344,In_1276,In_1147);
and U345 (N_345,N_150,In_290);
or U346 (N_346,In_1854,In_444);
and U347 (N_347,In_555,In_779);
or U348 (N_348,In_206,In_1447);
nand U349 (N_349,In_1084,In_2025);
nand U350 (N_350,In_868,In_1964);
and U351 (N_351,In_1318,In_1914);
nor U352 (N_352,In_391,In_131);
nor U353 (N_353,In_1372,In_2116);
and U354 (N_354,In_3,In_1557);
or U355 (N_355,In_703,In_439);
or U356 (N_356,In_355,In_989);
nand U357 (N_357,In_1202,In_842);
and U358 (N_358,In_809,N_126);
and U359 (N_359,In_2082,In_1295);
or U360 (N_360,In_1934,In_825);
or U361 (N_361,In_82,In_2110);
or U362 (N_362,In_1623,In_1238);
nand U363 (N_363,In_2138,In_1547);
and U364 (N_364,In_1077,In_2081);
nand U365 (N_365,In_815,In_2306);
xor U366 (N_366,In_1654,In_1663);
and U367 (N_367,In_2324,In_1826);
or U368 (N_368,In_826,In_2185);
nand U369 (N_369,In_2280,In_2240);
nor U370 (N_370,In_153,In_342);
nor U371 (N_371,In_1533,In_2394);
nand U372 (N_372,In_2099,In_221);
or U373 (N_373,In_1283,In_956);
and U374 (N_374,In_2137,In_1670);
or U375 (N_375,In_2199,In_2378);
or U376 (N_376,N_124,In_1567);
nor U377 (N_377,In_949,In_1201);
and U378 (N_378,In_1080,In_1636);
nand U379 (N_379,In_1943,In_881);
nor U380 (N_380,In_2460,In_1645);
nand U381 (N_381,In_2472,In_8);
and U382 (N_382,In_171,In_1750);
and U383 (N_383,In_1362,In_603);
and U384 (N_384,In_2178,In_1583);
and U385 (N_385,In_1959,In_2095);
and U386 (N_386,In_883,N_2);
or U387 (N_387,In_2463,In_1816);
nand U388 (N_388,In_2245,In_2367);
nand U389 (N_389,In_802,In_1186);
or U390 (N_390,In_2418,In_10);
and U391 (N_391,In_1481,In_1780);
nor U392 (N_392,In_155,N_190);
nand U393 (N_393,In_1359,In_488);
xnor U394 (N_394,In_1004,N_207);
nand U395 (N_395,In_607,In_1514);
nand U396 (N_396,In_1234,In_358);
or U397 (N_397,In_223,N_77);
or U398 (N_398,In_2462,In_1841);
or U399 (N_399,In_236,In_1389);
nand U400 (N_400,In_1064,N_249);
or U401 (N_401,In_1076,In_249);
or U402 (N_402,N_155,In_1809);
nor U403 (N_403,In_1151,In_1569);
or U404 (N_404,In_1167,In_1390);
or U405 (N_405,In_1397,In_634);
nor U406 (N_406,In_424,In_1633);
nor U407 (N_407,In_1460,In_2131);
and U408 (N_408,In_1957,In_43);
or U409 (N_409,In_245,In_2168);
nand U410 (N_410,In_1595,In_2456);
nor U411 (N_411,In_335,N_27);
or U412 (N_412,In_2393,N_169);
or U413 (N_413,In_84,In_1504);
nor U414 (N_414,In_1894,In_1215);
and U415 (N_415,In_263,In_1037);
or U416 (N_416,In_1091,N_50);
and U417 (N_417,N_52,N_200);
or U418 (N_418,In_950,N_82);
nand U419 (N_419,In_506,In_1285);
nor U420 (N_420,In_2402,N_99);
nor U421 (N_421,In_1734,In_925);
or U422 (N_422,In_846,N_43);
nand U423 (N_423,In_1111,In_1979);
nor U424 (N_424,In_2057,In_1528);
and U425 (N_425,In_867,In_390);
or U426 (N_426,In_1867,N_37);
or U427 (N_427,In_2338,In_1337);
nand U428 (N_428,N_242,In_1653);
nor U429 (N_429,In_917,In_573);
or U430 (N_430,In_797,In_685);
nor U431 (N_431,In_1096,In_708);
nand U432 (N_432,In_1794,In_1373);
or U433 (N_433,In_2007,In_1392);
nor U434 (N_434,In_304,In_987);
nand U435 (N_435,In_1269,In_34);
nand U436 (N_436,In_406,N_53);
nor U437 (N_437,In_1950,In_1742);
and U438 (N_438,In_2012,In_1484);
nor U439 (N_439,In_1274,N_221);
nor U440 (N_440,In_1244,In_2136);
nor U441 (N_441,N_10,In_1587);
or U442 (N_442,In_1700,In_1994);
nand U443 (N_443,In_1329,N_26);
nor U444 (N_444,In_1007,In_916);
and U445 (N_445,In_446,In_420);
and U446 (N_446,In_1297,In_887);
and U447 (N_447,In_33,In_188);
or U448 (N_448,In_1086,In_1466);
nor U449 (N_449,In_700,In_1340);
and U450 (N_450,In_1526,In_1344);
and U451 (N_451,In_365,In_556);
nand U452 (N_452,N_133,In_2003);
nor U453 (N_453,In_36,In_1270);
nand U454 (N_454,In_274,In_2205);
and U455 (N_455,In_597,In_1400);
nor U456 (N_456,In_2273,In_308);
nor U457 (N_457,In_1910,In_538);
nand U458 (N_458,In_747,In_1989);
and U459 (N_459,In_1594,In_2015);
nand U460 (N_460,In_695,N_215);
or U461 (N_461,N_4,In_1844);
or U462 (N_462,In_2254,In_2141);
or U463 (N_463,In_2291,In_24);
and U464 (N_464,In_1864,In_2180);
nand U465 (N_465,N_186,In_1477);
nor U466 (N_466,In_1592,In_1954);
and U467 (N_467,In_715,In_2429);
nand U468 (N_468,In_512,In_1560);
nand U469 (N_469,In_621,N_139);
and U470 (N_470,In_798,In_684);
nor U471 (N_471,In_2172,In_1748);
nand U472 (N_472,In_413,In_720);
nor U473 (N_473,N_180,In_738);
nand U474 (N_474,In_1657,In_492);
and U475 (N_475,In_1088,In_1647);
nand U476 (N_476,In_1635,In_1768);
nand U477 (N_477,In_2212,In_402);
nand U478 (N_478,In_1699,In_1247);
nand U479 (N_479,N_210,In_1981);
nand U480 (N_480,N_87,In_1242);
or U481 (N_481,In_1776,In_2431);
or U482 (N_482,In_1045,In_936);
and U483 (N_483,N_90,In_2331);
or U484 (N_484,In_1947,In_1893);
or U485 (N_485,In_2089,In_994);
or U486 (N_486,In_428,In_523);
nand U487 (N_487,In_1384,N_178);
and U488 (N_488,In_652,In_499);
or U489 (N_489,In_1706,N_195);
nand U490 (N_490,In_1068,In_203);
and U491 (N_491,In_114,In_2203);
and U492 (N_492,In_602,In_819);
nor U493 (N_493,In_1374,In_1323);
nor U494 (N_494,In_2476,In_2084);
nand U495 (N_495,In_1746,N_11);
nor U496 (N_496,In_22,In_522);
nor U497 (N_497,In_1079,In_2048);
and U498 (N_498,N_159,In_697);
and U499 (N_499,In_1554,In_1168);
nor U500 (N_500,In_755,In_125);
and U501 (N_501,In_1690,N_66);
and U502 (N_502,In_1757,In_157);
nand U503 (N_503,In_2400,In_1225);
and U504 (N_504,In_611,In_2494);
nor U505 (N_505,In_1226,N_483);
nor U506 (N_506,In_367,In_1192);
nand U507 (N_507,In_1525,In_2313);
or U508 (N_508,In_194,In_655);
nand U509 (N_509,N_161,In_1267);
and U510 (N_510,In_1858,N_166);
and U511 (N_511,In_1355,In_1115);
and U512 (N_512,In_2126,In_265);
nand U513 (N_513,In_1552,N_216);
or U514 (N_514,In_1599,N_315);
or U515 (N_515,In_2480,In_1324);
nor U516 (N_516,In_1575,In_450);
and U517 (N_517,In_1171,N_20);
and U518 (N_518,In_1872,In_1172);
and U519 (N_519,In_731,In_879);
nand U520 (N_520,In_2297,In_264);
nor U521 (N_521,In_1246,In_1665);
or U522 (N_522,In_180,In_2238);
and U523 (N_523,In_37,In_266);
and U524 (N_524,N_339,In_337);
and U525 (N_525,In_1524,In_2005);
nor U526 (N_526,N_110,In_61);
nand U527 (N_527,N_160,N_105);
nand U528 (N_528,In_1505,In_1775);
or U529 (N_529,In_571,In_2498);
nor U530 (N_530,N_205,In_666);
nand U531 (N_531,N_112,In_875);
or U532 (N_532,In_2318,In_2392);
nand U533 (N_533,In_2414,In_2023);
and U534 (N_534,In_1409,In_618);
or U535 (N_535,In_103,In_109);
nor U536 (N_536,In_1519,N_312);
nor U537 (N_537,In_1406,In_57);
and U538 (N_538,In_2488,In_1469);
and U539 (N_539,In_1607,In_2163);
and U540 (N_540,In_940,In_1048);
and U541 (N_541,In_1023,In_353);
and U542 (N_542,In_448,In_475);
xnor U543 (N_543,N_97,In_669);
nand U544 (N_544,N_464,In_1678);
nand U545 (N_545,In_1601,In_1616);
or U546 (N_546,In_287,In_1713);
nand U547 (N_547,In_1150,In_992);
and U548 (N_548,In_1236,In_2466);
and U549 (N_549,In_948,In_340);
and U550 (N_550,N_410,In_2492);
nand U551 (N_551,In_2202,In_1570);
nor U552 (N_552,In_1180,In_723);
nor U553 (N_553,In_2422,In_2158);
and U554 (N_554,N_74,In_1932);
or U555 (N_555,In_12,In_459);
and U556 (N_556,N_348,In_2432);
nand U557 (N_557,In_1313,N_293);
or U558 (N_558,In_639,In_2059);
or U559 (N_559,In_1629,In_646);
nor U560 (N_560,In_159,N_15);
nand U561 (N_561,In_2255,In_1637);
and U562 (N_562,In_117,N_344);
nand U563 (N_563,In_1643,In_1141);
or U564 (N_564,N_274,In_510);
nor U565 (N_565,In_1188,In_1148);
nand U566 (N_566,In_786,In_1221);
nand U567 (N_567,In_2395,In_1499);
nand U568 (N_568,In_2467,In_1237);
nand U569 (N_569,In_1728,In_189);
nor U570 (N_570,In_210,In_161);
nand U571 (N_571,In_2053,In_2469);
and U572 (N_572,N_229,In_1882);
nor U573 (N_573,In_2020,In_1454);
nand U574 (N_574,In_1778,In_1316);
nand U575 (N_575,In_1937,In_1632);
and U576 (N_576,In_129,N_404);
nor U577 (N_577,In_1440,In_300);
nor U578 (N_578,In_1912,In_1709);
nor U579 (N_579,In_1598,In_463);
nor U580 (N_580,In_1405,In_1871);
nand U581 (N_581,N_426,N_313);
and U582 (N_582,In_2380,In_1204);
nand U583 (N_583,N_146,In_1053);
or U584 (N_584,In_1157,In_2320);
and U585 (N_585,In_711,In_2237);
and U586 (N_586,In_2019,In_910);
nand U587 (N_587,In_662,N_488);
nand U588 (N_588,N_377,In_1581);
or U589 (N_589,In_1608,In_410);
and U590 (N_590,In_550,In_183);
nand U591 (N_591,In_1877,In_2063);
nor U592 (N_592,In_412,In_1888);
nor U593 (N_593,In_292,In_541);
nand U594 (N_594,In_1574,In_1969);
nor U595 (N_595,N_40,In_485);
nand U596 (N_596,In_2244,In_319);
and U597 (N_597,N_319,In_1245);
and U598 (N_598,In_191,In_2375);
or U599 (N_599,In_719,In_1307);
or U600 (N_600,In_2154,N_291);
nand U601 (N_601,In_1207,In_469);
or U602 (N_602,In_1443,In_2086);
or U603 (N_603,In_1056,In_1741);
or U604 (N_604,In_2434,In_2310);
or U605 (N_605,N_497,In_1103);
or U606 (N_606,In_1874,In_2224);
nand U607 (N_607,In_2461,In_2235);
and U608 (N_608,N_9,In_930);
nand U609 (N_609,In_1941,In_282);
or U610 (N_610,In_735,N_349);
nand U611 (N_611,In_316,In_1320);
and U612 (N_612,In_1876,In_2401);
nor U613 (N_613,N_5,N_417);
nor U614 (N_614,In_841,In_1089);
and U615 (N_615,In_2118,In_1811);
and U616 (N_616,N_384,N_199);
and U617 (N_617,In_1170,In_1177);
or U618 (N_618,In_2220,In_1027);
or U619 (N_619,In_839,In_172);
and U620 (N_620,In_89,N_309);
or U621 (N_621,In_880,In_235);
nand U622 (N_622,In_963,In_1293);
nand U623 (N_623,N_397,In_1511);
and U624 (N_624,In_2040,In_279);
nand U625 (N_625,In_1744,In_143);
nor U626 (N_626,In_850,In_788);
nand U627 (N_627,In_2061,In_401);
or U628 (N_628,In_1828,In_1074);
or U629 (N_629,In_516,N_362);
nand U630 (N_630,In_627,N_285);
or U631 (N_631,In_2423,In_1356);
nor U632 (N_632,In_1536,In_419);
nand U633 (N_633,In_661,In_302);
and U634 (N_634,In_1456,In_1411);
nand U635 (N_635,In_1273,N_296);
nand U636 (N_636,In_2408,N_6);
nand U637 (N_637,N_364,In_766);
and U638 (N_638,In_416,N_172);
nand U639 (N_639,N_423,In_168);
nor U640 (N_640,N_342,N_197);
xor U641 (N_641,In_1891,In_1235);
nand U642 (N_642,In_1849,N_22);
nand U643 (N_643,In_1548,N_374);
and U644 (N_644,N_301,N_103);
nand U645 (N_645,In_2156,In_293);
nand U646 (N_646,In_2210,N_367);
nor U647 (N_647,N_174,In_1217);
nor U648 (N_648,In_149,In_1184);
or U649 (N_649,In_138,In_2479);
and U650 (N_650,In_898,In_1986);
nand U651 (N_651,In_1462,N_85);
and U652 (N_652,In_1158,N_248);
nand U653 (N_653,N_101,In_2305);
and U654 (N_654,In_240,In_2342);
and U655 (N_655,In_1652,N_3);
and U656 (N_656,In_2115,In_1498);
or U657 (N_657,In_1673,In_437);
and U658 (N_658,In_108,In_1193);
and U659 (N_659,In_1624,In_127);
and U660 (N_660,In_1264,N_176);
and U661 (N_661,In_1719,N_388);
and U662 (N_662,N_496,In_2328);
or U663 (N_663,N_329,In_1062);
nor U664 (N_664,In_1280,In_1995);
nand U665 (N_665,In_540,In_1375);
or U666 (N_666,In_112,In_795);
or U667 (N_667,In_1565,In_692);
nand U668 (N_668,In_1510,N_380);
and U669 (N_669,In_78,In_1848);
and U670 (N_670,N_450,In_1319);
or U671 (N_671,In_1093,In_2074);
and U672 (N_672,In_1646,In_651);
nor U673 (N_673,In_997,In_73);
nand U674 (N_674,In_352,In_1046);
or U675 (N_675,In_2287,N_485);
or U676 (N_676,In_1294,In_248);
or U677 (N_677,In_2420,In_604);
or U678 (N_678,In_79,In_1082);
nor U679 (N_679,N_182,In_2117);
or U680 (N_680,In_858,In_2139);
or U681 (N_681,In_1102,In_496);
and U682 (N_682,In_2261,In_722);
nand U683 (N_683,In_237,In_1058);
or U684 (N_684,In_1991,In_1537);
or U685 (N_685,In_400,In_1913);
nor U686 (N_686,N_254,In_1026);
and U687 (N_687,In_1666,In_134);
or U688 (N_688,In_111,In_239);
nor U689 (N_689,N_225,In_1855);
and U690 (N_690,In_957,N_206);
nor U691 (N_691,In_790,In_1674);
nor U692 (N_692,In_1205,In_1732);
nor U693 (N_693,In_2317,In_1092);
nor U694 (N_694,In_1393,In_100);
and U695 (N_695,In_1335,In_1958);
nand U696 (N_696,In_2022,In_733);
or U697 (N_697,N_29,N_86);
or U698 (N_698,In_768,N_165);
nand U699 (N_699,In_2102,In_275);
or U700 (N_700,In_1368,In_53);
and U701 (N_701,In_442,In_1222);
and U702 (N_702,N_23,In_2206);
and U703 (N_703,N_7,In_1717);
and U704 (N_704,In_939,In_568);
or U705 (N_705,N_157,In_1782);
nand U706 (N_706,In_2027,In_1847);
nor U707 (N_707,In_2473,In_232);
nor U708 (N_708,In_2058,In_1600);
or U709 (N_709,In_1197,In_1261);
or U710 (N_710,In_2179,N_211);
nor U711 (N_711,In_306,In_961);
nand U712 (N_712,In_106,In_714);
or U713 (N_713,In_796,In_0);
nand U714 (N_714,In_549,N_34);
nor U715 (N_715,N_73,In_552);
and U716 (N_716,N_326,N_48);
or U717 (N_717,N_487,In_2169);
and U718 (N_718,In_941,In_2177);
nand U719 (N_719,In_320,N_484);
or U720 (N_720,N_454,N_435);
or U721 (N_721,In_986,N_36);
nor U722 (N_722,In_277,In_2491);
and U723 (N_723,In_610,N_212);
nand U724 (N_724,In_32,N_389);
nand U725 (N_725,In_2309,N_439);
nor U726 (N_726,In_2308,In_92);
and U727 (N_727,In_558,N_42);
and U728 (N_728,N_321,In_1210);
or U729 (N_729,In_51,In_1859);
nor U730 (N_730,In_574,In_2365);
nor U731 (N_731,In_1668,In_899);
or U732 (N_732,In_980,In_2192);
and U733 (N_733,N_456,N_420);
nor U734 (N_734,In_2149,In_2364);
and U735 (N_735,N_403,In_1306);
nand U736 (N_736,N_441,In_1041);
or U737 (N_737,In_1642,In_1692);
or U738 (N_738,In_544,In_2171);
nand U739 (N_739,In_295,In_2428);
nor U740 (N_740,In_1179,In_1655);
nor U741 (N_741,In_1438,In_35);
and U742 (N_742,In_2135,In_1707);
nor U743 (N_743,N_368,In_317);
xnor U744 (N_744,In_1465,In_2303);
or U745 (N_745,In_120,In_1880);
nand U746 (N_746,In_1824,In_1290);
nor U747 (N_747,N_267,In_760);
or U748 (N_748,In_1107,N_140);
nand U749 (N_749,In_864,N_239);
or U750 (N_750,In_314,N_705);
nor U751 (N_751,In_2078,N_76);
or U752 (N_752,In_491,N_350);
nor U753 (N_753,In_1976,N_709);
or U754 (N_754,N_578,In_2376);
nor U755 (N_755,In_230,In_2464);
and U756 (N_756,N_263,In_200);
or U757 (N_757,N_280,N_286);
and U758 (N_758,In_165,N_698);
nor U759 (N_759,In_2113,In_1243);
nand U760 (N_760,In_1131,In_2207);
nand U761 (N_761,N_638,In_1789);
or U762 (N_762,N_394,In_2153);
nor U763 (N_763,N_532,In_2165);
nand U764 (N_764,N_516,In_461);
nor U765 (N_765,In_135,In_1999);
and U766 (N_766,N_446,N_656);
or U767 (N_767,In_893,In_519);
nand U768 (N_768,In_85,In_58);
and U769 (N_769,N_398,In_915);
nand U770 (N_770,N_272,In_440);
or U771 (N_771,In_449,In_2133);
or U772 (N_772,In_962,In_833);
and U773 (N_773,In_1378,In_322);
or U774 (N_774,In_2271,N_524);
and U775 (N_775,In_1905,In_1227);
and U776 (N_776,N_575,In_169);
or U777 (N_777,N_565,N_259);
nand U778 (N_778,N_664,In_409);
or U779 (N_779,N_619,In_1669);
and U780 (N_780,In_1132,In_1819);
or U781 (N_781,In_47,In_2386);
nor U782 (N_782,In_2070,N_412);
nand U783 (N_783,In_2218,N_593);
nand U784 (N_784,N_651,In_789);
or U785 (N_785,In_1321,In_894);
nand U786 (N_786,N_655,In_115);
or U787 (N_787,In_821,In_2327);
nand U788 (N_788,In_1886,In_2193);
or U789 (N_789,N_277,In_1923);
nand U790 (N_790,N_151,N_71);
nor U791 (N_791,In_562,In_1833);
nor U792 (N_792,N_554,In_2215);
nand U793 (N_793,In_2354,In_1233);
or U794 (N_794,In_1672,In_681);
and U795 (N_795,In_83,In_508);
nand U796 (N_796,In_643,N_538);
or U797 (N_797,In_1684,In_1228);
nand U798 (N_798,In_2164,N_594);
nor U799 (N_799,N_588,In_2403);
or U800 (N_800,In_1946,N_503);
and U801 (N_801,In_2335,In_1363);
or U802 (N_802,N_617,In_1047);
and U803 (N_803,In_1211,In_330);
nand U804 (N_804,In_1843,In_69);
nor U805 (N_805,N_270,In_1101);
and U806 (N_806,In_1453,In_2299);
nor U807 (N_807,In_871,N_693);
or U808 (N_808,N_515,In_2362);
and U809 (N_809,N_741,In_1479);
and U810 (N_810,N_508,In_874);
or U811 (N_811,N_500,In_2497);
nand U812 (N_812,N_148,N_712);
nor U813 (N_813,N_678,In_1729);
nand U814 (N_814,In_1365,N_569);
nor U815 (N_815,N_455,N_611);
nand U816 (N_816,N_640,N_306);
xnor U817 (N_817,In_1842,N_391);
nor U818 (N_818,In_1118,In_923);
and U819 (N_819,N_231,N_616);
nor U820 (N_820,N_333,In_2487);
or U821 (N_821,In_170,In_1942);
or U822 (N_822,In_1446,N_316);
or U823 (N_823,N_490,In_141);
or U824 (N_824,N_252,In_581);
xnor U825 (N_825,In_479,N_580);
nor U826 (N_826,In_1116,In_28);
nor U827 (N_827,In_547,In_1945);
nor U828 (N_828,N_250,In_2024);
nand U829 (N_829,In_192,In_772);
nand U830 (N_830,N_223,In_1371);
xor U831 (N_831,N_521,N_537);
and U832 (N_832,In_589,N_662);
nor U833 (N_833,In_31,In_1901);
nand U834 (N_834,N_539,N_523);
nor U835 (N_835,N_445,In_1059);
or U836 (N_836,In_1259,In_2443);
nand U837 (N_837,In_1769,In_1579);
nand U838 (N_838,In_2159,In_873);
and U839 (N_839,In_654,N_224);
and U840 (N_840,In_1697,In_1562);
nor U841 (N_841,In_281,In_2493);
nand U842 (N_842,In_1347,N_675);
or U843 (N_843,In_151,In_178);
and U844 (N_844,In_2292,In_630);
and U845 (N_845,In_922,In_2014);
nor U846 (N_846,In_1032,N_354);
nand U847 (N_847,In_286,N_365);
nand U848 (N_848,In_1752,In_2276);
nand U849 (N_849,In_2259,In_1120);
xnor U850 (N_850,In_1928,In_1175);
nand U851 (N_851,In_1852,N_630);
nor U852 (N_852,In_39,In_2026);
nand U853 (N_853,N_191,In_2119);
nand U854 (N_854,In_1539,In_698);
nor U855 (N_855,In_2470,In_119);
nor U856 (N_856,N_620,In_234);
nor U857 (N_857,In_1651,N_748);
and U858 (N_858,In_104,In_1098);
or U859 (N_859,In_1766,In_1483);
nor U860 (N_860,N_89,N_560);
nand U861 (N_861,In_375,In_551);
nand U862 (N_862,In_806,In_1689);
nand U863 (N_863,In_27,In_665);
or U864 (N_864,In_1917,In_2174);
and U865 (N_865,In_313,In_1627);
and U866 (N_866,N_407,In_1576);
nand U867 (N_867,In_2060,N_722);
and U868 (N_868,In_1133,In_2439);
nand U869 (N_869,In_1922,N_577);
nand U870 (N_870,In_1626,In_190);
nand U871 (N_871,In_1921,N_311);
nand U872 (N_872,In_2097,In_2405);
nand U873 (N_873,N_147,N_720);
and U874 (N_874,In_699,N_547);
and U875 (N_875,In_503,N_444);
or U876 (N_876,In_599,In_2017);
nor U877 (N_877,In_520,N_305);
or U878 (N_878,N_715,In_781);
and U879 (N_879,In_2446,In_1558);
nand U880 (N_880,N_241,In_2004);
nor U881 (N_881,In_1610,In_934);
or U882 (N_882,In_2256,In_1305);
nor U883 (N_883,N_427,N_498);
nor U884 (N_884,N_647,In_793);
and U885 (N_885,In_341,N_41);
or U886 (N_886,In_1512,In_1006);
or U887 (N_887,In_2274,N_395);
nand U888 (N_888,In_658,In_1781);
and U889 (N_889,N_385,In_954);
nor U890 (N_890,In_408,In_374);
nand U891 (N_891,N_55,In_1617);
nand U892 (N_892,In_1899,In_588);
nor U893 (N_893,In_2246,N_240);
nand U894 (N_894,In_1836,In_754);
and U895 (N_895,N_24,N_727);
or U896 (N_896,N_94,In_656);
nor U897 (N_897,N_411,In_2227);
and U898 (N_898,In_1784,In_1182);
and U899 (N_899,In_537,In_557);
or U900 (N_900,In_489,In_1907);
nor U901 (N_901,In_1518,In_848);
and U902 (N_902,In_2300,N_453);
or U903 (N_903,N_54,In_1695);
nor U904 (N_904,N_665,In_584);
nor U905 (N_905,In_1470,N_1);
and U906 (N_906,N_409,In_417);
or U907 (N_907,N_134,In_1577);
nand U908 (N_908,N_589,N_265);
and U909 (N_909,In_622,In_1933);
nor U910 (N_910,In_1140,In_1455);
nor U911 (N_911,N_341,N_707);
and U912 (N_912,In_553,In_1350);
nor U913 (N_913,In_1325,In_564);
nand U914 (N_914,In_217,N_458);
nor U915 (N_915,In_484,In_198);
or U916 (N_916,In_468,In_927);
and U917 (N_917,In_1818,In_2387);
xnor U918 (N_918,In_693,In_1808);
nand U919 (N_919,N_230,In_1822);
and U920 (N_920,N_431,In_167);
and U921 (N_921,In_2412,In_2065);
nand U922 (N_922,In_2050,N_19);
or U923 (N_923,In_1687,In_1284);
or U924 (N_924,N_649,N_428);
and U925 (N_925,In_1366,In_2347);
or U926 (N_926,N_735,In_753);
nand U927 (N_927,In_1431,N_713);
xnor U928 (N_928,N_332,N_80);
xnor U929 (N_929,In_531,In_2352);
nor U930 (N_930,In_1834,N_213);
or U931 (N_931,N_448,In_339);
and U932 (N_932,N_300,N_227);
or U933 (N_933,N_38,In_2329);
or U934 (N_934,In_1801,N_466);
and U935 (N_935,In_828,In_1584);
nor U936 (N_936,N_360,In_2105);
nand U937 (N_937,N_196,In_1662);
nor U938 (N_938,In_1452,In_628);
nor U939 (N_939,N_452,In_1449);
nand U940 (N_940,In_2382,N_680);
xnor U941 (N_941,In_243,In_431);
and U942 (N_942,In_1659,N_728);
nand U943 (N_943,In_205,In_1582);
nor U944 (N_944,In_1181,In_1810);
xnor U945 (N_945,In_1155,In_75);
or U946 (N_946,N_615,In_379);
nor U947 (N_947,In_351,In_482);
and U948 (N_948,N_214,In_72);
nand U949 (N_949,N_257,N_408);
nor U950 (N_950,In_2419,N_607);
and U951 (N_951,N_461,In_1534);
or U952 (N_952,In_1063,In_88);
or U953 (N_953,In_241,In_1112);
or U954 (N_954,In_20,In_1503);
nand U955 (N_955,N_122,N_67);
or U956 (N_956,N_415,In_2445);
nor U957 (N_957,N_481,In_924);
nor U958 (N_958,N_232,In_1807);
or U959 (N_959,N_744,In_1232);
nand U960 (N_960,N_478,In_2134);
or U961 (N_961,In_947,In_1903);
nor U962 (N_962,In_388,In_533);
and U963 (N_963,N_108,N_299);
and U964 (N_964,In_1138,N_359);
or U965 (N_965,In_1190,N_123);
nand U966 (N_966,In_354,In_1275);
nand U967 (N_967,N_566,In_1395);
nor U968 (N_968,In_1779,N_708);
and U969 (N_969,In_1940,N_534);
or U970 (N_970,N_666,In_694);
and U971 (N_971,In_344,In_326);
or U972 (N_972,N_245,In_394);
nor U973 (N_973,N_609,N_702);
xor U974 (N_974,In_2421,In_777);
or U975 (N_975,In_2140,In_2262);
nor U976 (N_976,N_525,In_364);
or U977 (N_977,In_1545,In_2370);
or U978 (N_978,N_681,In_2336);
and U979 (N_979,N_46,In_1902);
nor U980 (N_980,N_472,In_445);
nor U981 (N_981,In_1054,In_2068);
and U982 (N_982,In_472,N_236);
nor U983 (N_983,N_235,In_1961);
nor U984 (N_984,N_266,In_247);
or U985 (N_985,In_1939,N_663);
and U986 (N_986,In_1992,In_474);
nor U987 (N_987,In_1428,In_1424);
or U988 (N_988,N_468,In_1938);
nand U989 (N_989,N_660,N_127);
nand U990 (N_990,N_184,In_1196);
or U991 (N_991,In_212,In_2103);
and U992 (N_992,In_1258,N_402);
nor U993 (N_993,In_2319,In_454);
nor U994 (N_994,In_177,N_533);
and U995 (N_995,In_2106,N_683);
nor U996 (N_996,N_204,N_202);
and U997 (N_997,N_512,N_401);
nand U998 (N_998,In_1821,In_1035);
nor U999 (N_999,In_382,N_320);
or U1000 (N_1000,N_691,In_216);
and U1001 (N_1001,In_673,N_883);
nand U1002 (N_1002,N_102,N_731);
and U1003 (N_1003,In_1213,In_1308);
nor U1004 (N_1004,In_2034,In_288);
or U1005 (N_1005,In_309,N_668);
or U1006 (N_1006,In_2247,N_429);
or U1007 (N_1007,In_490,In_870);
and U1008 (N_1008,In_769,In_2251);
nand U1009 (N_1009,In_1476,In_2243);
nor U1010 (N_1010,N_482,N_998);
nand U1011 (N_1011,N_657,N_430);
or U1012 (N_1012,In_845,In_613);
and U1013 (N_1013,In_2478,In_1771);
and U1014 (N_1014,N_279,In_1531);
nand U1015 (N_1015,In_2442,N_527);
nor U1016 (N_1016,N_701,In_186);
and U1017 (N_1017,In_1127,In_633);
nor U1018 (N_1018,In_2018,In_932);
or U1019 (N_1019,In_13,In_2011);
nand U1020 (N_1020,In_886,N_506);
and U1021 (N_1021,N_318,In_752);
nand U1022 (N_1022,In_460,N_171);
nor U1023 (N_1023,N_421,In_1383);
nor U1024 (N_1024,N_967,N_562);
nor U1025 (N_1025,N_872,N_473);
nand U1026 (N_1026,In_176,In_1738);
nor U1027 (N_1027,In_800,N_572);
nand U1028 (N_1028,In_629,N_298);
or U1029 (N_1029,N_70,In_128);
nor U1030 (N_1030,In_378,In_2073);
nand U1031 (N_1031,In_1521,In_822);
nand U1032 (N_1032,In_395,N_773);
or U1033 (N_1033,In_49,N_623);
and U1034 (N_1034,N_400,In_1915);
or U1035 (N_1035,In_179,N_81);
nand U1036 (N_1036,N_353,N_747);
nand U1037 (N_1037,N_813,N_697);
or U1038 (N_1038,In_2350,In_1418);
nor U1039 (N_1039,In_843,In_1589);
or U1040 (N_1040,N_564,In_582);
nand U1041 (N_1041,N_983,In_311);
nor U1042 (N_1042,In_1762,In_2435);
nor U1043 (N_1043,In_1920,N_672);
and U1044 (N_1044,N_757,N_625);
and U1045 (N_1045,N_938,In_687);
nand U1046 (N_1046,N_463,N_898);
or U1047 (N_1047,N_203,In_376);
nor U1048 (N_1048,In_415,N_966);
nor U1049 (N_1049,N_601,In_2161);
nor U1050 (N_1050,N_502,In_1884);
nor U1051 (N_1051,In_348,N_871);
xor U1052 (N_1052,N_810,N_778);
or U1053 (N_1053,N_600,N_626);
and U1054 (N_1054,In_592,In_888);
nor U1055 (N_1055,N_896,In_2142);
or U1056 (N_1056,In_734,N_958);
nor U1057 (N_1057,In_1224,N_476);
nor U1058 (N_1058,In_2121,N_686);
or U1059 (N_1059,In_150,N_803);
or U1060 (N_1060,In_1288,In_2152);
or U1061 (N_1061,In_911,N_219);
and U1062 (N_1062,N_923,In_2272);
nor U1063 (N_1063,N_694,N_642);
nand U1064 (N_1064,In_1364,N_598);
nand U1065 (N_1065,N_246,In_1802);
xor U1066 (N_1066,N_700,N_823);
and U1067 (N_1067,In_1840,In_1790);
nand U1068 (N_1068,In_914,In_452);
nor U1069 (N_1069,N_646,In_746);
or U1070 (N_1070,In_1568,In_1298);
nand U1071 (N_1071,In_196,N_866);
or U1072 (N_1072,N_836,In_756);
and U1073 (N_1073,In_1832,N_635);
and U1074 (N_1074,In_377,N_62);
or U1075 (N_1075,In_254,In_566);
and U1076 (N_1076,In_849,In_1529);
and U1077 (N_1077,N_807,In_2021);
or U1078 (N_1078,N_31,N_767);
or U1079 (N_1079,In_312,In_1277);
nand U1080 (N_1080,N_379,In_133);
nor U1081 (N_1081,N_605,N_338);
nor U1082 (N_1082,In_2111,In_2425);
or U1083 (N_1083,N_820,N_418);
nand U1084 (N_1084,N_158,N_844);
nand U1085 (N_1085,In_1691,In_466);
nor U1086 (N_1086,N_437,In_1918);
and U1087 (N_1087,In_2409,In_267);
nor U1088 (N_1088,In_737,In_1804);
and U1089 (N_1089,N_739,In_1073);
nand U1090 (N_1090,N_703,N_785);
nor U1091 (N_1091,In_2304,In_1538);
nand U1092 (N_1092,N_479,N_530);
or U1093 (N_1093,N_770,In_1441);
and U1094 (N_1094,N_121,N_927);
nor U1095 (N_1095,In_683,In_1733);
nand U1096 (N_1096,In_515,N_520);
nand U1097 (N_1097,N_835,In_1351);
and U1098 (N_1098,N_878,N_981);
and U1099 (N_1099,N_511,In_526);
nor U1100 (N_1100,In_2377,N_451);
nor U1101 (N_1101,In_1711,N_841);
and U1102 (N_1102,In_2253,N_854);
nand U1103 (N_1103,In_2150,In_517);
or U1104 (N_1104,N_969,In_252);
nor U1105 (N_1105,In_2013,N_874);
and U1106 (N_1106,In_2490,N_676);
nand U1107 (N_1107,In_706,N_509);
or U1108 (N_1108,In_1805,In_1788);
or U1109 (N_1109,In_2301,In_996);
and U1110 (N_1110,N_832,N_331);
and U1111 (N_1111,N_91,In_458);
nor U1112 (N_1112,In_2211,N_608);
or U1113 (N_1113,N_889,N_570);
or U1114 (N_1114,In_1813,N_779);
or U1115 (N_1115,In_892,In_1701);
nor U1116 (N_1116,In_1721,In_2388);
nand U1117 (N_1117,In_11,In_1);
nand U1118 (N_1118,In_2486,N_995);
nor U1119 (N_1119,In_2045,N_800);
or U1120 (N_1120,In_811,N_764);
nand U1121 (N_1121,In_1845,In_579);
or U1122 (N_1122,In_473,N_865);
and U1123 (N_1123,N_738,In_2316);
and U1124 (N_1124,In_1795,N_688);
nand U1125 (N_1125,In_2333,N_317);
and U1126 (N_1126,N_137,N_692);
nor U1127 (N_1127,In_988,In_1011);
and U1128 (N_1128,N_372,N_258);
nor U1129 (N_1129,In_1870,In_1095);
nand U1130 (N_1130,In_1520,In_1863);
nand U1131 (N_1131,In_2151,In_1430);
and U1132 (N_1132,In_2459,N_152);
and U1133 (N_1133,In_2384,In_1661);
or U1134 (N_1134,In_1260,N_732);
or U1135 (N_1135,In_54,N_677);
nor U1136 (N_1136,In_1763,N_128);
nand U1137 (N_1137,In_1798,In_2278);
nand U1138 (N_1138,In_1134,In_87);
nor U1139 (N_1139,N_330,N_812);
and U1140 (N_1140,N_993,In_90);
nor U1141 (N_1141,In_2038,In_2030);
and U1142 (N_1142,In_25,In_498);
nor U1143 (N_1143,In_1630,In_2085);
and U1144 (N_1144,N_730,In_2128);
or U1145 (N_1145,In_713,N_760);
nor U1146 (N_1146,N_432,In_2088);
nand U1147 (N_1147,N_13,In_1358);
and U1148 (N_1148,N_752,In_1869);
or U1149 (N_1149,In_1615,In_2155);
or U1150 (N_1150,In_1897,N_887);
or U1151 (N_1151,In_423,N_922);
and U1152 (N_1152,N_104,N_114);
nor U1153 (N_1153,In_575,In_765);
or U1154 (N_1154,In_1698,In_1254);
or U1155 (N_1155,In_1083,In_213);
nand U1156 (N_1156,In_1774,N_130);
xor U1157 (N_1157,N_495,In_2196);
or U1158 (N_1158,In_851,N_808);
and U1159 (N_1159,N_905,In_1725);
or U1160 (N_1160,N_858,In_1256);
or U1161 (N_1161,N_443,N_914);
nand U1162 (N_1162,In_1486,N_631);
or U1163 (N_1163,In_2090,N_136);
nand U1164 (N_1164,N_753,In_1812);
or U1165 (N_1165,In_2241,N_499);
and U1166 (N_1166,In_457,In_1977);
or U1167 (N_1167,In_2214,In_29);
or U1168 (N_1168,N_351,In_803);
or U1169 (N_1169,N_237,In_1241);
nor U1170 (N_1170,N_251,N_392);
nand U1171 (N_1171,In_1478,In_1722);
nand U1172 (N_1172,N_787,In_2266);
and U1173 (N_1173,N_295,In_164);
or U1174 (N_1174,In_2033,In_2268);
nand U1175 (N_1175,N_685,In_2357);
nand U1176 (N_1176,In_1124,In_678);
nand U1177 (N_1177,N_860,In_1487);
nor U1178 (N_1178,In_244,N_390);
and U1179 (N_1179,In_315,In_381);
nor U1180 (N_1180,In_832,In_371);
or U1181 (N_1181,In_906,N_774);
or U1182 (N_1182,In_1703,In_356);
and U1183 (N_1183,In_632,N_131);
or U1184 (N_1184,N_44,N_861);
nor U1185 (N_1185,In_667,N_602);
nor U1186 (N_1186,In_1281,N_422);
and U1187 (N_1187,In_717,In_1712);
nor U1188 (N_1188,In_2042,N_718);
and U1189 (N_1189,N_58,N_149);
and U1190 (N_1190,In_1508,In_1394);
nand U1191 (N_1191,In_688,In_783);
or U1192 (N_1192,N_209,N_228);
and U1193 (N_1193,In_1952,In_1573);
and U1194 (N_1194,In_619,N_624);
and U1195 (N_1195,In_1604,N_989);
nor U1196 (N_1196,In_784,In_447);
nor U1197 (N_1197,N_92,N_405);
nor U1198 (N_1198,In_1702,N_815);
nor U1199 (N_1199,N_763,In_2143);
or U1200 (N_1200,N_641,In_1580);
nor U1201 (N_1201,In_1906,N_590);
and U1202 (N_1202,In_953,N_937);
or U1203 (N_1203,In_743,In_1965);
nor U1204 (N_1204,N_749,In_1770);
nor U1205 (N_1205,In_1875,N_220);
nand U1206 (N_1206,In_2481,N_984);
nand U1207 (N_1207,N_775,N_352);
nor U1208 (N_1208,In_2436,N_491);
xnor U1209 (N_1209,In_2087,In_617);
nand U1210 (N_1210,N_175,In_1332);
and U1211 (N_1211,In_2129,N_838);
and U1212 (N_1212,In_1369,N_371);
or U1213 (N_1213,N_875,In_1302);
and U1214 (N_1214,N_754,N_991);
and U1215 (N_1215,In_435,In_1328);
or U1216 (N_1216,N_189,In_1025);
nor U1217 (N_1217,In_929,In_1553);
or U1218 (N_1218,In_620,In_527);
nand U1219 (N_1219,In_1900,N_964);
or U1220 (N_1220,In_1602,In_521);
and U1221 (N_1221,In_580,N_780);
or U1222 (N_1222,N_999,In_907);
or U1223 (N_1223,N_425,In_2194);
or U1224 (N_1224,In_535,In_1402);
and U1225 (N_1225,In_978,N_79);
nand U1226 (N_1226,N_936,In_705);
nand U1227 (N_1227,N_918,N_64);
and U1228 (N_1228,In_486,In_1404);
or U1229 (N_1229,In_640,In_467);
or U1230 (N_1230,In_1797,In_1987);
nand U1231 (N_1231,N_303,In_937);
nand U1232 (N_1232,In_1009,In_861);
nand U1233 (N_1233,In_638,In_981);
and U1234 (N_1234,In_763,N_113);
nand U1235 (N_1235,N_177,N_982);
nand U1236 (N_1236,N_143,In_1249);
or U1237 (N_1237,In_1904,N_335);
and U1238 (N_1238,In_855,N_262);
and U1239 (N_1239,In_2465,In_1551);
nor U1240 (N_1240,N_545,N_729);
and U1241 (N_1241,N_297,N_745);
and U1242 (N_1242,N_260,In_2353);
or U1243 (N_1243,In_193,N_83);
and U1244 (N_1244,In_1038,In_346);
nand U1245 (N_1245,In_598,In_1861);
nor U1246 (N_1246,In_2209,N_920);
nand U1247 (N_1247,In_2055,N_740);
or U1248 (N_1248,In_429,In_2144);
nand U1249 (N_1249,In_333,In_591);
and U1250 (N_1250,N_852,In_1482);
and U1251 (N_1251,N_217,N_567);
nor U1252 (N_1252,N_846,N_382);
and U1253 (N_1253,N_1116,In_1191);
nand U1254 (N_1254,N_18,N_1148);
nor U1255 (N_1255,N_959,In_2228);
and U1256 (N_1256,N_1064,N_542);
nand U1257 (N_1257,N_1082,N_921);
or U1258 (N_1258,N_1226,N_856);
nor U1259 (N_1259,In_132,N_867);
or U1260 (N_1260,In_1622,In_1078);
and U1261 (N_1261,In_80,In_1388);
nor U1262 (N_1262,In_1425,In_1457);
nand U1263 (N_1263,N_706,N_628);
nand U1264 (N_1264,N_1156,N_980);
nor U1265 (N_1265,N_762,In_840);
or U1266 (N_1266,N_1198,N_69);
and U1267 (N_1267,In_336,N_1246);
nand U1268 (N_1268,In_432,N_477);
or U1269 (N_1269,N_1038,N_1023);
nor U1270 (N_1270,N_973,N_1075);
nor U1271 (N_1271,In_869,N_1129);
or U1272 (N_1272,In_116,N_440);
and U1273 (N_1273,In_1911,N_1016);
nor U1274 (N_1274,In_1571,N_310);
nor U1275 (N_1275,N_802,In_830);
nor U1276 (N_1276,In_663,N_271);
and U1277 (N_1277,N_576,In_2410);
nand U1278 (N_1278,In_318,N_596);
nor U1279 (N_1279,In_1727,N_282);
and U1280 (N_1280,In_1881,N_862);
nor U1281 (N_1281,N_470,N_929);
nand U1282 (N_1282,N_1192,In_2334);
nand U1283 (N_1283,In_1399,N_737);
or U1284 (N_1284,N_47,N_1098);
nand U1285 (N_1285,N_908,N_904);
nor U1286 (N_1286,N_777,In_595);
or U1287 (N_1287,In_2263,N_789);
and U1288 (N_1288,N_373,In_2094);
and U1289 (N_1289,N_406,N_916);
and U1290 (N_1290,N_1242,N_1111);
nand U1291 (N_1291,N_386,In_2076);
or U1292 (N_1292,In_1052,In_105);
nor U1293 (N_1293,N_670,N_806);
nor U1294 (N_1294,N_939,N_897);
nand U1295 (N_1295,N_536,N_776);
and U1296 (N_1296,In_2100,N_932);
or U1297 (N_1297,N_449,N_264);
nand U1298 (N_1298,N_1110,N_154);
or U1299 (N_1299,In_2190,In_1398);
nor U1300 (N_1300,N_118,In_1605);
nor U1301 (N_1301,N_1041,N_1128);
or U1302 (N_1302,N_934,In_1413);
nand U1303 (N_1303,N_557,N_529);
nor U1304 (N_1304,In_296,In_1566);
and U1305 (N_1305,N_1208,In_1403);
nor U1306 (N_1306,In_970,In_1314);
and U1307 (N_1307,N_550,N_755);
nand U1308 (N_1308,N_571,N_1207);
nor U1309 (N_1309,N_1095,N_751);
nand U1310 (N_1310,N_986,N_383);
or U1311 (N_1311,N_208,N_911);
nor U1312 (N_1312,N_970,N_900);
nand U1313 (N_1313,N_535,N_1157);
and U1314 (N_1314,In_1751,N_1078);
and U1315 (N_1315,N_673,In_6);
nand U1316 (N_1316,In_299,N_416);
or U1317 (N_1317,In_1675,In_2290);
and U1318 (N_1318,N_1189,In_945);
nor U1319 (N_1319,N_1183,In_19);
and U1320 (N_1320,N_1169,In_596);
and U1321 (N_1321,In_497,In_1556);
and U1322 (N_1322,N_1074,N_857);
or U1323 (N_1323,In_66,N_1043);
nor U1324 (N_1324,In_570,In_96);
nand U1325 (N_1325,N_736,N_985);
nor U1326 (N_1326,In_1019,In_1951);
nor U1327 (N_1327,In_2072,N_307);
or U1328 (N_1328,In_1377,In_2332);
nand U1329 (N_1329,In_1427,In_2457);
nand U1330 (N_1330,In_2311,N_1240);
nor U1331 (N_1331,N_188,N_355);
nor U1332 (N_1332,In_2373,N_563);
or U1333 (N_1333,N_849,In_2208);
nand U1334 (N_1334,N_845,N_1049);
nor U1335 (N_1335,N_283,In_794);
nand U1336 (N_1336,In_332,N_334);
and U1337 (N_1337,In_2096,In_1144);
nor U1338 (N_1338,N_39,N_811);
nor U1339 (N_1339,In_1033,In_1799);
or U1340 (N_1340,N_1141,In_1603);
nand U1341 (N_1341,N_645,In_1206);
nand U1342 (N_1342,In_759,In_259);
and U1343 (N_1343,In_1352,N_1184);
nand U1344 (N_1344,N_1160,N_1040);
nand U1345 (N_1345,In_397,N_346);
nand U1346 (N_1346,N_783,In_91);
or U1347 (N_1347,In_890,In_600);
and U1348 (N_1348,N_1044,N_1006);
and U1349 (N_1349,N_558,In_2455);
nand U1350 (N_1350,N_1124,N_117);
nor U1351 (N_1351,N_514,In_740);
and U1352 (N_1352,In_976,In_1008);
or U1353 (N_1353,In_1451,In_966);
and U1354 (N_1354,In_2066,N_834);
or U1355 (N_1355,N_462,N_583);
nor U1356 (N_1356,N_304,In_1671);
nand U1357 (N_1357,N_797,In_2391);
and U1358 (N_1358,N_652,N_16);
nand U1359 (N_1359,In_1985,In_1506);
nand U1360 (N_1360,In_1165,N_486);
nor U1361 (N_1361,N_1212,N_325);
or U1362 (N_1362,N_1033,N_717);
or U1363 (N_1363,In_968,N_559);
or U1364 (N_1364,In_187,N_35);
and U1365 (N_1365,N_162,N_1176);
nor U1366 (N_1366,N_438,N_1232);
and U1367 (N_1367,In_2031,N_910);
and U1368 (N_1368,N_1138,N_796);
nor U1369 (N_1369,N_1134,N_494);
and U1370 (N_1370,N_591,In_1764);
nand U1371 (N_1371,N_132,In_2062);
nor U1372 (N_1372,In_751,In_399);
and U1373 (N_1373,N_1051,In_1060);
nand U1374 (N_1374,N_1060,In_524);
and U1375 (N_1375,N_1143,In_1838);
and U1376 (N_1376,N_977,N_1161);
or U1377 (N_1377,In_1341,N_1146);
or U1378 (N_1378,In_2122,In_534);
and U1379 (N_1379,In_1239,In_363);
nand U1380 (N_1380,N_951,In_902);
and U1381 (N_1381,In_1349,N_968);
and U1382 (N_1382,In_2160,N_1108);
and U1383 (N_1383,In_1346,N_870);
or U1384 (N_1384,N_671,N_507);
and U1385 (N_1385,In_707,In_744);
nand U1386 (N_1386,In_4,In_1973);
nor U1387 (N_1387,In_999,In_959);
or U1388 (N_1388,In_792,In_228);
or U1389 (N_1389,In_1220,In_284);
and U1390 (N_1390,N_843,In_30);
nand U1391 (N_1391,N_275,N_1114);
nand U1392 (N_1392,In_810,N_1021);
or U1393 (N_1393,N_192,In_918);
or U1394 (N_1394,In_567,In_1585);
or U1395 (N_1395,N_719,N_1015);
nand U1396 (N_1396,N_510,N_975);
nor U1397 (N_1397,N_480,In_1271);
and U1398 (N_1398,N_756,In_2326);
and U1399 (N_1399,N_1001,N_1027);
nand U1400 (N_1400,In_775,In_1694);
and U1401 (N_1401,In_1590,In_1360);
or U1402 (N_1402,In_2002,N_1080);
nand U1403 (N_1403,In_2181,N_1017);
and U1404 (N_1404,In_455,In_860);
or U1405 (N_1405,In_998,N_164);
and U1406 (N_1406,N_25,N_621);
nand U1407 (N_1407,N_743,N_1022);
and U1408 (N_1408,In_1415,N_1199);
nand U1409 (N_1409,N_961,N_1224);
nor U1410 (N_1410,N_290,In_2197);
nand U1411 (N_1411,N_1190,N_704);
nor U1412 (N_1412,N_637,In_2239);
and U1413 (N_1413,N_724,In_1747);
nand U1414 (N_1414,In_2277,N_599);
nand U1415 (N_1415,In_283,N_1222);
nand U1416 (N_1416,In_2186,In_350);
nor U1417 (N_1417,N_1197,N_644);
nor U1418 (N_1418,N_1019,In_1146);
nand U1419 (N_1419,In_995,N_1166);
and U1420 (N_1420,N_1237,N_1053);
nor U1421 (N_1421,N_460,In_921);
nand U1422 (N_1422,N_1058,N_1096);
xnor U1423 (N_1423,In_813,In_2296);
nand U1424 (N_1424,N_1070,In_2009);
and U1425 (N_1425,N_544,In_1357);
or U1426 (N_1426,In_2361,In_1013);
nor U1427 (N_1427,N_907,In_2343);
or U1428 (N_1428,N_1032,N_1187);
or U1429 (N_1429,N_1211,In_55);
nor U1430 (N_1430,N_1042,In_270);
and U1431 (N_1431,N_343,In_433);
and U1432 (N_1432,In_1492,In_271);
or U1433 (N_1433,N_859,In_1998);
and U1434 (N_1434,In_258,N_925);
or U1435 (N_1435,N_1135,In_2250);
and U1436 (N_1436,In_2234,N_1241);
and U1437 (N_1437,N_141,N_1085);
or U1438 (N_1438,N_100,N_884);
nor U1439 (N_1439,N_1028,N_475);
and U1440 (N_1440,In_59,N_1079);
nor U1441 (N_1441,In_971,N_667);
and U1442 (N_1442,N_179,In_71);
nor U1443 (N_1443,N_863,N_1093);
or U1444 (N_1444,N_643,In_1333);
nand U1445 (N_1445,N_531,N_1091);
nor U1446 (N_1446,N_839,N_1045);
and U1447 (N_1447,N_931,In_2383);
or U1448 (N_1448,In_1515,N_1238);
nand U1449 (N_1449,N_825,N_376);
nor U1450 (N_1450,N_30,N_1063);
or U1451 (N_1451,N_909,N_465);
and U1452 (N_1452,N_59,In_226);
nand U1453 (N_1453,In_530,In_616);
and U1454 (N_1454,N_261,N_888);
or U1455 (N_1455,In_321,N_879);
nand U1456 (N_1456,In_1336,N_1062);
and U1457 (N_1457,In_2282,In_94);
and U1458 (N_1458,In_542,In_1501);
nand U1459 (N_1459,In_2000,N_733);
nor U1460 (N_1460,N_892,In_1620);
nor U1461 (N_1461,In_836,N_328);
nor U1462 (N_1462,N_633,In_773);
nand U1463 (N_1463,In_2406,N_457);
or U1464 (N_1464,N_1054,In_1783);
nand U1465 (N_1465,In_278,In_1085);
nor U1466 (N_1466,In_2495,In_672);
nor U1467 (N_1467,In_1122,N_96);
or U1468 (N_1468,In_1286,In_1108);
nand U1469 (N_1469,N_772,N_1235);
nand U1470 (N_1470,N_622,N_65);
nor U1471 (N_1471,N_1159,In_1417);
and U1472 (N_1472,N_886,N_337);
and U1473 (N_1473,In_1000,N_842);
and U1474 (N_1474,In_1065,In_1296);
or U1475 (N_1475,In_1463,In_403);
and U1476 (N_1476,In_1385,N_513);
nor U1477 (N_1477,N_1057,N_1223);
or U1478 (N_1478,N_1002,N_109);
or U1479 (N_1479,In_1628,In_1472);
nand U1480 (N_1480,In_347,N_1228);
or U1481 (N_1481,In_2225,In_1983);
or U1482 (N_1482,In_838,In_289);
or U1483 (N_1483,In_1002,N_949);
or U1484 (N_1484,N_869,N_912);
or U1485 (N_1485,In_624,In_343);
nor U1486 (N_1486,N_952,In_438);
or U1487 (N_1487,In_389,In_1464);
nand U1488 (N_1488,In_2093,N_1059);
and U1489 (N_1489,In_2339,N_965);
nand U1490 (N_1490,In_2398,In_1461);
nor U1491 (N_1491,In_1704,N_72);
nor U1492 (N_1492,In_2450,In_101);
nor U1493 (N_1493,In_2195,In_955);
nand U1494 (N_1494,N_960,N_695);
and U1495 (N_1495,N_549,In_761);
and U1496 (N_1496,N_1034,In_126);
and U1497 (N_1497,N_1196,N_60);
nand U1498 (N_1498,In_1696,In_2204);
and U1499 (N_1499,In_2184,N_930);
nor U1500 (N_1500,N_1445,In_2371);
nand U1501 (N_1501,N_363,N_1039);
nor U1502 (N_1502,N_614,In_1322);
and U1503 (N_1503,N_1055,N_1398);
nand U1504 (N_1504,N_1067,N_586);
nand U1505 (N_1505,In_1853,In_931);
nor U1506 (N_1506,N_1408,N_582);
and U1507 (N_1507,In_2496,N_1460);
nand U1508 (N_1508,N_595,In_612);
or U1509 (N_1509,N_273,N_568);
and U1510 (N_1510,N_1417,N_433);
or U1511 (N_1511,N_1455,In_2267);
or U1512 (N_1512,N_1407,N_761);
nor U1513 (N_1513,In_2440,N_1331);
nor U1514 (N_1514,N_1492,N_1340);
or U1515 (N_1515,In_453,In_50);
and U1516 (N_1516,In_142,N_1274);
nand U1517 (N_1517,N_1444,In_1176);
and U1518 (N_1518,N_1188,N_1102);
nor U1519 (N_1519,N_501,N_1324);
nor U1520 (N_1520,In_494,N_1463);
nor U1521 (N_1521,In_370,N_1465);
and U1522 (N_1522,In_421,In_958);
and U1523 (N_1523,In_396,N_758);
and U1524 (N_1524,In_324,In_1485);
or U1525 (N_1525,N_1084,In_518);
and U1526 (N_1526,In_1223,N_654);
or U1527 (N_1527,In_1490,In_1301);
and U1528 (N_1528,N_1278,In_587);
nand U1529 (N_1529,N_436,N_634);
or U1530 (N_1530,N_893,N_684);
nor U1531 (N_1531,N_579,N_1037);
or U1532 (N_1532,N_1436,In_2396);
nor U1533 (N_1533,N_1269,N_1125);
nor U1534 (N_1534,In_46,N_459);
or U1535 (N_1535,N_361,N_1185);
and U1536 (N_1536,N_1103,In_1129);
and U1537 (N_1537,In_102,In_1507);
or U1538 (N_1538,N_1419,In_1513);
nor U1539 (N_1539,N_1259,N_794);
and U1540 (N_1540,In_2092,N_769);
nand U1541 (N_1541,In_1433,N_1003);
and U1542 (N_1542,N_1122,In_261);
nand U1543 (N_1543,In_65,N_281);
nand U1544 (N_1544,N_1451,N_679);
and U1545 (N_1545,N_393,N_948);
nand U1546 (N_1546,N_1256,In_2132);
and U1547 (N_1547,N_1420,In_1944);
or U1548 (N_1548,N_1025,N_244);
nand U1549 (N_1549,N_618,N_1231);
nor U1550 (N_1550,In_451,N_798);
nor U1551 (N_1551,In_1135,In_418);
nand U1552 (N_1552,N_1065,In_1974);
and U1553 (N_1553,In_1289,N_167);
or U1554 (N_1554,N_1258,N_1290);
nor U1555 (N_1555,N_1221,In_2483);
nand U1556 (N_1556,N_1266,In_1163);
nand U1557 (N_1557,N_1163,N_1477);
nand U1558 (N_1558,In_1028,N_1428);
nor U1559 (N_1559,N_541,In_2298);
xor U1560 (N_1560,N_791,In_2307);
and U1561 (N_1561,In_476,N_1081);
nor U1562 (N_1562,N_1356,N_1381);
nand U1563 (N_1563,N_768,In_1731);
nor U1564 (N_1564,In_933,N_1421);
nor U1565 (N_1565,N_766,N_1047);
nand U1566 (N_1566,N_824,N_1151);
or U1567 (N_1567,N_1391,N_1302);
or U1568 (N_1568,N_492,N_1387);
xor U1569 (N_1569,In_1123,In_107);
and U1570 (N_1570,N_356,N_551);
nor U1571 (N_1571,N_1397,N_1487);
nor U1572 (N_1572,N_1338,N_1355);
or U1573 (N_1573,N_1469,In_1471);
and U1574 (N_1574,N_28,In_201);
and U1575 (N_1575,N_366,In_2356);
or U1576 (N_1576,N_12,N_1195);
and U1577 (N_1577,N_1352,N_1326);
and U1578 (N_1578,N_163,In_647);
and U1579 (N_1579,N_1008,In_824);
or U1580 (N_1580,N_1403,N_1362);
and U1581 (N_1581,In_1015,N_1339);
or U1582 (N_1582,In_1055,In_52);
or U1583 (N_1583,In_2049,In_889);
and U1584 (N_1584,N_994,N_1225);
nand U1585 (N_1585,In_2006,N_1412);
and U1586 (N_1586,In_1419,N_1384);
or U1587 (N_1587,N_604,N_369);
or U1588 (N_1588,N_1099,N_750);
nor U1589 (N_1589,N_1337,N_553);
and U1590 (N_1590,N_1165,N_1485);
and U1591 (N_1591,In_1517,N_1264);
or U1592 (N_1592,In_990,N_288);
and U1593 (N_1593,N_1069,N_899);
and U1594 (N_1594,N_837,In_689);
nor U1595 (N_1595,N_901,N_322);
nor U1596 (N_1596,N_1435,N_945);
nor U1597 (N_1597,N_1254,In_67);
or U1598 (N_1598,N_1341,N_1430);
nor U1599 (N_1599,N_1117,N_1279);
nand U1600 (N_1600,In_2426,N_696);
and U1601 (N_1601,N_1348,N_1210);
nor U1602 (N_1602,N_1167,N_997);
nand U1603 (N_1603,In_1857,N_782);
xor U1604 (N_1604,In_1087,N_1181);
or U1605 (N_1605,N_1136,In_162);
and U1606 (N_1606,N_1346,N_826);
nor U1607 (N_1607,N_238,In_1423);
nor U1608 (N_1608,N_1380,In_1649);
and U1609 (N_1609,In_1846,In_509);
and U1610 (N_1610,N_340,N_917);
nand U1611 (N_1611,N_505,N_442);
nor U1612 (N_1612,N_243,N_1296);
and U1613 (N_1613,N_734,In_98);
nand U1614 (N_1614,N_976,N_950);
nand U1615 (N_1615,N_419,In_45);
nor U1616 (N_1616,N_721,N_1411);
and U1617 (N_1617,N_1205,N_1194);
or U1618 (N_1618,N_1314,In_1740);
and U1619 (N_1619,N_610,N_1105);
or U1620 (N_1620,N_1305,In_209);
and U1621 (N_1621,N_1478,N_1385);
or U1622 (N_1622,N_786,N_144);
and U1623 (N_1623,In_256,N_962);
nor U1624 (N_1624,In_1216,In_1830);
and U1625 (N_1625,N_1107,In_1081);
nand U1626 (N_1626,In_726,In_725);
or U1627 (N_1627,In_2315,N_1229);
nor U1628 (N_1628,N_1130,N_1206);
or U1629 (N_1629,N_850,In_2041);
nand U1630 (N_1630,N_1179,N_287);
or U1631 (N_1631,N_1209,N_518);
and U1632 (N_1632,In_645,N_1343);
or U1633 (N_1633,In_1495,N_1323);
and U1634 (N_1634,N_1393,In_1984);
nor U1635 (N_1635,N_1395,N_587);
nor U1636 (N_1636,N_1328,N_788);
or U1637 (N_1637,In_2477,N_795);
and U1638 (N_1638,N_1126,N_996);
nor U1639 (N_1639,N_821,N_1173);
nand U1640 (N_1640,In_93,N_1292);
nor U1641 (N_1641,In_1198,In_897);
and U1642 (N_1642,N_1404,N_585);
and U1643 (N_1643,N_1068,N_1248);
nand U1644 (N_1644,In_1153,N_1413);
and U1645 (N_1645,N_1350,In_366);
or U1646 (N_1646,In_2067,In_1745);
or U1647 (N_1647,N_759,N_1233);
or U1648 (N_1648,N_1140,N_1443);
or U1649 (N_1649,In_2231,N_833);
nand U1650 (N_1650,In_1927,N_1282);
or U1651 (N_1651,N_974,N_1088);
or U1652 (N_1652,N_714,In_493);
nand U1653 (N_1653,N_1371,N_1402);
or U1654 (N_1654,N_1330,In_593);
or U1655 (N_1655,In_741,In_195);
nor U1656 (N_1656,N_979,In_41);
or U1657 (N_1657,N_946,N_895);
nand U1658 (N_1658,In_121,In_866);
nand U1659 (N_1659,N_1171,N_1471);
nor U1660 (N_1660,N_1164,N_1466);
and U1661 (N_1661,N_1461,N_1334);
or U1662 (N_1662,N_765,N_971);
and U1663 (N_1663,N_424,N_1452);
or U1664 (N_1664,N_1448,N_1459);
nand U1665 (N_1665,N_801,N_873);
and U1666 (N_1666,In_1382,N_890);
nand U1667 (N_1667,N_804,N_771);
nor U1668 (N_1668,N_661,In_1354);
nand U1669 (N_1669,N_1046,N_447);
nor U1670 (N_1670,N_793,N_1429);
or U1671 (N_1671,In_659,N_1473);
or U1672 (N_1672,N_1300,N_115);
nand U1673 (N_1673,N_1158,In_1773);
or U1674 (N_1674,In_2341,In_1311);
nand U1675 (N_1675,In_1516,N_1342);
nor U1676 (N_1676,In_1137,N_357);
nand U1677 (N_1677,In_525,N_1215);
and U1678 (N_1678,N_1378,N_1457);
or U1679 (N_1679,N_742,In_787);
and U1680 (N_1680,In_1522,N_1200);
or U1681 (N_1681,N_1193,In_507);
nand U1682 (N_1682,N_504,In_1677);
and U1683 (N_1683,N_581,N_1145);
nand U1684 (N_1684,N_1447,N_1453);
nor U1685 (N_1685,N_302,N_1100);
or U1686 (N_1686,In_724,In_1003);
nand U1687 (N_1687,In_1029,N_881);
nor U1688 (N_1688,N_1312,N_1276);
nor U1689 (N_1689,N_1310,In_1837);
and U1690 (N_1690,N_1496,N_1147);
nor U1691 (N_1691,N_1012,In_1530);
nor U1692 (N_1692,N_853,In_908);
nor U1693 (N_1693,N_573,In_233);
nand U1694 (N_1694,N_817,N_540);
nand U1695 (N_1695,N_1319,N_1261);
nor U1696 (N_1696,In_251,N_1144);
or U1697 (N_1697,N_1036,N_1061);
nand U1698 (N_1698,N_474,In_2468);
nor U1699 (N_1699,N_639,In_1016);
nand U1700 (N_1700,N_1214,In_1978);
nand U1701 (N_1701,In_280,N_1441);
and U1702 (N_1702,N_1336,N_1050);
nand U1703 (N_1703,N_1345,N_687);
and U1704 (N_1704,In_1683,N_1382);
and U1705 (N_1705,In_757,N_792);
or U1706 (N_1706,N_1251,N_627);
and U1707 (N_1707,N_399,N_1243);
and U1708 (N_1708,N_75,N_682);
nor U1709 (N_1709,N_1244,N_1383);
or U1710 (N_1710,N_1472,In_649);
or U1711 (N_1711,In_1240,N_877);
nand U1712 (N_1712,N_387,N_324);
or U1713 (N_1713,In_1758,N_1366);
xnor U1714 (N_1714,N_1396,N_1335);
or U1715 (N_1715,In_2233,N_1142);
nand U1716 (N_1716,In_2283,N_1217);
or U1717 (N_1717,In_1644,In_1916);
and U1718 (N_1718,N_1123,In_1535);
and U1719 (N_1719,In_1739,N_548);
nand U1720 (N_1720,N_987,N_944);
or U1721 (N_1721,In_1057,N_1365);
nor U1722 (N_1722,N_1361,N_1320);
nand U1723 (N_1723,N_1120,In_2035);
nor U1724 (N_1724,N_1283,In_1024);
nand U1725 (N_1725,In_1650,In_2219);
and U1726 (N_1726,N_1066,N_222);
and U1727 (N_1727,N_603,N_1288);
and U1728 (N_1728,In_42,N_919);
nand U1729 (N_1729,In_1756,In_427);
and U1730 (N_1730,N_0,In_1755);
nor U1731 (N_1731,N_1307,N_526);
and U1732 (N_1732,N_1218,N_493);
or U1733 (N_1733,N_467,N_1092);
nand U1734 (N_1734,In_441,In_2390);
nor U1735 (N_1735,In_847,N_1056);
nand U1736 (N_1736,N_906,N_1267);
nand U1737 (N_1737,In_780,N_1048);
nand U1738 (N_1738,N_933,N_597);
nor U1739 (N_1739,N_880,In_1679);
nor U1740 (N_1740,N_1168,N_972);
nand U1741 (N_1741,N_819,In_2363);
nand U1742 (N_1742,In_767,In_615);
nand U1743 (N_1743,In_1621,N_1358);
or U1744 (N_1744,N_49,N_830);
and U1745 (N_1745,N_1468,N_1354);
nor U1746 (N_1746,N_689,In_1682);
and U1747 (N_1747,In_2091,N_1014);
nand U1748 (N_1748,N_1394,In_1926);
and U1749 (N_1749,In_854,N_1497);
nor U1750 (N_1750,N_1253,In_2366);
and U1751 (N_1751,N_1601,In_623);
xnor U1752 (N_1752,N_1665,In_1761);
and U1753 (N_1753,N_1191,N_201);
xnor U1754 (N_1754,N_1568,In_764);
or U1755 (N_1755,N_1203,N_1550);
and U1756 (N_1756,In_262,N_1632);
nor U1757 (N_1757,In_173,In_1593);
nand U1758 (N_1758,N_489,N_1293);
nor U1759 (N_1759,N_1585,In_1067);
nand U1760 (N_1760,N_1657,In_771);
or U1761 (N_1761,N_1559,N_1423);
or U1762 (N_1762,N_1359,N_1536);
and U1763 (N_1763,N_1257,N_1427);
and U1764 (N_1764,In_1203,N_1297);
nand U1765 (N_1765,N_1476,N_1462);
nand U1766 (N_1766,N_253,In_1012);
nand U1767 (N_1767,N_629,In_1543);
or U1768 (N_1768,N_1369,N_78);
nand U1769 (N_1769,N_1635,N_1586);
and U1770 (N_1770,In_303,N_928);
and U1771 (N_1771,N_1714,N_1608);
and U1772 (N_1772,N_1589,In_801);
and U1773 (N_1773,In_1218,N_1152);
or U1774 (N_1774,N_1557,N_1721);
nor U1775 (N_1775,N_284,In_361);
and U1776 (N_1776,N_990,N_840);
nor U1777 (N_1777,N_1628,N_1177);
or U1778 (N_1778,N_848,N_517);
or U1779 (N_1779,In_844,N_1534);
nor U1780 (N_1780,N_308,N_1375);
nor U1781 (N_1781,N_51,N_345);
and U1782 (N_1782,N_636,N_1491);
nand U1783 (N_1783,N_546,N_1071);
nand U1784 (N_1784,N_1437,N_1464);
or U1785 (N_1785,N_116,In_2447);
and U1786 (N_1786,N_1520,N_522);
or U1787 (N_1787,N_941,N_1101);
or U1788 (N_1788,N_1706,N_1584);
or U1789 (N_1789,N_1683,N_1654);
nand U1790 (N_1790,N_1119,N_56);
nor U1791 (N_1791,N_1400,N_1688);
and U1792 (N_1792,N_1741,N_947);
nor U1793 (N_1793,In_943,N_1554);
and U1794 (N_1794,N_1377,N_1623);
or U1795 (N_1795,In_357,In_77);
and U1796 (N_1796,N_1668,N_1510);
or U1797 (N_1797,In_979,In_739);
nor U1798 (N_1798,N_1127,In_749);
nand U1799 (N_1799,N_584,N_1650);
and U1800 (N_1800,N_1658,N_1137);
and U1801 (N_1801,N_8,N_1684);
xnor U1802 (N_1802,N_814,N_1370);
and U1803 (N_1803,In_1034,N_381);
and U1804 (N_1804,N_1679,N_1272);
or U1805 (N_1805,N_1527,N_1609);
and U1806 (N_1806,N_1097,N_659);
or U1807 (N_1807,N_1406,N_1720);
and U1808 (N_1808,N_710,N_1541);
and U1809 (N_1809,N_1013,In_965);
nand U1810 (N_1810,N_1599,N_847);
and U1811 (N_1811,N_1175,N_1303);
and U1812 (N_1812,In_231,N_1701);
and U1813 (N_1813,N_1739,N_1113);
or U1814 (N_1814,N_978,N_1667);
or U1815 (N_1815,N_1285,N_1693);
nor U1816 (N_1816,N_1484,N_145);
nand U1817 (N_1817,N_1549,In_1705);
and U1818 (N_1818,In_831,N_1664);
nand U1819 (N_1819,N_1422,N_1115);
nor U1820 (N_1820,N_953,N_1357);
or U1821 (N_1821,N_1268,N_1470);
or U1822 (N_1822,N_1317,N_1155);
and U1823 (N_1823,N_574,N_1640);
nand U1824 (N_1824,N_1029,N_1593);
or U1825 (N_1825,In_204,N_1732);
and U1826 (N_1826,N_1503,N_1704);
and U1827 (N_1827,N_1132,N_1271);
or U1828 (N_1828,N_1482,N_868);
and U1829 (N_1829,N_1728,In_1658);
or U1830 (N_1830,In_2052,In_139);
nand U1831 (N_1831,N_1219,N_1716);
nor U1832 (N_1832,N_1565,N_107);
and U1833 (N_1833,N_1695,In_829);
and U1834 (N_1834,N_1431,In_2001);
nor U1835 (N_1835,In_1422,N_1440);
nor U1836 (N_1836,In_1326,In_1022);
and U1837 (N_1837,N_1349,N_1133);
nor U1838 (N_1838,N_1446,N_1629);
nand U1839 (N_1839,In_1434,N_1474);
nor U1840 (N_1840,In_60,N_829);
nand U1841 (N_1841,In_1149,N_1551);
nor U1842 (N_1842,N_827,N_413);
nand U1843 (N_1843,In_1681,N_63);
and U1844 (N_1844,N_1479,N_1649);
and U1845 (N_1845,N_556,In_1414);
nand U1846 (N_1846,N_1090,N_1647);
nand U1847 (N_1847,N_1547,N_1634);
and U1848 (N_1848,N_653,N_669);
and U1849 (N_1849,N_1094,In_359);
and U1850 (N_1850,N_289,N_1501);
nor U1851 (N_1851,N_1611,N_1504);
and U1852 (N_1852,N_1700,N_1072);
or U1853 (N_1853,N_725,N_1594);
nor U1854 (N_1854,N_375,N_1562);
and U1855 (N_1855,N_1518,In_709);
and U1856 (N_1856,N_1576,N_1363);
nor U1857 (N_1857,N_1230,N_1630);
nand U1858 (N_1858,N_1104,N_1327);
or U1859 (N_1859,N_799,N_1368);
nand U1860 (N_1860,N_218,In_2188);
or U1861 (N_1861,N_1322,N_1291);
nor U1862 (N_1862,N_1710,N_746);
xnor U1863 (N_1863,N_1636,N_1392);
and U1864 (N_1864,N_125,N_1727);
nor U1865 (N_1865,N_1170,N_414);
or U1866 (N_1866,N_1519,N_1450);
nor U1867 (N_1867,N_1588,N_1597);
nor U1868 (N_1868,N_1390,N_1590);
or U1869 (N_1869,N_726,In_559);
or U1870 (N_1870,N_1626,In_2489);
nand U1871 (N_1871,N_1724,N_1743);
and U1872 (N_1872,N_1360,In_26);
or U1873 (N_1873,N_1410,N_347);
nand U1874 (N_1874,N_1619,N_327);
nand U1875 (N_1875,N_809,N_1605);
nand U1876 (N_1876,N_1737,N_1204);
nor U1877 (N_1877,N_278,N_552);
or U1878 (N_1878,N_255,N_1733);
nor U1879 (N_1879,N_855,N_790);
or U1880 (N_1880,N_1571,In_1136);
nand U1881 (N_1881,N_1415,In_110);
or U1882 (N_1882,N_45,N_1153);
and U1883 (N_1883,N_1575,In_118);
nand U1884 (N_1884,N_1592,In_1128);
and U1885 (N_1885,In_95,N_1494);
or U1886 (N_1886,N_1486,N_198);
and U1887 (N_1887,N_1625,N_1662);
and U1888 (N_1888,N_924,N_1388);
nor U1889 (N_1889,N_1682,N_1690);
nor U1890 (N_1890,N_1596,N_1475);
and U1891 (N_1891,N_1174,N_1073);
or U1892 (N_1892,N_1595,N_1449);
and U1893 (N_1893,In_2016,In_2064);
and U1894 (N_1894,N_956,N_1670);
or U1895 (N_1895,N_1675,N_1182);
and U1896 (N_1896,N_926,N_1216);
nor U1897 (N_1897,N_1432,N_831);
or U1898 (N_1898,N_1304,N_1089);
or U1899 (N_1899,N_1618,In_572);
nand U1900 (N_1900,N_1252,N_233);
or U1901 (N_1901,N_1602,In_144);
nand U1902 (N_1902,N_1511,N_314);
nor U1903 (N_1903,In_2399,N_1607);
nand U1904 (N_1904,N_1301,N_1631);
nor U1905 (N_1905,N_358,In_938);
or U1906 (N_1906,In_546,N_1483);
nor U1907 (N_1907,N_1582,N_1521);
nand U1908 (N_1908,N_1367,In_2279);
nand U1909 (N_1909,N_1121,N_1548);
nand U1910 (N_1910,N_1600,N_1656);
and U1911 (N_1911,N_1009,N_1622);
nor U1912 (N_1912,N_1500,N_1738);
nor U1913 (N_1913,N_1730,In_2051);
nand U1914 (N_1914,N_1633,N_1386);
nand U1915 (N_1915,N_1005,N_1162);
nor U1916 (N_1916,N_1522,In_543);
nand U1917 (N_1917,N_1747,N_1616);
nor U1918 (N_1918,N_1603,N_84);
and U1919 (N_1919,N_1506,In_257);
nand U1920 (N_1920,In_1263,N_784);
or U1921 (N_1921,N_1236,N_1220);
nor U1922 (N_1922,N_1718,N_1680);
nand U1923 (N_1923,N_1641,In_1117);
and U1924 (N_1924,N_1655,N_891);
nor U1925 (N_1925,N_276,N_1424);
nor U1926 (N_1926,N_1507,N_1713);
nor U1927 (N_1927,N_1213,In_554);
nand U1928 (N_1928,In_480,In_2374);
nand U1929 (N_1929,In_1162,N_851);
and U1930 (N_1930,N_1708,N_828);
and U1931 (N_1931,In_23,N_1530);
nand U1932 (N_1932,In_2032,N_818);
or U1933 (N_1933,N_1298,N_234);
or U1934 (N_1934,N_1250,In_876);
and U1935 (N_1935,N_1691,N_1287);
and U1936 (N_1936,N_1109,In_762);
nor U1937 (N_1937,N_1517,N_1531);
nor U1938 (N_1938,N_674,N_1481);
nor U1939 (N_1939,N_1726,N_1493);
and U1940 (N_1940,N_988,N_1260);
nand U1941 (N_1941,In_1785,N_1612);
nand U1942 (N_1942,N_1372,N_1627);
nand U1943 (N_1943,N_1458,In_1448);
nor U1944 (N_1944,N_1643,N_1638);
nand U1945 (N_1945,N_711,N_1673);
nand U1946 (N_1946,N_1513,In_1997);
and U1947 (N_1947,N_1717,N_1729);
or U1948 (N_1948,N_268,N_1544);
and U1949 (N_1949,N_1644,N_396);
nand U1950 (N_1950,N_1529,In_1895);
or U1951 (N_1951,N_1639,N_1454);
nor U1952 (N_1952,N_1566,In_1421);
and U1953 (N_1953,In_184,N_1433);
and U1954 (N_1954,N_471,N_1645);
or U1955 (N_1955,N_1344,In_2010);
and U1956 (N_1956,In_1042,In_44);
nor U1957 (N_1957,In_2288,N_942);
and U1958 (N_1958,N_1745,In_40);
and U1959 (N_1959,N_1694,In_1099);
nor U1960 (N_1960,N_1524,N_940);
or U1961 (N_1961,N_606,N_1698);
nand U1962 (N_1962,N_1004,N_1325);
or U1963 (N_1963,N_1674,N_543);
or U1964 (N_1964,N_1542,In_273);
and U1965 (N_1965,N_1676,In_2123);
and U1966 (N_1966,N_1648,N_1270);
nand U1967 (N_1967,N_1570,N_957);
nor U1968 (N_1968,N_370,In_373);
or U1969 (N_1969,N_1525,N_1748);
nor U1970 (N_1970,N_1262,N_1637);
and U1971 (N_1971,N_1553,N_1373);
nand U1972 (N_1972,N_1376,N_1569);
or U1973 (N_1973,N_699,In_1161);
or U1974 (N_1974,In_2413,N_1031);
nor U1975 (N_1975,N_1703,In_502);
nor U1976 (N_1976,N_1663,In_1250);
and U1977 (N_1977,N_1574,N_1495);
and U1978 (N_1978,In_1931,In_2120);
or U1979 (N_1979,N_1425,In_2029);
nand U1980 (N_1980,N_1545,In_1278);
xnor U1981 (N_1981,N_648,In_1017);
nor U1982 (N_1982,N_1567,N_943);
nor U1983 (N_1983,In_944,N_1523);
and U1984 (N_1984,N_256,N_1659);
nor U1985 (N_1985,N_1587,N_434);
nor U1986 (N_1986,N_1528,In_2358);
nand U1987 (N_1987,N_1315,N_1560);
and U1988 (N_1988,N_1715,N_1249);
or U1989 (N_1989,N_1653,N_1026);
nand U1990 (N_1990,In_1640,N_555);
or U1991 (N_1991,N_1516,In_1036);
or U1992 (N_1992,N_1488,In_1069);
or U1993 (N_1993,N_1052,N_1490);
and U1994 (N_1994,N_1000,N_1539);
nand U1995 (N_1995,In_398,N_1011);
nand U1996 (N_1996,N_1351,N_1512);
nand U1997 (N_1997,N_1178,N_1742);
and U1998 (N_1998,N_1672,N_915);
nand U1999 (N_1999,N_1020,In_2444);
or U2000 (N_2000,N_561,N_181);
and U2001 (N_2001,N_1709,N_142);
nand U2002 (N_2002,N_1572,N_1936);
and U2003 (N_2003,N_1150,N_1854);
nand U2004 (N_2004,N_1912,N_1910);
and U2005 (N_2005,N_1766,N_1943);
or U2006 (N_2006,N_1955,N_1857);
and U2007 (N_2007,N_1877,N_1961);
or U2008 (N_2008,N_1660,N_1131);
or U2009 (N_2009,N_1865,N_1830);
nor U2010 (N_2010,N_1273,N_1735);
or U2011 (N_2011,N_1870,N_1822);
and U2012 (N_2012,N_292,N_1818);
or U2013 (N_2013,N_1306,In_1631);
or U2014 (N_2014,N_1981,N_1467);
nand U2015 (N_2015,In_2294,N_1765);
nor U2016 (N_2016,N_1788,N_1940);
nand U2017 (N_2017,N_1883,N_1893);
nor U2018 (N_2018,N_1753,N_1891);
and U2019 (N_2019,N_864,N_1935);
or U2020 (N_2020,N_1800,N_1843);
nand U2021 (N_2021,N_1118,In_1255);
or U2022 (N_2022,N_1858,N_1389);
and U2023 (N_2023,N_690,N_1824);
or U2024 (N_2024,N_1862,N_1789);
nor U2025 (N_2025,N_1867,N_658);
or U2026 (N_2026,N_1901,N_1831);
or U2027 (N_2027,N_1887,N_1499);
nand U2028 (N_2028,N_1749,N_1884);
or U2029 (N_2029,N_1844,N_1797);
nand U2030 (N_2030,N_1332,In_214);
nand U2031 (N_2031,N_882,N_1968);
nor U2032 (N_2032,N_1234,N_469);
nor U2033 (N_2033,N_1149,N_1848);
or U2034 (N_2034,In_2372,N_1944);
or U2035 (N_2035,In_1878,N_1374);
nand U2036 (N_2036,N_1889,N_1613);
nor U2037 (N_2037,N_1930,N_1686);
nor U2038 (N_2038,N_528,N_1950);
and U2039 (N_2039,N_1767,N_1991);
or U2040 (N_2040,N_1806,N_1677);
nor U2041 (N_2041,In_253,N_1689);
nor U2042 (N_2042,N_1018,N_1722);
xnor U2043 (N_2043,N_1263,N_1010);
and U2044 (N_2044,N_1775,N_1847);
and U2045 (N_2045,N_1882,N_1932);
nor U2046 (N_2046,N_1505,In_1561);
and U2047 (N_2047,N_173,N_1927);
nand U2048 (N_2048,N_1578,N_1786);
and U2049 (N_2049,N_1646,In_1126);
and U2050 (N_2050,N_1439,N_1888);
nand U2051 (N_2051,N_1834,N_1681);
and U2052 (N_2052,N_1313,N_1836);
nand U2053 (N_2053,N_781,N_1974);
and U2054 (N_2054,N_1809,N_1591);
nor U2055 (N_2055,N_1414,N_894);
nor U2056 (N_2056,N_1364,N_1963);
nor U2057 (N_2057,N_1489,N_1416);
nor U2058 (N_2058,N_1418,N_1770);
and U2059 (N_2059,N_1139,N_1255);
or U2060 (N_2060,N_1699,N_1948);
nor U2061 (N_2061,N_1353,N_1172);
nand U2062 (N_2062,N_336,N_1881);
nand U2063 (N_2063,N_1087,N_1798);
or U2064 (N_2064,N_1438,N_1734);
and U2065 (N_2065,N_1908,In_807);
or U2066 (N_2066,N_816,N_1275);
nor U2067 (N_2067,N_1880,N_612);
or U2068 (N_2068,N_1872,N_1998);
xor U2069 (N_2069,N_1620,N_1960);
and U2070 (N_2070,N_1855,N_1868);
and U2071 (N_2071,In_2379,N_1347);
and U2072 (N_2072,N_1580,N_1980);
or U2073 (N_2073,In_578,In_2454);
or U2074 (N_2074,N_1083,N_14);
or U2075 (N_2075,N_1825,N_1856);
nor U2076 (N_2076,N_269,N_1719);
or U2077 (N_2077,N_1754,N_1763);
nor U2078 (N_2078,N_1086,N_1953);
nor U2079 (N_2079,N_1277,N_716);
and U2080 (N_2080,N_1860,N_1543);
nand U2081 (N_2081,In_2286,N_1617);
and U2082 (N_2082,N_1744,N_1964);
nor U2083 (N_2083,N_1816,N_1785);
nand U2084 (N_2084,N_1815,In_1391);
nor U2085 (N_2085,N_194,In_919);
nand U2086 (N_2086,N_1931,N_1907);
nand U2087 (N_2087,N_1939,N_1841);
or U2088 (N_2088,N_1509,N_1934);
or U2089 (N_2089,N_1740,N_1784);
or U2090 (N_2090,N_1711,N_1905);
and U2091 (N_2091,N_1966,N_1712);
and U2092 (N_2092,N_1379,N_1997);
nand U2093 (N_2093,N_1827,In_349);
and U2094 (N_2094,N_1915,N_1977);
nor U2095 (N_2095,N_1875,N_1035);
nor U2096 (N_2096,N_1946,N_1929);
or U2097 (N_2097,N_1614,N_1793);
or U2098 (N_2098,N_1918,In_1001);
nand U2099 (N_2099,N_1106,N_1820);
nand U2100 (N_2100,In_1714,N_1913);
and U2101 (N_2101,N_1661,N_1976);
nand U2102 (N_2102,N_1456,N_1971);
and U2103 (N_2103,In_1279,N_1994);
nor U2104 (N_2104,N_1725,N_1076);
nor U2105 (N_2105,N_1577,N_992);
nand U2106 (N_2106,N_1799,N_1780);
nand U2107 (N_2107,N_1409,N_138);
nor U2108 (N_2108,N_1928,N_1573);
and U2109 (N_2109,N_1794,N_1983);
nand U2110 (N_2110,In_857,N_1508);
and U2111 (N_2111,N_1898,N_1967);
and U2112 (N_2112,N_1919,N_1687);
or U2113 (N_2113,N_1666,N_1537);
nor U2114 (N_2114,N_935,In_2242);
or U2115 (N_2115,N_1838,N_1781);
or U2116 (N_2116,N_1876,In_576);
or U2117 (N_2117,N_1556,N_1762);
or U2118 (N_2118,N_1959,N_1952);
and U2119 (N_2119,N_1853,N_1988);
nor U2120 (N_2120,N_1757,N_1399);
nor U2121 (N_2121,N_1937,In_778);
or U2122 (N_2122,N_1900,N_1265);
and U2123 (N_2123,N_1957,N_1768);
nor U2124 (N_2124,N_1832,N_1999);
nor U2125 (N_2125,N_1864,N_1904);
nand U2126 (N_2126,N_1321,N_1869);
nor U2127 (N_2127,In_675,N_1546);
nand U2128 (N_2128,In_2046,N_1705);
nand U2129 (N_2129,N_1802,N_1917);
nor U2130 (N_2130,In_1955,N_885);
nor U2131 (N_2131,N_1984,N_1778);
nor U2132 (N_2132,N_1982,N_1792);
nor U2133 (N_2133,N_1828,N_1990);
and U2134 (N_2134,N_1286,N_1502);
nor U2135 (N_2135,N_1958,N_1989);
nor U2136 (N_2136,N_1895,N_1281);
and U2137 (N_2137,N_1986,N_1759);
and U2138 (N_2138,N_1924,N_1515);
or U2139 (N_2139,N_1859,N_1696);
and U2140 (N_2140,N_1906,N_1318);
and U2141 (N_2141,N_613,N_1851);
nand U2142 (N_2142,N_1558,N_1442);
nand U2143 (N_2143,N_1498,N_1922);
or U2144 (N_2144,N_1426,N_1678);
nand U2145 (N_2145,N_1311,N_294);
nand U2146 (N_2146,In_691,N_1902);
nand U2147 (N_2147,N_1030,N_95);
or U2148 (N_2148,N_592,N_1846);
nand U2149 (N_2149,N_1723,N_1892);
nand U2150 (N_2150,N_1923,N_1758);
and U2151 (N_2151,N_1951,N_1316);
or U2152 (N_2152,N_1813,N_1972);
nor U2153 (N_2153,N_1284,N_1890);
xor U2154 (N_2154,N_1801,N_1731);
nor U2155 (N_2155,N_1480,N_1810);
nor U2156 (N_2156,N_1850,N_1773);
or U2157 (N_2157,N_1909,N_1581);
and U2158 (N_2158,N_1007,N_1791);
xor U2159 (N_2159,N_1239,N_1692);
nand U2160 (N_2160,N_1651,N_1992);
nand U2161 (N_2161,N_1969,N_1985);
and U2162 (N_2162,N_1874,N_1610);
or U2163 (N_2163,In_1532,N_963);
nor U2164 (N_2164,N_1807,N_1604);
and U2165 (N_2165,N_1970,N_822);
nand U2166 (N_2166,N_1839,N_1947);
nor U2167 (N_2167,In_1815,N_1555);
or U2168 (N_2168,N_1840,N_1942);
and U2169 (N_2169,N_1996,N_1819);
or U2170 (N_2170,N_1774,N_1746);
nand U2171 (N_2171,In_1909,N_805);
nor U2172 (N_2172,N_1787,N_1814);
nor U2173 (N_2173,N_1642,N_1866);
nand U2174 (N_2174,N_1736,N_1772);
and U2175 (N_2175,In_967,N_1829);
nand U2176 (N_2176,N_1579,N_1837);
or U2177 (N_2177,N_1914,N_1776);
nand U2178 (N_2178,N_1697,N_185);
or U2179 (N_2179,N_1752,N_1790);
nand U2180 (N_2180,N_1978,N_1812);
or U2181 (N_2181,N_1871,N_1783);
nand U2182 (N_2182,In_2452,N_1624);
nor U2183 (N_2183,N_323,N_1777);
nand U2184 (N_2184,N_1563,N_1669);
or U2185 (N_2185,N_1945,In_425);
nor U2186 (N_2186,N_1552,N_1842);
nand U2187 (N_2187,N_913,N_1598);
or U2188 (N_2188,N_1540,N_1077);
or U2189 (N_2189,N_1804,N_1897);
nor U2190 (N_2190,N_1821,In_702);
or U2191 (N_2191,N_1795,N_1920);
nor U2192 (N_2192,N_1925,N_1606);
and U2193 (N_2193,N_1295,N_1202);
nor U2194 (N_2194,N_1299,N_1803);
and U2195 (N_2195,N_1561,N_1926);
or U2196 (N_2196,N_1878,N_1760);
nor U2197 (N_2197,N_1538,N_1916);
nand U2198 (N_2198,N_1975,N_903);
nand U2199 (N_2199,N_1621,N_1769);
nor U2200 (N_2200,In_561,N_1309);
xor U2201 (N_2201,N_1933,In_2322);
or U2202 (N_2202,N_1685,N_1956);
and U2203 (N_2203,N_1333,N_1845);
and U2204 (N_2204,N_1938,N_1671);
nand U2205 (N_2205,N_519,N_1751);
and U2206 (N_2206,N_1808,In_2176);
or U2207 (N_2207,N_1993,N_1849);
or U2208 (N_2208,N_1615,N_1899);
nor U2209 (N_2209,In_818,N_1535);
and U2210 (N_2210,N_88,N_876);
nor U2211 (N_2211,N_1247,N_1154);
nand U2212 (N_2212,N_1564,N_1405);
nand U2213 (N_2213,N_1583,N_1782);
nor U2214 (N_2214,N_1941,N_32);
nor U2215 (N_2215,N_1987,N_1852);
nor U2216 (N_2216,N_1755,N_1308);
nor U2217 (N_2217,N_1227,N_378);
or U2218 (N_2218,N_1896,N_1973);
nor U2219 (N_2219,N_1186,N_1894);
or U2220 (N_2220,N_1949,N_1863);
nor U2221 (N_2221,N_1434,N_1401);
nand U2222 (N_2222,N_1764,In_238);
and U2223 (N_2223,N_1879,N_1329);
nand U2224 (N_2224,N_1817,N_33);
nand U2225 (N_2225,N_1532,N_1965);
or U2226 (N_2226,N_1024,N_1652);
and U2227 (N_2227,N_1514,N_650);
or U2228 (N_2228,N_1886,N_723);
and U2229 (N_2229,N_1979,N_1112);
and U2230 (N_2230,N_1779,N_1805);
nor U2231 (N_2231,N_1921,N_902);
or U2232 (N_2232,In_2198,N_1995);
or U2233 (N_2233,N_1962,N_1526);
nand U2234 (N_2234,N_1201,In_456);
and U2235 (N_2235,In_1051,N_1954);
or U2236 (N_2236,N_1823,In_68);
or U2237 (N_2237,N_1294,N_1861);
nor U2238 (N_2238,N_954,N_1811);
or U2239 (N_2239,N_1245,N_1533);
nand U2240 (N_2240,N_1707,N_1702);
nor U2241 (N_2241,N_1771,N_1796);
nor U2242 (N_2242,N_1885,N_1835);
or U2243 (N_2243,N_1756,N_1761);
nor U2244 (N_2244,N_632,N_1911);
nand U2245 (N_2245,N_1280,N_1903);
nor U2246 (N_2246,N_1289,N_1826);
and U2247 (N_2247,N_1180,In_545);
or U2248 (N_2248,N_1873,N_1833);
and U2249 (N_2249,N_1750,N_955);
or U2250 (N_2250,N_2166,N_2216);
nand U2251 (N_2251,N_2180,N_2025);
nor U2252 (N_2252,N_2042,N_2191);
nand U2253 (N_2253,N_2044,N_2228);
and U2254 (N_2254,N_2196,N_2176);
or U2255 (N_2255,N_2005,N_2215);
nand U2256 (N_2256,N_2072,N_2199);
or U2257 (N_2257,N_2062,N_2186);
and U2258 (N_2258,N_2011,N_2245);
nor U2259 (N_2259,N_2134,N_2095);
or U2260 (N_2260,N_2087,N_2202);
nand U2261 (N_2261,N_2093,N_2084);
nor U2262 (N_2262,N_2157,N_2123);
or U2263 (N_2263,N_2117,N_2225);
or U2264 (N_2264,N_2097,N_2089);
and U2265 (N_2265,N_2231,N_2086);
and U2266 (N_2266,N_2066,N_2079);
nor U2267 (N_2267,N_2107,N_2161);
nand U2268 (N_2268,N_2001,N_2160);
nor U2269 (N_2269,N_2131,N_2125);
or U2270 (N_2270,N_2081,N_2187);
nand U2271 (N_2271,N_2047,N_2181);
and U2272 (N_2272,N_2092,N_2090);
or U2273 (N_2273,N_2221,N_2050);
or U2274 (N_2274,N_2068,N_2164);
xnor U2275 (N_2275,N_2034,N_2113);
nor U2276 (N_2276,N_2155,N_2008);
nor U2277 (N_2277,N_2061,N_2183);
nand U2278 (N_2278,N_2041,N_2153);
nand U2279 (N_2279,N_2003,N_2165);
nand U2280 (N_2280,N_2185,N_2060);
and U2281 (N_2281,N_2057,N_2067);
and U2282 (N_2282,N_2096,N_2237);
or U2283 (N_2283,N_2129,N_2082);
nor U2284 (N_2284,N_2158,N_2145);
and U2285 (N_2285,N_2031,N_2218);
and U2286 (N_2286,N_2065,N_2208);
nand U2287 (N_2287,N_2171,N_2154);
nand U2288 (N_2288,N_2249,N_2172);
or U2289 (N_2289,N_2136,N_2120);
nand U2290 (N_2290,N_2132,N_2207);
nand U2291 (N_2291,N_2007,N_2016);
and U2292 (N_2292,N_2211,N_2178);
nor U2293 (N_2293,N_2054,N_2053);
nand U2294 (N_2294,N_2233,N_2073);
or U2295 (N_2295,N_2106,N_2241);
and U2296 (N_2296,N_2023,N_2190);
or U2297 (N_2297,N_2217,N_2052);
and U2298 (N_2298,N_2204,N_2130);
nor U2299 (N_2299,N_2213,N_2243);
nor U2300 (N_2300,N_2116,N_2159);
nand U2301 (N_2301,N_2247,N_2197);
nor U2302 (N_2302,N_2017,N_2006);
nand U2303 (N_2303,N_2040,N_2173);
nand U2304 (N_2304,N_2142,N_2015);
nand U2305 (N_2305,N_2032,N_2019);
nand U2306 (N_2306,N_2168,N_2102);
nor U2307 (N_2307,N_2058,N_2140);
and U2308 (N_2308,N_2144,N_2021);
nor U2309 (N_2309,N_2198,N_2009);
and U2310 (N_2310,N_2075,N_2244);
nand U2311 (N_2311,N_2105,N_2056);
nand U2312 (N_2312,N_2012,N_2043);
or U2313 (N_2313,N_2045,N_2220);
or U2314 (N_2314,N_2020,N_2029);
nand U2315 (N_2315,N_2018,N_2000);
nand U2316 (N_2316,N_2030,N_2046);
or U2317 (N_2317,N_2163,N_2024);
nor U2318 (N_2318,N_2119,N_2078);
and U2319 (N_2319,N_2112,N_2088);
and U2320 (N_2320,N_2195,N_2010);
and U2321 (N_2321,N_2039,N_2121);
and U2322 (N_2322,N_2122,N_2246);
and U2323 (N_2323,N_2004,N_2169);
and U2324 (N_2324,N_2035,N_2242);
nor U2325 (N_2325,N_2209,N_2049);
nor U2326 (N_2326,N_2074,N_2110);
nand U2327 (N_2327,N_2222,N_2240);
or U2328 (N_2328,N_2126,N_2036);
or U2329 (N_2329,N_2149,N_2162);
or U2330 (N_2330,N_2192,N_2139);
or U2331 (N_2331,N_2177,N_2069);
or U2332 (N_2332,N_2064,N_2059);
and U2333 (N_2333,N_2238,N_2174);
nor U2334 (N_2334,N_2135,N_2170);
and U2335 (N_2335,N_2002,N_2219);
nor U2336 (N_2336,N_2234,N_2212);
and U2337 (N_2337,N_2103,N_2115);
or U2338 (N_2338,N_2137,N_2205);
and U2339 (N_2339,N_2227,N_2232);
nand U2340 (N_2340,N_2083,N_2239);
and U2341 (N_2341,N_2152,N_2055);
or U2342 (N_2342,N_2048,N_2108);
xnor U2343 (N_2343,N_2099,N_2114);
or U2344 (N_2344,N_2229,N_2070);
or U2345 (N_2345,N_2148,N_2167);
and U2346 (N_2346,N_2100,N_2098);
nor U2347 (N_2347,N_2013,N_2214);
or U2348 (N_2348,N_2193,N_2182);
and U2349 (N_2349,N_2014,N_2179);
nand U2350 (N_2350,N_2037,N_2194);
and U2351 (N_2351,N_2150,N_2080);
and U2352 (N_2352,N_2128,N_2071);
or U2353 (N_2353,N_2077,N_2210);
and U2354 (N_2354,N_2091,N_2141);
or U2355 (N_2355,N_2230,N_2184);
nand U2356 (N_2356,N_2203,N_2201);
and U2357 (N_2357,N_2111,N_2109);
nor U2358 (N_2358,N_2063,N_2189);
or U2359 (N_2359,N_2133,N_2101);
nand U2360 (N_2360,N_2188,N_2248);
nand U2361 (N_2361,N_2235,N_2156);
nor U2362 (N_2362,N_2027,N_2146);
and U2363 (N_2363,N_2200,N_2028);
and U2364 (N_2364,N_2033,N_2124);
nor U2365 (N_2365,N_2226,N_2118);
or U2366 (N_2366,N_2104,N_2138);
or U2367 (N_2367,N_2151,N_2175);
or U2368 (N_2368,N_2022,N_2206);
and U2369 (N_2369,N_2127,N_2143);
nand U2370 (N_2370,N_2147,N_2038);
or U2371 (N_2371,N_2076,N_2223);
and U2372 (N_2372,N_2026,N_2236);
nand U2373 (N_2373,N_2051,N_2224);
and U2374 (N_2374,N_2094,N_2085);
nor U2375 (N_2375,N_2222,N_2234);
nor U2376 (N_2376,N_2112,N_2076);
nor U2377 (N_2377,N_2014,N_2127);
nor U2378 (N_2378,N_2169,N_2107);
and U2379 (N_2379,N_2053,N_2222);
and U2380 (N_2380,N_2100,N_2114);
and U2381 (N_2381,N_2047,N_2218);
nand U2382 (N_2382,N_2209,N_2238);
or U2383 (N_2383,N_2180,N_2103);
xor U2384 (N_2384,N_2176,N_2089);
xnor U2385 (N_2385,N_2151,N_2002);
nand U2386 (N_2386,N_2181,N_2157);
or U2387 (N_2387,N_2242,N_2212);
or U2388 (N_2388,N_2076,N_2169);
nand U2389 (N_2389,N_2043,N_2144);
and U2390 (N_2390,N_2219,N_2218);
or U2391 (N_2391,N_2142,N_2086);
nand U2392 (N_2392,N_2037,N_2226);
nand U2393 (N_2393,N_2009,N_2027);
nand U2394 (N_2394,N_2178,N_2245);
or U2395 (N_2395,N_2114,N_2106);
and U2396 (N_2396,N_2014,N_2094);
or U2397 (N_2397,N_2240,N_2173);
and U2398 (N_2398,N_2066,N_2012);
and U2399 (N_2399,N_2214,N_2206);
nand U2400 (N_2400,N_2243,N_2140);
or U2401 (N_2401,N_2029,N_2031);
nand U2402 (N_2402,N_2062,N_2035);
nand U2403 (N_2403,N_2183,N_2113);
nor U2404 (N_2404,N_2184,N_2065);
nand U2405 (N_2405,N_2147,N_2135);
and U2406 (N_2406,N_2228,N_2156);
nor U2407 (N_2407,N_2183,N_2009);
xnor U2408 (N_2408,N_2190,N_2070);
and U2409 (N_2409,N_2006,N_2228);
nor U2410 (N_2410,N_2209,N_2080);
nor U2411 (N_2411,N_2051,N_2136);
nor U2412 (N_2412,N_2170,N_2226);
and U2413 (N_2413,N_2106,N_2148);
or U2414 (N_2414,N_2051,N_2205);
or U2415 (N_2415,N_2096,N_2011);
nor U2416 (N_2416,N_2187,N_2079);
nor U2417 (N_2417,N_2136,N_2188);
or U2418 (N_2418,N_2027,N_2144);
and U2419 (N_2419,N_2010,N_2015);
or U2420 (N_2420,N_2198,N_2196);
nand U2421 (N_2421,N_2066,N_2054);
and U2422 (N_2422,N_2141,N_2239);
nor U2423 (N_2423,N_2120,N_2173);
or U2424 (N_2424,N_2204,N_2076);
and U2425 (N_2425,N_2146,N_2060);
nand U2426 (N_2426,N_2114,N_2121);
and U2427 (N_2427,N_2194,N_2116);
nand U2428 (N_2428,N_2016,N_2179);
and U2429 (N_2429,N_2048,N_2172);
and U2430 (N_2430,N_2091,N_2195);
nor U2431 (N_2431,N_2136,N_2119);
nor U2432 (N_2432,N_2100,N_2235);
nand U2433 (N_2433,N_2238,N_2013);
nor U2434 (N_2434,N_2064,N_2107);
nand U2435 (N_2435,N_2137,N_2003);
nor U2436 (N_2436,N_2123,N_2220);
or U2437 (N_2437,N_2078,N_2018);
nor U2438 (N_2438,N_2245,N_2157);
nor U2439 (N_2439,N_2143,N_2016);
nand U2440 (N_2440,N_2212,N_2171);
nand U2441 (N_2441,N_2170,N_2174);
nand U2442 (N_2442,N_2205,N_2236);
nand U2443 (N_2443,N_2183,N_2241);
and U2444 (N_2444,N_2123,N_2101);
and U2445 (N_2445,N_2074,N_2089);
nor U2446 (N_2446,N_2075,N_2098);
nor U2447 (N_2447,N_2046,N_2248);
or U2448 (N_2448,N_2036,N_2133);
or U2449 (N_2449,N_2018,N_2047);
or U2450 (N_2450,N_2200,N_2064);
and U2451 (N_2451,N_2066,N_2002);
nand U2452 (N_2452,N_2138,N_2006);
or U2453 (N_2453,N_2240,N_2187);
nor U2454 (N_2454,N_2197,N_2160);
or U2455 (N_2455,N_2168,N_2195);
and U2456 (N_2456,N_2070,N_2072);
and U2457 (N_2457,N_2071,N_2069);
nor U2458 (N_2458,N_2181,N_2220);
and U2459 (N_2459,N_2182,N_2121);
and U2460 (N_2460,N_2095,N_2237);
nand U2461 (N_2461,N_2054,N_2213);
nor U2462 (N_2462,N_2151,N_2000);
or U2463 (N_2463,N_2029,N_2150);
or U2464 (N_2464,N_2230,N_2090);
or U2465 (N_2465,N_2028,N_2171);
nor U2466 (N_2466,N_2189,N_2135);
nand U2467 (N_2467,N_2064,N_2186);
or U2468 (N_2468,N_2115,N_2233);
nand U2469 (N_2469,N_2017,N_2203);
nand U2470 (N_2470,N_2007,N_2198);
and U2471 (N_2471,N_2057,N_2024);
nor U2472 (N_2472,N_2077,N_2023);
nor U2473 (N_2473,N_2144,N_2207);
nor U2474 (N_2474,N_2065,N_2115);
nand U2475 (N_2475,N_2224,N_2034);
nand U2476 (N_2476,N_2048,N_2144);
nor U2477 (N_2477,N_2044,N_2163);
or U2478 (N_2478,N_2187,N_2162);
and U2479 (N_2479,N_2210,N_2066);
xor U2480 (N_2480,N_2057,N_2003);
or U2481 (N_2481,N_2043,N_2193);
and U2482 (N_2482,N_2200,N_2196);
nand U2483 (N_2483,N_2245,N_2193);
and U2484 (N_2484,N_2224,N_2164);
nand U2485 (N_2485,N_2083,N_2045);
and U2486 (N_2486,N_2238,N_2242);
or U2487 (N_2487,N_2067,N_2092);
nor U2488 (N_2488,N_2186,N_2145);
nand U2489 (N_2489,N_2118,N_2057);
or U2490 (N_2490,N_2056,N_2144);
nor U2491 (N_2491,N_2072,N_2131);
nand U2492 (N_2492,N_2063,N_2117);
nand U2493 (N_2493,N_2118,N_2228);
nor U2494 (N_2494,N_2106,N_2160);
or U2495 (N_2495,N_2023,N_2043);
or U2496 (N_2496,N_2189,N_2181);
or U2497 (N_2497,N_2045,N_2211);
or U2498 (N_2498,N_2186,N_2198);
and U2499 (N_2499,N_2108,N_2089);
and U2500 (N_2500,N_2345,N_2462);
nand U2501 (N_2501,N_2370,N_2346);
or U2502 (N_2502,N_2453,N_2431);
nor U2503 (N_2503,N_2268,N_2418);
and U2504 (N_2504,N_2380,N_2467);
nor U2505 (N_2505,N_2296,N_2269);
or U2506 (N_2506,N_2434,N_2363);
or U2507 (N_2507,N_2419,N_2498);
or U2508 (N_2508,N_2396,N_2417);
nor U2509 (N_2509,N_2459,N_2320);
nor U2510 (N_2510,N_2339,N_2325);
and U2511 (N_2511,N_2415,N_2294);
and U2512 (N_2512,N_2482,N_2350);
nor U2513 (N_2513,N_2366,N_2272);
nand U2514 (N_2514,N_2359,N_2303);
nor U2515 (N_2515,N_2460,N_2440);
or U2516 (N_2516,N_2421,N_2435);
and U2517 (N_2517,N_2316,N_2284);
or U2518 (N_2518,N_2429,N_2321);
nand U2519 (N_2519,N_2483,N_2495);
and U2520 (N_2520,N_2331,N_2456);
nor U2521 (N_2521,N_2463,N_2376);
nand U2522 (N_2522,N_2414,N_2277);
nand U2523 (N_2523,N_2259,N_2281);
and U2524 (N_2524,N_2261,N_2494);
or U2525 (N_2525,N_2365,N_2478);
or U2526 (N_2526,N_2403,N_2423);
nand U2527 (N_2527,N_2258,N_2420);
nand U2528 (N_2528,N_2322,N_2445);
or U2529 (N_2529,N_2274,N_2323);
and U2530 (N_2530,N_2324,N_2471);
nor U2531 (N_2531,N_2399,N_2279);
xnor U2532 (N_2532,N_2355,N_2369);
nor U2533 (N_2533,N_2464,N_2298);
nor U2534 (N_2534,N_2338,N_2461);
nand U2535 (N_2535,N_2449,N_2314);
nor U2536 (N_2536,N_2476,N_2313);
nor U2537 (N_2537,N_2457,N_2254);
and U2538 (N_2538,N_2336,N_2477);
nand U2539 (N_2539,N_2319,N_2271);
and U2540 (N_2540,N_2291,N_2302);
or U2541 (N_2541,N_2406,N_2288);
nand U2542 (N_2542,N_2315,N_2264);
or U2543 (N_2543,N_2391,N_2489);
nand U2544 (N_2544,N_2437,N_2454);
nor U2545 (N_2545,N_2310,N_2341);
nor U2546 (N_2546,N_2260,N_2416);
nand U2547 (N_2547,N_2468,N_2424);
or U2548 (N_2548,N_2358,N_2330);
or U2549 (N_2549,N_2318,N_2446);
nand U2550 (N_2550,N_2308,N_2390);
nor U2551 (N_2551,N_2262,N_2295);
or U2552 (N_2552,N_2328,N_2436);
and U2553 (N_2553,N_2304,N_2250);
or U2554 (N_2554,N_2301,N_2401);
and U2555 (N_2555,N_2475,N_2356);
or U2556 (N_2556,N_2251,N_2493);
or U2557 (N_2557,N_2469,N_2388);
nand U2558 (N_2558,N_2337,N_2387);
nor U2559 (N_2559,N_2379,N_2381);
or U2560 (N_2560,N_2367,N_2492);
nor U2561 (N_2561,N_2427,N_2497);
or U2562 (N_2562,N_2344,N_2430);
nor U2563 (N_2563,N_2480,N_2293);
and U2564 (N_2564,N_2364,N_2486);
nor U2565 (N_2565,N_2299,N_2395);
nor U2566 (N_2566,N_2402,N_2317);
nor U2567 (N_2567,N_2253,N_2392);
or U2568 (N_2568,N_2394,N_2273);
and U2569 (N_2569,N_2263,N_2485);
nand U2570 (N_2570,N_2404,N_2428);
or U2571 (N_2571,N_2285,N_2289);
or U2572 (N_2572,N_2408,N_2479);
nand U2573 (N_2573,N_2373,N_2267);
nor U2574 (N_2574,N_2278,N_2466);
or U2575 (N_2575,N_2411,N_2342);
or U2576 (N_2576,N_2287,N_2286);
and U2577 (N_2577,N_2398,N_2487);
and U2578 (N_2578,N_2374,N_2305);
and U2579 (N_2579,N_2270,N_2362);
nand U2580 (N_2580,N_2306,N_2326);
or U2581 (N_2581,N_2265,N_2409);
nand U2582 (N_2582,N_2474,N_2333);
and U2583 (N_2583,N_2472,N_2451);
nand U2584 (N_2584,N_2255,N_2292);
and U2585 (N_2585,N_2389,N_2343);
nor U2586 (N_2586,N_2276,N_2443);
or U2587 (N_2587,N_2252,N_2332);
nor U2588 (N_2588,N_2432,N_2499);
nand U2589 (N_2589,N_2452,N_2385);
nor U2590 (N_2590,N_2307,N_2384);
nor U2591 (N_2591,N_2327,N_2282);
and U2592 (N_2592,N_2377,N_2257);
or U2593 (N_2593,N_2484,N_2439);
and U2594 (N_2594,N_2393,N_2256);
or U2595 (N_2595,N_2354,N_2300);
nor U2596 (N_2596,N_2349,N_2413);
or U2597 (N_2597,N_2351,N_2422);
or U2598 (N_2598,N_2496,N_2455);
or U2599 (N_2599,N_2378,N_2400);
and U2600 (N_2600,N_2371,N_2412);
nor U2601 (N_2601,N_2426,N_2386);
and U2602 (N_2602,N_2438,N_2410);
nand U2603 (N_2603,N_2481,N_2335);
xnor U2604 (N_2604,N_2357,N_2458);
and U2605 (N_2605,N_2447,N_2407);
nand U2606 (N_2606,N_2450,N_2340);
or U2607 (N_2607,N_2372,N_2353);
nand U2608 (N_2608,N_2329,N_2290);
nand U2609 (N_2609,N_2425,N_2441);
nand U2610 (N_2610,N_2311,N_2383);
and U2611 (N_2611,N_2334,N_2297);
or U2612 (N_2612,N_2442,N_2490);
or U2613 (N_2613,N_2382,N_2280);
or U2614 (N_2614,N_2312,N_2360);
nand U2615 (N_2615,N_2444,N_2465);
xor U2616 (N_2616,N_2347,N_2352);
or U2617 (N_2617,N_2266,N_2309);
and U2618 (N_2618,N_2375,N_2348);
nor U2619 (N_2619,N_2448,N_2275);
nor U2620 (N_2620,N_2397,N_2283);
and U2621 (N_2621,N_2368,N_2433);
or U2622 (N_2622,N_2405,N_2491);
nand U2623 (N_2623,N_2361,N_2470);
nand U2624 (N_2624,N_2488,N_2473);
and U2625 (N_2625,N_2261,N_2447);
and U2626 (N_2626,N_2365,N_2491);
and U2627 (N_2627,N_2265,N_2443);
nand U2628 (N_2628,N_2479,N_2462);
nor U2629 (N_2629,N_2291,N_2383);
and U2630 (N_2630,N_2360,N_2282);
or U2631 (N_2631,N_2339,N_2329);
and U2632 (N_2632,N_2332,N_2255);
or U2633 (N_2633,N_2273,N_2427);
nand U2634 (N_2634,N_2328,N_2404);
nand U2635 (N_2635,N_2363,N_2466);
nand U2636 (N_2636,N_2273,N_2379);
nand U2637 (N_2637,N_2456,N_2274);
or U2638 (N_2638,N_2287,N_2337);
nand U2639 (N_2639,N_2275,N_2270);
nand U2640 (N_2640,N_2416,N_2350);
nor U2641 (N_2641,N_2285,N_2318);
and U2642 (N_2642,N_2381,N_2289);
nand U2643 (N_2643,N_2446,N_2426);
xnor U2644 (N_2644,N_2399,N_2428);
nand U2645 (N_2645,N_2259,N_2326);
nand U2646 (N_2646,N_2277,N_2421);
nand U2647 (N_2647,N_2353,N_2340);
nand U2648 (N_2648,N_2458,N_2471);
nand U2649 (N_2649,N_2421,N_2272);
nor U2650 (N_2650,N_2312,N_2446);
or U2651 (N_2651,N_2417,N_2387);
and U2652 (N_2652,N_2468,N_2287);
nand U2653 (N_2653,N_2313,N_2478);
or U2654 (N_2654,N_2440,N_2312);
nor U2655 (N_2655,N_2366,N_2267);
nor U2656 (N_2656,N_2494,N_2445);
or U2657 (N_2657,N_2457,N_2389);
or U2658 (N_2658,N_2310,N_2277);
nand U2659 (N_2659,N_2446,N_2273);
nor U2660 (N_2660,N_2451,N_2262);
nand U2661 (N_2661,N_2335,N_2442);
nor U2662 (N_2662,N_2304,N_2471);
nand U2663 (N_2663,N_2499,N_2383);
nand U2664 (N_2664,N_2470,N_2350);
and U2665 (N_2665,N_2386,N_2251);
nand U2666 (N_2666,N_2411,N_2419);
or U2667 (N_2667,N_2298,N_2361);
or U2668 (N_2668,N_2450,N_2457);
or U2669 (N_2669,N_2479,N_2383);
and U2670 (N_2670,N_2496,N_2296);
and U2671 (N_2671,N_2325,N_2442);
nor U2672 (N_2672,N_2412,N_2260);
and U2673 (N_2673,N_2311,N_2442);
or U2674 (N_2674,N_2320,N_2285);
nor U2675 (N_2675,N_2498,N_2314);
and U2676 (N_2676,N_2254,N_2317);
nand U2677 (N_2677,N_2368,N_2423);
or U2678 (N_2678,N_2267,N_2325);
or U2679 (N_2679,N_2363,N_2338);
nor U2680 (N_2680,N_2349,N_2289);
nand U2681 (N_2681,N_2426,N_2398);
nor U2682 (N_2682,N_2427,N_2417);
nand U2683 (N_2683,N_2460,N_2259);
nand U2684 (N_2684,N_2332,N_2375);
or U2685 (N_2685,N_2319,N_2266);
nand U2686 (N_2686,N_2468,N_2484);
and U2687 (N_2687,N_2402,N_2311);
nor U2688 (N_2688,N_2340,N_2451);
nor U2689 (N_2689,N_2330,N_2452);
and U2690 (N_2690,N_2360,N_2256);
nand U2691 (N_2691,N_2341,N_2381);
nor U2692 (N_2692,N_2499,N_2483);
nand U2693 (N_2693,N_2434,N_2476);
or U2694 (N_2694,N_2351,N_2499);
or U2695 (N_2695,N_2285,N_2269);
nand U2696 (N_2696,N_2290,N_2412);
nand U2697 (N_2697,N_2367,N_2260);
and U2698 (N_2698,N_2328,N_2475);
nor U2699 (N_2699,N_2473,N_2446);
or U2700 (N_2700,N_2291,N_2388);
or U2701 (N_2701,N_2275,N_2428);
and U2702 (N_2702,N_2298,N_2325);
or U2703 (N_2703,N_2285,N_2315);
or U2704 (N_2704,N_2421,N_2314);
nor U2705 (N_2705,N_2332,N_2330);
nor U2706 (N_2706,N_2358,N_2354);
and U2707 (N_2707,N_2253,N_2350);
nand U2708 (N_2708,N_2313,N_2396);
nand U2709 (N_2709,N_2463,N_2250);
and U2710 (N_2710,N_2356,N_2404);
nor U2711 (N_2711,N_2376,N_2434);
or U2712 (N_2712,N_2283,N_2285);
nand U2713 (N_2713,N_2282,N_2332);
and U2714 (N_2714,N_2469,N_2459);
nand U2715 (N_2715,N_2482,N_2434);
nand U2716 (N_2716,N_2352,N_2426);
nand U2717 (N_2717,N_2400,N_2333);
nand U2718 (N_2718,N_2448,N_2393);
or U2719 (N_2719,N_2392,N_2280);
or U2720 (N_2720,N_2470,N_2267);
and U2721 (N_2721,N_2286,N_2432);
or U2722 (N_2722,N_2296,N_2386);
and U2723 (N_2723,N_2388,N_2472);
nor U2724 (N_2724,N_2253,N_2446);
or U2725 (N_2725,N_2347,N_2397);
nor U2726 (N_2726,N_2498,N_2397);
or U2727 (N_2727,N_2258,N_2418);
or U2728 (N_2728,N_2321,N_2308);
or U2729 (N_2729,N_2335,N_2463);
nand U2730 (N_2730,N_2436,N_2409);
and U2731 (N_2731,N_2433,N_2412);
or U2732 (N_2732,N_2319,N_2341);
nand U2733 (N_2733,N_2476,N_2294);
or U2734 (N_2734,N_2309,N_2430);
nor U2735 (N_2735,N_2445,N_2273);
or U2736 (N_2736,N_2299,N_2429);
or U2737 (N_2737,N_2316,N_2299);
or U2738 (N_2738,N_2344,N_2390);
or U2739 (N_2739,N_2487,N_2311);
nand U2740 (N_2740,N_2310,N_2484);
nand U2741 (N_2741,N_2309,N_2437);
nand U2742 (N_2742,N_2473,N_2346);
and U2743 (N_2743,N_2341,N_2462);
nand U2744 (N_2744,N_2274,N_2362);
nor U2745 (N_2745,N_2316,N_2457);
or U2746 (N_2746,N_2383,N_2271);
or U2747 (N_2747,N_2428,N_2309);
and U2748 (N_2748,N_2325,N_2381);
and U2749 (N_2749,N_2320,N_2252);
nor U2750 (N_2750,N_2626,N_2550);
and U2751 (N_2751,N_2599,N_2566);
nand U2752 (N_2752,N_2523,N_2624);
nand U2753 (N_2753,N_2597,N_2607);
nor U2754 (N_2754,N_2587,N_2501);
nand U2755 (N_2755,N_2743,N_2661);
and U2756 (N_2756,N_2514,N_2683);
or U2757 (N_2757,N_2533,N_2672);
nor U2758 (N_2758,N_2507,N_2530);
and U2759 (N_2759,N_2719,N_2736);
nor U2760 (N_2760,N_2679,N_2608);
nand U2761 (N_2761,N_2625,N_2724);
and U2762 (N_2762,N_2594,N_2572);
nand U2763 (N_2763,N_2521,N_2742);
nor U2764 (N_2764,N_2657,N_2706);
and U2765 (N_2765,N_2580,N_2637);
nor U2766 (N_2766,N_2729,N_2581);
and U2767 (N_2767,N_2583,N_2745);
nand U2768 (N_2768,N_2635,N_2524);
nor U2769 (N_2769,N_2603,N_2703);
and U2770 (N_2770,N_2554,N_2696);
nor U2771 (N_2771,N_2663,N_2713);
and U2772 (N_2772,N_2722,N_2548);
and U2773 (N_2773,N_2646,N_2668);
nor U2774 (N_2774,N_2666,N_2688);
nand U2775 (N_2775,N_2588,N_2670);
or U2776 (N_2776,N_2546,N_2552);
or U2777 (N_2777,N_2674,N_2553);
or U2778 (N_2778,N_2731,N_2676);
and U2779 (N_2779,N_2565,N_2701);
or U2780 (N_2780,N_2694,N_2601);
and U2781 (N_2781,N_2615,N_2623);
nor U2782 (N_2782,N_2611,N_2718);
and U2783 (N_2783,N_2658,N_2505);
and U2784 (N_2784,N_2631,N_2741);
or U2785 (N_2785,N_2629,N_2602);
nand U2786 (N_2786,N_2520,N_2700);
and U2787 (N_2787,N_2617,N_2705);
nand U2788 (N_2788,N_2544,N_2571);
and U2789 (N_2789,N_2606,N_2709);
nor U2790 (N_2790,N_2564,N_2695);
and U2791 (N_2791,N_2522,N_2515);
xor U2792 (N_2792,N_2728,N_2711);
and U2793 (N_2793,N_2538,N_2641);
nor U2794 (N_2794,N_2627,N_2585);
or U2795 (N_2795,N_2577,N_2567);
and U2796 (N_2796,N_2531,N_2690);
and U2797 (N_2797,N_2612,N_2734);
nand U2798 (N_2798,N_2730,N_2500);
nor U2799 (N_2799,N_2595,N_2662);
and U2800 (N_2800,N_2503,N_2532);
and U2801 (N_2801,N_2737,N_2687);
nor U2802 (N_2802,N_2526,N_2525);
nor U2803 (N_2803,N_2653,N_2575);
and U2804 (N_2804,N_2621,N_2632);
nor U2805 (N_2805,N_2638,N_2639);
or U2806 (N_2806,N_2513,N_2673);
nor U2807 (N_2807,N_2685,N_2746);
nand U2808 (N_2808,N_2568,N_2618);
nor U2809 (N_2809,N_2576,N_2504);
nor U2810 (N_2810,N_2691,N_2678);
or U2811 (N_2811,N_2593,N_2714);
or U2812 (N_2812,N_2682,N_2630);
nor U2813 (N_2813,N_2735,N_2622);
or U2814 (N_2814,N_2647,N_2535);
nor U2815 (N_2815,N_2508,N_2651);
nor U2816 (N_2816,N_2667,N_2697);
nand U2817 (N_2817,N_2640,N_2733);
or U2818 (N_2818,N_2652,N_2708);
or U2819 (N_2819,N_2675,N_2547);
and U2820 (N_2820,N_2726,N_2649);
nor U2821 (N_2821,N_2592,N_2720);
and U2822 (N_2822,N_2570,N_2738);
or U2823 (N_2823,N_2536,N_2616);
nor U2824 (N_2824,N_2613,N_2643);
or U2825 (N_2825,N_2671,N_2557);
nand U2826 (N_2826,N_2555,N_2702);
nand U2827 (N_2827,N_2528,N_2614);
or U2828 (N_2828,N_2739,N_2549);
nor U2829 (N_2829,N_2609,N_2744);
and U2830 (N_2830,N_2740,N_2534);
nand U2831 (N_2831,N_2610,N_2732);
nand U2832 (N_2832,N_2582,N_2749);
and U2833 (N_2833,N_2509,N_2656);
xor U2834 (N_2834,N_2655,N_2654);
nand U2835 (N_2835,N_2692,N_2681);
nand U2836 (N_2836,N_2727,N_2512);
and U2837 (N_2837,N_2619,N_2573);
nor U2838 (N_2838,N_2669,N_2605);
nor U2839 (N_2839,N_2644,N_2725);
and U2840 (N_2840,N_2551,N_2712);
nor U2841 (N_2841,N_2586,N_2707);
nand U2842 (N_2842,N_2541,N_2559);
nand U2843 (N_2843,N_2511,N_2529);
and U2844 (N_2844,N_2604,N_2715);
or U2845 (N_2845,N_2596,N_2589);
nand U2846 (N_2846,N_2636,N_2648);
nor U2847 (N_2847,N_2600,N_2628);
and U2848 (N_2848,N_2723,N_2693);
and U2849 (N_2849,N_2545,N_2689);
and U2850 (N_2850,N_2584,N_2516);
and U2851 (N_2851,N_2562,N_2716);
or U2852 (N_2852,N_2517,N_2699);
or U2853 (N_2853,N_2680,N_2748);
and U2854 (N_2854,N_2704,N_2634);
nor U2855 (N_2855,N_2558,N_2633);
or U2856 (N_2856,N_2502,N_2747);
and U2857 (N_2857,N_2506,N_2578);
nand U2858 (N_2858,N_2569,N_2560);
nor U2859 (N_2859,N_2518,N_2537);
or U2860 (N_2860,N_2543,N_2684);
or U2861 (N_2861,N_2642,N_2664);
or U2862 (N_2862,N_2519,N_2561);
and U2863 (N_2863,N_2645,N_2721);
nor U2864 (N_2864,N_2591,N_2527);
and U2865 (N_2865,N_2563,N_2717);
nor U2866 (N_2866,N_2556,N_2698);
or U2867 (N_2867,N_2542,N_2540);
or U2868 (N_2868,N_2510,N_2539);
nand U2869 (N_2869,N_2598,N_2650);
nand U2870 (N_2870,N_2590,N_2574);
or U2871 (N_2871,N_2579,N_2710);
or U2872 (N_2872,N_2659,N_2665);
nand U2873 (N_2873,N_2620,N_2686);
or U2874 (N_2874,N_2660,N_2677);
or U2875 (N_2875,N_2598,N_2725);
and U2876 (N_2876,N_2615,N_2710);
or U2877 (N_2877,N_2662,N_2741);
nor U2878 (N_2878,N_2617,N_2736);
nor U2879 (N_2879,N_2606,N_2735);
or U2880 (N_2880,N_2641,N_2577);
and U2881 (N_2881,N_2606,N_2511);
nor U2882 (N_2882,N_2605,N_2676);
nor U2883 (N_2883,N_2746,N_2706);
nand U2884 (N_2884,N_2600,N_2575);
xnor U2885 (N_2885,N_2724,N_2660);
and U2886 (N_2886,N_2597,N_2533);
nor U2887 (N_2887,N_2613,N_2550);
nand U2888 (N_2888,N_2520,N_2540);
nand U2889 (N_2889,N_2557,N_2740);
nand U2890 (N_2890,N_2653,N_2748);
nor U2891 (N_2891,N_2732,N_2605);
nor U2892 (N_2892,N_2686,N_2555);
nor U2893 (N_2893,N_2730,N_2648);
nand U2894 (N_2894,N_2634,N_2685);
or U2895 (N_2895,N_2535,N_2566);
or U2896 (N_2896,N_2672,N_2539);
and U2897 (N_2897,N_2580,N_2697);
nand U2898 (N_2898,N_2565,N_2698);
nor U2899 (N_2899,N_2593,N_2689);
or U2900 (N_2900,N_2645,N_2543);
and U2901 (N_2901,N_2660,N_2669);
nor U2902 (N_2902,N_2530,N_2536);
and U2903 (N_2903,N_2591,N_2700);
and U2904 (N_2904,N_2740,N_2735);
or U2905 (N_2905,N_2694,N_2684);
or U2906 (N_2906,N_2596,N_2709);
or U2907 (N_2907,N_2527,N_2674);
or U2908 (N_2908,N_2587,N_2685);
nor U2909 (N_2909,N_2740,N_2714);
or U2910 (N_2910,N_2572,N_2671);
or U2911 (N_2911,N_2739,N_2717);
or U2912 (N_2912,N_2704,N_2516);
nand U2913 (N_2913,N_2680,N_2601);
and U2914 (N_2914,N_2585,N_2593);
nor U2915 (N_2915,N_2721,N_2581);
nor U2916 (N_2916,N_2719,N_2660);
and U2917 (N_2917,N_2718,N_2693);
nand U2918 (N_2918,N_2534,N_2712);
and U2919 (N_2919,N_2732,N_2532);
nand U2920 (N_2920,N_2633,N_2586);
and U2921 (N_2921,N_2720,N_2581);
nand U2922 (N_2922,N_2703,N_2535);
or U2923 (N_2923,N_2557,N_2595);
nand U2924 (N_2924,N_2545,N_2669);
or U2925 (N_2925,N_2702,N_2587);
nor U2926 (N_2926,N_2528,N_2579);
nor U2927 (N_2927,N_2703,N_2700);
nor U2928 (N_2928,N_2691,N_2699);
and U2929 (N_2929,N_2511,N_2551);
nand U2930 (N_2930,N_2559,N_2725);
nand U2931 (N_2931,N_2547,N_2705);
nor U2932 (N_2932,N_2557,N_2694);
or U2933 (N_2933,N_2602,N_2661);
and U2934 (N_2934,N_2736,N_2667);
nand U2935 (N_2935,N_2655,N_2580);
nand U2936 (N_2936,N_2564,N_2559);
nand U2937 (N_2937,N_2518,N_2650);
and U2938 (N_2938,N_2546,N_2586);
or U2939 (N_2939,N_2561,N_2638);
or U2940 (N_2940,N_2531,N_2642);
nor U2941 (N_2941,N_2680,N_2686);
and U2942 (N_2942,N_2526,N_2599);
and U2943 (N_2943,N_2585,N_2545);
or U2944 (N_2944,N_2705,N_2740);
and U2945 (N_2945,N_2538,N_2693);
and U2946 (N_2946,N_2606,N_2541);
nor U2947 (N_2947,N_2568,N_2530);
nor U2948 (N_2948,N_2590,N_2514);
and U2949 (N_2949,N_2545,N_2562);
and U2950 (N_2950,N_2746,N_2735);
and U2951 (N_2951,N_2556,N_2689);
nor U2952 (N_2952,N_2524,N_2547);
nor U2953 (N_2953,N_2500,N_2641);
or U2954 (N_2954,N_2581,N_2737);
or U2955 (N_2955,N_2656,N_2686);
nand U2956 (N_2956,N_2640,N_2685);
and U2957 (N_2957,N_2602,N_2530);
nor U2958 (N_2958,N_2525,N_2557);
nor U2959 (N_2959,N_2541,N_2586);
nor U2960 (N_2960,N_2643,N_2660);
and U2961 (N_2961,N_2530,N_2626);
nor U2962 (N_2962,N_2589,N_2602);
nand U2963 (N_2963,N_2668,N_2679);
and U2964 (N_2964,N_2661,N_2741);
nor U2965 (N_2965,N_2711,N_2639);
nor U2966 (N_2966,N_2660,N_2728);
and U2967 (N_2967,N_2745,N_2503);
and U2968 (N_2968,N_2692,N_2727);
nand U2969 (N_2969,N_2747,N_2697);
and U2970 (N_2970,N_2668,N_2604);
nand U2971 (N_2971,N_2631,N_2658);
or U2972 (N_2972,N_2687,N_2518);
nor U2973 (N_2973,N_2586,N_2540);
or U2974 (N_2974,N_2744,N_2589);
or U2975 (N_2975,N_2648,N_2596);
and U2976 (N_2976,N_2566,N_2518);
nand U2977 (N_2977,N_2510,N_2535);
nand U2978 (N_2978,N_2653,N_2671);
nor U2979 (N_2979,N_2558,N_2648);
nand U2980 (N_2980,N_2730,N_2573);
and U2981 (N_2981,N_2595,N_2513);
nor U2982 (N_2982,N_2701,N_2625);
nand U2983 (N_2983,N_2678,N_2740);
and U2984 (N_2984,N_2546,N_2660);
nor U2985 (N_2985,N_2605,N_2580);
or U2986 (N_2986,N_2540,N_2554);
and U2987 (N_2987,N_2630,N_2711);
and U2988 (N_2988,N_2675,N_2740);
and U2989 (N_2989,N_2632,N_2633);
nor U2990 (N_2990,N_2695,N_2730);
and U2991 (N_2991,N_2501,N_2553);
or U2992 (N_2992,N_2706,N_2745);
and U2993 (N_2993,N_2548,N_2519);
or U2994 (N_2994,N_2561,N_2720);
nor U2995 (N_2995,N_2661,N_2528);
nand U2996 (N_2996,N_2592,N_2583);
and U2997 (N_2997,N_2605,N_2557);
nor U2998 (N_2998,N_2703,N_2659);
and U2999 (N_2999,N_2573,N_2701);
nor U3000 (N_3000,N_2867,N_2896);
nand U3001 (N_3001,N_2917,N_2970);
or U3002 (N_3002,N_2959,N_2990);
nand U3003 (N_3003,N_2761,N_2980);
or U3004 (N_3004,N_2784,N_2920);
nor U3005 (N_3005,N_2799,N_2885);
nand U3006 (N_3006,N_2822,N_2928);
nor U3007 (N_3007,N_2847,N_2931);
nor U3008 (N_3008,N_2901,N_2986);
nor U3009 (N_3009,N_2856,N_2786);
or U3010 (N_3010,N_2989,N_2825);
nand U3011 (N_3011,N_2956,N_2946);
or U3012 (N_3012,N_2880,N_2902);
and U3013 (N_3013,N_2978,N_2987);
and U3014 (N_3014,N_2783,N_2942);
and U3015 (N_3015,N_2889,N_2813);
nor U3016 (N_3016,N_2823,N_2875);
and U3017 (N_3017,N_2776,N_2953);
and U3018 (N_3018,N_2933,N_2979);
nand U3019 (N_3019,N_2963,N_2895);
and U3020 (N_3020,N_2801,N_2996);
and U3021 (N_3021,N_2992,N_2750);
or U3022 (N_3022,N_2891,N_2983);
nand U3023 (N_3023,N_2982,N_2976);
nor U3024 (N_3024,N_2914,N_2893);
and U3025 (N_3025,N_2812,N_2924);
nand U3026 (N_3026,N_2887,N_2851);
nand U3027 (N_3027,N_2998,N_2961);
nand U3028 (N_3028,N_2929,N_2829);
nor U3029 (N_3029,N_2997,N_2897);
and U3030 (N_3030,N_2848,N_2854);
nand U3031 (N_3031,N_2894,N_2771);
nand U3032 (N_3032,N_2918,N_2862);
nor U3033 (N_3033,N_2973,N_2780);
nor U3034 (N_3034,N_2947,N_2820);
or U3035 (N_3035,N_2949,N_2888);
nand U3036 (N_3036,N_2962,N_2922);
and U3037 (N_3037,N_2912,N_2814);
or U3038 (N_3038,N_2964,N_2951);
and U3039 (N_3039,N_2850,N_2868);
or U3040 (N_3040,N_2752,N_2878);
nand U3041 (N_3041,N_2826,N_2935);
nand U3042 (N_3042,N_2940,N_2797);
and U3043 (N_3043,N_2808,N_2919);
or U3044 (N_3044,N_2795,N_2916);
and U3045 (N_3045,N_2960,N_2939);
nor U3046 (N_3046,N_2802,N_2806);
or U3047 (N_3047,N_2882,N_2807);
or U3048 (N_3048,N_2762,N_2775);
or U3049 (N_3049,N_2787,N_2796);
and U3050 (N_3050,N_2846,N_2866);
and U3051 (N_3051,N_2890,N_2824);
nand U3052 (N_3052,N_2793,N_2899);
nor U3053 (N_3053,N_2810,N_2753);
nand U3054 (N_3054,N_2852,N_2816);
nor U3055 (N_3055,N_2871,N_2781);
nand U3056 (N_3056,N_2991,N_2981);
or U3057 (N_3057,N_2835,N_2766);
xnor U3058 (N_3058,N_2907,N_2790);
nor U3059 (N_3059,N_2758,N_2792);
or U3060 (N_3060,N_2840,N_2872);
nand U3061 (N_3061,N_2863,N_2827);
nor U3062 (N_3062,N_2849,N_2789);
nand U3063 (N_3063,N_2788,N_2772);
nor U3064 (N_3064,N_2955,N_2857);
nand U3065 (N_3065,N_2994,N_2967);
and U3066 (N_3066,N_2811,N_2845);
nor U3067 (N_3067,N_2965,N_2756);
nor U3068 (N_3068,N_2975,N_2817);
or U3069 (N_3069,N_2938,N_2774);
and U3070 (N_3070,N_2966,N_2832);
or U3071 (N_3071,N_2906,N_2937);
nor U3072 (N_3072,N_2958,N_2943);
or U3073 (N_3073,N_2974,N_2984);
and U3074 (N_3074,N_2969,N_2800);
and U3075 (N_3075,N_2833,N_2853);
nand U3076 (N_3076,N_2763,N_2841);
or U3077 (N_3077,N_2865,N_2945);
or U3078 (N_3078,N_2798,N_2768);
xnor U3079 (N_3079,N_2782,N_2873);
nor U3080 (N_3080,N_2844,N_2900);
or U3081 (N_3081,N_2886,N_2858);
nor U3082 (N_3082,N_2755,N_2954);
or U3083 (N_3083,N_2957,N_2836);
nor U3084 (N_3084,N_2769,N_2883);
nor U3085 (N_3085,N_2968,N_2831);
xor U3086 (N_3086,N_2874,N_2905);
nand U3087 (N_3087,N_2985,N_2778);
nand U3088 (N_3088,N_2877,N_2834);
or U3089 (N_3089,N_2767,N_2830);
nor U3090 (N_3090,N_2843,N_2764);
and U3091 (N_3091,N_2927,N_2870);
nor U3092 (N_3092,N_2932,N_2855);
or U3093 (N_3093,N_2842,N_2910);
nand U3094 (N_3094,N_2884,N_2930);
and U3095 (N_3095,N_2898,N_2926);
and U3096 (N_3096,N_2759,N_2803);
nor U3097 (N_3097,N_2760,N_2838);
or U3098 (N_3098,N_2915,N_2876);
and U3099 (N_3099,N_2999,N_2921);
and U3100 (N_3100,N_2821,N_2773);
nand U3101 (N_3101,N_2879,N_2864);
nand U3102 (N_3102,N_2804,N_2818);
nand U3103 (N_3103,N_2765,N_2909);
nor U3104 (N_3104,N_2977,N_2923);
and U3105 (N_3105,N_2936,N_2839);
nor U3106 (N_3106,N_2837,N_2815);
or U3107 (N_3107,N_2971,N_2881);
and U3108 (N_3108,N_2911,N_2952);
nor U3109 (N_3109,N_2785,N_2950);
nand U3110 (N_3110,N_2860,N_2757);
nand U3111 (N_3111,N_2904,N_2993);
or U3112 (N_3112,N_2794,N_2859);
and U3113 (N_3113,N_2972,N_2869);
or U3114 (N_3114,N_2770,N_2751);
and U3115 (N_3115,N_2892,N_2995);
and U3116 (N_3116,N_2925,N_2908);
nand U3117 (N_3117,N_2861,N_2791);
nor U3118 (N_3118,N_2819,N_2777);
nand U3119 (N_3119,N_2805,N_2779);
and U3120 (N_3120,N_2944,N_2988);
and U3121 (N_3121,N_2913,N_2948);
nor U3122 (N_3122,N_2828,N_2754);
or U3123 (N_3123,N_2941,N_2903);
nor U3124 (N_3124,N_2809,N_2934);
nand U3125 (N_3125,N_2977,N_2999);
or U3126 (N_3126,N_2775,N_2890);
nor U3127 (N_3127,N_2852,N_2757);
nand U3128 (N_3128,N_2970,N_2997);
or U3129 (N_3129,N_2889,N_2867);
nand U3130 (N_3130,N_2906,N_2954);
and U3131 (N_3131,N_2843,N_2888);
nor U3132 (N_3132,N_2901,N_2940);
and U3133 (N_3133,N_2791,N_2867);
and U3134 (N_3134,N_2891,N_2881);
nor U3135 (N_3135,N_2791,N_2930);
nor U3136 (N_3136,N_2860,N_2952);
and U3137 (N_3137,N_2898,N_2855);
and U3138 (N_3138,N_2936,N_2861);
or U3139 (N_3139,N_2938,N_2980);
or U3140 (N_3140,N_2978,N_2943);
nand U3141 (N_3141,N_2779,N_2961);
or U3142 (N_3142,N_2770,N_2812);
nor U3143 (N_3143,N_2791,N_2966);
nand U3144 (N_3144,N_2764,N_2880);
or U3145 (N_3145,N_2962,N_2865);
nor U3146 (N_3146,N_2796,N_2919);
or U3147 (N_3147,N_2968,N_2992);
or U3148 (N_3148,N_2777,N_2870);
or U3149 (N_3149,N_2920,N_2849);
nor U3150 (N_3150,N_2963,N_2837);
nor U3151 (N_3151,N_2848,N_2888);
and U3152 (N_3152,N_2779,N_2756);
nand U3153 (N_3153,N_2984,N_2959);
nand U3154 (N_3154,N_2912,N_2754);
nand U3155 (N_3155,N_2841,N_2830);
or U3156 (N_3156,N_2952,N_2884);
or U3157 (N_3157,N_2914,N_2944);
nor U3158 (N_3158,N_2984,N_2877);
nor U3159 (N_3159,N_2935,N_2768);
and U3160 (N_3160,N_2843,N_2813);
nor U3161 (N_3161,N_2900,N_2808);
and U3162 (N_3162,N_2885,N_2898);
and U3163 (N_3163,N_2878,N_2830);
and U3164 (N_3164,N_2819,N_2770);
and U3165 (N_3165,N_2943,N_2961);
nand U3166 (N_3166,N_2826,N_2907);
nor U3167 (N_3167,N_2937,N_2969);
nand U3168 (N_3168,N_2776,N_2932);
nor U3169 (N_3169,N_2769,N_2973);
nor U3170 (N_3170,N_2787,N_2818);
and U3171 (N_3171,N_2828,N_2870);
or U3172 (N_3172,N_2898,N_2931);
and U3173 (N_3173,N_2849,N_2817);
or U3174 (N_3174,N_2938,N_2802);
and U3175 (N_3175,N_2834,N_2995);
and U3176 (N_3176,N_2849,N_2868);
or U3177 (N_3177,N_2955,N_2875);
and U3178 (N_3178,N_2769,N_2909);
or U3179 (N_3179,N_2957,N_2872);
or U3180 (N_3180,N_2936,N_2927);
nor U3181 (N_3181,N_2832,N_2896);
or U3182 (N_3182,N_2872,N_2897);
and U3183 (N_3183,N_2822,N_2917);
and U3184 (N_3184,N_2836,N_2776);
or U3185 (N_3185,N_2924,N_2863);
nor U3186 (N_3186,N_2937,N_2820);
nor U3187 (N_3187,N_2768,N_2896);
nor U3188 (N_3188,N_2897,N_2817);
or U3189 (N_3189,N_2893,N_2822);
nand U3190 (N_3190,N_2885,N_2801);
and U3191 (N_3191,N_2928,N_2784);
nor U3192 (N_3192,N_2867,N_2890);
or U3193 (N_3193,N_2820,N_2785);
or U3194 (N_3194,N_2826,N_2857);
or U3195 (N_3195,N_2797,N_2915);
nor U3196 (N_3196,N_2975,N_2929);
nand U3197 (N_3197,N_2965,N_2917);
and U3198 (N_3198,N_2937,N_2785);
and U3199 (N_3199,N_2833,N_2760);
and U3200 (N_3200,N_2928,N_2778);
or U3201 (N_3201,N_2911,N_2852);
nand U3202 (N_3202,N_2804,N_2896);
nand U3203 (N_3203,N_2949,N_2802);
nand U3204 (N_3204,N_2930,N_2980);
or U3205 (N_3205,N_2883,N_2786);
nand U3206 (N_3206,N_2761,N_2893);
nor U3207 (N_3207,N_2897,N_2954);
and U3208 (N_3208,N_2929,N_2991);
or U3209 (N_3209,N_2885,N_2976);
nor U3210 (N_3210,N_2972,N_2755);
and U3211 (N_3211,N_2797,N_2815);
nor U3212 (N_3212,N_2832,N_2984);
nand U3213 (N_3213,N_2981,N_2885);
nor U3214 (N_3214,N_2855,N_2794);
or U3215 (N_3215,N_2847,N_2872);
and U3216 (N_3216,N_2860,N_2915);
or U3217 (N_3217,N_2869,N_2841);
or U3218 (N_3218,N_2802,N_2910);
nand U3219 (N_3219,N_2990,N_2947);
and U3220 (N_3220,N_2820,N_2968);
nor U3221 (N_3221,N_2756,N_2972);
nand U3222 (N_3222,N_2844,N_2845);
or U3223 (N_3223,N_2993,N_2986);
nand U3224 (N_3224,N_2913,N_2791);
or U3225 (N_3225,N_2959,N_2806);
nor U3226 (N_3226,N_2995,N_2792);
or U3227 (N_3227,N_2897,N_2948);
and U3228 (N_3228,N_2921,N_2787);
nand U3229 (N_3229,N_2886,N_2843);
nand U3230 (N_3230,N_2988,N_2758);
or U3231 (N_3231,N_2969,N_2761);
and U3232 (N_3232,N_2805,N_2766);
nand U3233 (N_3233,N_2839,N_2863);
and U3234 (N_3234,N_2814,N_2842);
or U3235 (N_3235,N_2969,N_2815);
nor U3236 (N_3236,N_2907,N_2836);
or U3237 (N_3237,N_2900,N_2805);
nand U3238 (N_3238,N_2972,N_2918);
or U3239 (N_3239,N_2773,N_2828);
nand U3240 (N_3240,N_2914,N_2891);
or U3241 (N_3241,N_2874,N_2940);
nor U3242 (N_3242,N_2796,N_2956);
or U3243 (N_3243,N_2790,N_2841);
nand U3244 (N_3244,N_2805,N_2812);
nand U3245 (N_3245,N_2866,N_2857);
nor U3246 (N_3246,N_2956,N_2788);
or U3247 (N_3247,N_2876,N_2813);
nor U3248 (N_3248,N_2811,N_2962);
and U3249 (N_3249,N_2816,N_2868);
nor U3250 (N_3250,N_3007,N_3231);
or U3251 (N_3251,N_3164,N_3205);
nor U3252 (N_3252,N_3131,N_3024);
nor U3253 (N_3253,N_3077,N_3213);
or U3254 (N_3254,N_3115,N_3095);
nor U3255 (N_3255,N_3038,N_3017);
and U3256 (N_3256,N_3093,N_3202);
and U3257 (N_3257,N_3244,N_3072);
nor U3258 (N_3258,N_3040,N_3178);
or U3259 (N_3259,N_3001,N_3111);
nor U3260 (N_3260,N_3041,N_3188);
nand U3261 (N_3261,N_3203,N_3224);
and U3262 (N_3262,N_3055,N_3125);
nor U3263 (N_3263,N_3218,N_3217);
nand U3264 (N_3264,N_3191,N_3216);
nand U3265 (N_3265,N_3158,N_3098);
or U3266 (N_3266,N_3239,N_3124);
or U3267 (N_3267,N_3154,N_3201);
nand U3268 (N_3268,N_3196,N_3094);
nor U3269 (N_3269,N_3019,N_3092);
and U3270 (N_3270,N_3054,N_3075);
or U3271 (N_3271,N_3233,N_3005);
and U3272 (N_3272,N_3241,N_3228);
or U3273 (N_3273,N_3086,N_3242);
or U3274 (N_3274,N_3078,N_3215);
nand U3275 (N_3275,N_3046,N_3056);
nor U3276 (N_3276,N_3129,N_3018);
and U3277 (N_3277,N_3186,N_3155);
nor U3278 (N_3278,N_3180,N_3166);
or U3279 (N_3279,N_3081,N_3004);
and U3280 (N_3280,N_3069,N_3099);
and U3281 (N_3281,N_3159,N_3084);
nand U3282 (N_3282,N_3235,N_3121);
and U3283 (N_3283,N_3130,N_3232);
and U3284 (N_3284,N_3179,N_3238);
and U3285 (N_3285,N_3057,N_3112);
nand U3286 (N_3286,N_3047,N_3199);
and U3287 (N_3287,N_3008,N_3137);
nand U3288 (N_3288,N_3144,N_3109);
or U3289 (N_3289,N_3101,N_3226);
nand U3290 (N_3290,N_3170,N_3212);
nand U3291 (N_3291,N_3010,N_3176);
nor U3292 (N_3292,N_3059,N_3100);
nand U3293 (N_3293,N_3211,N_3060);
nor U3294 (N_3294,N_3210,N_3229);
nand U3295 (N_3295,N_3066,N_3013);
nor U3296 (N_3296,N_3136,N_3135);
xor U3297 (N_3297,N_3167,N_3009);
nand U3298 (N_3298,N_3181,N_3117);
nor U3299 (N_3299,N_3068,N_3185);
nor U3300 (N_3300,N_3149,N_3134);
nor U3301 (N_3301,N_3189,N_3049);
nor U3302 (N_3302,N_3090,N_3208);
nand U3303 (N_3303,N_3160,N_3104);
or U3304 (N_3304,N_3119,N_3143);
or U3305 (N_3305,N_3048,N_3163);
nor U3306 (N_3306,N_3053,N_3067);
and U3307 (N_3307,N_3083,N_3247);
nor U3308 (N_3308,N_3114,N_3015);
nor U3309 (N_3309,N_3153,N_3165);
nand U3310 (N_3310,N_3102,N_3039);
or U3311 (N_3311,N_3120,N_3128);
nand U3312 (N_3312,N_3089,N_3036);
or U3313 (N_3313,N_3145,N_3230);
or U3314 (N_3314,N_3245,N_3044);
xnor U3315 (N_3315,N_3197,N_3157);
and U3316 (N_3316,N_3172,N_3194);
nand U3317 (N_3317,N_3022,N_3123);
nand U3318 (N_3318,N_3033,N_3193);
and U3319 (N_3319,N_3105,N_3248);
or U3320 (N_3320,N_3110,N_3195);
nand U3321 (N_3321,N_3225,N_3037);
nand U3322 (N_3322,N_3021,N_3204);
nor U3323 (N_3323,N_3070,N_3052);
nor U3324 (N_3324,N_3034,N_3209);
and U3325 (N_3325,N_3138,N_3139);
or U3326 (N_3326,N_3243,N_3107);
nor U3327 (N_3327,N_3088,N_3097);
nand U3328 (N_3328,N_3198,N_3192);
nor U3329 (N_3329,N_3071,N_3042);
nand U3330 (N_3330,N_3012,N_3026);
xor U3331 (N_3331,N_3222,N_3246);
and U3332 (N_3332,N_3237,N_3000);
and U3333 (N_3333,N_3087,N_3020);
and U3334 (N_3334,N_3062,N_3183);
or U3335 (N_3335,N_3106,N_3152);
nand U3336 (N_3336,N_3161,N_3006);
or U3337 (N_3337,N_3074,N_3169);
nor U3338 (N_3338,N_3184,N_3035);
nor U3339 (N_3339,N_3043,N_3002);
and U3340 (N_3340,N_3147,N_3063);
nand U3341 (N_3341,N_3076,N_3206);
nor U3342 (N_3342,N_3014,N_3168);
nand U3343 (N_3343,N_3142,N_3113);
or U3344 (N_3344,N_3187,N_3174);
nor U3345 (N_3345,N_3108,N_3079);
or U3346 (N_3346,N_3030,N_3171);
or U3347 (N_3347,N_3214,N_3073);
and U3348 (N_3348,N_3249,N_3223);
or U3349 (N_3349,N_3032,N_3080);
and U3350 (N_3350,N_3151,N_3029);
nand U3351 (N_3351,N_3240,N_3028);
and U3352 (N_3352,N_3175,N_3148);
and U3353 (N_3353,N_3132,N_3200);
and U3354 (N_3354,N_3126,N_3065);
and U3355 (N_3355,N_3116,N_3118);
nor U3356 (N_3356,N_3003,N_3061);
nor U3357 (N_3357,N_3085,N_3096);
or U3358 (N_3358,N_3133,N_3173);
and U3359 (N_3359,N_3190,N_3103);
or U3360 (N_3360,N_3177,N_3091);
nor U3361 (N_3361,N_3025,N_3016);
nor U3362 (N_3362,N_3140,N_3027);
and U3363 (N_3363,N_3150,N_3156);
and U3364 (N_3364,N_3234,N_3127);
nand U3365 (N_3365,N_3122,N_3236);
nor U3366 (N_3366,N_3162,N_3023);
nand U3367 (N_3367,N_3051,N_3031);
nand U3368 (N_3368,N_3045,N_3221);
and U3369 (N_3369,N_3227,N_3220);
nand U3370 (N_3370,N_3219,N_3064);
or U3371 (N_3371,N_3141,N_3182);
nand U3372 (N_3372,N_3082,N_3058);
nand U3373 (N_3373,N_3050,N_3146);
nand U3374 (N_3374,N_3011,N_3207);
nand U3375 (N_3375,N_3018,N_3020);
nor U3376 (N_3376,N_3190,N_3233);
nand U3377 (N_3377,N_3163,N_3230);
nand U3378 (N_3378,N_3183,N_3047);
and U3379 (N_3379,N_3115,N_3208);
or U3380 (N_3380,N_3206,N_3220);
or U3381 (N_3381,N_3130,N_3011);
nor U3382 (N_3382,N_3150,N_3163);
and U3383 (N_3383,N_3166,N_3020);
nand U3384 (N_3384,N_3106,N_3206);
or U3385 (N_3385,N_3043,N_3242);
nor U3386 (N_3386,N_3054,N_3153);
nor U3387 (N_3387,N_3063,N_3228);
nor U3388 (N_3388,N_3249,N_3105);
and U3389 (N_3389,N_3004,N_3063);
or U3390 (N_3390,N_3042,N_3154);
nor U3391 (N_3391,N_3154,N_3046);
and U3392 (N_3392,N_3168,N_3223);
nor U3393 (N_3393,N_3101,N_3003);
nand U3394 (N_3394,N_3129,N_3177);
and U3395 (N_3395,N_3233,N_3105);
nand U3396 (N_3396,N_3216,N_3048);
or U3397 (N_3397,N_3025,N_3080);
nand U3398 (N_3398,N_3119,N_3003);
and U3399 (N_3399,N_3236,N_3026);
nor U3400 (N_3400,N_3123,N_3246);
nor U3401 (N_3401,N_3199,N_3148);
and U3402 (N_3402,N_3226,N_3144);
and U3403 (N_3403,N_3196,N_3004);
and U3404 (N_3404,N_3061,N_3037);
and U3405 (N_3405,N_3036,N_3016);
or U3406 (N_3406,N_3202,N_3218);
and U3407 (N_3407,N_3225,N_3235);
nor U3408 (N_3408,N_3232,N_3095);
nor U3409 (N_3409,N_3068,N_3137);
nor U3410 (N_3410,N_3230,N_3220);
or U3411 (N_3411,N_3030,N_3211);
and U3412 (N_3412,N_3211,N_3122);
and U3413 (N_3413,N_3203,N_3042);
nor U3414 (N_3414,N_3176,N_3217);
nand U3415 (N_3415,N_3186,N_3152);
and U3416 (N_3416,N_3075,N_3205);
xnor U3417 (N_3417,N_3044,N_3198);
or U3418 (N_3418,N_3165,N_3054);
and U3419 (N_3419,N_3149,N_3036);
or U3420 (N_3420,N_3181,N_3039);
nor U3421 (N_3421,N_3212,N_3029);
and U3422 (N_3422,N_3219,N_3120);
nor U3423 (N_3423,N_3216,N_3120);
and U3424 (N_3424,N_3160,N_3001);
nand U3425 (N_3425,N_3083,N_3078);
or U3426 (N_3426,N_3133,N_3038);
nand U3427 (N_3427,N_3144,N_3029);
nand U3428 (N_3428,N_3089,N_3112);
nor U3429 (N_3429,N_3186,N_3008);
nor U3430 (N_3430,N_3173,N_3186);
xnor U3431 (N_3431,N_3162,N_3157);
nor U3432 (N_3432,N_3138,N_3214);
nand U3433 (N_3433,N_3055,N_3046);
nor U3434 (N_3434,N_3089,N_3022);
nor U3435 (N_3435,N_3131,N_3158);
nor U3436 (N_3436,N_3072,N_3210);
and U3437 (N_3437,N_3200,N_3082);
and U3438 (N_3438,N_3185,N_3143);
and U3439 (N_3439,N_3075,N_3062);
or U3440 (N_3440,N_3012,N_3238);
nand U3441 (N_3441,N_3019,N_3209);
nor U3442 (N_3442,N_3226,N_3008);
and U3443 (N_3443,N_3181,N_3089);
or U3444 (N_3444,N_3092,N_3016);
nor U3445 (N_3445,N_3213,N_3200);
nor U3446 (N_3446,N_3037,N_3143);
nor U3447 (N_3447,N_3153,N_3168);
nand U3448 (N_3448,N_3148,N_3084);
or U3449 (N_3449,N_3162,N_3177);
nor U3450 (N_3450,N_3172,N_3106);
or U3451 (N_3451,N_3140,N_3086);
and U3452 (N_3452,N_3163,N_3207);
nor U3453 (N_3453,N_3201,N_3117);
nor U3454 (N_3454,N_3024,N_3219);
and U3455 (N_3455,N_3205,N_3161);
and U3456 (N_3456,N_3118,N_3142);
and U3457 (N_3457,N_3110,N_3141);
nand U3458 (N_3458,N_3075,N_3233);
nand U3459 (N_3459,N_3005,N_3139);
nor U3460 (N_3460,N_3190,N_3005);
and U3461 (N_3461,N_3005,N_3125);
or U3462 (N_3462,N_3078,N_3024);
or U3463 (N_3463,N_3162,N_3087);
and U3464 (N_3464,N_3229,N_3062);
or U3465 (N_3465,N_3130,N_3218);
nand U3466 (N_3466,N_3130,N_3166);
nor U3467 (N_3467,N_3067,N_3156);
xnor U3468 (N_3468,N_3223,N_3208);
or U3469 (N_3469,N_3221,N_3177);
nor U3470 (N_3470,N_3011,N_3235);
nor U3471 (N_3471,N_3179,N_3016);
nand U3472 (N_3472,N_3114,N_3195);
nand U3473 (N_3473,N_3111,N_3000);
or U3474 (N_3474,N_3051,N_3135);
and U3475 (N_3475,N_3175,N_3242);
or U3476 (N_3476,N_3061,N_3246);
nor U3477 (N_3477,N_3223,N_3206);
and U3478 (N_3478,N_3011,N_3194);
and U3479 (N_3479,N_3145,N_3003);
nand U3480 (N_3480,N_3158,N_3195);
and U3481 (N_3481,N_3160,N_3142);
or U3482 (N_3482,N_3065,N_3014);
nand U3483 (N_3483,N_3155,N_3001);
or U3484 (N_3484,N_3248,N_3071);
nor U3485 (N_3485,N_3036,N_3020);
or U3486 (N_3486,N_3117,N_3082);
nand U3487 (N_3487,N_3145,N_3097);
nor U3488 (N_3488,N_3063,N_3093);
and U3489 (N_3489,N_3073,N_3035);
nor U3490 (N_3490,N_3243,N_3201);
or U3491 (N_3491,N_3122,N_3024);
nand U3492 (N_3492,N_3137,N_3098);
and U3493 (N_3493,N_3053,N_3012);
and U3494 (N_3494,N_3087,N_3150);
nand U3495 (N_3495,N_3118,N_3042);
nand U3496 (N_3496,N_3060,N_3089);
nor U3497 (N_3497,N_3180,N_3090);
nor U3498 (N_3498,N_3082,N_3024);
nor U3499 (N_3499,N_3154,N_3091);
nor U3500 (N_3500,N_3324,N_3356);
and U3501 (N_3501,N_3310,N_3400);
nand U3502 (N_3502,N_3452,N_3263);
or U3503 (N_3503,N_3455,N_3449);
nand U3504 (N_3504,N_3315,N_3294);
and U3505 (N_3505,N_3437,N_3375);
nand U3506 (N_3506,N_3312,N_3467);
nand U3507 (N_3507,N_3292,N_3280);
nor U3508 (N_3508,N_3451,N_3384);
nand U3509 (N_3509,N_3320,N_3394);
or U3510 (N_3510,N_3287,N_3306);
nand U3511 (N_3511,N_3440,N_3334);
and U3512 (N_3512,N_3409,N_3285);
xnor U3513 (N_3513,N_3266,N_3488);
or U3514 (N_3514,N_3460,N_3252);
or U3515 (N_3515,N_3420,N_3275);
and U3516 (N_3516,N_3344,N_3302);
or U3517 (N_3517,N_3380,N_3329);
or U3518 (N_3518,N_3381,N_3382);
nor U3519 (N_3519,N_3362,N_3260);
or U3520 (N_3520,N_3297,N_3379);
or U3521 (N_3521,N_3368,N_3256);
xnor U3522 (N_3522,N_3392,N_3354);
xnor U3523 (N_3523,N_3465,N_3357);
nor U3524 (N_3524,N_3326,N_3377);
or U3525 (N_3525,N_3401,N_3495);
nand U3526 (N_3526,N_3349,N_3339);
or U3527 (N_3527,N_3456,N_3270);
and U3528 (N_3528,N_3498,N_3333);
or U3529 (N_3529,N_3414,N_3250);
or U3530 (N_3530,N_3492,N_3459);
nor U3531 (N_3531,N_3436,N_3412);
nand U3532 (N_3532,N_3445,N_3469);
or U3533 (N_3533,N_3358,N_3262);
nand U3534 (N_3534,N_3376,N_3254);
nand U3535 (N_3535,N_3346,N_3336);
nor U3536 (N_3536,N_3341,N_3295);
nor U3537 (N_3537,N_3387,N_3353);
and U3538 (N_3538,N_3485,N_3385);
nor U3539 (N_3539,N_3276,N_3390);
or U3540 (N_3540,N_3416,N_3407);
nand U3541 (N_3541,N_3342,N_3408);
nand U3542 (N_3542,N_3421,N_3328);
nand U3543 (N_3543,N_3345,N_3423);
and U3544 (N_3544,N_3355,N_3444);
nand U3545 (N_3545,N_3337,N_3286);
nand U3546 (N_3546,N_3418,N_3251);
and U3547 (N_3547,N_3261,N_3494);
nand U3548 (N_3548,N_3417,N_3271);
or U3549 (N_3549,N_3352,N_3299);
and U3550 (N_3550,N_3428,N_3476);
nor U3551 (N_3551,N_3454,N_3330);
nor U3552 (N_3552,N_3278,N_3359);
or U3553 (N_3553,N_3325,N_3478);
xnor U3554 (N_3554,N_3473,N_3487);
nor U3555 (N_3555,N_3383,N_3338);
nand U3556 (N_3556,N_3374,N_3348);
and U3557 (N_3557,N_3396,N_3415);
or U3558 (N_3558,N_3288,N_3404);
and U3559 (N_3559,N_3433,N_3419);
nor U3560 (N_3560,N_3311,N_3483);
nand U3561 (N_3561,N_3489,N_3350);
nor U3562 (N_3562,N_3273,N_3443);
nand U3563 (N_3563,N_3486,N_3389);
xor U3564 (N_3564,N_3316,N_3448);
nand U3565 (N_3565,N_3468,N_3308);
nand U3566 (N_3566,N_3327,N_3309);
and U3567 (N_3567,N_3464,N_3411);
and U3568 (N_3568,N_3323,N_3447);
nand U3569 (N_3569,N_3291,N_3300);
and U3570 (N_3570,N_3397,N_3319);
or U3571 (N_3571,N_3474,N_3413);
or U3572 (N_3572,N_3466,N_3321);
nor U3573 (N_3573,N_3304,N_3259);
or U3574 (N_3574,N_3435,N_3430);
or U3575 (N_3575,N_3313,N_3284);
nor U3576 (N_3576,N_3391,N_3481);
nand U3577 (N_3577,N_3340,N_3386);
nor U3578 (N_3578,N_3395,N_3290);
and U3579 (N_3579,N_3264,N_3283);
nand U3580 (N_3580,N_3439,N_3277);
nand U3581 (N_3581,N_3393,N_3298);
nand U3582 (N_3582,N_3422,N_3438);
nor U3583 (N_3583,N_3429,N_3332);
and U3584 (N_3584,N_3406,N_3480);
and U3585 (N_3585,N_3446,N_3361);
nor U3586 (N_3586,N_3493,N_3462);
nor U3587 (N_3587,N_3373,N_3314);
or U3588 (N_3588,N_3365,N_3281);
and U3589 (N_3589,N_3363,N_3442);
or U3590 (N_3590,N_3399,N_3265);
or U3591 (N_3591,N_3497,N_3258);
or U3592 (N_3592,N_3491,N_3369);
nand U3593 (N_3593,N_3293,N_3424);
or U3594 (N_3594,N_3461,N_3410);
or U3595 (N_3595,N_3470,N_3335);
nand U3596 (N_3596,N_3274,N_3482);
and U3597 (N_3597,N_3269,N_3471);
and U3598 (N_3598,N_3305,N_3303);
nor U3599 (N_3599,N_3318,N_3296);
and U3600 (N_3600,N_3499,N_3272);
or U3601 (N_3601,N_3427,N_3372);
nand U3602 (N_3602,N_3351,N_3370);
nor U3603 (N_3603,N_3426,N_3367);
nor U3604 (N_3604,N_3279,N_3405);
nand U3605 (N_3605,N_3331,N_3450);
nor U3606 (N_3606,N_3484,N_3479);
nand U3607 (N_3607,N_3432,N_3398);
or U3608 (N_3608,N_3441,N_3475);
nand U3609 (N_3609,N_3253,N_3496);
nand U3610 (N_3610,N_3434,N_3402);
and U3611 (N_3611,N_3282,N_3463);
or U3612 (N_3612,N_3472,N_3490);
nand U3613 (N_3613,N_3307,N_3343);
nand U3614 (N_3614,N_3425,N_3360);
nand U3615 (N_3615,N_3347,N_3322);
nand U3616 (N_3616,N_3453,N_3431);
or U3617 (N_3617,N_3371,N_3364);
nand U3618 (N_3618,N_3289,N_3477);
nand U3619 (N_3619,N_3301,N_3257);
and U3620 (N_3620,N_3255,N_3457);
nand U3621 (N_3621,N_3267,N_3366);
or U3622 (N_3622,N_3388,N_3268);
and U3623 (N_3623,N_3378,N_3458);
nor U3624 (N_3624,N_3403,N_3317);
and U3625 (N_3625,N_3484,N_3300);
nor U3626 (N_3626,N_3449,N_3333);
nor U3627 (N_3627,N_3264,N_3438);
and U3628 (N_3628,N_3318,N_3469);
or U3629 (N_3629,N_3408,N_3384);
and U3630 (N_3630,N_3372,N_3360);
nand U3631 (N_3631,N_3282,N_3395);
nand U3632 (N_3632,N_3458,N_3354);
nand U3633 (N_3633,N_3411,N_3429);
nor U3634 (N_3634,N_3480,N_3435);
nor U3635 (N_3635,N_3494,N_3306);
nor U3636 (N_3636,N_3277,N_3342);
nand U3637 (N_3637,N_3348,N_3379);
or U3638 (N_3638,N_3357,N_3339);
nor U3639 (N_3639,N_3471,N_3343);
nand U3640 (N_3640,N_3297,N_3314);
and U3641 (N_3641,N_3420,N_3411);
and U3642 (N_3642,N_3378,N_3327);
nand U3643 (N_3643,N_3466,N_3356);
and U3644 (N_3644,N_3301,N_3281);
nand U3645 (N_3645,N_3380,N_3308);
nor U3646 (N_3646,N_3318,N_3443);
nand U3647 (N_3647,N_3375,N_3398);
or U3648 (N_3648,N_3392,N_3396);
nor U3649 (N_3649,N_3405,N_3350);
nand U3650 (N_3650,N_3274,N_3441);
nand U3651 (N_3651,N_3263,N_3418);
nor U3652 (N_3652,N_3408,N_3428);
nand U3653 (N_3653,N_3403,N_3384);
nor U3654 (N_3654,N_3281,N_3254);
and U3655 (N_3655,N_3361,N_3493);
or U3656 (N_3656,N_3412,N_3288);
nor U3657 (N_3657,N_3320,N_3466);
nor U3658 (N_3658,N_3353,N_3342);
nor U3659 (N_3659,N_3261,N_3399);
or U3660 (N_3660,N_3458,N_3365);
and U3661 (N_3661,N_3352,N_3425);
and U3662 (N_3662,N_3305,N_3450);
and U3663 (N_3663,N_3315,N_3417);
nand U3664 (N_3664,N_3421,N_3322);
and U3665 (N_3665,N_3417,N_3462);
xnor U3666 (N_3666,N_3348,N_3288);
and U3667 (N_3667,N_3298,N_3449);
nor U3668 (N_3668,N_3412,N_3419);
nor U3669 (N_3669,N_3478,N_3431);
nor U3670 (N_3670,N_3459,N_3385);
nand U3671 (N_3671,N_3282,N_3447);
nand U3672 (N_3672,N_3332,N_3284);
nor U3673 (N_3673,N_3458,N_3417);
nor U3674 (N_3674,N_3410,N_3277);
and U3675 (N_3675,N_3273,N_3302);
nand U3676 (N_3676,N_3340,N_3449);
nand U3677 (N_3677,N_3254,N_3391);
xnor U3678 (N_3678,N_3499,N_3400);
nand U3679 (N_3679,N_3320,N_3489);
or U3680 (N_3680,N_3361,N_3369);
nand U3681 (N_3681,N_3368,N_3406);
nor U3682 (N_3682,N_3482,N_3413);
or U3683 (N_3683,N_3299,N_3457);
nor U3684 (N_3684,N_3335,N_3486);
nor U3685 (N_3685,N_3278,N_3286);
and U3686 (N_3686,N_3365,N_3325);
or U3687 (N_3687,N_3376,N_3369);
and U3688 (N_3688,N_3285,N_3290);
nor U3689 (N_3689,N_3415,N_3288);
or U3690 (N_3690,N_3354,N_3341);
and U3691 (N_3691,N_3454,N_3376);
or U3692 (N_3692,N_3380,N_3429);
and U3693 (N_3693,N_3346,N_3487);
or U3694 (N_3694,N_3350,N_3494);
and U3695 (N_3695,N_3387,N_3485);
or U3696 (N_3696,N_3494,N_3317);
nor U3697 (N_3697,N_3408,N_3369);
and U3698 (N_3698,N_3413,N_3477);
or U3699 (N_3699,N_3408,N_3340);
nand U3700 (N_3700,N_3389,N_3443);
and U3701 (N_3701,N_3409,N_3273);
and U3702 (N_3702,N_3436,N_3263);
and U3703 (N_3703,N_3456,N_3271);
or U3704 (N_3704,N_3395,N_3450);
and U3705 (N_3705,N_3492,N_3345);
and U3706 (N_3706,N_3306,N_3423);
and U3707 (N_3707,N_3282,N_3394);
and U3708 (N_3708,N_3442,N_3423);
and U3709 (N_3709,N_3287,N_3298);
nand U3710 (N_3710,N_3297,N_3437);
nor U3711 (N_3711,N_3277,N_3395);
or U3712 (N_3712,N_3321,N_3440);
and U3713 (N_3713,N_3345,N_3270);
nor U3714 (N_3714,N_3439,N_3479);
nand U3715 (N_3715,N_3476,N_3266);
or U3716 (N_3716,N_3291,N_3450);
and U3717 (N_3717,N_3418,N_3327);
and U3718 (N_3718,N_3306,N_3257);
and U3719 (N_3719,N_3386,N_3270);
and U3720 (N_3720,N_3433,N_3412);
nor U3721 (N_3721,N_3387,N_3252);
nand U3722 (N_3722,N_3272,N_3495);
or U3723 (N_3723,N_3486,N_3498);
or U3724 (N_3724,N_3338,N_3452);
nand U3725 (N_3725,N_3302,N_3259);
and U3726 (N_3726,N_3428,N_3378);
or U3727 (N_3727,N_3313,N_3479);
nand U3728 (N_3728,N_3256,N_3273);
nor U3729 (N_3729,N_3382,N_3256);
or U3730 (N_3730,N_3320,N_3462);
and U3731 (N_3731,N_3253,N_3479);
nor U3732 (N_3732,N_3315,N_3277);
and U3733 (N_3733,N_3484,N_3454);
nor U3734 (N_3734,N_3309,N_3292);
nand U3735 (N_3735,N_3295,N_3272);
and U3736 (N_3736,N_3495,N_3261);
nor U3737 (N_3737,N_3385,N_3444);
or U3738 (N_3738,N_3367,N_3460);
nor U3739 (N_3739,N_3465,N_3388);
or U3740 (N_3740,N_3402,N_3310);
and U3741 (N_3741,N_3386,N_3384);
nand U3742 (N_3742,N_3452,N_3417);
nor U3743 (N_3743,N_3458,N_3471);
nor U3744 (N_3744,N_3375,N_3433);
nor U3745 (N_3745,N_3299,N_3368);
nand U3746 (N_3746,N_3364,N_3458);
or U3747 (N_3747,N_3261,N_3306);
nand U3748 (N_3748,N_3403,N_3341);
or U3749 (N_3749,N_3384,N_3374);
and U3750 (N_3750,N_3524,N_3520);
nand U3751 (N_3751,N_3528,N_3608);
nand U3752 (N_3752,N_3582,N_3589);
nand U3753 (N_3753,N_3707,N_3683);
nand U3754 (N_3754,N_3607,N_3747);
nand U3755 (N_3755,N_3651,N_3501);
nand U3756 (N_3756,N_3731,N_3543);
or U3757 (N_3757,N_3511,N_3685);
and U3758 (N_3758,N_3612,N_3690);
nand U3759 (N_3759,N_3661,N_3515);
and U3760 (N_3760,N_3539,N_3689);
nand U3761 (N_3761,N_3579,N_3548);
nor U3762 (N_3762,N_3638,N_3505);
or U3763 (N_3763,N_3565,N_3654);
and U3764 (N_3764,N_3704,N_3597);
nand U3765 (N_3765,N_3615,N_3713);
nand U3766 (N_3766,N_3610,N_3706);
or U3767 (N_3767,N_3547,N_3513);
nor U3768 (N_3768,N_3581,N_3556);
and U3769 (N_3769,N_3744,N_3641);
nand U3770 (N_3770,N_3561,N_3652);
and U3771 (N_3771,N_3630,N_3534);
and U3772 (N_3772,N_3600,N_3709);
and U3773 (N_3773,N_3507,N_3682);
nor U3774 (N_3774,N_3700,N_3719);
nor U3775 (N_3775,N_3724,N_3592);
and U3776 (N_3776,N_3650,N_3602);
nand U3777 (N_3777,N_3558,N_3523);
nor U3778 (N_3778,N_3504,N_3732);
nor U3779 (N_3779,N_3519,N_3563);
and U3780 (N_3780,N_3536,N_3730);
and U3781 (N_3781,N_3710,N_3684);
nor U3782 (N_3782,N_3551,N_3681);
and U3783 (N_3783,N_3555,N_3629);
and U3784 (N_3784,N_3532,N_3691);
nand U3785 (N_3785,N_3673,N_3699);
nor U3786 (N_3786,N_3668,N_3670);
and U3787 (N_3787,N_3735,N_3535);
nand U3788 (N_3788,N_3745,N_3617);
and U3789 (N_3789,N_3727,N_3571);
and U3790 (N_3790,N_3695,N_3632);
nor U3791 (N_3791,N_3593,N_3575);
and U3792 (N_3792,N_3733,N_3711);
or U3793 (N_3793,N_3687,N_3531);
or U3794 (N_3794,N_3648,N_3663);
nand U3795 (N_3795,N_3741,N_3658);
and U3796 (N_3796,N_3669,N_3509);
or U3797 (N_3797,N_3503,N_3739);
or U3798 (N_3798,N_3569,N_3559);
and U3799 (N_3799,N_3621,N_3742);
nand U3800 (N_3800,N_3637,N_3693);
or U3801 (N_3801,N_3667,N_3737);
and U3802 (N_3802,N_3740,N_3743);
nor U3803 (N_3803,N_3508,N_3665);
nand U3804 (N_3804,N_3553,N_3725);
nand U3805 (N_3805,N_3672,N_3573);
nor U3806 (N_3806,N_3609,N_3595);
nand U3807 (N_3807,N_3526,N_3623);
nor U3808 (N_3808,N_3676,N_3738);
nand U3809 (N_3809,N_3686,N_3678);
nor U3810 (N_3810,N_3562,N_3568);
nor U3811 (N_3811,N_3620,N_3702);
or U3812 (N_3812,N_3588,N_3675);
or U3813 (N_3813,N_3643,N_3622);
nor U3814 (N_3814,N_3703,N_3572);
or U3815 (N_3815,N_3574,N_3655);
nand U3816 (N_3816,N_3604,N_3577);
nor U3817 (N_3817,N_3522,N_3598);
or U3818 (N_3818,N_3510,N_3586);
and U3819 (N_3819,N_3611,N_3549);
or U3820 (N_3820,N_3715,N_3560);
or U3821 (N_3821,N_3587,N_3530);
nand U3822 (N_3822,N_3712,N_3506);
or U3823 (N_3823,N_3514,N_3613);
nand U3824 (N_3824,N_3601,N_3723);
nand U3825 (N_3825,N_3606,N_3627);
and U3826 (N_3826,N_3746,N_3599);
nand U3827 (N_3827,N_3578,N_3545);
or U3828 (N_3828,N_3500,N_3720);
nor U3829 (N_3829,N_3636,N_3583);
and U3830 (N_3830,N_3729,N_3640);
and U3831 (N_3831,N_3647,N_3546);
nand U3832 (N_3832,N_3674,N_3517);
or U3833 (N_3833,N_3584,N_3542);
and U3834 (N_3834,N_3540,N_3619);
or U3835 (N_3835,N_3516,N_3525);
nand U3836 (N_3836,N_3557,N_3644);
nand U3837 (N_3837,N_3585,N_3596);
nand U3838 (N_3838,N_3614,N_3576);
nor U3839 (N_3839,N_3659,N_3679);
nor U3840 (N_3840,N_3697,N_3716);
nand U3841 (N_3841,N_3554,N_3564);
and U3842 (N_3842,N_3749,N_3634);
and U3843 (N_3843,N_3656,N_3580);
and U3844 (N_3844,N_3705,N_3718);
and U3845 (N_3845,N_3714,N_3544);
or U3846 (N_3846,N_3657,N_3631);
nor U3847 (N_3847,N_3521,N_3728);
and U3848 (N_3848,N_3618,N_3533);
and U3849 (N_3849,N_3502,N_3701);
or U3850 (N_3850,N_3694,N_3527);
or U3851 (N_3851,N_3570,N_3590);
or U3852 (N_3852,N_3698,N_3734);
nand U3853 (N_3853,N_3717,N_3529);
or U3854 (N_3854,N_3639,N_3653);
and U3855 (N_3855,N_3624,N_3594);
or U3856 (N_3856,N_3566,N_3645);
or U3857 (N_3857,N_3537,N_3722);
nor U3858 (N_3858,N_3518,N_3708);
nor U3859 (N_3859,N_3541,N_3626);
and U3860 (N_3860,N_3616,N_3748);
and U3861 (N_3861,N_3538,N_3603);
and U3862 (N_3862,N_3677,N_3666);
nor U3863 (N_3863,N_3660,N_3662);
or U3864 (N_3864,N_3664,N_3605);
nand U3865 (N_3865,N_3649,N_3625);
xnor U3866 (N_3866,N_3696,N_3628);
and U3867 (N_3867,N_3567,N_3671);
nor U3868 (N_3868,N_3680,N_3646);
nand U3869 (N_3869,N_3550,N_3591);
nand U3870 (N_3870,N_3726,N_3688);
and U3871 (N_3871,N_3635,N_3692);
or U3872 (N_3872,N_3633,N_3721);
nand U3873 (N_3873,N_3642,N_3552);
and U3874 (N_3874,N_3736,N_3512);
or U3875 (N_3875,N_3564,N_3706);
or U3876 (N_3876,N_3548,N_3748);
nand U3877 (N_3877,N_3663,N_3519);
and U3878 (N_3878,N_3544,N_3576);
nor U3879 (N_3879,N_3537,N_3532);
nand U3880 (N_3880,N_3573,N_3631);
or U3881 (N_3881,N_3638,N_3535);
or U3882 (N_3882,N_3611,N_3675);
xor U3883 (N_3883,N_3736,N_3633);
nand U3884 (N_3884,N_3535,N_3740);
and U3885 (N_3885,N_3733,N_3727);
nor U3886 (N_3886,N_3688,N_3535);
or U3887 (N_3887,N_3635,N_3727);
and U3888 (N_3888,N_3544,N_3615);
nor U3889 (N_3889,N_3574,N_3570);
nor U3890 (N_3890,N_3630,N_3675);
or U3891 (N_3891,N_3565,N_3739);
xor U3892 (N_3892,N_3604,N_3590);
nand U3893 (N_3893,N_3745,N_3622);
and U3894 (N_3894,N_3728,N_3536);
or U3895 (N_3895,N_3683,N_3513);
nor U3896 (N_3896,N_3721,N_3584);
nand U3897 (N_3897,N_3519,N_3540);
nor U3898 (N_3898,N_3521,N_3671);
nor U3899 (N_3899,N_3684,N_3687);
or U3900 (N_3900,N_3568,N_3579);
and U3901 (N_3901,N_3507,N_3655);
nor U3902 (N_3902,N_3588,N_3566);
or U3903 (N_3903,N_3604,N_3515);
or U3904 (N_3904,N_3531,N_3583);
or U3905 (N_3905,N_3529,N_3595);
and U3906 (N_3906,N_3562,N_3565);
nand U3907 (N_3907,N_3615,N_3654);
or U3908 (N_3908,N_3632,N_3539);
or U3909 (N_3909,N_3565,N_3678);
nor U3910 (N_3910,N_3684,N_3624);
and U3911 (N_3911,N_3648,N_3619);
nor U3912 (N_3912,N_3562,N_3567);
nor U3913 (N_3913,N_3746,N_3667);
nor U3914 (N_3914,N_3521,N_3683);
and U3915 (N_3915,N_3628,N_3542);
nor U3916 (N_3916,N_3572,N_3630);
nor U3917 (N_3917,N_3564,N_3619);
nor U3918 (N_3918,N_3706,N_3606);
nor U3919 (N_3919,N_3541,N_3689);
nand U3920 (N_3920,N_3506,N_3695);
or U3921 (N_3921,N_3570,N_3533);
or U3922 (N_3922,N_3690,N_3502);
or U3923 (N_3923,N_3509,N_3501);
and U3924 (N_3924,N_3641,N_3726);
and U3925 (N_3925,N_3683,N_3700);
nand U3926 (N_3926,N_3557,N_3677);
nor U3927 (N_3927,N_3513,N_3662);
or U3928 (N_3928,N_3623,N_3632);
and U3929 (N_3929,N_3719,N_3697);
or U3930 (N_3930,N_3715,N_3702);
nor U3931 (N_3931,N_3622,N_3532);
and U3932 (N_3932,N_3693,N_3727);
and U3933 (N_3933,N_3587,N_3706);
nand U3934 (N_3934,N_3529,N_3657);
nand U3935 (N_3935,N_3718,N_3545);
or U3936 (N_3936,N_3736,N_3725);
nand U3937 (N_3937,N_3618,N_3702);
or U3938 (N_3938,N_3539,N_3600);
or U3939 (N_3939,N_3581,N_3543);
nand U3940 (N_3940,N_3508,N_3587);
and U3941 (N_3941,N_3593,N_3530);
nand U3942 (N_3942,N_3749,N_3547);
and U3943 (N_3943,N_3606,N_3684);
nand U3944 (N_3944,N_3551,N_3549);
and U3945 (N_3945,N_3621,N_3666);
nor U3946 (N_3946,N_3508,N_3628);
and U3947 (N_3947,N_3734,N_3554);
and U3948 (N_3948,N_3705,N_3749);
and U3949 (N_3949,N_3686,N_3503);
and U3950 (N_3950,N_3634,N_3519);
xnor U3951 (N_3951,N_3557,N_3692);
and U3952 (N_3952,N_3706,N_3714);
and U3953 (N_3953,N_3503,N_3703);
or U3954 (N_3954,N_3526,N_3592);
nand U3955 (N_3955,N_3622,N_3503);
or U3956 (N_3956,N_3615,N_3580);
nand U3957 (N_3957,N_3540,N_3534);
nor U3958 (N_3958,N_3505,N_3718);
or U3959 (N_3959,N_3619,N_3598);
or U3960 (N_3960,N_3547,N_3739);
and U3961 (N_3961,N_3688,N_3618);
nor U3962 (N_3962,N_3540,N_3672);
or U3963 (N_3963,N_3682,N_3630);
and U3964 (N_3964,N_3516,N_3565);
nor U3965 (N_3965,N_3575,N_3588);
nor U3966 (N_3966,N_3619,N_3717);
nand U3967 (N_3967,N_3678,N_3659);
or U3968 (N_3968,N_3729,N_3732);
and U3969 (N_3969,N_3695,N_3604);
and U3970 (N_3970,N_3587,N_3658);
nand U3971 (N_3971,N_3747,N_3589);
nor U3972 (N_3972,N_3714,N_3527);
or U3973 (N_3973,N_3528,N_3638);
nor U3974 (N_3974,N_3591,N_3689);
and U3975 (N_3975,N_3598,N_3672);
and U3976 (N_3976,N_3720,N_3555);
nor U3977 (N_3977,N_3521,N_3662);
or U3978 (N_3978,N_3741,N_3558);
and U3979 (N_3979,N_3625,N_3688);
or U3980 (N_3980,N_3501,N_3609);
nand U3981 (N_3981,N_3658,N_3699);
nor U3982 (N_3982,N_3628,N_3582);
nor U3983 (N_3983,N_3538,N_3703);
nand U3984 (N_3984,N_3713,N_3574);
nand U3985 (N_3985,N_3544,N_3636);
nand U3986 (N_3986,N_3652,N_3704);
or U3987 (N_3987,N_3710,N_3746);
or U3988 (N_3988,N_3623,N_3667);
xnor U3989 (N_3989,N_3586,N_3626);
nand U3990 (N_3990,N_3500,N_3608);
or U3991 (N_3991,N_3699,N_3628);
nor U3992 (N_3992,N_3637,N_3509);
or U3993 (N_3993,N_3704,N_3627);
or U3994 (N_3994,N_3597,N_3525);
or U3995 (N_3995,N_3699,N_3501);
nor U3996 (N_3996,N_3647,N_3687);
nand U3997 (N_3997,N_3613,N_3623);
or U3998 (N_3998,N_3658,N_3516);
nand U3999 (N_3999,N_3583,N_3682);
nor U4000 (N_4000,N_3771,N_3994);
nand U4001 (N_4001,N_3842,N_3997);
nand U4002 (N_4002,N_3859,N_3815);
nor U4003 (N_4003,N_3896,N_3784);
or U4004 (N_4004,N_3828,N_3750);
nand U4005 (N_4005,N_3865,N_3811);
xor U4006 (N_4006,N_3786,N_3819);
nor U4007 (N_4007,N_3777,N_3809);
and U4008 (N_4008,N_3803,N_3947);
and U4009 (N_4009,N_3894,N_3810);
and U4010 (N_4010,N_3876,N_3933);
nand U4011 (N_4011,N_3831,N_3808);
nand U4012 (N_4012,N_3818,N_3775);
or U4013 (N_4013,N_3821,N_3832);
nor U4014 (N_4014,N_3954,N_3908);
nand U4015 (N_4015,N_3812,N_3879);
and U4016 (N_4016,N_3797,N_3758);
and U4017 (N_4017,N_3878,N_3982);
nand U4018 (N_4018,N_3972,N_3945);
nor U4019 (N_4019,N_3943,N_3891);
and U4020 (N_4020,N_3970,N_3907);
or U4021 (N_4021,N_3886,N_3989);
nor U4022 (N_4022,N_3754,N_3902);
or U4023 (N_4023,N_3914,N_3930);
nand U4024 (N_4024,N_3778,N_3986);
nor U4025 (N_4025,N_3849,N_3981);
or U4026 (N_4026,N_3835,N_3780);
nand U4027 (N_4027,N_3976,N_3900);
and U4028 (N_4028,N_3925,N_3800);
and U4029 (N_4029,N_3949,N_3985);
xor U4030 (N_4030,N_3848,N_3841);
or U4031 (N_4031,N_3927,N_3998);
and U4032 (N_4032,N_3922,N_3988);
and U4033 (N_4033,N_3816,N_3763);
or U4034 (N_4034,N_3873,N_3843);
or U4035 (N_4035,N_3974,N_3958);
nor U4036 (N_4036,N_3804,N_3862);
nor U4037 (N_4037,N_3942,N_3991);
or U4038 (N_4038,N_3875,N_3906);
and U4039 (N_4039,N_3971,N_3996);
or U4040 (N_4040,N_3904,N_3987);
nor U4041 (N_4041,N_3992,N_3756);
nor U4042 (N_4042,N_3921,N_3926);
nor U4043 (N_4043,N_3788,N_3946);
and U4044 (N_4044,N_3980,N_3774);
nor U4045 (N_4045,N_3846,N_3779);
and U4046 (N_4046,N_3871,N_3787);
nand U4047 (N_4047,N_3755,N_3990);
or U4048 (N_4048,N_3884,N_3975);
nor U4049 (N_4049,N_3913,N_3941);
and U4050 (N_4050,N_3888,N_3932);
and U4051 (N_4051,N_3833,N_3957);
nand U4052 (N_4052,N_3937,N_3850);
nand U4053 (N_4053,N_3966,N_3887);
and U4054 (N_4054,N_3805,N_3924);
nor U4055 (N_4055,N_3752,N_3798);
nor U4056 (N_4056,N_3920,N_3829);
nand U4057 (N_4057,N_3911,N_3825);
or U4058 (N_4058,N_3993,N_3885);
nand U4059 (N_4059,N_3951,N_3918);
nor U4060 (N_4060,N_3844,N_3934);
nor U4061 (N_4061,N_3881,N_3965);
nand U4062 (N_4062,N_3867,N_3897);
nor U4063 (N_4063,N_3765,N_3802);
and U4064 (N_4064,N_3869,N_3963);
or U4065 (N_4065,N_3751,N_3772);
and U4066 (N_4066,N_3753,N_3880);
nand U4067 (N_4067,N_3764,N_3785);
nand U4068 (N_4068,N_3762,N_3757);
nand U4069 (N_4069,N_3955,N_3905);
nor U4070 (N_4070,N_3961,N_3826);
nand U4071 (N_4071,N_3768,N_3845);
nand U4072 (N_4072,N_3817,N_3890);
nor U4073 (N_4073,N_3834,N_3983);
and U4074 (N_4074,N_3767,N_3915);
and U4075 (N_4075,N_3794,N_3814);
and U4076 (N_4076,N_3919,N_3795);
or U4077 (N_4077,N_3909,N_3766);
and U4078 (N_4078,N_3916,N_3889);
or U4079 (N_4079,N_3944,N_3882);
or U4080 (N_4080,N_3855,N_3759);
nand U4081 (N_4081,N_3968,N_3813);
nor U4082 (N_4082,N_3903,N_3877);
and U4083 (N_4083,N_3979,N_3860);
or U4084 (N_4084,N_3861,N_3910);
and U4085 (N_4085,N_3928,N_3858);
nand U4086 (N_4086,N_3852,N_3984);
nor U4087 (N_4087,N_3801,N_3929);
nor U4088 (N_4088,N_3962,N_3854);
and U4089 (N_4089,N_3870,N_3792);
nand U4090 (N_4090,N_3838,N_3964);
nor U4091 (N_4091,N_3769,N_3953);
nand U4092 (N_4092,N_3836,N_3868);
and U4093 (N_4093,N_3847,N_3807);
nor U4094 (N_4094,N_3901,N_3893);
or U4095 (N_4095,N_3995,N_3864);
nor U4096 (N_4096,N_3857,N_3969);
and U4097 (N_4097,N_3761,N_3782);
nor U4098 (N_4098,N_3820,N_3760);
xor U4099 (N_4099,N_3960,N_3823);
and U4100 (N_4100,N_3899,N_3977);
nor U4101 (N_4101,N_3863,N_3898);
nand U4102 (N_4102,N_3776,N_3892);
xnor U4103 (N_4103,N_3912,N_3790);
nor U4104 (N_4104,N_3791,N_3789);
and U4105 (N_4105,N_3883,N_3895);
nand U4106 (N_4106,N_3866,N_3781);
nand U4107 (N_4107,N_3799,N_3999);
nand U4108 (N_4108,N_3967,N_3840);
and U4109 (N_4109,N_3936,N_3872);
and U4110 (N_4110,N_3956,N_3938);
nand U4111 (N_4111,N_3830,N_3856);
nor U4112 (N_4112,N_3806,N_3952);
nand U4113 (N_4113,N_3917,N_3822);
or U4114 (N_4114,N_3793,N_3839);
nor U4115 (N_4115,N_3837,N_3939);
nor U4116 (N_4116,N_3874,N_3851);
nand U4117 (N_4117,N_3770,N_3853);
nor U4118 (N_4118,N_3796,N_3783);
or U4119 (N_4119,N_3827,N_3978);
or U4120 (N_4120,N_3950,N_3940);
and U4121 (N_4121,N_3931,N_3923);
and U4122 (N_4122,N_3948,N_3935);
nor U4123 (N_4123,N_3773,N_3973);
nor U4124 (N_4124,N_3824,N_3959);
or U4125 (N_4125,N_3789,N_3981);
or U4126 (N_4126,N_3909,N_3927);
nor U4127 (N_4127,N_3824,N_3853);
and U4128 (N_4128,N_3828,N_3753);
and U4129 (N_4129,N_3807,N_3844);
or U4130 (N_4130,N_3779,N_3760);
nand U4131 (N_4131,N_3777,N_3914);
nor U4132 (N_4132,N_3844,N_3955);
nor U4133 (N_4133,N_3926,N_3993);
or U4134 (N_4134,N_3932,N_3848);
xnor U4135 (N_4135,N_3826,N_3780);
or U4136 (N_4136,N_3895,N_3892);
and U4137 (N_4137,N_3983,N_3857);
nor U4138 (N_4138,N_3809,N_3750);
xor U4139 (N_4139,N_3990,N_3792);
or U4140 (N_4140,N_3824,N_3860);
nand U4141 (N_4141,N_3989,N_3894);
nor U4142 (N_4142,N_3987,N_3968);
nor U4143 (N_4143,N_3872,N_3783);
nor U4144 (N_4144,N_3857,N_3824);
nor U4145 (N_4145,N_3961,N_3780);
or U4146 (N_4146,N_3842,N_3793);
nand U4147 (N_4147,N_3986,N_3751);
or U4148 (N_4148,N_3805,N_3984);
nand U4149 (N_4149,N_3967,N_3917);
nand U4150 (N_4150,N_3984,N_3985);
nor U4151 (N_4151,N_3790,N_3787);
or U4152 (N_4152,N_3858,N_3943);
and U4153 (N_4153,N_3895,N_3884);
nor U4154 (N_4154,N_3931,N_3995);
and U4155 (N_4155,N_3793,N_3919);
nand U4156 (N_4156,N_3853,N_3920);
nor U4157 (N_4157,N_3971,N_3793);
nor U4158 (N_4158,N_3796,N_3954);
nand U4159 (N_4159,N_3865,N_3922);
nand U4160 (N_4160,N_3913,N_3794);
nor U4161 (N_4161,N_3815,N_3756);
nor U4162 (N_4162,N_3903,N_3989);
and U4163 (N_4163,N_3812,N_3867);
or U4164 (N_4164,N_3851,N_3831);
nand U4165 (N_4165,N_3894,N_3838);
and U4166 (N_4166,N_3914,N_3980);
or U4167 (N_4167,N_3815,N_3979);
and U4168 (N_4168,N_3894,N_3831);
or U4169 (N_4169,N_3752,N_3940);
nand U4170 (N_4170,N_3847,N_3994);
nand U4171 (N_4171,N_3897,N_3873);
nand U4172 (N_4172,N_3815,N_3868);
nor U4173 (N_4173,N_3774,N_3826);
nand U4174 (N_4174,N_3790,N_3796);
nor U4175 (N_4175,N_3926,N_3879);
or U4176 (N_4176,N_3812,N_3918);
nand U4177 (N_4177,N_3894,N_3835);
nand U4178 (N_4178,N_3767,N_3914);
or U4179 (N_4179,N_3977,N_3771);
xor U4180 (N_4180,N_3891,N_3867);
or U4181 (N_4181,N_3855,N_3778);
or U4182 (N_4182,N_3863,N_3848);
nor U4183 (N_4183,N_3900,N_3790);
and U4184 (N_4184,N_3772,N_3915);
and U4185 (N_4185,N_3751,N_3981);
and U4186 (N_4186,N_3963,N_3823);
or U4187 (N_4187,N_3758,N_3922);
or U4188 (N_4188,N_3919,N_3938);
nor U4189 (N_4189,N_3839,N_3928);
or U4190 (N_4190,N_3837,N_3992);
and U4191 (N_4191,N_3877,N_3979);
nand U4192 (N_4192,N_3808,N_3829);
nand U4193 (N_4193,N_3885,N_3920);
and U4194 (N_4194,N_3845,N_3801);
or U4195 (N_4195,N_3952,N_3902);
nand U4196 (N_4196,N_3888,N_3957);
or U4197 (N_4197,N_3808,N_3816);
and U4198 (N_4198,N_3752,N_3967);
or U4199 (N_4199,N_3794,N_3795);
nand U4200 (N_4200,N_3753,N_3921);
and U4201 (N_4201,N_3902,N_3949);
or U4202 (N_4202,N_3986,N_3777);
or U4203 (N_4203,N_3930,N_3957);
nand U4204 (N_4204,N_3981,N_3822);
or U4205 (N_4205,N_3879,N_3781);
and U4206 (N_4206,N_3783,N_3908);
nand U4207 (N_4207,N_3768,N_3854);
nor U4208 (N_4208,N_3907,N_3961);
nor U4209 (N_4209,N_3814,N_3805);
nand U4210 (N_4210,N_3776,N_3753);
and U4211 (N_4211,N_3761,N_3974);
or U4212 (N_4212,N_3774,N_3929);
nand U4213 (N_4213,N_3898,N_3751);
or U4214 (N_4214,N_3880,N_3758);
nor U4215 (N_4215,N_3980,N_3849);
or U4216 (N_4216,N_3969,N_3932);
and U4217 (N_4217,N_3757,N_3768);
or U4218 (N_4218,N_3797,N_3994);
nor U4219 (N_4219,N_3801,N_3987);
or U4220 (N_4220,N_3907,N_3750);
and U4221 (N_4221,N_3877,N_3981);
and U4222 (N_4222,N_3963,N_3771);
nand U4223 (N_4223,N_3922,N_3800);
or U4224 (N_4224,N_3799,N_3764);
nand U4225 (N_4225,N_3801,N_3995);
and U4226 (N_4226,N_3908,N_3795);
nor U4227 (N_4227,N_3964,N_3802);
and U4228 (N_4228,N_3929,N_3975);
or U4229 (N_4229,N_3862,N_3948);
or U4230 (N_4230,N_3792,N_3778);
nand U4231 (N_4231,N_3907,N_3960);
or U4232 (N_4232,N_3780,N_3767);
or U4233 (N_4233,N_3912,N_3768);
nor U4234 (N_4234,N_3824,N_3900);
nor U4235 (N_4235,N_3838,N_3813);
xor U4236 (N_4236,N_3811,N_3920);
nor U4237 (N_4237,N_3966,N_3949);
nor U4238 (N_4238,N_3753,N_3769);
and U4239 (N_4239,N_3810,N_3951);
nand U4240 (N_4240,N_3960,N_3945);
and U4241 (N_4241,N_3986,N_3876);
and U4242 (N_4242,N_3879,N_3797);
and U4243 (N_4243,N_3875,N_3980);
and U4244 (N_4244,N_3935,N_3811);
nand U4245 (N_4245,N_3828,N_3876);
or U4246 (N_4246,N_3936,N_3836);
or U4247 (N_4247,N_3815,N_3841);
nor U4248 (N_4248,N_3996,N_3909);
nand U4249 (N_4249,N_3868,N_3880);
and U4250 (N_4250,N_4064,N_4189);
nand U4251 (N_4251,N_4092,N_4192);
nand U4252 (N_4252,N_4172,N_4188);
nor U4253 (N_4253,N_4021,N_4082);
nand U4254 (N_4254,N_4066,N_4099);
nor U4255 (N_4255,N_4232,N_4184);
nand U4256 (N_4256,N_4235,N_4054);
and U4257 (N_4257,N_4069,N_4149);
nand U4258 (N_4258,N_4114,N_4233);
nand U4259 (N_4259,N_4112,N_4013);
or U4260 (N_4260,N_4131,N_4146);
and U4261 (N_4261,N_4206,N_4191);
or U4262 (N_4262,N_4180,N_4138);
and U4263 (N_4263,N_4018,N_4070);
or U4264 (N_4264,N_4036,N_4014);
nor U4265 (N_4265,N_4074,N_4088);
or U4266 (N_4266,N_4212,N_4024);
nor U4267 (N_4267,N_4150,N_4121);
nand U4268 (N_4268,N_4104,N_4110);
nor U4269 (N_4269,N_4229,N_4041);
nand U4270 (N_4270,N_4198,N_4139);
nand U4271 (N_4271,N_4011,N_4096);
nand U4272 (N_4272,N_4239,N_4230);
nor U4273 (N_4273,N_4071,N_4141);
nor U4274 (N_4274,N_4095,N_4026);
nand U4275 (N_4275,N_4111,N_4193);
or U4276 (N_4276,N_4169,N_4032);
and U4277 (N_4277,N_4063,N_4202);
and U4278 (N_4278,N_4019,N_4120);
or U4279 (N_4279,N_4058,N_4025);
or U4280 (N_4280,N_4152,N_4143);
nor U4281 (N_4281,N_4001,N_4086);
and U4282 (N_4282,N_4196,N_4009);
or U4283 (N_4283,N_4243,N_4186);
or U4284 (N_4284,N_4119,N_4240);
xor U4285 (N_4285,N_4079,N_4052);
nand U4286 (N_4286,N_4136,N_4102);
or U4287 (N_4287,N_4008,N_4106);
or U4288 (N_4288,N_4050,N_4157);
nor U4289 (N_4289,N_4047,N_4090);
nor U4290 (N_4290,N_4030,N_4137);
nand U4291 (N_4291,N_4012,N_4238);
nor U4292 (N_4292,N_4003,N_4231);
and U4293 (N_4293,N_4101,N_4133);
nor U4294 (N_4294,N_4181,N_4098);
nand U4295 (N_4295,N_4144,N_4207);
nor U4296 (N_4296,N_4051,N_4155);
nand U4297 (N_4297,N_4228,N_4075);
nor U4298 (N_4298,N_4046,N_4147);
or U4299 (N_4299,N_4222,N_4195);
nand U4300 (N_4300,N_4134,N_4241);
nor U4301 (N_4301,N_4065,N_4130);
xnor U4302 (N_4302,N_4246,N_4037);
nand U4303 (N_4303,N_4145,N_4168);
nand U4304 (N_4304,N_4045,N_4227);
or U4305 (N_4305,N_4171,N_4016);
or U4306 (N_4306,N_4034,N_4044);
nor U4307 (N_4307,N_4201,N_4108);
and U4308 (N_4308,N_4091,N_4178);
nand U4309 (N_4309,N_4062,N_4153);
nand U4310 (N_4310,N_4087,N_4127);
or U4311 (N_4311,N_4199,N_4118);
nor U4312 (N_4312,N_4126,N_4213);
nand U4313 (N_4313,N_4103,N_4078);
or U4314 (N_4314,N_4100,N_4161);
nand U4315 (N_4315,N_4190,N_4038);
nand U4316 (N_4316,N_4125,N_4226);
and U4317 (N_4317,N_4000,N_4151);
nand U4318 (N_4318,N_4060,N_4214);
nand U4319 (N_4319,N_4218,N_4164);
nor U4320 (N_4320,N_4160,N_4061);
or U4321 (N_4321,N_4217,N_4223);
or U4322 (N_4322,N_4242,N_4107);
and U4323 (N_4323,N_4200,N_4234);
and U4324 (N_4324,N_4205,N_4128);
and U4325 (N_4325,N_4057,N_4221);
xnor U4326 (N_4326,N_4084,N_4209);
and U4327 (N_4327,N_4093,N_4005);
nor U4328 (N_4328,N_4176,N_4156);
and U4329 (N_4329,N_4163,N_4165);
nand U4330 (N_4330,N_4080,N_4208);
or U4331 (N_4331,N_4173,N_4236);
and U4332 (N_4332,N_4048,N_4017);
nand U4333 (N_4333,N_4170,N_4077);
nor U4334 (N_4334,N_4006,N_4224);
nand U4335 (N_4335,N_4166,N_4097);
nand U4336 (N_4336,N_4204,N_4249);
and U4337 (N_4337,N_4022,N_4055);
and U4338 (N_4338,N_4042,N_4072);
nor U4339 (N_4339,N_4142,N_4094);
xor U4340 (N_4340,N_4117,N_4076);
and U4341 (N_4341,N_4059,N_4179);
and U4342 (N_4342,N_4073,N_4031);
nor U4343 (N_4343,N_4248,N_4068);
nor U4344 (N_4344,N_4203,N_4113);
or U4345 (N_4345,N_4245,N_4085);
nand U4346 (N_4346,N_4175,N_4028);
nor U4347 (N_4347,N_4159,N_4089);
nand U4348 (N_4348,N_4162,N_4132);
and U4349 (N_4349,N_4220,N_4004);
and U4350 (N_4350,N_4105,N_4197);
or U4351 (N_4351,N_4148,N_4115);
nand U4352 (N_4352,N_4237,N_4039);
nand U4353 (N_4353,N_4185,N_4040);
or U4354 (N_4354,N_4027,N_4081);
nand U4355 (N_4355,N_4049,N_4158);
or U4356 (N_4356,N_4194,N_4174);
nand U4357 (N_4357,N_4154,N_4029);
nand U4358 (N_4358,N_4056,N_4122);
nor U4359 (N_4359,N_4002,N_4007);
or U4360 (N_4360,N_4123,N_4010);
nor U4361 (N_4361,N_4219,N_4109);
nand U4362 (N_4362,N_4211,N_4167);
and U4363 (N_4363,N_4187,N_4033);
nor U4364 (N_4364,N_4020,N_4210);
nor U4365 (N_4365,N_4053,N_4177);
or U4366 (N_4366,N_4043,N_4023);
xor U4367 (N_4367,N_4083,N_4216);
nand U4368 (N_4368,N_4247,N_4225);
and U4369 (N_4369,N_4135,N_4116);
nor U4370 (N_4370,N_4129,N_4035);
nor U4371 (N_4371,N_4215,N_4244);
and U4372 (N_4372,N_4124,N_4140);
or U4373 (N_4373,N_4015,N_4183);
and U4374 (N_4374,N_4067,N_4182);
or U4375 (N_4375,N_4138,N_4132);
or U4376 (N_4376,N_4236,N_4158);
or U4377 (N_4377,N_4197,N_4002);
nor U4378 (N_4378,N_4239,N_4179);
nand U4379 (N_4379,N_4160,N_4086);
nand U4380 (N_4380,N_4175,N_4123);
or U4381 (N_4381,N_4047,N_4074);
and U4382 (N_4382,N_4211,N_4045);
and U4383 (N_4383,N_4228,N_4160);
or U4384 (N_4384,N_4042,N_4180);
nand U4385 (N_4385,N_4138,N_4060);
or U4386 (N_4386,N_4224,N_4223);
nor U4387 (N_4387,N_4060,N_4080);
nand U4388 (N_4388,N_4085,N_4102);
or U4389 (N_4389,N_4248,N_4192);
nor U4390 (N_4390,N_4075,N_4168);
nor U4391 (N_4391,N_4203,N_4026);
and U4392 (N_4392,N_4066,N_4129);
or U4393 (N_4393,N_4139,N_4064);
nor U4394 (N_4394,N_4211,N_4115);
or U4395 (N_4395,N_4177,N_4071);
nor U4396 (N_4396,N_4205,N_4157);
nand U4397 (N_4397,N_4028,N_4161);
nor U4398 (N_4398,N_4214,N_4207);
and U4399 (N_4399,N_4007,N_4159);
and U4400 (N_4400,N_4078,N_4030);
or U4401 (N_4401,N_4036,N_4085);
or U4402 (N_4402,N_4123,N_4073);
nand U4403 (N_4403,N_4115,N_4010);
nor U4404 (N_4404,N_4021,N_4227);
or U4405 (N_4405,N_4121,N_4032);
or U4406 (N_4406,N_4119,N_4147);
nand U4407 (N_4407,N_4025,N_4042);
nand U4408 (N_4408,N_4240,N_4141);
and U4409 (N_4409,N_4074,N_4106);
and U4410 (N_4410,N_4142,N_4009);
or U4411 (N_4411,N_4163,N_4064);
or U4412 (N_4412,N_4105,N_4219);
and U4413 (N_4413,N_4127,N_4010);
nor U4414 (N_4414,N_4032,N_4081);
nor U4415 (N_4415,N_4114,N_4134);
or U4416 (N_4416,N_4055,N_4120);
and U4417 (N_4417,N_4110,N_4165);
and U4418 (N_4418,N_4049,N_4197);
and U4419 (N_4419,N_4171,N_4219);
or U4420 (N_4420,N_4247,N_4120);
or U4421 (N_4421,N_4220,N_4202);
and U4422 (N_4422,N_4230,N_4061);
and U4423 (N_4423,N_4103,N_4187);
nor U4424 (N_4424,N_4117,N_4036);
and U4425 (N_4425,N_4077,N_4075);
and U4426 (N_4426,N_4094,N_4133);
nand U4427 (N_4427,N_4015,N_4154);
and U4428 (N_4428,N_4075,N_4060);
nand U4429 (N_4429,N_4148,N_4154);
nor U4430 (N_4430,N_4124,N_4168);
and U4431 (N_4431,N_4124,N_4008);
and U4432 (N_4432,N_4058,N_4221);
or U4433 (N_4433,N_4195,N_4215);
xnor U4434 (N_4434,N_4143,N_4163);
nand U4435 (N_4435,N_4013,N_4096);
nand U4436 (N_4436,N_4242,N_4082);
nand U4437 (N_4437,N_4020,N_4227);
nand U4438 (N_4438,N_4135,N_4118);
and U4439 (N_4439,N_4029,N_4063);
nor U4440 (N_4440,N_4217,N_4247);
nand U4441 (N_4441,N_4222,N_4074);
or U4442 (N_4442,N_4084,N_4173);
or U4443 (N_4443,N_4152,N_4177);
or U4444 (N_4444,N_4217,N_4216);
nand U4445 (N_4445,N_4096,N_4228);
nand U4446 (N_4446,N_4203,N_4209);
or U4447 (N_4447,N_4117,N_4024);
nor U4448 (N_4448,N_4041,N_4213);
and U4449 (N_4449,N_4111,N_4209);
and U4450 (N_4450,N_4148,N_4072);
or U4451 (N_4451,N_4004,N_4070);
or U4452 (N_4452,N_4082,N_4118);
nor U4453 (N_4453,N_4223,N_4116);
or U4454 (N_4454,N_4204,N_4056);
and U4455 (N_4455,N_4173,N_4213);
and U4456 (N_4456,N_4113,N_4201);
xnor U4457 (N_4457,N_4243,N_4136);
and U4458 (N_4458,N_4160,N_4089);
or U4459 (N_4459,N_4051,N_4229);
nor U4460 (N_4460,N_4103,N_4111);
and U4461 (N_4461,N_4069,N_4106);
nor U4462 (N_4462,N_4178,N_4191);
or U4463 (N_4463,N_4163,N_4248);
nor U4464 (N_4464,N_4058,N_4083);
nand U4465 (N_4465,N_4106,N_4026);
nand U4466 (N_4466,N_4026,N_4153);
and U4467 (N_4467,N_4219,N_4019);
or U4468 (N_4468,N_4087,N_4157);
or U4469 (N_4469,N_4086,N_4095);
or U4470 (N_4470,N_4085,N_4150);
or U4471 (N_4471,N_4191,N_4220);
and U4472 (N_4472,N_4135,N_4175);
nand U4473 (N_4473,N_4210,N_4150);
or U4474 (N_4474,N_4064,N_4137);
nor U4475 (N_4475,N_4208,N_4238);
or U4476 (N_4476,N_4103,N_4231);
or U4477 (N_4477,N_4051,N_4142);
or U4478 (N_4478,N_4155,N_4221);
nor U4479 (N_4479,N_4094,N_4041);
nand U4480 (N_4480,N_4033,N_4110);
and U4481 (N_4481,N_4021,N_4177);
and U4482 (N_4482,N_4007,N_4198);
and U4483 (N_4483,N_4035,N_4104);
or U4484 (N_4484,N_4036,N_4230);
or U4485 (N_4485,N_4021,N_4225);
or U4486 (N_4486,N_4208,N_4241);
or U4487 (N_4487,N_4163,N_4131);
nand U4488 (N_4488,N_4187,N_4063);
nand U4489 (N_4489,N_4085,N_4211);
and U4490 (N_4490,N_4087,N_4000);
nor U4491 (N_4491,N_4238,N_4184);
nor U4492 (N_4492,N_4211,N_4037);
or U4493 (N_4493,N_4222,N_4224);
and U4494 (N_4494,N_4129,N_4041);
and U4495 (N_4495,N_4067,N_4211);
xor U4496 (N_4496,N_4009,N_4043);
nor U4497 (N_4497,N_4125,N_4138);
nor U4498 (N_4498,N_4039,N_4049);
nand U4499 (N_4499,N_4104,N_4091);
and U4500 (N_4500,N_4327,N_4273);
and U4501 (N_4501,N_4356,N_4498);
and U4502 (N_4502,N_4276,N_4308);
and U4503 (N_4503,N_4307,N_4321);
or U4504 (N_4504,N_4298,N_4335);
and U4505 (N_4505,N_4260,N_4350);
nor U4506 (N_4506,N_4394,N_4455);
and U4507 (N_4507,N_4410,N_4277);
nor U4508 (N_4508,N_4414,N_4300);
nor U4509 (N_4509,N_4415,N_4337);
nand U4510 (N_4510,N_4467,N_4281);
and U4511 (N_4511,N_4393,N_4351);
nor U4512 (N_4512,N_4326,N_4269);
nand U4513 (N_4513,N_4427,N_4383);
and U4514 (N_4514,N_4424,N_4405);
or U4515 (N_4515,N_4359,N_4460);
or U4516 (N_4516,N_4294,N_4271);
nor U4517 (N_4517,N_4272,N_4375);
and U4518 (N_4518,N_4317,N_4340);
or U4519 (N_4519,N_4329,N_4477);
nand U4520 (N_4520,N_4322,N_4270);
or U4521 (N_4521,N_4412,N_4313);
and U4522 (N_4522,N_4345,N_4333);
and U4523 (N_4523,N_4413,N_4443);
nand U4524 (N_4524,N_4399,N_4374);
and U4525 (N_4525,N_4334,N_4433);
and U4526 (N_4526,N_4320,N_4324);
and U4527 (N_4527,N_4278,N_4325);
or U4528 (N_4528,N_4445,N_4389);
or U4529 (N_4529,N_4316,N_4417);
and U4530 (N_4530,N_4396,N_4419);
nor U4531 (N_4531,N_4435,N_4478);
or U4532 (N_4532,N_4259,N_4457);
nor U4533 (N_4533,N_4341,N_4452);
nand U4534 (N_4534,N_4296,N_4252);
nand U4535 (N_4535,N_4456,N_4441);
and U4536 (N_4536,N_4297,N_4390);
and U4537 (N_4537,N_4357,N_4288);
nor U4538 (N_4538,N_4255,N_4482);
or U4539 (N_4539,N_4499,N_4309);
nand U4540 (N_4540,N_4280,N_4409);
and U4541 (N_4541,N_4497,N_4458);
nor U4542 (N_4542,N_4440,N_4379);
nand U4543 (N_4543,N_4385,N_4423);
nor U4544 (N_4544,N_4291,N_4481);
nand U4545 (N_4545,N_4444,N_4254);
nor U4546 (N_4546,N_4484,N_4369);
or U4547 (N_4547,N_4287,N_4446);
nand U4548 (N_4548,N_4268,N_4381);
xor U4549 (N_4549,N_4261,N_4432);
xnor U4550 (N_4550,N_4373,N_4358);
nand U4551 (N_4551,N_4464,N_4302);
nor U4552 (N_4552,N_4420,N_4489);
nor U4553 (N_4553,N_4403,N_4469);
xor U4554 (N_4554,N_4480,N_4279);
nor U4555 (N_4555,N_4392,N_4263);
and U4556 (N_4556,N_4372,N_4353);
nand U4557 (N_4557,N_4476,N_4496);
nand U4558 (N_4558,N_4306,N_4395);
or U4559 (N_4559,N_4336,N_4386);
and U4560 (N_4560,N_4311,N_4343);
nor U4561 (N_4561,N_4470,N_4371);
nand U4562 (N_4562,N_4338,N_4303);
xor U4563 (N_4563,N_4366,N_4267);
nor U4564 (N_4564,N_4284,N_4293);
and U4565 (N_4565,N_4407,N_4257);
nor U4566 (N_4566,N_4400,N_4384);
nand U4567 (N_4567,N_4376,N_4436);
nor U4568 (N_4568,N_4387,N_4348);
or U4569 (N_4569,N_4434,N_4398);
nand U4570 (N_4570,N_4354,N_4439);
and U4571 (N_4571,N_4422,N_4347);
nand U4572 (N_4572,N_4483,N_4490);
or U4573 (N_4573,N_4253,N_4388);
and U4574 (N_4574,N_4342,N_4431);
nor U4575 (N_4575,N_4262,N_4323);
and U4576 (N_4576,N_4266,N_4401);
nor U4577 (N_4577,N_4305,N_4404);
or U4578 (N_4578,N_4449,N_4377);
nand U4579 (N_4579,N_4304,N_4448);
nor U4580 (N_4580,N_4318,N_4428);
or U4581 (N_4581,N_4365,N_4397);
or U4582 (N_4582,N_4461,N_4474);
and U4583 (N_4583,N_4488,N_4391);
or U4584 (N_4584,N_4319,N_4364);
nor U4585 (N_4585,N_4264,N_4295);
and U4586 (N_4586,N_4416,N_4363);
nand U4587 (N_4587,N_4362,N_4402);
nor U4588 (N_4588,N_4465,N_4286);
or U4589 (N_4589,N_4450,N_4473);
nand U4590 (N_4590,N_4425,N_4312);
nor U4591 (N_4591,N_4494,N_4368);
nor U4592 (N_4592,N_4360,N_4486);
and U4593 (N_4593,N_4332,N_4437);
nand U4594 (N_4594,N_4468,N_4283);
nor U4595 (N_4595,N_4265,N_4282);
nor U4596 (N_4596,N_4274,N_4485);
and U4597 (N_4597,N_4361,N_4451);
or U4598 (N_4598,N_4355,N_4459);
nor U4599 (N_4599,N_4454,N_4453);
nand U4600 (N_4600,N_4479,N_4475);
nor U4601 (N_4601,N_4330,N_4382);
nor U4602 (N_4602,N_4349,N_4418);
nor U4603 (N_4603,N_4331,N_4442);
nand U4604 (N_4604,N_4438,N_4429);
nand U4605 (N_4605,N_4421,N_4370);
and U4606 (N_4606,N_4462,N_4367);
nand U4607 (N_4607,N_4406,N_4258);
and U4608 (N_4608,N_4430,N_4408);
or U4609 (N_4609,N_4314,N_4315);
nor U4610 (N_4610,N_4378,N_4301);
or U4611 (N_4611,N_4493,N_4411);
and U4612 (N_4612,N_4495,N_4492);
nor U4613 (N_4613,N_4491,N_4344);
and U4614 (N_4614,N_4250,N_4380);
or U4615 (N_4615,N_4352,N_4328);
nor U4616 (N_4616,N_4466,N_4285);
or U4617 (N_4617,N_4256,N_4339);
and U4618 (N_4618,N_4289,N_4275);
and U4619 (N_4619,N_4346,N_4310);
and U4620 (N_4620,N_4299,N_4472);
or U4621 (N_4621,N_4471,N_4487);
nor U4622 (N_4622,N_4290,N_4426);
or U4623 (N_4623,N_4447,N_4292);
xor U4624 (N_4624,N_4251,N_4463);
or U4625 (N_4625,N_4294,N_4361);
and U4626 (N_4626,N_4454,N_4477);
and U4627 (N_4627,N_4353,N_4290);
and U4628 (N_4628,N_4252,N_4328);
and U4629 (N_4629,N_4421,N_4348);
nor U4630 (N_4630,N_4364,N_4333);
nand U4631 (N_4631,N_4326,N_4268);
and U4632 (N_4632,N_4456,N_4332);
nand U4633 (N_4633,N_4290,N_4381);
nor U4634 (N_4634,N_4273,N_4386);
and U4635 (N_4635,N_4417,N_4296);
nor U4636 (N_4636,N_4429,N_4441);
or U4637 (N_4637,N_4251,N_4449);
nor U4638 (N_4638,N_4397,N_4494);
and U4639 (N_4639,N_4494,N_4256);
or U4640 (N_4640,N_4405,N_4463);
or U4641 (N_4641,N_4461,N_4457);
or U4642 (N_4642,N_4496,N_4341);
and U4643 (N_4643,N_4478,N_4476);
nand U4644 (N_4644,N_4358,N_4465);
and U4645 (N_4645,N_4327,N_4436);
or U4646 (N_4646,N_4337,N_4499);
nand U4647 (N_4647,N_4257,N_4286);
nor U4648 (N_4648,N_4304,N_4306);
nand U4649 (N_4649,N_4342,N_4308);
and U4650 (N_4650,N_4467,N_4418);
and U4651 (N_4651,N_4373,N_4406);
and U4652 (N_4652,N_4462,N_4414);
and U4653 (N_4653,N_4332,N_4307);
or U4654 (N_4654,N_4481,N_4428);
and U4655 (N_4655,N_4494,N_4462);
nor U4656 (N_4656,N_4312,N_4443);
nand U4657 (N_4657,N_4470,N_4294);
nand U4658 (N_4658,N_4278,N_4446);
nor U4659 (N_4659,N_4351,N_4308);
and U4660 (N_4660,N_4357,N_4323);
nor U4661 (N_4661,N_4335,N_4405);
nor U4662 (N_4662,N_4332,N_4368);
or U4663 (N_4663,N_4419,N_4449);
nor U4664 (N_4664,N_4468,N_4312);
nand U4665 (N_4665,N_4337,N_4315);
nand U4666 (N_4666,N_4400,N_4306);
nand U4667 (N_4667,N_4313,N_4426);
and U4668 (N_4668,N_4265,N_4357);
nand U4669 (N_4669,N_4302,N_4258);
nand U4670 (N_4670,N_4477,N_4258);
nor U4671 (N_4671,N_4439,N_4310);
and U4672 (N_4672,N_4436,N_4283);
and U4673 (N_4673,N_4348,N_4381);
nand U4674 (N_4674,N_4285,N_4429);
or U4675 (N_4675,N_4305,N_4458);
nand U4676 (N_4676,N_4419,N_4336);
or U4677 (N_4677,N_4403,N_4476);
nor U4678 (N_4678,N_4292,N_4334);
nor U4679 (N_4679,N_4320,N_4406);
nor U4680 (N_4680,N_4477,N_4261);
or U4681 (N_4681,N_4473,N_4490);
and U4682 (N_4682,N_4427,N_4377);
and U4683 (N_4683,N_4274,N_4296);
and U4684 (N_4684,N_4360,N_4297);
or U4685 (N_4685,N_4389,N_4301);
or U4686 (N_4686,N_4363,N_4429);
nand U4687 (N_4687,N_4303,N_4257);
and U4688 (N_4688,N_4417,N_4276);
nor U4689 (N_4689,N_4461,N_4420);
or U4690 (N_4690,N_4359,N_4462);
and U4691 (N_4691,N_4371,N_4285);
nor U4692 (N_4692,N_4408,N_4363);
nand U4693 (N_4693,N_4350,N_4277);
or U4694 (N_4694,N_4383,N_4476);
nand U4695 (N_4695,N_4419,N_4334);
and U4696 (N_4696,N_4274,N_4285);
nor U4697 (N_4697,N_4499,N_4384);
and U4698 (N_4698,N_4372,N_4367);
nand U4699 (N_4699,N_4295,N_4318);
nand U4700 (N_4700,N_4391,N_4254);
nand U4701 (N_4701,N_4375,N_4257);
nand U4702 (N_4702,N_4479,N_4389);
or U4703 (N_4703,N_4356,N_4322);
nor U4704 (N_4704,N_4307,N_4354);
or U4705 (N_4705,N_4263,N_4345);
and U4706 (N_4706,N_4358,N_4336);
or U4707 (N_4707,N_4283,N_4332);
nor U4708 (N_4708,N_4383,N_4251);
or U4709 (N_4709,N_4278,N_4478);
nand U4710 (N_4710,N_4265,N_4317);
nand U4711 (N_4711,N_4276,N_4355);
or U4712 (N_4712,N_4431,N_4389);
and U4713 (N_4713,N_4473,N_4478);
or U4714 (N_4714,N_4299,N_4273);
nor U4715 (N_4715,N_4389,N_4298);
nand U4716 (N_4716,N_4458,N_4360);
or U4717 (N_4717,N_4296,N_4316);
nand U4718 (N_4718,N_4283,N_4342);
or U4719 (N_4719,N_4380,N_4431);
or U4720 (N_4720,N_4336,N_4391);
nand U4721 (N_4721,N_4405,N_4436);
nand U4722 (N_4722,N_4407,N_4340);
nand U4723 (N_4723,N_4307,N_4498);
and U4724 (N_4724,N_4418,N_4340);
or U4725 (N_4725,N_4369,N_4414);
nand U4726 (N_4726,N_4379,N_4269);
and U4727 (N_4727,N_4435,N_4404);
nand U4728 (N_4728,N_4380,N_4488);
nand U4729 (N_4729,N_4265,N_4481);
xor U4730 (N_4730,N_4409,N_4497);
nor U4731 (N_4731,N_4348,N_4321);
or U4732 (N_4732,N_4313,N_4350);
or U4733 (N_4733,N_4339,N_4262);
nand U4734 (N_4734,N_4482,N_4293);
and U4735 (N_4735,N_4344,N_4497);
or U4736 (N_4736,N_4330,N_4396);
xor U4737 (N_4737,N_4463,N_4295);
or U4738 (N_4738,N_4272,N_4367);
nand U4739 (N_4739,N_4426,N_4398);
nand U4740 (N_4740,N_4310,N_4350);
or U4741 (N_4741,N_4432,N_4407);
and U4742 (N_4742,N_4389,N_4367);
nand U4743 (N_4743,N_4445,N_4363);
nand U4744 (N_4744,N_4374,N_4310);
or U4745 (N_4745,N_4265,N_4465);
and U4746 (N_4746,N_4358,N_4423);
or U4747 (N_4747,N_4254,N_4471);
and U4748 (N_4748,N_4443,N_4378);
nor U4749 (N_4749,N_4484,N_4294);
nor U4750 (N_4750,N_4749,N_4552);
nand U4751 (N_4751,N_4656,N_4734);
nor U4752 (N_4752,N_4592,N_4657);
nand U4753 (N_4753,N_4625,N_4745);
nor U4754 (N_4754,N_4722,N_4677);
and U4755 (N_4755,N_4744,N_4702);
nand U4756 (N_4756,N_4645,N_4743);
nor U4757 (N_4757,N_4723,N_4623);
or U4758 (N_4758,N_4616,N_4654);
and U4759 (N_4759,N_4539,N_4605);
or U4760 (N_4760,N_4530,N_4501);
nor U4761 (N_4761,N_4532,N_4538);
nor U4762 (N_4762,N_4600,N_4505);
or U4763 (N_4763,N_4737,N_4720);
and U4764 (N_4764,N_4606,N_4557);
and U4765 (N_4765,N_4621,N_4725);
and U4766 (N_4766,N_4670,N_4627);
or U4767 (N_4767,N_4551,N_4571);
nand U4768 (N_4768,N_4573,N_4578);
or U4769 (N_4769,N_4547,N_4746);
and U4770 (N_4770,N_4739,N_4643);
or U4771 (N_4771,N_4541,N_4611);
nor U4772 (N_4772,N_4704,N_4558);
nand U4773 (N_4773,N_4515,N_4663);
and U4774 (N_4774,N_4634,N_4700);
nand U4775 (N_4775,N_4672,N_4610);
nor U4776 (N_4776,N_4527,N_4597);
or U4777 (N_4777,N_4553,N_4651);
nand U4778 (N_4778,N_4554,N_4546);
or U4779 (N_4779,N_4686,N_4735);
or U4780 (N_4780,N_4537,N_4510);
or U4781 (N_4781,N_4563,N_4718);
nor U4782 (N_4782,N_4521,N_4646);
nor U4783 (N_4783,N_4727,N_4613);
nand U4784 (N_4784,N_4655,N_4642);
nand U4785 (N_4785,N_4580,N_4641);
nor U4786 (N_4786,N_4748,N_4639);
and U4787 (N_4787,N_4731,N_4703);
nor U4788 (N_4788,N_4583,N_4589);
nor U4789 (N_4789,N_4667,N_4518);
and U4790 (N_4790,N_4692,N_4635);
or U4791 (N_4791,N_4705,N_4526);
nor U4792 (N_4792,N_4716,N_4717);
and U4793 (N_4793,N_4682,N_4556);
nor U4794 (N_4794,N_4548,N_4649);
nand U4795 (N_4795,N_4564,N_4522);
and U4796 (N_4796,N_4650,N_4508);
and U4797 (N_4797,N_4601,N_4608);
and U4798 (N_4798,N_4624,N_4588);
or U4799 (N_4799,N_4685,N_4647);
nand U4800 (N_4800,N_4706,N_4579);
and U4801 (N_4801,N_4604,N_4586);
nor U4802 (N_4802,N_4721,N_4528);
nand U4803 (N_4803,N_4695,N_4545);
or U4804 (N_4804,N_4740,N_4659);
nand U4805 (N_4805,N_4535,N_4543);
nor U4806 (N_4806,N_4628,N_4559);
nand U4807 (N_4807,N_4509,N_4728);
nor U4808 (N_4808,N_4517,N_4617);
nand U4809 (N_4809,N_4512,N_4742);
nand U4810 (N_4810,N_4693,N_4637);
or U4811 (N_4811,N_4631,N_4507);
and U4812 (N_4812,N_4511,N_4683);
or U4813 (N_4813,N_4567,N_4697);
nand U4814 (N_4814,N_4719,N_4593);
or U4815 (N_4815,N_4555,N_4678);
nand U4816 (N_4816,N_4690,N_4688);
and U4817 (N_4817,N_4595,N_4500);
nor U4818 (N_4818,N_4569,N_4640);
nor U4819 (N_4819,N_4701,N_4529);
nand U4820 (N_4820,N_4707,N_4665);
nor U4821 (N_4821,N_4599,N_4536);
nor U4822 (N_4822,N_4738,N_4630);
or U4823 (N_4823,N_4516,N_4747);
or U4824 (N_4824,N_4615,N_4603);
nor U4825 (N_4825,N_4523,N_4503);
nor U4826 (N_4826,N_4575,N_4662);
nor U4827 (N_4827,N_4544,N_4542);
or U4828 (N_4828,N_4708,N_4561);
or U4829 (N_4829,N_4582,N_4609);
and U4830 (N_4830,N_4620,N_4562);
nor U4831 (N_4831,N_4712,N_4669);
or U4832 (N_4832,N_4596,N_4602);
and U4833 (N_4833,N_4622,N_4633);
and U4834 (N_4834,N_4591,N_4619);
nand U4835 (N_4835,N_4681,N_4698);
and U4836 (N_4836,N_4694,N_4713);
or U4837 (N_4837,N_4540,N_4676);
and U4838 (N_4838,N_4566,N_4671);
nor U4839 (N_4839,N_4724,N_4666);
nor U4840 (N_4840,N_4661,N_4581);
nor U4841 (N_4841,N_4560,N_4550);
nand U4842 (N_4842,N_4570,N_4715);
nor U4843 (N_4843,N_4587,N_4504);
nor U4844 (N_4844,N_4626,N_4574);
nand U4845 (N_4845,N_4520,N_4514);
and U4846 (N_4846,N_4733,N_4691);
or U4847 (N_4847,N_4644,N_4584);
and U4848 (N_4848,N_4699,N_4598);
and U4849 (N_4849,N_4668,N_4648);
nand U4850 (N_4850,N_4696,N_4709);
or U4851 (N_4851,N_4513,N_4632);
nor U4852 (N_4852,N_4629,N_4732);
nor U4853 (N_4853,N_4568,N_4687);
nor U4854 (N_4854,N_4652,N_4664);
or U4855 (N_4855,N_4590,N_4531);
nand U4856 (N_4856,N_4565,N_4660);
nor U4857 (N_4857,N_4638,N_4680);
and U4858 (N_4858,N_4711,N_4730);
or U4859 (N_4859,N_4736,N_4549);
nor U4860 (N_4860,N_4572,N_4506);
nor U4861 (N_4861,N_4533,N_4675);
nand U4862 (N_4862,N_4618,N_4534);
and U4863 (N_4863,N_4594,N_4714);
and U4864 (N_4864,N_4653,N_4689);
or U4865 (N_4865,N_4679,N_4612);
and U4866 (N_4866,N_4502,N_4726);
and U4867 (N_4867,N_4607,N_4576);
xnor U4868 (N_4868,N_4525,N_4577);
and U4869 (N_4869,N_4674,N_4729);
nand U4870 (N_4870,N_4519,N_4673);
or U4871 (N_4871,N_4585,N_4741);
or U4872 (N_4872,N_4524,N_4710);
nor U4873 (N_4873,N_4614,N_4636);
nor U4874 (N_4874,N_4684,N_4658);
nor U4875 (N_4875,N_4696,N_4708);
or U4876 (N_4876,N_4745,N_4640);
or U4877 (N_4877,N_4504,N_4663);
or U4878 (N_4878,N_4508,N_4645);
nand U4879 (N_4879,N_4515,N_4571);
nand U4880 (N_4880,N_4710,N_4630);
nand U4881 (N_4881,N_4655,N_4666);
and U4882 (N_4882,N_4585,N_4733);
or U4883 (N_4883,N_4621,N_4602);
and U4884 (N_4884,N_4653,N_4685);
or U4885 (N_4885,N_4622,N_4666);
nor U4886 (N_4886,N_4526,N_4570);
and U4887 (N_4887,N_4650,N_4628);
and U4888 (N_4888,N_4544,N_4618);
nor U4889 (N_4889,N_4513,N_4578);
nor U4890 (N_4890,N_4681,N_4694);
or U4891 (N_4891,N_4577,N_4712);
or U4892 (N_4892,N_4678,N_4688);
nand U4893 (N_4893,N_4704,N_4737);
and U4894 (N_4894,N_4682,N_4524);
and U4895 (N_4895,N_4542,N_4606);
xor U4896 (N_4896,N_4508,N_4666);
nand U4897 (N_4897,N_4706,N_4700);
and U4898 (N_4898,N_4582,N_4672);
nor U4899 (N_4899,N_4743,N_4644);
and U4900 (N_4900,N_4654,N_4734);
or U4901 (N_4901,N_4713,N_4600);
nor U4902 (N_4902,N_4628,N_4555);
nand U4903 (N_4903,N_4721,N_4658);
and U4904 (N_4904,N_4602,N_4699);
and U4905 (N_4905,N_4657,N_4699);
nor U4906 (N_4906,N_4650,N_4563);
nor U4907 (N_4907,N_4532,N_4731);
nor U4908 (N_4908,N_4535,N_4583);
nand U4909 (N_4909,N_4684,N_4686);
and U4910 (N_4910,N_4625,N_4510);
and U4911 (N_4911,N_4661,N_4649);
or U4912 (N_4912,N_4677,N_4573);
or U4913 (N_4913,N_4629,N_4611);
nor U4914 (N_4914,N_4504,N_4584);
or U4915 (N_4915,N_4735,N_4529);
nand U4916 (N_4916,N_4585,N_4572);
nor U4917 (N_4917,N_4728,N_4624);
or U4918 (N_4918,N_4695,N_4596);
nor U4919 (N_4919,N_4589,N_4543);
nor U4920 (N_4920,N_4633,N_4634);
nor U4921 (N_4921,N_4539,N_4690);
nor U4922 (N_4922,N_4643,N_4642);
nand U4923 (N_4923,N_4713,N_4515);
nand U4924 (N_4924,N_4518,N_4560);
and U4925 (N_4925,N_4518,N_4620);
and U4926 (N_4926,N_4556,N_4568);
nand U4927 (N_4927,N_4660,N_4728);
nor U4928 (N_4928,N_4718,N_4542);
nand U4929 (N_4929,N_4511,N_4716);
nor U4930 (N_4930,N_4571,N_4617);
nand U4931 (N_4931,N_4573,N_4545);
and U4932 (N_4932,N_4699,N_4668);
nand U4933 (N_4933,N_4719,N_4607);
or U4934 (N_4934,N_4634,N_4738);
or U4935 (N_4935,N_4679,N_4560);
nand U4936 (N_4936,N_4629,N_4548);
nand U4937 (N_4937,N_4700,N_4612);
or U4938 (N_4938,N_4575,N_4551);
nand U4939 (N_4939,N_4714,N_4679);
or U4940 (N_4940,N_4544,N_4634);
nor U4941 (N_4941,N_4537,N_4563);
and U4942 (N_4942,N_4582,N_4531);
nor U4943 (N_4943,N_4661,N_4601);
nor U4944 (N_4944,N_4575,N_4507);
and U4945 (N_4945,N_4671,N_4614);
nor U4946 (N_4946,N_4557,N_4550);
and U4947 (N_4947,N_4684,N_4538);
and U4948 (N_4948,N_4503,N_4513);
and U4949 (N_4949,N_4537,N_4559);
nor U4950 (N_4950,N_4687,N_4621);
nor U4951 (N_4951,N_4664,N_4676);
nand U4952 (N_4952,N_4588,N_4600);
nor U4953 (N_4953,N_4748,N_4680);
or U4954 (N_4954,N_4547,N_4674);
and U4955 (N_4955,N_4740,N_4568);
and U4956 (N_4956,N_4627,N_4631);
or U4957 (N_4957,N_4501,N_4748);
nor U4958 (N_4958,N_4512,N_4708);
nor U4959 (N_4959,N_4526,N_4614);
or U4960 (N_4960,N_4606,N_4643);
nand U4961 (N_4961,N_4744,N_4572);
or U4962 (N_4962,N_4626,N_4681);
or U4963 (N_4963,N_4612,N_4591);
nand U4964 (N_4964,N_4546,N_4665);
or U4965 (N_4965,N_4738,N_4726);
nor U4966 (N_4966,N_4698,N_4501);
nor U4967 (N_4967,N_4506,N_4682);
nor U4968 (N_4968,N_4745,N_4644);
and U4969 (N_4969,N_4578,N_4647);
nand U4970 (N_4970,N_4701,N_4619);
nand U4971 (N_4971,N_4739,N_4557);
nand U4972 (N_4972,N_4575,N_4606);
nand U4973 (N_4973,N_4727,N_4580);
nand U4974 (N_4974,N_4631,N_4596);
nand U4975 (N_4975,N_4702,N_4592);
nand U4976 (N_4976,N_4589,N_4630);
and U4977 (N_4977,N_4596,N_4661);
or U4978 (N_4978,N_4721,N_4539);
nand U4979 (N_4979,N_4713,N_4655);
nor U4980 (N_4980,N_4568,N_4720);
nor U4981 (N_4981,N_4717,N_4707);
and U4982 (N_4982,N_4747,N_4575);
and U4983 (N_4983,N_4516,N_4635);
and U4984 (N_4984,N_4707,N_4697);
nor U4985 (N_4985,N_4584,N_4681);
nand U4986 (N_4986,N_4544,N_4580);
or U4987 (N_4987,N_4683,N_4632);
or U4988 (N_4988,N_4684,N_4716);
nand U4989 (N_4989,N_4649,N_4662);
nor U4990 (N_4990,N_4599,N_4690);
nor U4991 (N_4991,N_4638,N_4624);
or U4992 (N_4992,N_4705,N_4561);
or U4993 (N_4993,N_4650,N_4562);
nand U4994 (N_4994,N_4638,N_4629);
and U4995 (N_4995,N_4709,N_4556);
or U4996 (N_4996,N_4620,N_4533);
nand U4997 (N_4997,N_4520,N_4691);
or U4998 (N_4998,N_4578,N_4710);
nor U4999 (N_4999,N_4719,N_4733);
nand U5000 (N_5000,N_4959,N_4769);
or U5001 (N_5001,N_4967,N_4816);
nand U5002 (N_5002,N_4779,N_4883);
or U5003 (N_5003,N_4940,N_4792);
nor U5004 (N_5004,N_4780,N_4810);
or U5005 (N_5005,N_4838,N_4938);
or U5006 (N_5006,N_4950,N_4818);
nor U5007 (N_5007,N_4970,N_4943);
nand U5008 (N_5008,N_4977,N_4922);
nor U5009 (N_5009,N_4806,N_4876);
nor U5010 (N_5010,N_4899,N_4781);
nor U5011 (N_5011,N_4969,N_4881);
or U5012 (N_5012,N_4912,N_4993);
nand U5013 (N_5013,N_4803,N_4962);
and U5014 (N_5014,N_4885,N_4917);
nand U5015 (N_5015,N_4773,N_4937);
and U5016 (N_5016,N_4907,N_4765);
nand U5017 (N_5017,N_4869,N_4985);
and U5018 (N_5018,N_4819,N_4889);
nand U5019 (N_5019,N_4972,N_4976);
or U5020 (N_5020,N_4960,N_4989);
nor U5021 (N_5021,N_4788,N_4915);
nand U5022 (N_5022,N_4975,N_4945);
and U5023 (N_5023,N_4790,N_4867);
nand U5024 (N_5024,N_4798,N_4903);
and U5025 (N_5025,N_4898,N_4764);
or U5026 (N_5026,N_4865,N_4956);
nor U5027 (N_5027,N_4766,N_4951);
and U5028 (N_5028,N_4952,N_4910);
nand U5029 (N_5029,N_4995,N_4758);
and U5030 (N_5030,N_4866,N_4813);
nand U5031 (N_5031,N_4785,N_4777);
nor U5032 (N_5032,N_4759,N_4942);
and U5033 (N_5033,N_4750,N_4856);
nor U5034 (N_5034,N_4795,N_4994);
and U5035 (N_5035,N_4913,N_4988);
nand U5036 (N_5036,N_4918,N_4770);
nand U5037 (N_5037,N_4939,N_4804);
nor U5038 (N_5038,N_4833,N_4776);
nor U5039 (N_5039,N_4891,N_4927);
nand U5040 (N_5040,N_4932,N_4986);
nor U5041 (N_5041,N_4755,N_4886);
or U5042 (N_5042,N_4973,N_4857);
and U5043 (N_5043,N_4829,N_4826);
and U5044 (N_5044,N_4812,N_4884);
nand U5045 (N_5045,N_4753,N_4895);
nand U5046 (N_5046,N_4793,N_4842);
and U5047 (N_5047,N_4957,N_4852);
and U5048 (N_5048,N_4953,N_4831);
or U5049 (N_5049,N_4999,N_4835);
and U5050 (N_5050,N_4958,N_4966);
nor U5051 (N_5051,N_4875,N_4862);
and U5052 (N_5052,N_4752,N_4944);
nand U5053 (N_5053,N_4815,N_4859);
nand U5054 (N_5054,N_4978,N_4871);
and U5055 (N_5055,N_4929,N_4787);
nand U5056 (N_5056,N_4968,N_4800);
and U5057 (N_5057,N_4822,N_4870);
and U5058 (N_5058,N_4981,N_4778);
nand U5059 (N_5059,N_4930,N_4897);
or U5060 (N_5060,N_4916,N_4820);
nand U5061 (N_5061,N_4955,N_4805);
nand U5062 (N_5062,N_4855,N_4762);
and U5063 (N_5063,N_4877,N_4823);
and U5064 (N_5064,N_4992,N_4987);
nand U5065 (N_5065,N_4980,N_4996);
nand U5066 (N_5066,N_4919,N_4757);
and U5067 (N_5067,N_4825,N_4754);
nand U5068 (N_5068,N_4834,N_4843);
nor U5069 (N_5069,N_4911,N_4900);
nor U5070 (N_5070,N_4828,N_4901);
nor U5071 (N_5071,N_4947,N_4783);
and U5072 (N_5072,N_4761,N_4832);
or U5073 (N_5073,N_4905,N_4896);
nand U5074 (N_5074,N_4914,N_4949);
nor U5075 (N_5075,N_4946,N_4873);
or U5076 (N_5076,N_4904,N_4814);
and U5077 (N_5077,N_4933,N_4979);
nor U5078 (N_5078,N_4909,N_4984);
xnor U5079 (N_5079,N_4850,N_4971);
nor U5080 (N_5080,N_4756,N_4880);
nand U5081 (N_5081,N_4954,N_4965);
or U5082 (N_5082,N_4768,N_4948);
or U5083 (N_5083,N_4854,N_4863);
and U5084 (N_5084,N_4796,N_4963);
and U5085 (N_5085,N_4990,N_4797);
nor U5086 (N_5086,N_4847,N_4921);
or U5087 (N_5087,N_4935,N_4827);
or U5088 (N_5088,N_4861,N_4771);
or U5089 (N_5089,N_4925,N_4974);
nand U5090 (N_5090,N_4821,N_4920);
nand U5091 (N_5091,N_4888,N_4936);
nor U5092 (N_5092,N_4786,N_4964);
and U5093 (N_5093,N_4961,N_4893);
and U5094 (N_5094,N_4928,N_4878);
and U5095 (N_5095,N_4851,N_4887);
nand U5096 (N_5096,N_4902,N_4845);
nand U5097 (N_5097,N_4794,N_4874);
nor U5098 (N_5098,N_4811,N_4890);
nand U5099 (N_5099,N_4848,N_4840);
and U5100 (N_5100,N_4791,N_4849);
nor U5101 (N_5101,N_4872,N_4983);
nand U5102 (N_5102,N_4751,N_4998);
nor U5103 (N_5103,N_4808,N_4908);
or U5104 (N_5104,N_4799,N_4894);
nor U5105 (N_5105,N_4824,N_4868);
or U5106 (N_5106,N_4892,N_4923);
or U5107 (N_5107,N_4846,N_4837);
or U5108 (N_5108,N_4882,N_4789);
nor U5109 (N_5109,N_4772,N_4844);
and U5110 (N_5110,N_4836,N_4767);
or U5111 (N_5111,N_4830,N_4941);
nand U5112 (N_5112,N_4760,N_4991);
nand U5113 (N_5113,N_4926,N_4782);
nor U5114 (N_5114,N_4982,N_4802);
nand U5115 (N_5115,N_4817,N_4763);
nand U5116 (N_5116,N_4774,N_4858);
nand U5117 (N_5117,N_4997,N_4784);
or U5118 (N_5118,N_4775,N_4853);
and U5119 (N_5119,N_4906,N_4879);
nor U5120 (N_5120,N_4841,N_4809);
nor U5121 (N_5121,N_4807,N_4839);
nor U5122 (N_5122,N_4801,N_4934);
or U5123 (N_5123,N_4931,N_4924);
and U5124 (N_5124,N_4864,N_4860);
and U5125 (N_5125,N_4940,N_4794);
nor U5126 (N_5126,N_4858,N_4766);
and U5127 (N_5127,N_4921,N_4826);
and U5128 (N_5128,N_4792,N_4910);
nand U5129 (N_5129,N_4763,N_4885);
nand U5130 (N_5130,N_4988,N_4934);
nor U5131 (N_5131,N_4829,N_4899);
or U5132 (N_5132,N_4756,N_4896);
or U5133 (N_5133,N_4848,N_4914);
nand U5134 (N_5134,N_4838,N_4986);
nand U5135 (N_5135,N_4863,N_4927);
nor U5136 (N_5136,N_4861,N_4970);
nor U5137 (N_5137,N_4890,N_4898);
nand U5138 (N_5138,N_4896,N_4992);
and U5139 (N_5139,N_4956,N_4913);
nor U5140 (N_5140,N_4771,N_4791);
or U5141 (N_5141,N_4890,N_4986);
and U5142 (N_5142,N_4757,N_4937);
nand U5143 (N_5143,N_4820,N_4833);
and U5144 (N_5144,N_4816,N_4800);
or U5145 (N_5145,N_4889,N_4774);
nor U5146 (N_5146,N_4966,N_4987);
nand U5147 (N_5147,N_4754,N_4780);
nor U5148 (N_5148,N_4835,N_4886);
and U5149 (N_5149,N_4759,N_4979);
nor U5150 (N_5150,N_4818,N_4988);
nor U5151 (N_5151,N_4872,N_4870);
nand U5152 (N_5152,N_4833,N_4926);
or U5153 (N_5153,N_4864,N_4945);
nand U5154 (N_5154,N_4970,N_4915);
or U5155 (N_5155,N_4953,N_4778);
nor U5156 (N_5156,N_4792,N_4935);
nand U5157 (N_5157,N_4768,N_4849);
or U5158 (N_5158,N_4998,N_4863);
nand U5159 (N_5159,N_4876,N_4909);
or U5160 (N_5160,N_4835,N_4983);
or U5161 (N_5161,N_4808,N_4851);
or U5162 (N_5162,N_4855,N_4992);
nor U5163 (N_5163,N_4851,N_4930);
nand U5164 (N_5164,N_4762,N_4934);
or U5165 (N_5165,N_4978,N_4824);
or U5166 (N_5166,N_4796,N_4804);
and U5167 (N_5167,N_4811,N_4842);
or U5168 (N_5168,N_4819,N_4781);
and U5169 (N_5169,N_4995,N_4762);
nor U5170 (N_5170,N_4973,N_4970);
or U5171 (N_5171,N_4901,N_4964);
nor U5172 (N_5172,N_4751,N_4975);
nand U5173 (N_5173,N_4751,N_4811);
nand U5174 (N_5174,N_4933,N_4872);
and U5175 (N_5175,N_4950,N_4889);
or U5176 (N_5176,N_4878,N_4839);
nor U5177 (N_5177,N_4901,N_4830);
nand U5178 (N_5178,N_4756,N_4891);
nor U5179 (N_5179,N_4873,N_4823);
nand U5180 (N_5180,N_4849,N_4890);
nor U5181 (N_5181,N_4970,N_4908);
or U5182 (N_5182,N_4917,N_4866);
and U5183 (N_5183,N_4899,N_4930);
nor U5184 (N_5184,N_4868,N_4818);
or U5185 (N_5185,N_4868,N_4886);
and U5186 (N_5186,N_4843,N_4990);
nor U5187 (N_5187,N_4874,N_4782);
or U5188 (N_5188,N_4886,N_4972);
or U5189 (N_5189,N_4857,N_4976);
and U5190 (N_5190,N_4972,N_4940);
or U5191 (N_5191,N_4915,N_4823);
nand U5192 (N_5192,N_4825,N_4991);
nor U5193 (N_5193,N_4796,N_4844);
nor U5194 (N_5194,N_4843,N_4825);
nand U5195 (N_5195,N_4831,N_4779);
nor U5196 (N_5196,N_4957,N_4973);
nand U5197 (N_5197,N_4894,N_4901);
nor U5198 (N_5198,N_4812,N_4967);
nand U5199 (N_5199,N_4751,N_4878);
nor U5200 (N_5200,N_4962,N_4867);
or U5201 (N_5201,N_4972,N_4900);
and U5202 (N_5202,N_4815,N_4964);
or U5203 (N_5203,N_4983,N_4869);
and U5204 (N_5204,N_4819,N_4780);
or U5205 (N_5205,N_4843,N_4936);
nand U5206 (N_5206,N_4790,N_4785);
or U5207 (N_5207,N_4849,N_4750);
or U5208 (N_5208,N_4818,N_4785);
and U5209 (N_5209,N_4920,N_4868);
or U5210 (N_5210,N_4928,N_4834);
and U5211 (N_5211,N_4986,N_4833);
nand U5212 (N_5212,N_4824,N_4888);
nor U5213 (N_5213,N_4836,N_4869);
or U5214 (N_5214,N_4777,N_4896);
nand U5215 (N_5215,N_4757,N_4968);
nor U5216 (N_5216,N_4853,N_4946);
nor U5217 (N_5217,N_4967,N_4996);
nor U5218 (N_5218,N_4943,N_4949);
nand U5219 (N_5219,N_4818,N_4975);
nand U5220 (N_5220,N_4855,N_4896);
and U5221 (N_5221,N_4824,N_4950);
nor U5222 (N_5222,N_4774,N_4986);
nor U5223 (N_5223,N_4947,N_4971);
and U5224 (N_5224,N_4878,N_4857);
nand U5225 (N_5225,N_4931,N_4980);
nand U5226 (N_5226,N_4908,N_4959);
or U5227 (N_5227,N_4951,N_4809);
and U5228 (N_5228,N_4967,N_4911);
and U5229 (N_5229,N_4840,N_4818);
nor U5230 (N_5230,N_4906,N_4857);
and U5231 (N_5231,N_4828,N_4910);
or U5232 (N_5232,N_4806,N_4987);
and U5233 (N_5233,N_4791,N_4781);
and U5234 (N_5234,N_4755,N_4783);
or U5235 (N_5235,N_4851,N_4852);
and U5236 (N_5236,N_4991,N_4933);
or U5237 (N_5237,N_4941,N_4918);
or U5238 (N_5238,N_4814,N_4765);
and U5239 (N_5239,N_4869,N_4777);
or U5240 (N_5240,N_4785,N_4753);
or U5241 (N_5241,N_4985,N_4829);
nand U5242 (N_5242,N_4764,N_4941);
nand U5243 (N_5243,N_4771,N_4951);
and U5244 (N_5244,N_4852,N_4862);
nand U5245 (N_5245,N_4900,N_4969);
and U5246 (N_5246,N_4802,N_4949);
or U5247 (N_5247,N_4764,N_4899);
or U5248 (N_5248,N_4885,N_4990);
nand U5249 (N_5249,N_4805,N_4819);
and U5250 (N_5250,N_5154,N_5007);
nand U5251 (N_5251,N_5220,N_5199);
and U5252 (N_5252,N_5004,N_5071);
nand U5253 (N_5253,N_5018,N_5129);
nor U5254 (N_5254,N_5001,N_5140);
and U5255 (N_5255,N_5157,N_5052);
or U5256 (N_5256,N_5170,N_5248);
nor U5257 (N_5257,N_5247,N_5207);
nand U5258 (N_5258,N_5091,N_5108);
and U5259 (N_5259,N_5229,N_5069);
and U5260 (N_5260,N_5147,N_5133);
or U5261 (N_5261,N_5121,N_5060);
nand U5262 (N_5262,N_5160,N_5130);
nor U5263 (N_5263,N_5212,N_5137);
or U5264 (N_5264,N_5092,N_5187);
or U5265 (N_5265,N_5036,N_5010);
nor U5266 (N_5266,N_5233,N_5003);
or U5267 (N_5267,N_5245,N_5169);
or U5268 (N_5268,N_5019,N_5043);
and U5269 (N_5269,N_5230,N_5066);
and U5270 (N_5270,N_5041,N_5242);
or U5271 (N_5271,N_5006,N_5005);
nand U5272 (N_5272,N_5163,N_5132);
and U5273 (N_5273,N_5135,N_5032);
nand U5274 (N_5274,N_5072,N_5175);
and U5275 (N_5275,N_5030,N_5167);
nand U5276 (N_5276,N_5144,N_5081);
nand U5277 (N_5277,N_5090,N_5008);
or U5278 (N_5278,N_5044,N_5115);
nor U5279 (N_5279,N_5033,N_5200);
nand U5280 (N_5280,N_5075,N_5240);
or U5281 (N_5281,N_5011,N_5182);
or U5282 (N_5282,N_5151,N_5078);
nand U5283 (N_5283,N_5020,N_5225);
or U5284 (N_5284,N_5236,N_5101);
nor U5285 (N_5285,N_5205,N_5249);
nor U5286 (N_5286,N_5062,N_5150);
nor U5287 (N_5287,N_5246,N_5067);
nand U5288 (N_5288,N_5038,N_5219);
nor U5289 (N_5289,N_5215,N_5244);
and U5290 (N_5290,N_5166,N_5149);
or U5291 (N_5291,N_5145,N_5012);
or U5292 (N_5292,N_5055,N_5158);
and U5293 (N_5293,N_5234,N_5123);
nor U5294 (N_5294,N_5024,N_5107);
and U5295 (N_5295,N_5079,N_5028);
nor U5296 (N_5296,N_5180,N_5177);
nor U5297 (N_5297,N_5085,N_5088);
nor U5298 (N_5298,N_5102,N_5161);
or U5299 (N_5299,N_5217,N_5156);
nand U5300 (N_5300,N_5174,N_5098);
nor U5301 (N_5301,N_5216,N_5082);
and U5302 (N_5302,N_5164,N_5031);
nor U5303 (N_5303,N_5083,N_5226);
and U5304 (N_5304,N_5143,N_5221);
and U5305 (N_5305,N_5025,N_5027);
and U5306 (N_5306,N_5209,N_5112);
and U5307 (N_5307,N_5224,N_5086);
and U5308 (N_5308,N_5120,N_5077);
nand U5309 (N_5309,N_5204,N_5218);
and U5310 (N_5310,N_5022,N_5045);
or U5311 (N_5311,N_5124,N_5070);
nand U5312 (N_5312,N_5184,N_5089);
and U5313 (N_5313,N_5100,N_5047);
or U5314 (N_5314,N_5119,N_5165);
nand U5315 (N_5315,N_5073,N_5065);
and U5316 (N_5316,N_5015,N_5155);
nor U5317 (N_5317,N_5168,N_5017);
and U5318 (N_5318,N_5105,N_5223);
or U5319 (N_5319,N_5189,N_5197);
nor U5320 (N_5320,N_5040,N_5064);
and U5321 (N_5321,N_5099,N_5152);
nor U5322 (N_5322,N_5059,N_5111);
nand U5323 (N_5323,N_5171,N_5113);
or U5324 (N_5324,N_5231,N_5185);
and U5325 (N_5325,N_5153,N_5178);
or U5326 (N_5326,N_5035,N_5176);
nand U5327 (N_5327,N_5116,N_5138);
nor U5328 (N_5328,N_5181,N_5014);
nand U5329 (N_5329,N_5068,N_5084);
and U5330 (N_5330,N_5106,N_5002);
xor U5331 (N_5331,N_5211,N_5037);
and U5332 (N_5332,N_5188,N_5227);
nand U5333 (N_5333,N_5114,N_5186);
nand U5334 (N_5334,N_5162,N_5243);
nand U5335 (N_5335,N_5080,N_5048);
nor U5336 (N_5336,N_5009,N_5029);
and U5337 (N_5337,N_5054,N_5093);
nand U5338 (N_5338,N_5046,N_5183);
and U5339 (N_5339,N_5050,N_5125);
and U5340 (N_5340,N_5238,N_5104);
xor U5341 (N_5341,N_5016,N_5173);
and U5342 (N_5342,N_5237,N_5201);
or U5343 (N_5343,N_5023,N_5131);
nor U5344 (N_5344,N_5159,N_5203);
or U5345 (N_5345,N_5128,N_5039);
and U5346 (N_5346,N_5206,N_5214);
nand U5347 (N_5347,N_5076,N_5042);
nor U5348 (N_5348,N_5061,N_5192);
nand U5349 (N_5349,N_5056,N_5136);
nor U5350 (N_5350,N_5122,N_5095);
or U5351 (N_5351,N_5117,N_5026);
nor U5352 (N_5352,N_5097,N_5094);
nand U5353 (N_5353,N_5146,N_5110);
and U5354 (N_5354,N_5142,N_5208);
nor U5355 (N_5355,N_5058,N_5109);
nor U5356 (N_5356,N_5049,N_5103);
nand U5357 (N_5357,N_5126,N_5213);
and U5358 (N_5358,N_5196,N_5190);
and U5359 (N_5359,N_5051,N_5063);
nand U5360 (N_5360,N_5118,N_5053);
nor U5361 (N_5361,N_5127,N_5148);
nand U5362 (N_5362,N_5000,N_5134);
or U5363 (N_5363,N_5235,N_5193);
or U5364 (N_5364,N_5191,N_5232);
nor U5365 (N_5365,N_5195,N_5087);
and U5366 (N_5366,N_5074,N_5179);
nand U5367 (N_5367,N_5241,N_5210);
nor U5368 (N_5368,N_5194,N_5139);
nand U5369 (N_5369,N_5034,N_5096);
and U5370 (N_5370,N_5239,N_5228);
xor U5371 (N_5371,N_5021,N_5013);
and U5372 (N_5372,N_5222,N_5141);
nand U5373 (N_5373,N_5057,N_5202);
nand U5374 (N_5374,N_5198,N_5172);
or U5375 (N_5375,N_5082,N_5116);
nor U5376 (N_5376,N_5053,N_5112);
and U5377 (N_5377,N_5185,N_5232);
or U5378 (N_5378,N_5152,N_5014);
xor U5379 (N_5379,N_5232,N_5089);
and U5380 (N_5380,N_5076,N_5032);
nor U5381 (N_5381,N_5166,N_5154);
nand U5382 (N_5382,N_5031,N_5229);
or U5383 (N_5383,N_5160,N_5185);
nor U5384 (N_5384,N_5229,N_5160);
or U5385 (N_5385,N_5227,N_5092);
nand U5386 (N_5386,N_5142,N_5246);
nand U5387 (N_5387,N_5234,N_5226);
and U5388 (N_5388,N_5095,N_5021);
nor U5389 (N_5389,N_5174,N_5208);
or U5390 (N_5390,N_5248,N_5178);
and U5391 (N_5391,N_5239,N_5170);
and U5392 (N_5392,N_5127,N_5139);
and U5393 (N_5393,N_5181,N_5153);
nor U5394 (N_5394,N_5061,N_5212);
nor U5395 (N_5395,N_5210,N_5032);
nand U5396 (N_5396,N_5164,N_5150);
or U5397 (N_5397,N_5130,N_5122);
nand U5398 (N_5398,N_5200,N_5119);
and U5399 (N_5399,N_5133,N_5196);
nor U5400 (N_5400,N_5024,N_5207);
nor U5401 (N_5401,N_5134,N_5186);
or U5402 (N_5402,N_5112,N_5248);
or U5403 (N_5403,N_5212,N_5020);
nor U5404 (N_5404,N_5229,N_5086);
and U5405 (N_5405,N_5155,N_5216);
nor U5406 (N_5406,N_5006,N_5094);
nor U5407 (N_5407,N_5064,N_5010);
and U5408 (N_5408,N_5037,N_5187);
and U5409 (N_5409,N_5023,N_5106);
or U5410 (N_5410,N_5213,N_5215);
nand U5411 (N_5411,N_5142,N_5034);
nor U5412 (N_5412,N_5044,N_5166);
and U5413 (N_5413,N_5030,N_5175);
and U5414 (N_5414,N_5212,N_5095);
nor U5415 (N_5415,N_5171,N_5048);
nor U5416 (N_5416,N_5130,N_5102);
and U5417 (N_5417,N_5013,N_5060);
or U5418 (N_5418,N_5074,N_5195);
and U5419 (N_5419,N_5080,N_5068);
xor U5420 (N_5420,N_5211,N_5149);
nor U5421 (N_5421,N_5093,N_5012);
nor U5422 (N_5422,N_5141,N_5185);
and U5423 (N_5423,N_5146,N_5084);
nor U5424 (N_5424,N_5105,N_5245);
or U5425 (N_5425,N_5072,N_5008);
nor U5426 (N_5426,N_5053,N_5091);
or U5427 (N_5427,N_5054,N_5207);
nand U5428 (N_5428,N_5116,N_5006);
or U5429 (N_5429,N_5230,N_5063);
and U5430 (N_5430,N_5060,N_5048);
nor U5431 (N_5431,N_5103,N_5191);
nand U5432 (N_5432,N_5179,N_5079);
nand U5433 (N_5433,N_5201,N_5068);
or U5434 (N_5434,N_5101,N_5215);
nor U5435 (N_5435,N_5125,N_5066);
nor U5436 (N_5436,N_5170,N_5114);
nor U5437 (N_5437,N_5130,N_5191);
and U5438 (N_5438,N_5171,N_5192);
nor U5439 (N_5439,N_5142,N_5071);
nand U5440 (N_5440,N_5035,N_5033);
and U5441 (N_5441,N_5136,N_5020);
nand U5442 (N_5442,N_5190,N_5007);
xor U5443 (N_5443,N_5022,N_5167);
nor U5444 (N_5444,N_5168,N_5100);
nand U5445 (N_5445,N_5130,N_5224);
nor U5446 (N_5446,N_5246,N_5189);
or U5447 (N_5447,N_5156,N_5079);
or U5448 (N_5448,N_5239,N_5110);
and U5449 (N_5449,N_5153,N_5109);
and U5450 (N_5450,N_5099,N_5043);
and U5451 (N_5451,N_5238,N_5217);
nor U5452 (N_5452,N_5173,N_5241);
or U5453 (N_5453,N_5172,N_5011);
nand U5454 (N_5454,N_5160,N_5017);
and U5455 (N_5455,N_5172,N_5130);
and U5456 (N_5456,N_5117,N_5162);
and U5457 (N_5457,N_5099,N_5212);
and U5458 (N_5458,N_5214,N_5232);
and U5459 (N_5459,N_5113,N_5199);
or U5460 (N_5460,N_5088,N_5136);
nor U5461 (N_5461,N_5123,N_5191);
or U5462 (N_5462,N_5050,N_5102);
and U5463 (N_5463,N_5059,N_5094);
nand U5464 (N_5464,N_5182,N_5080);
nand U5465 (N_5465,N_5230,N_5185);
and U5466 (N_5466,N_5028,N_5164);
or U5467 (N_5467,N_5157,N_5022);
nor U5468 (N_5468,N_5039,N_5151);
and U5469 (N_5469,N_5226,N_5055);
or U5470 (N_5470,N_5031,N_5220);
and U5471 (N_5471,N_5055,N_5234);
nor U5472 (N_5472,N_5153,N_5201);
nand U5473 (N_5473,N_5115,N_5099);
or U5474 (N_5474,N_5021,N_5216);
nor U5475 (N_5475,N_5128,N_5179);
or U5476 (N_5476,N_5032,N_5064);
or U5477 (N_5477,N_5192,N_5163);
or U5478 (N_5478,N_5181,N_5144);
nand U5479 (N_5479,N_5040,N_5191);
nand U5480 (N_5480,N_5081,N_5186);
and U5481 (N_5481,N_5092,N_5243);
and U5482 (N_5482,N_5159,N_5197);
or U5483 (N_5483,N_5026,N_5150);
nand U5484 (N_5484,N_5099,N_5225);
nand U5485 (N_5485,N_5058,N_5033);
and U5486 (N_5486,N_5228,N_5180);
nor U5487 (N_5487,N_5057,N_5142);
and U5488 (N_5488,N_5112,N_5162);
nand U5489 (N_5489,N_5208,N_5108);
or U5490 (N_5490,N_5081,N_5236);
nor U5491 (N_5491,N_5146,N_5161);
nand U5492 (N_5492,N_5136,N_5222);
xor U5493 (N_5493,N_5117,N_5180);
nor U5494 (N_5494,N_5243,N_5158);
and U5495 (N_5495,N_5237,N_5115);
or U5496 (N_5496,N_5069,N_5070);
nand U5497 (N_5497,N_5191,N_5238);
nor U5498 (N_5498,N_5061,N_5132);
nor U5499 (N_5499,N_5025,N_5174);
and U5500 (N_5500,N_5250,N_5381);
and U5501 (N_5501,N_5305,N_5266);
nor U5502 (N_5502,N_5499,N_5370);
and U5503 (N_5503,N_5409,N_5419);
or U5504 (N_5504,N_5449,N_5358);
nor U5505 (N_5505,N_5425,N_5487);
and U5506 (N_5506,N_5453,N_5447);
nor U5507 (N_5507,N_5377,N_5379);
and U5508 (N_5508,N_5495,N_5307);
and U5509 (N_5509,N_5461,N_5394);
nor U5510 (N_5510,N_5348,N_5433);
or U5511 (N_5511,N_5304,N_5411);
nand U5512 (N_5512,N_5300,N_5317);
xnor U5513 (N_5513,N_5363,N_5439);
or U5514 (N_5514,N_5260,N_5459);
nand U5515 (N_5515,N_5486,N_5391);
nor U5516 (N_5516,N_5410,N_5422);
nor U5517 (N_5517,N_5493,N_5268);
nand U5518 (N_5518,N_5415,N_5421);
and U5519 (N_5519,N_5265,N_5443);
or U5520 (N_5520,N_5445,N_5314);
nand U5521 (N_5521,N_5429,N_5401);
or U5522 (N_5522,N_5418,N_5452);
nand U5523 (N_5523,N_5367,N_5446);
or U5524 (N_5524,N_5286,N_5320);
or U5525 (N_5525,N_5389,N_5349);
and U5526 (N_5526,N_5273,N_5342);
nand U5527 (N_5527,N_5426,N_5364);
or U5528 (N_5528,N_5292,N_5492);
nand U5529 (N_5529,N_5489,N_5458);
nand U5530 (N_5530,N_5340,N_5472);
nor U5531 (N_5531,N_5413,N_5269);
nor U5532 (N_5532,N_5420,N_5442);
nor U5533 (N_5533,N_5466,N_5395);
or U5534 (N_5534,N_5339,N_5270);
nor U5535 (N_5535,N_5326,N_5297);
or U5536 (N_5536,N_5322,N_5276);
and U5537 (N_5537,N_5464,N_5319);
nand U5538 (N_5538,N_5456,N_5385);
nor U5539 (N_5539,N_5480,N_5479);
nor U5540 (N_5540,N_5295,N_5404);
or U5541 (N_5541,N_5325,N_5274);
and U5542 (N_5542,N_5259,N_5283);
or U5543 (N_5543,N_5428,N_5275);
and U5544 (N_5544,N_5468,N_5312);
nand U5545 (N_5545,N_5255,N_5465);
nor U5546 (N_5546,N_5457,N_5455);
nor U5547 (N_5547,N_5336,N_5288);
and U5548 (N_5548,N_5347,N_5403);
nand U5549 (N_5549,N_5316,N_5406);
and U5550 (N_5550,N_5359,N_5373);
nand U5551 (N_5551,N_5258,N_5460);
and U5552 (N_5552,N_5372,N_5328);
or U5553 (N_5553,N_5397,N_5343);
nand U5554 (N_5554,N_5463,N_5431);
and U5555 (N_5555,N_5400,N_5393);
or U5556 (N_5556,N_5263,N_5365);
or U5557 (N_5557,N_5306,N_5374);
nand U5558 (N_5558,N_5388,N_5285);
nand U5559 (N_5559,N_5416,N_5454);
nand U5560 (N_5560,N_5251,N_5462);
nor U5561 (N_5561,N_5301,N_5490);
nand U5562 (N_5562,N_5444,N_5488);
and U5563 (N_5563,N_5254,N_5256);
nor U5564 (N_5564,N_5396,N_5323);
and U5565 (N_5565,N_5272,N_5375);
nor U5566 (N_5566,N_5282,N_5337);
and U5567 (N_5567,N_5281,N_5277);
and U5568 (N_5568,N_5289,N_5354);
and U5569 (N_5569,N_5332,N_5484);
nand U5570 (N_5570,N_5369,N_5308);
nor U5571 (N_5571,N_5262,N_5423);
and U5572 (N_5572,N_5253,N_5334);
nand U5573 (N_5573,N_5296,N_5496);
or U5574 (N_5574,N_5310,N_5284);
and U5575 (N_5575,N_5384,N_5353);
and U5576 (N_5576,N_5318,N_5427);
or U5577 (N_5577,N_5346,N_5360);
or U5578 (N_5578,N_5405,N_5287);
nand U5579 (N_5579,N_5437,N_5441);
and U5580 (N_5580,N_5264,N_5478);
nor U5581 (N_5581,N_5473,N_5371);
or U5582 (N_5582,N_5430,N_5475);
nand U5583 (N_5583,N_5436,N_5414);
nor U5584 (N_5584,N_5257,N_5481);
nor U5585 (N_5585,N_5331,N_5376);
nor U5586 (N_5586,N_5378,N_5355);
nand U5587 (N_5587,N_5361,N_5344);
nor U5588 (N_5588,N_5327,N_5470);
and U5589 (N_5589,N_5280,N_5387);
nor U5590 (N_5590,N_5482,N_5380);
and U5591 (N_5591,N_5350,N_5483);
nand U5592 (N_5592,N_5345,N_5313);
nor U5593 (N_5593,N_5491,N_5356);
and U5594 (N_5594,N_5485,N_5278);
or U5595 (N_5595,N_5474,N_5290);
and U5596 (N_5596,N_5412,N_5335);
nand U5597 (N_5597,N_5351,N_5324);
and U5598 (N_5598,N_5338,N_5362);
nand U5599 (N_5599,N_5271,N_5329);
and U5600 (N_5600,N_5448,N_5498);
nor U5601 (N_5601,N_5279,N_5333);
nand U5602 (N_5602,N_5298,N_5471);
nor U5603 (N_5603,N_5311,N_5469);
or U5604 (N_5604,N_5451,N_5368);
nor U5605 (N_5605,N_5294,N_5467);
nor U5606 (N_5606,N_5252,N_5438);
nand U5607 (N_5607,N_5440,N_5267);
or U5608 (N_5608,N_5302,N_5450);
and U5609 (N_5609,N_5382,N_5386);
or U5610 (N_5610,N_5494,N_5293);
and U5611 (N_5611,N_5392,N_5299);
nand U5612 (N_5612,N_5407,N_5390);
or U5613 (N_5613,N_5497,N_5435);
or U5614 (N_5614,N_5303,N_5261);
nor U5615 (N_5615,N_5477,N_5309);
nor U5616 (N_5616,N_5352,N_5476);
nand U5617 (N_5617,N_5330,N_5434);
or U5618 (N_5618,N_5398,N_5383);
and U5619 (N_5619,N_5341,N_5357);
nand U5620 (N_5620,N_5432,N_5408);
nor U5621 (N_5621,N_5402,N_5315);
or U5622 (N_5622,N_5417,N_5399);
or U5623 (N_5623,N_5321,N_5424);
nor U5624 (N_5624,N_5366,N_5291);
and U5625 (N_5625,N_5350,N_5266);
and U5626 (N_5626,N_5287,N_5387);
nand U5627 (N_5627,N_5422,N_5255);
or U5628 (N_5628,N_5410,N_5427);
nor U5629 (N_5629,N_5298,N_5338);
nand U5630 (N_5630,N_5340,N_5285);
nand U5631 (N_5631,N_5417,N_5461);
and U5632 (N_5632,N_5490,N_5437);
nand U5633 (N_5633,N_5382,N_5366);
or U5634 (N_5634,N_5297,N_5408);
or U5635 (N_5635,N_5325,N_5470);
and U5636 (N_5636,N_5477,N_5479);
or U5637 (N_5637,N_5270,N_5345);
nand U5638 (N_5638,N_5420,N_5450);
or U5639 (N_5639,N_5371,N_5282);
nor U5640 (N_5640,N_5479,N_5274);
and U5641 (N_5641,N_5273,N_5332);
xor U5642 (N_5642,N_5489,N_5368);
nand U5643 (N_5643,N_5426,N_5475);
nor U5644 (N_5644,N_5434,N_5350);
and U5645 (N_5645,N_5378,N_5421);
and U5646 (N_5646,N_5315,N_5296);
and U5647 (N_5647,N_5268,N_5298);
and U5648 (N_5648,N_5346,N_5265);
or U5649 (N_5649,N_5312,N_5279);
or U5650 (N_5650,N_5493,N_5317);
or U5651 (N_5651,N_5365,N_5402);
nand U5652 (N_5652,N_5487,N_5370);
or U5653 (N_5653,N_5463,N_5279);
or U5654 (N_5654,N_5460,N_5423);
or U5655 (N_5655,N_5435,N_5324);
or U5656 (N_5656,N_5316,N_5381);
or U5657 (N_5657,N_5296,N_5417);
and U5658 (N_5658,N_5345,N_5394);
or U5659 (N_5659,N_5295,N_5417);
nor U5660 (N_5660,N_5256,N_5399);
or U5661 (N_5661,N_5294,N_5390);
nand U5662 (N_5662,N_5395,N_5402);
nand U5663 (N_5663,N_5431,N_5437);
nand U5664 (N_5664,N_5429,N_5426);
nand U5665 (N_5665,N_5496,N_5351);
or U5666 (N_5666,N_5308,N_5410);
nand U5667 (N_5667,N_5345,N_5285);
or U5668 (N_5668,N_5346,N_5405);
and U5669 (N_5669,N_5279,N_5406);
nand U5670 (N_5670,N_5327,N_5375);
nand U5671 (N_5671,N_5456,N_5257);
and U5672 (N_5672,N_5429,N_5330);
nor U5673 (N_5673,N_5431,N_5465);
nand U5674 (N_5674,N_5285,N_5387);
nand U5675 (N_5675,N_5289,N_5291);
nand U5676 (N_5676,N_5321,N_5367);
nor U5677 (N_5677,N_5421,N_5437);
nor U5678 (N_5678,N_5318,N_5404);
nand U5679 (N_5679,N_5338,N_5386);
or U5680 (N_5680,N_5328,N_5292);
nand U5681 (N_5681,N_5495,N_5385);
or U5682 (N_5682,N_5277,N_5434);
nand U5683 (N_5683,N_5250,N_5283);
nand U5684 (N_5684,N_5284,N_5352);
or U5685 (N_5685,N_5268,N_5338);
nor U5686 (N_5686,N_5405,N_5461);
or U5687 (N_5687,N_5314,N_5416);
nor U5688 (N_5688,N_5273,N_5282);
or U5689 (N_5689,N_5433,N_5490);
nor U5690 (N_5690,N_5297,N_5409);
nor U5691 (N_5691,N_5260,N_5487);
or U5692 (N_5692,N_5309,N_5308);
nand U5693 (N_5693,N_5427,N_5345);
nor U5694 (N_5694,N_5471,N_5250);
and U5695 (N_5695,N_5270,N_5395);
nand U5696 (N_5696,N_5369,N_5290);
nand U5697 (N_5697,N_5349,N_5393);
nor U5698 (N_5698,N_5347,N_5475);
nor U5699 (N_5699,N_5485,N_5269);
and U5700 (N_5700,N_5329,N_5256);
nor U5701 (N_5701,N_5485,N_5408);
or U5702 (N_5702,N_5383,N_5342);
and U5703 (N_5703,N_5351,N_5410);
nor U5704 (N_5704,N_5300,N_5354);
and U5705 (N_5705,N_5292,N_5403);
nor U5706 (N_5706,N_5289,N_5396);
and U5707 (N_5707,N_5417,N_5425);
and U5708 (N_5708,N_5497,N_5476);
nor U5709 (N_5709,N_5445,N_5272);
and U5710 (N_5710,N_5384,N_5428);
nand U5711 (N_5711,N_5450,N_5368);
and U5712 (N_5712,N_5279,N_5348);
or U5713 (N_5713,N_5471,N_5332);
and U5714 (N_5714,N_5366,N_5293);
nor U5715 (N_5715,N_5292,N_5376);
nand U5716 (N_5716,N_5349,N_5421);
nor U5717 (N_5717,N_5312,N_5330);
or U5718 (N_5718,N_5428,N_5298);
nor U5719 (N_5719,N_5266,N_5402);
nand U5720 (N_5720,N_5316,N_5351);
nor U5721 (N_5721,N_5315,N_5299);
or U5722 (N_5722,N_5410,N_5473);
nand U5723 (N_5723,N_5333,N_5346);
nor U5724 (N_5724,N_5338,N_5461);
or U5725 (N_5725,N_5383,N_5293);
and U5726 (N_5726,N_5334,N_5258);
nor U5727 (N_5727,N_5481,N_5451);
nor U5728 (N_5728,N_5287,N_5432);
nand U5729 (N_5729,N_5429,N_5300);
nand U5730 (N_5730,N_5493,N_5369);
or U5731 (N_5731,N_5479,N_5262);
nor U5732 (N_5732,N_5460,N_5370);
nor U5733 (N_5733,N_5430,N_5484);
and U5734 (N_5734,N_5496,N_5481);
and U5735 (N_5735,N_5368,N_5259);
nor U5736 (N_5736,N_5309,N_5368);
nand U5737 (N_5737,N_5385,N_5415);
nor U5738 (N_5738,N_5478,N_5366);
and U5739 (N_5739,N_5483,N_5438);
or U5740 (N_5740,N_5349,N_5377);
and U5741 (N_5741,N_5491,N_5353);
nand U5742 (N_5742,N_5293,N_5430);
nand U5743 (N_5743,N_5376,N_5425);
or U5744 (N_5744,N_5283,N_5464);
nand U5745 (N_5745,N_5309,N_5259);
nor U5746 (N_5746,N_5431,N_5305);
nor U5747 (N_5747,N_5455,N_5388);
or U5748 (N_5748,N_5496,N_5291);
nand U5749 (N_5749,N_5431,N_5356);
nand U5750 (N_5750,N_5647,N_5522);
nor U5751 (N_5751,N_5711,N_5531);
and U5752 (N_5752,N_5576,N_5582);
nor U5753 (N_5753,N_5651,N_5639);
nor U5754 (N_5754,N_5714,N_5657);
or U5755 (N_5755,N_5700,N_5743);
or U5756 (N_5756,N_5595,N_5593);
and U5757 (N_5757,N_5678,N_5554);
and U5758 (N_5758,N_5702,N_5506);
nand U5759 (N_5759,N_5697,N_5588);
nor U5760 (N_5760,N_5590,N_5517);
nand U5761 (N_5761,N_5514,N_5545);
nand U5762 (N_5762,N_5612,N_5656);
or U5763 (N_5763,N_5699,N_5726);
and U5764 (N_5764,N_5586,N_5694);
and U5765 (N_5765,N_5605,N_5601);
nor U5766 (N_5766,N_5616,N_5515);
and U5767 (N_5767,N_5630,N_5553);
or U5768 (N_5768,N_5672,N_5661);
and U5769 (N_5769,N_5730,N_5525);
nand U5770 (N_5770,N_5505,N_5716);
or U5771 (N_5771,N_5537,N_5544);
nand U5772 (N_5772,N_5589,N_5562);
nand U5773 (N_5773,N_5645,N_5653);
nor U5774 (N_5774,N_5655,N_5527);
nand U5775 (N_5775,N_5561,N_5611);
nor U5776 (N_5776,N_5592,N_5633);
xor U5777 (N_5777,N_5705,N_5691);
nand U5778 (N_5778,N_5523,N_5543);
or U5779 (N_5779,N_5568,N_5721);
nand U5780 (N_5780,N_5631,N_5646);
and U5781 (N_5781,N_5583,N_5731);
and U5782 (N_5782,N_5529,N_5629);
nor U5783 (N_5783,N_5689,N_5572);
and U5784 (N_5784,N_5680,N_5692);
or U5785 (N_5785,N_5548,N_5613);
and U5786 (N_5786,N_5737,N_5528);
or U5787 (N_5787,N_5650,N_5503);
and U5788 (N_5788,N_5677,N_5546);
nand U5789 (N_5789,N_5742,N_5557);
nor U5790 (N_5790,N_5728,N_5695);
and U5791 (N_5791,N_5564,N_5608);
nand U5792 (N_5792,N_5693,N_5539);
or U5793 (N_5793,N_5683,N_5644);
or U5794 (N_5794,N_5508,N_5634);
nand U5795 (N_5795,N_5674,N_5501);
and U5796 (N_5796,N_5635,N_5615);
or U5797 (N_5797,N_5690,N_5717);
or U5798 (N_5798,N_5641,N_5524);
and U5799 (N_5799,N_5602,N_5533);
and U5800 (N_5800,N_5587,N_5526);
or U5801 (N_5801,N_5547,N_5622);
nor U5802 (N_5802,N_5570,N_5624);
or U5803 (N_5803,N_5607,N_5504);
nor U5804 (N_5804,N_5735,N_5500);
nand U5805 (N_5805,N_5620,N_5549);
nor U5806 (N_5806,N_5706,N_5738);
or U5807 (N_5807,N_5625,N_5540);
nor U5808 (N_5808,N_5746,N_5687);
or U5809 (N_5809,N_5732,N_5667);
nor U5810 (N_5810,N_5676,N_5718);
nor U5811 (N_5811,N_5573,N_5575);
nor U5812 (N_5812,N_5555,N_5708);
nand U5813 (N_5813,N_5686,N_5623);
xnor U5814 (N_5814,N_5669,N_5679);
or U5815 (N_5815,N_5654,N_5671);
nand U5816 (N_5816,N_5560,N_5534);
and U5817 (N_5817,N_5556,N_5668);
nand U5818 (N_5818,N_5617,N_5532);
nor U5819 (N_5819,N_5518,N_5535);
nand U5820 (N_5820,N_5530,N_5739);
nand U5821 (N_5821,N_5720,N_5510);
or U5822 (N_5822,N_5642,N_5606);
nand U5823 (N_5823,N_5538,N_5591);
or U5824 (N_5824,N_5638,N_5727);
nand U5825 (N_5825,N_5599,N_5652);
nor U5826 (N_5826,N_5659,N_5621);
and U5827 (N_5827,N_5709,N_5675);
or U5828 (N_5828,N_5574,N_5609);
and U5829 (N_5829,N_5660,N_5596);
and U5830 (N_5830,N_5551,N_5744);
nand U5831 (N_5831,N_5600,N_5502);
and U5832 (N_5832,N_5640,N_5628);
nor U5833 (N_5833,N_5627,N_5729);
nor U5834 (N_5834,N_5724,N_5741);
nor U5835 (N_5835,N_5698,N_5666);
or U5836 (N_5836,N_5673,N_5703);
or U5837 (N_5837,N_5521,N_5585);
nor U5838 (N_5838,N_5567,N_5707);
and U5839 (N_5839,N_5748,N_5559);
or U5840 (N_5840,N_5519,N_5632);
nor U5841 (N_5841,N_5665,N_5662);
nor U5842 (N_5842,N_5619,N_5747);
nor U5843 (N_5843,N_5563,N_5719);
or U5844 (N_5844,N_5740,N_5701);
nand U5845 (N_5845,N_5636,N_5710);
nor U5846 (N_5846,N_5648,N_5663);
and U5847 (N_5847,N_5597,N_5542);
or U5848 (N_5848,N_5626,N_5618);
and U5849 (N_5849,N_5713,N_5658);
or U5850 (N_5850,N_5566,N_5664);
nor U5851 (N_5851,N_5581,N_5688);
or U5852 (N_5852,N_5685,N_5704);
nand U5853 (N_5853,N_5736,N_5614);
nor U5854 (N_5854,N_5511,N_5552);
nand U5855 (N_5855,N_5598,N_5745);
or U5856 (N_5856,N_5649,N_5513);
nor U5857 (N_5857,N_5594,N_5565);
nor U5858 (N_5858,N_5696,N_5684);
or U5859 (N_5859,N_5578,N_5509);
and U5860 (N_5860,N_5733,N_5670);
nor U5861 (N_5861,N_5584,N_5541);
nand U5862 (N_5862,N_5734,N_5579);
nand U5863 (N_5863,N_5682,N_5725);
nand U5864 (N_5864,N_5749,N_5643);
nand U5865 (N_5865,N_5571,N_5507);
nor U5866 (N_5866,N_5603,N_5516);
nor U5867 (N_5867,N_5681,N_5712);
nor U5868 (N_5868,N_5604,N_5520);
and U5869 (N_5869,N_5580,N_5550);
and U5870 (N_5870,N_5610,N_5577);
and U5871 (N_5871,N_5536,N_5715);
or U5872 (N_5872,N_5512,N_5569);
nand U5873 (N_5873,N_5558,N_5723);
or U5874 (N_5874,N_5637,N_5722);
or U5875 (N_5875,N_5577,N_5661);
or U5876 (N_5876,N_5613,N_5641);
nand U5877 (N_5877,N_5665,N_5611);
nor U5878 (N_5878,N_5610,N_5639);
nand U5879 (N_5879,N_5607,N_5667);
or U5880 (N_5880,N_5577,N_5549);
or U5881 (N_5881,N_5591,N_5540);
or U5882 (N_5882,N_5535,N_5524);
or U5883 (N_5883,N_5504,N_5659);
nor U5884 (N_5884,N_5738,N_5560);
nand U5885 (N_5885,N_5527,N_5540);
and U5886 (N_5886,N_5616,N_5730);
and U5887 (N_5887,N_5504,N_5623);
and U5888 (N_5888,N_5549,N_5748);
nand U5889 (N_5889,N_5643,N_5642);
nand U5890 (N_5890,N_5625,N_5704);
xnor U5891 (N_5891,N_5690,N_5510);
and U5892 (N_5892,N_5547,N_5669);
nand U5893 (N_5893,N_5549,N_5504);
nand U5894 (N_5894,N_5644,N_5669);
nor U5895 (N_5895,N_5581,N_5503);
and U5896 (N_5896,N_5739,N_5685);
nor U5897 (N_5897,N_5520,N_5651);
nor U5898 (N_5898,N_5631,N_5686);
and U5899 (N_5899,N_5711,N_5559);
or U5900 (N_5900,N_5598,N_5704);
nor U5901 (N_5901,N_5700,N_5614);
or U5902 (N_5902,N_5634,N_5641);
or U5903 (N_5903,N_5634,N_5542);
nor U5904 (N_5904,N_5595,N_5665);
nand U5905 (N_5905,N_5703,N_5526);
nor U5906 (N_5906,N_5730,N_5675);
or U5907 (N_5907,N_5649,N_5736);
nor U5908 (N_5908,N_5679,N_5711);
and U5909 (N_5909,N_5621,N_5642);
nor U5910 (N_5910,N_5562,N_5687);
and U5911 (N_5911,N_5502,N_5625);
nand U5912 (N_5912,N_5575,N_5666);
nand U5913 (N_5913,N_5679,N_5545);
nand U5914 (N_5914,N_5718,N_5638);
and U5915 (N_5915,N_5558,N_5514);
nand U5916 (N_5916,N_5585,N_5616);
nor U5917 (N_5917,N_5741,N_5557);
nand U5918 (N_5918,N_5517,N_5725);
nand U5919 (N_5919,N_5673,N_5666);
nand U5920 (N_5920,N_5679,N_5712);
nand U5921 (N_5921,N_5711,N_5601);
or U5922 (N_5922,N_5549,N_5714);
or U5923 (N_5923,N_5575,N_5528);
nor U5924 (N_5924,N_5634,N_5541);
nand U5925 (N_5925,N_5555,N_5512);
or U5926 (N_5926,N_5746,N_5674);
nor U5927 (N_5927,N_5749,N_5698);
and U5928 (N_5928,N_5574,N_5713);
nor U5929 (N_5929,N_5546,N_5641);
nand U5930 (N_5930,N_5686,N_5661);
nand U5931 (N_5931,N_5656,N_5719);
and U5932 (N_5932,N_5589,N_5685);
nor U5933 (N_5933,N_5534,N_5555);
nand U5934 (N_5934,N_5666,N_5606);
nor U5935 (N_5935,N_5536,N_5562);
nor U5936 (N_5936,N_5526,N_5592);
or U5937 (N_5937,N_5614,N_5726);
nand U5938 (N_5938,N_5562,N_5685);
or U5939 (N_5939,N_5701,N_5535);
or U5940 (N_5940,N_5681,N_5705);
nor U5941 (N_5941,N_5571,N_5575);
and U5942 (N_5942,N_5586,N_5557);
nand U5943 (N_5943,N_5646,N_5540);
nor U5944 (N_5944,N_5734,N_5635);
nor U5945 (N_5945,N_5564,N_5607);
nand U5946 (N_5946,N_5517,N_5510);
and U5947 (N_5947,N_5514,N_5580);
nor U5948 (N_5948,N_5593,N_5611);
or U5949 (N_5949,N_5636,N_5560);
nand U5950 (N_5950,N_5538,N_5732);
nand U5951 (N_5951,N_5637,N_5697);
and U5952 (N_5952,N_5696,N_5520);
nand U5953 (N_5953,N_5727,N_5736);
nor U5954 (N_5954,N_5740,N_5603);
and U5955 (N_5955,N_5660,N_5521);
nor U5956 (N_5956,N_5545,N_5579);
nand U5957 (N_5957,N_5672,N_5526);
nand U5958 (N_5958,N_5516,N_5730);
and U5959 (N_5959,N_5539,N_5547);
nor U5960 (N_5960,N_5553,N_5595);
nand U5961 (N_5961,N_5633,N_5659);
nand U5962 (N_5962,N_5556,N_5728);
and U5963 (N_5963,N_5747,N_5680);
and U5964 (N_5964,N_5606,N_5646);
nand U5965 (N_5965,N_5534,N_5612);
nand U5966 (N_5966,N_5631,N_5589);
nor U5967 (N_5967,N_5693,N_5743);
nand U5968 (N_5968,N_5610,N_5657);
nor U5969 (N_5969,N_5618,N_5595);
and U5970 (N_5970,N_5617,N_5713);
nor U5971 (N_5971,N_5696,N_5507);
and U5972 (N_5972,N_5583,N_5538);
nor U5973 (N_5973,N_5730,N_5570);
nor U5974 (N_5974,N_5636,N_5717);
nor U5975 (N_5975,N_5735,N_5699);
nand U5976 (N_5976,N_5654,N_5667);
nor U5977 (N_5977,N_5551,N_5656);
nor U5978 (N_5978,N_5617,N_5529);
nor U5979 (N_5979,N_5525,N_5627);
or U5980 (N_5980,N_5624,N_5734);
nand U5981 (N_5981,N_5547,N_5568);
and U5982 (N_5982,N_5511,N_5526);
nand U5983 (N_5983,N_5580,N_5512);
and U5984 (N_5984,N_5718,N_5679);
xnor U5985 (N_5985,N_5747,N_5631);
nor U5986 (N_5986,N_5702,N_5612);
nor U5987 (N_5987,N_5505,N_5513);
and U5988 (N_5988,N_5616,N_5674);
nor U5989 (N_5989,N_5670,N_5612);
and U5990 (N_5990,N_5662,N_5595);
and U5991 (N_5991,N_5695,N_5571);
nor U5992 (N_5992,N_5587,N_5628);
nor U5993 (N_5993,N_5500,N_5608);
nor U5994 (N_5994,N_5737,N_5600);
nor U5995 (N_5995,N_5505,N_5595);
and U5996 (N_5996,N_5683,N_5515);
nor U5997 (N_5997,N_5625,N_5684);
nand U5998 (N_5998,N_5690,N_5556);
or U5999 (N_5999,N_5589,N_5564);
or U6000 (N_6000,N_5804,N_5892);
xor U6001 (N_6001,N_5881,N_5763);
nand U6002 (N_6002,N_5931,N_5983);
and U6003 (N_6003,N_5995,N_5758);
and U6004 (N_6004,N_5962,N_5832);
and U6005 (N_6005,N_5996,N_5753);
nand U6006 (N_6006,N_5992,N_5954);
or U6007 (N_6007,N_5999,N_5915);
or U6008 (N_6008,N_5961,N_5784);
and U6009 (N_6009,N_5979,N_5938);
nand U6010 (N_6010,N_5880,N_5842);
or U6011 (N_6011,N_5792,N_5887);
and U6012 (N_6012,N_5821,N_5827);
nor U6013 (N_6013,N_5928,N_5893);
or U6014 (N_6014,N_5861,N_5933);
or U6015 (N_6015,N_5815,N_5754);
and U6016 (N_6016,N_5896,N_5799);
and U6017 (N_6017,N_5762,N_5869);
and U6018 (N_6018,N_5910,N_5774);
or U6019 (N_6019,N_5994,N_5820);
nand U6020 (N_6020,N_5872,N_5850);
xor U6021 (N_6021,N_5908,N_5889);
or U6022 (N_6022,N_5807,N_5845);
nor U6023 (N_6023,N_5855,N_5953);
nor U6024 (N_6024,N_5858,N_5773);
and U6025 (N_6025,N_5835,N_5787);
nand U6026 (N_6026,N_5822,N_5756);
and U6027 (N_6027,N_5883,N_5897);
and U6028 (N_6028,N_5851,N_5932);
nor U6029 (N_6029,N_5806,N_5919);
nor U6030 (N_6030,N_5975,N_5761);
nor U6031 (N_6031,N_5906,N_5970);
xor U6032 (N_6032,N_5788,N_5865);
nor U6033 (N_6033,N_5768,N_5884);
and U6034 (N_6034,N_5830,N_5843);
nor U6035 (N_6035,N_5966,N_5789);
and U6036 (N_6036,N_5902,N_5952);
nand U6037 (N_6037,N_5793,N_5885);
nor U6038 (N_6038,N_5967,N_5790);
or U6039 (N_6039,N_5907,N_5987);
nor U6040 (N_6040,N_5779,N_5819);
and U6041 (N_6041,N_5947,N_5782);
nand U6042 (N_6042,N_5825,N_5911);
and U6043 (N_6043,N_5873,N_5755);
and U6044 (N_6044,N_5760,N_5847);
nand U6045 (N_6045,N_5963,N_5921);
nor U6046 (N_6046,N_5844,N_5795);
or U6047 (N_6047,N_5859,N_5955);
or U6048 (N_6048,N_5904,N_5991);
or U6049 (N_6049,N_5759,N_5870);
and U6050 (N_6050,N_5917,N_5837);
nand U6051 (N_6051,N_5794,N_5791);
nand U6052 (N_6052,N_5934,N_5778);
nand U6053 (N_6053,N_5866,N_5882);
and U6054 (N_6054,N_5848,N_5803);
xnor U6055 (N_6055,N_5752,N_5985);
or U6056 (N_6056,N_5783,N_5964);
or U6057 (N_6057,N_5800,N_5875);
and U6058 (N_6058,N_5998,N_5831);
or U6059 (N_6059,N_5940,N_5960);
nor U6060 (N_6060,N_5878,N_5901);
and U6061 (N_6061,N_5863,N_5909);
or U6062 (N_6062,N_5856,N_5988);
nand U6063 (N_6063,N_5945,N_5939);
nand U6064 (N_6064,N_5879,N_5854);
nand U6065 (N_6065,N_5974,N_5786);
and U6066 (N_6066,N_5944,N_5886);
nor U6067 (N_6067,N_5809,N_5898);
or U6068 (N_6068,N_5982,N_5853);
or U6069 (N_6069,N_5929,N_5905);
and U6070 (N_6070,N_5968,N_5922);
nand U6071 (N_6071,N_5834,N_5775);
or U6072 (N_6072,N_5770,N_5972);
nor U6073 (N_6073,N_5984,N_5941);
and U6074 (N_6074,N_5918,N_5958);
nand U6075 (N_6075,N_5813,N_5950);
nor U6076 (N_6076,N_5937,N_5757);
nand U6077 (N_6077,N_5969,N_5816);
or U6078 (N_6078,N_5942,N_5891);
nand U6079 (N_6079,N_5797,N_5899);
nand U6080 (N_6080,N_5777,N_5924);
or U6081 (N_6081,N_5903,N_5976);
or U6082 (N_6082,N_5956,N_5798);
nor U6083 (N_6083,N_5936,N_5767);
or U6084 (N_6084,N_5838,N_5890);
and U6085 (N_6085,N_5867,N_5895);
nand U6086 (N_6086,N_5852,N_5860);
nand U6087 (N_6087,N_5776,N_5957);
nand U6088 (N_6088,N_5833,N_5841);
and U6089 (N_6089,N_5888,N_5930);
and U6090 (N_6090,N_5993,N_5814);
or U6091 (N_6091,N_5949,N_5874);
nand U6092 (N_6092,N_5959,N_5971);
and U6093 (N_6093,N_5780,N_5925);
nand U6094 (N_6094,N_5801,N_5810);
nor U6095 (N_6095,N_5785,N_5965);
nand U6096 (N_6096,N_5868,N_5823);
nor U6097 (N_6097,N_5764,N_5923);
and U6098 (N_6098,N_5990,N_5840);
nand U6099 (N_6099,N_5828,N_5876);
and U6100 (N_6100,N_5916,N_5818);
nand U6101 (N_6101,N_5751,N_5977);
nand U6102 (N_6102,N_5771,N_5951);
nand U6103 (N_6103,N_5920,N_5948);
and U6104 (N_6104,N_5981,N_5912);
nor U6105 (N_6105,N_5864,N_5914);
and U6106 (N_6106,N_5772,N_5769);
nand U6107 (N_6107,N_5849,N_5817);
or U6108 (N_6108,N_5824,N_5894);
or U6109 (N_6109,N_5836,N_5808);
or U6110 (N_6110,N_5900,N_5811);
and U6111 (N_6111,N_5750,N_5826);
nor U6112 (N_6112,N_5812,N_5877);
nand U6113 (N_6113,N_5997,N_5926);
or U6114 (N_6114,N_5946,N_5978);
nand U6115 (N_6115,N_5935,N_5973);
or U6116 (N_6116,N_5989,N_5871);
nor U6117 (N_6117,N_5846,N_5805);
xnor U6118 (N_6118,N_5796,N_5857);
nand U6119 (N_6119,N_5839,N_5913);
or U6120 (N_6120,N_5829,N_5927);
nor U6121 (N_6121,N_5781,N_5802);
nor U6122 (N_6122,N_5766,N_5943);
nor U6123 (N_6123,N_5980,N_5986);
and U6124 (N_6124,N_5765,N_5862);
nand U6125 (N_6125,N_5992,N_5893);
nor U6126 (N_6126,N_5958,N_5945);
and U6127 (N_6127,N_5882,N_5967);
and U6128 (N_6128,N_5820,N_5827);
nor U6129 (N_6129,N_5931,N_5771);
and U6130 (N_6130,N_5894,N_5853);
nand U6131 (N_6131,N_5792,N_5901);
nor U6132 (N_6132,N_5816,N_5960);
nor U6133 (N_6133,N_5932,N_5783);
and U6134 (N_6134,N_5807,N_5753);
nand U6135 (N_6135,N_5958,N_5857);
nor U6136 (N_6136,N_5841,N_5840);
nor U6137 (N_6137,N_5837,N_5899);
nand U6138 (N_6138,N_5942,N_5961);
nand U6139 (N_6139,N_5898,N_5865);
and U6140 (N_6140,N_5750,N_5909);
nand U6141 (N_6141,N_5932,N_5876);
nor U6142 (N_6142,N_5827,N_5939);
and U6143 (N_6143,N_5881,N_5849);
nand U6144 (N_6144,N_5867,N_5816);
or U6145 (N_6145,N_5828,N_5924);
or U6146 (N_6146,N_5985,N_5932);
and U6147 (N_6147,N_5992,N_5920);
or U6148 (N_6148,N_5816,N_5998);
nand U6149 (N_6149,N_5807,N_5969);
or U6150 (N_6150,N_5919,N_5927);
nor U6151 (N_6151,N_5871,N_5921);
or U6152 (N_6152,N_5890,N_5778);
nor U6153 (N_6153,N_5781,N_5832);
nand U6154 (N_6154,N_5952,N_5997);
nand U6155 (N_6155,N_5758,N_5832);
nor U6156 (N_6156,N_5893,N_5790);
nor U6157 (N_6157,N_5818,N_5836);
or U6158 (N_6158,N_5957,N_5775);
and U6159 (N_6159,N_5861,N_5955);
nand U6160 (N_6160,N_5804,N_5854);
nand U6161 (N_6161,N_5889,N_5795);
or U6162 (N_6162,N_5871,N_5906);
or U6163 (N_6163,N_5920,N_5898);
or U6164 (N_6164,N_5866,N_5873);
and U6165 (N_6165,N_5808,N_5759);
nand U6166 (N_6166,N_5807,N_5868);
nor U6167 (N_6167,N_5807,N_5818);
and U6168 (N_6168,N_5974,N_5994);
or U6169 (N_6169,N_5903,N_5808);
and U6170 (N_6170,N_5810,N_5916);
and U6171 (N_6171,N_5981,N_5773);
or U6172 (N_6172,N_5854,N_5770);
nand U6173 (N_6173,N_5830,N_5942);
nand U6174 (N_6174,N_5916,N_5921);
nand U6175 (N_6175,N_5900,N_5844);
or U6176 (N_6176,N_5993,N_5802);
nand U6177 (N_6177,N_5825,N_5879);
nand U6178 (N_6178,N_5918,N_5861);
and U6179 (N_6179,N_5837,N_5977);
nand U6180 (N_6180,N_5973,N_5946);
xnor U6181 (N_6181,N_5899,N_5936);
nand U6182 (N_6182,N_5869,N_5764);
nor U6183 (N_6183,N_5909,N_5814);
nand U6184 (N_6184,N_5826,N_5813);
and U6185 (N_6185,N_5926,N_5899);
and U6186 (N_6186,N_5751,N_5750);
and U6187 (N_6187,N_5780,N_5765);
nor U6188 (N_6188,N_5878,N_5864);
and U6189 (N_6189,N_5840,N_5765);
and U6190 (N_6190,N_5841,N_5838);
nand U6191 (N_6191,N_5902,N_5780);
nand U6192 (N_6192,N_5824,N_5872);
nor U6193 (N_6193,N_5878,N_5757);
and U6194 (N_6194,N_5986,N_5828);
nor U6195 (N_6195,N_5804,N_5945);
nand U6196 (N_6196,N_5750,N_5857);
and U6197 (N_6197,N_5948,N_5817);
nand U6198 (N_6198,N_5828,N_5989);
or U6199 (N_6199,N_5765,N_5899);
and U6200 (N_6200,N_5953,N_5762);
nor U6201 (N_6201,N_5926,N_5919);
nand U6202 (N_6202,N_5771,N_5862);
nand U6203 (N_6203,N_5825,N_5823);
nand U6204 (N_6204,N_5838,N_5786);
nor U6205 (N_6205,N_5953,N_5905);
nand U6206 (N_6206,N_5867,N_5906);
xor U6207 (N_6207,N_5848,N_5938);
nor U6208 (N_6208,N_5777,N_5870);
nor U6209 (N_6209,N_5930,N_5830);
or U6210 (N_6210,N_5780,N_5766);
nor U6211 (N_6211,N_5795,N_5977);
and U6212 (N_6212,N_5820,N_5963);
nor U6213 (N_6213,N_5843,N_5752);
or U6214 (N_6214,N_5845,N_5961);
or U6215 (N_6215,N_5799,N_5882);
nor U6216 (N_6216,N_5940,N_5782);
or U6217 (N_6217,N_5964,N_5823);
and U6218 (N_6218,N_5988,N_5862);
or U6219 (N_6219,N_5936,N_5996);
or U6220 (N_6220,N_5786,N_5985);
and U6221 (N_6221,N_5934,N_5921);
and U6222 (N_6222,N_5804,N_5765);
nand U6223 (N_6223,N_5935,N_5925);
and U6224 (N_6224,N_5857,N_5992);
or U6225 (N_6225,N_5918,N_5950);
and U6226 (N_6226,N_5881,N_5987);
nor U6227 (N_6227,N_5789,N_5808);
or U6228 (N_6228,N_5803,N_5818);
nand U6229 (N_6229,N_5917,N_5961);
or U6230 (N_6230,N_5872,N_5888);
nand U6231 (N_6231,N_5976,N_5918);
or U6232 (N_6232,N_5754,N_5938);
nand U6233 (N_6233,N_5834,N_5810);
nor U6234 (N_6234,N_5821,N_5826);
nor U6235 (N_6235,N_5765,N_5822);
nor U6236 (N_6236,N_5854,N_5764);
nor U6237 (N_6237,N_5945,N_5920);
nand U6238 (N_6238,N_5868,N_5787);
or U6239 (N_6239,N_5771,N_5789);
and U6240 (N_6240,N_5959,N_5878);
nor U6241 (N_6241,N_5825,N_5898);
nand U6242 (N_6242,N_5846,N_5894);
nand U6243 (N_6243,N_5936,N_5902);
nor U6244 (N_6244,N_5999,N_5860);
or U6245 (N_6245,N_5927,N_5844);
and U6246 (N_6246,N_5934,N_5789);
nand U6247 (N_6247,N_5941,N_5977);
nor U6248 (N_6248,N_5882,N_5831);
nor U6249 (N_6249,N_5886,N_5906);
nand U6250 (N_6250,N_6210,N_6211);
or U6251 (N_6251,N_6154,N_6179);
and U6252 (N_6252,N_6164,N_6085);
nand U6253 (N_6253,N_6066,N_6076);
or U6254 (N_6254,N_6081,N_6220);
or U6255 (N_6255,N_6141,N_6244);
or U6256 (N_6256,N_6124,N_6065);
nor U6257 (N_6257,N_6127,N_6032);
nand U6258 (N_6258,N_6194,N_6005);
nand U6259 (N_6259,N_6018,N_6185);
or U6260 (N_6260,N_6083,N_6198);
nand U6261 (N_6261,N_6174,N_6205);
or U6262 (N_6262,N_6117,N_6017);
or U6263 (N_6263,N_6231,N_6110);
nor U6264 (N_6264,N_6126,N_6043);
nor U6265 (N_6265,N_6125,N_6193);
and U6266 (N_6266,N_6173,N_6049);
nand U6267 (N_6267,N_6213,N_6138);
or U6268 (N_6268,N_6040,N_6008);
nand U6269 (N_6269,N_6137,N_6200);
nand U6270 (N_6270,N_6218,N_6063);
and U6271 (N_6271,N_6191,N_6216);
nor U6272 (N_6272,N_6132,N_6229);
nor U6273 (N_6273,N_6007,N_6190);
and U6274 (N_6274,N_6109,N_6222);
or U6275 (N_6275,N_6009,N_6012);
nand U6276 (N_6276,N_6036,N_6054);
nand U6277 (N_6277,N_6115,N_6037);
nor U6278 (N_6278,N_6170,N_6055);
and U6279 (N_6279,N_6142,N_6071);
or U6280 (N_6280,N_6165,N_6230);
and U6281 (N_6281,N_6177,N_6228);
or U6282 (N_6282,N_6241,N_6082);
nor U6283 (N_6283,N_6099,N_6148);
and U6284 (N_6284,N_6143,N_6105);
nand U6285 (N_6285,N_6070,N_6206);
nor U6286 (N_6286,N_6161,N_6106);
nor U6287 (N_6287,N_6225,N_6038);
or U6288 (N_6288,N_6239,N_6006);
nand U6289 (N_6289,N_6156,N_6059);
nand U6290 (N_6290,N_6157,N_6107);
nand U6291 (N_6291,N_6031,N_6045);
or U6292 (N_6292,N_6175,N_6204);
or U6293 (N_6293,N_6247,N_6217);
nor U6294 (N_6294,N_6022,N_6183);
nand U6295 (N_6295,N_6145,N_6118);
nand U6296 (N_6296,N_6245,N_6015);
nor U6297 (N_6297,N_6176,N_6025);
xnor U6298 (N_6298,N_6130,N_6069);
nor U6299 (N_6299,N_6016,N_6114);
nor U6300 (N_6300,N_6122,N_6086);
and U6301 (N_6301,N_6238,N_6098);
nand U6302 (N_6302,N_6075,N_6196);
nand U6303 (N_6303,N_6046,N_6112);
nor U6304 (N_6304,N_6027,N_6167);
nor U6305 (N_6305,N_6095,N_6158);
nand U6306 (N_6306,N_6020,N_6003);
or U6307 (N_6307,N_6101,N_6026);
nand U6308 (N_6308,N_6236,N_6197);
and U6309 (N_6309,N_6226,N_6062);
nand U6310 (N_6310,N_6171,N_6068);
and U6311 (N_6311,N_6094,N_6155);
or U6312 (N_6312,N_6052,N_6084);
nor U6313 (N_6313,N_6151,N_6030);
and U6314 (N_6314,N_6004,N_6203);
nor U6315 (N_6315,N_6144,N_6188);
or U6316 (N_6316,N_6235,N_6093);
nor U6317 (N_6317,N_6123,N_6134);
nor U6318 (N_6318,N_6088,N_6240);
nor U6319 (N_6319,N_6202,N_6140);
and U6320 (N_6320,N_6146,N_6195);
and U6321 (N_6321,N_6135,N_6139);
nor U6322 (N_6322,N_6061,N_6047);
nor U6323 (N_6323,N_6136,N_6149);
or U6324 (N_6324,N_6091,N_6078);
and U6325 (N_6325,N_6249,N_6248);
nor U6326 (N_6326,N_6207,N_6182);
and U6327 (N_6327,N_6057,N_6067);
and U6328 (N_6328,N_6237,N_6242);
or U6329 (N_6329,N_6000,N_6187);
nor U6330 (N_6330,N_6100,N_6234);
nand U6331 (N_6331,N_6064,N_6212);
nand U6332 (N_6332,N_6192,N_6189);
and U6333 (N_6333,N_6060,N_6219);
nand U6334 (N_6334,N_6221,N_6172);
nand U6335 (N_6335,N_6050,N_6131);
nand U6336 (N_6336,N_6181,N_6111);
nor U6337 (N_6337,N_6199,N_6224);
nand U6338 (N_6338,N_6053,N_6024);
nand U6339 (N_6339,N_6133,N_6090);
or U6340 (N_6340,N_6058,N_6034);
nor U6341 (N_6341,N_6201,N_6243);
and U6342 (N_6342,N_6041,N_6214);
nor U6343 (N_6343,N_6232,N_6180);
and U6344 (N_6344,N_6014,N_6169);
nor U6345 (N_6345,N_6023,N_6233);
nor U6346 (N_6346,N_6087,N_6092);
or U6347 (N_6347,N_6178,N_6010);
nor U6348 (N_6348,N_6162,N_6089);
or U6349 (N_6349,N_6186,N_6150);
nor U6350 (N_6350,N_6035,N_6223);
or U6351 (N_6351,N_6044,N_6184);
or U6352 (N_6352,N_6042,N_6056);
nand U6353 (N_6353,N_6128,N_6159);
and U6354 (N_6354,N_6227,N_6048);
nand U6355 (N_6355,N_6119,N_6152);
nor U6356 (N_6356,N_6096,N_6097);
nand U6357 (N_6357,N_6074,N_6013);
or U6358 (N_6358,N_6147,N_6113);
and U6359 (N_6359,N_6163,N_6153);
or U6360 (N_6360,N_6120,N_6011);
nand U6361 (N_6361,N_6080,N_6001);
nand U6362 (N_6362,N_6209,N_6208);
and U6363 (N_6363,N_6021,N_6039);
or U6364 (N_6364,N_6129,N_6077);
nor U6365 (N_6365,N_6079,N_6160);
nand U6366 (N_6366,N_6029,N_6073);
nand U6367 (N_6367,N_6033,N_6108);
nand U6368 (N_6368,N_6116,N_6072);
and U6369 (N_6369,N_6102,N_6002);
and U6370 (N_6370,N_6103,N_6246);
nand U6371 (N_6371,N_6121,N_6168);
or U6372 (N_6372,N_6215,N_6051);
nor U6373 (N_6373,N_6028,N_6166);
nand U6374 (N_6374,N_6104,N_6019);
nand U6375 (N_6375,N_6202,N_6032);
nand U6376 (N_6376,N_6011,N_6000);
nand U6377 (N_6377,N_6230,N_6059);
nor U6378 (N_6378,N_6141,N_6229);
nor U6379 (N_6379,N_6119,N_6076);
nand U6380 (N_6380,N_6187,N_6061);
nor U6381 (N_6381,N_6157,N_6009);
nand U6382 (N_6382,N_6248,N_6075);
nand U6383 (N_6383,N_6243,N_6168);
and U6384 (N_6384,N_6195,N_6170);
nand U6385 (N_6385,N_6232,N_6041);
nand U6386 (N_6386,N_6212,N_6100);
and U6387 (N_6387,N_6177,N_6055);
nor U6388 (N_6388,N_6099,N_6137);
nand U6389 (N_6389,N_6018,N_6030);
and U6390 (N_6390,N_6125,N_6132);
or U6391 (N_6391,N_6140,N_6023);
nand U6392 (N_6392,N_6106,N_6159);
xor U6393 (N_6393,N_6205,N_6194);
and U6394 (N_6394,N_6091,N_6109);
nand U6395 (N_6395,N_6028,N_6053);
nor U6396 (N_6396,N_6047,N_6189);
nor U6397 (N_6397,N_6183,N_6162);
and U6398 (N_6398,N_6220,N_6113);
nand U6399 (N_6399,N_6100,N_6079);
or U6400 (N_6400,N_6144,N_6108);
and U6401 (N_6401,N_6006,N_6030);
nand U6402 (N_6402,N_6138,N_6199);
and U6403 (N_6403,N_6210,N_6104);
nand U6404 (N_6404,N_6007,N_6078);
nand U6405 (N_6405,N_6067,N_6111);
nand U6406 (N_6406,N_6188,N_6077);
and U6407 (N_6407,N_6155,N_6213);
and U6408 (N_6408,N_6115,N_6137);
nor U6409 (N_6409,N_6213,N_6034);
nand U6410 (N_6410,N_6110,N_6085);
nand U6411 (N_6411,N_6017,N_6025);
nor U6412 (N_6412,N_6104,N_6009);
and U6413 (N_6413,N_6225,N_6192);
or U6414 (N_6414,N_6028,N_6021);
nor U6415 (N_6415,N_6037,N_6001);
nor U6416 (N_6416,N_6002,N_6066);
and U6417 (N_6417,N_6101,N_6141);
or U6418 (N_6418,N_6120,N_6012);
nor U6419 (N_6419,N_6225,N_6128);
or U6420 (N_6420,N_6094,N_6185);
or U6421 (N_6421,N_6152,N_6142);
nor U6422 (N_6422,N_6172,N_6242);
and U6423 (N_6423,N_6032,N_6087);
nand U6424 (N_6424,N_6071,N_6115);
or U6425 (N_6425,N_6033,N_6161);
and U6426 (N_6426,N_6170,N_6119);
nand U6427 (N_6427,N_6097,N_6086);
nor U6428 (N_6428,N_6183,N_6249);
nand U6429 (N_6429,N_6201,N_6160);
and U6430 (N_6430,N_6238,N_6074);
and U6431 (N_6431,N_6131,N_6091);
nand U6432 (N_6432,N_6000,N_6093);
and U6433 (N_6433,N_6045,N_6034);
nor U6434 (N_6434,N_6231,N_6062);
nand U6435 (N_6435,N_6005,N_6140);
and U6436 (N_6436,N_6213,N_6122);
and U6437 (N_6437,N_6220,N_6030);
nand U6438 (N_6438,N_6073,N_6009);
nor U6439 (N_6439,N_6011,N_6224);
nand U6440 (N_6440,N_6091,N_6158);
and U6441 (N_6441,N_6249,N_6075);
nor U6442 (N_6442,N_6170,N_6081);
nor U6443 (N_6443,N_6246,N_6159);
or U6444 (N_6444,N_6234,N_6095);
nand U6445 (N_6445,N_6083,N_6163);
or U6446 (N_6446,N_6163,N_6178);
or U6447 (N_6447,N_6126,N_6052);
and U6448 (N_6448,N_6071,N_6057);
nand U6449 (N_6449,N_6223,N_6190);
and U6450 (N_6450,N_6107,N_6020);
nand U6451 (N_6451,N_6188,N_6091);
or U6452 (N_6452,N_6209,N_6013);
or U6453 (N_6453,N_6119,N_6166);
or U6454 (N_6454,N_6070,N_6199);
or U6455 (N_6455,N_6077,N_6235);
nor U6456 (N_6456,N_6192,N_6158);
xor U6457 (N_6457,N_6184,N_6133);
nand U6458 (N_6458,N_6167,N_6159);
or U6459 (N_6459,N_6096,N_6163);
or U6460 (N_6460,N_6106,N_6062);
or U6461 (N_6461,N_6034,N_6062);
or U6462 (N_6462,N_6153,N_6087);
nor U6463 (N_6463,N_6107,N_6004);
or U6464 (N_6464,N_6216,N_6046);
nor U6465 (N_6465,N_6081,N_6248);
or U6466 (N_6466,N_6144,N_6237);
nor U6467 (N_6467,N_6045,N_6000);
or U6468 (N_6468,N_6201,N_6075);
nand U6469 (N_6469,N_6050,N_6116);
xnor U6470 (N_6470,N_6034,N_6018);
nand U6471 (N_6471,N_6122,N_6248);
nand U6472 (N_6472,N_6042,N_6234);
and U6473 (N_6473,N_6013,N_6055);
and U6474 (N_6474,N_6050,N_6071);
xnor U6475 (N_6475,N_6080,N_6046);
nand U6476 (N_6476,N_6102,N_6039);
or U6477 (N_6477,N_6090,N_6004);
nor U6478 (N_6478,N_6150,N_6107);
or U6479 (N_6479,N_6185,N_6121);
or U6480 (N_6480,N_6231,N_6187);
nor U6481 (N_6481,N_6015,N_6089);
nand U6482 (N_6482,N_6188,N_6153);
xnor U6483 (N_6483,N_6013,N_6185);
nor U6484 (N_6484,N_6234,N_6046);
nand U6485 (N_6485,N_6130,N_6101);
and U6486 (N_6486,N_6126,N_6166);
nand U6487 (N_6487,N_6199,N_6051);
nand U6488 (N_6488,N_6140,N_6075);
nand U6489 (N_6489,N_6234,N_6178);
nor U6490 (N_6490,N_6227,N_6168);
nand U6491 (N_6491,N_6206,N_6143);
nor U6492 (N_6492,N_6075,N_6215);
and U6493 (N_6493,N_6207,N_6057);
or U6494 (N_6494,N_6038,N_6054);
nor U6495 (N_6495,N_6160,N_6178);
nand U6496 (N_6496,N_6028,N_6222);
nand U6497 (N_6497,N_6205,N_6212);
nor U6498 (N_6498,N_6246,N_6087);
nand U6499 (N_6499,N_6041,N_6026);
nand U6500 (N_6500,N_6350,N_6348);
nand U6501 (N_6501,N_6368,N_6283);
nor U6502 (N_6502,N_6498,N_6468);
and U6503 (N_6503,N_6440,N_6407);
nor U6504 (N_6504,N_6391,N_6353);
nand U6505 (N_6505,N_6397,N_6262);
or U6506 (N_6506,N_6413,N_6433);
nand U6507 (N_6507,N_6434,N_6321);
nor U6508 (N_6508,N_6362,N_6320);
nor U6509 (N_6509,N_6340,N_6437);
or U6510 (N_6510,N_6270,N_6250);
nor U6511 (N_6511,N_6357,N_6483);
nor U6512 (N_6512,N_6431,N_6343);
and U6513 (N_6513,N_6354,N_6490);
nand U6514 (N_6514,N_6332,N_6421);
nand U6515 (N_6515,N_6331,N_6478);
and U6516 (N_6516,N_6319,N_6288);
nand U6517 (N_6517,N_6312,N_6449);
or U6518 (N_6518,N_6374,N_6306);
or U6519 (N_6519,N_6417,N_6268);
nor U6520 (N_6520,N_6394,N_6361);
nand U6521 (N_6521,N_6435,N_6359);
nand U6522 (N_6522,N_6488,N_6410);
nand U6523 (N_6523,N_6495,N_6304);
and U6524 (N_6524,N_6323,N_6390);
and U6525 (N_6525,N_6257,N_6396);
nor U6526 (N_6526,N_6302,N_6479);
nand U6527 (N_6527,N_6461,N_6252);
or U6528 (N_6528,N_6423,N_6327);
or U6529 (N_6529,N_6475,N_6356);
nand U6530 (N_6530,N_6378,N_6265);
nand U6531 (N_6531,N_6403,N_6412);
nand U6532 (N_6532,N_6287,N_6363);
xnor U6533 (N_6533,N_6339,N_6454);
nand U6534 (N_6534,N_6254,N_6464);
and U6535 (N_6535,N_6281,N_6429);
nor U6536 (N_6536,N_6329,N_6261);
or U6537 (N_6537,N_6451,N_6467);
nor U6538 (N_6538,N_6263,N_6290);
nand U6539 (N_6539,N_6486,N_6352);
and U6540 (N_6540,N_6401,N_6355);
nand U6541 (N_6541,N_6484,N_6346);
nand U6542 (N_6542,N_6317,N_6489);
and U6543 (N_6543,N_6476,N_6322);
and U6544 (N_6544,N_6389,N_6453);
nand U6545 (N_6545,N_6497,N_6289);
nand U6546 (N_6546,N_6485,N_6274);
nand U6547 (N_6547,N_6406,N_6324);
nand U6548 (N_6548,N_6336,N_6446);
or U6549 (N_6549,N_6482,N_6430);
and U6550 (N_6550,N_6445,N_6441);
nor U6551 (N_6551,N_6291,N_6309);
nand U6552 (N_6552,N_6258,N_6259);
nor U6553 (N_6553,N_6272,N_6305);
nor U6554 (N_6554,N_6293,N_6427);
nand U6555 (N_6555,N_6408,N_6360);
nand U6556 (N_6556,N_6448,N_6299);
nor U6557 (N_6557,N_6379,N_6260);
or U6558 (N_6558,N_6428,N_6269);
nor U6559 (N_6559,N_6499,N_6480);
and U6560 (N_6560,N_6273,N_6481);
nor U6561 (N_6561,N_6436,N_6316);
nand U6562 (N_6562,N_6298,N_6381);
nor U6563 (N_6563,N_6347,N_6251);
nand U6564 (N_6564,N_6366,N_6314);
and U6565 (N_6565,N_6395,N_6307);
nand U6566 (N_6566,N_6494,N_6473);
nand U6567 (N_6567,N_6458,N_6383);
nand U6568 (N_6568,N_6400,N_6333);
nor U6569 (N_6569,N_6328,N_6364);
nor U6570 (N_6570,N_6295,N_6308);
nand U6571 (N_6571,N_6402,N_6267);
nor U6572 (N_6572,N_6369,N_6470);
and U6573 (N_6573,N_6438,N_6424);
nor U6574 (N_6574,N_6469,N_6326);
nand U6575 (N_6575,N_6371,N_6447);
nor U6576 (N_6576,N_6455,N_6393);
nor U6577 (N_6577,N_6315,N_6418);
or U6578 (N_6578,N_6341,N_6384);
nand U6579 (N_6579,N_6313,N_6330);
or U6580 (N_6580,N_6422,N_6286);
nor U6581 (N_6581,N_6386,N_6474);
nor U6582 (N_6582,N_6277,N_6432);
nand U6583 (N_6583,N_6452,N_6491);
and U6584 (N_6584,N_6414,N_6275);
or U6585 (N_6585,N_6310,N_6311);
nand U6586 (N_6586,N_6344,N_6318);
nand U6587 (N_6587,N_6292,N_6325);
nand U6588 (N_6588,N_6377,N_6460);
nor U6589 (N_6589,N_6493,N_6337);
nor U6590 (N_6590,N_6496,N_6405);
or U6591 (N_6591,N_6375,N_6399);
nand U6592 (N_6592,N_6465,N_6284);
and U6593 (N_6593,N_6297,N_6444);
or U6594 (N_6594,N_6450,N_6463);
and U6595 (N_6595,N_6338,N_6459);
or U6596 (N_6596,N_6279,N_6342);
nor U6597 (N_6597,N_6349,N_6278);
and U6598 (N_6598,N_6276,N_6285);
nor U6599 (N_6599,N_6255,N_6398);
and U6600 (N_6600,N_6466,N_6351);
and U6601 (N_6601,N_6425,N_6380);
nand U6602 (N_6602,N_6388,N_6471);
nand U6603 (N_6603,N_6370,N_6294);
or U6604 (N_6604,N_6457,N_6385);
nand U6605 (N_6605,N_6303,N_6426);
or U6606 (N_6606,N_6492,N_6300);
or U6607 (N_6607,N_6472,N_6365);
nand U6608 (N_6608,N_6253,N_6266);
xor U6609 (N_6609,N_6392,N_6264);
nor U6610 (N_6610,N_6456,N_6409);
or U6611 (N_6611,N_6335,N_6271);
nand U6612 (N_6612,N_6372,N_6439);
or U6613 (N_6613,N_6256,N_6404);
nor U6614 (N_6614,N_6420,N_6415);
and U6615 (N_6615,N_6296,N_6442);
nand U6616 (N_6616,N_6416,N_6334);
and U6617 (N_6617,N_6387,N_6443);
nand U6618 (N_6618,N_6367,N_6358);
or U6619 (N_6619,N_6373,N_6376);
or U6620 (N_6620,N_6282,N_6487);
nor U6621 (N_6621,N_6462,N_6382);
nor U6622 (N_6622,N_6345,N_6411);
nand U6623 (N_6623,N_6301,N_6477);
and U6624 (N_6624,N_6419,N_6280);
xor U6625 (N_6625,N_6495,N_6488);
or U6626 (N_6626,N_6439,N_6450);
nor U6627 (N_6627,N_6388,N_6321);
or U6628 (N_6628,N_6425,N_6315);
nand U6629 (N_6629,N_6384,N_6332);
or U6630 (N_6630,N_6352,N_6359);
or U6631 (N_6631,N_6449,N_6472);
nand U6632 (N_6632,N_6430,N_6300);
and U6633 (N_6633,N_6297,N_6320);
and U6634 (N_6634,N_6327,N_6273);
nand U6635 (N_6635,N_6310,N_6329);
nand U6636 (N_6636,N_6283,N_6254);
or U6637 (N_6637,N_6410,N_6306);
or U6638 (N_6638,N_6473,N_6474);
and U6639 (N_6639,N_6470,N_6289);
or U6640 (N_6640,N_6295,N_6348);
or U6641 (N_6641,N_6323,N_6374);
or U6642 (N_6642,N_6368,N_6470);
and U6643 (N_6643,N_6481,N_6493);
or U6644 (N_6644,N_6350,N_6412);
nor U6645 (N_6645,N_6480,N_6421);
nor U6646 (N_6646,N_6438,N_6365);
nand U6647 (N_6647,N_6456,N_6253);
nand U6648 (N_6648,N_6481,N_6431);
and U6649 (N_6649,N_6397,N_6403);
nor U6650 (N_6650,N_6424,N_6472);
nor U6651 (N_6651,N_6418,N_6401);
nor U6652 (N_6652,N_6421,N_6424);
or U6653 (N_6653,N_6257,N_6377);
nand U6654 (N_6654,N_6256,N_6293);
nand U6655 (N_6655,N_6472,N_6490);
nor U6656 (N_6656,N_6330,N_6472);
nor U6657 (N_6657,N_6411,N_6253);
or U6658 (N_6658,N_6470,N_6294);
or U6659 (N_6659,N_6306,N_6477);
or U6660 (N_6660,N_6462,N_6378);
and U6661 (N_6661,N_6421,N_6428);
nor U6662 (N_6662,N_6451,N_6338);
or U6663 (N_6663,N_6440,N_6465);
nand U6664 (N_6664,N_6321,N_6443);
or U6665 (N_6665,N_6344,N_6435);
nor U6666 (N_6666,N_6495,N_6279);
and U6667 (N_6667,N_6445,N_6425);
nor U6668 (N_6668,N_6493,N_6385);
nor U6669 (N_6669,N_6285,N_6308);
nand U6670 (N_6670,N_6294,N_6324);
or U6671 (N_6671,N_6309,N_6321);
or U6672 (N_6672,N_6299,N_6453);
or U6673 (N_6673,N_6440,N_6307);
nor U6674 (N_6674,N_6345,N_6361);
or U6675 (N_6675,N_6381,N_6400);
or U6676 (N_6676,N_6319,N_6447);
nand U6677 (N_6677,N_6328,N_6472);
or U6678 (N_6678,N_6347,N_6385);
nor U6679 (N_6679,N_6386,N_6365);
nand U6680 (N_6680,N_6375,N_6313);
and U6681 (N_6681,N_6340,N_6355);
nor U6682 (N_6682,N_6481,N_6393);
and U6683 (N_6683,N_6321,N_6442);
nand U6684 (N_6684,N_6469,N_6307);
nand U6685 (N_6685,N_6446,N_6361);
and U6686 (N_6686,N_6293,N_6466);
or U6687 (N_6687,N_6376,N_6267);
nand U6688 (N_6688,N_6301,N_6455);
nor U6689 (N_6689,N_6492,N_6372);
nand U6690 (N_6690,N_6256,N_6357);
or U6691 (N_6691,N_6493,N_6387);
nor U6692 (N_6692,N_6352,N_6399);
and U6693 (N_6693,N_6341,N_6487);
or U6694 (N_6694,N_6493,N_6362);
nand U6695 (N_6695,N_6262,N_6377);
nand U6696 (N_6696,N_6404,N_6494);
nor U6697 (N_6697,N_6435,N_6450);
or U6698 (N_6698,N_6432,N_6288);
nor U6699 (N_6699,N_6266,N_6444);
and U6700 (N_6700,N_6376,N_6344);
nor U6701 (N_6701,N_6285,N_6419);
nand U6702 (N_6702,N_6304,N_6441);
nand U6703 (N_6703,N_6409,N_6437);
or U6704 (N_6704,N_6383,N_6382);
and U6705 (N_6705,N_6486,N_6350);
nor U6706 (N_6706,N_6458,N_6448);
or U6707 (N_6707,N_6385,N_6299);
and U6708 (N_6708,N_6363,N_6468);
and U6709 (N_6709,N_6439,N_6484);
or U6710 (N_6710,N_6424,N_6401);
nand U6711 (N_6711,N_6383,N_6401);
and U6712 (N_6712,N_6356,N_6295);
and U6713 (N_6713,N_6342,N_6404);
and U6714 (N_6714,N_6299,N_6482);
or U6715 (N_6715,N_6330,N_6357);
nand U6716 (N_6716,N_6465,N_6300);
and U6717 (N_6717,N_6268,N_6332);
nand U6718 (N_6718,N_6384,N_6263);
nor U6719 (N_6719,N_6319,N_6279);
nor U6720 (N_6720,N_6476,N_6343);
and U6721 (N_6721,N_6303,N_6382);
and U6722 (N_6722,N_6438,N_6272);
or U6723 (N_6723,N_6309,N_6417);
nor U6724 (N_6724,N_6427,N_6266);
or U6725 (N_6725,N_6404,N_6487);
and U6726 (N_6726,N_6398,N_6430);
nor U6727 (N_6727,N_6357,N_6393);
or U6728 (N_6728,N_6367,N_6331);
or U6729 (N_6729,N_6319,N_6326);
and U6730 (N_6730,N_6356,N_6464);
or U6731 (N_6731,N_6383,N_6334);
and U6732 (N_6732,N_6431,N_6319);
nand U6733 (N_6733,N_6358,N_6331);
nand U6734 (N_6734,N_6383,N_6317);
and U6735 (N_6735,N_6286,N_6291);
nand U6736 (N_6736,N_6421,N_6306);
nand U6737 (N_6737,N_6416,N_6384);
nor U6738 (N_6738,N_6349,N_6375);
nor U6739 (N_6739,N_6343,N_6366);
and U6740 (N_6740,N_6392,N_6365);
nor U6741 (N_6741,N_6344,N_6434);
nor U6742 (N_6742,N_6475,N_6260);
nand U6743 (N_6743,N_6418,N_6286);
nand U6744 (N_6744,N_6428,N_6444);
nand U6745 (N_6745,N_6447,N_6379);
and U6746 (N_6746,N_6308,N_6264);
xor U6747 (N_6747,N_6355,N_6351);
or U6748 (N_6748,N_6299,N_6356);
or U6749 (N_6749,N_6436,N_6305);
or U6750 (N_6750,N_6631,N_6572);
nor U6751 (N_6751,N_6629,N_6677);
and U6752 (N_6752,N_6684,N_6526);
nand U6753 (N_6753,N_6720,N_6636);
or U6754 (N_6754,N_6537,N_6669);
or U6755 (N_6755,N_6657,N_6639);
nor U6756 (N_6756,N_6571,N_6606);
nor U6757 (N_6757,N_6617,N_6730);
xor U6758 (N_6758,N_6687,N_6627);
nor U6759 (N_6759,N_6524,N_6634);
or U6760 (N_6760,N_6717,N_6530);
or U6761 (N_6761,N_6541,N_6696);
or U6762 (N_6762,N_6690,N_6500);
and U6763 (N_6763,N_6678,N_6722);
nand U6764 (N_6764,N_6507,N_6664);
xnor U6765 (N_6765,N_6551,N_6651);
nor U6766 (N_6766,N_6719,N_6726);
and U6767 (N_6767,N_6591,N_6703);
and U6768 (N_6768,N_6540,N_6577);
nor U6769 (N_6769,N_6580,N_6748);
or U6770 (N_6770,N_6701,N_6638);
nor U6771 (N_6771,N_6565,N_6501);
nand U6772 (N_6772,N_6645,N_6536);
nand U6773 (N_6773,N_6525,N_6532);
nor U6774 (N_6774,N_6714,N_6584);
or U6775 (N_6775,N_6670,N_6588);
or U6776 (N_6776,N_6517,N_6610);
nand U6777 (N_6777,N_6665,N_6566);
nor U6778 (N_6778,N_6693,N_6502);
nor U6779 (N_6779,N_6550,N_6522);
nor U6780 (N_6780,N_6582,N_6555);
or U6781 (N_6781,N_6688,N_6643);
nand U6782 (N_6782,N_6534,N_6734);
or U6783 (N_6783,N_6652,N_6671);
and U6784 (N_6784,N_6718,N_6654);
and U6785 (N_6785,N_6563,N_6663);
or U6786 (N_6786,N_6589,N_6595);
and U6787 (N_6787,N_6535,N_6647);
nor U6788 (N_6788,N_6587,N_6689);
nand U6789 (N_6789,N_6613,N_6641);
or U6790 (N_6790,N_6543,N_6523);
nand U6791 (N_6791,N_6650,N_6609);
nand U6792 (N_6792,N_6552,N_6620);
and U6793 (N_6793,N_6586,N_6702);
and U6794 (N_6794,N_6600,N_6708);
nand U6795 (N_6795,N_6527,N_6683);
nor U6796 (N_6796,N_6637,N_6542);
and U6797 (N_6797,N_6656,N_6642);
or U6798 (N_6798,N_6605,N_6632);
or U6799 (N_6799,N_6608,N_6731);
and U6800 (N_6800,N_6510,N_6514);
nor U6801 (N_6801,N_6668,N_6557);
or U6802 (N_6802,N_6594,N_6529);
nand U6803 (N_6803,N_6559,N_6513);
or U6804 (N_6804,N_6581,N_6685);
or U6805 (N_6805,N_6700,N_6698);
or U6806 (N_6806,N_6674,N_6503);
or U6807 (N_6807,N_6575,N_6635);
or U6808 (N_6808,N_6672,N_6622);
nor U6809 (N_6809,N_6679,N_6640);
or U6810 (N_6810,N_6740,N_6599);
nand U6811 (N_6811,N_6564,N_6604);
or U6812 (N_6812,N_6707,N_6603);
nor U6813 (N_6813,N_6616,N_6597);
and U6814 (N_6814,N_6583,N_6704);
and U6815 (N_6815,N_6625,N_6713);
nor U6816 (N_6816,N_6744,N_6621);
and U6817 (N_6817,N_6735,N_6697);
and U6818 (N_6818,N_6709,N_6662);
and U6819 (N_6819,N_6749,N_6691);
nor U6820 (N_6820,N_6607,N_6560);
or U6821 (N_6821,N_6729,N_6723);
nor U6822 (N_6822,N_6538,N_6711);
and U6823 (N_6823,N_6653,N_6661);
nor U6824 (N_6824,N_6633,N_6743);
and U6825 (N_6825,N_6533,N_6699);
nor U6826 (N_6826,N_6660,N_6673);
and U6827 (N_6827,N_6554,N_6547);
nor U6828 (N_6828,N_6515,N_6576);
and U6829 (N_6829,N_6738,N_6568);
nand U6830 (N_6830,N_6676,N_6614);
and U6831 (N_6831,N_6516,N_6659);
nor U6832 (N_6832,N_6686,N_6590);
or U6833 (N_6833,N_6544,N_6724);
nand U6834 (N_6834,N_6710,N_6742);
or U6835 (N_6835,N_6546,N_6624);
or U6836 (N_6836,N_6648,N_6585);
nand U6837 (N_6837,N_6509,N_6570);
nand U6838 (N_6838,N_6562,N_6666);
or U6839 (N_6839,N_6611,N_6528);
nand U6840 (N_6840,N_6721,N_6539);
or U6841 (N_6841,N_6618,N_6505);
nand U6842 (N_6842,N_6630,N_6695);
or U6843 (N_6843,N_6574,N_6593);
or U6844 (N_6844,N_6519,N_6692);
nand U6845 (N_6845,N_6553,N_6601);
or U6846 (N_6846,N_6705,N_6715);
or U6847 (N_6847,N_6682,N_6520);
nand U6848 (N_6848,N_6733,N_6619);
nand U6849 (N_6849,N_6579,N_6556);
or U6850 (N_6850,N_6626,N_6549);
nor U6851 (N_6851,N_6598,N_6747);
nand U6852 (N_6852,N_6578,N_6521);
nor U6853 (N_6853,N_6596,N_6667);
nor U6854 (N_6854,N_6739,N_6545);
nor U6855 (N_6855,N_6725,N_6658);
nand U6856 (N_6856,N_6741,N_6518);
nand U6857 (N_6857,N_6706,N_6716);
nor U6858 (N_6858,N_6649,N_6737);
or U6859 (N_6859,N_6628,N_6569);
or U6860 (N_6860,N_6592,N_6644);
nand U6861 (N_6861,N_6508,N_6615);
and U6862 (N_6862,N_6612,N_6623);
and U6863 (N_6863,N_6602,N_6506);
nor U6864 (N_6864,N_6531,N_6558);
nor U6865 (N_6865,N_6655,N_6745);
nor U6866 (N_6866,N_6680,N_6675);
nor U6867 (N_6867,N_6567,N_6728);
or U6868 (N_6868,N_6548,N_6504);
or U6869 (N_6869,N_6646,N_6512);
nand U6870 (N_6870,N_6746,N_6681);
nand U6871 (N_6871,N_6694,N_6573);
nor U6872 (N_6872,N_6561,N_6511);
and U6873 (N_6873,N_6727,N_6736);
nor U6874 (N_6874,N_6732,N_6712);
nand U6875 (N_6875,N_6551,N_6541);
and U6876 (N_6876,N_6575,N_6724);
nand U6877 (N_6877,N_6577,N_6710);
or U6878 (N_6878,N_6639,N_6744);
or U6879 (N_6879,N_6668,N_6542);
or U6880 (N_6880,N_6661,N_6654);
or U6881 (N_6881,N_6633,N_6582);
nand U6882 (N_6882,N_6555,N_6636);
and U6883 (N_6883,N_6609,N_6671);
and U6884 (N_6884,N_6710,N_6606);
nand U6885 (N_6885,N_6607,N_6635);
nand U6886 (N_6886,N_6623,N_6504);
and U6887 (N_6887,N_6658,N_6728);
and U6888 (N_6888,N_6660,N_6603);
or U6889 (N_6889,N_6549,N_6545);
nor U6890 (N_6890,N_6747,N_6501);
or U6891 (N_6891,N_6505,N_6549);
or U6892 (N_6892,N_6553,N_6580);
or U6893 (N_6893,N_6662,N_6552);
and U6894 (N_6894,N_6610,N_6529);
or U6895 (N_6895,N_6528,N_6602);
and U6896 (N_6896,N_6645,N_6610);
nor U6897 (N_6897,N_6738,N_6729);
nor U6898 (N_6898,N_6620,N_6643);
and U6899 (N_6899,N_6728,N_6632);
or U6900 (N_6900,N_6561,N_6582);
nor U6901 (N_6901,N_6689,N_6584);
nand U6902 (N_6902,N_6507,N_6569);
nor U6903 (N_6903,N_6517,N_6749);
nor U6904 (N_6904,N_6561,N_6595);
or U6905 (N_6905,N_6553,N_6747);
nand U6906 (N_6906,N_6597,N_6595);
or U6907 (N_6907,N_6655,N_6623);
or U6908 (N_6908,N_6518,N_6576);
nor U6909 (N_6909,N_6589,N_6564);
and U6910 (N_6910,N_6618,N_6515);
or U6911 (N_6911,N_6525,N_6714);
or U6912 (N_6912,N_6587,N_6743);
or U6913 (N_6913,N_6735,N_6541);
or U6914 (N_6914,N_6588,N_6625);
or U6915 (N_6915,N_6517,N_6633);
or U6916 (N_6916,N_6549,N_6667);
nor U6917 (N_6917,N_6630,N_6648);
nand U6918 (N_6918,N_6655,N_6538);
nand U6919 (N_6919,N_6647,N_6656);
nand U6920 (N_6920,N_6728,N_6637);
or U6921 (N_6921,N_6740,N_6687);
nand U6922 (N_6922,N_6612,N_6582);
and U6923 (N_6923,N_6585,N_6531);
or U6924 (N_6924,N_6630,N_6680);
nand U6925 (N_6925,N_6690,N_6645);
nor U6926 (N_6926,N_6651,N_6609);
or U6927 (N_6927,N_6627,N_6532);
nand U6928 (N_6928,N_6533,N_6559);
nor U6929 (N_6929,N_6740,N_6558);
nor U6930 (N_6930,N_6524,N_6607);
and U6931 (N_6931,N_6554,N_6571);
and U6932 (N_6932,N_6656,N_6578);
nand U6933 (N_6933,N_6674,N_6628);
and U6934 (N_6934,N_6619,N_6584);
xnor U6935 (N_6935,N_6533,N_6679);
and U6936 (N_6936,N_6675,N_6676);
nand U6937 (N_6937,N_6727,N_6733);
or U6938 (N_6938,N_6533,N_6627);
or U6939 (N_6939,N_6662,N_6633);
nor U6940 (N_6940,N_6698,N_6735);
or U6941 (N_6941,N_6511,N_6548);
and U6942 (N_6942,N_6516,N_6685);
and U6943 (N_6943,N_6679,N_6665);
nand U6944 (N_6944,N_6716,N_6721);
or U6945 (N_6945,N_6594,N_6735);
or U6946 (N_6946,N_6591,N_6520);
or U6947 (N_6947,N_6634,N_6654);
or U6948 (N_6948,N_6617,N_6568);
nor U6949 (N_6949,N_6695,N_6718);
nand U6950 (N_6950,N_6728,N_6696);
or U6951 (N_6951,N_6670,N_6663);
and U6952 (N_6952,N_6716,N_6665);
and U6953 (N_6953,N_6517,N_6564);
nand U6954 (N_6954,N_6561,N_6725);
nor U6955 (N_6955,N_6692,N_6593);
nand U6956 (N_6956,N_6704,N_6598);
or U6957 (N_6957,N_6510,N_6615);
nor U6958 (N_6958,N_6600,N_6520);
or U6959 (N_6959,N_6532,N_6531);
nand U6960 (N_6960,N_6712,N_6592);
nand U6961 (N_6961,N_6674,N_6720);
and U6962 (N_6962,N_6512,N_6589);
and U6963 (N_6963,N_6579,N_6599);
nor U6964 (N_6964,N_6723,N_6618);
and U6965 (N_6965,N_6674,N_6526);
and U6966 (N_6966,N_6716,N_6705);
nand U6967 (N_6967,N_6742,N_6535);
nand U6968 (N_6968,N_6711,N_6626);
nor U6969 (N_6969,N_6741,N_6635);
or U6970 (N_6970,N_6575,N_6596);
nor U6971 (N_6971,N_6662,N_6539);
nor U6972 (N_6972,N_6625,N_6548);
and U6973 (N_6973,N_6643,N_6590);
or U6974 (N_6974,N_6688,N_6526);
and U6975 (N_6975,N_6735,N_6642);
nand U6976 (N_6976,N_6569,N_6687);
nor U6977 (N_6977,N_6522,N_6732);
or U6978 (N_6978,N_6572,N_6603);
nand U6979 (N_6979,N_6635,N_6639);
and U6980 (N_6980,N_6520,N_6683);
and U6981 (N_6981,N_6583,N_6738);
nor U6982 (N_6982,N_6727,N_6587);
nand U6983 (N_6983,N_6525,N_6597);
nand U6984 (N_6984,N_6507,N_6554);
and U6985 (N_6985,N_6642,N_6514);
nand U6986 (N_6986,N_6658,N_6748);
nand U6987 (N_6987,N_6723,N_6731);
nand U6988 (N_6988,N_6584,N_6558);
or U6989 (N_6989,N_6627,N_6510);
nand U6990 (N_6990,N_6660,N_6690);
or U6991 (N_6991,N_6595,N_6549);
nand U6992 (N_6992,N_6539,N_6592);
or U6993 (N_6993,N_6597,N_6564);
nand U6994 (N_6994,N_6644,N_6667);
nand U6995 (N_6995,N_6613,N_6700);
nor U6996 (N_6996,N_6716,N_6587);
nand U6997 (N_6997,N_6659,N_6554);
nand U6998 (N_6998,N_6646,N_6525);
or U6999 (N_6999,N_6670,N_6692);
and U7000 (N_7000,N_6950,N_6750);
and U7001 (N_7001,N_6899,N_6829);
and U7002 (N_7002,N_6849,N_6973);
or U7003 (N_7003,N_6777,N_6954);
nand U7004 (N_7004,N_6904,N_6959);
and U7005 (N_7005,N_6864,N_6772);
and U7006 (N_7006,N_6969,N_6768);
nor U7007 (N_7007,N_6886,N_6916);
nand U7008 (N_7008,N_6977,N_6798);
and U7009 (N_7009,N_6919,N_6868);
nand U7010 (N_7010,N_6958,N_6957);
nor U7011 (N_7011,N_6811,N_6927);
nor U7012 (N_7012,N_6804,N_6932);
or U7013 (N_7013,N_6752,N_6862);
nor U7014 (N_7014,N_6838,N_6913);
or U7015 (N_7015,N_6826,N_6908);
nor U7016 (N_7016,N_6970,N_6762);
and U7017 (N_7017,N_6808,N_6814);
or U7018 (N_7018,N_6955,N_6924);
or U7019 (N_7019,N_6876,N_6931);
nor U7020 (N_7020,N_6995,N_6930);
or U7021 (N_7021,N_6994,N_6833);
and U7022 (N_7022,N_6902,N_6940);
nand U7023 (N_7023,N_6906,N_6914);
or U7024 (N_7024,N_6816,N_6929);
and U7025 (N_7025,N_6870,N_6837);
or U7026 (N_7026,N_6776,N_6810);
nor U7027 (N_7027,N_6791,N_6907);
nand U7028 (N_7028,N_6836,N_6821);
nand U7029 (N_7029,N_6892,N_6786);
and U7030 (N_7030,N_6858,N_6866);
nand U7031 (N_7031,N_6967,N_6872);
and U7032 (N_7032,N_6962,N_6869);
xnor U7033 (N_7033,N_6935,N_6765);
or U7034 (N_7034,N_6852,N_6889);
or U7035 (N_7035,N_6880,N_6802);
and U7036 (N_7036,N_6900,N_6767);
or U7037 (N_7037,N_6921,N_6897);
nand U7038 (N_7038,N_6839,N_6757);
and U7039 (N_7039,N_6953,N_6946);
or U7040 (N_7040,N_6778,N_6912);
and U7041 (N_7041,N_6817,N_6830);
or U7042 (N_7042,N_6846,N_6915);
nor U7043 (N_7043,N_6783,N_6766);
or U7044 (N_7044,N_6827,N_6898);
nor U7045 (N_7045,N_6853,N_6854);
or U7046 (N_7046,N_6999,N_6961);
nand U7047 (N_7047,N_6980,N_6834);
nor U7048 (N_7048,N_6806,N_6865);
nor U7049 (N_7049,N_6781,N_6945);
nand U7050 (N_7050,N_6888,N_6799);
and U7051 (N_7051,N_6943,N_6877);
or U7052 (N_7052,N_6797,N_6843);
nand U7053 (N_7053,N_6928,N_6990);
and U7054 (N_7054,N_6785,N_6784);
nor U7055 (N_7055,N_6754,N_6891);
or U7056 (N_7056,N_6769,N_6763);
or U7057 (N_7057,N_6947,N_6989);
or U7058 (N_7058,N_6795,N_6918);
and U7059 (N_7059,N_6993,N_6847);
nand U7060 (N_7060,N_6890,N_6857);
nand U7061 (N_7061,N_6801,N_6984);
nand U7062 (N_7062,N_6760,N_6911);
or U7063 (N_7063,N_6761,N_6972);
or U7064 (N_7064,N_6774,N_6780);
nand U7065 (N_7065,N_6922,N_6822);
or U7066 (N_7066,N_6820,N_6788);
nor U7067 (N_7067,N_6831,N_6963);
or U7068 (N_7068,N_6964,N_6985);
nand U7069 (N_7069,N_6818,N_6775);
nand U7070 (N_7070,N_6859,N_6867);
nand U7071 (N_7071,N_6812,N_6782);
nor U7072 (N_7072,N_6960,N_6895);
nand U7073 (N_7073,N_6986,N_6923);
or U7074 (N_7074,N_6988,N_6764);
nand U7075 (N_7075,N_6875,N_6840);
nor U7076 (N_7076,N_6809,N_6893);
and U7077 (N_7077,N_6910,N_6793);
nand U7078 (N_7078,N_6997,N_6887);
nand U7079 (N_7079,N_6753,N_6796);
or U7080 (N_7080,N_6894,N_6987);
nor U7081 (N_7081,N_6758,N_6825);
and U7082 (N_7082,N_6828,N_6979);
and U7083 (N_7083,N_6873,N_6934);
nand U7084 (N_7084,N_6882,N_6998);
or U7085 (N_7085,N_6982,N_6850);
nand U7086 (N_7086,N_6805,N_6884);
nand U7087 (N_7087,N_6878,N_6794);
and U7088 (N_7088,N_6759,N_6779);
or U7089 (N_7089,N_6917,N_6855);
nor U7090 (N_7090,N_6789,N_6991);
nand U7091 (N_7091,N_6815,N_6813);
or U7092 (N_7092,N_6936,N_6860);
and U7093 (N_7093,N_6926,N_6771);
nand U7094 (N_7094,N_6966,N_6863);
nor U7095 (N_7095,N_6905,N_6944);
or U7096 (N_7096,N_6787,N_6819);
or U7097 (N_7097,N_6832,N_6939);
and U7098 (N_7098,N_6976,N_6874);
nor U7099 (N_7099,N_6951,N_6844);
and U7100 (N_7100,N_6965,N_6755);
or U7101 (N_7101,N_6807,N_6903);
or U7102 (N_7102,N_6751,N_6835);
nor U7103 (N_7103,N_6861,N_6949);
or U7104 (N_7104,N_6823,N_6942);
nor U7105 (N_7105,N_6920,N_6845);
nor U7106 (N_7106,N_6790,N_6773);
or U7107 (N_7107,N_6971,N_6925);
nor U7108 (N_7108,N_6978,N_6933);
nor U7109 (N_7109,N_6848,N_6974);
or U7110 (N_7110,N_6871,N_6851);
nor U7111 (N_7111,N_6952,N_6879);
or U7112 (N_7112,N_6975,N_6981);
and U7113 (N_7113,N_6883,N_6770);
nor U7114 (N_7114,N_6938,N_6803);
and U7115 (N_7115,N_6996,N_6756);
or U7116 (N_7116,N_6992,N_6800);
nor U7117 (N_7117,N_6885,N_6881);
and U7118 (N_7118,N_6909,N_6841);
and U7119 (N_7119,N_6956,N_6937);
nor U7120 (N_7120,N_6968,N_6948);
nor U7121 (N_7121,N_6824,N_6842);
nand U7122 (N_7122,N_6941,N_6792);
and U7123 (N_7123,N_6983,N_6901);
or U7124 (N_7124,N_6896,N_6856);
nand U7125 (N_7125,N_6965,N_6948);
nor U7126 (N_7126,N_6834,N_6845);
and U7127 (N_7127,N_6775,N_6887);
nor U7128 (N_7128,N_6958,N_6826);
nor U7129 (N_7129,N_6995,N_6783);
or U7130 (N_7130,N_6990,N_6786);
nor U7131 (N_7131,N_6825,N_6904);
nand U7132 (N_7132,N_6765,N_6990);
nand U7133 (N_7133,N_6874,N_6997);
or U7134 (N_7134,N_6893,N_6916);
nor U7135 (N_7135,N_6854,N_6759);
nor U7136 (N_7136,N_6802,N_6966);
or U7137 (N_7137,N_6827,N_6952);
and U7138 (N_7138,N_6937,N_6907);
and U7139 (N_7139,N_6891,N_6752);
and U7140 (N_7140,N_6946,N_6870);
nor U7141 (N_7141,N_6898,N_6878);
and U7142 (N_7142,N_6925,N_6905);
nand U7143 (N_7143,N_6848,N_6895);
and U7144 (N_7144,N_6852,N_6878);
nand U7145 (N_7145,N_6957,N_6900);
nor U7146 (N_7146,N_6923,N_6783);
xnor U7147 (N_7147,N_6842,N_6928);
or U7148 (N_7148,N_6933,N_6783);
nand U7149 (N_7149,N_6946,N_6811);
nand U7150 (N_7150,N_6974,N_6840);
nand U7151 (N_7151,N_6990,N_6822);
and U7152 (N_7152,N_6985,N_6972);
nand U7153 (N_7153,N_6831,N_6882);
nor U7154 (N_7154,N_6813,N_6797);
nor U7155 (N_7155,N_6999,N_6811);
and U7156 (N_7156,N_6999,N_6998);
and U7157 (N_7157,N_6980,N_6967);
nand U7158 (N_7158,N_6792,N_6765);
nand U7159 (N_7159,N_6849,N_6980);
nand U7160 (N_7160,N_6889,N_6787);
or U7161 (N_7161,N_6902,N_6926);
and U7162 (N_7162,N_6957,N_6924);
or U7163 (N_7163,N_6965,N_6944);
and U7164 (N_7164,N_6901,N_6889);
nor U7165 (N_7165,N_6831,N_6909);
and U7166 (N_7166,N_6759,N_6910);
and U7167 (N_7167,N_6795,N_6762);
and U7168 (N_7168,N_6967,N_6838);
and U7169 (N_7169,N_6824,N_6884);
and U7170 (N_7170,N_6859,N_6761);
nand U7171 (N_7171,N_6909,N_6770);
nand U7172 (N_7172,N_6799,N_6932);
or U7173 (N_7173,N_6959,N_6950);
nand U7174 (N_7174,N_6833,N_6953);
nand U7175 (N_7175,N_6988,N_6807);
or U7176 (N_7176,N_6907,N_6780);
or U7177 (N_7177,N_6903,N_6806);
or U7178 (N_7178,N_6964,N_6814);
and U7179 (N_7179,N_6768,N_6811);
and U7180 (N_7180,N_6924,N_6862);
nand U7181 (N_7181,N_6936,N_6927);
and U7182 (N_7182,N_6979,N_6844);
or U7183 (N_7183,N_6924,N_6882);
nor U7184 (N_7184,N_6899,N_6865);
or U7185 (N_7185,N_6868,N_6821);
nand U7186 (N_7186,N_6812,N_6876);
nand U7187 (N_7187,N_6839,N_6834);
or U7188 (N_7188,N_6962,N_6955);
or U7189 (N_7189,N_6936,N_6757);
nand U7190 (N_7190,N_6841,N_6760);
nand U7191 (N_7191,N_6820,N_6758);
and U7192 (N_7192,N_6995,N_6934);
nor U7193 (N_7193,N_6860,N_6975);
and U7194 (N_7194,N_6763,N_6760);
nor U7195 (N_7195,N_6791,N_6879);
and U7196 (N_7196,N_6966,N_6906);
or U7197 (N_7197,N_6764,N_6934);
nor U7198 (N_7198,N_6926,N_6817);
nand U7199 (N_7199,N_6994,N_6956);
and U7200 (N_7200,N_6811,N_6952);
or U7201 (N_7201,N_6751,N_6928);
nor U7202 (N_7202,N_6983,N_6904);
or U7203 (N_7203,N_6827,N_6946);
or U7204 (N_7204,N_6944,N_6881);
nor U7205 (N_7205,N_6875,N_6878);
and U7206 (N_7206,N_6817,N_6984);
and U7207 (N_7207,N_6848,N_6752);
and U7208 (N_7208,N_6767,N_6793);
and U7209 (N_7209,N_6878,N_6808);
and U7210 (N_7210,N_6895,N_6797);
nor U7211 (N_7211,N_6770,N_6911);
nor U7212 (N_7212,N_6795,N_6988);
and U7213 (N_7213,N_6817,N_6815);
nor U7214 (N_7214,N_6922,N_6908);
and U7215 (N_7215,N_6870,N_6933);
nand U7216 (N_7216,N_6957,N_6940);
nor U7217 (N_7217,N_6865,N_6889);
or U7218 (N_7218,N_6800,N_6889);
or U7219 (N_7219,N_6982,N_6844);
nand U7220 (N_7220,N_6985,N_6850);
and U7221 (N_7221,N_6915,N_6918);
nand U7222 (N_7222,N_6999,N_6812);
nor U7223 (N_7223,N_6886,N_6803);
nand U7224 (N_7224,N_6891,N_6815);
and U7225 (N_7225,N_6786,N_6773);
nand U7226 (N_7226,N_6926,N_6892);
nand U7227 (N_7227,N_6942,N_6818);
and U7228 (N_7228,N_6944,N_6864);
or U7229 (N_7229,N_6830,N_6849);
or U7230 (N_7230,N_6894,N_6771);
nor U7231 (N_7231,N_6828,N_6925);
nand U7232 (N_7232,N_6811,N_6960);
nor U7233 (N_7233,N_6934,N_6761);
and U7234 (N_7234,N_6759,N_6911);
and U7235 (N_7235,N_6962,N_6902);
nand U7236 (N_7236,N_6984,N_6846);
nor U7237 (N_7237,N_6795,N_6946);
or U7238 (N_7238,N_6883,N_6974);
nand U7239 (N_7239,N_6858,N_6763);
nand U7240 (N_7240,N_6850,N_6793);
and U7241 (N_7241,N_6816,N_6906);
nand U7242 (N_7242,N_6882,N_6875);
or U7243 (N_7243,N_6853,N_6795);
nor U7244 (N_7244,N_6804,N_6955);
and U7245 (N_7245,N_6755,N_6938);
nand U7246 (N_7246,N_6816,N_6782);
or U7247 (N_7247,N_6823,N_6756);
nor U7248 (N_7248,N_6753,N_6829);
or U7249 (N_7249,N_6822,N_6940);
xor U7250 (N_7250,N_7066,N_7165);
and U7251 (N_7251,N_7164,N_7246);
and U7252 (N_7252,N_7052,N_7200);
or U7253 (N_7253,N_7069,N_7145);
and U7254 (N_7254,N_7082,N_7088);
nand U7255 (N_7255,N_7089,N_7056);
nand U7256 (N_7256,N_7199,N_7023);
or U7257 (N_7257,N_7085,N_7074);
or U7258 (N_7258,N_7133,N_7060);
or U7259 (N_7259,N_7059,N_7180);
nand U7260 (N_7260,N_7214,N_7243);
nor U7261 (N_7261,N_7135,N_7095);
nand U7262 (N_7262,N_7004,N_7010);
or U7263 (N_7263,N_7012,N_7048);
nor U7264 (N_7264,N_7031,N_7249);
or U7265 (N_7265,N_7072,N_7077);
and U7266 (N_7266,N_7049,N_7104);
or U7267 (N_7267,N_7197,N_7203);
nor U7268 (N_7268,N_7212,N_7114);
and U7269 (N_7269,N_7171,N_7054);
nor U7270 (N_7270,N_7020,N_7144);
nand U7271 (N_7271,N_7198,N_7110);
and U7272 (N_7272,N_7011,N_7018);
or U7273 (N_7273,N_7157,N_7235);
and U7274 (N_7274,N_7136,N_7134);
nand U7275 (N_7275,N_7227,N_7099);
nor U7276 (N_7276,N_7219,N_7042);
nand U7277 (N_7277,N_7016,N_7075);
or U7278 (N_7278,N_7087,N_7137);
nor U7279 (N_7279,N_7143,N_7106);
and U7280 (N_7280,N_7209,N_7167);
or U7281 (N_7281,N_7067,N_7131);
nand U7282 (N_7282,N_7022,N_7037);
nand U7283 (N_7283,N_7228,N_7027);
and U7284 (N_7284,N_7210,N_7116);
or U7285 (N_7285,N_7166,N_7148);
nor U7286 (N_7286,N_7040,N_7242);
or U7287 (N_7287,N_7097,N_7083);
and U7288 (N_7288,N_7140,N_7240);
nor U7289 (N_7289,N_7124,N_7035);
nor U7290 (N_7290,N_7008,N_7232);
nor U7291 (N_7291,N_7221,N_7001);
nand U7292 (N_7292,N_7032,N_7194);
nand U7293 (N_7293,N_7147,N_7019);
or U7294 (N_7294,N_7046,N_7247);
nor U7295 (N_7295,N_7244,N_7039);
nand U7296 (N_7296,N_7123,N_7142);
or U7297 (N_7297,N_7113,N_7132);
or U7298 (N_7298,N_7120,N_7204);
nand U7299 (N_7299,N_7026,N_7101);
nor U7300 (N_7300,N_7150,N_7160);
or U7301 (N_7301,N_7055,N_7118);
nand U7302 (N_7302,N_7217,N_7159);
and U7303 (N_7303,N_7156,N_7183);
nand U7304 (N_7304,N_7090,N_7080);
nand U7305 (N_7305,N_7182,N_7061);
or U7306 (N_7306,N_7102,N_7107);
nor U7307 (N_7307,N_7126,N_7108);
or U7308 (N_7308,N_7201,N_7216);
nand U7309 (N_7309,N_7234,N_7062);
nor U7310 (N_7310,N_7033,N_7236);
or U7311 (N_7311,N_7015,N_7245);
xnor U7312 (N_7312,N_7161,N_7051);
nand U7313 (N_7313,N_7076,N_7154);
or U7314 (N_7314,N_7112,N_7237);
or U7315 (N_7315,N_7231,N_7025);
nor U7316 (N_7316,N_7172,N_7014);
nand U7317 (N_7317,N_7065,N_7169);
xor U7318 (N_7318,N_7153,N_7206);
or U7319 (N_7319,N_7239,N_7207);
and U7320 (N_7320,N_7000,N_7128);
and U7321 (N_7321,N_7196,N_7050);
nor U7322 (N_7322,N_7189,N_7129);
nor U7323 (N_7323,N_7086,N_7092);
or U7324 (N_7324,N_7096,N_7175);
and U7325 (N_7325,N_7127,N_7007);
nor U7326 (N_7326,N_7173,N_7105);
and U7327 (N_7327,N_7111,N_7178);
nor U7328 (N_7328,N_7071,N_7091);
and U7329 (N_7329,N_7146,N_7229);
or U7330 (N_7330,N_7094,N_7079);
or U7331 (N_7331,N_7058,N_7177);
nand U7332 (N_7332,N_7130,N_7029);
or U7333 (N_7333,N_7036,N_7081);
nor U7334 (N_7334,N_7225,N_7176);
or U7335 (N_7335,N_7230,N_7045);
nor U7336 (N_7336,N_7041,N_7034);
or U7337 (N_7337,N_7070,N_7005);
nand U7338 (N_7338,N_7002,N_7179);
nand U7339 (N_7339,N_7125,N_7241);
nor U7340 (N_7340,N_7226,N_7195);
or U7341 (N_7341,N_7044,N_7047);
or U7342 (N_7342,N_7205,N_7248);
and U7343 (N_7343,N_7053,N_7238);
nand U7344 (N_7344,N_7155,N_7218);
or U7345 (N_7345,N_7163,N_7006);
or U7346 (N_7346,N_7003,N_7109);
or U7347 (N_7347,N_7030,N_7185);
and U7348 (N_7348,N_7220,N_7170);
or U7349 (N_7349,N_7028,N_7117);
nand U7350 (N_7350,N_7013,N_7038);
or U7351 (N_7351,N_7187,N_7119);
nand U7352 (N_7352,N_7139,N_7202);
and U7353 (N_7353,N_7138,N_7186);
nor U7354 (N_7354,N_7224,N_7098);
or U7355 (N_7355,N_7057,N_7115);
and U7356 (N_7356,N_7024,N_7215);
nor U7357 (N_7357,N_7168,N_7190);
nand U7358 (N_7358,N_7188,N_7093);
nor U7359 (N_7359,N_7223,N_7213);
nand U7360 (N_7360,N_7149,N_7084);
nor U7361 (N_7361,N_7151,N_7158);
or U7362 (N_7362,N_7233,N_7193);
or U7363 (N_7363,N_7141,N_7184);
nand U7364 (N_7364,N_7100,N_7017);
and U7365 (N_7365,N_7078,N_7211);
and U7366 (N_7366,N_7021,N_7121);
and U7367 (N_7367,N_7068,N_7181);
nor U7368 (N_7368,N_7162,N_7208);
nand U7369 (N_7369,N_7043,N_7122);
xnor U7370 (N_7370,N_7103,N_7192);
nand U7371 (N_7371,N_7073,N_7174);
nor U7372 (N_7372,N_7064,N_7009);
and U7373 (N_7373,N_7191,N_7063);
nor U7374 (N_7374,N_7152,N_7222);
and U7375 (N_7375,N_7093,N_7064);
nor U7376 (N_7376,N_7169,N_7141);
and U7377 (N_7377,N_7167,N_7085);
nor U7378 (N_7378,N_7212,N_7148);
nand U7379 (N_7379,N_7161,N_7038);
nor U7380 (N_7380,N_7200,N_7016);
and U7381 (N_7381,N_7007,N_7199);
and U7382 (N_7382,N_7136,N_7122);
or U7383 (N_7383,N_7161,N_7227);
and U7384 (N_7384,N_7083,N_7138);
and U7385 (N_7385,N_7138,N_7132);
nand U7386 (N_7386,N_7009,N_7033);
and U7387 (N_7387,N_7100,N_7153);
or U7388 (N_7388,N_7119,N_7148);
nand U7389 (N_7389,N_7196,N_7121);
nor U7390 (N_7390,N_7234,N_7070);
nor U7391 (N_7391,N_7022,N_7152);
nor U7392 (N_7392,N_7109,N_7002);
nor U7393 (N_7393,N_7144,N_7042);
and U7394 (N_7394,N_7237,N_7176);
or U7395 (N_7395,N_7022,N_7118);
nand U7396 (N_7396,N_7071,N_7185);
or U7397 (N_7397,N_7085,N_7131);
nand U7398 (N_7398,N_7017,N_7039);
nor U7399 (N_7399,N_7059,N_7137);
or U7400 (N_7400,N_7098,N_7088);
and U7401 (N_7401,N_7051,N_7088);
nor U7402 (N_7402,N_7001,N_7121);
nand U7403 (N_7403,N_7203,N_7086);
nor U7404 (N_7404,N_7087,N_7074);
or U7405 (N_7405,N_7204,N_7084);
nor U7406 (N_7406,N_7157,N_7184);
or U7407 (N_7407,N_7233,N_7060);
nor U7408 (N_7408,N_7211,N_7225);
nor U7409 (N_7409,N_7147,N_7068);
or U7410 (N_7410,N_7043,N_7218);
nand U7411 (N_7411,N_7086,N_7141);
nand U7412 (N_7412,N_7074,N_7145);
nand U7413 (N_7413,N_7052,N_7114);
nand U7414 (N_7414,N_7243,N_7235);
nand U7415 (N_7415,N_7029,N_7135);
nor U7416 (N_7416,N_7045,N_7130);
and U7417 (N_7417,N_7102,N_7097);
nor U7418 (N_7418,N_7222,N_7025);
nor U7419 (N_7419,N_7064,N_7181);
nor U7420 (N_7420,N_7032,N_7015);
nand U7421 (N_7421,N_7247,N_7148);
or U7422 (N_7422,N_7155,N_7010);
nand U7423 (N_7423,N_7171,N_7044);
nor U7424 (N_7424,N_7139,N_7095);
nand U7425 (N_7425,N_7144,N_7226);
nor U7426 (N_7426,N_7126,N_7023);
nor U7427 (N_7427,N_7042,N_7093);
or U7428 (N_7428,N_7145,N_7174);
or U7429 (N_7429,N_7086,N_7201);
nand U7430 (N_7430,N_7195,N_7160);
nand U7431 (N_7431,N_7051,N_7225);
or U7432 (N_7432,N_7017,N_7071);
or U7433 (N_7433,N_7198,N_7246);
and U7434 (N_7434,N_7095,N_7212);
nor U7435 (N_7435,N_7201,N_7126);
or U7436 (N_7436,N_7083,N_7062);
nor U7437 (N_7437,N_7080,N_7118);
and U7438 (N_7438,N_7011,N_7036);
or U7439 (N_7439,N_7061,N_7074);
and U7440 (N_7440,N_7123,N_7092);
nor U7441 (N_7441,N_7174,N_7229);
nand U7442 (N_7442,N_7081,N_7055);
or U7443 (N_7443,N_7034,N_7046);
or U7444 (N_7444,N_7150,N_7069);
nor U7445 (N_7445,N_7097,N_7121);
nor U7446 (N_7446,N_7221,N_7064);
or U7447 (N_7447,N_7105,N_7068);
nor U7448 (N_7448,N_7171,N_7236);
nand U7449 (N_7449,N_7158,N_7198);
or U7450 (N_7450,N_7092,N_7229);
or U7451 (N_7451,N_7078,N_7027);
and U7452 (N_7452,N_7108,N_7127);
nand U7453 (N_7453,N_7024,N_7225);
nand U7454 (N_7454,N_7011,N_7204);
and U7455 (N_7455,N_7213,N_7046);
nand U7456 (N_7456,N_7058,N_7089);
or U7457 (N_7457,N_7207,N_7119);
nand U7458 (N_7458,N_7097,N_7198);
or U7459 (N_7459,N_7135,N_7053);
nand U7460 (N_7460,N_7161,N_7131);
and U7461 (N_7461,N_7059,N_7139);
nand U7462 (N_7462,N_7094,N_7237);
or U7463 (N_7463,N_7248,N_7080);
nand U7464 (N_7464,N_7229,N_7134);
nand U7465 (N_7465,N_7036,N_7031);
nor U7466 (N_7466,N_7085,N_7222);
nor U7467 (N_7467,N_7183,N_7063);
nand U7468 (N_7468,N_7243,N_7147);
and U7469 (N_7469,N_7097,N_7148);
nor U7470 (N_7470,N_7028,N_7045);
or U7471 (N_7471,N_7106,N_7156);
nand U7472 (N_7472,N_7035,N_7141);
and U7473 (N_7473,N_7125,N_7075);
nor U7474 (N_7474,N_7132,N_7167);
nand U7475 (N_7475,N_7063,N_7156);
and U7476 (N_7476,N_7114,N_7099);
or U7477 (N_7477,N_7057,N_7111);
nor U7478 (N_7478,N_7236,N_7201);
or U7479 (N_7479,N_7122,N_7163);
nor U7480 (N_7480,N_7105,N_7046);
or U7481 (N_7481,N_7194,N_7184);
or U7482 (N_7482,N_7091,N_7155);
nor U7483 (N_7483,N_7024,N_7008);
or U7484 (N_7484,N_7081,N_7109);
or U7485 (N_7485,N_7245,N_7011);
or U7486 (N_7486,N_7162,N_7137);
nand U7487 (N_7487,N_7235,N_7002);
nor U7488 (N_7488,N_7203,N_7206);
and U7489 (N_7489,N_7166,N_7076);
and U7490 (N_7490,N_7238,N_7086);
nor U7491 (N_7491,N_7159,N_7197);
xor U7492 (N_7492,N_7248,N_7036);
nor U7493 (N_7493,N_7080,N_7096);
nor U7494 (N_7494,N_7052,N_7034);
nand U7495 (N_7495,N_7220,N_7066);
nor U7496 (N_7496,N_7032,N_7031);
nand U7497 (N_7497,N_7025,N_7216);
and U7498 (N_7498,N_7247,N_7042);
nor U7499 (N_7499,N_7014,N_7065);
and U7500 (N_7500,N_7370,N_7439);
nand U7501 (N_7501,N_7498,N_7483);
or U7502 (N_7502,N_7292,N_7276);
and U7503 (N_7503,N_7307,N_7329);
nand U7504 (N_7504,N_7466,N_7308);
nor U7505 (N_7505,N_7476,N_7350);
nand U7506 (N_7506,N_7458,N_7294);
and U7507 (N_7507,N_7260,N_7290);
and U7508 (N_7508,N_7358,N_7306);
or U7509 (N_7509,N_7264,N_7461);
nor U7510 (N_7510,N_7443,N_7356);
nand U7511 (N_7511,N_7398,N_7481);
nand U7512 (N_7512,N_7420,N_7313);
and U7513 (N_7513,N_7499,N_7257);
nand U7514 (N_7514,N_7451,N_7280);
and U7515 (N_7515,N_7359,N_7427);
or U7516 (N_7516,N_7312,N_7347);
and U7517 (N_7517,N_7365,N_7395);
and U7518 (N_7518,N_7304,N_7343);
and U7519 (N_7519,N_7409,N_7465);
nor U7520 (N_7520,N_7303,N_7385);
or U7521 (N_7521,N_7445,N_7273);
nand U7522 (N_7522,N_7418,N_7277);
nand U7523 (N_7523,N_7255,N_7386);
or U7524 (N_7524,N_7421,N_7298);
and U7525 (N_7525,N_7301,N_7355);
and U7526 (N_7526,N_7402,N_7423);
or U7527 (N_7527,N_7468,N_7340);
or U7528 (N_7528,N_7253,N_7442);
or U7529 (N_7529,N_7318,N_7413);
or U7530 (N_7530,N_7474,N_7464);
nand U7531 (N_7531,N_7414,N_7394);
nor U7532 (N_7532,N_7361,N_7428);
and U7533 (N_7533,N_7497,N_7388);
or U7534 (N_7534,N_7315,N_7486);
nand U7535 (N_7535,N_7422,N_7351);
and U7536 (N_7536,N_7339,N_7256);
nand U7537 (N_7537,N_7321,N_7327);
or U7538 (N_7538,N_7432,N_7455);
xnor U7539 (N_7539,N_7381,N_7462);
nor U7540 (N_7540,N_7281,N_7447);
nor U7541 (N_7541,N_7289,N_7478);
nor U7542 (N_7542,N_7396,N_7407);
and U7543 (N_7543,N_7285,N_7334);
and U7544 (N_7544,N_7267,N_7263);
and U7545 (N_7545,N_7283,N_7410);
nor U7546 (N_7546,N_7317,N_7484);
nor U7547 (N_7547,N_7332,N_7282);
nor U7548 (N_7548,N_7341,N_7374);
or U7549 (N_7549,N_7431,N_7363);
nand U7550 (N_7550,N_7411,N_7252);
and U7551 (N_7551,N_7324,N_7390);
or U7552 (N_7552,N_7380,N_7275);
or U7553 (N_7553,N_7446,N_7258);
nor U7554 (N_7554,N_7482,N_7412);
nor U7555 (N_7555,N_7354,N_7477);
nor U7556 (N_7556,N_7438,N_7251);
or U7557 (N_7557,N_7357,N_7314);
and U7558 (N_7558,N_7373,N_7371);
and U7559 (N_7559,N_7403,N_7353);
and U7560 (N_7560,N_7435,N_7364);
nand U7561 (N_7561,N_7459,N_7261);
and U7562 (N_7562,N_7299,N_7408);
and U7563 (N_7563,N_7378,N_7489);
or U7564 (N_7564,N_7453,N_7325);
or U7565 (N_7565,N_7291,N_7367);
or U7566 (N_7566,N_7425,N_7316);
nor U7567 (N_7567,N_7473,N_7470);
nor U7568 (N_7568,N_7479,N_7405);
or U7569 (N_7569,N_7360,N_7415);
or U7570 (N_7570,N_7288,N_7310);
or U7571 (N_7571,N_7436,N_7254);
or U7572 (N_7572,N_7467,N_7305);
or U7573 (N_7573,N_7495,N_7278);
nor U7574 (N_7574,N_7399,N_7469);
xnor U7575 (N_7575,N_7491,N_7487);
and U7576 (N_7576,N_7279,N_7384);
nand U7577 (N_7577,N_7377,N_7322);
nand U7578 (N_7578,N_7349,N_7492);
nand U7579 (N_7579,N_7393,N_7320);
nand U7580 (N_7580,N_7488,N_7426);
and U7581 (N_7581,N_7284,N_7366);
or U7582 (N_7582,N_7379,N_7406);
or U7583 (N_7583,N_7429,N_7480);
and U7584 (N_7584,N_7401,N_7452);
nor U7585 (N_7585,N_7392,N_7376);
nand U7586 (N_7586,N_7293,N_7419);
or U7587 (N_7587,N_7404,N_7433);
nor U7588 (N_7588,N_7493,N_7262);
or U7589 (N_7589,N_7272,N_7463);
nor U7590 (N_7590,N_7300,N_7485);
nand U7591 (N_7591,N_7330,N_7372);
and U7592 (N_7592,N_7297,N_7400);
nor U7593 (N_7593,N_7430,N_7424);
and U7594 (N_7594,N_7450,N_7259);
and U7595 (N_7595,N_7490,N_7335);
nand U7596 (N_7596,N_7397,N_7440);
nand U7597 (N_7597,N_7369,N_7302);
nand U7598 (N_7598,N_7270,N_7268);
nor U7599 (N_7599,N_7323,N_7391);
and U7600 (N_7600,N_7417,N_7348);
or U7601 (N_7601,N_7265,N_7271);
or U7602 (N_7602,N_7250,N_7326);
nand U7603 (N_7603,N_7416,N_7449);
nand U7604 (N_7604,N_7287,N_7383);
or U7605 (N_7605,N_7328,N_7266);
and U7606 (N_7606,N_7333,N_7382);
and U7607 (N_7607,N_7286,N_7496);
or U7608 (N_7608,N_7269,N_7274);
or U7609 (N_7609,N_7296,N_7441);
nor U7610 (N_7610,N_7342,N_7389);
and U7611 (N_7611,N_7494,N_7475);
or U7612 (N_7612,N_7346,N_7387);
nand U7613 (N_7613,N_7472,N_7344);
and U7614 (N_7614,N_7295,N_7460);
nor U7615 (N_7615,N_7471,N_7457);
nor U7616 (N_7616,N_7352,N_7434);
nand U7617 (N_7617,N_7345,N_7319);
and U7618 (N_7618,N_7437,N_7337);
nor U7619 (N_7619,N_7444,N_7309);
nand U7620 (N_7620,N_7362,N_7331);
and U7621 (N_7621,N_7368,N_7456);
nor U7622 (N_7622,N_7336,N_7375);
or U7623 (N_7623,N_7454,N_7311);
or U7624 (N_7624,N_7338,N_7448);
or U7625 (N_7625,N_7376,N_7486);
nand U7626 (N_7626,N_7278,N_7296);
xor U7627 (N_7627,N_7289,N_7459);
or U7628 (N_7628,N_7373,N_7447);
nand U7629 (N_7629,N_7256,N_7330);
nor U7630 (N_7630,N_7257,N_7350);
and U7631 (N_7631,N_7374,N_7475);
and U7632 (N_7632,N_7470,N_7353);
and U7633 (N_7633,N_7415,N_7268);
nand U7634 (N_7634,N_7488,N_7484);
nand U7635 (N_7635,N_7495,N_7498);
nor U7636 (N_7636,N_7314,N_7351);
nand U7637 (N_7637,N_7473,N_7351);
nand U7638 (N_7638,N_7315,N_7337);
and U7639 (N_7639,N_7333,N_7269);
nand U7640 (N_7640,N_7405,N_7442);
or U7641 (N_7641,N_7367,N_7458);
xnor U7642 (N_7642,N_7366,N_7270);
and U7643 (N_7643,N_7369,N_7379);
nor U7644 (N_7644,N_7386,N_7475);
xnor U7645 (N_7645,N_7352,N_7401);
nor U7646 (N_7646,N_7483,N_7468);
and U7647 (N_7647,N_7264,N_7403);
or U7648 (N_7648,N_7494,N_7258);
nand U7649 (N_7649,N_7347,N_7412);
or U7650 (N_7650,N_7364,N_7329);
and U7651 (N_7651,N_7266,N_7386);
nor U7652 (N_7652,N_7469,N_7296);
nor U7653 (N_7653,N_7285,N_7307);
nor U7654 (N_7654,N_7489,N_7490);
and U7655 (N_7655,N_7423,N_7290);
nor U7656 (N_7656,N_7494,N_7486);
and U7657 (N_7657,N_7312,N_7410);
or U7658 (N_7658,N_7426,N_7250);
nand U7659 (N_7659,N_7265,N_7423);
and U7660 (N_7660,N_7258,N_7487);
or U7661 (N_7661,N_7348,N_7457);
and U7662 (N_7662,N_7494,N_7328);
and U7663 (N_7663,N_7405,N_7424);
nor U7664 (N_7664,N_7402,N_7383);
nor U7665 (N_7665,N_7281,N_7310);
or U7666 (N_7666,N_7271,N_7404);
nand U7667 (N_7667,N_7282,N_7353);
or U7668 (N_7668,N_7348,N_7282);
nor U7669 (N_7669,N_7486,N_7354);
and U7670 (N_7670,N_7276,N_7338);
nand U7671 (N_7671,N_7457,N_7439);
nand U7672 (N_7672,N_7354,N_7363);
or U7673 (N_7673,N_7276,N_7413);
nand U7674 (N_7674,N_7488,N_7302);
or U7675 (N_7675,N_7313,N_7485);
and U7676 (N_7676,N_7376,N_7368);
and U7677 (N_7677,N_7335,N_7372);
nor U7678 (N_7678,N_7354,N_7467);
nand U7679 (N_7679,N_7404,N_7414);
nand U7680 (N_7680,N_7382,N_7413);
nor U7681 (N_7681,N_7387,N_7292);
and U7682 (N_7682,N_7273,N_7267);
or U7683 (N_7683,N_7310,N_7394);
and U7684 (N_7684,N_7360,N_7287);
or U7685 (N_7685,N_7387,N_7315);
xor U7686 (N_7686,N_7326,N_7417);
nand U7687 (N_7687,N_7411,N_7251);
nor U7688 (N_7688,N_7253,N_7499);
and U7689 (N_7689,N_7395,N_7466);
nand U7690 (N_7690,N_7371,N_7296);
or U7691 (N_7691,N_7482,N_7490);
or U7692 (N_7692,N_7255,N_7457);
nand U7693 (N_7693,N_7284,N_7293);
nand U7694 (N_7694,N_7391,N_7306);
and U7695 (N_7695,N_7285,N_7415);
nor U7696 (N_7696,N_7454,N_7363);
nor U7697 (N_7697,N_7351,N_7316);
and U7698 (N_7698,N_7428,N_7453);
nor U7699 (N_7699,N_7364,N_7288);
and U7700 (N_7700,N_7294,N_7269);
and U7701 (N_7701,N_7366,N_7399);
nand U7702 (N_7702,N_7478,N_7265);
nor U7703 (N_7703,N_7266,N_7312);
nand U7704 (N_7704,N_7311,N_7440);
nor U7705 (N_7705,N_7268,N_7414);
and U7706 (N_7706,N_7404,N_7284);
nor U7707 (N_7707,N_7389,N_7450);
and U7708 (N_7708,N_7450,N_7485);
and U7709 (N_7709,N_7477,N_7291);
nor U7710 (N_7710,N_7421,N_7305);
and U7711 (N_7711,N_7356,N_7350);
or U7712 (N_7712,N_7394,N_7487);
or U7713 (N_7713,N_7308,N_7350);
nand U7714 (N_7714,N_7391,N_7439);
or U7715 (N_7715,N_7276,N_7358);
or U7716 (N_7716,N_7429,N_7252);
nor U7717 (N_7717,N_7463,N_7447);
nor U7718 (N_7718,N_7494,N_7320);
nand U7719 (N_7719,N_7403,N_7271);
and U7720 (N_7720,N_7277,N_7307);
nor U7721 (N_7721,N_7433,N_7335);
and U7722 (N_7722,N_7444,N_7400);
nor U7723 (N_7723,N_7283,N_7284);
nor U7724 (N_7724,N_7283,N_7342);
or U7725 (N_7725,N_7384,N_7412);
xor U7726 (N_7726,N_7310,N_7429);
nor U7727 (N_7727,N_7449,N_7470);
or U7728 (N_7728,N_7293,N_7344);
or U7729 (N_7729,N_7292,N_7455);
and U7730 (N_7730,N_7251,N_7418);
or U7731 (N_7731,N_7419,N_7252);
or U7732 (N_7732,N_7337,N_7308);
and U7733 (N_7733,N_7493,N_7311);
xnor U7734 (N_7734,N_7386,N_7470);
nand U7735 (N_7735,N_7375,N_7268);
nand U7736 (N_7736,N_7493,N_7294);
nor U7737 (N_7737,N_7336,N_7444);
nand U7738 (N_7738,N_7475,N_7492);
and U7739 (N_7739,N_7423,N_7443);
and U7740 (N_7740,N_7280,N_7464);
or U7741 (N_7741,N_7333,N_7483);
or U7742 (N_7742,N_7250,N_7377);
or U7743 (N_7743,N_7344,N_7482);
nand U7744 (N_7744,N_7456,N_7390);
nand U7745 (N_7745,N_7270,N_7403);
and U7746 (N_7746,N_7486,N_7311);
or U7747 (N_7747,N_7456,N_7349);
or U7748 (N_7748,N_7450,N_7333);
or U7749 (N_7749,N_7385,N_7452);
and U7750 (N_7750,N_7660,N_7639);
or U7751 (N_7751,N_7681,N_7637);
nor U7752 (N_7752,N_7705,N_7718);
or U7753 (N_7753,N_7563,N_7539);
nand U7754 (N_7754,N_7500,N_7561);
nand U7755 (N_7755,N_7601,N_7590);
or U7756 (N_7756,N_7679,N_7710);
and U7757 (N_7757,N_7592,N_7525);
and U7758 (N_7758,N_7701,N_7613);
nand U7759 (N_7759,N_7565,N_7627);
nand U7760 (N_7760,N_7723,N_7519);
or U7761 (N_7761,N_7673,N_7547);
nor U7762 (N_7762,N_7657,N_7595);
nor U7763 (N_7763,N_7686,N_7618);
or U7764 (N_7764,N_7584,N_7650);
nor U7765 (N_7765,N_7535,N_7581);
and U7766 (N_7766,N_7505,N_7544);
nor U7767 (N_7767,N_7739,N_7645);
nand U7768 (N_7768,N_7576,N_7514);
and U7769 (N_7769,N_7522,N_7672);
and U7770 (N_7770,N_7731,N_7633);
xor U7771 (N_7771,N_7702,N_7588);
nor U7772 (N_7772,N_7598,N_7564);
or U7773 (N_7773,N_7740,N_7502);
nand U7774 (N_7774,N_7724,N_7720);
nand U7775 (N_7775,N_7621,N_7693);
or U7776 (N_7776,N_7506,N_7725);
nand U7777 (N_7777,N_7518,N_7680);
and U7778 (N_7778,N_7537,N_7741);
nor U7779 (N_7779,N_7512,N_7656);
or U7780 (N_7780,N_7682,N_7596);
nor U7781 (N_7781,N_7623,N_7735);
nor U7782 (N_7782,N_7714,N_7593);
nand U7783 (N_7783,N_7675,N_7520);
nor U7784 (N_7784,N_7614,N_7607);
nor U7785 (N_7785,N_7662,N_7635);
or U7786 (N_7786,N_7553,N_7638);
nor U7787 (N_7787,N_7580,N_7556);
nor U7788 (N_7788,N_7669,N_7634);
nand U7789 (N_7789,N_7543,N_7533);
nor U7790 (N_7790,N_7515,N_7549);
or U7791 (N_7791,N_7600,N_7641);
and U7792 (N_7792,N_7732,N_7636);
and U7793 (N_7793,N_7659,N_7610);
or U7794 (N_7794,N_7625,N_7670);
or U7795 (N_7795,N_7643,N_7713);
or U7796 (N_7796,N_7524,N_7697);
nor U7797 (N_7797,N_7632,N_7742);
or U7798 (N_7798,N_7619,N_7729);
nand U7799 (N_7799,N_7716,N_7648);
or U7800 (N_7800,N_7726,N_7651);
nor U7801 (N_7801,N_7616,N_7597);
and U7802 (N_7802,N_7738,N_7579);
nand U7803 (N_7803,N_7568,N_7667);
nor U7804 (N_7804,N_7622,N_7575);
and U7805 (N_7805,N_7583,N_7629);
nand U7806 (N_7806,N_7604,N_7691);
or U7807 (N_7807,N_7715,N_7699);
nor U7808 (N_7808,N_7559,N_7717);
and U7809 (N_7809,N_7586,N_7507);
nand U7810 (N_7810,N_7552,N_7516);
nand U7811 (N_7811,N_7501,N_7671);
or U7812 (N_7812,N_7529,N_7689);
or U7813 (N_7813,N_7571,N_7570);
and U7814 (N_7814,N_7737,N_7555);
or U7815 (N_7815,N_7644,N_7599);
and U7816 (N_7816,N_7594,N_7646);
and U7817 (N_7817,N_7708,N_7608);
nand U7818 (N_7818,N_7676,N_7719);
nand U7819 (N_7819,N_7692,N_7655);
or U7820 (N_7820,N_7538,N_7626);
and U7821 (N_7821,N_7589,N_7558);
or U7822 (N_7822,N_7703,N_7749);
nor U7823 (N_7823,N_7508,N_7711);
and U7824 (N_7824,N_7536,N_7678);
and U7825 (N_7825,N_7513,N_7747);
nor U7826 (N_7826,N_7523,N_7569);
or U7827 (N_7827,N_7685,N_7603);
nand U7828 (N_7828,N_7652,N_7649);
and U7829 (N_7829,N_7542,N_7688);
or U7830 (N_7830,N_7728,N_7540);
nand U7831 (N_7831,N_7528,N_7521);
and U7832 (N_7832,N_7574,N_7527);
nor U7833 (N_7833,N_7609,N_7587);
nand U7834 (N_7834,N_7577,N_7628);
nor U7835 (N_7835,N_7695,N_7606);
or U7836 (N_7836,N_7722,N_7712);
or U7837 (N_7837,N_7582,N_7630);
nand U7838 (N_7838,N_7698,N_7510);
and U7839 (N_7839,N_7530,N_7677);
and U7840 (N_7840,N_7545,N_7642);
and U7841 (N_7841,N_7572,N_7504);
and U7842 (N_7842,N_7707,N_7709);
and U7843 (N_7843,N_7573,N_7548);
or U7844 (N_7844,N_7663,N_7733);
nor U7845 (N_7845,N_7605,N_7744);
nand U7846 (N_7846,N_7509,N_7661);
nor U7847 (N_7847,N_7531,N_7612);
nor U7848 (N_7848,N_7578,N_7700);
or U7849 (N_7849,N_7541,N_7734);
or U7850 (N_7850,N_7684,N_7551);
or U7851 (N_7851,N_7666,N_7664);
and U7852 (N_7852,N_7550,N_7745);
and U7853 (N_7853,N_7727,N_7591);
nor U7854 (N_7854,N_7736,N_7746);
nor U7855 (N_7855,N_7503,N_7654);
nor U7856 (N_7856,N_7585,N_7721);
and U7857 (N_7857,N_7694,N_7687);
or U7858 (N_7858,N_7706,N_7532);
nor U7859 (N_7859,N_7730,N_7631);
and U7860 (N_7860,N_7704,N_7658);
and U7861 (N_7861,N_7640,N_7611);
or U7862 (N_7862,N_7567,N_7511);
nand U7863 (N_7863,N_7560,N_7534);
and U7864 (N_7864,N_7554,N_7624);
or U7865 (N_7865,N_7615,N_7647);
and U7866 (N_7866,N_7696,N_7562);
and U7867 (N_7867,N_7617,N_7743);
nand U7868 (N_7868,N_7602,N_7690);
or U7869 (N_7869,N_7668,N_7674);
nor U7870 (N_7870,N_7683,N_7546);
or U7871 (N_7871,N_7517,N_7665);
or U7872 (N_7872,N_7620,N_7748);
nor U7873 (N_7873,N_7526,N_7566);
nand U7874 (N_7874,N_7653,N_7557);
and U7875 (N_7875,N_7678,N_7745);
nor U7876 (N_7876,N_7603,N_7716);
and U7877 (N_7877,N_7736,N_7690);
nand U7878 (N_7878,N_7677,N_7703);
and U7879 (N_7879,N_7578,N_7702);
or U7880 (N_7880,N_7654,N_7599);
nand U7881 (N_7881,N_7527,N_7532);
and U7882 (N_7882,N_7519,N_7510);
or U7883 (N_7883,N_7684,N_7614);
nand U7884 (N_7884,N_7690,N_7604);
nor U7885 (N_7885,N_7708,N_7690);
and U7886 (N_7886,N_7602,N_7715);
nor U7887 (N_7887,N_7528,N_7602);
nand U7888 (N_7888,N_7565,N_7609);
nor U7889 (N_7889,N_7722,N_7718);
nand U7890 (N_7890,N_7554,N_7555);
nand U7891 (N_7891,N_7662,N_7667);
and U7892 (N_7892,N_7604,N_7637);
nand U7893 (N_7893,N_7511,N_7537);
and U7894 (N_7894,N_7599,N_7699);
nand U7895 (N_7895,N_7670,N_7513);
and U7896 (N_7896,N_7580,N_7684);
or U7897 (N_7897,N_7671,N_7607);
and U7898 (N_7898,N_7591,N_7613);
and U7899 (N_7899,N_7600,N_7700);
nor U7900 (N_7900,N_7699,N_7504);
or U7901 (N_7901,N_7580,N_7523);
xor U7902 (N_7902,N_7722,N_7671);
or U7903 (N_7903,N_7717,N_7516);
nor U7904 (N_7904,N_7641,N_7631);
or U7905 (N_7905,N_7579,N_7630);
and U7906 (N_7906,N_7600,N_7689);
nor U7907 (N_7907,N_7748,N_7557);
or U7908 (N_7908,N_7670,N_7616);
and U7909 (N_7909,N_7676,N_7574);
nor U7910 (N_7910,N_7626,N_7725);
nand U7911 (N_7911,N_7568,N_7642);
nor U7912 (N_7912,N_7542,N_7538);
nand U7913 (N_7913,N_7530,N_7612);
and U7914 (N_7914,N_7720,N_7521);
nand U7915 (N_7915,N_7713,N_7690);
nand U7916 (N_7916,N_7622,N_7609);
and U7917 (N_7917,N_7510,N_7623);
nor U7918 (N_7918,N_7688,N_7673);
or U7919 (N_7919,N_7624,N_7507);
nor U7920 (N_7920,N_7613,N_7639);
nor U7921 (N_7921,N_7745,N_7505);
or U7922 (N_7922,N_7729,N_7552);
nor U7923 (N_7923,N_7582,N_7605);
nor U7924 (N_7924,N_7718,N_7720);
and U7925 (N_7925,N_7647,N_7518);
nand U7926 (N_7926,N_7677,N_7604);
nor U7927 (N_7927,N_7725,N_7736);
or U7928 (N_7928,N_7550,N_7669);
nand U7929 (N_7929,N_7521,N_7612);
or U7930 (N_7930,N_7535,N_7651);
nor U7931 (N_7931,N_7593,N_7719);
nor U7932 (N_7932,N_7691,N_7616);
or U7933 (N_7933,N_7539,N_7704);
nand U7934 (N_7934,N_7651,N_7599);
nand U7935 (N_7935,N_7731,N_7503);
or U7936 (N_7936,N_7626,N_7621);
nor U7937 (N_7937,N_7693,N_7500);
xor U7938 (N_7938,N_7662,N_7733);
and U7939 (N_7939,N_7533,N_7664);
nand U7940 (N_7940,N_7684,N_7675);
and U7941 (N_7941,N_7540,N_7518);
or U7942 (N_7942,N_7653,N_7741);
and U7943 (N_7943,N_7725,N_7568);
and U7944 (N_7944,N_7618,N_7644);
nor U7945 (N_7945,N_7682,N_7709);
nor U7946 (N_7946,N_7662,N_7525);
or U7947 (N_7947,N_7726,N_7538);
nor U7948 (N_7948,N_7606,N_7555);
nor U7949 (N_7949,N_7740,N_7573);
and U7950 (N_7950,N_7692,N_7560);
xnor U7951 (N_7951,N_7641,N_7652);
and U7952 (N_7952,N_7525,N_7504);
nand U7953 (N_7953,N_7636,N_7662);
and U7954 (N_7954,N_7568,N_7744);
and U7955 (N_7955,N_7633,N_7595);
nor U7956 (N_7956,N_7669,N_7583);
nand U7957 (N_7957,N_7654,N_7543);
or U7958 (N_7958,N_7682,N_7623);
or U7959 (N_7959,N_7684,N_7628);
xnor U7960 (N_7960,N_7579,N_7590);
nand U7961 (N_7961,N_7597,N_7613);
and U7962 (N_7962,N_7618,N_7612);
nor U7963 (N_7963,N_7512,N_7573);
xnor U7964 (N_7964,N_7728,N_7605);
nor U7965 (N_7965,N_7505,N_7510);
nor U7966 (N_7966,N_7635,N_7735);
nand U7967 (N_7967,N_7657,N_7682);
and U7968 (N_7968,N_7683,N_7607);
and U7969 (N_7969,N_7510,N_7693);
or U7970 (N_7970,N_7676,N_7577);
or U7971 (N_7971,N_7515,N_7703);
and U7972 (N_7972,N_7651,N_7517);
or U7973 (N_7973,N_7566,N_7580);
or U7974 (N_7974,N_7701,N_7587);
or U7975 (N_7975,N_7748,N_7664);
nor U7976 (N_7976,N_7612,N_7716);
nand U7977 (N_7977,N_7634,N_7525);
nand U7978 (N_7978,N_7682,N_7553);
or U7979 (N_7979,N_7702,N_7617);
or U7980 (N_7980,N_7549,N_7659);
nor U7981 (N_7981,N_7610,N_7661);
or U7982 (N_7982,N_7702,N_7546);
or U7983 (N_7983,N_7688,N_7575);
or U7984 (N_7984,N_7530,N_7667);
nor U7985 (N_7985,N_7546,N_7649);
xor U7986 (N_7986,N_7709,N_7640);
and U7987 (N_7987,N_7673,N_7517);
nor U7988 (N_7988,N_7517,N_7568);
nor U7989 (N_7989,N_7502,N_7646);
and U7990 (N_7990,N_7534,N_7743);
and U7991 (N_7991,N_7658,N_7713);
nor U7992 (N_7992,N_7584,N_7660);
nand U7993 (N_7993,N_7648,N_7531);
and U7994 (N_7994,N_7717,N_7694);
nor U7995 (N_7995,N_7682,N_7614);
or U7996 (N_7996,N_7653,N_7702);
and U7997 (N_7997,N_7640,N_7627);
and U7998 (N_7998,N_7598,N_7606);
nand U7999 (N_7999,N_7527,N_7657);
nand U8000 (N_8000,N_7841,N_7902);
or U8001 (N_8001,N_7949,N_7942);
and U8002 (N_8002,N_7907,N_7803);
nor U8003 (N_8003,N_7926,N_7781);
nand U8004 (N_8004,N_7912,N_7786);
and U8005 (N_8005,N_7915,N_7764);
nand U8006 (N_8006,N_7796,N_7779);
nand U8007 (N_8007,N_7819,N_7852);
nand U8008 (N_8008,N_7883,N_7989);
nand U8009 (N_8009,N_7999,N_7800);
and U8010 (N_8010,N_7821,N_7900);
nand U8011 (N_8011,N_7775,N_7817);
and U8012 (N_8012,N_7911,N_7863);
or U8013 (N_8013,N_7997,N_7771);
or U8014 (N_8014,N_7832,N_7901);
and U8015 (N_8015,N_7801,N_7844);
nand U8016 (N_8016,N_7857,N_7904);
nand U8017 (N_8017,N_7964,N_7856);
nor U8018 (N_8018,N_7979,N_7908);
nor U8019 (N_8019,N_7961,N_7892);
or U8020 (N_8020,N_7935,N_7778);
or U8021 (N_8021,N_7957,N_7939);
nand U8022 (N_8022,N_7797,N_7916);
nor U8023 (N_8023,N_7931,N_7820);
and U8024 (N_8024,N_7766,N_7898);
nor U8025 (N_8025,N_7816,N_7962);
nor U8026 (N_8026,N_7885,N_7802);
or U8027 (N_8027,N_7910,N_7823);
and U8028 (N_8028,N_7763,N_7891);
and U8029 (N_8029,N_7782,N_7993);
or U8030 (N_8030,N_7808,N_7991);
nor U8031 (N_8031,N_7869,N_7897);
nand U8032 (N_8032,N_7947,N_7861);
nand U8033 (N_8033,N_7970,N_7951);
and U8034 (N_8034,N_7813,N_7804);
and U8035 (N_8035,N_7758,N_7812);
nor U8036 (N_8036,N_7944,N_7965);
or U8037 (N_8037,N_7868,N_7994);
nor U8038 (N_8038,N_7762,N_7930);
and U8039 (N_8039,N_7793,N_7811);
nand U8040 (N_8040,N_7756,N_7806);
and U8041 (N_8041,N_7919,N_7855);
nor U8042 (N_8042,N_7822,N_7995);
or U8043 (N_8043,N_7848,N_7975);
and U8044 (N_8044,N_7952,N_7825);
nand U8045 (N_8045,N_7946,N_7830);
and U8046 (N_8046,N_7770,N_7966);
and U8047 (N_8047,N_7988,N_7978);
nor U8048 (N_8048,N_7838,N_7909);
nand U8049 (N_8049,N_7761,N_7789);
nand U8050 (N_8050,N_7923,N_7788);
nand U8051 (N_8051,N_7889,N_7750);
nand U8052 (N_8052,N_7887,N_7953);
nor U8053 (N_8053,N_7851,N_7794);
or U8054 (N_8054,N_7922,N_7928);
or U8055 (N_8055,N_7847,N_7877);
nor U8056 (N_8056,N_7974,N_7850);
or U8057 (N_8057,N_7876,N_7914);
nand U8058 (N_8058,N_7780,N_7809);
nor U8059 (N_8059,N_7945,N_7969);
and U8060 (N_8060,N_7843,N_7878);
xnor U8061 (N_8061,N_7867,N_7872);
or U8062 (N_8062,N_7906,N_7984);
nand U8063 (N_8063,N_7996,N_7846);
or U8064 (N_8064,N_7772,N_7929);
and U8065 (N_8065,N_7981,N_7829);
nand U8066 (N_8066,N_7774,N_7977);
and U8067 (N_8067,N_7976,N_7913);
nand U8068 (N_8068,N_7893,N_7888);
and U8069 (N_8069,N_7757,N_7986);
and U8070 (N_8070,N_7787,N_7955);
nor U8071 (N_8071,N_7769,N_7881);
and U8072 (N_8072,N_7920,N_7840);
nand U8073 (N_8073,N_7973,N_7783);
nand U8074 (N_8074,N_7784,N_7870);
or U8075 (N_8075,N_7773,N_7948);
nand U8076 (N_8076,N_7814,N_7862);
and U8077 (N_8077,N_7836,N_7776);
and U8078 (N_8078,N_7983,N_7967);
nand U8079 (N_8079,N_7932,N_7925);
nand U8080 (N_8080,N_7968,N_7858);
nand U8081 (N_8081,N_7890,N_7971);
nand U8082 (N_8082,N_7859,N_7799);
nand U8083 (N_8083,N_7835,N_7972);
and U8084 (N_8084,N_7950,N_7767);
or U8085 (N_8085,N_7864,N_7818);
nand U8086 (N_8086,N_7815,N_7755);
or U8087 (N_8087,N_7896,N_7936);
nand U8088 (N_8088,N_7791,N_7751);
and U8089 (N_8089,N_7954,N_7826);
or U8090 (N_8090,N_7894,N_7866);
nand U8091 (N_8091,N_7798,N_7795);
and U8092 (N_8092,N_7886,N_7963);
and U8093 (N_8093,N_7845,N_7992);
and U8094 (N_8094,N_7768,N_7918);
and U8095 (N_8095,N_7760,N_7985);
and U8096 (N_8096,N_7927,N_7940);
or U8097 (N_8097,N_7810,N_7871);
nor U8098 (N_8098,N_7873,N_7837);
nor U8099 (N_8099,N_7934,N_7792);
nand U8100 (N_8100,N_7941,N_7924);
and U8101 (N_8101,N_7938,N_7827);
or U8102 (N_8102,N_7880,N_7754);
or U8103 (N_8103,N_7853,N_7865);
nand U8104 (N_8104,N_7958,N_7960);
or U8105 (N_8105,N_7903,N_7839);
nor U8106 (N_8106,N_7785,N_7842);
and U8107 (N_8107,N_7882,N_7854);
and U8108 (N_8108,N_7759,N_7752);
and U8109 (N_8109,N_7753,N_7921);
nand U8110 (N_8110,N_7805,N_7982);
nor U8111 (N_8111,N_7875,N_7895);
and U8112 (N_8112,N_7849,N_7943);
nor U8113 (N_8113,N_7874,N_7998);
and U8114 (N_8114,N_7765,N_7990);
nor U8115 (N_8115,N_7833,N_7956);
nand U8116 (N_8116,N_7824,N_7980);
and U8117 (N_8117,N_7905,N_7831);
and U8118 (N_8118,N_7937,N_7879);
nor U8119 (N_8119,N_7834,N_7860);
and U8120 (N_8120,N_7933,N_7777);
or U8121 (N_8121,N_7828,N_7790);
or U8122 (N_8122,N_7917,N_7899);
and U8123 (N_8123,N_7959,N_7884);
nor U8124 (N_8124,N_7987,N_7807);
nand U8125 (N_8125,N_7814,N_7882);
nor U8126 (N_8126,N_7858,N_7880);
or U8127 (N_8127,N_7792,N_7785);
nor U8128 (N_8128,N_7867,N_7799);
and U8129 (N_8129,N_7798,N_7962);
or U8130 (N_8130,N_7827,N_7977);
nand U8131 (N_8131,N_7787,N_7927);
nand U8132 (N_8132,N_7803,N_7983);
nand U8133 (N_8133,N_7808,N_7969);
nand U8134 (N_8134,N_7902,N_7839);
nand U8135 (N_8135,N_7964,N_7817);
nor U8136 (N_8136,N_7856,N_7762);
and U8137 (N_8137,N_7814,N_7917);
or U8138 (N_8138,N_7935,N_7762);
and U8139 (N_8139,N_7981,N_7797);
and U8140 (N_8140,N_7881,N_7820);
nor U8141 (N_8141,N_7974,N_7961);
nor U8142 (N_8142,N_7903,N_7850);
or U8143 (N_8143,N_7995,N_7946);
nor U8144 (N_8144,N_7860,N_7762);
and U8145 (N_8145,N_7927,N_7917);
nand U8146 (N_8146,N_7971,N_7921);
or U8147 (N_8147,N_7844,N_7897);
nor U8148 (N_8148,N_7960,N_7822);
or U8149 (N_8149,N_7995,N_7910);
nand U8150 (N_8150,N_7796,N_7910);
nand U8151 (N_8151,N_7761,N_7891);
or U8152 (N_8152,N_7768,N_7985);
or U8153 (N_8153,N_7905,N_7859);
nand U8154 (N_8154,N_7981,N_7951);
and U8155 (N_8155,N_7796,N_7917);
and U8156 (N_8156,N_7806,N_7771);
or U8157 (N_8157,N_7785,N_7789);
nor U8158 (N_8158,N_7765,N_7924);
nor U8159 (N_8159,N_7798,N_7988);
nand U8160 (N_8160,N_7775,N_7871);
and U8161 (N_8161,N_7922,N_7967);
or U8162 (N_8162,N_7954,N_7977);
nand U8163 (N_8163,N_7968,N_7800);
nor U8164 (N_8164,N_7774,N_7938);
nand U8165 (N_8165,N_7824,N_7773);
nor U8166 (N_8166,N_7929,N_7763);
or U8167 (N_8167,N_7811,N_7787);
nor U8168 (N_8168,N_7860,N_7957);
xor U8169 (N_8169,N_7824,N_7791);
and U8170 (N_8170,N_7754,N_7926);
nor U8171 (N_8171,N_7803,N_7856);
nor U8172 (N_8172,N_7805,N_7838);
nor U8173 (N_8173,N_7977,N_7825);
nand U8174 (N_8174,N_7917,N_7863);
nor U8175 (N_8175,N_7975,N_7822);
nand U8176 (N_8176,N_7842,N_7997);
and U8177 (N_8177,N_7970,N_7947);
xnor U8178 (N_8178,N_7903,N_7920);
nor U8179 (N_8179,N_7898,N_7829);
and U8180 (N_8180,N_7967,N_7923);
nor U8181 (N_8181,N_7817,N_7848);
and U8182 (N_8182,N_7913,N_7793);
nand U8183 (N_8183,N_7891,N_7931);
or U8184 (N_8184,N_7965,N_7797);
nand U8185 (N_8185,N_7846,N_7839);
and U8186 (N_8186,N_7884,N_7753);
or U8187 (N_8187,N_7781,N_7892);
and U8188 (N_8188,N_7924,N_7915);
nor U8189 (N_8189,N_7816,N_7909);
or U8190 (N_8190,N_7968,N_7814);
nor U8191 (N_8191,N_7906,N_7879);
nand U8192 (N_8192,N_7927,N_7831);
nor U8193 (N_8193,N_7949,N_7960);
and U8194 (N_8194,N_7866,N_7951);
and U8195 (N_8195,N_7853,N_7920);
or U8196 (N_8196,N_7784,N_7817);
nand U8197 (N_8197,N_7847,N_7971);
nor U8198 (N_8198,N_7868,N_7921);
nor U8199 (N_8199,N_7998,N_7836);
nor U8200 (N_8200,N_7903,N_7935);
or U8201 (N_8201,N_7786,N_7799);
and U8202 (N_8202,N_7891,N_7756);
or U8203 (N_8203,N_7888,N_7973);
nand U8204 (N_8204,N_7828,N_7781);
or U8205 (N_8205,N_7934,N_7774);
nor U8206 (N_8206,N_7750,N_7976);
or U8207 (N_8207,N_7843,N_7890);
and U8208 (N_8208,N_7755,N_7974);
nor U8209 (N_8209,N_7947,N_7881);
and U8210 (N_8210,N_7811,N_7893);
and U8211 (N_8211,N_7774,N_7762);
nor U8212 (N_8212,N_7962,N_7957);
nor U8213 (N_8213,N_7802,N_7977);
or U8214 (N_8214,N_7779,N_7996);
or U8215 (N_8215,N_7958,N_7929);
nor U8216 (N_8216,N_7853,N_7841);
nor U8217 (N_8217,N_7884,N_7954);
nand U8218 (N_8218,N_7832,N_7885);
or U8219 (N_8219,N_7753,N_7880);
nor U8220 (N_8220,N_7898,N_7875);
or U8221 (N_8221,N_7976,N_7828);
nor U8222 (N_8222,N_7778,N_7967);
nor U8223 (N_8223,N_7812,N_7926);
nor U8224 (N_8224,N_7788,N_7818);
nor U8225 (N_8225,N_7976,N_7818);
and U8226 (N_8226,N_7888,N_7787);
and U8227 (N_8227,N_7752,N_7903);
nand U8228 (N_8228,N_7851,N_7953);
or U8229 (N_8229,N_7800,N_7825);
nor U8230 (N_8230,N_7759,N_7959);
nand U8231 (N_8231,N_7952,N_7843);
nand U8232 (N_8232,N_7769,N_7892);
and U8233 (N_8233,N_7999,N_7965);
and U8234 (N_8234,N_7777,N_7840);
or U8235 (N_8235,N_7792,N_7905);
or U8236 (N_8236,N_7982,N_7845);
nor U8237 (N_8237,N_7839,N_7813);
and U8238 (N_8238,N_7846,N_7874);
nand U8239 (N_8239,N_7798,N_7991);
nand U8240 (N_8240,N_7806,N_7818);
and U8241 (N_8241,N_7907,N_7994);
and U8242 (N_8242,N_7811,N_7937);
and U8243 (N_8243,N_7911,N_7930);
nand U8244 (N_8244,N_7971,N_7767);
nand U8245 (N_8245,N_7878,N_7914);
or U8246 (N_8246,N_7819,N_7833);
and U8247 (N_8247,N_7999,N_7783);
or U8248 (N_8248,N_7998,N_7869);
nand U8249 (N_8249,N_7960,N_7961);
nand U8250 (N_8250,N_8237,N_8096);
nor U8251 (N_8251,N_8236,N_8067);
and U8252 (N_8252,N_8156,N_8186);
nand U8253 (N_8253,N_8053,N_8111);
nor U8254 (N_8254,N_8235,N_8201);
nand U8255 (N_8255,N_8182,N_8208);
and U8256 (N_8256,N_8195,N_8026);
or U8257 (N_8257,N_8037,N_8017);
or U8258 (N_8258,N_8179,N_8152);
nand U8259 (N_8259,N_8183,N_8242);
or U8260 (N_8260,N_8094,N_8046);
nand U8261 (N_8261,N_8103,N_8151);
and U8262 (N_8262,N_8014,N_8131);
and U8263 (N_8263,N_8013,N_8097);
or U8264 (N_8264,N_8190,N_8185);
nor U8265 (N_8265,N_8114,N_8052);
or U8266 (N_8266,N_8064,N_8089);
or U8267 (N_8267,N_8104,N_8193);
nor U8268 (N_8268,N_8184,N_8132);
and U8269 (N_8269,N_8044,N_8091);
nor U8270 (N_8270,N_8061,N_8161);
and U8271 (N_8271,N_8233,N_8115);
nor U8272 (N_8272,N_8088,N_8136);
nor U8273 (N_8273,N_8058,N_8194);
nor U8274 (N_8274,N_8117,N_8125);
nand U8275 (N_8275,N_8055,N_8139);
nand U8276 (N_8276,N_8138,N_8223);
and U8277 (N_8277,N_8134,N_8234);
nand U8278 (N_8278,N_8015,N_8051);
or U8279 (N_8279,N_8016,N_8215);
or U8280 (N_8280,N_8021,N_8245);
or U8281 (N_8281,N_8042,N_8227);
and U8282 (N_8282,N_8027,N_8118);
nor U8283 (N_8283,N_8168,N_8098);
or U8284 (N_8284,N_8011,N_8211);
nor U8285 (N_8285,N_8188,N_8174);
nor U8286 (N_8286,N_8084,N_8028);
and U8287 (N_8287,N_8248,N_8197);
and U8288 (N_8288,N_8191,N_8092);
or U8289 (N_8289,N_8126,N_8112);
or U8290 (N_8290,N_8203,N_8080);
nor U8291 (N_8291,N_8169,N_8085);
or U8292 (N_8292,N_8124,N_8229);
or U8293 (N_8293,N_8217,N_8108);
nor U8294 (N_8294,N_8231,N_8249);
nand U8295 (N_8295,N_8012,N_8214);
or U8296 (N_8296,N_8207,N_8110);
nand U8297 (N_8297,N_8120,N_8142);
or U8298 (N_8298,N_8130,N_8218);
or U8299 (N_8299,N_8150,N_8005);
nand U8300 (N_8300,N_8222,N_8240);
and U8301 (N_8301,N_8070,N_8004);
and U8302 (N_8302,N_8057,N_8221);
or U8303 (N_8303,N_8119,N_8239);
or U8304 (N_8304,N_8153,N_8060);
nor U8305 (N_8305,N_8148,N_8128);
and U8306 (N_8306,N_8204,N_8178);
xnor U8307 (N_8307,N_8047,N_8025);
or U8308 (N_8308,N_8228,N_8009);
or U8309 (N_8309,N_8087,N_8160);
nor U8310 (N_8310,N_8083,N_8166);
or U8311 (N_8311,N_8145,N_8196);
nand U8312 (N_8312,N_8158,N_8045);
and U8313 (N_8313,N_8140,N_8069);
nor U8314 (N_8314,N_8147,N_8225);
nand U8315 (N_8315,N_8090,N_8059);
nor U8316 (N_8316,N_8146,N_8036);
nor U8317 (N_8317,N_8020,N_8007);
and U8318 (N_8318,N_8238,N_8167);
and U8319 (N_8319,N_8056,N_8206);
nand U8320 (N_8320,N_8181,N_8008);
nand U8321 (N_8321,N_8212,N_8122);
nand U8322 (N_8322,N_8006,N_8003);
and U8323 (N_8323,N_8241,N_8200);
nor U8324 (N_8324,N_8062,N_8162);
nor U8325 (N_8325,N_8232,N_8127);
and U8326 (N_8326,N_8081,N_8086);
nor U8327 (N_8327,N_8198,N_8116);
nor U8328 (N_8328,N_8244,N_8077);
nand U8329 (N_8329,N_8010,N_8105);
nand U8330 (N_8330,N_8023,N_8187);
and U8331 (N_8331,N_8192,N_8068);
nand U8332 (N_8332,N_8209,N_8079);
and U8333 (N_8333,N_8071,N_8177);
or U8334 (N_8334,N_8101,N_8219);
nand U8335 (N_8335,N_8180,N_8173);
or U8336 (N_8336,N_8199,N_8159);
nor U8337 (N_8337,N_8135,N_8246);
and U8338 (N_8338,N_8141,N_8066);
nand U8339 (N_8339,N_8022,N_8106);
xor U8340 (N_8340,N_8018,N_8076);
or U8341 (N_8341,N_8082,N_8224);
or U8342 (N_8342,N_8247,N_8073);
or U8343 (N_8343,N_8133,N_8107);
and U8344 (N_8344,N_8202,N_8001);
nand U8345 (N_8345,N_8048,N_8050);
and U8346 (N_8346,N_8220,N_8170);
nor U8347 (N_8347,N_8034,N_8129);
nand U8348 (N_8348,N_8172,N_8109);
and U8349 (N_8349,N_8137,N_8230);
or U8350 (N_8350,N_8155,N_8176);
and U8351 (N_8351,N_8019,N_8039);
and U8352 (N_8352,N_8024,N_8210);
or U8353 (N_8353,N_8075,N_8226);
nor U8354 (N_8354,N_8033,N_8093);
nand U8355 (N_8355,N_8165,N_8002);
or U8356 (N_8356,N_8175,N_8030);
nor U8357 (N_8357,N_8157,N_8078);
or U8358 (N_8358,N_8035,N_8205);
or U8359 (N_8359,N_8100,N_8243);
and U8360 (N_8360,N_8063,N_8032);
nand U8361 (N_8361,N_8095,N_8163);
nor U8362 (N_8362,N_8121,N_8031);
or U8363 (N_8363,N_8041,N_8149);
nand U8364 (N_8364,N_8154,N_8000);
nor U8365 (N_8365,N_8171,N_8040);
nand U8366 (N_8366,N_8123,N_8144);
nor U8367 (N_8367,N_8065,N_8074);
nand U8368 (N_8368,N_8099,N_8213);
nand U8369 (N_8369,N_8038,N_8189);
or U8370 (N_8370,N_8029,N_8216);
and U8371 (N_8371,N_8049,N_8043);
nor U8372 (N_8372,N_8164,N_8113);
nand U8373 (N_8373,N_8143,N_8102);
or U8374 (N_8374,N_8072,N_8054);
nor U8375 (N_8375,N_8223,N_8120);
nand U8376 (N_8376,N_8083,N_8122);
nor U8377 (N_8377,N_8134,N_8059);
and U8378 (N_8378,N_8069,N_8061);
and U8379 (N_8379,N_8239,N_8096);
or U8380 (N_8380,N_8178,N_8160);
nor U8381 (N_8381,N_8003,N_8117);
nand U8382 (N_8382,N_8062,N_8233);
or U8383 (N_8383,N_8120,N_8112);
nand U8384 (N_8384,N_8227,N_8044);
nand U8385 (N_8385,N_8126,N_8166);
and U8386 (N_8386,N_8097,N_8191);
or U8387 (N_8387,N_8105,N_8075);
nand U8388 (N_8388,N_8002,N_8162);
nor U8389 (N_8389,N_8110,N_8223);
and U8390 (N_8390,N_8059,N_8011);
or U8391 (N_8391,N_8191,N_8025);
nand U8392 (N_8392,N_8132,N_8106);
and U8393 (N_8393,N_8160,N_8162);
nor U8394 (N_8394,N_8178,N_8013);
nand U8395 (N_8395,N_8056,N_8077);
or U8396 (N_8396,N_8167,N_8197);
and U8397 (N_8397,N_8075,N_8130);
and U8398 (N_8398,N_8247,N_8077);
nor U8399 (N_8399,N_8205,N_8145);
nand U8400 (N_8400,N_8210,N_8145);
nand U8401 (N_8401,N_8119,N_8122);
or U8402 (N_8402,N_8185,N_8036);
or U8403 (N_8403,N_8160,N_8012);
nand U8404 (N_8404,N_8019,N_8162);
nand U8405 (N_8405,N_8070,N_8039);
and U8406 (N_8406,N_8163,N_8205);
and U8407 (N_8407,N_8069,N_8126);
nor U8408 (N_8408,N_8189,N_8030);
or U8409 (N_8409,N_8184,N_8090);
and U8410 (N_8410,N_8116,N_8076);
and U8411 (N_8411,N_8087,N_8021);
or U8412 (N_8412,N_8096,N_8193);
and U8413 (N_8413,N_8109,N_8166);
nor U8414 (N_8414,N_8110,N_8193);
nand U8415 (N_8415,N_8238,N_8091);
nand U8416 (N_8416,N_8114,N_8170);
and U8417 (N_8417,N_8229,N_8201);
nand U8418 (N_8418,N_8197,N_8210);
and U8419 (N_8419,N_8126,N_8188);
or U8420 (N_8420,N_8016,N_8047);
and U8421 (N_8421,N_8100,N_8084);
nand U8422 (N_8422,N_8197,N_8159);
nor U8423 (N_8423,N_8018,N_8012);
or U8424 (N_8424,N_8085,N_8221);
nor U8425 (N_8425,N_8100,N_8063);
or U8426 (N_8426,N_8222,N_8049);
nor U8427 (N_8427,N_8141,N_8214);
nand U8428 (N_8428,N_8052,N_8227);
nor U8429 (N_8429,N_8122,N_8053);
nor U8430 (N_8430,N_8079,N_8099);
nand U8431 (N_8431,N_8121,N_8101);
nor U8432 (N_8432,N_8228,N_8186);
nor U8433 (N_8433,N_8060,N_8058);
nor U8434 (N_8434,N_8105,N_8061);
and U8435 (N_8435,N_8218,N_8072);
and U8436 (N_8436,N_8127,N_8002);
nand U8437 (N_8437,N_8233,N_8133);
and U8438 (N_8438,N_8033,N_8122);
and U8439 (N_8439,N_8240,N_8025);
nor U8440 (N_8440,N_8065,N_8195);
nor U8441 (N_8441,N_8227,N_8134);
nor U8442 (N_8442,N_8206,N_8078);
or U8443 (N_8443,N_8180,N_8161);
nor U8444 (N_8444,N_8038,N_8160);
and U8445 (N_8445,N_8108,N_8070);
nor U8446 (N_8446,N_8160,N_8179);
nand U8447 (N_8447,N_8137,N_8075);
nor U8448 (N_8448,N_8237,N_8166);
and U8449 (N_8449,N_8215,N_8157);
nor U8450 (N_8450,N_8185,N_8133);
or U8451 (N_8451,N_8215,N_8119);
or U8452 (N_8452,N_8026,N_8174);
nor U8453 (N_8453,N_8043,N_8102);
or U8454 (N_8454,N_8081,N_8196);
and U8455 (N_8455,N_8043,N_8232);
nor U8456 (N_8456,N_8153,N_8152);
nor U8457 (N_8457,N_8057,N_8044);
nor U8458 (N_8458,N_8184,N_8148);
nand U8459 (N_8459,N_8056,N_8104);
nor U8460 (N_8460,N_8078,N_8052);
nand U8461 (N_8461,N_8190,N_8202);
nand U8462 (N_8462,N_8184,N_8129);
nand U8463 (N_8463,N_8061,N_8079);
nor U8464 (N_8464,N_8084,N_8121);
or U8465 (N_8465,N_8076,N_8204);
and U8466 (N_8466,N_8004,N_8096);
or U8467 (N_8467,N_8011,N_8062);
nor U8468 (N_8468,N_8202,N_8244);
or U8469 (N_8469,N_8024,N_8103);
or U8470 (N_8470,N_8203,N_8209);
nand U8471 (N_8471,N_8237,N_8004);
nand U8472 (N_8472,N_8044,N_8035);
nor U8473 (N_8473,N_8058,N_8011);
nor U8474 (N_8474,N_8134,N_8157);
or U8475 (N_8475,N_8049,N_8068);
nor U8476 (N_8476,N_8035,N_8063);
and U8477 (N_8477,N_8182,N_8054);
and U8478 (N_8478,N_8070,N_8020);
nand U8479 (N_8479,N_8134,N_8166);
nand U8480 (N_8480,N_8067,N_8009);
and U8481 (N_8481,N_8130,N_8028);
and U8482 (N_8482,N_8174,N_8233);
and U8483 (N_8483,N_8020,N_8016);
nand U8484 (N_8484,N_8069,N_8028);
or U8485 (N_8485,N_8068,N_8044);
or U8486 (N_8486,N_8113,N_8026);
nand U8487 (N_8487,N_8118,N_8046);
and U8488 (N_8488,N_8116,N_8235);
or U8489 (N_8489,N_8018,N_8064);
nor U8490 (N_8490,N_8137,N_8059);
nand U8491 (N_8491,N_8025,N_8100);
nor U8492 (N_8492,N_8070,N_8019);
or U8493 (N_8493,N_8046,N_8197);
nand U8494 (N_8494,N_8071,N_8007);
nor U8495 (N_8495,N_8071,N_8185);
or U8496 (N_8496,N_8177,N_8022);
nor U8497 (N_8497,N_8028,N_8117);
nand U8498 (N_8498,N_8021,N_8246);
nand U8499 (N_8499,N_8230,N_8005);
and U8500 (N_8500,N_8446,N_8364);
nand U8501 (N_8501,N_8318,N_8424);
and U8502 (N_8502,N_8469,N_8412);
nand U8503 (N_8503,N_8254,N_8397);
or U8504 (N_8504,N_8325,N_8336);
or U8505 (N_8505,N_8487,N_8294);
and U8506 (N_8506,N_8283,N_8423);
and U8507 (N_8507,N_8261,N_8298);
and U8508 (N_8508,N_8402,N_8489);
nand U8509 (N_8509,N_8281,N_8428);
and U8510 (N_8510,N_8253,N_8410);
or U8511 (N_8511,N_8356,N_8416);
nand U8512 (N_8512,N_8435,N_8250);
nor U8513 (N_8513,N_8386,N_8321);
or U8514 (N_8514,N_8484,N_8494);
nand U8515 (N_8515,N_8429,N_8344);
or U8516 (N_8516,N_8417,N_8268);
nand U8517 (N_8517,N_8251,N_8404);
or U8518 (N_8518,N_8300,N_8384);
nor U8519 (N_8519,N_8312,N_8320);
or U8520 (N_8520,N_8441,N_8473);
nand U8521 (N_8521,N_8290,N_8358);
or U8522 (N_8522,N_8490,N_8483);
and U8523 (N_8523,N_8276,N_8496);
and U8524 (N_8524,N_8476,N_8335);
or U8525 (N_8525,N_8324,N_8448);
or U8526 (N_8526,N_8273,N_8352);
or U8527 (N_8527,N_8420,N_8415);
or U8528 (N_8528,N_8319,N_8296);
and U8529 (N_8529,N_8439,N_8345);
and U8530 (N_8530,N_8289,N_8332);
or U8531 (N_8531,N_8431,N_8427);
nor U8532 (N_8532,N_8278,N_8495);
nor U8533 (N_8533,N_8414,N_8308);
nor U8534 (N_8534,N_8493,N_8337);
nand U8535 (N_8535,N_8387,N_8301);
nor U8536 (N_8536,N_8465,N_8349);
or U8537 (N_8537,N_8316,N_8376);
and U8538 (N_8538,N_8383,N_8492);
nor U8539 (N_8539,N_8295,N_8449);
or U8540 (N_8540,N_8292,N_8421);
or U8541 (N_8541,N_8348,N_8381);
nor U8542 (N_8542,N_8280,N_8432);
or U8543 (N_8543,N_8440,N_8470);
nor U8544 (N_8544,N_8329,N_8365);
or U8545 (N_8545,N_8355,N_8486);
nand U8546 (N_8546,N_8390,N_8371);
or U8547 (N_8547,N_8363,N_8311);
nand U8548 (N_8548,N_8272,N_8498);
or U8549 (N_8549,N_8310,N_8370);
nor U8550 (N_8550,N_8475,N_8453);
and U8551 (N_8551,N_8480,N_8451);
and U8552 (N_8552,N_8482,N_8454);
nand U8553 (N_8553,N_8455,N_8372);
or U8554 (N_8554,N_8357,N_8293);
nor U8555 (N_8555,N_8401,N_8360);
nand U8556 (N_8556,N_8422,N_8399);
and U8557 (N_8557,N_8256,N_8317);
or U8558 (N_8558,N_8291,N_8438);
and U8559 (N_8559,N_8460,N_8269);
or U8560 (N_8560,N_8327,N_8459);
and U8561 (N_8561,N_8443,N_8334);
or U8562 (N_8562,N_8340,N_8464);
and U8563 (N_8563,N_8343,N_8395);
nor U8564 (N_8564,N_8323,N_8382);
or U8565 (N_8565,N_8252,N_8391);
nor U8566 (N_8566,N_8347,N_8354);
nand U8567 (N_8567,N_8388,N_8413);
nor U8568 (N_8568,N_8419,N_8462);
or U8569 (N_8569,N_8458,N_8373);
nor U8570 (N_8570,N_8333,N_8457);
and U8571 (N_8571,N_8411,N_8375);
or U8572 (N_8572,N_8463,N_8369);
and U8573 (N_8573,N_8271,N_8418);
and U8574 (N_8574,N_8258,N_8367);
nand U8575 (N_8575,N_8409,N_8346);
nand U8576 (N_8576,N_8479,N_8270);
or U8577 (N_8577,N_8262,N_8275);
nor U8578 (N_8578,N_8468,N_8497);
nand U8579 (N_8579,N_8304,N_8485);
nand U8580 (N_8580,N_8408,N_8481);
nand U8581 (N_8581,N_8359,N_8339);
nor U8582 (N_8582,N_8499,N_8442);
xor U8583 (N_8583,N_8331,N_8313);
xnor U8584 (N_8584,N_8477,N_8287);
nand U8585 (N_8585,N_8315,N_8306);
or U8586 (N_8586,N_8342,N_8350);
nor U8587 (N_8587,N_8392,N_8263);
nand U8588 (N_8588,N_8466,N_8341);
nor U8589 (N_8589,N_8305,N_8378);
nor U8590 (N_8590,N_8456,N_8302);
or U8591 (N_8591,N_8377,N_8303);
and U8592 (N_8592,N_8405,N_8379);
nand U8593 (N_8593,N_8474,N_8403);
or U8594 (N_8594,N_8472,N_8307);
nand U8595 (N_8595,N_8297,N_8394);
and U8596 (N_8596,N_8282,N_8444);
nor U8597 (N_8597,N_8284,N_8445);
nor U8598 (N_8598,N_8380,N_8393);
or U8599 (N_8599,N_8368,N_8266);
and U8600 (N_8600,N_8361,N_8436);
nand U8601 (N_8601,N_8277,N_8362);
nand U8602 (N_8602,N_8264,N_8267);
or U8603 (N_8603,N_8326,N_8434);
or U8604 (N_8604,N_8353,N_8433);
and U8605 (N_8605,N_8450,N_8471);
and U8606 (N_8606,N_8255,N_8426);
and U8607 (N_8607,N_8491,N_8259);
nand U8608 (N_8608,N_8330,N_8406);
nand U8609 (N_8609,N_8257,N_8279);
nand U8610 (N_8610,N_8425,N_8400);
and U8611 (N_8611,N_8398,N_8430);
nor U8612 (N_8612,N_8385,N_8285);
or U8613 (N_8613,N_8260,N_8286);
nand U8614 (N_8614,N_8274,N_8309);
nor U8615 (N_8615,N_8299,N_8407);
or U8616 (N_8616,N_8452,N_8437);
and U8617 (N_8617,N_8366,N_8314);
nor U8618 (N_8618,N_8389,N_8265);
nor U8619 (N_8619,N_8461,N_8447);
or U8620 (N_8620,N_8288,N_8338);
nand U8621 (N_8621,N_8328,N_8488);
or U8622 (N_8622,N_8396,N_8467);
and U8623 (N_8623,N_8322,N_8351);
and U8624 (N_8624,N_8478,N_8374);
and U8625 (N_8625,N_8352,N_8305);
and U8626 (N_8626,N_8473,N_8480);
and U8627 (N_8627,N_8383,N_8345);
nand U8628 (N_8628,N_8257,N_8428);
nor U8629 (N_8629,N_8293,N_8498);
nand U8630 (N_8630,N_8432,N_8377);
and U8631 (N_8631,N_8467,N_8413);
nand U8632 (N_8632,N_8273,N_8434);
and U8633 (N_8633,N_8280,N_8452);
nand U8634 (N_8634,N_8330,N_8401);
nand U8635 (N_8635,N_8260,N_8433);
nand U8636 (N_8636,N_8423,N_8359);
nand U8637 (N_8637,N_8431,N_8477);
or U8638 (N_8638,N_8266,N_8414);
nand U8639 (N_8639,N_8482,N_8265);
or U8640 (N_8640,N_8269,N_8480);
or U8641 (N_8641,N_8439,N_8251);
nand U8642 (N_8642,N_8335,N_8327);
nor U8643 (N_8643,N_8263,N_8303);
and U8644 (N_8644,N_8271,N_8401);
or U8645 (N_8645,N_8470,N_8465);
and U8646 (N_8646,N_8459,N_8466);
and U8647 (N_8647,N_8254,N_8338);
or U8648 (N_8648,N_8254,N_8360);
nand U8649 (N_8649,N_8313,N_8464);
and U8650 (N_8650,N_8405,N_8371);
nor U8651 (N_8651,N_8274,N_8464);
nand U8652 (N_8652,N_8498,N_8318);
and U8653 (N_8653,N_8388,N_8255);
nand U8654 (N_8654,N_8495,N_8470);
nor U8655 (N_8655,N_8432,N_8489);
nor U8656 (N_8656,N_8254,N_8262);
or U8657 (N_8657,N_8285,N_8449);
nor U8658 (N_8658,N_8261,N_8370);
nor U8659 (N_8659,N_8412,N_8452);
nor U8660 (N_8660,N_8354,N_8461);
and U8661 (N_8661,N_8345,N_8385);
nor U8662 (N_8662,N_8322,N_8359);
and U8663 (N_8663,N_8297,N_8299);
and U8664 (N_8664,N_8351,N_8309);
nand U8665 (N_8665,N_8472,N_8499);
nand U8666 (N_8666,N_8369,N_8373);
or U8667 (N_8667,N_8348,N_8341);
nand U8668 (N_8668,N_8316,N_8373);
and U8669 (N_8669,N_8448,N_8342);
or U8670 (N_8670,N_8282,N_8261);
or U8671 (N_8671,N_8326,N_8491);
and U8672 (N_8672,N_8339,N_8348);
and U8673 (N_8673,N_8472,N_8308);
or U8674 (N_8674,N_8408,N_8452);
nor U8675 (N_8675,N_8339,N_8387);
and U8676 (N_8676,N_8301,N_8276);
nor U8677 (N_8677,N_8465,N_8479);
and U8678 (N_8678,N_8313,N_8429);
nand U8679 (N_8679,N_8385,N_8275);
or U8680 (N_8680,N_8321,N_8474);
nand U8681 (N_8681,N_8273,N_8442);
and U8682 (N_8682,N_8439,N_8265);
nor U8683 (N_8683,N_8362,N_8406);
or U8684 (N_8684,N_8343,N_8456);
nor U8685 (N_8685,N_8344,N_8251);
nand U8686 (N_8686,N_8340,N_8270);
nand U8687 (N_8687,N_8461,N_8266);
or U8688 (N_8688,N_8459,N_8474);
xor U8689 (N_8689,N_8287,N_8408);
nand U8690 (N_8690,N_8340,N_8415);
nor U8691 (N_8691,N_8339,N_8287);
and U8692 (N_8692,N_8396,N_8474);
nor U8693 (N_8693,N_8273,N_8451);
nand U8694 (N_8694,N_8258,N_8368);
and U8695 (N_8695,N_8493,N_8432);
and U8696 (N_8696,N_8445,N_8490);
or U8697 (N_8697,N_8307,N_8319);
or U8698 (N_8698,N_8393,N_8455);
nand U8699 (N_8699,N_8322,N_8424);
and U8700 (N_8700,N_8255,N_8300);
nand U8701 (N_8701,N_8289,N_8274);
and U8702 (N_8702,N_8327,N_8443);
and U8703 (N_8703,N_8381,N_8475);
nand U8704 (N_8704,N_8298,N_8349);
or U8705 (N_8705,N_8360,N_8397);
nand U8706 (N_8706,N_8389,N_8444);
and U8707 (N_8707,N_8413,N_8262);
nor U8708 (N_8708,N_8320,N_8315);
and U8709 (N_8709,N_8372,N_8496);
and U8710 (N_8710,N_8459,N_8321);
nor U8711 (N_8711,N_8318,N_8304);
or U8712 (N_8712,N_8250,N_8262);
and U8713 (N_8713,N_8483,N_8446);
nand U8714 (N_8714,N_8481,N_8452);
nor U8715 (N_8715,N_8484,N_8251);
nor U8716 (N_8716,N_8286,N_8414);
or U8717 (N_8717,N_8439,N_8281);
nor U8718 (N_8718,N_8443,N_8442);
or U8719 (N_8719,N_8288,N_8453);
or U8720 (N_8720,N_8382,N_8483);
or U8721 (N_8721,N_8369,N_8275);
nor U8722 (N_8722,N_8269,N_8441);
nand U8723 (N_8723,N_8270,N_8453);
nand U8724 (N_8724,N_8392,N_8428);
and U8725 (N_8725,N_8360,N_8474);
nor U8726 (N_8726,N_8354,N_8479);
and U8727 (N_8727,N_8476,N_8329);
or U8728 (N_8728,N_8343,N_8312);
and U8729 (N_8729,N_8399,N_8387);
and U8730 (N_8730,N_8484,N_8312);
nand U8731 (N_8731,N_8376,N_8394);
and U8732 (N_8732,N_8498,N_8322);
nor U8733 (N_8733,N_8477,N_8447);
nand U8734 (N_8734,N_8458,N_8268);
or U8735 (N_8735,N_8360,N_8368);
nor U8736 (N_8736,N_8294,N_8491);
or U8737 (N_8737,N_8341,N_8406);
and U8738 (N_8738,N_8382,N_8286);
nor U8739 (N_8739,N_8370,N_8324);
or U8740 (N_8740,N_8284,N_8431);
and U8741 (N_8741,N_8365,N_8392);
or U8742 (N_8742,N_8420,N_8448);
nand U8743 (N_8743,N_8425,N_8299);
nor U8744 (N_8744,N_8443,N_8488);
nor U8745 (N_8745,N_8489,N_8389);
nor U8746 (N_8746,N_8345,N_8498);
or U8747 (N_8747,N_8334,N_8277);
and U8748 (N_8748,N_8338,N_8392);
or U8749 (N_8749,N_8303,N_8477);
nor U8750 (N_8750,N_8541,N_8640);
nor U8751 (N_8751,N_8522,N_8543);
and U8752 (N_8752,N_8675,N_8501);
and U8753 (N_8753,N_8670,N_8612);
and U8754 (N_8754,N_8538,N_8738);
nand U8755 (N_8755,N_8588,N_8546);
nor U8756 (N_8756,N_8608,N_8733);
nor U8757 (N_8757,N_8651,N_8745);
and U8758 (N_8758,N_8658,N_8527);
nor U8759 (N_8759,N_8578,N_8652);
or U8760 (N_8760,N_8526,N_8564);
or U8761 (N_8761,N_8684,N_8679);
or U8762 (N_8762,N_8596,N_8532);
or U8763 (N_8763,N_8719,N_8537);
and U8764 (N_8764,N_8595,N_8562);
and U8765 (N_8765,N_8683,N_8568);
and U8766 (N_8766,N_8749,N_8587);
and U8767 (N_8767,N_8566,N_8731);
or U8768 (N_8768,N_8744,N_8603);
or U8769 (N_8769,N_8604,N_8613);
nor U8770 (N_8770,N_8539,N_8708);
or U8771 (N_8771,N_8669,N_8580);
and U8772 (N_8772,N_8736,N_8748);
and U8773 (N_8773,N_8556,N_8648);
nand U8774 (N_8774,N_8726,N_8552);
nand U8775 (N_8775,N_8691,N_8617);
nand U8776 (N_8776,N_8607,N_8703);
and U8777 (N_8777,N_8665,N_8505);
or U8778 (N_8778,N_8629,N_8545);
nand U8779 (N_8779,N_8506,N_8540);
and U8780 (N_8780,N_8746,N_8618);
nor U8781 (N_8781,N_8710,N_8517);
and U8782 (N_8782,N_8729,N_8686);
or U8783 (N_8783,N_8649,N_8525);
and U8784 (N_8784,N_8591,N_8689);
and U8785 (N_8785,N_8730,N_8645);
or U8786 (N_8786,N_8698,N_8633);
or U8787 (N_8787,N_8531,N_8561);
and U8788 (N_8788,N_8605,N_8668);
nand U8789 (N_8789,N_8586,N_8739);
nand U8790 (N_8790,N_8616,N_8671);
or U8791 (N_8791,N_8575,N_8567);
or U8792 (N_8792,N_8666,N_8519);
nand U8793 (N_8793,N_8592,N_8622);
and U8794 (N_8794,N_8542,N_8626);
or U8795 (N_8795,N_8523,N_8634);
or U8796 (N_8796,N_8712,N_8700);
and U8797 (N_8797,N_8643,N_8694);
and U8798 (N_8798,N_8535,N_8530);
nor U8799 (N_8799,N_8747,N_8641);
nor U8800 (N_8800,N_8687,N_8662);
and U8801 (N_8801,N_8601,N_8609);
nor U8802 (N_8802,N_8724,N_8685);
or U8803 (N_8803,N_8515,N_8695);
and U8804 (N_8804,N_8699,N_8598);
nor U8805 (N_8805,N_8620,N_8516);
nand U8806 (N_8806,N_8570,N_8565);
nor U8807 (N_8807,N_8690,N_8682);
nor U8808 (N_8808,N_8602,N_8674);
nand U8809 (N_8809,N_8741,N_8646);
nand U8810 (N_8810,N_8625,N_8637);
or U8811 (N_8811,N_8692,N_8705);
and U8812 (N_8812,N_8619,N_8585);
nand U8813 (N_8813,N_8707,N_8611);
nand U8814 (N_8814,N_8718,N_8632);
nor U8815 (N_8815,N_8696,N_8599);
nand U8816 (N_8816,N_8630,N_8732);
or U8817 (N_8817,N_8597,N_8569);
or U8818 (N_8818,N_8709,N_8704);
nand U8819 (N_8819,N_8742,N_8503);
or U8820 (N_8820,N_8717,N_8582);
or U8821 (N_8821,N_8560,N_8550);
nand U8822 (N_8822,N_8576,N_8688);
nand U8823 (N_8823,N_8728,N_8508);
and U8824 (N_8824,N_8635,N_8697);
nand U8825 (N_8825,N_8727,N_8593);
and U8826 (N_8826,N_8528,N_8715);
nand U8827 (N_8827,N_8614,N_8507);
nand U8828 (N_8828,N_8524,N_8638);
and U8829 (N_8829,N_8706,N_8521);
and U8830 (N_8830,N_8513,N_8702);
and U8831 (N_8831,N_8536,N_8714);
xor U8832 (N_8832,N_8577,N_8661);
nor U8833 (N_8833,N_8520,N_8636);
and U8834 (N_8834,N_8610,N_8627);
nand U8835 (N_8835,N_8594,N_8504);
and U8836 (N_8836,N_8500,N_8589);
and U8837 (N_8837,N_8659,N_8737);
nor U8838 (N_8838,N_8642,N_8555);
nor U8839 (N_8839,N_8548,N_8502);
nor U8840 (N_8840,N_8663,N_8529);
and U8841 (N_8841,N_8600,N_8650);
nor U8842 (N_8842,N_8557,N_8681);
nand U8843 (N_8843,N_8584,N_8680);
or U8844 (N_8844,N_8631,N_8701);
or U8845 (N_8845,N_8720,N_8558);
xor U8846 (N_8846,N_8572,N_8664);
nor U8847 (N_8847,N_8734,N_8721);
nor U8848 (N_8848,N_8660,N_8563);
or U8849 (N_8849,N_8624,N_8514);
nor U8850 (N_8850,N_8672,N_8615);
and U8851 (N_8851,N_8655,N_8647);
nor U8852 (N_8852,N_8544,N_8559);
and U8853 (N_8853,N_8667,N_8623);
nand U8854 (N_8854,N_8581,N_8628);
and U8855 (N_8855,N_8735,N_8654);
nand U8856 (N_8856,N_8740,N_8574);
nor U8857 (N_8857,N_8657,N_8579);
nand U8858 (N_8858,N_8554,N_8518);
nor U8859 (N_8859,N_8743,N_8606);
nand U8860 (N_8860,N_8673,N_8573);
nor U8861 (N_8861,N_8722,N_8725);
xor U8862 (N_8862,N_8571,N_8534);
or U8863 (N_8863,N_8509,N_8678);
nor U8864 (N_8864,N_8639,N_8512);
or U8865 (N_8865,N_8723,N_8676);
nor U8866 (N_8866,N_8533,N_8510);
nor U8867 (N_8867,N_8711,N_8716);
nor U8868 (N_8868,N_8511,N_8693);
or U8869 (N_8869,N_8656,N_8621);
nor U8870 (N_8870,N_8547,N_8583);
nand U8871 (N_8871,N_8677,N_8713);
nor U8872 (N_8872,N_8590,N_8549);
nor U8873 (N_8873,N_8644,N_8553);
nor U8874 (N_8874,N_8551,N_8653);
or U8875 (N_8875,N_8629,N_8546);
xnor U8876 (N_8876,N_8569,N_8589);
nand U8877 (N_8877,N_8586,N_8713);
and U8878 (N_8878,N_8532,N_8702);
and U8879 (N_8879,N_8507,N_8652);
or U8880 (N_8880,N_8524,N_8666);
or U8881 (N_8881,N_8564,N_8561);
nor U8882 (N_8882,N_8505,N_8515);
and U8883 (N_8883,N_8576,N_8510);
nand U8884 (N_8884,N_8668,N_8742);
and U8885 (N_8885,N_8667,N_8601);
and U8886 (N_8886,N_8604,N_8558);
and U8887 (N_8887,N_8656,N_8650);
and U8888 (N_8888,N_8527,N_8744);
nor U8889 (N_8889,N_8522,N_8529);
or U8890 (N_8890,N_8722,N_8508);
or U8891 (N_8891,N_8722,N_8606);
nand U8892 (N_8892,N_8739,N_8531);
and U8893 (N_8893,N_8623,N_8521);
and U8894 (N_8894,N_8707,N_8742);
or U8895 (N_8895,N_8645,N_8509);
nand U8896 (N_8896,N_8568,N_8523);
nand U8897 (N_8897,N_8532,N_8565);
or U8898 (N_8898,N_8560,N_8534);
nor U8899 (N_8899,N_8626,N_8500);
or U8900 (N_8900,N_8564,N_8705);
and U8901 (N_8901,N_8524,N_8535);
and U8902 (N_8902,N_8569,N_8727);
or U8903 (N_8903,N_8548,N_8681);
and U8904 (N_8904,N_8533,N_8562);
nand U8905 (N_8905,N_8568,N_8591);
and U8906 (N_8906,N_8600,N_8727);
and U8907 (N_8907,N_8547,N_8654);
or U8908 (N_8908,N_8741,N_8658);
and U8909 (N_8909,N_8534,N_8556);
nand U8910 (N_8910,N_8509,N_8677);
nand U8911 (N_8911,N_8646,N_8723);
and U8912 (N_8912,N_8640,N_8628);
or U8913 (N_8913,N_8555,N_8745);
nand U8914 (N_8914,N_8680,N_8608);
nand U8915 (N_8915,N_8620,N_8651);
or U8916 (N_8916,N_8675,N_8747);
nand U8917 (N_8917,N_8674,N_8673);
nor U8918 (N_8918,N_8661,N_8649);
nor U8919 (N_8919,N_8656,N_8520);
nand U8920 (N_8920,N_8657,N_8610);
or U8921 (N_8921,N_8673,N_8534);
nand U8922 (N_8922,N_8748,N_8508);
or U8923 (N_8923,N_8724,N_8630);
and U8924 (N_8924,N_8508,N_8545);
nand U8925 (N_8925,N_8740,N_8691);
or U8926 (N_8926,N_8580,N_8611);
xor U8927 (N_8927,N_8599,N_8569);
or U8928 (N_8928,N_8520,N_8525);
nand U8929 (N_8929,N_8747,N_8698);
and U8930 (N_8930,N_8726,N_8542);
or U8931 (N_8931,N_8697,N_8740);
nand U8932 (N_8932,N_8682,N_8620);
nand U8933 (N_8933,N_8749,N_8721);
and U8934 (N_8934,N_8711,N_8591);
or U8935 (N_8935,N_8537,N_8714);
xnor U8936 (N_8936,N_8641,N_8617);
nor U8937 (N_8937,N_8507,N_8597);
or U8938 (N_8938,N_8510,N_8679);
and U8939 (N_8939,N_8638,N_8702);
nand U8940 (N_8940,N_8600,N_8678);
and U8941 (N_8941,N_8547,N_8541);
xnor U8942 (N_8942,N_8608,N_8704);
nand U8943 (N_8943,N_8667,N_8556);
nor U8944 (N_8944,N_8575,N_8643);
nand U8945 (N_8945,N_8746,N_8572);
nand U8946 (N_8946,N_8524,N_8655);
nand U8947 (N_8947,N_8549,N_8646);
or U8948 (N_8948,N_8728,N_8622);
nand U8949 (N_8949,N_8628,N_8501);
xnor U8950 (N_8950,N_8696,N_8529);
nand U8951 (N_8951,N_8625,N_8600);
nor U8952 (N_8952,N_8614,N_8709);
and U8953 (N_8953,N_8677,N_8581);
nor U8954 (N_8954,N_8644,N_8523);
nand U8955 (N_8955,N_8632,N_8682);
or U8956 (N_8956,N_8691,N_8728);
and U8957 (N_8957,N_8677,N_8604);
or U8958 (N_8958,N_8746,N_8716);
and U8959 (N_8959,N_8646,N_8511);
or U8960 (N_8960,N_8748,N_8634);
and U8961 (N_8961,N_8731,N_8546);
nand U8962 (N_8962,N_8747,N_8741);
nor U8963 (N_8963,N_8733,N_8645);
or U8964 (N_8964,N_8537,N_8502);
nor U8965 (N_8965,N_8613,N_8618);
and U8966 (N_8966,N_8500,N_8631);
nand U8967 (N_8967,N_8662,N_8713);
or U8968 (N_8968,N_8543,N_8678);
nand U8969 (N_8969,N_8700,N_8630);
nor U8970 (N_8970,N_8519,N_8650);
or U8971 (N_8971,N_8662,N_8621);
nor U8972 (N_8972,N_8580,N_8506);
nand U8973 (N_8973,N_8557,N_8636);
or U8974 (N_8974,N_8651,N_8536);
nor U8975 (N_8975,N_8539,N_8563);
or U8976 (N_8976,N_8533,N_8550);
or U8977 (N_8977,N_8544,N_8716);
nand U8978 (N_8978,N_8519,N_8641);
or U8979 (N_8979,N_8529,N_8538);
or U8980 (N_8980,N_8519,N_8703);
xnor U8981 (N_8981,N_8702,N_8650);
or U8982 (N_8982,N_8620,N_8622);
nand U8983 (N_8983,N_8559,N_8578);
or U8984 (N_8984,N_8671,N_8682);
and U8985 (N_8985,N_8566,N_8544);
or U8986 (N_8986,N_8724,N_8687);
or U8987 (N_8987,N_8736,N_8515);
or U8988 (N_8988,N_8665,N_8547);
nor U8989 (N_8989,N_8726,N_8504);
or U8990 (N_8990,N_8669,N_8683);
nor U8991 (N_8991,N_8628,N_8621);
and U8992 (N_8992,N_8556,N_8660);
nor U8993 (N_8993,N_8715,N_8722);
xor U8994 (N_8994,N_8646,N_8607);
xnor U8995 (N_8995,N_8591,N_8708);
nand U8996 (N_8996,N_8509,N_8724);
nand U8997 (N_8997,N_8557,N_8714);
and U8998 (N_8998,N_8715,N_8537);
or U8999 (N_8999,N_8644,N_8682);
nor U9000 (N_9000,N_8967,N_8962);
nor U9001 (N_9001,N_8880,N_8765);
nand U9002 (N_9002,N_8862,N_8943);
or U9003 (N_9003,N_8755,N_8953);
or U9004 (N_9004,N_8936,N_8822);
nor U9005 (N_9005,N_8792,N_8828);
nor U9006 (N_9006,N_8964,N_8754);
nor U9007 (N_9007,N_8857,N_8836);
and U9008 (N_9008,N_8850,N_8753);
nor U9009 (N_9009,N_8934,N_8948);
or U9010 (N_9010,N_8994,N_8979);
or U9011 (N_9011,N_8832,N_8767);
and U9012 (N_9012,N_8879,N_8838);
nor U9013 (N_9013,N_8801,N_8788);
nor U9014 (N_9014,N_8961,N_8963);
or U9015 (N_9015,N_8995,N_8893);
nor U9016 (N_9016,N_8906,N_8927);
or U9017 (N_9017,N_8797,N_8899);
or U9018 (N_9018,N_8888,N_8777);
nor U9019 (N_9019,N_8892,N_8835);
nor U9020 (N_9020,N_8972,N_8853);
nor U9021 (N_9021,N_8837,N_8989);
or U9022 (N_9022,N_8846,N_8965);
and U9023 (N_9023,N_8816,N_8773);
nand U9024 (N_9024,N_8900,N_8954);
and U9025 (N_9025,N_8809,N_8774);
xor U9026 (N_9026,N_8870,N_8891);
nor U9027 (N_9027,N_8912,N_8895);
or U9028 (N_9028,N_8819,N_8908);
or U9029 (N_9029,N_8883,N_8750);
and U9030 (N_9030,N_8821,N_8863);
nand U9031 (N_9031,N_8849,N_8919);
nand U9032 (N_9032,N_8826,N_8763);
nand U9033 (N_9033,N_8882,N_8806);
and U9034 (N_9034,N_8905,N_8983);
and U9035 (N_9035,N_8896,N_8988);
nand U9036 (N_9036,N_8876,N_8847);
or U9037 (N_9037,N_8901,N_8966);
nand U9038 (N_9038,N_8910,N_8907);
xnor U9039 (N_9039,N_8769,N_8981);
nand U9040 (N_9040,N_8851,N_8920);
nor U9041 (N_9041,N_8782,N_8868);
or U9042 (N_9042,N_8808,N_8968);
xor U9043 (N_9043,N_8783,N_8772);
and U9044 (N_9044,N_8815,N_8974);
and U9045 (N_9045,N_8798,N_8766);
or U9046 (N_9046,N_8976,N_8844);
and U9047 (N_9047,N_8940,N_8776);
nor U9048 (N_9048,N_8894,N_8759);
nor U9049 (N_9049,N_8793,N_8761);
or U9050 (N_9050,N_8771,N_8827);
and U9051 (N_9051,N_8830,N_8993);
nand U9052 (N_9052,N_8984,N_8947);
and U9053 (N_9053,N_8817,N_8818);
nand U9054 (N_9054,N_8887,N_8824);
nand U9055 (N_9055,N_8952,N_8939);
and U9056 (N_9056,N_8871,N_8904);
nand U9057 (N_9057,N_8790,N_8752);
nor U9058 (N_9058,N_8855,N_8758);
nor U9059 (N_9059,N_8834,N_8903);
nor U9060 (N_9060,N_8987,N_8926);
and U9061 (N_9061,N_8878,N_8959);
nor U9062 (N_9062,N_8866,N_8794);
nor U9063 (N_9063,N_8820,N_8751);
and U9064 (N_9064,N_8889,N_8779);
and U9065 (N_9065,N_8760,N_8898);
nor U9066 (N_9066,N_8781,N_8829);
and U9067 (N_9067,N_8881,N_8823);
nor U9068 (N_9068,N_8999,N_8950);
and U9069 (N_9069,N_8922,N_8825);
nand U9070 (N_9070,N_8803,N_8897);
nor U9071 (N_9071,N_8840,N_8977);
or U9072 (N_9072,N_8852,N_8884);
nor U9073 (N_9073,N_8872,N_8924);
nand U9074 (N_9074,N_8998,N_8789);
or U9075 (N_9075,N_8831,N_8944);
or U9076 (N_9076,N_8784,N_8929);
and U9077 (N_9077,N_8869,N_8909);
nor U9078 (N_9078,N_8973,N_8970);
or U9079 (N_9079,N_8957,N_8860);
and U9080 (N_9080,N_8842,N_8938);
nor U9081 (N_9081,N_8902,N_8833);
nand U9082 (N_9082,N_8982,N_8786);
nand U9083 (N_9083,N_8800,N_8854);
nor U9084 (N_9084,N_8757,N_8810);
or U9085 (N_9085,N_8756,N_8875);
and U9086 (N_9086,N_8978,N_8796);
nand U9087 (N_9087,N_8787,N_8941);
or U9088 (N_9088,N_8861,N_8937);
or U9089 (N_9089,N_8848,N_8942);
nand U9090 (N_9090,N_8935,N_8864);
and U9091 (N_9091,N_8958,N_8932);
nor U9092 (N_9092,N_8992,N_8811);
nor U9093 (N_9093,N_8807,N_8991);
or U9094 (N_9094,N_8928,N_8770);
nor U9095 (N_9095,N_8949,N_8839);
or U9096 (N_9096,N_8980,N_8877);
and U9097 (N_9097,N_8996,N_8985);
or U9098 (N_9098,N_8799,N_8914);
or U9099 (N_9099,N_8841,N_8867);
and U9100 (N_9100,N_8780,N_8802);
nand U9101 (N_9101,N_8960,N_8921);
nor U9102 (N_9102,N_8762,N_8930);
or U9103 (N_9103,N_8915,N_8886);
nor U9104 (N_9104,N_8843,N_8946);
or U9105 (N_9105,N_8791,N_8885);
nor U9106 (N_9106,N_8805,N_8874);
nand U9107 (N_9107,N_8858,N_8918);
or U9108 (N_9108,N_8986,N_8911);
nand U9109 (N_9109,N_8925,N_8951);
nand U9110 (N_9110,N_8990,N_8804);
or U9111 (N_9111,N_8916,N_8814);
nor U9112 (N_9112,N_8971,N_8795);
or U9113 (N_9113,N_8813,N_8923);
or U9114 (N_9114,N_8785,N_8873);
and U9115 (N_9115,N_8975,N_8945);
nor U9116 (N_9116,N_8933,N_8768);
or U9117 (N_9117,N_8955,N_8917);
nand U9118 (N_9118,N_8812,N_8775);
nor U9119 (N_9119,N_8969,N_8856);
nor U9120 (N_9120,N_8997,N_8778);
and U9121 (N_9121,N_8956,N_8865);
or U9122 (N_9122,N_8764,N_8913);
or U9123 (N_9123,N_8845,N_8859);
or U9124 (N_9124,N_8931,N_8890);
nand U9125 (N_9125,N_8908,N_8973);
or U9126 (N_9126,N_8939,N_8915);
or U9127 (N_9127,N_8978,N_8901);
or U9128 (N_9128,N_8768,N_8803);
or U9129 (N_9129,N_8807,N_8889);
nor U9130 (N_9130,N_8842,N_8916);
nor U9131 (N_9131,N_8920,N_8966);
nand U9132 (N_9132,N_8882,N_8763);
nand U9133 (N_9133,N_8865,N_8883);
and U9134 (N_9134,N_8905,N_8751);
and U9135 (N_9135,N_8892,N_8807);
and U9136 (N_9136,N_8839,N_8934);
and U9137 (N_9137,N_8942,N_8842);
nor U9138 (N_9138,N_8901,N_8907);
and U9139 (N_9139,N_8965,N_8924);
nor U9140 (N_9140,N_8765,N_8774);
nand U9141 (N_9141,N_8774,N_8811);
nor U9142 (N_9142,N_8861,N_8978);
nor U9143 (N_9143,N_8844,N_8818);
nor U9144 (N_9144,N_8864,N_8915);
nand U9145 (N_9145,N_8797,N_8926);
or U9146 (N_9146,N_8975,N_8809);
or U9147 (N_9147,N_8803,N_8766);
nand U9148 (N_9148,N_8775,N_8867);
and U9149 (N_9149,N_8844,N_8796);
and U9150 (N_9150,N_8974,N_8978);
or U9151 (N_9151,N_8977,N_8812);
nand U9152 (N_9152,N_8899,N_8820);
nor U9153 (N_9153,N_8998,N_8996);
nand U9154 (N_9154,N_8867,N_8998);
nor U9155 (N_9155,N_8959,N_8946);
nor U9156 (N_9156,N_8912,N_8866);
nor U9157 (N_9157,N_8964,N_8973);
or U9158 (N_9158,N_8781,N_8964);
nand U9159 (N_9159,N_8856,N_8896);
and U9160 (N_9160,N_8820,N_8765);
and U9161 (N_9161,N_8855,N_8933);
and U9162 (N_9162,N_8930,N_8936);
nand U9163 (N_9163,N_8933,N_8970);
or U9164 (N_9164,N_8964,N_8808);
and U9165 (N_9165,N_8827,N_8782);
or U9166 (N_9166,N_8757,N_8775);
and U9167 (N_9167,N_8868,N_8806);
or U9168 (N_9168,N_8863,N_8909);
nor U9169 (N_9169,N_8792,N_8812);
nor U9170 (N_9170,N_8853,N_8830);
nor U9171 (N_9171,N_8851,N_8865);
nand U9172 (N_9172,N_8928,N_8788);
and U9173 (N_9173,N_8785,N_8934);
or U9174 (N_9174,N_8887,N_8872);
or U9175 (N_9175,N_8969,N_8834);
nand U9176 (N_9176,N_8988,N_8915);
nand U9177 (N_9177,N_8797,N_8967);
nor U9178 (N_9178,N_8768,N_8807);
and U9179 (N_9179,N_8995,N_8856);
and U9180 (N_9180,N_8991,N_8823);
and U9181 (N_9181,N_8867,N_8799);
nor U9182 (N_9182,N_8889,N_8966);
nor U9183 (N_9183,N_8924,N_8919);
and U9184 (N_9184,N_8844,N_8927);
and U9185 (N_9185,N_8984,N_8959);
nand U9186 (N_9186,N_8910,N_8881);
nand U9187 (N_9187,N_8774,N_8913);
or U9188 (N_9188,N_8836,N_8819);
nor U9189 (N_9189,N_8774,N_8950);
or U9190 (N_9190,N_8870,N_8872);
nor U9191 (N_9191,N_8980,N_8842);
or U9192 (N_9192,N_8794,N_8950);
nand U9193 (N_9193,N_8759,N_8828);
or U9194 (N_9194,N_8858,N_8975);
nor U9195 (N_9195,N_8988,N_8861);
xnor U9196 (N_9196,N_8899,N_8900);
or U9197 (N_9197,N_8851,N_8757);
and U9198 (N_9198,N_8882,N_8886);
or U9199 (N_9199,N_8986,N_8856);
or U9200 (N_9200,N_8819,N_8820);
or U9201 (N_9201,N_8806,N_8939);
nand U9202 (N_9202,N_8914,N_8845);
or U9203 (N_9203,N_8829,N_8815);
nand U9204 (N_9204,N_8884,N_8758);
or U9205 (N_9205,N_8990,N_8956);
or U9206 (N_9206,N_8947,N_8982);
and U9207 (N_9207,N_8763,N_8956);
nor U9208 (N_9208,N_8900,N_8975);
or U9209 (N_9209,N_8999,N_8987);
nand U9210 (N_9210,N_8780,N_8763);
and U9211 (N_9211,N_8882,N_8762);
nand U9212 (N_9212,N_8958,N_8842);
nor U9213 (N_9213,N_8814,N_8879);
nor U9214 (N_9214,N_8891,N_8776);
nand U9215 (N_9215,N_8832,N_8966);
or U9216 (N_9216,N_8800,N_8809);
and U9217 (N_9217,N_8852,N_8828);
and U9218 (N_9218,N_8893,N_8767);
and U9219 (N_9219,N_8978,N_8986);
and U9220 (N_9220,N_8936,N_8855);
nand U9221 (N_9221,N_8951,N_8853);
nor U9222 (N_9222,N_8890,N_8785);
and U9223 (N_9223,N_8868,N_8893);
and U9224 (N_9224,N_8786,N_8855);
and U9225 (N_9225,N_8960,N_8757);
xnor U9226 (N_9226,N_8934,N_8756);
nand U9227 (N_9227,N_8953,N_8979);
and U9228 (N_9228,N_8905,N_8857);
or U9229 (N_9229,N_8978,N_8964);
nor U9230 (N_9230,N_8756,N_8793);
and U9231 (N_9231,N_8824,N_8855);
nor U9232 (N_9232,N_8854,N_8912);
or U9233 (N_9233,N_8921,N_8840);
nor U9234 (N_9234,N_8760,N_8921);
nand U9235 (N_9235,N_8862,N_8790);
nor U9236 (N_9236,N_8854,N_8929);
or U9237 (N_9237,N_8781,N_8914);
nand U9238 (N_9238,N_8770,N_8863);
nor U9239 (N_9239,N_8784,N_8933);
and U9240 (N_9240,N_8935,N_8896);
and U9241 (N_9241,N_8792,N_8880);
nor U9242 (N_9242,N_8787,N_8971);
or U9243 (N_9243,N_8819,N_8862);
or U9244 (N_9244,N_8847,N_8998);
or U9245 (N_9245,N_8884,N_8763);
or U9246 (N_9246,N_8838,N_8949);
nor U9247 (N_9247,N_8926,N_8856);
nor U9248 (N_9248,N_8770,N_8979);
nor U9249 (N_9249,N_8964,N_8986);
and U9250 (N_9250,N_9014,N_9212);
and U9251 (N_9251,N_9102,N_9146);
nor U9252 (N_9252,N_9003,N_9184);
and U9253 (N_9253,N_9164,N_9093);
nor U9254 (N_9254,N_9183,N_9158);
xnor U9255 (N_9255,N_9217,N_9225);
nor U9256 (N_9256,N_9203,N_9037);
nand U9257 (N_9257,N_9244,N_9055);
nor U9258 (N_9258,N_9230,N_9169);
nand U9259 (N_9259,N_9043,N_9181);
or U9260 (N_9260,N_9130,N_9009);
nor U9261 (N_9261,N_9126,N_9010);
nor U9262 (N_9262,N_9232,N_9088);
nand U9263 (N_9263,N_9028,N_9165);
and U9264 (N_9264,N_9054,N_9188);
or U9265 (N_9265,N_9019,N_9198);
and U9266 (N_9266,N_9153,N_9180);
nor U9267 (N_9267,N_9100,N_9117);
or U9268 (N_9268,N_9066,N_9096);
and U9269 (N_9269,N_9053,N_9175);
nor U9270 (N_9270,N_9029,N_9012);
and U9271 (N_9271,N_9024,N_9087);
or U9272 (N_9272,N_9199,N_9155);
or U9273 (N_9273,N_9196,N_9177);
and U9274 (N_9274,N_9119,N_9125);
or U9275 (N_9275,N_9056,N_9101);
or U9276 (N_9276,N_9033,N_9161);
nor U9277 (N_9277,N_9190,N_9006);
or U9278 (N_9278,N_9071,N_9157);
and U9279 (N_9279,N_9191,N_9209);
nor U9280 (N_9280,N_9240,N_9204);
nor U9281 (N_9281,N_9160,N_9152);
nor U9282 (N_9282,N_9243,N_9247);
nor U9283 (N_9283,N_9151,N_9085);
nor U9284 (N_9284,N_9064,N_9110);
or U9285 (N_9285,N_9229,N_9038);
or U9286 (N_9286,N_9048,N_9142);
nand U9287 (N_9287,N_9002,N_9045);
and U9288 (N_9288,N_9178,N_9156);
and U9289 (N_9289,N_9228,N_9201);
and U9290 (N_9290,N_9219,N_9026);
nor U9291 (N_9291,N_9216,N_9001);
or U9292 (N_9292,N_9246,N_9097);
or U9293 (N_9293,N_9074,N_9089);
nand U9294 (N_9294,N_9124,N_9020);
or U9295 (N_9295,N_9154,N_9103);
and U9296 (N_9296,N_9138,N_9150);
or U9297 (N_9297,N_9215,N_9098);
nor U9298 (N_9298,N_9176,N_9236);
nor U9299 (N_9299,N_9017,N_9116);
or U9300 (N_9300,N_9141,N_9106);
and U9301 (N_9301,N_9172,N_9113);
or U9302 (N_9302,N_9131,N_9245);
nand U9303 (N_9303,N_9075,N_9070);
or U9304 (N_9304,N_9221,N_9210);
nor U9305 (N_9305,N_9111,N_9086);
nor U9306 (N_9306,N_9135,N_9025);
nor U9307 (N_9307,N_9227,N_9092);
or U9308 (N_9308,N_9051,N_9162);
and U9309 (N_9309,N_9249,N_9171);
nor U9310 (N_9310,N_9222,N_9005);
nand U9311 (N_9311,N_9076,N_9032);
nor U9312 (N_9312,N_9039,N_9205);
or U9313 (N_9313,N_9238,N_9062);
and U9314 (N_9314,N_9174,N_9213);
nor U9315 (N_9315,N_9067,N_9140);
nor U9316 (N_9316,N_9139,N_9134);
nand U9317 (N_9317,N_9036,N_9011);
or U9318 (N_9318,N_9211,N_9136);
and U9319 (N_9319,N_9104,N_9073);
and U9320 (N_9320,N_9046,N_9034);
nand U9321 (N_9321,N_9168,N_9091);
xor U9322 (N_9322,N_9173,N_9042);
or U9323 (N_9323,N_9109,N_9059);
nor U9324 (N_9324,N_9061,N_9200);
and U9325 (N_9325,N_9082,N_9069);
and U9326 (N_9326,N_9159,N_9118);
nand U9327 (N_9327,N_9233,N_9187);
and U9328 (N_9328,N_9099,N_9008);
nor U9329 (N_9329,N_9120,N_9015);
nor U9330 (N_9330,N_9114,N_9193);
nand U9331 (N_9331,N_9084,N_9237);
nor U9332 (N_9332,N_9148,N_9145);
and U9333 (N_9333,N_9133,N_9195);
nand U9334 (N_9334,N_9049,N_9128);
or U9335 (N_9335,N_9027,N_9081);
and U9336 (N_9336,N_9202,N_9063);
or U9337 (N_9337,N_9021,N_9018);
nor U9338 (N_9338,N_9224,N_9000);
or U9339 (N_9339,N_9013,N_9189);
nor U9340 (N_9340,N_9107,N_9129);
or U9341 (N_9341,N_9065,N_9223);
xor U9342 (N_9342,N_9231,N_9090);
and U9343 (N_9343,N_9208,N_9239);
or U9344 (N_9344,N_9248,N_9016);
nand U9345 (N_9345,N_9127,N_9207);
nor U9346 (N_9346,N_9078,N_9047);
and U9347 (N_9347,N_9242,N_9052);
nor U9348 (N_9348,N_9058,N_9004);
or U9349 (N_9349,N_9115,N_9234);
and U9350 (N_9350,N_9241,N_9040);
nor U9351 (N_9351,N_9060,N_9022);
nor U9352 (N_9352,N_9192,N_9112);
nand U9353 (N_9353,N_9094,N_9057);
nand U9354 (N_9354,N_9144,N_9031);
nand U9355 (N_9355,N_9149,N_9105);
nand U9356 (N_9356,N_9179,N_9220);
nand U9357 (N_9357,N_9123,N_9077);
xnor U9358 (N_9358,N_9182,N_9137);
nor U9359 (N_9359,N_9122,N_9166);
and U9360 (N_9360,N_9170,N_9030);
or U9361 (N_9361,N_9121,N_9235);
nor U9362 (N_9362,N_9143,N_9035);
nand U9363 (N_9363,N_9214,N_9068);
or U9364 (N_9364,N_9007,N_9072);
or U9365 (N_9365,N_9041,N_9147);
nand U9366 (N_9366,N_9095,N_9197);
and U9367 (N_9367,N_9083,N_9079);
and U9368 (N_9368,N_9080,N_9194);
or U9369 (N_9369,N_9186,N_9050);
or U9370 (N_9370,N_9167,N_9226);
nand U9371 (N_9371,N_9218,N_9163);
nor U9372 (N_9372,N_9044,N_9206);
nor U9373 (N_9373,N_9132,N_9108);
nand U9374 (N_9374,N_9185,N_9023);
or U9375 (N_9375,N_9027,N_9199);
nand U9376 (N_9376,N_9152,N_9213);
and U9377 (N_9377,N_9045,N_9140);
and U9378 (N_9378,N_9174,N_9240);
nand U9379 (N_9379,N_9160,N_9031);
or U9380 (N_9380,N_9019,N_9193);
nor U9381 (N_9381,N_9234,N_9135);
nand U9382 (N_9382,N_9162,N_9074);
nor U9383 (N_9383,N_9074,N_9001);
nand U9384 (N_9384,N_9234,N_9095);
nor U9385 (N_9385,N_9035,N_9090);
and U9386 (N_9386,N_9249,N_9147);
nand U9387 (N_9387,N_9047,N_9208);
nand U9388 (N_9388,N_9205,N_9011);
nor U9389 (N_9389,N_9137,N_9248);
nor U9390 (N_9390,N_9176,N_9048);
and U9391 (N_9391,N_9181,N_9136);
nand U9392 (N_9392,N_9129,N_9239);
nor U9393 (N_9393,N_9110,N_9042);
and U9394 (N_9394,N_9211,N_9134);
nor U9395 (N_9395,N_9004,N_9237);
nor U9396 (N_9396,N_9120,N_9130);
and U9397 (N_9397,N_9212,N_9038);
and U9398 (N_9398,N_9094,N_9190);
nor U9399 (N_9399,N_9218,N_9024);
nand U9400 (N_9400,N_9142,N_9123);
and U9401 (N_9401,N_9206,N_9082);
nand U9402 (N_9402,N_9099,N_9209);
or U9403 (N_9403,N_9003,N_9120);
or U9404 (N_9404,N_9199,N_9039);
nand U9405 (N_9405,N_9189,N_9009);
and U9406 (N_9406,N_9099,N_9204);
and U9407 (N_9407,N_9246,N_9184);
nand U9408 (N_9408,N_9078,N_9145);
nor U9409 (N_9409,N_9167,N_9066);
nor U9410 (N_9410,N_9053,N_9120);
and U9411 (N_9411,N_9238,N_9206);
and U9412 (N_9412,N_9180,N_9241);
or U9413 (N_9413,N_9220,N_9134);
or U9414 (N_9414,N_9217,N_9014);
and U9415 (N_9415,N_9056,N_9029);
and U9416 (N_9416,N_9206,N_9133);
or U9417 (N_9417,N_9001,N_9142);
or U9418 (N_9418,N_9217,N_9119);
and U9419 (N_9419,N_9178,N_9059);
nor U9420 (N_9420,N_9075,N_9137);
nor U9421 (N_9421,N_9013,N_9057);
and U9422 (N_9422,N_9247,N_9093);
or U9423 (N_9423,N_9131,N_9011);
nand U9424 (N_9424,N_9121,N_9056);
nor U9425 (N_9425,N_9158,N_9216);
nand U9426 (N_9426,N_9200,N_9047);
nor U9427 (N_9427,N_9096,N_9215);
or U9428 (N_9428,N_9143,N_9163);
or U9429 (N_9429,N_9066,N_9174);
nor U9430 (N_9430,N_9060,N_9040);
and U9431 (N_9431,N_9104,N_9111);
and U9432 (N_9432,N_9161,N_9113);
or U9433 (N_9433,N_9120,N_9001);
nor U9434 (N_9434,N_9130,N_9053);
or U9435 (N_9435,N_9138,N_9113);
nor U9436 (N_9436,N_9014,N_9194);
and U9437 (N_9437,N_9168,N_9046);
nand U9438 (N_9438,N_9123,N_9032);
nand U9439 (N_9439,N_9222,N_9244);
nor U9440 (N_9440,N_9093,N_9249);
xor U9441 (N_9441,N_9024,N_9164);
xor U9442 (N_9442,N_9103,N_9041);
nor U9443 (N_9443,N_9069,N_9215);
nand U9444 (N_9444,N_9027,N_9188);
and U9445 (N_9445,N_9027,N_9212);
nor U9446 (N_9446,N_9193,N_9215);
or U9447 (N_9447,N_9048,N_9173);
and U9448 (N_9448,N_9005,N_9113);
nand U9449 (N_9449,N_9077,N_9089);
nand U9450 (N_9450,N_9033,N_9149);
nand U9451 (N_9451,N_9103,N_9204);
nor U9452 (N_9452,N_9089,N_9075);
nor U9453 (N_9453,N_9001,N_9143);
nor U9454 (N_9454,N_9069,N_9077);
nor U9455 (N_9455,N_9197,N_9153);
nor U9456 (N_9456,N_9025,N_9120);
and U9457 (N_9457,N_9134,N_9239);
or U9458 (N_9458,N_9029,N_9024);
nor U9459 (N_9459,N_9068,N_9054);
nor U9460 (N_9460,N_9145,N_9016);
or U9461 (N_9461,N_9227,N_9149);
nor U9462 (N_9462,N_9001,N_9047);
or U9463 (N_9463,N_9155,N_9084);
and U9464 (N_9464,N_9016,N_9046);
xnor U9465 (N_9465,N_9035,N_9071);
nand U9466 (N_9466,N_9214,N_9218);
and U9467 (N_9467,N_9244,N_9123);
or U9468 (N_9468,N_9187,N_9072);
nand U9469 (N_9469,N_9178,N_9150);
and U9470 (N_9470,N_9150,N_9249);
nor U9471 (N_9471,N_9124,N_9045);
nor U9472 (N_9472,N_9227,N_9072);
or U9473 (N_9473,N_9072,N_9082);
nor U9474 (N_9474,N_9015,N_9105);
nand U9475 (N_9475,N_9240,N_9209);
or U9476 (N_9476,N_9076,N_9185);
or U9477 (N_9477,N_9028,N_9145);
or U9478 (N_9478,N_9195,N_9015);
or U9479 (N_9479,N_9205,N_9076);
nor U9480 (N_9480,N_9095,N_9238);
nor U9481 (N_9481,N_9161,N_9003);
nor U9482 (N_9482,N_9227,N_9055);
nor U9483 (N_9483,N_9234,N_9195);
or U9484 (N_9484,N_9165,N_9214);
or U9485 (N_9485,N_9227,N_9148);
and U9486 (N_9486,N_9239,N_9041);
xor U9487 (N_9487,N_9069,N_9179);
and U9488 (N_9488,N_9101,N_9020);
or U9489 (N_9489,N_9126,N_9033);
nor U9490 (N_9490,N_9204,N_9066);
or U9491 (N_9491,N_9086,N_9249);
and U9492 (N_9492,N_9079,N_9013);
or U9493 (N_9493,N_9230,N_9049);
nor U9494 (N_9494,N_9182,N_9018);
and U9495 (N_9495,N_9031,N_9119);
and U9496 (N_9496,N_9143,N_9140);
nand U9497 (N_9497,N_9175,N_9084);
or U9498 (N_9498,N_9211,N_9000);
and U9499 (N_9499,N_9152,N_9165);
nand U9500 (N_9500,N_9279,N_9403);
and U9501 (N_9501,N_9309,N_9344);
or U9502 (N_9502,N_9289,N_9383);
nand U9503 (N_9503,N_9276,N_9400);
or U9504 (N_9504,N_9469,N_9385);
or U9505 (N_9505,N_9356,N_9430);
nand U9506 (N_9506,N_9277,N_9267);
or U9507 (N_9507,N_9419,N_9411);
nand U9508 (N_9508,N_9278,N_9372);
and U9509 (N_9509,N_9432,N_9451);
and U9510 (N_9510,N_9358,N_9449);
or U9511 (N_9511,N_9284,N_9417);
nor U9512 (N_9512,N_9465,N_9416);
and U9513 (N_9513,N_9326,N_9260);
nor U9514 (N_9514,N_9397,N_9257);
and U9515 (N_9515,N_9497,N_9299);
and U9516 (N_9516,N_9334,N_9335);
and U9517 (N_9517,N_9450,N_9448);
and U9518 (N_9518,N_9423,N_9280);
nor U9519 (N_9519,N_9368,N_9393);
nand U9520 (N_9520,N_9376,N_9458);
or U9521 (N_9521,N_9412,N_9434);
and U9522 (N_9522,N_9336,N_9271);
nor U9523 (N_9523,N_9371,N_9441);
or U9524 (N_9524,N_9351,N_9360);
nor U9525 (N_9525,N_9477,N_9338);
nand U9526 (N_9526,N_9459,N_9380);
nor U9527 (N_9527,N_9253,N_9475);
and U9528 (N_9528,N_9395,N_9377);
xnor U9529 (N_9529,N_9345,N_9300);
nor U9530 (N_9530,N_9487,N_9259);
or U9531 (N_9531,N_9270,N_9387);
nand U9532 (N_9532,N_9355,N_9386);
nor U9533 (N_9533,N_9298,N_9457);
xor U9534 (N_9534,N_9341,N_9327);
nor U9535 (N_9535,N_9404,N_9282);
and U9536 (N_9536,N_9323,N_9476);
nor U9537 (N_9537,N_9491,N_9373);
nor U9538 (N_9538,N_9264,N_9367);
nor U9539 (N_9539,N_9409,N_9408);
nor U9540 (N_9540,N_9443,N_9472);
and U9541 (N_9541,N_9346,N_9399);
nor U9542 (N_9542,N_9440,N_9274);
and U9543 (N_9543,N_9402,N_9486);
nand U9544 (N_9544,N_9405,N_9428);
nand U9545 (N_9545,N_9357,N_9384);
nor U9546 (N_9546,N_9406,N_9349);
and U9547 (N_9547,N_9281,N_9347);
nor U9548 (N_9548,N_9414,N_9366);
nand U9549 (N_9549,N_9410,N_9392);
nand U9550 (N_9550,N_9488,N_9452);
nand U9551 (N_9551,N_9471,N_9389);
nand U9552 (N_9552,N_9263,N_9467);
nor U9553 (N_9553,N_9314,N_9313);
or U9554 (N_9554,N_9401,N_9333);
nand U9555 (N_9555,N_9444,N_9375);
or U9556 (N_9556,N_9292,N_9424);
nand U9557 (N_9557,N_9268,N_9407);
nor U9558 (N_9558,N_9363,N_9311);
nor U9559 (N_9559,N_9287,N_9272);
and U9560 (N_9560,N_9258,N_9342);
nor U9561 (N_9561,N_9316,N_9302);
nor U9562 (N_9562,N_9413,N_9461);
or U9563 (N_9563,N_9446,N_9261);
and U9564 (N_9564,N_9285,N_9481);
nand U9565 (N_9565,N_9463,N_9331);
or U9566 (N_9566,N_9445,N_9330);
and U9567 (N_9567,N_9437,N_9421);
and U9568 (N_9568,N_9493,N_9466);
nor U9569 (N_9569,N_9297,N_9329);
nor U9570 (N_9570,N_9304,N_9391);
or U9571 (N_9571,N_9359,N_9352);
or U9572 (N_9572,N_9398,N_9462);
or U9573 (N_9573,N_9374,N_9431);
xor U9574 (N_9574,N_9381,N_9328);
nor U9575 (N_9575,N_9332,N_9254);
and U9576 (N_9576,N_9269,N_9483);
and U9577 (N_9577,N_9456,N_9301);
nor U9578 (N_9578,N_9353,N_9343);
and U9579 (N_9579,N_9256,N_9339);
nand U9580 (N_9580,N_9415,N_9265);
nor U9581 (N_9581,N_9422,N_9464);
nor U9582 (N_9582,N_9266,N_9418);
and U9583 (N_9583,N_9317,N_9482);
nand U9584 (N_9584,N_9354,N_9286);
nor U9585 (N_9585,N_9290,N_9273);
nand U9586 (N_9586,N_9315,N_9251);
or U9587 (N_9587,N_9480,N_9447);
nand U9588 (N_9588,N_9291,N_9453);
nand U9589 (N_9589,N_9474,N_9460);
nand U9590 (N_9590,N_9425,N_9348);
nand U9591 (N_9591,N_9365,N_9484);
and U9592 (N_9592,N_9396,N_9433);
nand U9593 (N_9593,N_9490,N_9296);
nor U9594 (N_9594,N_9420,N_9324);
nor U9595 (N_9595,N_9283,N_9435);
and U9596 (N_9596,N_9485,N_9288);
nand U9597 (N_9597,N_9306,N_9494);
and U9598 (N_9598,N_9320,N_9489);
nor U9599 (N_9599,N_9255,N_9322);
nor U9600 (N_9600,N_9496,N_9379);
or U9601 (N_9601,N_9340,N_9250);
nand U9602 (N_9602,N_9388,N_9439);
nand U9603 (N_9603,N_9455,N_9473);
or U9604 (N_9604,N_9495,N_9252);
nor U9605 (N_9605,N_9307,N_9454);
or U9606 (N_9606,N_9370,N_9275);
nor U9607 (N_9607,N_9390,N_9382);
nand U9608 (N_9608,N_9369,N_9378);
nor U9609 (N_9609,N_9294,N_9318);
and U9610 (N_9610,N_9310,N_9350);
and U9611 (N_9611,N_9325,N_9499);
nor U9612 (N_9612,N_9321,N_9312);
or U9613 (N_9613,N_9262,N_9426);
or U9614 (N_9614,N_9308,N_9337);
or U9615 (N_9615,N_9492,N_9293);
nor U9616 (N_9616,N_9438,N_9479);
nand U9617 (N_9617,N_9429,N_9468);
and U9618 (N_9618,N_9394,N_9470);
nor U9619 (N_9619,N_9364,N_9362);
nor U9620 (N_9620,N_9319,N_9295);
nor U9621 (N_9621,N_9361,N_9498);
or U9622 (N_9622,N_9305,N_9442);
nand U9623 (N_9623,N_9303,N_9478);
and U9624 (N_9624,N_9436,N_9427);
nor U9625 (N_9625,N_9350,N_9430);
nand U9626 (N_9626,N_9421,N_9372);
nand U9627 (N_9627,N_9406,N_9347);
or U9628 (N_9628,N_9408,N_9344);
nand U9629 (N_9629,N_9397,N_9363);
nor U9630 (N_9630,N_9462,N_9439);
or U9631 (N_9631,N_9421,N_9397);
nor U9632 (N_9632,N_9288,N_9389);
or U9633 (N_9633,N_9484,N_9483);
nor U9634 (N_9634,N_9352,N_9394);
nand U9635 (N_9635,N_9409,N_9286);
or U9636 (N_9636,N_9431,N_9254);
nand U9637 (N_9637,N_9262,N_9442);
nand U9638 (N_9638,N_9271,N_9360);
and U9639 (N_9639,N_9293,N_9366);
xnor U9640 (N_9640,N_9431,N_9436);
or U9641 (N_9641,N_9462,N_9314);
nor U9642 (N_9642,N_9496,N_9350);
and U9643 (N_9643,N_9393,N_9486);
nor U9644 (N_9644,N_9463,N_9326);
and U9645 (N_9645,N_9254,N_9360);
or U9646 (N_9646,N_9480,N_9430);
or U9647 (N_9647,N_9279,N_9472);
nand U9648 (N_9648,N_9421,N_9434);
nor U9649 (N_9649,N_9453,N_9394);
nand U9650 (N_9650,N_9317,N_9410);
and U9651 (N_9651,N_9389,N_9419);
or U9652 (N_9652,N_9324,N_9274);
and U9653 (N_9653,N_9337,N_9253);
and U9654 (N_9654,N_9288,N_9270);
or U9655 (N_9655,N_9308,N_9475);
or U9656 (N_9656,N_9316,N_9476);
nor U9657 (N_9657,N_9256,N_9451);
and U9658 (N_9658,N_9326,N_9319);
and U9659 (N_9659,N_9258,N_9257);
nand U9660 (N_9660,N_9483,N_9433);
and U9661 (N_9661,N_9453,N_9492);
or U9662 (N_9662,N_9428,N_9317);
or U9663 (N_9663,N_9447,N_9423);
or U9664 (N_9664,N_9460,N_9423);
nor U9665 (N_9665,N_9259,N_9316);
and U9666 (N_9666,N_9285,N_9303);
nor U9667 (N_9667,N_9352,N_9297);
nor U9668 (N_9668,N_9375,N_9415);
nor U9669 (N_9669,N_9446,N_9330);
nand U9670 (N_9670,N_9266,N_9351);
nor U9671 (N_9671,N_9341,N_9256);
and U9672 (N_9672,N_9321,N_9411);
or U9673 (N_9673,N_9439,N_9484);
and U9674 (N_9674,N_9360,N_9442);
and U9675 (N_9675,N_9327,N_9332);
and U9676 (N_9676,N_9300,N_9426);
nor U9677 (N_9677,N_9428,N_9309);
or U9678 (N_9678,N_9434,N_9343);
or U9679 (N_9679,N_9283,N_9449);
nor U9680 (N_9680,N_9367,N_9320);
and U9681 (N_9681,N_9255,N_9387);
or U9682 (N_9682,N_9402,N_9326);
or U9683 (N_9683,N_9278,N_9425);
and U9684 (N_9684,N_9359,N_9276);
nor U9685 (N_9685,N_9287,N_9344);
nand U9686 (N_9686,N_9442,N_9353);
or U9687 (N_9687,N_9395,N_9402);
nor U9688 (N_9688,N_9467,N_9392);
nand U9689 (N_9689,N_9346,N_9332);
nor U9690 (N_9690,N_9490,N_9342);
nor U9691 (N_9691,N_9441,N_9252);
nor U9692 (N_9692,N_9376,N_9260);
xnor U9693 (N_9693,N_9420,N_9419);
or U9694 (N_9694,N_9367,N_9333);
and U9695 (N_9695,N_9300,N_9483);
nand U9696 (N_9696,N_9302,N_9289);
or U9697 (N_9697,N_9402,N_9456);
nor U9698 (N_9698,N_9303,N_9350);
nand U9699 (N_9699,N_9369,N_9422);
and U9700 (N_9700,N_9277,N_9397);
and U9701 (N_9701,N_9453,N_9373);
nor U9702 (N_9702,N_9445,N_9474);
or U9703 (N_9703,N_9378,N_9293);
nor U9704 (N_9704,N_9451,N_9448);
and U9705 (N_9705,N_9365,N_9428);
nor U9706 (N_9706,N_9387,N_9367);
and U9707 (N_9707,N_9345,N_9411);
nand U9708 (N_9708,N_9435,N_9406);
nor U9709 (N_9709,N_9284,N_9476);
or U9710 (N_9710,N_9262,N_9381);
and U9711 (N_9711,N_9390,N_9352);
or U9712 (N_9712,N_9486,N_9345);
nand U9713 (N_9713,N_9263,N_9342);
nor U9714 (N_9714,N_9343,N_9403);
nand U9715 (N_9715,N_9360,N_9343);
and U9716 (N_9716,N_9454,N_9368);
and U9717 (N_9717,N_9452,N_9329);
and U9718 (N_9718,N_9326,N_9344);
or U9719 (N_9719,N_9455,N_9252);
nand U9720 (N_9720,N_9415,N_9259);
nand U9721 (N_9721,N_9466,N_9388);
nand U9722 (N_9722,N_9404,N_9262);
and U9723 (N_9723,N_9328,N_9406);
and U9724 (N_9724,N_9318,N_9366);
nand U9725 (N_9725,N_9330,N_9266);
and U9726 (N_9726,N_9260,N_9273);
nand U9727 (N_9727,N_9305,N_9461);
and U9728 (N_9728,N_9354,N_9279);
nand U9729 (N_9729,N_9363,N_9375);
nor U9730 (N_9730,N_9316,N_9291);
or U9731 (N_9731,N_9317,N_9304);
or U9732 (N_9732,N_9461,N_9330);
nor U9733 (N_9733,N_9439,N_9312);
nor U9734 (N_9734,N_9257,N_9489);
and U9735 (N_9735,N_9332,N_9278);
nand U9736 (N_9736,N_9398,N_9426);
nor U9737 (N_9737,N_9396,N_9463);
or U9738 (N_9738,N_9402,N_9442);
nand U9739 (N_9739,N_9362,N_9355);
nor U9740 (N_9740,N_9435,N_9293);
nand U9741 (N_9741,N_9498,N_9337);
nand U9742 (N_9742,N_9447,N_9450);
or U9743 (N_9743,N_9289,N_9449);
or U9744 (N_9744,N_9364,N_9255);
and U9745 (N_9745,N_9354,N_9274);
nor U9746 (N_9746,N_9329,N_9390);
nand U9747 (N_9747,N_9468,N_9405);
or U9748 (N_9748,N_9369,N_9461);
nor U9749 (N_9749,N_9258,N_9428);
and U9750 (N_9750,N_9700,N_9653);
nand U9751 (N_9751,N_9735,N_9610);
nor U9752 (N_9752,N_9508,N_9705);
xor U9753 (N_9753,N_9711,N_9509);
or U9754 (N_9754,N_9746,N_9635);
nor U9755 (N_9755,N_9687,N_9545);
nand U9756 (N_9756,N_9520,N_9590);
nand U9757 (N_9757,N_9578,N_9633);
and U9758 (N_9758,N_9692,N_9629);
and U9759 (N_9759,N_9522,N_9531);
nand U9760 (N_9760,N_9555,N_9521);
nand U9761 (N_9761,N_9631,N_9693);
and U9762 (N_9762,N_9706,N_9716);
nand U9763 (N_9763,N_9533,N_9729);
nor U9764 (N_9764,N_9618,N_9564);
or U9765 (N_9765,N_9620,N_9734);
nand U9766 (N_9766,N_9641,N_9669);
nand U9767 (N_9767,N_9503,N_9595);
nand U9768 (N_9768,N_9501,N_9624);
and U9769 (N_9769,N_9690,N_9698);
nand U9770 (N_9770,N_9607,N_9621);
nand U9771 (N_9771,N_9684,N_9748);
nor U9772 (N_9772,N_9625,N_9691);
or U9773 (N_9773,N_9630,N_9699);
or U9774 (N_9774,N_9666,N_9683);
nand U9775 (N_9775,N_9540,N_9542);
nand U9776 (N_9776,N_9726,N_9642);
nand U9777 (N_9777,N_9678,N_9601);
and U9778 (N_9778,N_9737,N_9597);
or U9779 (N_9779,N_9728,N_9743);
nand U9780 (N_9780,N_9636,N_9619);
or U9781 (N_9781,N_9710,N_9697);
nand U9782 (N_9782,N_9722,N_9721);
nor U9783 (N_9783,N_9534,N_9626);
or U9784 (N_9784,N_9557,N_9550);
and U9785 (N_9785,N_9732,N_9613);
nand U9786 (N_9786,N_9675,N_9541);
nand U9787 (N_9787,N_9548,N_9702);
nand U9788 (N_9788,N_9745,N_9556);
nand U9789 (N_9789,N_9720,N_9696);
nand U9790 (N_9790,N_9530,N_9739);
nor U9791 (N_9791,N_9731,N_9718);
nor U9792 (N_9792,N_9504,N_9709);
or U9793 (N_9793,N_9519,N_9671);
and U9794 (N_9794,N_9615,N_9563);
nand U9795 (N_9795,N_9685,N_9516);
or U9796 (N_9796,N_9525,N_9559);
or U9797 (N_9797,N_9637,N_9688);
or U9798 (N_9798,N_9535,N_9606);
and U9799 (N_9799,N_9605,N_9528);
nor U9800 (N_9800,N_9573,N_9659);
nor U9801 (N_9801,N_9676,N_9612);
nor U9802 (N_9802,N_9565,N_9518);
or U9803 (N_9803,N_9648,N_9523);
or U9804 (N_9804,N_9609,N_9581);
nand U9805 (N_9805,N_9572,N_9713);
nand U9806 (N_9806,N_9513,N_9661);
and U9807 (N_9807,N_9539,N_9517);
and U9808 (N_9808,N_9526,N_9596);
nor U9809 (N_9809,N_9622,N_9674);
and U9810 (N_9810,N_9584,N_9672);
nand U9811 (N_9811,N_9561,N_9667);
or U9812 (N_9812,N_9647,N_9507);
or U9813 (N_9813,N_9547,N_9554);
or U9814 (N_9814,N_9695,N_9591);
or U9815 (N_9815,N_9723,N_9510);
and U9816 (N_9816,N_9654,N_9543);
nand U9817 (N_9817,N_9725,N_9538);
nor U9818 (N_9818,N_9512,N_9511);
nor U9819 (N_9819,N_9611,N_9663);
and U9820 (N_9820,N_9592,N_9657);
or U9821 (N_9821,N_9529,N_9575);
or U9822 (N_9822,N_9680,N_9703);
nand U9823 (N_9823,N_9594,N_9623);
nand U9824 (N_9824,N_9599,N_9682);
nor U9825 (N_9825,N_9727,N_9701);
or U9826 (N_9826,N_9714,N_9640);
nor U9827 (N_9827,N_9740,N_9544);
nand U9828 (N_9828,N_9536,N_9665);
or U9829 (N_9829,N_9562,N_9608);
or U9830 (N_9830,N_9733,N_9628);
nand U9831 (N_9831,N_9558,N_9744);
or U9832 (N_9832,N_9502,N_9662);
nor U9833 (N_9833,N_9668,N_9741);
and U9834 (N_9834,N_9598,N_9579);
xor U9835 (N_9835,N_9551,N_9651);
nand U9836 (N_9836,N_9515,N_9738);
nor U9837 (N_9837,N_9645,N_9566);
or U9838 (N_9838,N_9537,N_9634);
nor U9839 (N_9839,N_9583,N_9664);
or U9840 (N_9840,N_9736,N_9638);
and U9841 (N_9841,N_9712,N_9627);
nor U9842 (N_9842,N_9694,N_9660);
and U9843 (N_9843,N_9603,N_9686);
or U9844 (N_9844,N_9614,N_9724);
and U9845 (N_9845,N_9658,N_9505);
or U9846 (N_9846,N_9719,N_9639);
or U9847 (N_9847,N_9704,N_9589);
nor U9848 (N_9848,N_9587,N_9552);
or U9849 (N_9849,N_9568,N_9707);
or U9850 (N_9850,N_9715,N_9500);
xnor U9851 (N_9851,N_9616,N_9649);
nand U9852 (N_9852,N_9679,N_9546);
and U9853 (N_9853,N_9650,N_9656);
and U9854 (N_9854,N_9532,N_9749);
nand U9855 (N_9855,N_9717,N_9574);
and U9856 (N_9856,N_9646,N_9582);
or U9857 (N_9857,N_9689,N_9553);
or U9858 (N_9858,N_9567,N_9569);
or U9859 (N_9859,N_9708,N_9580);
nor U9860 (N_9860,N_9681,N_9600);
nor U9861 (N_9861,N_9570,N_9643);
and U9862 (N_9862,N_9673,N_9585);
nor U9863 (N_9863,N_9560,N_9506);
or U9864 (N_9864,N_9742,N_9604);
nand U9865 (N_9865,N_9730,N_9670);
and U9866 (N_9866,N_9576,N_9524);
nand U9867 (N_9867,N_9514,N_9602);
and U9868 (N_9868,N_9652,N_9617);
or U9869 (N_9869,N_9571,N_9549);
nand U9870 (N_9870,N_9644,N_9632);
nor U9871 (N_9871,N_9747,N_9527);
and U9872 (N_9872,N_9577,N_9586);
nor U9873 (N_9873,N_9655,N_9593);
nor U9874 (N_9874,N_9677,N_9588);
nor U9875 (N_9875,N_9637,N_9685);
and U9876 (N_9876,N_9512,N_9642);
nand U9877 (N_9877,N_9689,N_9598);
nor U9878 (N_9878,N_9531,N_9640);
nor U9879 (N_9879,N_9504,N_9542);
or U9880 (N_9880,N_9640,N_9649);
or U9881 (N_9881,N_9598,N_9655);
nor U9882 (N_9882,N_9548,N_9697);
nand U9883 (N_9883,N_9728,N_9614);
nor U9884 (N_9884,N_9648,N_9733);
nand U9885 (N_9885,N_9554,N_9585);
nand U9886 (N_9886,N_9683,N_9664);
and U9887 (N_9887,N_9732,N_9700);
nand U9888 (N_9888,N_9502,N_9650);
or U9889 (N_9889,N_9538,N_9552);
and U9890 (N_9890,N_9733,N_9536);
nor U9891 (N_9891,N_9515,N_9624);
nand U9892 (N_9892,N_9730,N_9635);
or U9893 (N_9893,N_9553,N_9589);
and U9894 (N_9894,N_9517,N_9530);
and U9895 (N_9895,N_9736,N_9688);
nor U9896 (N_9896,N_9633,N_9672);
and U9897 (N_9897,N_9667,N_9627);
nor U9898 (N_9898,N_9666,N_9655);
or U9899 (N_9899,N_9599,N_9747);
and U9900 (N_9900,N_9650,N_9595);
or U9901 (N_9901,N_9517,N_9673);
and U9902 (N_9902,N_9531,N_9570);
nand U9903 (N_9903,N_9506,N_9718);
nor U9904 (N_9904,N_9696,N_9587);
nor U9905 (N_9905,N_9551,N_9693);
and U9906 (N_9906,N_9516,N_9557);
nand U9907 (N_9907,N_9595,N_9724);
and U9908 (N_9908,N_9693,N_9586);
and U9909 (N_9909,N_9709,N_9609);
nor U9910 (N_9910,N_9632,N_9555);
and U9911 (N_9911,N_9625,N_9743);
and U9912 (N_9912,N_9515,N_9592);
nand U9913 (N_9913,N_9630,N_9575);
nor U9914 (N_9914,N_9625,N_9685);
nand U9915 (N_9915,N_9597,N_9748);
and U9916 (N_9916,N_9684,N_9572);
or U9917 (N_9917,N_9600,N_9654);
and U9918 (N_9918,N_9606,N_9652);
nand U9919 (N_9919,N_9713,N_9626);
and U9920 (N_9920,N_9718,N_9676);
or U9921 (N_9921,N_9585,N_9544);
and U9922 (N_9922,N_9638,N_9558);
nand U9923 (N_9923,N_9630,N_9690);
or U9924 (N_9924,N_9655,N_9569);
or U9925 (N_9925,N_9586,N_9553);
and U9926 (N_9926,N_9654,N_9684);
nand U9927 (N_9927,N_9585,N_9665);
nand U9928 (N_9928,N_9691,N_9650);
and U9929 (N_9929,N_9518,N_9735);
nor U9930 (N_9930,N_9639,N_9721);
nand U9931 (N_9931,N_9737,N_9720);
or U9932 (N_9932,N_9747,N_9601);
nor U9933 (N_9933,N_9609,N_9642);
nand U9934 (N_9934,N_9614,N_9531);
nand U9935 (N_9935,N_9628,N_9621);
nor U9936 (N_9936,N_9588,N_9713);
nor U9937 (N_9937,N_9504,N_9731);
nand U9938 (N_9938,N_9568,N_9534);
or U9939 (N_9939,N_9623,N_9663);
nor U9940 (N_9940,N_9680,N_9621);
nand U9941 (N_9941,N_9512,N_9668);
or U9942 (N_9942,N_9641,N_9719);
or U9943 (N_9943,N_9654,N_9659);
nor U9944 (N_9944,N_9616,N_9680);
nor U9945 (N_9945,N_9554,N_9660);
and U9946 (N_9946,N_9695,N_9615);
nand U9947 (N_9947,N_9671,N_9640);
nand U9948 (N_9948,N_9673,N_9653);
nor U9949 (N_9949,N_9559,N_9660);
nand U9950 (N_9950,N_9549,N_9739);
nand U9951 (N_9951,N_9621,N_9682);
xor U9952 (N_9952,N_9681,N_9663);
or U9953 (N_9953,N_9612,N_9539);
nor U9954 (N_9954,N_9511,N_9525);
nand U9955 (N_9955,N_9626,N_9607);
or U9956 (N_9956,N_9588,N_9676);
and U9957 (N_9957,N_9543,N_9689);
nand U9958 (N_9958,N_9664,N_9576);
and U9959 (N_9959,N_9700,N_9585);
nor U9960 (N_9960,N_9543,N_9675);
and U9961 (N_9961,N_9621,N_9544);
nand U9962 (N_9962,N_9518,N_9647);
and U9963 (N_9963,N_9629,N_9564);
nor U9964 (N_9964,N_9710,N_9736);
or U9965 (N_9965,N_9608,N_9530);
and U9966 (N_9966,N_9694,N_9629);
nand U9967 (N_9967,N_9545,N_9588);
and U9968 (N_9968,N_9628,N_9645);
or U9969 (N_9969,N_9730,N_9651);
nand U9970 (N_9970,N_9571,N_9664);
nor U9971 (N_9971,N_9580,N_9730);
or U9972 (N_9972,N_9515,N_9708);
and U9973 (N_9973,N_9508,N_9696);
nand U9974 (N_9974,N_9647,N_9629);
or U9975 (N_9975,N_9531,N_9508);
nand U9976 (N_9976,N_9513,N_9533);
nor U9977 (N_9977,N_9554,N_9558);
or U9978 (N_9978,N_9567,N_9659);
or U9979 (N_9979,N_9553,N_9699);
or U9980 (N_9980,N_9591,N_9526);
nor U9981 (N_9981,N_9711,N_9556);
nand U9982 (N_9982,N_9618,N_9512);
nor U9983 (N_9983,N_9519,N_9722);
nor U9984 (N_9984,N_9550,N_9706);
or U9985 (N_9985,N_9689,N_9644);
and U9986 (N_9986,N_9588,N_9598);
nor U9987 (N_9987,N_9512,N_9546);
or U9988 (N_9988,N_9613,N_9664);
nand U9989 (N_9989,N_9537,N_9728);
nand U9990 (N_9990,N_9579,N_9660);
xnor U9991 (N_9991,N_9611,N_9667);
nand U9992 (N_9992,N_9671,N_9606);
nand U9993 (N_9993,N_9700,N_9705);
and U9994 (N_9994,N_9541,N_9734);
and U9995 (N_9995,N_9735,N_9569);
and U9996 (N_9996,N_9724,N_9572);
or U9997 (N_9997,N_9523,N_9557);
and U9998 (N_9998,N_9667,N_9721);
nand U9999 (N_9999,N_9590,N_9514);
nor U10000 (N_10000,N_9899,N_9817);
and U10001 (N_10001,N_9815,N_9757);
nor U10002 (N_10002,N_9845,N_9987);
nor U10003 (N_10003,N_9751,N_9909);
nand U10004 (N_10004,N_9996,N_9814);
nand U10005 (N_10005,N_9758,N_9787);
or U10006 (N_10006,N_9847,N_9761);
nor U10007 (N_10007,N_9916,N_9795);
and U10008 (N_10008,N_9828,N_9753);
or U10009 (N_10009,N_9980,N_9784);
or U10010 (N_10010,N_9781,N_9999);
nor U10011 (N_10011,N_9837,N_9906);
and U10012 (N_10012,N_9914,N_9908);
nand U10013 (N_10013,N_9883,N_9913);
xor U10014 (N_10014,N_9963,N_9968);
and U10015 (N_10015,N_9919,N_9940);
and U10016 (N_10016,N_9953,N_9839);
nand U10017 (N_10017,N_9827,N_9907);
and U10018 (N_10018,N_9918,N_9971);
and U10019 (N_10019,N_9994,N_9863);
or U10020 (N_10020,N_9892,N_9820);
and U10021 (N_10021,N_9951,N_9886);
nand U10022 (N_10022,N_9850,N_9796);
nor U10023 (N_10023,N_9838,N_9920);
nand U10024 (N_10024,N_9842,N_9976);
or U10025 (N_10025,N_9860,N_9959);
or U10026 (N_10026,N_9877,N_9912);
nor U10027 (N_10027,N_9865,N_9923);
or U10028 (N_10028,N_9969,N_9970);
and U10029 (N_10029,N_9788,N_9926);
or U10030 (N_10030,N_9864,N_9823);
nor U10031 (N_10031,N_9754,N_9997);
and U10032 (N_10032,N_9874,N_9779);
nor U10033 (N_10033,N_9786,N_9873);
nand U10034 (N_10034,N_9986,N_9775);
and U10035 (N_10035,N_9856,N_9984);
nor U10036 (N_10036,N_9910,N_9879);
and U10037 (N_10037,N_9958,N_9843);
or U10038 (N_10038,N_9866,N_9898);
nand U10039 (N_10039,N_9915,N_9922);
or U10040 (N_10040,N_9891,N_9948);
nor U10041 (N_10041,N_9861,N_9844);
nor U10042 (N_10042,N_9790,N_9826);
or U10043 (N_10043,N_9871,N_9981);
or U10044 (N_10044,N_9966,N_9943);
or U10045 (N_10045,N_9887,N_9832);
or U10046 (N_10046,N_9936,N_9835);
and U10047 (N_10047,N_9829,N_9840);
and U10048 (N_10048,N_9851,N_9917);
and U10049 (N_10049,N_9854,N_9962);
nor U10050 (N_10050,N_9858,N_9880);
or U10051 (N_10051,N_9799,N_9950);
and U10052 (N_10052,N_9807,N_9960);
or U10053 (N_10053,N_9965,N_9768);
or U10054 (N_10054,N_9763,N_9766);
nand U10055 (N_10055,N_9830,N_9804);
or U10056 (N_10056,N_9805,N_9993);
and U10057 (N_10057,N_9872,N_9957);
nor U10058 (N_10058,N_9985,N_9777);
nand U10059 (N_10059,N_9895,N_9875);
and U10060 (N_10060,N_9927,N_9961);
nor U10061 (N_10061,N_9888,N_9822);
and U10062 (N_10062,N_9897,N_9789);
nor U10063 (N_10063,N_9780,N_9982);
nand U10064 (N_10064,N_9989,N_9932);
nand U10065 (N_10065,N_9811,N_9983);
and U10066 (N_10066,N_9855,N_9939);
nand U10067 (N_10067,N_9967,N_9785);
or U10068 (N_10068,N_9988,N_9764);
nand U10069 (N_10069,N_9849,N_9806);
and U10070 (N_10070,N_9762,N_9931);
nor U10071 (N_10071,N_9778,N_9797);
nand U10072 (N_10072,N_9769,N_9995);
or U10073 (N_10073,N_9890,N_9870);
nand U10074 (N_10074,N_9972,N_9824);
or U10075 (N_10075,N_9848,N_9859);
and U10076 (N_10076,N_9798,N_9928);
or U10077 (N_10077,N_9938,N_9801);
nand U10078 (N_10078,N_9752,N_9750);
or U10079 (N_10079,N_9770,N_9974);
nor U10080 (N_10080,N_9867,N_9911);
nor U10081 (N_10081,N_9760,N_9954);
nor U10082 (N_10082,N_9808,N_9852);
and U10083 (N_10083,N_9925,N_9884);
nor U10084 (N_10084,N_9782,N_9944);
nor U10085 (N_10085,N_9949,N_9836);
and U10086 (N_10086,N_9952,N_9862);
nand U10087 (N_10087,N_9929,N_9973);
or U10088 (N_10088,N_9809,N_9755);
or U10089 (N_10089,N_9990,N_9978);
nor U10090 (N_10090,N_9846,N_9889);
and U10091 (N_10091,N_9885,N_9869);
and U10092 (N_10092,N_9937,N_9825);
or U10093 (N_10093,N_9853,N_9765);
nor U10094 (N_10094,N_9813,N_9818);
nand U10095 (N_10095,N_9904,N_9894);
and U10096 (N_10096,N_9902,N_9810);
nor U10097 (N_10097,N_9868,N_9771);
or U10098 (N_10098,N_9945,N_9900);
or U10099 (N_10099,N_9774,N_9794);
nor U10100 (N_10100,N_9924,N_9776);
and U10101 (N_10101,N_9800,N_9882);
and U10102 (N_10102,N_9756,N_9930);
nand U10103 (N_10103,N_9992,N_9921);
nor U10104 (N_10104,N_9956,N_9792);
or U10105 (N_10105,N_9979,N_9975);
or U10106 (N_10106,N_9881,N_9772);
nor U10107 (N_10107,N_9998,N_9964);
and U10108 (N_10108,N_9935,N_9841);
nand U10109 (N_10109,N_9802,N_9947);
and U10110 (N_10110,N_9783,N_9803);
or U10111 (N_10111,N_9934,N_9791);
and U10112 (N_10112,N_9773,N_9905);
nor U10113 (N_10113,N_9821,N_9876);
nand U10114 (N_10114,N_9896,N_9878);
nand U10115 (N_10115,N_9903,N_9834);
or U10116 (N_10116,N_9816,N_9941);
nand U10117 (N_10117,N_9942,N_9812);
or U10118 (N_10118,N_9831,N_9946);
and U10119 (N_10119,N_9977,N_9819);
or U10120 (N_10120,N_9901,N_9955);
nor U10121 (N_10121,N_9893,N_9991);
and U10122 (N_10122,N_9793,N_9767);
and U10123 (N_10123,N_9833,N_9759);
nor U10124 (N_10124,N_9933,N_9857);
and U10125 (N_10125,N_9874,N_9843);
and U10126 (N_10126,N_9996,N_9778);
nor U10127 (N_10127,N_9882,N_9865);
nor U10128 (N_10128,N_9823,N_9989);
nor U10129 (N_10129,N_9752,N_9969);
nand U10130 (N_10130,N_9997,N_9753);
or U10131 (N_10131,N_9797,N_9962);
nor U10132 (N_10132,N_9982,N_9892);
nand U10133 (N_10133,N_9902,N_9758);
or U10134 (N_10134,N_9750,N_9764);
and U10135 (N_10135,N_9909,N_9904);
nor U10136 (N_10136,N_9829,N_9831);
nand U10137 (N_10137,N_9843,N_9852);
nand U10138 (N_10138,N_9920,N_9876);
or U10139 (N_10139,N_9790,N_9916);
nand U10140 (N_10140,N_9781,N_9906);
nand U10141 (N_10141,N_9889,N_9989);
nand U10142 (N_10142,N_9907,N_9824);
or U10143 (N_10143,N_9926,N_9770);
nand U10144 (N_10144,N_9948,N_9803);
nor U10145 (N_10145,N_9931,N_9889);
and U10146 (N_10146,N_9939,N_9787);
and U10147 (N_10147,N_9781,N_9828);
nand U10148 (N_10148,N_9882,N_9804);
nand U10149 (N_10149,N_9996,N_9965);
nor U10150 (N_10150,N_9990,N_9956);
or U10151 (N_10151,N_9822,N_9885);
nand U10152 (N_10152,N_9937,N_9770);
nor U10153 (N_10153,N_9864,N_9918);
or U10154 (N_10154,N_9780,N_9950);
and U10155 (N_10155,N_9966,N_9837);
and U10156 (N_10156,N_9910,N_9817);
or U10157 (N_10157,N_9801,N_9911);
and U10158 (N_10158,N_9762,N_9857);
or U10159 (N_10159,N_9801,N_9889);
nand U10160 (N_10160,N_9808,N_9886);
or U10161 (N_10161,N_9845,N_9849);
nor U10162 (N_10162,N_9880,N_9879);
nor U10163 (N_10163,N_9937,N_9816);
nand U10164 (N_10164,N_9901,N_9927);
nor U10165 (N_10165,N_9959,N_9908);
nand U10166 (N_10166,N_9750,N_9760);
nand U10167 (N_10167,N_9787,N_9782);
nand U10168 (N_10168,N_9904,N_9771);
nand U10169 (N_10169,N_9931,N_9783);
and U10170 (N_10170,N_9981,N_9797);
and U10171 (N_10171,N_9818,N_9982);
and U10172 (N_10172,N_9870,N_9961);
or U10173 (N_10173,N_9904,N_9984);
nand U10174 (N_10174,N_9753,N_9820);
or U10175 (N_10175,N_9916,N_9862);
nor U10176 (N_10176,N_9869,N_9999);
nand U10177 (N_10177,N_9975,N_9930);
nor U10178 (N_10178,N_9827,N_9882);
nand U10179 (N_10179,N_9882,N_9758);
and U10180 (N_10180,N_9890,N_9887);
nand U10181 (N_10181,N_9964,N_9921);
nor U10182 (N_10182,N_9947,N_9878);
xnor U10183 (N_10183,N_9874,N_9891);
nand U10184 (N_10184,N_9781,N_9924);
and U10185 (N_10185,N_9971,N_9830);
and U10186 (N_10186,N_9903,N_9847);
nor U10187 (N_10187,N_9967,N_9831);
and U10188 (N_10188,N_9895,N_9927);
and U10189 (N_10189,N_9958,N_9841);
nor U10190 (N_10190,N_9925,N_9814);
nand U10191 (N_10191,N_9793,N_9927);
nand U10192 (N_10192,N_9850,N_9768);
or U10193 (N_10193,N_9810,N_9968);
nor U10194 (N_10194,N_9871,N_9786);
nor U10195 (N_10195,N_9951,N_9814);
and U10196 (N_10196,N_9994,N_9846);
nor U10197 (N_10197,N_9965,N_9840);
and U10198 (N_10198,N_9881,N_9861);
nand U10199 (N_10199,N_9880,N_9899);
or U10200 (N_10200,N_9816,N_9883);
or U10201 (N_10201,N_9950,N_9905);
and U10202 (N_10202,N_9785,N_9842);
nand U10203 (N_10203,N_9791,N_9991);
and U10204 (N_10204,N_9763,N_9905);
or U10205 (N_10205,N_9990,N_9860);
nor U10206 (N_10206,N_9839,N_9984);
nand U10207 (N_10207,N_9781,N_9752);
and U10208 (N_10208,N_9882,N_9854);
nand U10209 (N_10209,N_9765,N_9832);
and U10210 (N_10210,N_9919,N_9929);
nand U10211 (N_10211,N_9984,N_9913);
or U10212 (N_10212,N_9838,N_9855);
and U10213 (N_10213,N_9929,N_9803);
or U10214 (N_10214,N_9874,N_9774);
and U10215 (N_10215,N_9886,N_9781);
or U10216 (N_10216,N_9886,N_9841);
nor U10217 (N_10217,N_9893,N_9964);
and U10218 (N_10218,N_9850,N_9861);
or U10219 (N_10219,N_9788,N_9898);
nor U10220 (N_10220,N_9914,N_9809);
and U10221 (N_10221,N_9797,N_9872);
or U10222 (N_10222,N_9772,N_9890);
or U10223 (N_10223,N_9925,N_9931);
and U10224 (N_10224,N_9818,N_9856);
or U10225 (N_10225,N_9766,N_9899);
nand U10226 (N_10226,N_9793,N_9979);
nor U10227 (N_10227,N_9967,N_9864);
nor U10228 (N_10228,N_9769,N_9815);
and U10229 (N_10229,N_9803,N_9765);
xor U10230 (N_10230,N_9900,N_9777);
or U10231 (N_10231,N_9987,N_9985);
and U10232 (N_10232,N_9861,N_9998);
nand U10233 (N_10233,N_9984,N_9831);
nand U10234 (N_10234,N_9829,N_9940);
or U10235 (N_10235,N_9791,N_9966);
nor U10236 (N_10236,N_9966,N_9959);
or U10237 (N_10237,N_9804,N_9972);
and U10238 (N_10238,N_9955,N_9935);
nor U10239 (N_10239,N_9927,N_9750);
and U10240 (N_10240,N_9911,N_9835);
nor U10241 (N_10241,N_9801,N_9920);
nor U10242 (N_10242,N_9844,N_9773);
nand U10243 (N_10243,N_9879,N_9918);
nor U10244 (N_10244,N_9758,N_9996);
or U10245 (N_10245,N_9760,N_9762);
or U10246 (N_10246,N_9813,N_9770);
nor U10247 (N_10247,N_9774,N_9827);
nor U10248 (N_10248,N_9983,N_9952);
and U10249 (N_10249,N_9863,N_9846);
nand U10250 (N_10250,N_10095,N_10135);
nand U10251 (N_10251,N_10166,N_10069);
nand U10252 (N_10252,N_10220,N_10131);
or U10253 (N_10253,N_10128,N_10205);
and U10254 (N_10254,N_10134,N_10045);
nand U10255 (N_10255,N_10017,N_10203);
and U10256 (N_10256,N_10155,N_10225);
and U10257 (N_10257,N_10013,N_10178);
nand U10258 (N_10258,N_10073,N_10190);
and U10259 (N_10259,N_10014,N_10108);
nor U10260 (N_10260,N_10080,N_10103);
or U10261 (N_10261,N_10026,N_10195);
and U10262 (N_10262,N_10099,N_10194);
nor U10263 (N_10263,N_10024,N_10201);
or U10264 (N_10264,N_10081,N_10027);
nand U10265 (N_10265,N_10188,N_10023);
nor U10266 (N_10266,N_10115,N_10151);
nand U10267 (N_10267,N_10010,N_10158);
and U10268 (N_10268,N_10067,N_10143);
and U10269 (N_10269,N_10210,N_10110);
and U10270 (N_10270,N_10226,N_10048);
nand U10271 (N_10271,N_10041,N_10053);
nand U10272 (N_10272,N_10090,N_10156);
nor U10273 (N_10273,N_10047,N_10102);
nor U10274 (N_10274,N_10167,N_10025);
nand U10275 (N_10275,N_10062,N_10022);
nor U10276 (N_10276,N_10057,N_10191);
and U10277 (N_10277,N_10060,N_10239);
nor U10278 (N_10278,N_10176,N_10211);
nor U10279 (N_10279,N_10231,N_10005);
xor U10280 (N_10280,N_10170,N_10089);
nand U10281 (N_10281,N_10147,N_10182);
and U10282 (N_10282,N_10165,N_10033);
or U10283 (N_10283,N_10198,N_10031);
nand U10284 (N_10284,N_10145,N_10177);
nor U10285 (N_10285,N_10181,N_10248);
nor U10286 (N_10286,N_10002,N_10237);
nand U10287 (N_10287,N_10107,N_10127);
nor U10288 (N_10288,N_10240,N_10034);
nand U10289 (N_10289,N_10228,N_10119);
and U10290 (N_10290,N_10111,N_10114);
and U10291 (N_10291,N_10121,N_10079);
nand U10292 (N_10292,N_10000,N_10233);
or U10293 (N_10293,N_10172,N_10137);
nor U10294 (N_10294,N_10008,N_10097);
nand U10295 (N_10295,N_10243,N_10153);
or U10296 (N_10296,N_10179,N_10072);
nor U10297 (N_10297,N_10019,N_10204);
or U10298 (N_10298,N_10193,N_10049);
nor U10299 (N_10299,N_10154,N_10076);
nor U10300 (N_10300,N_10174,N_10219);
nor U10301 (N_10301,N_10068,N_10140);
nor U10302 (N_10302,N_10052,N_10037);
nand U10303 (N_10303,N_10015,N_10215);
nand U10304 (N_10304,N_10106,N_10206);
nand U10305 (N_10305,N_10104,N_10249);
or U10306 (N_10306,N_10118,N_10163);
nand U10307 (N_10307,N_10141,N_10035);
nand U10308 (N_10308,N_10087,N_10064);
and U10309 (N_10309,N_10180,N_10032);
and U10310 (N_10310,N_10112,N_10075);
nand U10311 (N_10311,N_10117,N_10105);
and U10312 (N_10312,N_10244,N_10129);
or U10313 (N_10313,N_10171,N_10161);
and U10314 (N_10314,N_10085,N_10186);
and U10315 (N_10315,N_10217,N_10216);
and U10316 (N_10316,N_10212,N_10199);
or U10317 (N_10317,N_10150,N_10036);
and U10318 (N_10318,N_10044,N_10184);
nand U10319 (N_10319,N_10120,N_10149);
nand U10320 (N_10320,N_10020,N_10222);
and U10321 (N_10321,N_10055,N_10189);
nand U10322 (N_10322,N_10230,N_10098);
or U10323 (N_10323,N_10007,N_10183);
or U10324 (N_10324,N_10058,N_10218);
and U10325 (N_10325,N_10136,N_10246);
nand U10326 (N_10326,N_10046,N_10051);
or U10327 (N_10327,N_10175,N_10125);
nor U10328 (N_10328,N_10030,N_10213);
and U10329 (N_10329,N_10078,N_10004);
nand U10330 (N_10330,N_10133,N_10234);
nand U10331 (N_10331,N_10071,N_10096);
and U10332 (N_10332,N_10227,N_10202);
or U10333 (N_10333,N_10245,N_10235);
nor U10334 (N_10334,N_10092,N_10223);
or U10335 (N_10335,N_10187,N_10113);
nor U10336 (N_10336,N_10192,N_10162);
and U10337 (N_10337,N_10148,N_10061);
nand U10338 (N_10338,N_10232,N_10159);
or U10339 (N_10339,N_10006,N_10039);
or U10340 (N_10340,N_10050,N_10021);
or U10341 (N_10341,N_10056,N_10146);
nand U10342 (N_10342,N_10157,N_10173);
nand U10343 (N_10343,N_10065,N_10236);
nor U10344 (N_10344,N_10139,N_10241);
nand U10345 (N_10345,N_10042,N_10238);
nand U10346 (N_10346,N_10082,N_10001);
nor U10347 (N_10347,N_10028,N_10130);
nor U10348 (N_10348,N_10091,N_10122);
nand U10349 (N_10349,N_10208,N_10088);
nor U10350 (N_10350,N_10063,N_10038);
nand U10351 (N_10351,N_10164,N_10074);
and U10352 (N_10352,N_10054,N_10040);
or U10353 (N_10353,N_10168,N_10160);
and U10354 (N_10354,N_10066,N_10242);
or U10355 (N_10355,N_10116,N_10123);
or U10356 (N_10356,N_10138,N_10221);
nor U10357 (N_10357,N_10209,N_10124);
or U10358 (N_10358,N_10200,N_10016);
and U10359 (N_10359,N_10207,N_10083);
and U10360 (N_10360,N_10101,N_10003);
xnor U10361 (N_10361,N_10012,N_10185);
or U10362 (N_10362,N_10093,N_10011);
and U10363 (N_10363,N_10077,N_10018);
nand U10364 (N_10364,N_10094,N_10152);
and U10365 (N_10365,N_10169,N_10214);
nand U10366 (N_10366,N_10142,N_10197);
and U10367 (N_10367,N_10144,N_10247);
nand U10368 (N_10368,N_10132,N_10229);
nor U10369 (N_10369,N_10109,N_10059);
nor U10370 (N_10370,N_10086,N_10029);
or U10371 (N_10371,N_10100,N_10196);
or U10372 (N_10372,N_10126,N_10009);
nand U10373 (N_10373,N_10043,N_10084);
nor U10374 (N_10374,N_10070,N_10224);
and U10375 (N_10375,N_10095,N_10066);
or U10376 (N_10376,N_10072,N_10039);
nor U10377 (N_10377,N_10111,N_10168);
nor U10378 (N_10378,N_10224,N_10105);
and U10379 (N_10379,N_10225,N_10107);
or U10380 (N_10380,N_10077,N_10082);
and U10381 (N_10381,N_10084,N_10204);
nor U10382 (N_10382,N_10002,N_10231);
and U10383 (N_10383,N_10127,N_10000);
and U10384 (N_10384,N_10019,N_10157);
nand U10385 (N_10385,N_10156,N_10037);
nand U10386 (N_10386,N_10154,N_10089);
and U10387 (N_10387,N_10157,N_10135);
and U10388 (N_10388,N_10247,N_10083);
or U10389 (N_10389,N_10134,N_10165);
and U10390 (N_10390,N_10088,N_10129);
nor U10391 (N_10391,N_10120,N_10188);
and U10392 (N_10392,N_10210,N_10125);
nor U10393 (N_10393,N_10005,N_10098);
nor U10394 (N_10394,N_10004,N_10007);
or U10395 (N_10395,N_10159,N_10077);
nand U10396 (N_10396,N_10249,N_10227);
or U10397 (N_10397,N_10078,N_10096);
and U10398 (N_10398,N_10098,N_10160);
nor U10399 (N_10399,N_10155,N_10198);
nor U10400 (N_10400,N_10009,N_10197);
and U10401 (N_10401,N_10110,N_10064);
nor U10402 (N_10402,N_10002,N_10141);
nor U10403 (N_10403,N_10177,N_10021);
or U10404 (N_10404,N_10152,N_10040);
or U10405 (N_10405,N_10045,N_10169);
nor U10406 (N_10406,N_10099,N_10166);
and U10407 (N_10407,N_10086,N_10020);
or U10408 (N_10408,N_10195,N_10192);
xor U10409 (N_10409,N_10096,N_10196);
and U10410 (N_10410,N_10145,N_10064);
nand U10411 (N_10411,N_10152,N_10011);
nor U10412 (N_10412,N_10194,N_10219);
nor U10413 (N_10413,N_10181,N_10199);
or U10414 (N_10414,N_10077,N_10024);
and U10415 (N_10415,N_10004,N_10061);
nand U10416 (N_10416,N_10150,N_10097);
nor U10417 (N_10417,N_10245,N_10103);
nor U10418 (N_10418,N_10134,N_10205);
nor U10419 (N_10419,N_10213,N_10241);
or U10420 (N_10420,N_10114,N_10227);
and U10421 (N_10421,N_10067,N_10058);
nor U10422 (N_10422,N_10197,N_10018);
and U10423 (N_10423,N_10143,N_10208);
and U10424 (N_10424,N_10206,N_10027);
or U10425 (N_10425,N_10214,N_10094);
nand U10426 (N_10426,N_10117,N_10081);
nand U10427 (N_10427,N_10226,N_10068);
and U10428 (N_10428,N_10168,N_10029);
nor U10429 (N_10429,N_10190,N_10067);
and U10430 (N_10430,N_10111,N_10165);
nand U10431 (N_10431,N_10138,N_10192);
nor U10432 (N_10432,N_10112,N_10237);
or U10433 (N_10433,N_10101,N_10005);
or U10434 (N_10434,N_10079,N_10235);
nor U10435 (N_10435,N_10152,N_10068);
nor U10436 (N_10436,N_10097,N_10135);
or U10437 (N_10437,N_10122,N_10092);
nor U10438 (N_10438,N_10040,N_10149);
and U10439 (N_10439,N_10152,N_10247);
or U10440 (N_10440,N_10024,N_10208);
or U10441 (N_10441,N_10126,N_10071);
or U10442 (N_10442,N_10065,N_10074);
and U10443 (N_10443,N_10200,N_10067);
and U10444 (N_10444,N_10101,N_10026);
nand U10445 (N_10445,N_10024,N_10202);
and U10446 (N_10446,N_10078,N_10104);
nand U10447 (N_10447,N_10217,N_10240);
or U10448 (N_10448,N_10008,N_10131);
or U10449 (N_10449,N_10119,N_10125);
nor U10450 (N_10450,N_10180,N_10057);
and U10451 (N_10451,N_10248,N_10190);
and U10452 (N_10452,N_10062,N_10123);
nor U10453 (N_10453,N_10189,N_10006);
nand U10454 (N_10454,N_10185,N_10247);
nand U10455 (N_10455,N_10232,N_10198);
or U10456 (N_10456,N_10240,N_10060);
nand U10457 (N_10457,N_10202,N_10076);
nor U10458 (N_10458,N_10187,N_10066);
xnor U10459 (N_10459,N_10231,N_10000);
or U10460 (N_10460,N_10031,N_10151);
or U10461 (N_10461,N_10005,N_10064);
nor U10462 (N_10462,N_10013,N_10029);
nand U10463 (N_10463,N_10207,N_10092);
and U10464 (N_10464,N_10079,N_10027);
nor U10465 (N_10465,N_10052,N_10225);
nand U10466 (N_10466,N_10148,N_10048);
nor U10467 (N_10467,N_10127,N_10098);
and U10468 (N_10468,N_10075,N_10187);
nor U10469 (N_10469,N_10075,N_10065);
nor U10470 (N_10470,N_10089,N_10093);
nand U10471 (N_10471,N_10236,N_10095);
and U10472 (N_10472,N_10009,N_10205);
nor U10473 (N_10473,N_10124,N_10202);
nor U10474 (N_10474,N_10003,N_10055);
nand U10475 (N_10475,N_10210,N_10107);
nand U10476 (N_10476,N_10067,N_10082);
and U10477 (N_10477,N_10248,N_10026);
nand U10478 (N_10478,N_10153,N_10037);
and U10479 (N_10479,N_10030,N_10023);
nand U10480 (N_10480,N_10014,N_10217);
or U10481 (N_10481,N_10210,N_10002);
and U10482 (N_10482,N_10164,N_10179);
and U10483 (N_10483,N_10121,N_10099);
nand U10484 (N_10484,N_10107,N_10001);
nand U10485 (N_10485,N_10219,N_10213);
and U10486 (N_10486,N_10218,N_10038);
nor U10487 (N_10487,N_10034,N_10044);
nor U10488 (N_10488,N_10037,N_10214);
nand U10489 (N_10489,N_10033,N_10105);
and U10490 (N_10490,N_10138,N_10124);
nor U10491 (N_10491,N_10159,N_10012);
or U10492 (N_10492,N_10025,N_10191);
nand U10493 (N_10493,N_10227,N_10211);
nor U10494 (N_10494,N_10039,N_10247);
nor U10495 (N_10495,N_10026,N_10024);
or U10496 (N_10496,N_10192,N_10014);
or U10497 (N_10497,N_10207,N_10157);
and U10498 (N_10498,N_10062,N_10104);
nand U10499 (N_10499,N_10013,N_10193);
nand U10500 (N_10500,N_10353,N_10289);
and U10501 (N_10501,N_10448,N_10252);
and U10502 (N_10502,N_10413,N_10326);
nand U10503 (N_10503,N_10327,N_10317);
or U10504 (N_10504,N_10393,N_10320);
nand U10505 (N_10505,N_10277,N_10390);
nor U10506 (N_10506,N_10485,N_10375);
and U10507 (N_10507,N_10286,N_10358);
nor U10508 (N_10508,N_10492,N_10355);
or U10509 (N_10509,N_10288,N_10481);
xnor U10510 (N_10510,N_10444,N_10278);
nand U10511 (N_10511,N_10346,N_10428);
xor U10512 (N_10512,N_10308,N_10285);
and U10513 (N_10513,N_10426,N_10356);
and U10514 (N_10514,N_10360,N_10334);
or U10515 (N_10515,N_10427,N_10385);
and U10516 (N_10516,N_10420,N_10298);
nand U10517 (N_10517,N_10363,N_10330);
nand U10518 (N_10518,N_10272,N_10409);
or U10519 (N_10519,N_10265,N_10387);
nand U10520 (N_10520,N_10386,N_10279);
or U10521 (N_10521,N_10379,N_10264);
nor U10522 (N_10522,N_10318,N_10276);
nand U10523 (N_10523,N_10435,N_10496);
and U10524 (N_10524,N_10497,N_10486);
nor U10525 (N_10525,N_10433,N_10395);
and U10526 (N_10526,N_10484,N_10449);
or U10527 (N_10527,N_10431,N_10441);
nor U10528 (N_10528,N_10365,N_10401);
nor U10529 (N_10529,N_10478,N_10464);
or U10530 (N_10530,N_10407,N_10312);
or U10531 (N_10531,N_10302,N_10342);
nand U10532 (N_10532,N_10383,N_10488);
or U10533 (N_10533,N_10324,N_10367);
nor U10534 (N_10534,N_10335,N_10479);
or U10535 (N_10535,N_10414,N_10362);
and U10536 (N_10536,N_10472,N_10344);
nor U10537 (N_10537,N_10493,N_10377);
or U10538 (N_10538,N_10260,N_10301);
nor U10539 (N_10539,N_10352,N_10261);
or U10540 (N_10540,N_10354,N_10452);
and U10541 (N_10541,N_10253,N_10439);
or U10542 (N_10542,N_10305,N_10349);
nor U10543 (N_10543,N_10384,N_10462);
and U10544 (N_10544,N_10477,N_10376);
nor U10545 (N_10545,N_10315,N_10474);
and U10546 (N_10546,N_10311,N_10434);
or U10547 (N_10547,N_10406,N_10307);
nand U10548 (N_10548,N_10498,N_10491);
nand U10549 (N_10549,N_10371,N_10469);
nand U10550 (N_10550,N_10259,N_10430);
nor U10551 (N_10551,N_10490,N_10391);
nand U10552 (N_10552,N_10350,N_10471);
and U10553 (N_10553,N_10304,N_10299);
nand U10554 (N_10554,N_10446,N_10382);
or U10555 (N_10555,N_10399,N_10280);
nor U10556 (N_10556,N_10411,N_10432);
nand U10557 (N_10557,N_10313,N_10389);
or U10558 (N_10558,N_10332,N_10348);
and U10559 (N_10559,N_10329,N_10268);
and U10560 (N_10560,N_10297,N_10405);
or U10561 (N_10561,N_10270,N_10489);
and U10562 (N_10562,N_10412,N_10416);
nand U10563 (N_10563,N_10467,N_10321);
nor U10564 (N_10564,N_10293,N_10404);
nor U10565 (N_10565,N_10263,N_10480);
and U10566 (N_10566,N_10473,N_10392);
and U10567 (N_10567,N_10372,N_10456);
nand U10568 (N_10568,N_10423,N_10408);
nor U10569 (N_10569,N_10368,N_10262);
nor U10570 (N_10570,N_10410,N_10458);
and U10571 (N_10571,N_10457,N_10400);
or U10572 (N_10572,N_10338,N_10483);
nor U10573 (N_10573,N_10466,N_10257);
nor U10574 (N_10574,N_10361,N_10269);
nor U10575 (N_10575,N_10255,N_10316);
and U10576 (N_10576,N_10380,N_10282);
nand U10577 (N_10577,N_10419,N_10374);
or U10578 (N_10578,N_10397,N_10254);
nor U10579 (N_10579,N_10422,N_10266);
and U10580 (N_10580,N_10442,N_10396);
nor U10581 (N_10581,N_10284,N_10487);
nor U10582 (N_10582,N_10323,N_10463);
and U10583 (N_10583,N_10271,N_10455);
or U10584 (N_10584,N_10388,N_10429);
nor U10585 (N_10585,N_10369,N_10402);
and U10586 (N_10586,N_10461,N_10283);
and U10587 (N_10587,N_10443,N_10476);
or U10588 (N_10588,N_10294,N_10394);
nand U10589 (N_10589,N_10273,N_10447);
or U10590 (N_10590,N_10341,N_10303);
and U10591 (N_10591,N_10359,N_10291);
nand U10592 (N_10592,N_10495,N_10425);
and U10593 (N_10593,N_10421,N_10281);
and U10594 (N_10594,N_10418,N_10251);
nand U10595 (N_10595,N_10424,N_10328);
nor U10596 (N_10596,N_10314,N_10296);
nand U10597 (N_10597,N_10440,N_10470);
nor U10598 (N_10598,N_10322,N_10373);
xor U10599 (N_10599,N_10347,N_10459);
nor U10600 (N_10600,N_10287,N_10465);
nor U10601 (N_10601,N_10319,N_10290);
and U10602 (N_10602,N_10364,N_10494);
and U10603 (N_10603,N_10445,N_10258);
nor U10604 (N_10604,N_10436,N_10460);
and U10605 (N_10605,N_10453,N_10450);
and U10606 (N_10606,N_10300,N_10468);
and U10607 (N_10607,N_10482,N_10345);
nand U10608 (N_10608,N_10398,N_10357);
or U10609 (N_10609,N_10370,N_10339);
or U10610 (N_10610,N_10310,N_10454);
nand U10611 (N_10611,N_10267,N_10351);
nand U10612 (N_10612,N_10306,N_10250);
and U10613 (N_10613,N_10337,N_10274);
and U10614 (N_10614,N_10331,N_10415);
and U10615 (N_10615,N_10451,N_10340);
and U10616 (N_10616,N_10275,N_10378);
and U10617 (N_10617,N_10333,N_10336);
nor U10618 (N_10618,N_10475,N_10417);
and U10619 (N_10619,N_10499,N_10256);
nor U10620 (N_10620,N_10437,N_10292);
or U10621 (N_10621,N_10381,N_10325);
nor U10622 (N_10622,N_10403,N_10343);
nand U10623 (N_10623,N_10295,N_10309);
nor U10624 (N_10624,N_10366,N_10438);
and U10625 (N_10625,N_10333,N_10337);
or U10626 (N_10626,N_10378,N_10398);
and U10627 (N_10627,N_10355,N_10259);
nor U10628 (N_10628,N_10463,N_10321);
nand U10629 (N_10629,N_10306,N_10353);
nor U10630 (N_10630,N_10267,N_10454);
and U10631 (N_10631,N_10473,N_10368);
or U10632 (N_10632,N_10252,N_10362);
nor U10633 (N_10633,N_10454,N_10327);
or U10634 (N_10634,N_10359,N_10297);
nand U10635 (N_10635,N_10482,N_10422);
nand U10636 (N_10636,N_10284,N_10455);
and U10637 (N_10637,N_10409,N_10422);
nand U10638 (N_10638,N_10369,N_10463);
and U10639 (N_10639,N_10265,N_10455);
and U10640 (N_10640,N_10376,N_10451);
nor U10641 (N_10641,N_10419,N_10400);
nand U10642 (N_10642,N_10397,N_10316);
and U10643 (N_10643,N_10347,N_10350);
or U10644 (N_10644,N_10321,N_10478);
and U10645 (N_10645,N_10392,N_10317);
and U10646 (N_10646,N_10451,N_10390);
nand U10647 (N_10647,N_10315,N_10355);
nand U10648 (N_10648,N_10372,N_10388);
or U10649 (N_10649,N_10481,N_10306);
or U10650 (N_10650,N_10483,N_10321);
nand U10651 (N_10651,N_10319,N_10279);
nor U10652 (N_10652,N_10474,N_10312);
and U10653 (N_10653,N_10344,N_10302);
or U10654 (N_10654,N_10424,N_10287);
nor U10655 (N_10655,N_10485,N_10432);
or U10656 (N_10656,N_10373,N_10351);
and U10657 (N_10657,N_10321,N_10437);
nor U10658 (N_10658,N_10367,N_10448);
nor U10659 (N_10659,N_10252,N_10270);
and U10660 (N_10660,N_10308,N_10426);
nor U10661 (N_10661,N_10318,N_10437);
and U10662 (N_10662,N_10268,N_10384);
and U10663 (N_10663,N_10294,N_10444);
nor U10664 (N_10664,N_10424,N_10266);
nand U10665 (N_10665,N_10320,N_10455);
nor U10666 (N_10666,N_10329,N_10497);
nand U10667 (N_10667,N_10384,N_10301);
or U10668 (N_10668,N_10257,N_10433);
xor U10669 (N_10669,N_10318,N_10396);
and U10670 (N_10670,N_10291,N_10284);
and U10671 (N_10671,N_10268,N_10340);
nand U10672 (N_10672,N_10284,N_10253);
or U10673 (N_10673,N_10271,N_10488);
nor U10674 (N_10674,N_10344,N_10369);
nor U10675 (N_10675,N_10349,N_10422);
or U10676 (N_10676,N_10278,N_10308);
nand U10677 (N_10677,N_10329,N_10350);
nand U10678 (N_10678,N_10310,N_10251);
or U10679 (N_10679,N_10320,N_10275);
nand U10680 (N_10680,N_10292,N_10431);
nand U10681 (N_10681,N_10384,N_10385);
or U10682 (N_10682,N_10467,N_10266);
or U10683 (N_10683,N_10479,N_10344);
and U10684 (N_10684,N_10438,N_10313);
nand U10685 (N_10685,N_10398,N_10325);
nor U10686 (N_10686,N_10467,N_10372);
nand U10687 (N_10687,N_10462,N_10472);
and U10688 (N_10688,N_10452,N_10365);
or U10689 (N_10689,N_10318,N_10268);
nor U10690 (N_10690,N_10273,N_10407);
or U10691 (N_10691,N_10402,N_10258);
and U10692 (N_10692,N_10414,N_10440);
nor U10693 (N_10693,N_10413,N_10382);
nand U10694 (N_10694,N_10369,N_10357);
nand U10695 (N_10695,N_10302,N_10300);
nor U10696 (N_10696,N_10386,N_10355);
or U10697 (N_10697,N_10443,N_10298);
nand U10698 (N_10698,N_10428,N_10322);
nand U10699 (N_10699,N_10461,N_10475);
or U10700 (N_10700,N_10324,N_10262);
nor U10701 (N_10701,N_10388,N_10443);
nand U10702 (N_10702,N_10425,N_10492);
or U10703 (N_10703,N_10467,N_10466);
nor U10704 (N_10704,N_10387,N_10487);
nor U10705 (N_10705,N_10399,N_10457);
nor U10706 (N_10706,N_10282,N_10267);
nor U10707 (N_10707,N_10275,N_10269);
nor U10708 (N_10708,N_10374,N_10459);
nand U10709 (N_10709,N_10304,N_10339);
or U10710 (N_10710,N_10493,N_10403);
or U10711 (N_10711,N_10438,N_10345);
nand U10712 (N_10712,N_10417,N_10481);
or U10713 (N_10713,N_10402,N_10435);
or U10714 (N_10714,N_10464,N_10473);
or U10715 (N_10715,N_10341,N_10282);
and U10716 (N_10716,N_10291,N_10427);
or U10717 (N_10717,N_10367,N_10360);
and U10718 (N_10718,N_10439,N_10322);
and U10719 (N_10719,N_10436,N_10393);
or U10720 (N_10720,N_10267,N_10330);
and U10721 (N_10721,N_10447,N_10490);
nand U10722 (N_10722,N_10344,N_10305);
or U10723 (N_10723,N_10282,N_10272);
nor U10724 (N_10724,N_10429,N_10282);
nand U10725 (N_10725,N_10459,N_10445);
and U10726 (N_10726,N_10273,N_10403);
nand U10727 (N_10727,N_10403,N_10460);
or U10728 (N_10728,N_10430,N_10470);
nand U10729 (N_10729,N_10292,N_10306);
and U10730 (N_10730,N_10369,N_10270);
and U10731 (N_10731,N_10495,N_10295);
nand U10732 (N_10732,N_10304,N_10364);
nor U10733 (N_10733,N_10345,N_10387);
nand U10734 (N_10734,N_10267,N_10328);
nor U10735 (N_10735,N_10494,N_10448);
and U10736 (N_10736,N_10417,N_10482);
nor U10737 (N_10737,N_10275,N_10261);
or U10738 (N_10738,N_10355,N_10379);
nand U10739 (N_10739,N_10254,N_10281);
nor U10740 (N_10740,N_10445,N_10302);
nor U10741 (N_10741,N_10416,N_10482);
or U10742 (N_10742,N_10324,N_10327);
or U10743 (N_10743,N_10378,N_10499);
nor U10744 (N_10744,N_10487,N_10358);
nor U10745 (N_10745,N_10320,N_10484);
or U10746 (N_10746,N_10359,N_10255);
or U10747 (N_10747,N_10379,N_10338);
nand U10748 (N_10748,N_10357,N_10466);
nor U10749 (N_10749,N_10294,N_10460);
and U10750 (N_10750,N_10604,N_10714);
nand U10751 (N_10751,N_10600,N_10742);
and U10752 (N_10752,N_10655,N_10623);
nand U10753 (N_10753,N_10612,N_10534);
and U10754 (N_10754,N_10730,N_10706);
nand U10755 (N_10755,N_10522,N_10658);
and U10756 (N_10756,N_10628,N_10682);
or U10757 (N_10757,N_10713,N_10544);
nor U10758 (N_10758,N_10716,N_10618);
or U10759 (N_10759,N_10694,N_10577);
nor U10760 (N_10760,N_10509,N_10624);
xor U10761 (N_10761,N_10698,N_10657);
or U10762 (N_10762,N_10631,N_10603);
nor U10763 (N_10763,N_10681,N_10507);
or U10764 (N_10764,N_10661,N_10591);
nor U10765 (N_10765,N_10506,N_10725);
xor U10766 (N_10766,N_10527,N_10526);
and U10767 (N_10767,N_10503,N_10584);
or U10768 (N_10768,N_10557,N_10643);
nor U10769 (N_10769,N_10673,N_10552);
and U10770 (N_10770,N_10626,N_10668);
and U10771 (N_10771,N_10546,N_10662);
and U10772 (N_10772,N_10633,N_10564);
and U10773 (N_10773,N_10656,N_10708);
and U10774 (N_10774,N_10531,N_10639);
or U10775 (N_10775,N_10644,N_10518);
or U10776 (N_10776,N_10563,N_10501);
nor U10777 (N_10777,N_10703,N_10724);
and U10778 (N_10778,N_10739,N_10620);
nor U10779 (N_10779,N_10717,N_10660);
and U10780 (N_10780,N_10685,N_10671);
or U10781 (N_10781,N_10593,N_10736);
and U10782 (N_10782,N_10561,N_10636);
or U10783 (N_10783,N_10590,N_10523);
nor U10784 (N_10784,N_10511,N_10516);
nand U10785 (N_10785,N_10740,N_10621);
or U10786 (N_10786,N_10615,N_10539);
nor U10787 (N_10787,N_10700,N_10529);
or U10788 (N_10788,N_10635,N_10535);
and U10789 (N_10789,N_10687,N_10719);
or U10790 (N_10790,N_10568,N_10670);
xnor U10791 (N_10791,N_10537,N_10723);
nand U10792 (N_10792,N_10689,N_10630);
nand U10793 (N_10793,N_10517,N_10669);
or U10794 (N_10794,N_10744,N_10536);
nand U10795 (N_10795,N_10582,N_10560);
nor U10796 (N_10796,N_10596,N_10580);
and U10797 (N_10797,N_10602,N_10638);
or U10798 (N_10798,N_10553,N_10570);
and U10799 (N_10799,N_10665,N_10538);
nor U10800 (N_10800,N_10699,N_10543);
or U10801 (N_10801,N_10693,N_10556);
nand U10802 (N_10802,N_10540,N_10542);
and U10803 (N_10803,N_10521,N_10738);
and U10804 (N_10804,N_10586,N_10504);
or U10805 (N_10805,N_10711,N_10675);
and U10806 (N_10806,N_10663,N_10550);
or U10807 (N_10807,N_10642,N_10674);
nor U10808 (N_10808,N_10562,N_10734);
and U10809 (N_10809,N_10705,N_10571);
nor U10810 (N_10810,N_10667,N_10599);
nand U10811 (N_10811,N_10619,N_10710);
nand U10812 (N_10812,N_10555,N_10709);
or U10813 (N_10813,N_10745,N_10651);
nor U10814 (N_10814,N_10650,N_10525);
or U10815 (N_10815,N_10608,N_10583);
or U10816 (N_10816,N_10659,N_10541);
nor U10817 (N_10817,N_10653,N_10721);
nand U10818 (N_10818,N_10566,N_10647);
nand U10819 (N_10819,N_10545,N_10614);
and U10820 (N_10820,N_10679,N_10569);
nor U10821 (N_10821,N_10722,N_10617);
nor U10822 (N_10822,N_10533,N_10733);
nor U10823 (N_10823,N_10585,N_10601);
and U10824 (N_10824,N_10688,N_10524);
nor U10825 (N_10825,N_10718,N_10589);
nor U10826 (N_10826,N_10575,N_10735);
or U10827 (N_10827,N_10666,N_10567);
or U10828 (N_10828,N_10727,N_10677);
or U10829 (N_10829,N_10747,N_10547);
nand U10830 (N_10830,N_10640,N_10696);
nand U10831 (N_10831,N_10729,N_10587);
nand U10832 (N_10832,N_10559,N_10512);
nor U10833 (N_10833,N_10737,N_10672);
nand U10834 (N_10834,N_10548,N_10692);
nand U10835 (N_10835,N_10519,N_10707);
nand U10836 (N_10836,N_10500,N_10572);
nor U10837 (N_10837,N_10678,N_10588);
nor U10838 (N_10838,N_10549,N_10578);
or U10839 (N_10839,N_10664,N_10554);
nor U10840 (N_10840,N_10610,N_10646);
nand U10841 (N_10841,N_10625,N_10513);
or U10842 (N_10842,N_10613,N_10505);
and U10843 (N_10843,N_10690,N_10607);
and U10844 (N_10844,N_10715,N_10514);
nand U10845 (N_10845,N_10712,N_10605);
or U10846 (N_10846,N_10528,N_10592);
or U10847 (N_10847,N_10691,N_10728);
or U10848 (N_10848,N_10627,N_10576);
or U10849 (N_10849,N_10530,N_10520);
nand U10850 (N_10850,N_10558,N_10641);
nand U10851 (N_10851,N_10684,N_10743);
or U10852 (N_10852,N_10574,N_10749);
nor U10853 (N_10853,N_10616,N_10573);
or U10854 (N_10854,N_10702,N_10532);
and U10855 (N_10855,N_10579,N_10697);
or U10856 (N_10856,N_10649,N_10510);
nor U10857 (N_10857,N_10508,N_10645);
or U10858 (N_10858,N_10606,N_10720);
nor U10859 (N_10859,N_10732,N_10680);
nor U10860 (N_10860,N_10632,N_10611);
nand U10861 (N_10861,N_10648,N_10598);
and U10862 (N_10862,N_10634,N_10551);
nand U10863 (N_10863,N_10637,N_10695);
or U10864 (N_10864,N_10741,N_10622);
xor U10865 (N_10865,N_10683,N_10597);
nand U10866 (N_10866,N_10676,N_10731);
and U10867 (N_10867,N_10652,N_10515);
and U10868 (N_10868,N_10726,N_10686);
or U10869 (N_10869,N_10609,N_10746);
and U10870 (N_10870,N_10502,N_10701);
or U10871 (N_10871,N_10748,N_10594);
nor U10872 (N_10872,N_10704,N_10595);
nor U10873 (N_10873,N_10654,N_10581);
and U10874 (N_10874,N_10629,N_10565);
nand U10875 (N_10875,N_10644,N_10706);
nand U10876 (N_10876,N_10668,N_10602);
and U10877 (N_10877,N_10667,N_10715);
nor U10878 (N_10878,N_10518,N_10673);
nand U10879 (N_10879,N_10701,N_10686);
or U10880 (N_10880,N_10596,N_10531);
or U10881 (N_10881,N_10519,N_10711);
and U10882 (N_10882,N_10555,N_10595);
nor U10883 (N_10883,N_10691,N_10651);
and U10884 (N_10884,N_10707,N_10590);
or U10885 (N_10885,N_10621,N_10577);
nand U10886 (N_10886,N_10516,N_10609);
and U10887 (N_10887,N_10668,N_10747);
nand U10888 (N_10888,N_10688,N_10644);
or U10889 (N_10889,N_10721,N_10549);
or U10890 (N_10890,N_10731,N_10562);
and U10891 (N_10891,N_10669,N_10702);
nor U10892 (N_10892,N_10557,N_10628);
and U10893 (N_10893,N_10662,N_10689);
nor U10894 (N_10894,N_10649,N_10626);
and U10895 (N_10895,N_10545,N_10528);
nand U10896 (N_10896,N_10552,N_10581);
and U10897 (N_10897,N_10538,N_10742);
nor U10898 (N_10898,N_10632,N_10679);
or U10899 (N_10899,N_10515,N_10575);
nand U10900 (N_10900,N_10566,N_10706);
nand U10901 (N_10901,N_10535,N_10500);
and U10902 (N_10902,N_10692,N_10699);
and U10903 (N_10903,N_10568,N_10732);
and U10904 (N_10904,N_10739,N_10691);
or U10905 (N_10905,N_10566,N_10628);
or U10906 (N_10906,N_10511,N_10685);
or U10907 (N_10907,N_10638,N_10521);
nor U10908 (N_10908,N_10529,N_10721);
nand U10909 (N_10909,N_10596,N_10588);
or U10910 (N_10910,N_10643,N_10608);
or U10911 (N_10911,N_10644,N_10585);
or U10912 (N_10912,N_10557,N_10598);
nor U10913 (N_10913,N_10566,N_10658);
or U10914 (N_10914,N_10736,N_10569);
nor U10915 (N_10915,N_10517,N_10676);
nor U10916 (N_10916,N_10581,N_10507);
nand U10917 (N_10917,N_10644,N_10720);
and U10918 (N_10918,N_10514,N_10508);
and U10919 (N_10919,N_10535,N_10538);
or U10920 (N_10920,N_10608,N_10563);
and U10921 (N_10921,N_10554,N_10568);
nor U10922 (N_10922,N_10519,N_10565);
and U10923 (N_10923,N_10722,N_10624);
nand U10924 (N_10924,N_10712,N_10720);
nor U10925 (N_10925,N_10673,N_10701);
or U10926 (N_10926,N_10646,N_10519);
or U10927 (N_10927,N_10638,N_10641);
nor U10928 (N_10928,N_10522,N_10648);
nand U10929 (N_10929,N_10742,N_10577);
and U10930 (N_10930,N_10725,N_10568);
nor U10931 (N_10931,N_10701,N_10600);
or U10932 (N_10932,N_10500,N_10544);
nor U10933 (N_10933,N_10704,N_10598);
or U10934 (N_10934,N_10630,N_10519);
or U10935 (N_10935,N_10608,N_10531);
or U10936 (N_10936,N_10562,N_10692);
xor U10937 (N_10937,N_10614,N_10685);
or U10938 (N_10938,N_10503,N_10695);
or U10939 (N_10939,N_10618,N_10632);
or U10940 (N_10940,N_10537,N_10613);
nand U10941 (N_10941,N_10537,N_10639);
and U10942 (N_10942,N_10604,N_10525);
nand U10943 (N_10943,N_10666,N_10539);
or U10944 (N_10944,N_10509,N_10690);
and U10945 (N_10945,N_10699,N_10670);
or U10946 (N_10946,N_10601,N_10708);
or U10947 (N_10947,N_10562,N_10694);
and U10948 (N_10948,N_10690,N_10683);
and U10949 (N_10949,N_10582,N_10747);
nor U10950 (N_10950,N_10576,N_10746);
nand U10951 (N_10951,N_10513,N_10615);
nor U10952 (N_10952,N_10600,N_10559);
nand U10953 (N_10953,N_10626,N_10524);
nand U10954 (N_10954,N_10509,N_10718);
nand U10955 (N_10955,N_10676,N_10524);
nor U10956 (N_10956,N_10734,N_10561);
nor U10957 (N_10957,N_10640,N_10723);
and U10958 (N_10958,N_10511,N_10558);
nor U10959 (N_10959,N_10634,N_10507);
nor U10960 (N_10960,N_10603,N_10724);
and U10961 (N_10961,N_10745,N_10678);
nor U10962 (N_10962,N_10705,N_10550);
nor U10963 (N_10963,N_10525,N_10655);
and U10964 (N_10964,N_10507,N_10524);
nand U10965 (N_10965,N_10692,N_10514);
nand U10966 (N_10966,N_10701,N_10694);
xor U10967 (N_10967,N_10575,N_10707);
and U10968 (N_10968,N_10690,N_10640);
and U10969 (N_10969,N_10557,N_10702);
nor U10970 (N_10970,N_10676,N_10513);
nand U10971 (N_10971,N_10524,N_10596);
nor U10972 (N_10972,N_10525,N_10573);
nor U10973 (N_10973,N_10707,N_10581);
nor U10974 (N_10974,N_10662,N_10702);
nand U10975 (N_10975,N_10558,N_10646);
nor U10976 (N_10976,N_10711,N_10545);
nand U10977 (N_10977,N_10595,N_10541);
nand U10978 (N_10978,N_10668,N_10557);
or U10979 (N_10979,N_10741,N_10645);
nand U10980 (N_10980,N_10599,N_10681);
and U10981 (N_10981,N_10553,N_10500);
nor U10982 (N_10982,N_10737,N_10682);
or U10983 (N_10983,N_10514,N_10645);
nand U10984 (N_10984,N_10687,N_10710);
and U10985 (N_10985,N_10590,N_10745);
and U10986 (N_10986,N_10708,N_10591);
nor U10987 (N_10987,N_10558,N_10612);
nand U10988 (N_10988,N_10652,N_10739);
and U10989 (N_10989,N_10632,N_10597);
or U10990 (N_10990,N_10524,N_10527);
and U10991 (N_10991,N_10611,N_10539);
nor U10992 (N_10992,N_10622,N_10637);
nor U10993 (N_10993,N_10679,N_10648);
and U10994 (N_10994,N_10588,N_10713);
nor U10995 (N_10995,N_10595,N_10625);
nand U10996 (N_10996,N_10582,N_10717);
nand U10997 (N_10997,N_10714,N_10537);
nand U10998 (N_10998,N_10652,N_10577);
nor U10999 (N_10999,N_10566,N_10518);
and U11000 (N_11000,N_10826,N_10882);
nand U11001 (N_11001,N_10953,N_10888);
nor U11002 (N_11002,N_10768,N_10968);
nand U11003 (N_11003,N_10774,N_10755);
nand U11004 (N_11004,N_10947,N_10944);
nor U11005 (N_11005,N_10868,N_10884);
nand U11006 (N_11006,N_10941,N_10853);
nor U11007 (N_11007,N_10756,N_10914);
nor U11008 (N_11008,N_10913,N_10872);
nor U11009 (N_11009,N_10759,N_10804);
or U11010 (N_11010,N_10843,N_10906);
nand U11011 (N_11011,N_10835,N_10790);
and U11012 (N_11012,N_10878,N_10877);
nand U11013 (N_11013,N_10943,N_10919);
and U11014 (N_11014,N_10827,N_10809);
nor U11015 (N_11015,N_10824,N_10945);
and U11016 (N_11016,N_10891,N_10963);
or U11017 (N_11017,N_10829,N_10795);
or U11018 (N_11018,N_10987,N_10840);
or U11019 (N_11019,N_10848,N_10846);
and U11020 (N_11020,N_10983,N_10787);
and U11021 (N_11021,N_10961,N_10937);
nand U11022 (N_11022,N_10907,N_10808);
and U11023 (N_11023,N_10917,N_10817);
nor U11024 (N_11024,N_10856,N_10793);
nand U11025 (N_11025,N_10926,N_10858);
nand U11026 (N_11026,N_10940,N_10973);
or U11027 (N_11027,N_10845,N_10777);
and U11028 (N_11028,N_10839,N_10874);
and U11029 (N_11029,N_10875,N_10933);
nand U11030 (N_11030,N_10936,N_10828);
and U11031 (N_11031,N_10986,N_10866);
and U11032 (N_11032,N_10977,N_10960);
or U11033 (N_11033,N_10908,N_10894);
nand U11034 (N_11034,N_10762,N_10818);
or U11035 (N_11035,N_10763,N_10964);
and U11036 (N_11036,N_10922,N_10863);
and U11037 (N_11037,N_10772,N_10887);
nor U11038 (N_11038,N_10816,N_10991);
nand U11039 (N_11039,N_10970,N_10998);
nand U11040 (N_11040,N_10813,N_10903);
nand U11041 (N_11041,N_10912,N_10844);
or U11042 (N_11042,N_10796,N_10916);
nor U11043 (N_11043,N_10832,N_10948);
nor U11044 (N_11044,N_10957,N_10938);
and U11045 (N_11045,N_10930,N_10880);
nor U11046 (N_11046,N_10847,N_10904);
and U11047 (N_11047,N_10834,N_10852);
nor U11048 (N_11048,N_10886,N_10988);
and U11049 (N_11049,N_10995,N_10867);
nor U11050 (N_11050,N_10982,N_10897);
and U11051 (N_11051,N_10879,N_10791);
nor U11052 (N_11052,N_10905,N_10876);
nand U11053 (N_11053,N_10931,N_10929);
nand U11054 (N_11054,N_10965,N_10767);
nand U11055 (N_11055,N_10836,N_10918);
and U11056 (N_11056,N_10859,N_10994);
or U11057 (N_11057,N_10924,N_10902);
and U11058 (N_11058,N_10959,N_10927);
nor U11059 (N_11059,N_10925,N_10911);
and U11060 (N_11060,N_10823,N_10934);
nor U11061 (N_11061,N_10871,N_10942);
nor U11062 (N_11062,N_10923,N_10939);
nor U11063 (N_11063,N_10990,N_10788);
nor U11064 (N_11064,N_10833,N_10900);
and U11065 (N_11065,N_10864,N_10785);
nand U11066 (N_11066,N_10773,N_10792);
nand U11067 (N_11067,N_10811,N_10869);
nor U11068 (N_11068,N_10889,N_10985);
and U11069 (N_11069,N_10805,N_10975);
nor U11070 (N_11070,N_10758,N_10753);
nand U11071 (N_11071,N_10781,N_10801);
or U11072 (N_11072,N_10849,N_10831);
nand U11073 (N_11073,N_10760,N_10855);
nor U11074 (N_11074,N_10800,N_10954);
xnor U11075 (N_11075,N_10783,N_10861);
and U11076 (N_11076,N_10949,N_10842);
nor U11077 (N_11077,N_10766,N_10896);
or U11078 (N_11078,N_10819,N_10799);
and U11079 (N_11079,N_10771,N_10993);
and U11080 (N_11080,N_10780,N_10898);
nand U11081 (N_11081,N_10794,N_10893);
and U11082 (N_11082,N_10892,N_10857);
or U11083 (N_11083,N_10761,N_10976);
nor U11084 (N_11084,N_10946,N_10950);
nor U11085 (N_11085,N_10769,N_10757);
or U11086 (N_11086,N_10822,N_10786);
or U11087 (N_11087,N_10978,N_10776);
and U11088 (N_11088,N_10765,N_10971);
and U11089 (N_11089,N_10810,N_10992);
nor U11090 (N_11090,N_10750,N_10881);
nor U11091 (N_11091,N_10807,N_10873);
nand U11092 (N_11092,N_10782,N_10751);
nor U11093 (N_11093,N_10979,N_10920);
nor U11094 (N_11094,N_10915,N_10981);
nand U11095 (N_11095,N_10797,N_10806);
or U11096 (N_11096,N_10865,N_10837);
and U11097 (N_11097,N_10972,N_10784);
xor U11098 (N_11098,N_10984,N_10958);
and U11099 (N_11099,N_10870,N_10770);
nor U11100 (N_11100,N_10838,N_10798);
nor U11101 (N_11101,N_10996,N_10775);
nand U11102 (N_11102,N_10778,N_10779);
or U11103 (N_11103,N_10830,N_10921);
nor U11104 (N_11104,N_10928,N_10812);
or U11105 (N_11105,N_10754,N_10862);
nor U11106 (N_11106,N_10969,N_10899);
or U11107 (N_11107,N_10752,N_10989);
nand U11108 (N_11108,N_10821,N_10901);
nor U11109 (N_11109,N_10850,N_10890);
nor U11110 (N_11110,N_10895,N_10883);
nor U11111 (N_11111,N_10789,N_10999);
and U11112 (N_11112,N_10825,N_10851);
or U11113 (N_11113,N_10909,N_10966);
or U11114 (N_11114,N_10841,N_10820);
or U11115 (N_11115,N_10997,N_10802);
and U11116 (N_11116,N_10962,N_10951);
or U11117 (N_11117,N_10967,N_10860);
nand U11118 (N_11118,N_10764,N_10815);
nand U11119 (N_11119,N_10956,N_10910);
nand U11120 (N_11120,N_10932,N_10854);
nand U11121 (N_11121,N_10955,N_10814);
and U11122 (N_11122,N_10952,N_10885);
or U11123 (N_11123,N_10980,N_10803);
nand U11124 (N_11124,N_10974,N_10935);
or U11125 (N_11125,N_10839,N_10807);
or U11126 (N_11126,N_10972,N_10777);
or U11127 (N_11127,N_10910,N_10759);
nand U11128 (N_11128,N_10857,N_10885);
and U11129 (N_11129,N_10752,N_10926);
or U11130 (N_11130,N_10837,N_10960);
and U11131 (N_11131,N_10818,N_10820);
nand U11132 (N_11132,N_10934,N_10804);
nand U11133 (N_11133,N_10802,N_10999);
and U11134 (N_11134,N_10900,N_10966);
nor U11135 (N_11135,N_10869,N_10958);
nor U11136 (N_11136,N_10884,N_10923);
nor U11137 (N_11137,N_10797,N_10945);
nand U11138 (N_11138,N_10931,N_10987);
and U11139 (N_11139,N_10878,N_10973);
and U11140 (N_11140,N_10761,N_10752);
nand U11141 (N_11141,N_10755,N_10883);
and U11142 (N_11142,N_10756,N_10818);
nand U11143 (N_11143,N_10918,N_10792);
nand U11144 (N_11144,N_10871,N_10907);
nand U11145 (N_11145,N_10955,N_10795);
nand U11146 (N_11146,N_10822,N_10833);
nand U11147 (N_11147,N_10892,N_10887);
nor U11148 (N_11148,N_10957,N_10764);
nor U11149 (N_11149,N_10885,N_10946);
and U11150 (N_11150,N_10815,N_10951);
and U11151 (N_11151,N_10752,N_10956);
and U11152 (N_11152,N_10895,N_10751);
and U11153 (N_11153,N_10990,N_10917);
and U11154 (N_11154,N_10995,N_10807);
nor U11155 (N_11155,N_10936,N_10994);
or U11156 (N_11156,N_10839,N_10895);
nand U11157 (N_11157,N_10959,N_10899);
nor U11158 (N_11158,N_10846,N_10764);
or U11159 (N_11159,N_10857,N_10809);
nor U11160 (N_11160,N_10759,N_10882);
or U11161 (N_11161,N_10884,N_10842);
or U11162 (N_11162,N_10928,N_10862);
nor U11163 (N_11163,N_10955,N_10970);
nand U11164 (N_11164,N_10840,N_10918);
nand U11165 (N_11165,N_10813,N_10898);
nor U11166 (N_11166,N_10767,N_10890);
nand U11167 (N_11167,N_10774,N_10859);
and U11168 (N_11168,N_10754,N_10963);
nand U11169 (N_11169,N_10950,N_10930);
and U11170 (N_11170,N_10804,N_10985);
nand U11171 (N_11171,N_10862,N_10770);
nand U11172 (N_11172,N_10778,N_10887);
nand U11173 (N_11173,N_10846,N_10947);
or U11174 (N_11174,N_10831,N_10812);
nand U11175 (N_11175,N_10939,N_10835);
and U11176 (N_11176,N_10908,N_10858);
nor U11177 (N_11177,N_10836,N_10916);
nor U11178 (N_11178,N_10922,N_10855);
nand U11179 (N_11179,N_10864,N_10890);
nand U11180 (N_11180,N_10941,N_10862);
and U11181 (N_11181,N_10881,N_10793);
nand U11182 (N_11182,N_10904,N_10891);
and U11183 (N_11183,N_10984,N_10848);
nor U11184 (N_11184,N_10965,N_10802);
or U11185 (N_11185,N_10922,N_10850);
nor U11186 (N_11186,N_10942,N_10887);
or U11187 (N_11187,N_10952,N_10908);
nor U11188 (N_11188,N_10991,N_10984);
or U11189 (N_11189,N_10967,N_10767);
or U11190 (N_11190,N_10958,N_10994);
nand U11191 (N_11191,N_10886,N_10856);
or U11192 (N_11192,N_10813,N_10775);
nand U11193 (N_11193,N_10810,N_10941);
and U11194 (N_11194,N_10866,N_10823);
and U11195 (N_11195,N_10854,N_10909);
nor U11196 (N_11196,N_10757,N_10957);
or U11197 (N_11197,N_10808,N_10878);
or U11198 (N_11198,N_10751,N_10750);
or U11199 (N_11199,N_10964,N_10797);
and U11200 (N_11200,N_10871,N_10857);
or U11201 (N_11201,N_10914,N_10975);
nand U11202 (N_11202,N_10831,N_10931);
or U11203 (N_11203,N_10959,N_10753);
or U11204 (N_11204,N_10867,N_10930);
and U11205 (N_11205,N_10841,N_10770);
nand U11206 (N_11206,N_10782,N_10986);
xor U11207 (N_11207,N_10843,N_10918);
and U11208 (N_11208,N_10855,N_10971);
nor U11209 (N_11209,N_10903,N_10867);
and U11210 (N_11210,N_10890,N_10787);
nor U11211 (N_11211,N_10898,N_10930);
xor U11212 (N_11212,N_10828,N_10756);
or U11213 (N_11213,N_10910,N_10999);
or U11214 (N_11214,N_10769,N_10942);
nor U11215 (N_11215,N_10757,N_10838);
nand U11216 (N_11216,N_10989,N_10977);
and U11217 (N_11217,N_10938,N_10865);
and U11218 (N_11218,N_10778,N_10901);
or U11219 (N_11219,N_10809,N_10901);
nor U11220 (N_11220,N_10946,N_10872);
or U11221 (N_11221,N_10789,N_10821);
nand U11222 (N_11222,N_10953,N_10833);
nand U11223 (N_11223,N_10947,N_10913);
and U11224 (N_11224,N_10888,N_10833);
nor U11225 (N_11225,N_10794,N_10879);
or U11226 (N_11226,N_10786,N_10779);
nand U11227 (N_11227,N_10988,N_10923);
nand U11228 (N_11228,N_10775,N_10911);
nand U11229 (N_11229,N_10902,N_10852);
nand U11230 (N_11230,N_10768,N_10909);
nand U11231 (N_11231,N_10935,N_10896);
and U11232 (N_11232,N_10951,N_10769);
nor U11233 (N_11233,N_10935,N_10899);
or U11234 (N_11234,N_10935,N_10772);
or U11235 (N_11235,N_10848,N_10770);
nand U11236 (N_11236,N_10932,N_10943);
nand U11237 (N_11237,N_10769,N_10768);
nor U11238 (N_11238,N_10880,N_10764);
nor U11239 (N_11239,N_10846,N_10984);
and U11240 (N_11240,N_10778,N_10859);
or U11241 (N_11241,N_10758,N_10755);
nand U11242 (N_11242,N_10756,N_10792);
or U11243 (N_11243,N_10834,N_10830);
nand U11244 (N_11244,N_10863,N_10908);
nand U11245 (N_11245,N_10877,N_10939);
nor U11246 (N_11246,N_10952,N_10977);
nor U11247 (N_11247,N_10991,N_10983);
nor U11248 (N_11248,N_10788,N_10913);
nor U11249 (N_11249,N_10831,N_10844);
nand U11250 (N_11250,N_11235,N_11056);
or U11251 (N_11251,N_11188,N_11106);
nand U11252 (N_11252,N_11226,N_11040);
or U11253 (N_11253,N_11086,N_11103);
nor U11254 (N_11254,N_11098,N_11121);
or U11255 (N_11255,N_11233,N_11085);
or U11256 (N_11256,N_11060,N_11037);
or U11257 (N_11257,N_11109,N_11142);
and U11258 (N_11258,N_11127,N_11216);
and U11259 (N_11259,N_11072,N_11028);
and U11260 (N_11260,N_11027,N_11120);
nor U11261 (N_11261,N_11137,N_11044);
nor U11262 (N_11262,N_11001,N_11196);
and U11263 (N_11263,N_11140,N_11202);
and U11264 (N_11264,N_11064,N_11069);
and U11265 (N_11265,N_11249,N_11020);
nor U11266 (N_11266,N_11143,N_11110);
nand U11267 (N_11267,N_11212,N_11095);
nor U11268 (N_11268,N_11013,N_11186);
nor U11269 (N_11269,N_11192,N_11038);
or U11270 (N_11270,N_11088,N_11003);
and U11271 (N_11271,N_11172,N_11117);
or U11272 (N_11272,N_11146,N_11042);
or U11273 (N_11273,N_11070,N_11191);
nor U11274 (N_11274,N_11144,N_11234);
and U11275 (N_11275,N_11023,N_11148);
or U11276 (N_11276,N_11031,N_11141);
nand U11277 (N_11277,N_11217,N_11162);
nor U11278 (N_11278,N_11169,N_11091);
nand U11279 (N_11279,N_11006,N_11164);
nor U11280 (N_11280,N_11017,N_11077);
xor U11281 (N_11281,N_11225,N_11094);
nor U11282 (N_11282,N_11016,N_11168);
nand U11283 (N_11283,N_11223,N_11171);
nand U11284 (N_11284,N_11097,N_11247);
and U11285 (N_11285,N_11151,N_11015);
and U11286 (N_11286,N_11182,N_11167);
or U11287 (N_11287,N_11032,N_11124);
or U11288 (N_11288,N_11068,N_11089);
and U11289 (N_11289,N_11238,N_11000);
or U11290 (N_11290,N_11046,N_11065);
nor U11291 (N_11291,N_11149,N_11138);
and U11292 (N_11292,N_11232,N_11227);
and U11293 (N_11293,N_11105,N_11183);
and U11294 (N_11294,N_11035,N_11011);
nor U11295 (N_11295,N_11055,N_11067);
nor U11296 (N_11296,N_11054,N_11123);
and U11297 (N_11297,N_11215,N_11156);
nor U11298 (N_11298,N_11181,N_11236);
nor U11299 (N_11299,N_11136,N_11048);
nor U11300 (N_11300,N_11066,N_11047);
or U11301 (N_11301,N_11240,N_11132);
nand U11302 (N_11302,N_11050,N_11159);
nor U11303 (N_11303,N_11173,N_11203);
xor U11304 (N_11304,N_11062,N_11214);
or U11305 (N_11305,N_11099,N_11219);
nand U11306 (N_11306,N_11152,N_11150);
and U11307 (N_11307,N_11176,N_11153);
nor U11308 (N_11308,N_11083,N_11134);
and U11309 (N_11309,N_11177,N_11058);
and U11310 (N_11310,N_11102,N_11005);
nor U11311 (N_11311,N_11248,N_11087);
or U11312 (N_11312,N_11145,N_11084);
nand U11313 (N_11313,N_11170,N_11108);
nand U11314 (N_11314,N_11004,N_11116);
nand U11315 (N_11315,N_11185,N_11113);
and U11316 (N_11316,N_11245,N_11158);
and U11317 (N_11317,N_11074,N_11201);
nor U11318 (N_11318,N_11049,N_11241);
nor U11319 (N_11319,N_11043,N_11165);
or U11320 (N_11320,N_11024,N_11114);
or U11321 (N_11321,N_11200,N_11092);
nand U11322 (N_11322,N_11107,N_11130);
nand U11323 (N_11323,N_11204,N_11218);
or U11324 (N_11324,N_11075,N_11008);
or U11325 (N_11325,N_11051,N_11039);
nor U11326 (N_11326,N_11007,N_11100);
nor U11327 (N_11327,N_11157,N_11045);
and U11328 (N_11328,N_11209,N_11224);
nor U11329 (N_11329,N_11071,N_11199);
and U11330 (N_11330,N_11229,N_11211);
and U11331 (N_11331,N_11187,N_11115);
or U11332 (N_11332,N_11198,N_11010);
and U11333 (N_11333,N_11222,N_11228);
nand U11334 (N_11334,N_11026,N_11025);
nand U11335 (N_11335,N_11154,N_11205);
or U11336 (N_11336,N_11161,N_11128);
nand U11337 (N_11337,N_11021,N_11030);
nor U11338 (N_11338,N_11053,N_11189);
nor U11339 (N_11339,N_11213,N_11081);
and U11340 (N_11340,N_11009,N_11197);
or U11341 (N_11341,N_11194,N_11131);
and U11342 (N_11342,N_11111,N_11082);
and U11343 (N_11343,N_11119,N_11160);
nor U11344 (N_11344,N_11125,N_11220);
nor U11345 (N_11345,N_11052,N_11029);
or U11346 (N_11346,N_11244,N_11175);
nand U11347 (N_11347,N_11112,N_11133);
nand U11348 (N_11348,N_11206,N_11193);
or U11349 (N_11349,N_11155,N_11178);
nor U11350 (N_11350,N_11080,N_11118);
and U11351 (N_11351,N_11012,N_11014);
nand U11352 (N_11352,N_11139,N_11179);
nand U11353 (N_11353,N_11073,N_11104);
or U11354 (N_11354,N_11090,N_11122);
or U11355 (N_11355,N_11231,N_11079);
and U11356 (N_11356,N_11126,N_11208);
or U11357 (N_11357,N_11166,N_11034);
or U11358 (N_11358,N_11061,N_11174);
nand U11359 (N_11359,N_11230,N_11018);
nand U11360 (N_11360,N_11033,N_11147);
or U11361 (N_11361,N_11237,N_11246);
or U11362 (N_11362,N_11190,N_11184);
or U11363 (N_11363,N_11243,N_11207);
nor U11364 (N_11364,N_11221,N_11057);
or U11365 (N_11365,N_11135,N_11242);
or U11366 (N_11366,N_11180,N_11195);
or U11367 (N_11367,N_11210,N_11002);
or U11368 (N_11368,N_11078,N_11129);
or U11369 (N_11369,N_11096,N_11063);
or U11370 (N_11370,N_11041,N_11163);
nand U11371 (N_11371,N_11059,N_11093);
or U11372 (N_11372,N_11022,N_11101);
or U11373 (N_11373,N_11076,N_11019);
or U11374 (N_11374,N_11239,N_11036);
and U11375 (N_11375,N_11161,N_11021);
and U11376 (N_11376,N_11112,N_11240);
and U11377 (N_11377,N_11243,N_11022);
and U11378 (N_11378,N_11229,N_11091);
and U11379 (N_11379,N_11209,N_11244);
and U11380 (N_11380,N_11053,N_11157);
or U11381 (N_11381,N_11001,N_11192);
nand U11382 (N_11382,N_11009,N_11156);
and U11383 (N_11383,N_11055,N_11128);
and U11384 (N_11384,N_11138,N_11178);
nor U11385 (N_11385,N_11195,N_11060);
and U11386 (N_11386,N_11049,N_11208);
and U11387 (N_11387,N_11176,N_11075);
or U11388 (N_11388,N_11107,N_11234);
and U11389 (N_11389,N_11168,N_11205);
or U11390 (N_11390,N_11096,N_11247);
nand U11391 (N_11391,N_11118,N_11206);
nor U11392 (N_11392,N_11046,N_11042);
nor U11393 (N_11393,N_11029,N_11231);
nor U11394 (N_11394,N_11011,N_11038);
nand U11395 (N_11395,N_11108,N_11195);
and U11396 (N_11396,N_11098,N_11046);
nor U11397 (N_11397,N_11170,N_11058);
or U11398 (N_11398,N_11233,N_11205);
and U11399 (N_11399,N_11193,N_11045);
nand U11400 (N_11400,N_11086,N_11101);
nor U11401 (N_11401,N_11012,N_11170);
and U11402 (N_11402,N_11061,N_11014);
and U11403 (N_11403,N_11069,N_11066);
nand U11404 (N_11404,N_11247,N_11138);
and U11405 (N_11405,N_11165,N_11212);
or U11406 (N_11406,N_11220,N_11131);
xor U11407 (N_11407,N_11031,N_11203);
or U11408 (N_11408,N_11228,N_11044);
nand U11409 (N_11409,N_11227,N_11193);
nand U11410 (N_11410,N_11204,N_11092);
nand U11411 (N_11411,N_11232,N_11163);
nand U11412 (N_11412,N_11105,N_11094);
nor U11413 (N_11413,N_11026,N_11246);
and U11414 (N_11414,N_11177,N_11088);
nand U11415 (N_11415,N_11090,N_11185);
and U11416 (N_11416,N_11072,N_11088);
or U11417 (N_11417,N_11025,N_11190);
nor U11418 (N_11418,N_11239,N_11099);
or U11419 (N_11419,N_11230,N_11086);
nor U11420 (N_11420,N_11059,N_11143);
nand U11421 (N_11421,N_11053,N_11070);
and U11422 (N_11422,N_11042,N_11161);
nor U11423 (N_11423,N_11000,N_11176);
nor U11424 (N_11424,N_11024,N_11001);
or U11425 (N_11425,N_11036,N_11204);
nor U11426 (N_11426,N_11198,N_11146);
nor U11427 (N_11427,N_11172,N_11108);
and U11428 (N_11428,N_11115,N_11178);
nor U11429 (N_11429,N_11166,N_11100);
or U11430 (N_11430,N_11192,N_11214);
nand U11431 (N_11431,N_11041,N_11130);
or U11432 (N_11432,N_11095,N_11246);
nor U11433 (N_11433,N_11024,N_11013);
nor U11434 (N_11434,N_11193,N_11106);
nand U11435 (N_11435,N_11144,N_11032);
nand U11436 (N_11436,N_11034,N_11051);
nand U11437 (N_11437,N_11019,N_11219);
nor U11438 (N_11438,N_11170,N_11038);
nand U11439 (N_11439,N_11078,N_11091);
or U11440 (N_11440,N_11165,N_11054);
or U11441 (N_11441,N_11082,N_11094);
nor U11442 (N_11442,N_11140,N_11000);
and U11443 (N_11443,N_11173,N_11023);
nand U11444 (N_11444,N_11100,N_11044);
or U11445 (N_11445,N_11106,N_11101);
or U11446 (N_11446,N_11022,N_11196);
and U11447 (N_11447,N_11056,N_11041);
or U11448 (N_11448,N_11069,N_11098);
and U11449 (N_11449,N_11126,N_11052);
and U11450 (N_11450,N_11241,N_11116);
nor U11451 (N_11451,N_11035,N_11079);
nand U11452 (N_11452,N_11213,N_11154);
nand U11453 (N_11453,N_11012,N_11217);
and U11454 (N_11454,N_11219,N_11129);
and U11455 (N_11455,N_11085,N_11098);
nand U11456 (N_11456,N_11120,N_11156);
or U11457 (N_11457,N_11015,N_11091);
and U11458 (N_11458,N_11127,N_11037);
nor U11459 (N_11459,N_11006,N_11063);
and U11460 (N_11460,N_11021,N_11212);
nand U11461 (N_11461,N_11125,N_11210);
or U11462 (N_11462,N_11087,N_11081);
and U11463 (N_11463,N_11023,N_11137);
nand U11464 (N_11464,N_11187,N_11047);
nand U11465 (N_11465,N_11184,N_11032);
or U11466 (N_11466,N_11208,N_11090);
or U11467 (N_11467,N_11132,N_11136);
or U11468 (N_11468,N_11051,N_11093);
nor U11469 (N_11469,N_11190,N_11051);
nand U11470 (N_11470,N_11017,N_11146);
and U11471 (N_11471,N_11074,N_11228);
or U11472 (N_11472,N_11109,N_11242);
nor U11473 (N_11473,N_11053,N_11042);
and U11474 (N_11474,N_11157,N_11058);
nor U11475 (N_11475,N_11077,N_11054);
and U11476 (N_11476,N_11100,N_11187);
or U11477 (N_11477,N_11131,N_11187);
nor U11478 (N_11478,N_11108,N_11129);
or U11479 (N_11479,N_11035,N_11051);
or U11480 (N_11480,N_11001,N_11098);
or U11481 (N_11481,N_11096,N_11020);
or U11482 (N_11482,N_11066,N_11045);
nor U11483 (N_11483,N_11231,N_11102);
or U11484 (N_11484,N_11034,N_11138);
and U11485 (N_11485,N_11176,N_11236);
nand U11486 (N_11486,N_11234,N_11079);
or U11487 (N_11487,N_11216,N_11116);
nand U11488 (N_11488,N_11163,N_11201);
and U11489 (N_11489,N_11242,N_11164);
or U11490 (N_11490,N_11244,N_11043);
nor U11491 (N_11491,N_11066,N_11247);
nor U11492 (N_11492,N_11238,N_11110);
and U11493 (N_11493,N_11030,N_11062);
nor U11494 (N_11494,N_11003,N_11011);
nor U11495 (N_11495,N_11208,N_11018);
or U11496 (N_11496,N_11047,N_11125);
or U11497 (N_11497,N_11162,N_11197);
and U11498 (N_11498,N_11009,N_11050);
nand U11499 (N_11499,N_11247,N_11225);
and U11500 (N_11500,N_11266,N_11378);
nor U11501 (N_11501,N_11317,N_11308);
nand U11502 (N_11502,N_11343,N_11442);
nand U11503 (N_11503,N_11283,N_11480);
nor U11504 (N_11504,N_11484,N_11334);
nand U11505 (N_11505,N_11447,N_11417);
nand U11506 (N_11506,N_11454,N_11420);
nand U11507 (N_11507,N_11279,N_11367);
nor U11508 (N_11508,N_11281,N_11310);
and U11509 (N_11509,N_11290,N_11437);
nor U11510 (N_11510,N_11315,N_11455);
or U11511 (N_11511,N_11405,N_11320);
and U11512 (N_11512,N_11386,N_11295);
or U11513 (N_11513,N_11297,N_11460);
nand U11514 (N_11514,N_11493,N_11462);
nor U11515 (N_11515,N_11273,N_11394);
and U11516 (N_11516,N_11381,N_11424);
or U11517 (N_11517,N_11401,N_11443);
and U11518 (N_11518,N_11348,N_11285);
nor U11519 (N_11519,N_11411,N_11450);
nand U11520 (N_11520,N_11483,N_11364);
xnor U11521 (N_11521,N_11339,N_11467);
nand U11522 (N_11522,N_11444,N_11469);
and U11523 (N_11523,N_11413,N_11466);
nor U11524 (N_11524,N_11250,N_11313);
and U11525 (N_11525,N_11341,N_11457);
nor U11526 (N_11526,N_11287,N_11270);
or U11527 (N_11527,N_11468,N_11463);
nor U11528 (N_11528,N_11387,N_11464);
or U11529 (N_11529,N_11395,N_11358);
and U11530 (N_11530,N_11421,N_11372);
nor U11531 (N_11531,N_11402,N_11436);
nand U11532 (N_11532,N_11403,N_11440);
nand U11533 (N_11533,N_11361,N_11498);
or U11534 (N_11534,N_11471,N_11353);
nor U11535 (N_11535,N_11311,N_11268);
nor U11536 (N_11536,N_11423,N_11300);
nor U11537 (N_11537,N_11446,N_11298);
nor U11538 (N_11538,N_11292,N_11370);
nand U11539 (N_11539,N_11330,N_11408);
or U11540 (N_11540,N_11284,N_11289);
nor U11541 (N_11541,N_11333,N_11303);
nor U11542 (N_11542,N_11261,N_11346);
and U11543 (N_11543,N_11384,N_11276);
and U11544 (N_11544,N_11286,N_11404);
or U11545 (N_11545,N_11355,N_11301);
nor U11546 (N_11546,N_11258,N_11280);
or U11547 (N_11547,N_11352,N_11407);
nand U11548 (N_11548,N_11327,N_11374);
nor U11549 (N_11549,N_11495,N_11337);
nand U11550 (N_11550,N_11269,N_11336);
nand U11551 (N_11551,N_11312,N_11487);
nand U11552 (N_11552,N_11377,N_11326);
nand U11553 (N_11553,N_11351,N_11476);
or U11554 (N_11554,N_11475,N_11438);
nor U11555 (N_11555,N_11272,N_11329);
xnor U11556 (N_11556,N_11251,N_11309);
and U11557 (N_11557,N_11415,N_11492);
or U11558 (N_11558,N_11332,N_11445);
or U11559 (N_11559,N_11429,N_11485);
nand U11560 (N_11560,N_11252,N_11254);
nor U11561 (N_11561,N_11465,N_11359);
nand U11562 (N_11562,N_11322,N_11418);
and U11563 (N_11563,N_11426,N_11323);
nand U11564 (N_11564,N_11388,N_11452);
nand U11565 (N_11565,N_11274,N_11441);
and U11566 (N_11566,N_11393,N_11306);
nand U11567 (N_11567,N_11494,N_11419);
or U11568 (N_11568,N_11479,N_11390);
or U11569 (N_11569,N_11499,N_11344);
and U11570 (N_11570,N_11391,N_11294);
nand U11571 (N_11571,N_11319,N_11253);
or U11572 (N_11572,N_11365,N_11278);
or U11573 (N_11573,N_11449,N_11347);
and U11574 (N_11574,N_11356,N_11324);
and U11575 (N_11575,N_11360,N_11260);
nand U11576 (N_11576,N_11321,N_11304);
nor U11577 (N_11577,N_11428,N_11345);
and U11578 (N_11578,N_11357,N_11267);
nor U11579 (N_11579,N_11262,N_11488);
nand U11580 (N_11580,N_11265,N_11416);
and U11581 (N_11581,N_11383,N_11368);
nor U11582 (N_11582,N_11427,N_11433);
nand U11583 (N_11583,N_11482,N_11496);
or U11584 (N_11584,N_11382,N_11461);
nor U11585 (N_11585,N_11422,N_11293);
nand U11586 (N_11586,N_11430,N_11296);
nand U11587 (N_11587,N_11439,N_11473);
and U11588 (N_11588,N_11314,N_11414);
or U11589 (N_11589,N_11478,N_11328);
nor U11590 (N_11590,N_11456,N_11481);
or U11591 (N_11591,N_11256,N_11335);
and U11592 (N_11592,N_11331,N_11435);
and U11593 (N_11593,N_11373,N_11474);
nor U11594 (N_11594,N_11362,N_11472);
nor U11595 (N_11595,N_11263,N_11257);
nor U11596 (N_11596,N_11397,N_11318);
and U11597 (N_11597,N_11282,N_11369);
nand U11598 (N_11598,N_11380,N_11307);
or U11599 (N_11599,N_11486,N_11410);
nand U11600 (N_11600,N_11354,N_11259);
or U11601 (N_11601,N_11271,N_11490);
nand U11602 (N_11602,N_11470,N_11448);
nand U11603 (N_11603,N_11491,N_11477);
and U11604 (N_11604,N_11451,N_11350);
or U11605 (N_11605,N_11376,N_11305);
nor U11606 (N_11606,N_11363,N_11316);
nand U11607 (N_11607,N_11431,N_11325);
nor U11608 (N_11608,N_11497,N_11375);
nor U11609 (N_11609,N_11398,N_11338);
or U11610 (N_11610,N_11389,N_11288);
and U11611 (N_11611,N_11371,N_11291);
nand U11612 (N_11612,N_11406,N_11264);
nand U11613 (N_11613,N_11453,N_11255);
nand U11614 (N_11614,N_11412,N_11349);
nor U11615 (N_11615,N_11277,N_11459);
and U11616 (N_11616,N_11400,N_11489);
nand U11617 (N_11617,N_11302,N_11379);
nor U11618 (N_11618,N_11409,N_11432);
and U11619 (N_11619,N_11366,N_11385);
nand U11620 (N_11620,N_11425,N_11275);
nand U11621 (N_11621,N_11342,N_11396);
nand U11622 (N_11622,N_11340,N_11399);
and U11623 (N_11623,N_11392,N_11434);
nor U11624 (N_11624,N_11458,N_11299);
nand U11625 (N_11625,N_11448,N_11432);
nor U11626 (N_11626,N_11428,N_11471);
and U11627 (N_11627,N_11409,N_11379);
or U11628 (N_11628,N_11377,N_11430);
or U11629 (N_11629,N_11486,N_11419);
nor U11630 (N_11630,N_11424,N_11437);
or U11631 (N_11631,N_11447,N_11406);
nand U11632 (N_11632,N_11429,N_11350);
nand U11633 (N_11633,N_11296,N_11498);
and U11634 (N_11634,N_11490,N_11357);
nor U11635 (N_11635,N_11488,N_11254);
nor U11636 (N_11636,N_11472,N_11379);
and U11637 (N_11637,N_11329,N_11355);
and U11638 (N_11638,N_11279,N_11479);
and U11639 (N_11639,N_11395,N_11322);
and U11640 (N_11640,N_11406,N_11395);
and U11641 (N_11641,N_11360,N_11263);
or U11642 (N_11642,N_11262,N_11491);
and U11643 (N_11643,N_11435,N_11433);
nand U11644 (N_11644,N_11482,N_11438);
or U11645 (N_11645,N_11315,N_11297);
nand U11646 (N_11646,N_11278,N_11260);
and U11647 (N_11647,N_11492,N_11377);
nor U11648 (N_11648,N_11442,N_11474);
and U11649 (N_11649,N_11332,N_11314);
nor U11650 (N_11650,N_11446,N_11337);
nor U11651 (N_11651,N_11257,N_11293);
nand U11652 (N_11652,N_11401,N_11431);
and U11653 (N_11653,N_11408,N_11380);
and U11654 (N_11654,N_11339,N_11337);
or U11655 (N_11655,N_11480,N_11365);
nand U11656 (N_11656,N_11432,N_11414);
or U11657 (N_11657,N_11351,N_11337);
and U11658 (N_11658,N_11300,N_11484);
nor U11659 (N_11659,N_11399,N_11289);
or U11660 (N_11660,N_11394,N_11424);
nand U11661 (N_11661,N_11292,N_11456);
and U11662 (N_11662,N_11401,N_11384);
and U11663 (N_11663,N_11371,N_11377);
or U11664 (N_11664,N_11351,N_11344);
nand U11665 (N_11665,N_11299,N_11359);
nand U11666 (N_11666,N_11371,N_11335);
nor U11667 (N_11667,N_11399,N_11421);
nand U11668 (N_11668,N_11497,N_11261);
nor U11669 (N_11669,N_11339,N_11366);
and U11670 (N_11670,N_11431,N_11413);
and U11671 (N_11671,N_11362,N_11400);
nor U11672 (N_11672,N_11273,N_11270);
nor U11673 (N_11673,N_11351,N_11310);
or U11674 (N_11674,N_11487,N_11285);
or U11675 (N_11675,N_11290,N_11250);
and U11676 (N_11676,N_11297,N_11436);
or U11677 (N_11677,N_11398,N_11298);
or U11678 (N_11678,N_11360,N_11477);
nand U11679 (N_11679,N_11337,N_11342);
nand U11680 (N_11680,N_11385,N_11314);
nand U11681 (N_11681,N_11315,N_11343);
nor U11682 (N_11682,N_11389,N_11279);
nand U11683 (N_11683,N_11431,N_11275);
and U11684 (N_11684,N_11419,N_11357);
or U11685 (N_11685,N_11311,N_11274);
and U11686 (N_11686,N_11292,N_11290);
nor U11687 (N_11687,N_11327,N_11367);
or U11688 (N_11688,N_11475,N_11288);
or U11689 (N_11689,N_11343,N_11451);
nor U11690 (N_11690,N_11363,N_11366);
or U11691 (N_11691,N_11419,N_11299);
nand U11692 (N_11692,N_11369,N_11280);
or U11693 (N_11693,N_11419,N_11408);
and U11694 (N_11694,N_11429,N_11472);
or U11695 (N_11695,N_11412,N_11327);
or U11696 (N_11696,N_11390,N_11303);
nand U11697 (N_11697,N_11355,N_11406);
nand U11698 (N_11698,N_11344,N_11390);
and U11699 (N_11699,N_11463,N_11374);
nand U11700 (N_11700,N_11329,N_11274);
or U11701 (N_11701,N_11310,N_11416);
nand U11702 (N_11702,N_11449,N_11483);
and U11703 (N_11703,N_11360,N_11410);
and U11704 (N_11704,N_11382,N_11467);
nor U11705 (N_11705,N_11461,N_11423);
nor U11706 (N_11706,N_11347,N_11466);
or U11707 (N_11707,N_11370,N_11431);
nor U11708 (N_11708,N_11418,N_11401);
or U11709 (N_11709,N_11255,N_11487);
xnor U11710 (N_11710,N_11278,N_11327);
nand U11711 (N_11711,N_11362,N_11422);
nor U11712 (N_11712,N_11469,N_11483);
nand U11713 (N_11713,N_11309,N_11310);
nand U11714 (N_11714,N_11431,N_11389);
or U11715 (N_11715,N_11269,N_11287);
and U11716 (N_11716,N_11331,N_11370);
nor U11717 (N_11717,N_11267,N_11339);
nand U11718 (N_11718,N_11413,N_11370);
xnor U11719 (N_11719,N_11440,N_11317);
nand U11720 (N_11720,N_11439,N_11399);
and U11721 (N_11721,N_11421,N_11280);
or U11722 (N_11722,N_11333,N_11330);
and U11723 (N_11723,N_11317,N_11385);
nor U11724 (N_11724,N_11285,N_11330);
and U11725 (N_11725,N_11256,N_11321);
and U11726 (N_11726,N_11364,N_11270);
and U11727 (N_11727,N_11298,N_11254);
nand U11728 (N_11728,N_11441,N_11311);
nand U11729 (N_11729,N_11401,N_11397);
or U11730 (N_11730,N_11488,N_11299);
and U11731 (N_11731,N_11389,N_11299);
nand U11732 (N_11732,N_11329,N_11357);
nor U11733 (N_11733,N_11325,N_11282);
and U11734 (N_11734,N_11278,N_11434);
nor U11735 (N_11735,N_11322,N_11384);
and U11736 (N_11736,N_11386,N_11412);
nor U11737 (N_11737,N_11254,N_11335);
or U11738 (N_11738,N_11378,N_11389);
and U11739 (N_11739,N_11403,N_11466);
or U11740 (N_11740,N_11444,N_11378);
or U11741 (N_11741,N_11261,N_11441);
or U11742 (N_11742,N_11485,N_11382);
nor U11743 (N_11743,N_11366,N_11318);
nand U11744 (N_11744,N_11374,N_11299);
and U11745 (N_11745,N_11400,N_11421);
nand U11746 (N_11746,N_11498,N_11292);
nand U11747 (N_11747,N_11482,N_11271);
nor U11748 (N_11748,N_11323,N_11354);
or U11749 (N_11749,N_11400,N_11457);
nor U11750 (N_11750,N_11722,N_11721);
and U11751 (N_11751,N_11515,N_11577);
and U11752 (N_11752,N_11537,N_11669);
nand U11753 (N_11753,N_11518,N_11731);
nand U11754 (N_11754,N_11663,N_11573);
and U11755 (N_11755,N_11733,N_11605);
xnor U11756 (N_11756,N_11588,N_11625);
nor U11757 (N_11757,N_11504,N_11640);
nand U11758 (N_11758,N_11735,N_11525);
or U11759 (N_11759,N_11520,N_11576);
nand U11760 (N_11760,N_11665,N_11559);
and U11761 (N_11761,N_11614,N_11709);
nand U11762 (N_11762,N_11700,N_11686);
or U11763 (N_11763,N_11681,N_11521);
nand U11764 (N_11764,N_11601,N_11684);
nor U11765 (N_11765,N_11547,N_11553);
nor U11766 (N_11766,N_11581,N_11740);
nand U11767 (N_11767,N_11703,N_11526);
and U11768 (N_11768,N_11685,N_11619);
nor U11769 (N_11769,N_11742,N_11666);
nor U11770 (N_11770,N_11594,N_11710);
or U11771 (N_11771,N_11678,N_11551);
nand U11772 (N_11772,N_11599,N_11734);
nor U11773 (N_11773,N_11568,N_11554);
nor U11774 (N_11774,N_11562,N_11720);
or U11775 (N_11775,N_11566,N_11602);
and U11776 (N_11776,N_11749,N_11745);
or U11777 (N_11777,N_11719,N_11657);
nor U11778 (N_11778,N_11536,N_11617);
nor U11779 (N_11779,N_11592,N_11743);
nand U11780 (N_11780,N_11716,N_11688);
or U11781 (N_11781,N_11560,N_11634);
and U11782 (N_11782,N_11699,N_11712);
or U11783 (N_11783,N_11590,N_11694);
or U11784 (N_11784,N_11682,N_11642);
and U11785 (N_11785,N_11607,N_11557);
or U11786 (N_11786,N_11546,N_11654);
nand U11787 (N_11787,N_11571,N_11664);
or U11788 (N_11788,N_11725,N_11500);
xnor U11789 (N_11789,N_11628,N_11556);
or U11790 (N_11790,N_11726,N_11652);
or U11791 (N_11791,N_11711,N_11727);
and U11792 (N_11792,N_11570,N_11639);
and U11793 (N_11793,N_11655,N_11502);
or U11794 (N_11794,N_11717,N_11693);
and U11795 (N_11795,N_11532,N_11616);
or U11796 (N_11796,N_11608,N_11680);
and U11797 (N_11797,N_11505,N_11552);
nor U11798 (N_11798,N_11569,N_11535);
nand U11799 (N_11799,N_11732,N_11512);
nand U11800 (N_11800,N_11503,N_11623);
or U11801 (N_11801,N_11530,N_11705);
nor U11802 (N_11802,N_11630,N_11656);
and U11803 (N_11803,N_11638,N_11741);
and U11804 (N_11804,N_11519,N_11713);
nor U11805 (N_11805,N_11683,N_11631);
and U11806 (N_11806,N_11689,N_11620);
or U11807 (N_11807,N_11615,N_11604);
nor U11808 (N_11808,N_11501,N_11645);
nand U11809 (N_11809,N_11544,N_11627);
nor U11810 (N_11810,N_11729,N_11509);
or U11811 (N_11811,N_11540,N_11578);
and U11812 (N_11812,N_11701,N_11609);
and U11813 (N_11813,N_11738,N_11648);
nor U11814 (N_11814,N_11548,N_11511);
nand U11815 (N_11815,N_11718,N_11730);
or U11816 (N_11816,N_11565,N_11633);
or U11817 (N_11817,N_11600,N_11517);
and U11818 (N_11818,N_11549,N_11618);
nor U11819 (N_11819,N_11651,N_11510);
nor U11820 (N_11820,N_11567,N_11507);
and U11821 (N_11821,N_11668,N_11690);
or U11822 (N_11822,N_11587,N_11583);
or U11823 (N_11823,N_11574,N_11555);
and U11824 (N_11824,N_11646,N_11586);
and U11825 (N_11825,N_11527,N_11637);
xnor U11826 (N_11826,N_11516,N_11533);
or U11827 (N_11827,N_11550,N_11653);
nor U11828 (N_11828,N_11675,N_11606);
nor U11829 (N_11829,N_11538,N_11528);
or U11830 (N_11830,N_11529,N_11674);
nand U11831 (N_11831,N_11728,N_11724);
nor U11832 (N_11832,N_11522,N_11695);
and U11833 (N_11833,N_11696,N_11621);
or U11834 (N_11834,N_11534,N_11589);
or U11835 (N_11835,N_11612,N_11622);
and U11836 (N_11836,N_11748,N_11692);
nand U11837 (N_11837,N_11603,N_11514);
nor U11838 (N_11838,N_11597,N_11659);
or U11839 (N_11839,N_11704,N_11658);
and U11840 (N_11840,N_11613,N_11593);
xnor U11841 (N_11841,N_11698,N_11611);
nor U11842 (N_11842,N_11708,N_11660);
or U11843 (N_11843,N_11596,N_11671);
nand U11844 (N_11844,N_11541,N_11723);
or U11845 (N_11845,N_11561,N_11673);
or U11846 (N_11846,N_11706,N_11575);
nand U11847 (N_11847,N_11524,N_11670);
or U11848 (N_11848,N_11580,N_11697);
nor U11849 (N_11849,N_11508,N_11513);
nor U11850 (N_11850,N_11636,N_11747);
nor U11851 (N_11851,N_11635,N_11545);
nand U11852 (N_11852,N_11629,N_11563);
or U11853 (N_11853,N_11595,N_11543);
nand U11854 (N_11854,N_11523,N_11715);
and U11855 (N_11855,N_11702,N_11641);
or U11856 (N_11856,N_11584,N_11624);
nor U11857 (N_11857,N_11676,N_11679);
or U11858 (N_11858,N_11632,N_11647);
and U11859 (N_11859,N_11506,N_11582);
nor U11860 (N_11860,N_11739,N_11585);
or U11861 (N_11861,N_11714,N_11542);
or U11862 (N_11862,N_11564,N_11649);
nor U11863 (N_11863,N_11610,N_11672);
nor U11864 (N_11864,N_11746,N_11667);
nand U11865 (N_11865,N_11591,N_11598);
nand U11866 (N_11866,N_11736,N_11572);
and U11867 (N_11867,N_11579,N_11744);
or U11868 (N_11868,N_11643,N_11687);
and U11869 (N_11869,N_11691,N_11539);
or U11870 (N_11870,N_11626,N_11644);
or U11871 (N_11871,N_11707,N_11650);
and U11872 (N_11872,N_11662,N_11677);
nand U11873 (N_11873,N_11737,N_11558);
nand U11874 (N_11874,N_11661,N_11531);
or U11875 (N_11875,N_11675,N_11510);
nor U11876 (N_11876,N_11728,N_11655);
xnor U11877 (N_11877,N_11721,N_11599);
nor U11878 (N_11878,N_11653,N_11533);
and U11879 (N_11879,N_11666,N_11649);
and U11880 (N_11880,N_11686,N_11691);
or U11881 (N_11881,N_11521,N_11700);
nor U11882 (N_11882,N_11646,N_11601);
nand U11883 (N_11883,N_11631,N_11620);
nand U11884 (N_11884,N_11601,N_11720);
and U11885 (N_11885,N_11546,N_11738);
nand U11886 (N_11886,N_11632,N_11566);
and U11887 (N_11887,N_11614,N_11524);
nand U11888 (N_11888,N_11542,N_11601);
or U11889 (N_11889,N_11524,N_11650);
or U11890 (N_11890,N_11648,N_11511);
or U11891 (N_11891,N_11504,N_11538);
nand U11892 (N_11892,N_11734,N_11501);
nor U11893 (N_11893,N_11745,N_11629);
nand U11894 (N_11894,N_11610,N_11695);
or U11895 (N_11895,N_11643,N_11650);
or U11896 (N_11896,N_11683,N_11538);
or U11897 (N_11897,N_11743,N_11666);
or U11898 (N_11898,N_11618,N_11732);
or U11899 (N_11899,N_11690,N_11736);
and U11900 (N_11900,N_11560,N_11506);
nor U11901 (N_11901,N_11626,N_11703);
nand U11902 (N_11902,N_11515,N_11597);
or U11903 (N_11903,N_11675,N_11699);
or U11904 (N_11904,N_11646,N_11597);
or U11905 (N_11905,N_11689,N_11632);
and U11906 (N_11906,N_11653,N_11561);
nand U11907 (N_11907,N_11681,N_11682);
or U11908 (N_11908,N_11502,N_11515);
nor U11909 (N_11909,N_11605,N_11525);
nor U11910 (N_11910,N_11720,N_11736);
nand U11911 (N_11911,N_11623,N_11510);
or U11912 (N_11912,N_11547,N_11627);
and U11913 (N_11913,N_11747,N_11638);
or U11914 (N_11914,N_11720,N_11600);
nand U11915 (N_11915,N_11577,N_11538);
nand U11916 (N_11916,N_11648,N_11506);
and U11917 (N_11917,N_11605,N_11671);
and U11918 (N_11918,N_11658,N_11503);
or U11919 (N_11919,N_11641,N_11516);
nor U11920 (N_11920,N_11551,N_11704);
nor U11921 (N_11921,N_11623,N_11749);
or U11922 (N_11922,N_11657,N_11619);
or U11923 (N_11923,N_11504,N_11586);
or U11924 (N_11924,N_11660,N_11625);
nor U11925 (N_11925,N_11647,N_11601);
and U11926 (N_11926,N_11659,N_11718);
or U11927 (N_11927,N_11613,N_11546);
nor U11928 (N_11928,N_11659,N_11695);
and U11929 (N_11929,N_11668,N_11615);
xnor U11930 (N_11930,N_11597,N_11513);
and U11931 (N_11931,N_11534,N_11615);
and U11932 (N_11932,N_11683,N_11741);
or U11933 (N_11933,N_11731,N_11503);
or U11934 (N_11934,N_11555,N_11580);
or U11935 (N_11935,N_11612,N_11627);
and U11936 (N_11936,N_11555,N_11619);
or U11937 (N_11937,N_11687,N_11523);
nor U11938 (N_11938,N_11714,N_11708);
nor U11939 (N_11939,N_11696,N_11637);
and U11940 (N_11940,N_11636,N_11608);
nor U11941 (N_11941,N_11562,N_11735);
nor U11942 (N_11942,N_11574,N_11588);
nand U11943 (N_11943,N_11578,N_11681);
and U11944 (N_11944,N_11585,N_11588);
nor U11945 (N_11945,N_11600,N_11686);
or U11946 (N_11946,N_11576,N_11515);
or U11947 (N_11947,N_11595,N_11502);
nor U11948 (N_11948,N_11618,N_11584);
and U11949 (N_11949,N_11688,N_11649);
nor U11950 (N_11950,N_11576,N_11743);
nor U11951 (N_11951,N_11613,N_11633);
and U11952 (N_11952,N_11598,N_11538);
nor U11953 (N_11953,N_11718,N_11635);
nor U11954 (N_11954,N_11681,N_11534);
nor U11955 (N_11955,N_11533,N_11515);
or U11956 (N_11956,N_11695,N_11615);
nand U11957 (N_11957,N_11578,N_11668);
nor U11958 (N_11958,N_11710,N_11528);
and U11959 (N_11959,N_11518,N_11568);
nand U11960 (N_11960,N_11694,N_11631);
and U11961 (N_11961,N_11740,N_11712);
nand U11962 (N_11962,N_11637,N_11599);
or U11963 (N_11963,N_11716,N_11574);
or U11964 (N_11964,N_11676,N_11727);
or U11965 (N_11965,N_11582,N_11540);
or U11966 (N_11966,N_11612,N_11722);
and U11967 (N_11967,N_11550,N_11614);
nor U11968 (N_11968,N_11688,N_11584);
or U11969 (N_11969,N_11643,N_11686);
nand U11970 (N_11970,N_11658,N_11544);
and U11971 (N_11971,N_11693,N_11724);
nand U11972 (N_11972,N_11503,N_11654);
nand U11973 (N_11973,N_11575,N_11748);
nand U11974 (N_11974,N_11731,N_11727);
nand U11975 (N_11975,N_11710,N_11537);
or U11976 (N_11976,N_11748,N_11722);
nand U11977 (N_11977,N_11696,N_11694);
and U11978 (N_11978,N_11554,N_11571);
or U11979 (N_11979,N_11747,N_11629);
nand U11980 (N_11980,N_11733,N_11746);
nand U11981 (N_11981,N_11648,N_11731);
or U11982 (N_11982,N_11528,N_11675);
nand U11983 (N_11983,N_11667,N_11719);
and U11984 (N_11984,N_11527,N_11665);
or U11985 (N_11985,N_11619,N_11745);
nand U11986 (N_11986,N_11524,N_11507);
nor U11987 (N_11987,N_11668,N_11665);
or U11988 (N_11988,N_11709,N_11643);
nor U11989 (N_11989,N_11688,N_11732);
and U11990 (N_11990,N_11691,N_11606);
nand U11991 (N_11991,N_11713,N_11708);
or U11992 (N_11992,N_11566,N_11720);
or U11993 (N_11993,N_11683,N_11635);
nor U11994 (N_11994,N_11692,N_11658);
nor U11995 (N_11995,N_11645,N_11525);
nand U11996 (N_11996,N_11532,N_11633);
or U11997 (N_11997,N_11551,N_11540);
nand U11998 (N_11998,N_11537,N_11562);
and U11999 (N_11999,N_11510,N_11559);
nor U12000 (N_12000,N_11860,N_11987);
nor U12001 (N_12001,N_11796,N_11857);
or U12002 (N_12002,N_11958,N_11880);
nand U12003 (N_12003,N_11787,N_11955);
nor U12004 (N_12004,N_11844,N_11895);
or U12005 (N_12005,N_11891,N_11798);
or U12006 (N_12006,N_11992,N_11766);
or U12007 (N_12007,N_11756,N_11911);
and U12008 (N_12008,N_11882,N_11863);
or U12009 (N_12009,N_11791,N_11840);
nor U12010 (N_12010,N_11765,N_11754);
xor U12011 (N_12011,N_11918,N_11817);
and U12012 (N_12012,N_11977,N_11776);
xor U12013 (N_12013,N_11871,N_11964);
and U12014 (N_12014,N_11973,N_11782);
and U12015 (N_12015,N_11949,N_11897);
nor U12016 (N_12016,N_11957,N_11861);
nor U12017 (N_12017,N_11773,N_11874);
xor U12018 (N_12018,N_11947,N_11758);
nor U12019 (N_12019,N_11953,N_11984);
and U12020 (N_12020,N_11907,N_11997);
and U12021 (N_12021,N_11944,N_11780);
and U12022 (N_12022,N_11757,N_11785);
and U12023 (N_12023,N_11981,N_11793);
and U12024 (N_12024,N_11879,N_11774);
nand U12025 (N_12025,N_11872,N_11956);
nand U12026 (N_12026,N_11814,N_11959);
and U12027 (N_12027,N_11760,N_11925);
nor U12028 (N_12028,N_11779,N_11873);
or U12029 (N_12029,N_11883,N_11930);
nor U12030 (N_12030,N_11846,N_11941);
and U12031 (N_12031,N_11762,N_11750);
or U12032 (N_12032,N_11868,N_11994);
nand U12033 (N_12033,N_11795,N_11892);
nand U12034 (N_12034,N_11838,N_11881);
and U12035 (N_12035,N_11853,N_11832);
or U12036 (N_12036,N_11858,N_11917);
or U12037 (N_12037,N_11970,N_11940);
nor U12038 (N_12038,N_11971,N_11811);
or U12039 (N_12039,N_11886,N_11968);
xnor U12040 (N_12040,N_11806,N_11933);
or U12041 (N_12041,N_11797,N_11979);
or U12042 (N_12042,N_11996,N_11915);
nand U12043 (N_12043,N_11781,N_11904);
and U12044 (N_12044,N_11835,N_11764);
and U12045 (N_12045,N_11829,N_11922);
and U12046 (N_12046,N_11908,N_11923);
or U12047 (N_12047,N_11901,N_11928);
nor U12048 (N_12048,N_11768,N_11753);
nand U12049 (N_12049,N_11802,N_11805);
and U12050 (N_12050,N_11788,N_11910);
nor U12051 (N_12051,N_11885,N_11951);
nand U12052 (N_12052,N_11999,N_11914);
nor U12053 (N_12053,N_11842,N_11893);
nand U12054 (N_12054,N_11896,N_11841);
nand U12055 (N_12055,N_11986,N_11899);
or U12056 (N_12056,N_11920,N_11943);
nor U12057 (N_12057,N_11852,N_11913);
nand U12058 (N_12058,N_11831,N_11888);
nand U12059 (N_12059,N_11794,N_11761);
or U12060 (N_12060,N_11803,N_11804);
or U12061 (N_12061,N_11869,N_11813);
nand U12062 (N_12062,N_11890,N_11812);
nand U12063 (N_12063,N_11849,N_11902);
or U12064 (N_12064,N_11822,N_11837);
nand U12065 (N_12065,N_11755,N_11909);
or U12066 (N_12066,N_11998,N_11912);
nor U12067 (N_12067,N_11966,N_11942);
nor U12068 (N_12068,N_11786,N_11752);
nor U12069 (N_12069,N_11789,N_11865);
and U12070 (N_12070,N_11825,N_11900);
or U12071 (N_12071,N_11801,N_11939);
or U12072 (N_12072,N_11894,N_11839);
nor U12073 (N_12073,N_11887,N_11830);
nand U12074 (N_12074,N_11864,N_11969);
and U12075 (N_12075,N_11763,N_11936);
nand U12076 (N_12076,N_11870,N_11967);
nor U12077 (N_12077,N_11995,N_11989);
or U12078 (N_12078,N_11961,N_11851);
and U12079 (N_12079,N_11905,N_11772);
nor U12080 (N_12080,N_11937,N_11847);
or U12081 (N_12081,N_11916,N_11862);
and U12082 (N_12082,N_11921,N_11935);
or U12083 (N_12083,N_11821,N_11827);
xor U12084 (N_12084,N_11898,N_11850);
and U12085 (N_12085,N_11990,N_11972);
nor U12086 (N_12086,N_11924,N_11978);
or U12087 (N_12087,N_11878,N_11819);
nor U12088 (N_12088,N_11783,N_11919);
nor U12089 (N_12089,N_11867,N_11884);
nand U12090 (N_12090,N_11877,N_11843);
nand U12091 (N_12091,N_11963,N_11960);
nor U12092 (N_12092,N_11751,N_11775);
or U12093 (N_12093,N_11770,N_11815);
nand U12094 (N_12094,N_11962,N_11906);
nor U12095 (N_12095,N_11808,N_11982);
nor U12096 (N_12096,N_11771,N_11777);
and U12097 (N_12097,N_11809,N_11927);
and U12098 (N_12098,N_11816,N_11988);
nor U12099 (N_12099,N_11845,N_11950);
and U12100 (N_12100,N_11820,N_11934);
nor U12101 (N_12101,N_11929,N_11800);
nand U12102 (N_12102,N_11903,N_11856);
and U12103 (N_12103,N_11790,N_11759);
nand U12104 (N_12104,N_11807,N_11965);
nor U12105 (N_12105,N_11866,N_11859);
nand U12106 (N_12106,N_11784,N_11932);
and U12107 (N_12107,N_11945,N_11792);
and U12108 (N_12108,N_11799,N_11833);
and U12109 (N_12109,N_11855,N_11875);
nor U12110 (N_12110,N_11931,N_11767);
and U12111 (N_12111,N_11976,N_11938);
or U12112 (N_12112,N_11854,N_11848);
nor U12113 (N_12113,N_11983,N_11769);
and U12114 (N_12114,N_11974,N_11889);
or U12115 (N_12115,N_11810,N_11948);
and U12116 (N_12116,N_11991,N_11954);
and U12117 (N_12117,N_11876,N_11818);
nor U12118 (N_12118,N_11778,N_11993);
nor U12119 (N_12119,N_11975,N_11834);
and U12120 (N_12120,N_11836,N_11824);
nor U12121 (N_12121,N_11946,N_11823);
and U12122 (N_12122,N_11926,N_11952);
or U12123 (N_12123,N_11980,N_11826);
nand U12124 (N_12124,N_11828,N_11985);
nand U12125 (N_12125,N_11773,N_11877);
nand U12126 (N_12126,N_11833,N_11986);
and U12127 (N_12127,N_11917,N_11880);
or U12128 (N_12128,N_11922,N_11860);
or U12129 (N_12129,N_11988,N_11917);
nor U12130 (N_12130,N_11941,N_11979);
nor U12131 (N_12131,N_11922,N_11911);
or U12132 (N_12132,N_11880,N_11865);
or U12133 (N_12133,N_11771,N_11825);
or U12134 (N_12134,N_11815,N_11938);
or U12135 (N_12135,N_11880,N_11871);
and U12136 (N_12136,N_11993,N_11791);
nand U12137 (N_12137,N_11886,N_11939);
or U12138 (N_12138,N_11900,N_11911);
or U12139 (N_12139,N_11807,N_11990);
or U12140 (N_12140,N_11761,N_11934);
and U12141 (N_12141,N_11913,N_11915);
nand U12142 (N_12142,N_11787,N_11862);
or U12143 (N_12143,N_11865,N_11901);
nor U12144 (N_12144,N_11879,N_11779);
or U12145 (N_12145,N_11979,N_11807);
nor U12146 (N_12146,N_11849,N_11839);
or U12147 (N_12147,N_11958,N_11965);
or U12148 (N_12148,N_11795,N_11992);
nand U12149 (N_12149,N_11761,N_11832);
and U12150 (N_12150,N_11856,N_11936);
and U12151 (N_12151,N_11771,N_11967);
nor U12152 (N_12152,N_11973,N_11955);
nor U12153 (N_12153,N_11810,N_11988);
nor U12154 (N_12154,N_11851,N_11818);
and U12155 (N_12155,N_11868,N_11864);
nand U12156 (N_12156,N_11913,N_11870);
or U12157 (N_12157,N_11981,N_11863);
or U12158 (N_12158,N_11907,N_11756);
and U12159 (N_12159,N_11787,N_11918);
and U12160 (N_12160,N_11979,N_11769);
nor U12161 (N_12161,N_11765,N_11797);
nand U12162 (N_12162,N_11925,N_11915);
and U12163 (N_12163,N_11810,N_11792);
and U12164 (N_12164,N_11881,N_11969);
nor U12165 (N_12165,N_11966,N_11909);
xnor U12166 (N_12166,N_11757,N_11767);
nand U12167 (N_12167,N_11886,N_11883);
or U12168 (N_12168,N_11846,N_11870);
nand U12169 (N_12169,N_11853,N_11838);
or U12170 (N_12170,N_11965,N_11756);
and U12171 (N_12171,N_11919,N_11915);
and U12172 (N_12172,N_11920,N_11854);
or U12173 (N_12173,N_11961,N_11924);
nor U12174 (N_12174,N_11937,N_11806);
or U12175 (N_12175,N_11833,N_11885);
nand U12176 (N_12176,N_11788,N_11994);
nor U12177 (N_12177,N_11918,N_11798);
nand U12178 (N_12178,N_11838,N_11992);
or U12179 (N_12179,N_11824,N_11932);
and U12180 (N_12180,N_11945,N_11855);
nor U12181 (N_12181,N_11815,N_11867);
or U12182 (N_12182,N_11921,N_11793);
nand U12183 (N_12183,N_11858,N_11818);
nand U12184 (N_12184,N_11806,N_11965);
or U12185 (N_12185,N_11977,N_11945);
nand U12186 (N_12186,N_11904,N_11777);
or U12187 (N_12187,N_11879,N_11759);
and U12188 (N_12188,N_11900,N_11850);
nand U12189 (N_12189,N_11869,N_11843);
nor U12190 (N_12190,N_11930,N_11769);
or U12191 (N_12191,N_11918,N_11991);
xnor U12192 (N_12192,N_11949,N_11772);
and U12193 (N_12193,N_11760,N_11870);
nor U12194 (N_12194,N_11824,N_11989);
or U12195 (N_12195,N_11772,N_11892);
nor U12196 (N_12196,N_11818,N_11886);
and U12197 (N_12197,N_11809,N_11942);
nor U12198 (N_12198,N_11974,N_11841);
nor U12199 (N_12199,N_11949,N_11905);
or U12200 (N_12200,N_11850,N_11911);
or U12201 (N_12201,N_11860,N_11948);
nand U12202 (N_12202,N_11806,N_11975);
and U12203 (N_12203,N_11845,N_11993);
or U12204 (N_12204,N_11974,N_11921);
nor U12205 (N_12205,N_11932,N_11882);
nor U12206 (N_12206,N_11750,N_11910);
and U12207 (N_12207,N_11963,N_11921);
and U12208 (N_12208,N_11973,N_11810);
nor U12209 (N_12209,N_11875,N_11877);
and U12210 (N_12210,N_11878,N_11952);
xor U12211 (N_12211,N_11932,N_11827);
nand U12212 (N_12212,N_11926,N_11902);
or U12213 (N_12213,N_11935,N_11979);
and U12214 (N_12214,N_11920,N_11879);
or U12215 (N_12215,N_11922,N_11857);
or U12216 (N_12216,N_11880,N_11817);
nor U12217 (N_12217,N_11898,N_11800);
and U12218 (N_12218,N_11782,N_11910);
and U12219 (N_12219,N_11932,N_11815);
or U12220 (N_12220,N_11791,N_11925);
or U12221 (N_12221,N_11947,N_11908);
nor U12222 (N_12222,N_11986,N_11992);
nand U12223 (N_12223,N_11995,N_11820);
nor U12224 (N_12224,N_11765,N_11821);
and U12225 (N_12225,N_11894,N_11906);
nand U12226 (N_12226,N_11905,N_11759);
and U12227 (N_12227,N_11950,N_11965);
and U12228 (N_12228,N_11953,N_11936);
nand U12229 (N_12229,N_11786,N_11789);
and U12230 (N_12230,N_11826,N_11874);
and U12231 (N_12231,N_11980,N_11808);
or U12232 (N_12232,N_11852,N_11988);
nor U12233 (N_12233,N_11962,N_11774);
nand U12234 (N_12234,N_11760,N_11983);
nand U12235 (N_12235,N_11956,N_11772);
nor U12236 (N_12236,N_11773,N_11886);
or U12237 (N_12237,N_11944,N_11805);
and U12238 (N_12238,N_11972,N_11962);
or U12239 (N_12239,N_11958,N_11843);
or U12240 (N_12240,N_11964,N_11963);
nor U12241 (N_12241,N_11954,N_11987);
or U12242 (N_12242,N_11957,N_11960);
and U12243 (N_12243,N_11829,N_11808);
and U12244 (N_12244,N_11975,N_11836);
nor U12245 (N_12245,N_11811,N_11888);
and U12246 (N_12246,N_11955,N_11767);
nor U12247 (N_12247,N_11915,N_11783);
nand U12248 (N_12248,N_11814,N_11952);
nand U12249 (N_12249,N_11826,N_11914);
nand U12250 (N_12250,N_12179,N_12099);
or U12251 (N_12251,N_12203,N_12228);
nor U12252 (N_12252,N_12006,N_12157);
and U12253 (N_12253,N_12005,N_12026);
nand U12254 (N_12254,N_12130,N_12218);
nand U12255 (N_12255,N_12231,N_12238);
and U12256 (N_12256,N_12193,N_12212);
or U12257 (N_12257,N_12014,N_12198);
nor U12258 (N_12258,N_12143,N_12201);
nand U12259 (N_12259,N_12145,N_12183);
or U12260 (N_12260,N_12223,N_12046);
nor U12261 (N_12261,N_12182,N_12208);
or U12262 (N_12262,N_12122,N_12091);
nor U12263 (N_12263,N_12108,N_12103);
and U12264 (N_12264,N_12170,N_12040);
nand U12265 (N_12265,N_12055,N_12081);
or U12266 (N_12266,N_12037,N_12042);
or U12267 (N_12267,N_12032,N_12050);
or U12268 (N_12268,N_12067,N_12240);
nand U12269 (N_12269,N_12142,N_12036);
and U12270 (N_12270,N_12071,N_12158);
and U12271 (N_12271,N_12059,N_12215);
and U12272 (N_12272,N_12156,N_12237);
or U12273 (N_12273,N_12126,N_12074);
nor U12274 (N_12274,N_12008,N_12069);
and U12275 (N_12275,N_12093,N_12058);
nor U12276 (N_12276,N_12001,N_12186);
nor U12277 (N_12277,N_12017,N_12100);
and U12278 (N_12278,N_12094,N_12111);
and U12279 (N_12279,N_12248,N_12224);
nor U12280 (N_12280,N_12194,N_12018);
nand U12281 (N_12281,N_12211,N_12233);
nand U12282 (N_12282,N_12209,N_12173);
and U12283 (N_12283,N_12084,N_12022);
or U12284 (N_12284,N_12129,N_12172);
or U12285 (N_12285,N_12159,N_12007);
nor U12286 (N_12286,N_12025,N_12035);
or U12287 (N_12287,N_12216,N_12119);
nand U12288 (N_12288,N_12152,N_12196);
nand U12289 (N_12289,N_12180,N_12095);
or U12290 (N_12290,N_12057,N_12160);
nand U12291 (N_12291,N_12167,N_12213);
and U12292 (N_12292,N_12133,N_12062);
nand U12293 (N_12293,N_12128,N_12056);
nand U12294 (N_12294,N_12181,N_12178);
and U12295 (N_12295,N_12221,N_12077);
nor U12296 (N_12296,N_12088,N_12080);
and U12297 (N_12297,N_12227,N_12051);
or U12298 (N_12298,N_12150,N_12054);
nand U12299 (N_12299,N_12117,N_12184);
nor U12300 (N_12300,N_12048,N_12086);
nand U12301 (N_12301,N_12164,N_12033);
and U12302 (N_12302,N_12161,N_12245);
nand U12303 (N_12303,N_12134,N_12202);
nor U12304 (N_12304,N_12024,N_12010);
and U12305 (N_12305,N_12234,N_12023);
or U12306 (N_12306,N_12019,N_12235);
and U12307 (N_12307,N_12098,N_12242);
or U12308 (N_12308,N_12174,N_12043);
and U12309 (N_12309,N_12028,N_12169);
nand U12310 (N_12310,N_12092,N_12020);
or U12311 (N_12311,N_12229,N_12105);
or U12312 (N_12312,N_12096,N_12073);
or U12313 (N_12313,N_12244,N_12197);
and U12314 (N_12314,N_12061,N_12199);
nor U12315 (N_12315,N_12038,N_12247);
xor U12316 (N_12316,N_12112,N_12192);
nand U12317 (N_12317,N_12082,N_12226);
nand U12318 (N_12318,N_12187,N_12002);
nand U12319 (N_12319,N_12188,N_12176);
and U12320 (N_12320,N_12041,N_12148);
nor U12321 (N_12321,N_12249,N_12230);
or U12322 (N_12322,N_12149,N_12016);
nor U12323 (N_12323,N_12189,N_12168);
and U12324 (N_12324,N_12217,N_12200);
or U12325 (N_12325,N_12144,N_12047);
nand U12326 (N_12326,N_12232,N_12120);
and U12327 (N_12327,N_12013,N_12075);
nor U12328 (N_12328,N_12078,N_12015);
nand U12329 (N_12329,N_12177,N_12190);
and U12330 (N_12330,N_12021,N_12085);
nor U12331 (N_12331,N_12039,N_12027);
nand U12332 (N_12332,N_12205,N_12243);
or U12333 (N_12333,N_12009,N_12004);
nand U12334 (N_12334,N_12204,N_12139);
and U12335 (N_12335,N_12166,N_12060);
nor U12336 (N_12336,N_12125,N_12011);
or U12337 (N_12337,N_12191,N_12109);
nor U12338 (N_12338,N_12163,N_12153);
nand U12339 (N_12339,N_12155,N_12070);
nor U12340 (N_12340,N_12135,N_12045);
nor U12341 (N_12341,N_12000,N_12171);
xnor U12342 (N_12342,N_12137,N_12131);
or U12343 (N_12343,N_12101,N_12031);
nor U12344 (N_12344,N_12003,N_12102);
xor U12345 (N_12345,N_12123,N_12034);
nor U12346 (N_12346,N_12151,N_12147);
or U12347 (N_12347,N_12063,N_12175);
nand U12348 (N_12348,N_12110,N_12210);
nand U12349 (N_12349,N_12104,N_12089);
and U12350 (N_12350,N_12165,N_12049);
or U12351 (N_12351,N_12053,N_12116);
and U12352 (N_12352,N_12124,N_12207);
or U12353 (N_12353,N_12107,N_12138);
nand U12354 (N_12354,N_12206,N_12114);
or U12355 (N_12355,N_12044,N_12185);
or U12356 (N_12356,N_12141,N_12090);
or U12357 (N_12357,N_12065,N_12064);
or U12358 (N_12358,N_12072,N_12136);
and U12359 (N_12359,N_12236,N_12083);
nand U12360 (N_12360,N_12162,N_12146);
or U12361 (N_12361,N_12079,N_12030);
nand U12362 (N_12362,N_12068,N_12118);
or U12363 (N_12363,N_12115,N_12241);
and U12364 (N_12364,N_12012,N_12140);
or U12365 (N_12365,N_12214,N_12195);
nand U12366 (N_12366,N_12220,N_12097);
and U12367 (N_12367,N_12127,N_12087);
and U12368 (N_12368,N_12246,N_12106);
and U12369 (N_12369,N_12076,N_12225);
nor U12370 (N_12370,N_12219,N_12029);
nand U12371 (N_12371,N_12052,N_12239);
and U12372 (N_12372,N_12154,N_12066);
or U12373 (N_12373,N_12121,N_12132);
nand U12374 (N_12374,N_12113,N_12222);
and U12375 (N_12375,N_12118,N_12099);
nor U12376 (N_12376,N_12175,N_12104);
and U12377 (N_12377,N_12043,N_12138);
and U12378 (N_12378,N_12066,N_12199);
nand U12379 (N_12379,N_12090,N_12243);
nand U12380 (N_12380,N_12000,N_12032);
nand U12381 (N_12381,N_12223,N_12106);
or U12382 (N_12382,N_12245,N_12122);
or U12383 (N_12383,N_12188,N_12029);
and U12384 (N_12384,N_12159,N_12066);
nor U12385 (N_12385,N_12230,N_12208);
and U12386 (N_12386,N_12116,N_12001);
nor U12387 (N_12387,N_12200,N_12013);
and U12388 (N_12388,N_12128,N_12157);
and U12389 (N_12389,N_12035,N_12010);
or U12390 (N_12390,N_12154,N_12111);
nand U12391 (N_12391,N_12131,N_12041);
nor U12392 (N_12392,N_12019,N_12098);
or U12393 (N_12393,N_12195,N_12166);
nor U12394 (N_12394,N_12239,N_12203);
or U12395 (N_12395,N_12202,N_12063);
nand U12396 (N_12396,N_12166,N_12130);
nor U12397 (N_12397,N_12123,N_12017);
and U12398 (N_12398,N_12124,N_12012);
nor U12399 (N_12399,N_12133,N_12247);
or U12400 (N_12400,N_12183,N_12012);
and U12401 (N_12401,N_12161,N_12194);
nand U12402 (N_12402,N_12078,N_12128);
or U12403 (N_12403,N_12052,N_12247);
and U12404 (N_12404,N_12148,N_12187);
and U12405 (N_12405,N_12094,N_12144);
nor U12406 (N_12406,N_12198,N_12059);
nor U12407 (N_12407,N_12023,N_12197);
or U12408 (N_12408,N_12040,N_12111);
or U12409 (N_12409,N_12168,N_12084);
or U12410 (N_12410,N_12244,N_12220);
nor U12411 (N_12411,N_12243,N_12151);
nand U12412 (N_12412,N_12222,N_12073);
and U12413 (N_12413,N_12003,N_12025);
and U12414 (N_12414,N_12100,N_12194);
nand U12415 (N_12415,N_12034,N_12028);
or U12416 (N_12416,N_12093,N_12088);
nand U12417 (N_12417,N_12064,N_12155);
nor U12418 (N_12418,N_12195,N_12237);
or U12419 (N_12419,N_12076,N_12031);
nand U12420 (N_12420,N_12231,N_12076);
or U12421 (N_12421,N_12109,N_12158);
nor U12422 (N_12422,N_12160,N_12064);
and U12423 (N_12423,N_12054,N_12061);
nor U12424 (N_12424,N_12084,N_12040);
and U12425 (N_12425,N_12066,N_12185);
and U12426 (N_12426,N_12067,N_12172);
and U12427 (N_12427,N_12247,N_12150);
or U12428 (N_12428,N_12085,N_12204);
or U12429 (N_12429,N_12222,N_12038);
nand U12430 (N_12430,N_12083,N_12005);
nand U12431 (N_12431,N_12010,N_12051);
nor U12432 (N_12432,N_12148,N_12105);
and U12433 (N_12433,N_12138,N_12140);
nand U12434 (N_12434,N_12014,N_12193);
nand U12435 (N_12435,N_12176,N_12237);
or U12436 (N_12436,N_12210,N_12038);
nor U12437 (N_12437,N_12248,N_12078);
nor U12438 (N_12438,N_12170,N_12147);
nand U12439 (N_12439,N_12227,N_12091);
and U12440 (N_12440,N_12060,N_12154);
or U12441 (N_12441,N_12188,N_12198);
or U12442 (N_12442,N_12010,N_12167);
nor U12443 (N_12443,N_12098,N_12216);
or U12444 (N_12444,N_12170,N_12182);
nor U12445 (N_12445,N_12132,N_12048);
nand U12446 (N_12446,N_12164,N_12145);
nor U12447 (N_12447,N_12233,N_12140);
nand U12448 (N_12448,N_12072,N_12126);
or U12449 (N_12449,N_12124,N_12089);
nand U12450 (N_12450,N_12106,N_12075);
and U12451 (N_12451,N_12136,N_12109);
nor U12452 (N_12452,N_12003,N_12213);
or U12453 (N_12453,N_12091,N_12139);
or U12454 (N_12454,N_12061,N_12111);
and U12455 (N_12455,N_12141,N_12202);
and U12456 (N_12456,N_12125,N_12222);
nand U12457 (N_12457,N_12127,N_12115);
and U12458 (N_12458,N_12085,N_12193);
nor U12459 (N_12459,N_12058,N_12051);
nand U12460 (N_12460,N_12172,N_12140);
nand U12461 (N_12461,N_12190,N_12000);
nor U12462 (N_12462,N_12079,N_12041);
nand U12463 (N_12463,N_12081,N_12173);
and U12464 (N_12464,N_12150,N_12240);
nand U12465 (N_12465,N_12058,N_12198);
or U12466 (N_12466,N_12095,N_12221);
and U12467 (N_12467,N_12045,N_12241);
or U12468 (N_12468,N_12166,N_12199);
nand U12469 (N_12469,N_12173,N_12181);
and U12470 (N_12470,N_12142,N_12099);
nor U12471 (N_12471,N_12232,N_12239);
nand U12472 (N_12472,N_12075,N_12244);
nor U12473 (N_12473,N_12173,N_12247);
nand U12474 (N_12474,N_12065,N_12067);
xor U12475 (N_12475,N_12137,N_12123);
nor U12476 (N_12476,N_12224,N_12209);
nor U12477 (N_12477,N_12165,N_12215);
or U12478 (N_12478,N_12174,N_12234);
or U12479 (N_12479,N_12065,N_12076);
nor U12480 (N_12480,N_12134,N_12100);
nand U12481 (N_12481,N_12090,N_12003);
or U12482 (N_12482,N_12036,N_12038);
and U12483 (N_12483,N_12102,N_12038);
and U12484 (N_12484,N_12244,N_12228);
nor U12485 (N_12485,N_12202,N_12028);
or U12486 (N_12486,N_12093,N_12226);
or U12487 (N_12487,N_12030,N_12048);
nand U12488 (N_12488,N_12124,N_12053);
nor U12489 (N_12489,N_12188,N_12220);
nor U12490 (N_12490,N_12209,N_12097);
nor U12491 (N_12491,N_12076,N_12226);
nor U12492 (N_12492,N_12136,N_12247);
and U12493 (N_12493,N_12189,N_12093);
nor U12494 (N_12494,N_12238,N_12203);
or U12495 (N_12495,N_12203,N_12029);
nor U12496 (N_12496,N_12089,N_12152);
nand U12497 (N_12497,N_12209,N_12093);
and U12498 (N_12498,N_12130,N_12131);
or U12499 (N_12499,N_12192,N_12156);
nand U12500 (N_12500,N_12430,N_12290);
or U12501 (N_12501,N_12255,N_12335);
and U12502 (N_12502,N_12317,N_12341);
and U12503 (N_12503,N_12372,N_12411);
nand U12504 (N_12504,N_12497,N_12428);
nor U12505 (N_12505,N_12443,N_12307);
nor U12506 (N_12506,N_12412,N_12304);
nor U12507 (N_12507,N_12362,N_12333);
nand U12508 (N_12508,N_12297,N_12293);
and U12509 (N_12509,N_12311,N_12262);
or U12510 (N_12510,N_12295,N_12254);
or U12511 (N_12511,N_12298,N_12488);
nand U12512 (N_12512,N_12460,N_12259);
nor U12513 (N_12513,N_12442,N_12452);
or U12514 (N_12514,N_12466,N_12356);
nand U12515 (N_12515,N_12454,N_12332);
nand U12516 (N_12516,N_12257,N_12338);
or U12517 (N_12517,N_12449,N_12274);
or U12518 (N_12518,N_12376,N_12471);
nor U12519 (N_12519,N_12263,N_12331);
or U12520 (N_12520,N_12299,N_12380);
nor U12521 (N_12521,N_12432,N_12426);
and U12522 (N_12522,N_12374,N_12422);
nor U12523 (N_12523,N_12472,N_12327);
nand U12524 (N_12524,N_12282,N_12347);
and U12525 (N_12525,N_12403,N_12370);
nand U12526 (N_12526,N_12277,N_12379);
nor U12527 (N_12527,N_12389,N_12294);
nand U12528 (N_12528,N_12283,N_12339);
nand U12529 (N_12529,N_12387,N_12336);
or U12530 (N_12530,N_12324,N_12329);
or U12531 (N_12531,N_12400,N_12289);
or U12532 (N_12532,N_12318,N_12438);
nor U12533 (N_12533,N_12477,N_12425);
nor U12534 (N_12534,N_12482,N_12485);
nor U12535 (N_12535,N_12349,N_12463);
or U12536 (N_12536,N_12405,N_12490);
and U12537 (N_12537,N_12384,N_12258);
and U12538 (N_12538,N_12351,N_12366);
or U12539 (N_12539,N_12253,N_12433);
or U12540 (N_12540,N_12291,N_12325);
or U12541 (N_12541,N_12464,N_12365);
or U12542 (N_12542,N_12421,N_12462);
nor U12543 (N_12543,N_12413,N_12252);
or U12544 (N_12544,N_12381,N_12456);
nor U12545 (N_12545,N_12267,N_12494);
nand U12546 (N_12546,N_12355,N_12396);
nand U12547 (N_12547,N_12260,N_12371);
nor U12548 (N_12548,N_12358,N_12489);
nand U12549 (N_12549,N_12447,N_12465);
nand U12550 (N_12550,N_12314,N_12306);
nor U12551 (N_12551,N_12352,N_12315);
or U12552 (N_12552,N_12287,N_12266);
nor U12553 (N_12553,N_12278,N_12346);
and U12554 (N_12554,N_12394,N_12469);
or U12555 (N_12555,N_12491,N_12303);
and U12556 (N_12556,N_12264,N_12367);
nor U12557 (N_12557,N_12453,N_12310);
nand U12558 (N_12558,N_12328,N_12334);
nor U12559 (N_12559,N_12281,N_12495);
nor U12560 (N_12560,N_12431,N_12316);
and U12561 (N_12561,N_12340,N_12499);
or U12562 (N_12562,N_12417,N_12312);
and U12563 (N_12563,N_12269,N_12300);
nor U12564 (N_12564,N_12343,N_12481);
or U12565 (N_12565,N_12437,N_12345);
nand U12566 (N_12566,N_12302,N_12377);
nand U12567 (N_12567,N_12492,N_12368);
and U12568 (N_12568,N_12418,N_12326);
nand U12569 (N_12569,N_12439,N_12448);
or U12570 (N_12570,N_12383,N_12408);
and U12571 (N_12571,N_12409,N_12280);
nand U12572 (N_12572,N_12450,N_12251);
and U12573 (N_12573,N_12475,N_12385);
and U12574 (N_12574,N_12313,N_12458);
and U12575 (N_12575,N_12480,N_12423);
nand U12576 (N_12576,N_12434,N_12342);
and U12577 (N_12577,N_12440,N_12337);
and U12578 (N_12578,N_12271,N_12410);
nor U12579 (N_12579,N_12470,N_12415);
nand U12580 (N_12580,N_12323,N_12395);
and U12581 (N_12581,N_12397,N_12373);
and U12582 (N_12582,N_12375,N_12436);
or U12583 (N_12583,N_12451,N_12445);
and U12584 (N_12584,N_12364,N_12479);
and U12585 (N_12585,N_12406,N_12285);
nor U12586 (N_12586,N_12378,N_12399);
and U12587 (N_12587,N_12476,N_12392);
nand U12588 (N_12588,N_12292,N_12390);
nor U12589 (N_12589,N_12330,N_12478);
and U12590 (N_12590,N_12435,N_12286);
nand U12591 (N_12591,N_12359,N_12461);
and U12592 (N_12592,N_12350,N_12496);
and U12593 (N_12593,N_12270,N_12401);
and U12594 (N_12594,N_12484,N_12427);
nor U12595 (N_12595,N_12361,N_12309);
or U12596 (N_12596,N_12357,N_12473);
nand U12597 (N_12597,N_12275,N_12429);
or U12598 (N_12598,N_12256,N_12288);
nor U12599 (N_12599,N_12322,N_12321);
nor U12600 (N_12600,N_12402,N_12414);
or U12601 (N_12601,N_12360,N_12457);
or U12602 (N_12602,N_12424,N_12261);
or U12603 (N_12603,N_12455,N_12284);
or U12604 (N_12604,N_12301,N_12474);
and U12605 (N_12605,N_12363,N_12268);
and U12606 (N_12606,N_12369,N_12483);
nor U12607 (N_12607,N_12420,N_12441);
xnor U12608 (N_12608,N_12498,N_12446);
nor U12609 (N_12609,N_12386,N_12250);
nor U12610 (N_12610,N_12404,N_12305);
or U12611 (N_12611,N_12272,N_12468);
and U12612 (N_12612,N_12416,N_12354);
nor U12613 (N_12613,N_12388,N_12486);
or U12614 (N_12614,N_12487,N_12320);
nor U12615 (N_12615,N_12344,N_12419);
nand U12616 (N_12616,N_12493,N_12393);
nor U12617 (N_12617,N_12296,N_12398);
or U12618 (N_12618,N_12276,N_12444);
nand U12619 (N_12619,N_12353,N_12279);
nand U12620 (N_12620,N_12265,N_12273);
nand U12621 (N_12621,N_12391,N_12348);
nand U12622 (N_12622,N_12467,N_12308);
and U12623 (N_12623,N_12382,N_12319);
nor U12624 (N_12624,N_12459,N_12407);
or U12625 (N_12625,N_12436,N_12392);
and U12626 (N_12626,N_12420,N_12282);
nor U12627 (N_12627,N_12403,N_12266);
nor U12628 (N_12628,N_12471,N_12367);
nand U12629 (N_12629,N_12435,N_12415);
or U12630 (N_12630,N_12348,N_12400);
or U12631 (N_12631,N_12409,N_12331);
nor U12632 (N_12632,N_12286,N_12481);
xnor U12633 (N_12633,N_12410,N_12476);
nand U12634 (N_12634,N_12475,N_12462);
nand U12635 (N_12635,N_12374,N_12383);
nand U12636 (N_12636,N_12347,N_12435);
nor U12637 (N_12637,N_12278,N_12384);
nand U12638 (N_12638,N_12471,N_12277);
nand U12639 (N_12639,N_12285,N_12334);
nor U12640 (N_12640,N_12252,N_12495);
or U12641 (N_12641,N_12478,N_12371);
and U12642 (N_12642,N_12479,N_12353);
nor U12643 (N_12643,N_12338,N_12396);
xnor U12644 (N_12644,N_12346,N_12303);
nand U12645 (N_12645,N_12342,N_12294);
nor U12646 (N_12646,N_12324,N_12404);
nor U12647 (N_12647,N_12383,N_12291);
nor U12648 (N_12648,N_12462,N_12425);
or U12649 (N_12649,N_12316,N_12346);
or U12650 (N_12650,N_12254,N_12285);
and U12651 (N_12651,N_12297,N_12405);
nor U12652 (N_12652,N_12483,N_12373);
or U12653 (N_12653,N_12382,N_12442);
or U12654 (N_12654,N_12272,N_12259);
nor U12655 (N_12655,N_12265,N_12305);
nand U12656 (N_12656,N_12339,N_12354);
nand U12657 (N_12657,N_12426,N_12260);
nor U12658 (N_12658,N_12397,N_12358);
nor U12659 (N_12659,N_12399,N_12302);
and U12660 (N_12660,N_12443,N_12421);
nand U12661 (N_12661,N_12433,N_12295);
xor U12662 (N_12662,N_12352,N_12263);
and U12663 (N_12663,N_12425,N_12402);
or U12664 (N_12664,N_12267,N_12250);
nand U12665 (N_12665,N_12489,N_12459);
and U12666 (N_12666,N_12476,N_12268);
nor U12667 (N_12667,N_12497,N_12493);
or U12668 (N_12668,N_12400,N_12380);
nor U12669 (N_12669,N_12416,N_12467);
and U12670 (N_12670,N_12330,N_12267);
and U12671 (N_12671,N_12417,N_12481);
nor U12672 (N_12672,N_12346,N_12342);
or U12673 (N_12673,N_12328,N_12407);
or U12674 (N_12674,N_12375,N_12340);
and U12675 (N_12675,N_12349,N_12419);
and U12676 (N_12676,N_12486,N_12310);
nor U12677 (N_12677,N_12364,N_12450);
or U12678 (N_12678,N_12471,N_12278);
and U12679 (N_12679,N_12290,N_12376);
and U12680 (N_12680,N_12433,N_12416);
nand U12681 (N_12681,N_12497,N_12461);
nand U12682 (N_12682,N_12491,N_12305);
or U12683 (N_12683,N_12292,N_12407);
or U12684 (N_12684,N_12290,N_12490);
or U12685 (N_12685,N_12348,N_12444);
nor U12686 (N_12686,N_12394,N_12360);
xor U12687 (N_12687,N_12433,N_12463);
or U12688 (N_12688,N_12251,N_12449);
nor U12689 (N_12689,N_12433,N_12280);
or U12690 (N_12690,N_12433,N_12426);
and U12691 (N_12691,N_12448,N_12499);
or U12692 (N_12692,N_12320,N_12383);
nor U12693 (N_12693,N_12317,N_12453);
nand U12694 (N_12694,N_12294,N_12280);
or U12695 (N_12695,N_12417,N_12421);
nor U12696 (N_12696,N_12302,N_12464);
or U12697 (N_12697,N_12428,N_12382);
or U12698 (N_12698,N_12458,N_12433);
nand U12699 (N_12699,N_12366,N_12414);
xnor U12700 (N_12700,N_12333,N_12295);
nor U12701 (N_12701,N_12381,N_12379);
or U12702 (N_12702,N_12339,N_12325);
and U12703 (N_12703,N_12371,N_12369);
or U12704 (N_12704,N_12378,N_12452);
nor U12705 (N_12705,N_12327,N_12386);
and U12706 (N_12706,N_12411,N_12492);
nand U12707 (N_12707,N_12293,N_12394);
nor U12708 (N_12708,N_12300,N_12265);
or U12709 (N_12709,N_12459,N_12306);
xor U12710 (N_12710,N_12293,N_12445);
and U12711 (N_12711,N_12348,N_12471);
and U12712 (N_12712,N_12408,N_12380);
or U12713 (N_12713,N_12306,N_12328);
or U12714 (N_12714,N_12449,N_12460);
and U12715 (N_12715,N_12416,N_12317);
and U12716 (N_12716,N_12337,N_12267);
nor U12717 (N_12717,N_12415,N_12392);
or U12718 (N_12718,N_12362,N_12411);
and U12719 (N_12719,N_12368,N_12384);
nand U12720 (N_12720,N_12444,N_12369);
nor U12721 (N_12721,N_12386,N_12457);
and U12722 (N_12722,N_12272,N_12258);
nor U12723 (N_12723,N_12438,N_12489);
nand U12724 (N_12724,N_12467,N_12327);
and U12725 (N_12725,N_12478,N_12360);
or U12726 (N_12726,N_12468,N_12408);
nand U12727 (N_12727,N_12298,N_12348);
nor U12728 (N_12728,N_12392,N_12383);
or U12729 (N_12729,N_12392,N_12343);
nand U12730 (N_12730,N_12337,N_12364);
and U12731 (N_12731,N_12370,N_12322);
nor U12732 (N_12732,N_12287,N_12411);
nor U12733 (N_12733,N_12473,N_12460);
or U12734 (N_12734,N_12387,N_12369);
and U12735 (N_12735,N_12429,N_12335);
and U12736 (N_12736,N_12337,N_12316);
and U12737 (N_12737,N_12345,N_12391);
or U12738 (N_12738,N_12432,N_12403);
nor U12739 (N_12739,N_12287,N_12391);
and U12740 (N_12740,N_12314,N_12393);
nor U12741 (N_12741,N_12457,N_12305);
nor U12742 (N_12742,N_12392,N_12420);
or U12743 (N_12743,N_12354,N_12397);
nor U12744 (N_12744,N_12439,N_12290);
nand U12745 (N_12745,N_12391,N_12449);
nand U12746 (N_12746,N_12444,N_12337);
and U12747 (N_12747,N_12487,N_12272);
nor U12748 (N_12748,N_12307,N_12263);
and U12749 (N_12749,N_12340,N_12323);
and U12750 (N_12750,N_12659,N_12625);
and U12751 (N_12751,N_12613,N_12538);
nand U12752 (N_12752,N_12656,N_12629);
nor U12753 (N_12753,N_12627,N_12644);
or U12754 (N_12754,N_12621,N_12559);
nand U12755 (N_12755,N_12636,N_12679);
nand U12756 (N_12756,N_12558,N_12686);
nand U12757 (N_12757,N_12556,N_12557);
nand U12758 (N_12758,N_12716,N_12701);
nor U12759 (N_12759,N_12631,N_12544);
and U12760 (N_12760,N_12720,N_12535);
and U12761 (N_12761,N_12733,N_12746);
or U12762 (N_12762,N_12622,N_12591);
nor U12763 (N_12763,N_12582,N_12673);
or U12764 (N_12764,N_12642,N_12731);
nor U12765 (N_12765,N_12569,N_12587);
and U12766 (N_12766,N_12518,N_12522);
or U12767 (N_12767,N_12732,N_12648);
and U12768 (N_12768,N_12555,N_12657);
and U12769 (N_12769,N_12708,N_12521);
or U12770 (N_12770,N_12712,N_12566);
nand U12771 (N_12771,N_12589,N_12570);
nor U12772 (N_12772,N_12601,N_12743);
nand U12773 (N_12773,N_12660,N_12742);
nor U12774 (N_12774,N_12586,N_12704);
nor U12775 (N_12775,N_12689,N_12501);
nor U12776 (N_12776,N_12547,N_12663);
and U12777 (N_12777,N_12635,N_12739);
and U12778 (N_12778,N_12724,N_12576);
or U12779 (N_12779,N_12696,N_12548);
or U12780 (N_12780,N_12740,N_12513);
or U12781 (N_12781,N_12512,N_12706);
nand U12782 (N_12782,N_12605,N_12700);
nand U12783 (N_12783,N_12607,N_12585);
or U12784 (N_12784,N_12718,N_12672);
or U12785 (N_12785,N_12667,N_12614);
or U12786 (N_12786,N_12617,N_12530);
nor U12787 (N_12787,N_12736,N_12647);
nor U12788 (N_12788,N_12688,N_12502);
nor U12789 (N_12789,N_12705,N_12504);
and U12790 (N_12790,N_12514,N_12674);
and U12791 (N_12791,N_12537,N_12630);
or U12792 (N_12792,N_12602,N_12722);
and U12793 (N_12793,N_12598,N_12577);
nand U12794 (N_12794,N_12632,N_12580);
or U12795 (N_12795,N_12610,N_12734);
or U12796 (N_12796,N_12531,N_12568);
nand U12797 (N_12797,N_12562,N_12620);
nand U12798 (N_12798,N_12594,N_12600);
and U12799 (N_12799,N_12729,N_12698);
nand U12800 (N_12800,N_12626,N_12539);
or U12801 (N_12801,N_12633,N_12721);
and U12802 (N_12802,N_12683,N_12572);
nand U12803 (N_12803,N_12609,N_12714);
and U12804 (N_12804,N_12578,N_12552);
or U12805 (N_12805,N_12604,N_12678);
or U12806 (N_12806,N_12612,N_12677);
nand U12807 (N_12807,N_12618,N_12575);
or U12808 (N_12808,N_12694,N_12643);
and U12809 (N_12809,N_12608,N_12709);
nor U12810 (N_12810,N_12713,N_12682);
or U12811 (N_12811,N_12534,N_12654);
nor U12812 (N_12812,N_12543,N_12540);
nor U12813 (N_12813,N_12728,N_12524);
or U12814 (N_12814,N_12662,N_12615);
nand U12815 (N_12815,N_12549,N_12503);
and U12816 (N_12816,N_12671,N_12588);
nor U12817 (N_12817,N_12645,N_12745);
and U12818 (N_12818,N_12520,N_12687);
nor U12819 (N_12819,N_12695,N_12725);
nor U12820 (N_12820,N_12646,N_12699);
nor U12821 (N_12821,N_12596,N_12649);
and U12822 (N_12822,N_12655,N_12541);
nand U12823 (N_12823,N_12639,N_12691);
nor U12824 (N_12824,N_12545,N_12719);
or U12825 (N_12825,N_12510,N_12593);
xnor U12826 (N_12826,N_12542,N_12500);
nand U12827 (N_12827,N_12685,N_12737);
and U12828 (N_12828,N_12669,N_12507);
nand U12829 (N_12829,N_12567,N_12735);
nor U12830 (N_12830,N_12707,N_12525);
nand U12831 (N_12831,N_12564,N_12628);
nor U12832 (N_12832,N_12563,N_12550);
nor U12833 (N_12833,N_12527,N_12595);
nand U12834 (N_12834,N_12748,N_12658);
and U12835 (N_12835,N_12711,N_12738);
or U12836 (N_12836,N_12680,N_12692);
nor U12837 (N_12837,N_12505,N_12747);
nand U12838 (N_12838,N_12515,N_12681);
nor U12839 (N_12839,N_12560,N_12710);
nand U12840 (N_12840,N_12693,N_12641);
and U12841 (N_12841,N_12611,N_12727);
nor U12842 (N_12842,N_12652,N_12638);
and U12843 (N_12843,N_12616,N_12551);
nand U12844 (N_12844,N_12583,N_12623);
and U12845 (N_12845,N_12508,N_12670);
or U12846 (N_12846,N_12723,N_12573);
nor U12847 (N_12847,N_12690,N_12624);
and U12848 (N_12848,N_12592,N_12697);
nand U12849 (N_12849,N_12553,N_12581);
nand U12850 (N_12850,N_12509,N_12741);
or U12851 (N_12851,N_12634,N_12717);
nor U12852 (N_12852,N_12715,N_12651);
nor U12853 (N_12853,N_12619,N_12640);
or U12854 (N_12854,N_12726,N_12584);
nand U12855 (N_12855,N_12650,N_12599);
nand U12856 (N_12856,N_12561,N_12675);
and U12857 (N_12857,N_12637,N_12653);
and U12858 (N_12858,N_12511,N_12532);
nor U12859 (N_12859,N_12661,N_12668);
xnor U12860 (N_12860,N_12536,N_12506);
nand U12861 (N_12861,N_12590,N_12519);
or U12862 (N_12862,N_12603,N_12529);
or U12863 (N_12863,N_12554,N_12528);
nor U12864 (N_12864,N_12749,N_12664);
nor U12865 (N_12865,N_12684,N_12574);
or U12866 (N_12866,N_12730,N_12565);
nor U12867 (N_12867,N_12702,N_12579);
and U12868 (N_12868,N_12516,N_12533);
and U12869 (N_12869,N_12546,N_12571);
nor U12870 (N_12870,N_12526,N_12517);
nor U12871 (N_12871,N_12523,N_12744);
and U12872 (N_12872,N_12597,N_12665);
nand U12873 (N_12873,N_12703,N_12606);
nor U12874 (N_12874,N_12666,N_12676);
or U12875 (N_12875,N_12640,N_12520);
and U12876 (N_12876,N_12510,N_12620);
nor U12877 (N_12877,N_12562,N_12678);
nand U12878 (N_12878,N_12510,N_12635);
and U12879 (N_12879,N_12699,N_12632);
nor U12880 (N_12880,N_12589,N_12569);
or U12881 (N_12881,N_12699,N_12623);
nor U12882 (N_12882,N_12652,N_12738);
or U12883 (N_12883,N_12561,N_12646);
or U12884 (N_12884,N_12587,N_12696);
or U12885 (N_12885,N_12742,N_12697);
nand U12886 (N_12886,N_12647,N_12656);
nand U12887 (N_12887,N_12534,N_12696);
and U12888 (N_12888,N_12749,N_12527);
nand U12889 (N_12889,N_12709,N_12518);
nor U12890 (N_12890,N_12509,N_12557);
or U12891 (N_12891,N_12683,N_12739);
or U12892 (N_12892,N_12654,N_12606);
and U12893 (N_12893,N_12711,N_12619);
nand U12894 (N_12894,N_12684,N_12736);
or U12895 (N_12895,N_12622,N_12681);
and U12896 (N_12896,N_12744,N_12702);
nand U12897 (N_12897,N_12527,N_12660);
or U12898 (N_12898,N_12695,N_12500);
nand U12899 (N_12899,N_12743,N_12568);
or U12900 (N_12900,N_12677,N_12732);
nand U12901 (N_12901,N_12720,N_12578);
nor U12902 (N_12902,N_12723,N_12734);
or U12903 (N_12903,N_12504,N_12528);
or U12904 (N_12904,N_12665,N_12549);
nor U12905 (N_12905,N_12520,N_12578);
nand U12906 (N_12906,N_12728,N_12573);
or U12907 (N_12907,N_12640,N_12677);
nor U12908 (N_12908,N_12614,N_12592);
nor U12909 (N_12909,N_12631,N_12723);
or U12910 (N_12910,N_12647,N_12534);
and U12911 (N_12911,N_12719,N_12747);
nand U12912 (N_12912,N_12746,N_12514);
or U12913 (N_12913,N_12669,N_12674);
nor U12914 (N_12914,N_12587,N_12727);
and U12915 (N_12915,N_12571,N_12724);
or U12916 (N_12916,N_12714,N_12692);
or U12917 (N_12917,N_12693,N_12611);
and U12918 (N_12918,N_12510,N_12656);
and U12919 (N_12919,N_12503,N_12664);
nand U12920 (N_12920,N_12705,N_12586);
nand U12921 (N_12921,N_12593,N_12582);
or U12922 (N_12922,N_12706,N_12518);
or U12923 (N_12923,N_12537,N_12541);
or U12924 (N_12924,N_12688,N_12724);
nor U12925 (N_12925,N_12664,N_12655);
and U12926 (N_12926,N_12502,N_12632);
nor U12927 (N_12927,N_12631,N_12564);
and U12928 (N_12928,N_12641,N_12661);
nor U12929 (N_12929,N_12726,N_12723);
or U12930 (N_12930,N_12713,N_12692);
nand U12931 (N_12931,N_12611,N_12729);
or U12932 (N_12932,N_12652,N_12605);
or U12933 (N_12933,N_12748,N_12737);
nor U12934 (N_12934,N_12638,N_12728);
or U12935 (N_12935,N_12712,N_12690);
and U12936 (N_12936,N_12577,N_12574);
nand U12937 (N_12937,N_12748,N_12703);
and U12938 (N_12938,N_12726,N_12531);
or U12939 (N_12939,N_12566,N_12646);
and U12940 (N_12940,N_12653,N_12575);
and U12941 (N_12941,N_12749,N_12685);
nand U12942 (N_12942,N_12644,N_12652);
or U12943 (N_12943,N_12740,N_12697);
xnor U12944 (N_12944,N_12606,N_12504);
and U12945 (N_12945,N_12673,N_12597);
nor U12946 (N_12946,N_12659,N_12573);
nand U12947 (N_12947,N_12530,N_12668);
nand U12948 (N_12948,N_12737,N_12614);
nor U12949 (N_12949,N_12687,N_12583);
nand U12950 (N_12950,N_12649,N_12633);
and U12951 (N_12951,N_12509,N_12572);
nand U12952 (N_12952,N_12557,N_12743);
and U12953 (N_12953,N_12720,N_12666);
or U12954 (N_12954,N_12505,N_12650);
and U12955 (N_12955,N_12558,N_12633);
or U12956 (N_12956,N_12597,N_12565);
and U12957 (N_12957,N_12504,N_12648);
or U12958 (N_12958,N_12504,N_12634);
or U12959 (N_12959,N_12598,N_12737);
and U12960 (N_12960,N_12720,N_12576);
nand U12961 (N_12961,N_12578,N_12591);
and U12962 (N_12962,N_12660,N_12666);
nor U12963 (N_12963,N_12612,N_12724);
nor U12964 (N_12964,N_12580,N_12563);
nand U12965 (N_12965,N_12677,N_12725);
xor U12966 (N_12966,N_12747,N_12718);
and U12967 (N_12967,N_12534,N_12571);
or U12968 (N_12968,N_12633,N_12538);
nand U12969 (N_12969,N_12653,N_12549);
or U12970 (N_12970,N_12531,N_12557);
and U12971 (N_12971,N_12728,N_12515);
nand U12972 (N_12972,N_12627,N_12734);
or U12973 (N_12973,N_12570,N_12695);
and U12974 (N_12974,N_12652,N_12527);
and U12975 (N_12975,N_12685,N_12546);
and U12976 (N_12976,N_12664,N_12519);
and U12977 (N_12977,N_12585,N_12706);
and U12978 (N_12978,N_12657,N_12741);
and U12979 (N_12979,N_12741,N_12648);
or U12980 (N_12980,N_12694,N_12540);
nor U12981 (N_12981,N_12620,N_12653);
and U12982 (N_12982,N_12524,N_12748);
nand U12983 (N_12983,N_12578,N_12645);
and U12984 (N_12984,N_12698,N_12526);
nor U12985 (N_12985,N_12607,N_12722);
and U12986 (N_12986,N_12552,N_12543);
nor U12987 (N_12987,N_12637,N_12730);
and U12988 (N_12988,N_12538,N_12636);
or U12989 (N_12989,N_12512,N_12546);
nand U12990 (N_12990,N_12544,N_12652);
nand U12991 (N_12991,N_12510,N_12742);
nor U12992 (N_12992,N_12530,N_12527);
and U12993 (N_12993,N_12746,N_12609);
nand U12994 (N_12994,N_12549,N_12612);
nor U12995 (N_12995,N_12673,N_12596);
and U12996 (N_12996,N_12560,N_12663);
nor U12997 (N_12997,N_12658,N_12552);
and U12998 (N_12998,N_12532,N_12614);
and U12999 (N_12999,N_12652,N_12637);
nor U13000 (N_13000,N_12800,N_12857);
and U13001 (N_13001,N_12924,N_12834);
nor U13002 (N_13002,N_12768,N_12883);
or U13003 (N_13003,N_12959,N_12961);
or U13004 (N_13004,N_12986,N_12958);
or U13005 (N_13005,N_12921,N_12782);
or U13006 (N_13006,N_12901,N_12797);
nand U13007 (N_13007,N_12822,N_12990);
nor U13008 (N_13008,N_12933,N_12848);
nand U13009 (N_13009,N_12871,N_12981);
nor U13010 (N_13010,N_12855,N_12950);
and U13011 (N_13011,N_12931,N_12932);
nand U13012 (N_13012,N_12841,N_12983);
nor U13013 (N_13013,N_12973,N_12905);
nor U13014 (N_13014,N_12878,N_12977);
or U13015 (N_13015,N_12819,N_12862);
nand U13016 (N_13016,N_12927,N_12964);
nand U13017 (N_13017,N_12787,N_12972);
nor U13018 (N_13018,N_12777,N_12962);
nor U13019 (N_13019,N_12966,N_12791);
nand U13020 (N_13020,N_12827,N_12910);
and U13021 (N_13021,N_12850,N_12849);
nand U13022 (N_13022,N_12833,N_12788);
or U13023 (N_13023,N_12876,N_12913);
nand U13024 (N_13024,N_12836,N_12815);
and U13025 (N_13025,N_12916,N_12997);
nand U13026 (N_13026,N_12999,N_12784);
nor U13027 (N_13027,N_12807,N_12989);
or U13028 (N_13028,N_12953,N_12873);
nor U13029 (N_13029,N_12774,N_12976);
nor U13030 (N_13030,N_12891,N_12904);
or U13031 (N_13031,N_12949,N_12754);
xor U13032 (N_13032,N_12821,N_12914);
or U13033 (N_13033,N_12840,N_12861);
nor U13034 (N_13034,N_12808,N_12872);
nor U13035 (N_13035,N_12847,N_12813);
nor U13036 (N_13036,N_12957,N_12867);
and U13037 (N_13037,N_12943,N_12877);
or U13038 (N_13038,N_12756,N_12942);
and U13039 (N_13039,N_12939,N_12955);
and U13040 (N_13040,N_12929,N_12825);
and U13041 (N_13041,N_12866,N_12810);
nor U13042 (N_13042,N_12856,N_12818);
and U13043 (N_13043,N_12969,N_12900);
nand U13044 (N_13044,N_12814,N_12837);
nand U13045 (N_13045,N_12975,N_12980);
or U13046 (N_13046,N_12766,N_12898);
and U13047 (N_13047,N_12994,N_12895);
nand U13048 (N_13048,N_12824,N_12886);
and U13049 (N_13049,N_12903,N_12854);
nor U13050 (N_13050,N_12792,N_12755);
and U13051 (N_13051,N_12875,N_12859);
nor U13052 (N_13052,N_12770,N_12760);
and U13053 (N_13053,N_12798,N_12993);
nand U13054 (N_13054,N_12839,N_12934);
nor U13055 (N_13055,N_12758,N_12930);
nor U13056 (N_13056,N_12963,N_12965);
nor U13057 (N_13057,N_12759,N_12764);
or U13058 (N_13058,N_12845,N_12945);
and U13059 (N_13059,N_12790,N_12960);
or U13060 (N_13060,N_12820,N_12864);
and U13061 (N_13061,N_12778,N_12796);
nand U13062 (N_13062,N_12880,N_12896);
nor U13063 (N_13063,N_12775,N_12912);
nor U13064 (N_13064,N_12786,N_12938);
or U13065 (N_13065,N_12829,N_12806);
and U13066 (N_13066,N_12885,N_12794);
xnor U13067 (N_13067,N_12751,N_12874);
or U13068 (N_13068,N_12776,N_12893);
nand U13069 (N_13069,N_12838,N_12887);
nand U13070 (N_13070,N_12805,N_12954);
and U13071 (N_13071,N_12920,N_12863);
nor U13072 (N_13072,N_12985,N_12936);
nor U13073 (N_13073,N_12987,N_12998);
or U13074 (N_13074,N_12988,N_12809);
and U13075 (N_13075,N_12982,N_12793);
or U13076 (N_13076,N_12843,N_12851);
nand U13077 (N_13077,N_12889,N_12978);
xnor U13078 (N_13078,N_12860,N_12974);
and U13079 (N_13079,N_12911,N_12937);
or U13080 (N_13080,N_12868,N_12881);
nand U13081 (N_13081,N_12769,N_12923);
nor U13082 (N_13082,N_12842,N_12779);
or U13083 (N_13083,N_12869,N_12879);
or U13084 (N_13084,N_12757,N_12783);
or U13085 (N_13085,N_12795,N_12902);
nand U13086 (N_13086,N_12884,N_12992);
nor U13087 (N_13087,N_12894,N_12811);
or U13088 (N_13088,N_12785,N_12970);
nor U13089 (N_13089,N_12762,N_12773);
nand U13090 (N_13090,N_12812,N_12897);
or U13091 (N_13091,N_12753,N_12832);
nand U13092 (N_13092,N_12761,N_12946);
and U13093 (N_13093,N_12858,N_12804);
and U13094 (N_13094,N_12763,N_12948);
nand U13095 (N_13095,N_12906,N_12853);
nand U13096 (N_13096,N_12951,N_12925);
or U13097 (N_13097,N_12991,N_12908);
nand U13098 (N_13098,N_12928,N_12944);
or U13099 (N_13099,N_12817,N_12940);
and U13100 (N_13100,N_12952,N_12870);
nand U13101 (N_13101,N_12979,N_12967);
nor U13102 (N_13102,N_12899,N_12828);
or U13103 (N_13103,N_12926,N_12802);
or U13104 (N_13104,N_12765,N_12984);
or U13105 (N_13105,N_12772,N_12892);
nor U13106 (N_13106,N_12781,N_12918);
nor U13107 (N_13107,N_12831,N_12907);
nor U13108 (N_13108,N_12780,N_12882);
and U13109 (N_13109,N_12865,N_12995);
nor U13110 (N_13110,N_12844,N_12935);
nor U13111 (N_13111,N_12956,N_12771);
or U13112 (N_13112,N_12852,N_12915);
or U13113 (N_13113,N_12823,N_12917);
and U13114 (N_13114,N_12801,N_12996);
nand U13115 (N_13115,N_12789,N_12767);
or U13116 (N_13116,N_12752,N_12888);
nand U13117 (N_13117,N_12968,N_12830);
xor U13118 (N_13118,N_12816,N_12890);
nor U13119 (N_13119,N_12826,N_12909);
nor U13120 (N_13120,N_12750,N_12922);
nor U13121 (N_13121,N_12803,N_12941);
and U13122 (N_13122,N_12799,N_12971);
nor U13123 (N_13123,N_12947,N_12835);
and U13124 (N_13124,N_12846,N_12919);
nor U13125 (N_13125,N_12823,N_12811);
nor U13126 (N_13126,N_12950,N_12807);
nor U13127 (N_13127,N_12912,N_12942);
and U13128 (N_13128,N_12753,N_12929);
nor U13129 (N_13129,N_12753,N_12785);
nor U13130 (N_13130,N_12846,N_12787);
nor U13131 (N_13131,N_12790,N_12820);
and U13132 (N_13132,N_12995,N_12843);
nor U13133 (N_13133,N_12999,N_12762);
or U13134 (N_13134,N_12784,N_12913);
nor U13135 (N_13135,N_12826,N_12957);
or U13136 (N_13136,N_12895,N_12922);
nand U13137 (N_13137,N_12813,N_12979);
nor U13138 (N_13138,N_12868,N_12871);
or U13139 (N_13139,N_12999,N_12943);
nor U13140 (N_13140,N_12917,N_12797);
nand U13141 (N_13141,N_12771,N_12955);
and U13142 (N_13142,N_12815,N_12847);
nor U13143 (N_13143,N_12887,N_12961);
nand U13144 (N_13144,N_12923,N_12946);
and U13145 (N_13145,N_12906,N_12880);
nor U13146 (N_13146,N_12865,N_12850);
or U13147 (N_13147,N_12922,N_12870);
nor U13148 (N_13148,N_12756,N_12928);
nand U13149 (N_13149,N_12928,N_12765);
nand U13150 (N_13150,N_12929,N_12882);
and U13151 (N_13151,N_12875,N_12861);
nor U13152 (N_13152,N_12965,N_12958);
and U13153 (N_13153,N_12957,N_12990);
nand U13154 (N_13154,N_12865,N_12878);
nor U13155 (N_13155,N_12954,N_12959);
and U13156 (N_13156,N_12936,N_12834);
or U13157 (N_13157,N_12944,N_12958);
or U13158 (N_13158,N_12856,N_12961);
or U13159 (N_13159,N_12802,N_12819);
or U13160 (N_13160,N_12964,N_12962);
or U13161 (N_13161,N_12959,N_12790);
or U13162 (N_13162,N_12983,N_12765);
and U13163 (N_13163,N_12975,N_12751);
or U13164 (N_13164,N_12986,N_12811);
or U13165 (N_13165,N_12804,N_12952);
nand U13166 (N_13166,N_12904,N_12883);
nand U13167 (N_13167,N_12980,N_12781);
nor U13168 (N_13168,N_12902,N_12895);
nand U13169 (N_13169,N_12922,N_12802);
nor U13170 (N_13170,N_12993,N_12808);
nand U13171 (N_13171,N_12892,N_12950);
and U13172 (N_13172,N_12861,N_12761);
nor U13173 (N_13173,N_12783,N_12777);
and U13174 (N_13174,N_12854,N_12821);
and U13175 (N_13175,N_12968,N_12983);
or U13176 (N_13176,N_12837,N_12922);
and U13177 (N_13177,N_12956,N_12801);
or U13178 (N_13178,N_12812,N_12925);
nor U13179 (N_13179,N_12911,N_12793);
nand U13180 (N_13180,N_12971,N_12960);
nor U13181 (N_13181,N_12831,N_12783);
nand U13182 (N_13182,N_12877,N_12909);
and U13183 (N_13183,N_12894,N_12769);
nand U13184 (N_13184,N_12934,N_12950);
or U13185 (N_13185,N_12945,N_12870);
or U13186 (N_13186,N_12983,N_12758);
or U13187 (N_13187,N_12926,N_12782);
or U13188 (N_13188,N_12927,N_12992);
or U13189 (N_13189,N_12871,N_12960);
nor U13190 (N_13190,N_12762,N_12796);
and U13191 (N_13191,N_12862,N_12965);
and U13192 (N_13192,N_12844,N_12987);
and U13193 (N_13193,N_12761,N_12963);
and U13194 (N_13194,N_12924,N_12922);
nor U13195 (N_13195,N_12841,N_12902);
nand U13196 (N_13196,N_12802,N_12848);
or U13197 (N_13197,N_12837,N_12954);
nor U13198 (N_13198,N_12848,N_12761);
nor U13199 (N_13199,N_12833,N_12752);
nand U13200 (N_13200,N_12829,N_12939);
or U13201 (N_13201,N_12945,N_12847);
or U13202 (N_13202,N_12890,N_12914);
nor U13203 (N_13203,N_12801,N_12786);
nand U13204 (N_13204,N_12901,N_12808);
and U13205 (N_13205,N_12897,N_12924);
or U13206 (N_13206,N_12881,N_12758);
nand U13207 (N_13207,N_12885,N_12978);
nor U13208 (N_13208,N_12763,N_12756);
and U13209 (N_13209,N_12862,N_12943);
or U13210 (N_13210,N_12949,N_12898);
or U13211 (N_13211,N_12965,N_12797);
nand U13212 (N_13212,N_12905,N_12930);
and U13213 (N_13213,N_12758,N_12850);
and U13214 (N_13214,N_12757,N_12814);
or U13215 (N_13215,N_12901,N_12822);
or U13216 (N_13216,N_12786,N_12869);
or U13217 (N_13217,N_12894,N_12775);
nor U13218 (N_13218,N_12907,N_12931);
and U13219 (N_13219,N_12836,N_12958);
xnor U13220 (N_13220,N_12815,N_12951);
or U13221 (N_13221,N_12937,N_12824);
nand U13222 (N_13222,N_12939,N_12920);
or U13223 (N_13223,N_12754,N_12923);
nand U13224 (N_13224,N_12862,N_12892);
nand U13225 (N_13225,N_12944,N_12964);
and U13226 (N_13226,N_12893,N_12931);
nor U13227 (N_13227,N_12764,N_12969);
nand U13228 (N_13228,N_12757,N_12867);
and U13229 (N_13229,N_12830,N_12776);
or U13230 (N_13230,N_12930,N_12845);
nor U13231 (N_13231,N_12864,N_12774);
nor U13232 (N_13232,N_12932,N_12923);
or U13233 (N_13233,N_12969,N_12880);
and U13234 (N_13234,N_12789,N_12832);
and U13235 (N_13235,N_12899,N_12915);
and U13236 (N_13236,N_12935,N_12869);
nand U13237 (N_13237,N_12810,N_12794);
and U13238 (N_13238,N_12858,N_12773);
or U13239 (N_13239,N_12973,N_12940);
nor U13240 (N_13240,N_12907,N_12947);
nand U13241 (N_13241,N_12851,N_12908);
xnor U13242 (N_13242,N_12841,N_12979);
nand U13243 (N_13243,N_12822,N_12881);
nor U13244 (N_13244,N_12852,N_12909);
and U13245 (N_13245,N_12925,N_12827);
or U13246 (N_13246,N_12891,N_12825);
nor U13247 (N_13247,N_12819,N_12794);
nor U13248 (N_13248,N_12816,N_12804);
nor U13249 (N_13249,N_12760,N_12887);
and U13250 (N_13250,N_13088,N_13193);
nor U13251 (N_13251,N_13008,N_13199);
and U13252 (N_13252,N_13047,N_13112);
nand U13253 (N_13253,N_13023,N_13078);
or U13254 (N_13254,N_13198,N_13173);
nand U13255 (N_13255,N_13016,N_13242);
or U13256 (N_13256,N_13048,N_13085);
nand U13257 (N_13257,N_13089,N_13209);
or U13258 (N_13258,N_13208,N_13010);
nand U13259 (N_13259,N_13218,N_13144);
nand U13260 (N_13260,N_13015,N_13145);
nand U13261 (N_13261,N_13094,N_13012);
nor U13262 (N_13262,N_13081,N_13196);
nand U13263 (N_13263,N_13003,N_13160);
nand U13264 (N_13264,N_13107,N_13235);
nand U13265 (N_13265,N_13150,N_13245);
or U13266 (N_13266,N_13125,N_13243);
nand U13267 (N_13267,N_13104,N_13131);
or U13268 (N_13268,N_13065,N_13223);
or U13269 (N_13269,N_13040,N_13185);
nand U13270 (N_13270,N_13149,N_13014);
and U13271 (N_13271,N_13049,N_13136);
nand U13272 (N_13272,N_13158,N_13076);
nor U13273 (N_13273,N_13056,N_13117);
nand U13274 (N_13274,N_13063,N_13041);
nand U13275 (N_13275,N_13236,N_13215);
and U13276 (N_13276,N_13122,N_13099);
nor U13277 (N_13277,N_13146,N_13036);
and U13278 (N_13278,N_13133,N_13230);
or U13279 (N_13279,N_13109,N_13226);
and U13280 (N_13280,N_13051,N_13163);
nand U13281 (N_13281,N_13224,N_13046);
or U13282 (N_13282,N_13028,N_13135);
or U13283 (N_13283,N_13141,N_13092);
nand U13284 (N_13284,N_13219,N_13073);
or U13285 (N_13285,N_13210,N_13098);
nand U13286 (N_13286,N_13027,N_13216);
nor U13287 (N_13287,N_13093,N_13152);
nor U13288 (N_13288,N_13241,N_13175);
nand U13289 (N_13289,N_13207,N_13186);
or U13290 (N_13290,N_13102,N_13080);
nor U13291 (N_13291,N_13083,N_13211);
nand U13292 (N_13292,N_13038,N_13164);
nand U13293 (N_13293,N_13134,N_13239);
nor U13294 (N_13294,N_13075,N_13004);
xnor U13295 (N_13295,N_13197,N_13084);
nand U13296 (N_13296,N_13123,N_13189);
nand U13297 (N_13297,N_13222,N_13229);
or U13298 (N_13298,N_13100,N_13184);
nand U13299 (N_13299,N_13037,N_13126);
or U13300 (N_13300,N_13039,N_13113);
nand U13301 (N_13301,N_13005,N_13227);
nand U13302 (N_13302,N_13180,N_13203);
and U13303 (N_13303,N_13139,N_13191);
nand U13304 (N_13304,N_13090,N_13155);
nor U13305 (N_13305,N_13143,N_13082);
nand U13306 (N_13306,N_13029,N_13057);
and U13307 (N_13307,N_13062,N_13194);
nand U13308 (N_13308,N_13086,N_13153);
nor U13309 (N_13309,N_13055,N_13069);
nor U13310 (N_13310,N_13035,N_13032);
nand U13311 (N_13311,N_13238,N_13017);
or U13312 (N_13312,N_13120,N_13091);
nand U13313 (N_13313,N_13240,N_13064);
or U13314 (N_13314,N_13248,N_13244);
nand U13315 (N_13315,N_13011,N_13110);
nor U13316 (N_13316,N_13172,N_13130);
nand U13317 (N_13317,N_13221,N_13054);
or U13318 (N_13318,N_13204,N_13151);
or U13319 (N_13319,N_13116,N_13097);
nand U13320 (N_13320,N_13105,N_13192);
or U13321 (N_13321,N_13019,N_13031);
or U13322 (N_13322,N_13066,N_13181);
nor U13323 (N_13323,N_13095,N_13006);
or U13324 (N_13324,N_13074,N_13231);
or U13325 (N_13325,N_13137,N_13108);
or U13326 (N_13326,N_13068,N_13111);
or U13327 (N_13327,N_13007,N_13161);
nand U13328 (N_13328,N_13079,N_13142);
nand U13329 (N_13329,N_13045,N_13000);
or U13330 (N_13330,N_13183,N_13171);
nand U13331 (N_13331,N_13179,N_13247);
nor U13332 (N_13332,N_13121,N_13138);
and U13333 (N_13333,N_13050,N_13176);
or U13334 (N_13334,N_13106,N_13087);
and U13335 (N_13335,N_13202,N_13170);
nand U13336 (N_13336,N_13190,N_13002);
or U13337 (N_13337,N_13177,N_13220);
and U13338 (N_13338,N_13025,N_13103);
and U13339 (N_13339,N_13234,N_13140);
nand U13340 (N_13340,N_13058,N_13042);
nand U13341 (N_13341,N_13178,N_13206);
and U13342 (N_13342,N_13053,N_13157);
nor U13343 (N_13343,N_13127,N_13043);
nor U13344 (N_13344,N_13059,N_13174);
nand U13345 (N_13345,N_13021,N_13118);
or U13346 (N_13346,N_13115,N_13156);
nand U13347 (N_13347,N_13067,N_13212);
nor U13348 (N_13348,N_13205,N_13060);
or U13349 (N_13349,N_13233,N_13072);
and U13350 (N_13350,N_13132,N_13201);
nand U13351 (N_13351,N_13061,N_13249);
nand U13352 (N_13352,N_13070,N_13148);
nor U13353 (N_13353,N_13165,N_13213);
nand U13354 (N_13354,N_13200,N_13167);
and U13355 (N_13355,N_13217,N_13044);
and U13356 (N_13356,N_13009,N_13147);
and U13357 (N_13357,N_13159,N_13052);
nor U13358 (N_13358,N_13195,N_13071);
and U13359 (N_13359,N_13001,N_13034);
nand U13360 (N_13360,N_13232,N_13214);
nor U13361 (N_13361,N_13182,N_13228);
and U13362 (N_13362,N_13018,N_13129);
and U13363 (N_13363,N_13166,N_13024);
nor U13364 (N_13364,N_13246,N_13237);
nand U13365 (N_13365,N_13101,N_13162);
nand U13366 (N_13366,N_13114,N_13077);
nand U13367 (N_13367,N_13013,N_13188);
or U13368 (N_13368,N_13124,N_13020);
nor U13369 (N_13369,N_13033,N_13154);
xor U13370 (N_13370,N_13022,N_13030);
or U13371 (N_13371,N_13096,N_13187);
nor U13372 (N_13372,N_13026,N_13225);
or U13373 (N_13373,N_13128,N_13169);
nand U13374 (N_13374,N_13168,N_13119);
nor U13375 (N_13375,N_13136,N_13143);
nand U13376 (N_13376,N_13047,N_13170);
nand U13377 (N_13377,N_13231,N_13066);
and U13378 (N_13378,N_13194,N_13065);
nand U13379 (N_13379,N_13095,N_13069);
nor U13380 (N_13380,N_13231,N_13203);
or U13381 (N_13381,N_13151,N_13237);
xnor U13382 (N_13382,N_13036,N_13094);
nor U13383 (N_13383,N_13238,N_13041);
or U13384 (N_13384,N_13160,N_13057);
nor U13385 (N_13385,N_13097,N_13058);
or U13386 (N_13386,N_13190,N_13071);
and U13387 (N_13387,N_13077,N_13116);
nor U13388 (N_13388,N_13206,N_13171);
or U13389 (N_13389,N_13182,N_13177);
nand U13390 (N_13390,N_13146,N_13006);
nor U13391 (N_13391,N_13070,N_13102);
or U13392 (N_13392,N_13142,N_13180);
and U13393 (N_13393,N_13242,N_13109);
nor U13394 (N_13394,N_13211,N_13055);
or U13395 (N_13395,N_13046,N_13003);
or U13396 (N_13396,N_13122,N_13038);
nand U13397 (N_13397,N_13116,N_13178);
nand U13398 (N_13398,N_13195,N_13236);
nor U13399 (N_13399,N_13027,N_13003);
and U13400 (N_13400,N_13054,N_13071);
or U13401 (N_13401,N_13085,N_13151);
nand U13402 (N_13402,N_13028,N_13105);
nor U13403 (N_13403,N_13226,N_13093);
nand U13404 (N_13404,N_13124,N_13162);
nand U13405 (N_13405,N_13057,N_13021);
nand U13406 (N_13406,N_13004,N_13020);
or U13407 (N_13407,N_13150,N_13142);
and U13408 (N_13408,N_13012,N_13183);
or U13409 (N_13409,N_13208,N_13089);
nor U13410 (N_13410,N_13032,N_13034);
nand U13411 (N_13411,N_13114,N_13162);
nor U13412 (N_13412,N_13066,N_13247);
or U13413 (N_13413,N_13066,N_13077);
or U13414 (N_13414,N_13039,N_13092);
or U13415 (N_13415,N_13123,N_13180);
or U13416 (N_13416,N_13102,N_13137);
nor U13417 (N_13417,N_13045,N_13105);
or U13418 (N_13418,N_13016,N_13229);
nand U13419 (N_13419,N_13228,N_13072);
or U13420 (N_13420,N_13055,N_13173);
nand U13421 (N_13421,N_13208,N_13154);
xor U13422 (N_13422,N_13087,N_13093);
nand U13423 (N_13423,N_13074,N_13058);
nor U13424 (N_13424,N_13004,N_13138);
nor U13425 (N_13425,N_13191,N_13096);
nand U13426 (N_13426,N_13022,N_13010);
nor U13427 (N_13427,N_13108,N_13075);
nor U13428 (N_13428,N_13042,N_13121);
and U13429 (N_13429,N_13161,N_13077);
nand U13430 (N_13430,N_13070,N_13014);
or U13431 (N_13431,N_13078,N_13235);
or U13432 (N_13432,N_13085,N_13159);
nand U13433 (N_13433,N_13118,N_13084);
nor U13434 (N_13434,N_13014,N_13154);
nor U13435 (N_13435,N_13112,N_13037);
and U13436 (N_13436,N_13142,N_13146);
or U13437 (N_13437,N_13020,N_13119);
or U13438 (N_13438,N_13224,N_13013);
nor U13439 (N_13439,N_13245,N_13241);
nor U13440 (N_13440,N_13067,N_13122);
nand U13441 (N_13441,N_13221,N_13028);
nand U13442 (N_13442,N_13091,N_13070);
nor U13443 (N_13443,N_13245,N_13133);
nand U13444 (N_13444,N_13019,N_13207);
or U13445 (N_13445,N_13091,N_13185);
nor U13446 (N_13446,N_13076,N_13014);
xnor U13447 (N_13447,N_13015,N_13045);
or U13448 (N_13448,N_13238,N_13175);
xnor U13449 (N_13449,N_13121,N_13031);
and U13450 (N_13450,N_13242,N_13005);
or U13451 (N_13451,N_13003,N_13080);
or U13452 (N_13452,N_13104,N_13241);
nand U13453 (N_13453,N_13033,N_13125);
nand U13454 (N_13454,N_13164,N_13094);
nor U13455 (N_13455,N_13029,N_13085);
nor U13456 (N_13456,N_13110,N_13187);
or U13457 (N_13457,N_13110,N_13125);
or U13458 (N_13458,N_13079,N_13087);
nand U13459 (N_13459,N_13141,N_13245);
and U13460 (N_13460,N_13008,N_13198);
nand U13461 (N_13461,N_13016,N_13033);
nor U13462 (N_13462,N_13002,N_13014);
and U13463 (N_13463,N_13111,N_13027);
nand U13464 (N_13464,N_13130,N_13218);
or U13465 (N_13465,N_13111,N_13127);
and U13466 (N_13466,N_13044,N_13049);
and U13467 (N_13467,N_13158,N_13235);
and U13468 (N_13468,N_13021,N_13025);
nor U13469 (N_13469,N_13124,N_13104);
nor U13470 (N_13470,N_13247,N_13021);
or U13471 (N_13471,N_13191,N_13015);
nor U13472 (N_13472,N_13057,N_13177);
nor U13473 (N_13473,N_13208,N_13235);
or U13474 (N_13474,N_13162,N_13126);
nand U13475 (N_13475,N_13201,N_13188);
and U13476 (N_13476,N_13096,N_13188);
nand U13477 (N_13477,N_13237,N_13075);
or U13478 (N_13478,N_13215,N_13246);
or U13479 (N_13479,N_13031,N_13240);
and U13480 (N_13480,N_13023,N_13006);
or U13481 (N_13481,N_13086,N_13240);
or U13482 (N_13482,N_13102,N_13111);
or U13483 (N_13483,N_13249,N_13248);
and U13484 (N_13484,N_13243,N_13070);
or U13485 (N_13485,N_13054,N_13098);
and U13486 (N_13486,N_13133,N_13187);
nand U13487 (N_13487,N_13154,N_13020);
nand U13488 (N_13488,N_13066,N_13221);
nand U13489 (N_13489,N_13098,N_13172);
and U13490 (N_13490,N_13026,N_13094);
and U13491 (N_13491,N_13078,N_13217);
or U13492 (N_13492,N_13211,N_13077);
nand U13493 (N_13493,N_13200,N_13248);
or U13494 (N_13494,N_13230,N_13195);
and U13495 (N_13495,N_13219,N_13070);
nor U13496 (N_13496,N_13192,N_13138);
or U13497 (N_13497,N_13084,N_13243);
and U13498 (N_13498,N_13103,N_13134);
nor U13499 (N_13499,N_13086,N_13182);
or U13500 (N_13500,N_13274,N_13482);
or U13501 (N_13501,N_13343,N_13497);
and U13502 (N_13502,N_13448,N_13469);
and U13503 (N_13503,N_13321,N_13403);
nand U13504 (N_13504,N_13349,N_13487);
nor U13505 (N_13505,N_13474,N_13422);
nand U13506 (N_13506,N_13444,N_13264);
nand U13507 (N_13507,N_13255,N_13364);
nor U13508 (N_13508,N_13253,N_13362);
nand U13509 (N_13509,N_13367,N_13402);
or U13510 (N_13510,N_13468,N_13436);
nor U13511 (N_13511,N_13407,N_13293);
nor U13512 (N_13512,N_13276,N_13263);
and U13513 (N_13513,N_13479,N_13459);
nand U13514 (N_13514,N_13388,N_13291);
and U13515 (N_13515,N_13330,N_13456);
nor U13516 (N_13516,N_13333,N_13396);
nand U13517 (N_13517,N_13381,N_13438);
nand U13518 (N_13518,N_13372,N_13356);
nor U13519 (N_13519,N_13268,N_13279);
and U13520 (N_13520,N_13376,N_13421);
xor U13521 (N_13521,N_13427,N_13314);
and U13522 (N_13522,N_13383,N_13322);
and U13523 (N_13523,N_13294,N_13281);
nor U13524 (N_13524,N_13411,N_13269);
and U13525 (N_13525,N_13414,N_13347);
and U13526 (N_13526,N_13345,N_13361);
and U13527 (N_13527,N_13471,N_13329);
nand U13528 (N_13528,N_13357,N_13295);
or U13529 (N_13529,N_13405,N_13316);
nor U13530 (N_13530,N_13341,N_13466);
and U13531 (N_13531,N_13297,N_13283);
nor U13532 (N_13532,N_13413,N_13432);
nor U13533 (N_13533,N_13445,N_13284);
or U13534 (N_13534,N_13325,N_13336);
and U13535 (N_13535,N_13429,N_13453);
nor U13536 (N_13536,N_13258,N_13256);
and U13537 (N_13537,N_13373,N_13326);
or U13538 (N_13538,N_13299,N_13420);
nand U13539 (N_13539,N_13398,N_13308);
nor U13540 (N_13540,N_13351,N_13289);
nand U13541 (N_13541,N_13406,N_13476);
or U13542 (N_13542,N_13386,N_13350);
or U13543 (N_13543,N_13337,N_13490);
nor U13544 (N_13544,N_13454,N_13369);
nand U13545 (N_13545,N_13252,N_13491);
nand U13546 (N_13546,N_13377,N_13486);
and U13547 (N_13547,N_13328,N_13404);
or U13548 (N_13548,N_13318,N_13277);
or U13549 (N_13549,N_13465,N_13475);
nand U13550 (N_13550,N_13488,N_13344);
nor U13551 (N_13551,N_13423,N_13495);
nand U13552 (N_13552,N_13499,N_13278);
nor U13553 (N_13553,N_13437,N_13300);
and U13554 (N_13554,N_13484,N_13451);
or U13555 (N_13555,N_13311,N_13266);
and U13556 (N_13556,N_13265,N_13272);
and U13557 (N_13557,N_13287,N_13340);
or U13558 (N_13558,N_13412,N_13324);
nor U13559 (N_13559,N_13320,N_13371);
nand U13560 (N_13560,N_13397,N_13359);
and U13561 (N_13561,N_13342,N_13280);
nand U13562 (N_13562,N_13251,N_13435);
nor U13563 (N_13563,N_13261,N_13393);
nor U13564 (N_13564,N_13260,N_13391);
and U13565 (N_13565,N_13472,N_13307);
nor U13566 (N_13566,N_13313,N_13439);
nand U13567 (N_13567,N_13358,N_13385);
nand U13568 (N_13568,N_13498,N_13494);
nor U13569 (N_13569,N_13426,N_13375);
nand U13570 (N_13570,N_13401,N_13478);
or U13571 (N_13571,N_13262,N_13493);
or U13572 (N_13572,N_13408,N_13433);
nand U13573 (N_13573,N_13400,N_13390);
nor U13574 (N_13574,N_13352,N_13399);
nand U13575 (N_13575,N_13309,N_13440);
or U13576 (N_13576,N_13380,N_13470);
nand U13577 (N_13577,N_13430,N_13424);
or U13578 (N_13578,N_13355,N_13431);
nand U13579 (N_13579,N_13332,N_13441);
or U13580 (N_13580,N_13288,N_13416);
nand U13581 (N_13581,N_13310,N_13461);
or U13582 (N_13582,N_13370,N_13292);
or U13583 (N_13583,N_13473,N_13410);
or U13584 (N_13584,N_13298,N_13374);
nand U13585 (N_13585,N_13418,N_13348);
or U13586 (N_13586,N_13339,N_13387);
nor U13587 (N_13587,N_13346,N_13428);
or U13588 (N_13588,N_13334,N_13290);
and U13589 (N_13589,N_13273,N_13271);
and U13590 (N_13590,N_13389,N_13319);
and U13591 (N_13591,N_13460,N_13382);
or U13592 (N_13592,N_13463,N_13480);
or U13593 (N_13593,N_13306,N_13270);
and U13594 (N_13594,N_13467,N_13312);
or U13595 (N_13595,N_13452,N_13458);
nor U13596 (N_13596,N_13259,N_13415);
or U13597 (N_13597,N_13481,N_13384);
nand U13598 (N_13598,N_13417,N_13305);
or U13599 (N_13599,N_13250,N_13353);
or U13600 (N_13600,N_13483,N_13457);
or U13601 (N_13601,N_13296,N_13363);
and U13602 (N_13602,N_13395,N_13327);
or U13603 (N_13603,N_13378,N_13409);
and U13604 (N_13604,N_13282,N_13335);
or U13605 (N_13605,N_13394,N_13267);
and U13606 (N_13606,N_13323,N_13285);
nor U13607 (N_13607,N_13485,N_13317);
or U13608 (N_13608,N_13489,N_13366);
nor U13609 (N_13609,N_13492,N_13257);
and U13610 (N_13610,N_13419,N_13455);
nand U13611 (N_13611,N_13434,N_13443);
nor U13612 (N_13612,N_13331,N_13360);
nand U13613 (N_13613,N_13450,N_13254);
nor U13614 (N_13614,N_13442,N_13462);
nor U13615 (N_13615,N_13464,N_13379);
and U13616 (N_13616,N_13304,N_13302);
nand U13617 (N_13617,N_13425,N_13392);
nor U13618 (N_13618,N_13368,N_13365);
and U13619 (N_13619,N_13301,N_13303);
or U13620 (N_13620,N_13286,N_13275);
and U13621 (N_13621,N_13354,N_13447);
or U13622 (N_13622,N_13449,N_13338);
or U13623 (N_13623,N_13315,N_13496);
or U13624 (N_13624,N_13477,N_13446);
and U13625 (N_13625,N_13479,N_13367);
nand U13626 (N_13626,N_13377,N_13493);
nor U13627 (N_13627,N_13416,N_13321);
or U13628 (N_13628,N_13274,N_13358);
and U13629 (N_13629,N_13404,N_13449);
or U13630 (N_13630,N_13387,N_13367);
nand U13631 (N_13631,N_13328,N_13335);
or U13632 (N_13632,N_13278,N_13354);
and U13633 (N_13633,N_13317,N_13256);
and U13634 (N_13634,N_13280,N_13408);
nor U13635 (N_13635,N_13485,N_13266);
nor U13636 (N_13636,N_13349,N_13483);
or U13637 (N_13637,N_13417,N_13250);
and U13638 (N_13638,N_13397,N_13264);
and U13639 (N_13639,N_13417,N_13458);
or U13640 (N_13640,N_13348,N_13434);
nor U13641 (N_13641,N_13413,N_13315);
and U13642 (N_13642,N_13455,N_13346);
and U13643 (N_13643,N_13459,N_13381);
and U13644 (N_13644,N_13491,N_13322);
nor U13645 (N_13645,N_13442,N_13259);
and U13646 (N_13646,N_13387,N_13419);
nor U13647 (N_13647,N_13338,N_13286);
or U13648 (N_13648,N_13327,N_13485);
nand U13649 (N_13649,N_13481,N_13296);
or U13650 (N_13650,N_13269,N_13258);
and U13651 (N_13651,N_13485,N_13482);
or U13652 (N_13652,N_13446,N_13493);
or U13653 (N_13653,N_13336,N_13405);
nand U13654 (N_13654,N_13484,N_13380);
nand U13655 (N_13655,N_13443,N_13470);
nand U13656 (N_13656,N_13257,N_13402);
or U13657 (N_13657,N_13375,N_13438);
or U13658 (N_13658,N_13252,N_13272);
xnor U13659 (N_13659,N_13408,N_13288);
and U13660 (N_13660,N_13304,N_13441);
nor U13661 (N_13661,N_13381,N_13367);
xor U13662 (N_13662,N_13490,N_13397);
and U13663 (N_13663,N_13492,N_13414);
nand U13664 (N_13664,N_13499,N_13497);
or U13665 (N_13665,N_13494,N_13264);
nand U13666 (N_13666,N_13324,N_13408);
or U13667 (N_13667,N_13459,N_13366);
nor U13668 (N_13668,N_13351,N_13379);
or U13669 (N_13669,N_13481,N_13257);
or U13670 (N_13670,N_13396,N_13411);
nand U13671 (N_13671,N_13472,N_13355);
nor U13672 (N_13672,N_13496,N_13266);
and U13673 (N_13673,N_13340,N_13289);
nor U13674 (N_13674,N_13464,N_13376);
nand U13675 (N_13675,N_13386,N_13419);
nand U13676 (N_13676,N_13437,N_13431);
nand U13677 (N_13677,N_13426,N_13311);
or U13678 (N_13678,N_13396,N_13480);
or U13679 (N_13679,N_13339,N_13424);
or U13680 (N_13680,N_13324,N_13396);
xor U13681 (N_13681,N_13475,N_13492);
and U13682 (N_13682,N_13285,N_13286);
nor U13683 (N_13683,N_13370,N_13468);
or U13684 (N_13684,N_13351,N_13294);
nor U13685 (N_13685,N_13282,N_13265);
or U13686 (N_13686,N_13338,N_13446);
or U13687 (N_13687,N_13499,N_13332);
nor U13688 (N_13688,N_13399,N_13335);
nand U13689 (N_13689,N_13390,N_13381);
or U13690 (N_13690,N_13409,N_13396);
or U13691 (N_13691,N_13387,N_13481);
and U13692 (N_13692,N_13367,N_13394);
nand U13693 (N_13693,N_13401,N_13316);
and U13694 (N_13694,N_13491,N_13395);
nor U13695 (N_13695,N_13402,N_13356);
and U13696 (N_13696,N_13319,N_13467);
nor U13697 (N_13697,N_13253,N_13475);
and U13698 (N_13698,N_13419,N_13293);
or U13699 (N_13699,N_13278,N_13298);
or U13700 (N_13700,N_13485,N_13359);
nand U13701 (N_13701,N_13492,N_13285);
and U13702 (N_13702,N_13371,N_13410);
nand U13703 (N_13703,N_13406,N_13483);
nand U13704 (N_13704,N_13319,N_13272);
and U13705 (N_13705,N_13289,N_13256);
or U13706 (N_13706,N_13312,N_13419);
nand U13707 (N_13707,N_13323,N_13387);
or U13708 (N_13708,N_13392,N_13489);
nand U13709 (N_13709,N_13444,N_13408);
and U13710 (N_13710,N_13277,N_13448);
or U13711 (N_13711,N_13308,N_13456);
nand U13712 (N_13712,N_13350,N_13315);
and U13713 (N_13713,N_13450,N_13329);
nand U13714 (N_13714,N_13463,N_13499);
and U13715 (N_13715,N_13457,N_13400);
or U13716 (N_13716,N_13470,N_13367);
nor U13717 (N_13717,N_13489,N_13263);
or U13718 (N_13718,N_13349,N_13276);
nor U13719 (N_13719,N_13300,N_13464);
nand U13720 (N_13720,N_13415,N_13278);
nand U13721 (N_13721,N_13442,N_13418);
nor U13722 (N_13722,N_13440,N_13414);
nor U13723 (N_13723,N_13494,N_13280);
nand U13724 (N_13724,N_13321,N_13445);
nand U13725 (N_13725,N_13253,N_13428);
nand U13726 (N_13726,N_13306,N_13272);
nor U13727 (N_13727,N_13367,N_13459);
nand U13728 (N_13728,N_13298,N_13385);
and U13729 (N_13729,N_13375,N_13308);
nand U13730 (N_13730,N_13269,N_13421);
or U13731 (N_13731,N_13495,N_13438);
nand U13732 (N_13732,N_13275,N_13475);
nand U13733 (N_13733,N_13488,N_13448);
nor U13734 (N_13734,N_13278,N_13327);
nand U13735 (N_13735,N_13265,N_13425);
nor U13736 (N_13736,N_13370,N_13427);
nand U13737 (N_13737,N_13352,N_13322);
and U13738 (N_13738,N_13481,N_13458);
and U13739 (N_13739,N_13252,N_13356);
nand U13740 (N_13740,N_13461,N_13428);
and U13741 (N_13741,N_13495,N_13289);
nand U13742 (N_13742,N_13281,N_13443);
nor U13743 (N_13743,N_13411,N_13267);
nor U13744 (N_13744,N_13415,N_13340);
nor U13745 (N_13745,N_13475,N_13252);
nand U13746 (N_13746,N_13291,N_13496);
and U13747 (N_13747,N_13435,N_13290);
or U13748 (N_13748,N_13440,N_13317);
and U13749 (N_13749,N_13439,N_13443);
and U13750 (N_13750,N_13677,N_13748);
and U13751 (N_13751,N_13543,N_13615);
or U13752 (N_13752,N_13676,N_13704);
and U13753 (N_13753,N_13643,N_13728);
and U13754 (N_13754,N_13611,N_13576);
nand U13755 (N_13755,N_13743,N_13687);
nor U13756 (N_13756,N_13563,N_13737);
and U13757 (N_13757,N_13667,N_13551);
or U13758 (N_13758,N_13695,N_13587);
nand U13759 (N_13759,N_13683,N_13568);
nand U13760 (N_13760,N_13678,N_13688);
or U13761 (N_13761,N_13518,N_13719);
nand U13762 (N_13762,N_13682,N_13745);
or U13763 (N_13763,N_13646,N_13545);
or U13764 (N_13764,N_13699,N_13630);
or U13765 (N_13765,N_13685,N_13606);
and U13766 (N_13766,N_13527,N_13625);
nand U13767 (N_13767,N_13746,N_13536);
or U13768 (N_13768,N_13608,N_13555);
or U13769 (N_13769,N_13662,N_13723);
or U13770 (N_13770,N_13668,N_13599);
nand U13771 (N_13771,N_13680,N_13648);
or U13772 (N_13772,N_13727,N_13529);
nor U13773 (N_13773,N_13562,N_13622);
nor U13774 (N_13774,N_13596,N_13550);
or U13775 (N_13775,N_13564,N_13635);
nor U13776 (N_13776,N_13707,N_13526);
and U13777 (N_13777,N_13724,N_13739);
nor U13778 (N_13778,N_13696,N_13552);
and U13779 (N_13779,N_13725,N_13503);
nand U13780 (N_13780,N_13519,N_13560);
and U13781 (N_13781,N_13540,N_13607);
nor U13782 (N_13782,N_13742,N_13617);
nand U13783 (N_13783,N_13506,N_13738);
xor U13784 (N_13784,N_13732,N_13580);
and U13785 (N_13785,N_13525,N_13570);
and U13786 (N_13786,N_13669,N_13666);
or U13787 (N_13787,N_13590,N_13616);
and U13788 (N_13788,N_13722,N_13644);
or U13789 (N_13789,N_13524,N_13647);
nor U13790 (N_13790,N_13694,N_13710);
nor U13791 (N_13791,N_13730,N_13597);
and U13792 (N_13792,N_13749,N_13547);
nor U13793 (N_13793,N_13649,N_13675);
nand U13794 (N_13794,N_13645,N_13595);
and U13795 (N_13795,N_13566,N_13589);
nand U13796 (N_13796,N_13508,N_13631);
and U13797 (N_13797,N_13532,N_13533);
nand U13798 (N_13798,N_13672,N_13714);
nand U13799 (N_13799,N_13613,N_13600);
nor U13800 (N_13800,N_13511,N_13747);
nand U13801 (N_13801,N_13558,N_13656);
and U13802 (N_13802,N_13690,N_13534);
and U13803 (N_13803,N_13548,N_13567);
or U13804 (N_13804,N_13502,N_13627);
and U13805 (N_13805,N_13574,N_13654);
and U13806 (N_13806,N_13584,N_13659);
and U13807 (N_13807,N_13500,N_13740);
and U13808 (N_13808,N_13535,N_13528);
nor U13809 (N_13809,N_13598,N_13701);
and U13810 (N_13810,N_13618,N_13711);
and U13811 (N_13811,N_13572,N_13541);
nand U13812 (N_13812,N_13709,N_13638);
or U13813 (N_13813,N_13619,N_13539);
or U13814 (N_13814,N_13712,N_13542);
nor U13815 (N_13815,N_13544,N_13731);
nor U13816 (N_13816,N_13610,N_13679);
or U13817 (N_13817,N_13639,N_13665);
and U13818 (N_13818,N_13583,N_13706);
nand U13819 (N_13819,N_13593,N_13691);
xnor U13820 (N_13820,N_13581,N_13673);
nor U13821 (N_13821,N_13661,N_13601);
nand U13822 (N_13822,N_13514,N_13650);
and U13823 (N_13823,N_13642,N_13604);
nor U13824 (N_13824,N_13717,N_13605);
and U13825 (N_13825,N_13612,N_13684);
or U13826 (N_13826,N_13586,N_13671);
and U13827 (N_13827,N_13554,N_13523);
nand U13828 (N_13828,N_13674,N_13620);
or U13829 (N_13829,N_13521,N_13693);
nor U13830 (N_13830,N_13628,N_13670);
and U13831 (N_13831,N_13579,N_13713);
and U13832 (N_13832,N_13512,N_13509);
or U13833 (N_13833,N_13556,N_13653);
and U13834 (N_13834,N_13735,N_13708);
nand U13835 (N_13835,N_13741,N_13505);
nor U13836 (N_13836,N_13517,N_13614);
and U13837 (N_13837,N_13510,N_13681);
nor U13838 (N_13838,N_13703,N_13626);
nand U13839 (N_13839,N_13702,N_13507);
or U13840 (N_13840,N_13546,N_13501);
nor U13841 (N_13841,N_13663,N_13522);
nand U13842 (N_13842,N_13585,N_13504);
or U13843 (N_13843,N_13655,N_13591);
and U13844 (N_13844,N_13716,N_13686);
or U13845 (N_13845,N_13515,N_13734);
or U13846 (N_13846,N_13520,N_13603);
nor U13847 (N_13847,N_13629,N_13651);
and U13848 (N_13848,N_13530,N_13559);
and U13849 (N_13849,N_13592,N_13537);
and U13850 (N_13850,N_13729,N_13640);
nand U13851 (N_13851,N_13577,N_13582);
nor U13852 (N_13852,N_13634,N_13652);
nor U13853 (N_13853,N_13633,N_13636);
nand U13854 (N_13854,N_13575,N_13561);
or U13855 (N_13855,N_13573,N_13571);
nor U13856 (N_13856,N_13689,N_13657);
or U13857 (N_13857,N_13538,N_13736);
or U13858 (N_13858,N_13602,N_13660);
or U13859 (N_13859,N_13637,N_13609);
and U13860 (N_13860,N_13733,N_13516);
and U13861 (N_13861,N_13623,N_13692);
nor U13862 (N_13862,N_13594,N_13715);
or U13863 (N_13863,N_13578,N_13744);
nor U13864 (N_13864,N_13698,N_13697);
or U13865 (N_13865,N_13700,N_13588);
nor U13866 (N_13866,N_13726,N_13720);
or U13867 (N_13867,N_13664,N_13705);
nand U13868 (N_13868,N_13624,N_13549);
nor U13869 (N_13869,N_13721,N_13658);
nand U13870 (N_13870,N_13621,N_13569);
or U13871 (N_13871,N_13531,N_13553);
or U13872 (N_13872,N_13565,N_13632);
nor U13873 (N_13873,N_13641,N_13557);
nand U13874 (N_13874,N_13513,N_13718);
xnor U13875 (N_13875,N_13632,N_13621);
or U13876 (N_13876,N_13538,N_13748);
nand U13877 (N_13877,N_13538,N_13637);
or U13878 (N_13878,N_13643,N_13714);
nor U13879 (N_13879,N_13657,N_13717);
nor U13880 (N_13880,N_13603,N_13569);
and U13881 (N_13881,N_13615,N_13561);
nand U13882 (N_13882,N_13617,N_13520);
or U13883 (N_13883,N_13688,N_13536);
nand U13884 (N_13884,N_13555,N_13547);
or U13885 (N_13885,N_13584,N_13743);
nand U13886 (N_13886,N_13624,N_13746);
and U13887 (N_13887,N_13587,N_13690);
and U13888 (N_13888,N_13534,N_13588);
and U13889 (N_13889,N_13665,N_13560);
nor U13890 (N_13890,N_13590,N_13562);
and U13891 (N_13891,N_13616,N_13619);
or U13892 (N_13892,N_13667,N_13660);
and U13893 (N_13893,N_13738,N_13719);
or U13894 (N_13894,N_13677,N_13531);
nand U13895 (N_13895,N_13602,N_13540);
nor U13896 (N_13896,N_13513,N_13573);
nor U13897 (N_13897,N_13590,N_13733);
nand U13898 (N_13898,N_13605,N_13615);
nor U13899 (N_13899,N_13670,N_13500);
nor U13900 (N_13900,N_13675,N_13664);
and U13901 (N_13901,N_13708,N_13630);
nand U13902 (N_13902,N_13697,N_13689);
or U13903 (N_13903,N_13524,N_13666);
nand U13904 (N_13904,N_13648,N_13543);
nand U13905 (N_13905,N_13522,N_13744);
nand U13906 (N_13906,N_13613,N_13719);
and U13907 (N_13907,N_13674,N_13673);
nand U13908 (N_13908,N_13743,N_13574);
or U13909 (N_13909,N_13734,N_13636);
xor U13910 (N_13910,N_13699,N_13745);
and U13911 (N_13911,N_13638,N_13687);
or U13912 (N_13912,N_13542,N_13591);
or U13913 (N_13913,N_13566,N_13730);
nand U13914 (N_13914,N_13622,N_13711);
or U13915 (N_13915,N_13627,N_13739);
and U13916 (N_13916,N_13521,N_13600);
nor U13917 (N_13917,N_13616,N_13594);
and U13918 (N_13918,N_13507,N_13720);
nand U13919 (N_13919,N_13596,N_13701);
nand U13920 (N_13920,N_13692,N_13603);
or U13921 (N_13921,N_13662,N_13713);
and U13922 (N_13922,N_13722,N_13567);
nand U13923 (N_13923,N_13747,N_13717);
nor U13924 (N_13924,N_13744,N_13524);
or U13925 (N_13925,N_13621,N_13534);
nor U13926 (N_13926,N_13708,N_13529);
nor U13927 (N_13927,N_13694,N_13531);
nand U13928 (N_13928,N_13559,N_13543);
nor U13929 (N_13929,N_13723,N_13559);
and U13930 (N_13930,N_13578,N_13594);
nor U13931 (N_13931,N_13718,N_13554);
and U13932 (N_13932,N_13712,N_13637);
nand U13933 (N_13933,N_13515,N_13555);
nand U13934 (N_13934,N_13715,N_13565);
nand U13935 (N_13935,N_13600,N_13726);
nand U13936 (N_13936,N_13616,N_13681);
or U13937 (N_13937,N_13720,N_13724);
and U13938 (N_13938,N_13627,N_13677);
nor U13939 (N_13939,N_13548,N_13602);
nand U13940 (N_13940,N_13723,N_13659);
nand U13941 (N_13941,N_13624,N_13530);
and U13942 (N_13942,N_13566,N_13599);
or U13943 (N_13943,N_13711,N_13673);
or U13944 (N_13944,N_13525,N_13625);
or U13945 (N_13945,N_13663,N_13719);
and U13946 (N_13946,N_13663,N_13656);
or U13947 (N_13947,N_13607,N_13723);
and U13948 (N_13948,N_13516,N_13726);
and U13949 (N_13949,N_13743,N_13677);
nor U13950 (N_13950,N_13651,N_13632);
nor U13951 (N_13951,N_13516,N_13536);
nand U13952 (N_13952,N_13740,N_13737);
nand U13953 (N_13953,N_13676,N_13679);
or U13954 (N_13954,N_13716,N_13628);
nand U13955 (N_13955,N_13559,N_13574);
and U13956 (N_13956,N_13656,N_13639);
nor U13957 (N_13957,N_13738,N_13729);
and U13958 (N_13958,N_13571,N_13567);
xor U13959 (N_13959,N_13737,N_13709);
nor U13960 (N_13960,N_13630,N_13511);
and U13961 (N_13961,N_13562,N_13654);
xor U13962 (N_13962,N_13513,N_13548);
nor U13963 (N_13963,N_13600,N_13657);
and U13964 (N_13964,N_13720,N_13566);
and U13965 (N_13965,N_13617,N_13527);
nand U13966 (N_13966,N_13577,N_13624);
nor U13967 (N_13967,N_13563,N_13717);
nand U13968 (N_13968,N_13724,N_13584);
and U13969 (N_13969,N_13586,N_13514);
or U13970 (N_13970,N_13728,N_13618);
and U13971 (N_13971,N_13571,N_13640);
nand U13972 (N_13972,N_13601,N_13682);
and U13973 (N_13973,N_13720,N_13575);
nand U13974 (N_13974,N_13640,N_13602);
nand U13975 (N_13975,N_13554,N_13649);
and U13976 (N_13976,N_13511,N_13612);
xnor U13977 (N_13977,N_13649,N_13526);
or U13978 (N_13978,N_13637,N_13610);
nand U13979 (N_13979,N_13588,N_13558);
or U13980 (N_13980,N_13622,N_13637);
nand U13981 (N_13981,N_13730,N_13729);
nor U13982 (N_13982,N_13515,N_13657);
nand U13983 (N_13983,N_13682,N_13533);
nand U13984 (N_13984,N_13591,N_13671);
nor U13985 (N_13985,N_13610,N_13531);
or U13986 (N_13986,N_13681,N_13579);
nand U13987 (N_13987,N_13660,N_13683);
or U13988 (N_13988,N_13659,N_13749);
nor U13989 (N_13989,N_13603,N_13522);
nor U13990 (N_13990,N_13536,N_13669);
or U13991 (N_13991,N_13596,N_13710);
nor U13992 (N_13992,N_13690,N_13551);
and U13993 (N_13993,N_13652,N_13621);
and U13994 (N_13994,N_13746,N_13602);
nand U13995 (N_13995,N_13597,N_13552);
nand U13996 (N_13996,N_13690,N_13602);
nor U13997 (N_13997,N_13736,N_13583);
nand U13998 (N_13998,N_13625,N_13629);
nand U13999 (N_13999,N_13682,N_13634);
and U14000 (N_14000,N_13933,N_13848);
and U14001 (N_14001,N_13942,N_13982);
nand U14002 (N_14002,N_13914,N_13964);
and U14003 (N_14003,N_13824,N_13817);
nor U14004 (N_14004,N_13873,N_13918);
nand U14005 (N_14005,N_13758,N_13781);
nand U14006 (N_14006,N_13981,N_13826);
and U14007 (N_14007,N_13892,N_13967);
nand U14008 (N_14008,N_13825,N_13976);
and U14009 (N_14009,N_13943,N_13954);
nor U14010 (N_14010,N_13860,N_13917);
or U14011 (N_14011,N_13957,N_13863);
nor U14012 (N_14012,N_13968,N_13839);
or U14013 (N_14013,N_13805,N_13978);
nor U14014 (N_14014,N_13815,N_13830);
nand U14015 (N_14015,N_13881,N_13799);
and U14016 (N_14016,N_13835,N_13938);
or U14017 (N_14017,N_13973,N_13885);
nand U14018 (N_14018,N_13949,N_13776);
nor U14019 (N_14019,N_13782,N_13762);
or U14020 (N_14020,N_13790,N_13779);
and U14021 (N_14021,N_13864,N_13798);
nand U14022 (N_14022,N_13970,N_13890);
or U14023 (N_14023,N_13979,N_13769);
nor U14024 (N_14024,N_13871,N_13813);
nor U14025 (N_14025,N_13874,N_13834);
nor U14026 (N_14026,N_13953,N_13757);
or U14027 (N_14027,N_13894,N_13876);
and U14028 (N_14028,N_13794,N_13856);
or U14029 (N_14029,N_13906,N_13941);
nand U14030 (N_14030,N_13920,N_13983);
or U14031 (N_14031,N_13755,N_13987);
and U14032 (N_14032,N_13752,N_13924);
nor U14033 (N_14033,N_13935,N_13937);
and U14034 (N_14034,N_13849,N_13851);
nand U14035 (N_14035,N_13930,N_13887);
and U14036 (N_14036,N_13974,N_13903);
nand U14037 (N_14037,N_13934,N_13827);
nor U14038 (N_14038,N_13771,N_13972);
or U14039 (N_14039,N_13988,N_13902);
xor U14040 (N_14040,N_13792,N_13754);
nor U14041 (N_14041,N_13886,N_13785);
nand U14042 (N_14042,N_13872,N_13803);
nor U14043 (N_14043,N_13904,N_13761);
nand U14044 (N_14044,N_13811,N_13927);
and U14045 (N_14045,N_13852,N_13992);
nor U14046 (N_14046,N_13910,N_13801);
nor U14047 (N_14047,N_13911,N_13945);
or U14048 (N_14048,N_13858,N_13932);
xnor U14049 (N_14049,N_13905,N_13908);
or U14050 (N_14050,N_13994,N_13916);
nand U14051 (N_14051,N_13850,N_13922);
nor U14052 (N_14052,N_13763,N_13944);
and U14053 (N_14053,N_13804,N_13962);
nor U14054 (N_14054,N_13808,N_13828);
nor U14055 (N_14055,N_13841,N_13773);
nand U14056 (N_14056,N_13778,N_13888);
and U14057 (N_14057,N_13996,N_13926);
or U14058 (N_14058,N_13961,N_13816);
nand U14059 (N_14059,N_13915,N_13759);
nand U14060 (N_14060,N_13853,N_13931);
nand U14061 (N_14061,N_13950,N_13870);
nand U14062 (N_14062,N_13818,N_13891);
nor U14063 (N_14063,N_13845,N_13963);
nand U14064 (N_14064,N_13819,N_13770);
and U14065 (N_14065,N_13875,N_13907);
and U14066 (N_14066,N_13939,N_13895);
nor U14067 (N_14067,N_13837,N_13857);
or U14068 (N_14068,N_13984,N_13788);
or U14069 (N_14069,N_13766,N_13750);
and U14070 (N_14070,N_13823,N_13767);
and U14071 (N_14071,N_13806,N_13940);
nand U14072 (N_14072,N_13877,N_13847);
and U14073 (N_14073,N_13909,N_13952);
xnor U14074 (N_14074,N_13893,N_13928);
or U14075 (N_14075,N_13969,N_13919);
nand U14076 (N_14076,N_13832,N_13993);
or U14077 (N_14077,N_13786,N_13966);
nand U14078 (N_14078,N_13859,N_13751);
nand U14079 (N_14079,N_13925,N_13768);
and U14080 (N_14080,N_13896,N_13854);
nand U14081 (N_14081,N_13838,N_13866);
nor U14082 (N_14082,N_13772,N_13980);
or U14083 (N_14083,N_13843,N_13884);
nand U14084 (N_14084,N_13869,N_13989);
nand U14085 (N_14085,N_13784,N_13814);
nor U14086 (N_14086,N_13936,N_13883);
or U14087 (N_14087,N_13971,N_13855);
or U14088 (N_14088,N_13990,N_13955);
or U14089 (N_14089,N_13793,N_13946);
nor U14090 (N_14090,N_13960,N_13822);
nor U14091 (N_14091,N_13880,N_13861);
nor U14092 (N_14092,N_13867,N_13956);
or U14093 (N_14093,N_13789,N_13991);
or U14094 (N_14094,N_13878,N_13780);
nor U14095 (N_14095,N_13900,N_13846);
xor U14096 (N_14096,N_13844,N_13840);
and U14097 (N_14097,N_13810,N_13796);
nor U14098 (N_14098,N_13787,N_13842);
nand U14099 (N_14099,N_13901,N_13913);
or U14100 (N_14100,N_13783,N_13897);
nor U14101 (N_14101,N_13929,N_13836);
nor U14102 (N_14102,N_13807,N_13868);
and U14103 (N_14103,N_13753,N_13795);
and U14104 (N_14104,N_13879,N_13948);
nand U14105 (N_14105,N_13882,N_13809);
or U14106 (N_14106,N_13764,N_13898);
nor U14107 (N_14107,N_13862,N_13889);
nor U14108 (N_14108,N_13899,N_13831);
nand U14109 (N_14109,N_13821,N_13923);
nand U14110 (N_14110,N_13958,N_13997);
or U14111 (N_14111,N_13995,N_13777);
or U14112 (N_14112,N_13797,N_13959);
and U14113 (N_14113,N_13985,N_13951);
and U14114 (N_14114,N_13912,N_13965);
or U14115 (N_14115,N_13829,N_13791);
and U14116 (N_14116,N_13775,N_13760);
nor U14117 (N_14117,N_13802,N_13833);
or U14118 (N_14118,N_13975,N_13977);
nor U14119 (N_14119,N_13921,N_13998);
or U14120 (N_14120,N_13812,N_13999);
or U14121 (N_14121,N_13774,N_13986);
nand U14122 (N_14122,N_13947,N_13865);
nor U14123 (N_14123,N_13800,N_13756);
and U14124 (N_14124,N_13765,N_13820);
nand U14125 (N_14125,N_13757,N_13917);
or U14126 (N_14126,N_13860,N_13812);
nor U14127 (N_14127,N_13901,N_13994);
or U14128 (N_14128,N_13768,N_13796);
nand U14129 (N_14129,N_13941,N_13938);
or U14130 (N_14130,N_13776,N_13886);
or U14131 (N_14131,N_13840,N_13935);
nor U14132 (N_14132,N_13846,N_13946);
nor U14133 (N_14133,N_13764,N_13847);
or U14134 (N_14134,N_13764,N_13896);
or U14135 (N_14135,N_13842,N_13941);
or U14136 (N_14136,N_13913,N_13778);
nor U14137 (N_14137,N_13941,N_13781);
nand U14138 (N_14138,N_13755,N_13819);
and U14139 (N_14139,N_13845,N_13842);
nand U14140 (N_14140,N_13764,N_13913);
nand U14141 (N_14141,N_13838,N_13886);
and U14142 (N_14142,N_13831,N_13992);
nor U14143 (N_14143,N_13889,N_13865);
and U14144 (N_14144,N_13861,N_13909);
or U14145 (N_14145,N_13779,N_13914);
and U14146 (N_14146,N_13916,N_13833);
or U14147 (N_14147,N_13857,N_13940);
nor U14148 (N_14148,N_13982,N_13761);
nand U14149 (N_14149,N_13949,N_13940);
or U14150 (N_14150,N_13853,N_13935);
nand U14151 (N_14151,N_13815,N_13905);
and U14152 (N_14152,N_13936,N_13753);
nand U14153 (N_14153,N_13811,N_13842);
nand U14154 (N_14154,N_13982,N_13824);
or U14155 (N_14155,N_13947,N_13931);
nor U14156 (N_14156,N_13924,N_13994);
nand U14157 (N_14157,N_13949,N_13827);
and U14158 (N_14158,N_13827,N_13990);
nand U14159 (N_14159,N_13878,N_13854);
and U14160 (N_14160,N_13824,N_13976);
and U14161 (N_14161,N_13926,N_13877);
or U14162 (N_14162,N_13942,N_13886);
xnor U14163 (N_14163,N_13839,N_13905);
and U14164 (N_14164,N_13999,N_13874);
and U14165 (N_14165,N_13958,N_13992);
and U14166 (N_14166,N_13826,N_13759);
nand U14167 (N_14167,N_13912,N_13829);
nand U14168 (N_14168,N_13750,N_13940);
nand U14169 (N_14169,N_13851,N_13889);
nor U14170 (N_14170,N_13814,N_13988);
nand U14171 (N_14171,N_13798,N_13794);
and U14172 (N_14172,N_13885,N_13768);
and U14173 (N_14173,N_13851,N_13987);
nor U14174 (N_14174,N_13933,N_13898);
and U14175 (N_14175,N_13913,N_13864);
nand U14176 (N_14176,N_13853,N_13920);
nand U14177 (N_14177,N_13800,N_13842);
nor U14178 (N_14178,N_13771,N_13868);
nor U14179 (N_14179,N_13839,N_13860);
nor U14180 (N_14180,N_13813,N_13892);
xnor U14181 (N_14181,N_13952,N_13904);
nor U14182 (N_14182,N_13899,N_13876);
or U14183 (N_14183,N_13938,N_13951);
or U14184 (N_14184,N_13838,N_13970);
and U14185 (N_14185,N_13960,N_13973);
and U14186 (N_14186,N_13892,N_13811);
nand U14187 (N_14187,N_13766,N_13832);
or U14188 (N_14188,N_13762,N_13860);
and U14189 (N_14189,N_13880,N_13796);
or U14190 (N_14190,N_13890,N_13886);
and U14191 (N_14191,N_13980,N_13777);
or U14192 (N_14192,N_13814,N_13817);
or U14193 (N_14193,N_13755,N_13809);
nand U14194 (N_14194,N_13998,N_13896);
and U14195 (N_14195,N_13901,N_13947);
nand U14196 (N_14196,N_13859,N_13997);
nor U14197 (N_14197,N_13992,N_13757);
xnor U14198 (N_14198,N_13981,N_13775);
xor U14199 (N_14199,N_13838,N_13948);
and U14200 (N_14200,N_13817,N_13978);
and U14201 (N_14201,N_13933,N_13880);
and U14202 (N_14202,N_13863,N_13882);
and U14203 (N_14203,N_13769,N_13949);
or U14204 (N_14204,N_13768,N_13923);
and U14205 (N_14205,N_13765,N_13863);
nand U14206 (N_14206,N_13789,N_13936);
nor U14207 (N_14207,N_13889,N_13876);
nor U14208 (N_14208,N_13804,N_13974);
nor U14209 (N_14209,N_13780,N_13999);
or U14210 (N_14210,N_13888,N_13905);
nor U14211 (N_14211,N_13858,N_13907);
and U14212 (N_14212,N_13765,N_13968);
and U14213 (N_14213,N_13995,N_13955);
nor U14214 (N_14214,N_13860,N_13863);
nand U14215 (N_14215,N_13869,N_13876);
nor U14216 (N_14216,N_13755,N_13797);
or U14217 (N_14217,N_13897,N_13928);
nand U14218 (N_14218,N_13947,N_13838);
and U14219 (N_14219,N_13777,N_13779);
nand U14220 (N_14220,N_13848,N_13908);
xor U14221 (N_14221,N_13894,N_13828);
or U14222 (N_14222,N_13956,N_13969);
or U14223 (N_14223,N_13937,N_13871);
or U14224 (N_14224,N_13930,N_13799);
nand U14225 (N_14225,N_13755,N_13991);
nor U14226 (N_14226,N_13966,N_13764);
nand U14227 (N_14227,N_13992,N_13892);
nand U14228 (N_14228,N_13764,N_13809);
nor U14229 (N_14229,N_13853,N_13896);
nor U14230 (N_14230,N_13944,N_13777);
or U14231 (N_14231,N_13985,N_13982);
nor U14232 (N_14232,N_13803,N_13796);
nor U14233 (N_14233,N_13812,N_13824);
nor U14234 (N_14234,N_13955,N_13758);
or U14235 (N_14235,N_13891,N_13895);
nand U14236 (N_14236,N_13883,N_13853);
nor U14237 (N_14237,N_13967,N_13877);
nor U14238 (N_14238,N_13984,N_13935);
or U14239 (N_14239,N_13952,N_13757);
or U14240 (N_14240,N_13999,N_13792);
or U14241 (N_14241,N_13852,N_13954);
or U14242 (N_14242,N_13989,N_13852);
nand U14243 (N_14243,N_13819,N_13756);
or U14244 (N_14244,N_13926,N_13979);
nor U14245 (N_14245,N_13840,N_13948);
and U14246 (N_14246,N_13900,N_13779);
nor U14247 (N_14247,N_13834,N_13846);
and U14248 (N_14248,N_13958,N_13887);
or U14249 (N_14249,N_13830,N_13993);
and U14250 (N_14250,N_14185,N_14196);
and U14251 (N_14251,N_14164,N_14184);
and U14252 (N_14252,N_14205,N_14135);
nand U14253 (N_14253,N_14062,N_14230);
nand U14254 (N_14254,N_14109,N_14031);
nor U14255 (N_14255,N_14066,N_14040);
or U14256 (N_14256,N_14224,N_14226);
xnor U14257 (N_14257,N_14092,N_14200);
and U14258 (N_14258,N_14064,N_14042);
nand U14259 (N_14259,N_14228,N_14059);
or U14260 (N_14260,N_14005,N_14156);
and U14261 (N_14261,N_14246,N_14094);
and U14262 (N_14262,N_14247,N_14098);
nand U14263 (N_14263,N_14133,N_14089);
or U14264 (N_14264,N_14183,N_14151);
nor U14265 (N_14265,N_14242,N_14145);
nand U14266 (N_14266,N_14154,N_14087);
nand U14267 (N_14267,N_14063,N_14174);
nand U14268 (N_14268,N_14225,N_14248);
nor U14269 (N_14269,N_14188,N_14144);
or U14270 (N_14270,N_14061,N_14152);
nor U14271 (N_14271,N_14167,N_14049);
or U14272 (N_14272,N_14020,N_14051);
and U14273 (N_14273,N_14153,N_14060);
xnor U14274 (N_14274,N_14065,N_14026);
and U14275 (N_14275,N_14025,N_14076);
nand U14276 (N_14276,N_14028,N_14068);
nand U14277 (N_14277,N_14053,N_14155);
xnor U14278 (N_14278,N_14018,N_14198);
or U14279 (N_14279,N_14127,N_14004);
or U14280 (N_14280,N_14173,N_14084);
nor U14281 (N_14281,N_14107,N_14178);
nand U14282 (N_14282,N_14123,N_14052);
nand U14283 (N_14283,N_14180,N_14222);
nor U14284 (N_14284,N_14148,N_14176);
nand U14285 (N_14285,N_14027,N_14234);
nand U14286 (N_14286,N_14015,N_14012);
and U14287 (N_14287,N_14067,N_14044);
nor U14288 (N_14288,N_14146,N_14165);
and U14289 (N_14289,N_14050,N_14209);
nor U14290 (N_14290,N_14233,N_14172);
and U14291 (N_14291,N_14048,N_14116);
or U14292 (N_14292,N_14002,N_14022);
or U14293 (N_14293,N_14217,N_14216);
nor U14294 (N_14294,N_14212,N_14021);
nor U14295 (N_14295,N_14079,N_14006);
nor U14296 (N_14296,N_14083,N_14220);
nor U14297 (N_14297,N_14110,N_14097);
and U14298 (N_14298,N_14124,N_14175);
nand U14299 (N_14299,N_14128,N_14186);
and U14300 (N_14300,N_14147,N_14204);
nand U14301 (N_14301,N_14125,N_14088);
and U14302 (N_14302,N_14126,N_14150);
nand U14303 (N_14303,N_14108,N_14029);
nand U14304 (N_14304,N_14041,N_14137);
nor U14305 (N_14305,N_14010,N_14192);
nand U14306 (N_14306,N_14245,N_14101);
and U14307 (N_14307,N_14111,N_14009);
and U14308 (N_14308,N_14170,N_14054);
or U14309 (N_14309,N_14055,N_14160);
and U14310 (N_14310,N_14240,N_14117);
nor U14311 (N_14311,N_14078,N_14187);
nand U14312 (N_14312,N_14034,N_14007);
nand U14313 (N_14313,N_14115,N_14024);
and U14314 (N_14314,N_14077,N_14102);
nand U14315 (N_14315,N_14195,N_14096);
nand U14316 (N_14316,N_14249,N_14139);
nor U14317 (N_14317,N_14001,N_14014);
and U14318 (N_14318,N_14000,N_14043);
or U14319 (N_14319,N_14073,N_14169);
nand U14320 (N_14320,N_14244,N_14243);
or U14321 (N_14321,N_14069,N_14210);
nor U14322 (N_14322,N_14238,N_14016);
and U14323 (N_14323,N_14211,N_14229);
and U14324 (N_14324,N_14072,N_14219);
and U14325 (N_14325,N_14231,N_14189);
nand U14326 (N_14326,N_14168,N_14190);
and U14327 (N_14327,N_14100,N_14104);
nor U14328 (N_14328,N_14199,N_14038);
or U14329 (N_14329,N_14112,N_14149);
nor U14330 (N_14330,N_14213,N_14138);
and U14331 (N_14331,N_14099,N_14120);
nor U14332 (N_14332,N_14207,N_14227);
nor U14333 (N_14333,N_14134,N_14136);
nor U14334 (N_14334,N_14235,N_14118);
or U14335 (N_14335,N_14241,N_14158);
nand U14336 (N_14336,N_14141,N_14106);
and U14337 (N_14337,N_14159,N_14223);
or U14338 (N_14338,N_14208,N_14019);
nor U14339 (N_14339,N_14215,N_14103);
nand U14340 (N_14340,N_14030,N_14131);
nor U14341 (N_14341,N_14095,N_14003);
nand U14342 (N_14342,N_14203,N_14157);
and U14343 (N_14343,N_14114,N_14090);
nand U14344 (N_14344,N_14194,N_14070);
and U14345 (N_14345,N_14237,N_14129);
or U14346 (N_14346,N_14082,N_14075);
nor U14347 (N_14347,N_14023,N_14093);
and U14348 (N_14348,N_14011,N_14081);
or U14349 (N_14349,N_14085,N_14056);
or U14350 (N_14350,N_14197,N_14166);
or U14351 (N_14351,N_14130,N_14140);
nand U14352 (N_14352,N_14119,N_14091);
and U14353 (N_14353,N_14037,N_14163);
and U14354 (N_14354,N_14218,N_14071);
nor U14355 (N_14355,N_14142,N_14013);
nand U14356 (N_14356,N_14161,N_14171);
and U14357 (N_14357,N_14201,N_14121);
and U14358 (N_14358,N_14105,N_14177);
or U14359 (N_14359,N_14008,N_14143);
nand U14360 (N_14360,N_14221,N_14057);
nor U14361 (N_14361,N_14179,N_14113);
nand U14362 (N_14362,N_14047,N_14086);
and U14363 (N_14363,N_14046,N_14191);
nand U14364 (N_14364,N_14239,N_14039);
or U14365 (N_14365,N_14162,N_14182);
or U14366 (N_14366,N_14045,N_14035);
nor U14367 (N_14367,N_14181,N_14033);
and U14368 (N_14368,N_14058,N_14232);
or U14369 (N_14369,N_14032,N_14132);
nand U14370 (N_14370,N_14193,N_14202);
nor U14371 (N_14371,N_14074,N_14080);
nor U14372 (N_14372,N_14214,N_14206);
nand U14373 (N_14373,N_14017,N_14036);
nand U14374 (N_14374,N_14236,N_14122);
or U14375 (N_14375,N_14030,N_14214);
nor U14376 (N_14376,N_14130,N_14025);
or U14377 (N_14377,N_14022,N_14015);
nor U14378 (N_14378,N_14008,N_14081);
and U14379 (N_14379,N_14032,N_14228);
nor U14380 (N_14380,N_14080,N_14014);
nand U14381 (N_14381,N_14023,N_14152);
nor U14382 (N_14382,N_14226,N_14117);
or U14383 (N_14383,N_14210,N_14096);
nand U14384 (N_14384,N_14183,N_14198);
or U14385 (N_14385,N_14215,N_14115);
or U14386 (N_14386,N_14127,N_14171);
or U14387 (N_14387,N_14233,N_14053);
nor U14388 (N_14388,N_14034,N_14053);
and U14389 (N_14389,N_14080,N_14127);
nor U14390 (N_14390,N_14065,N_14145);
or U14391 (N_14391,N_14166,N_14233);
and U14392 (N_14392,N_14243,N_14235);
and U14393 (N_14393,N_14021,N_14147);
or U14394 (N_14394,N_14049,N_14215);
or U14395 (N_14395,N_14132,N_14161);
or U14396 (N_14396,N_14207,N_14223);
nor U14397 (N_14397,N_14222,N_14138);
or U14398 (N_14398,N_14165,N_14169);
nor U14399 (N_14399,N_14227,N_14217);
and U14400 (N_14400,N_14220,N_14143);
nor U14401 (N_14401,N_14244,N_14034);
or U14402 (N_14402,N_14079,N_14179);
nand U14403 (N_14403,N_14144,N_14242);
or U14404 (N_14404,N_14162,N_14061);
or U14405 (N_14405,N_14177,N_14166);
or U14406 (N_14406,N_14233,N_14005);
nor U14407 (N_14407,N_14008,N_14134);
nor U14408 (N_14408,N_14013,N_14164);
xor U14409 (N_14409,N_14211,N_14055);
or U14410 (N_14410,N_14210,N_14101);
nand U14411 (N_14411,N_14221,N_14123);
nand U14412 (N_14412,N_14054,N_14179);
xnor U14413 (N_14413,N_14161,N_14124);
and U14414 (N_14414,N_14044,N_14051);
or U14415 (N_14415,N_14165,N_14084);
or U14416 (N_14416,N_14096,N_14017);
nand U14417 (N_14417,N_14170,N_14114);
nand U14418 (N_14418,N_14240,N_14036);
nand U14419 (N_14419,N_14171,N_14049);
nor U14420 (N_14420,N_14098,N_14024);
nor U14421 (N_14421,N_14040,N_14003);
and U14422 (N_14422,N_14082,N_14021);
and U14423 (N_14423,N_14059,N_14171);
nor U14424 (N_14424,N_14217,N_14155);
nand U14425 (N_14425,N_14150,N_14211);
nand U14426 (N_14426,N_14079,N_14243);
or U14427 (N_14427,N_14214,N_14084);
nor U14428 (N_14428,N_14119,N_14227);
or U14429 (N_14429,N_14016,N_14079);
nand U14430 (N_14430,N_14174,N_14098);
nor U14431 (N_14431,N_14025,N_14221);
or U14432 (N_14432,N_14023,N_14248);
xor U14433 (N_14433,N_14050,N_14084);
or U14434 (N_14434,N_14048,N_14247);
nand U14435 (N_14435,N_14085,N_14039);
nor U14436 (N_14436,N_14191,N_14144);
xnor U14437 (N_14437,N_14028,N_14029);
and U14438 (N_14438,N_14036,N_14142);
and U14439 (N_14439,N_14053,N_14100);
nand U14440 (N_14440,N_14124,N_14230);
nand U14441 (N_14441,N_14208,N_14197);
and U14442 (N_14442,N_14011,N_14019);
or U14443 (N_14443,N_14020,N_14093);
nand U14444 (N_14444,N_14120,N_14004);
nand U14445 (N_14445,N_14166,N_14173);
nand U14446 (N_14446,N_14104,N_14114);
or U14447 (N_14447,N_14171,N_14091);
and U14448 (N_14448,N_14249,N_14060);
and U14449 (N_14449,N_14169,N_14023);
nor U14450 (N_14450,N_14062,N_14057);
xnor U14451 (N_14451,N_14030,N_14046);
or U14452 (N_14452,N_14094,N_14089);
and U14453 (N_14453,N_14121,N_14051);
nor U14454 (N_14454,N_14221,N_14237);
nand U14455 (N_14455,N_14085,N_14185);
nor U14456 (N_14456,N_14188,N_14243);
and U14457 (N_14457,N_14114,N_14164);
and U14458 (N_14458,N_14187,N_14237);
and U14459 (N_14459,N_14177,N_14107);
nand U14460 (N_14460,N_14130,N_14191);
or U14461 (N_14461,N_14178,N_14093);
nand U14462 (N_14462,N_14211,N_14136);
nor U14463 (N_14463,N_14163,N_14190);
nor U14464 (N_14464,N_14199,N_14246);
nor U14465 (N_14465,N_14060,N_14121);
nand U14466 (N_14466,N_14160,N_14065);
and U14467 (N_14467,N_14051,N_14058);
nand U14468 (N_14468,N_14053,N_14104);
nand U14469 (N_14469,N_14165,N_14143);
nand U14470 (N_14470,N_14107,N_14048);
or U14471 (N_14471,N_14184,N_14226);
and U14472 (N_14472,N_14235,N_14023);
and U14473 (N_14473,N_14187,N_14208);
or U14474 (N_14474,N_14140,N_14129);
or U14475 (N_14475,N_14008,N_14068);
nand U14476 (N_14476,N_14019,N_14213);
or U14477 (N_14477,N_14176,N_14011);
nand U14478 (N_14478,N_14163,N_14140);
or U14479 (N_14479,N_14165,N_14038);
or U14480 (N_14480,N_14184,N_14035);
nand U14481 (N_14481,N_14155,N_14168);
and U14482 (N_14482,N_14202,N_14207);
nand U14483 (N_14483,N_14239,N_14001);
nand U14484 (N_14484,N_14148,N_14069);
nand U14485 (N_14485,N_14043,N_14040);
nor U14486 (N_14486,N_14080,N_14175);
and U14487 (N_14487,N_14107,N_14157);
and U14488 (N_14488,N_14135,N_14038);
or U14489 (N_14489,N_14107,N_14074);
and U14490 (N_14490,N_14050,N_14069);
nand U14491 (N_14491,N_14199,N_14216);
nor U14492 (N_14492,N_14053,N_14179);
nor U14493 (N_14493,N_14111,N_14002);
nand U14494 (N_14494,N_14049,N_14045);
nand U14495 (N_14495,N_14167,N_14229);
or U14496 (N_14496,N_14066,N_14097);
or U14497 (N_14497,N_14234,N_14219);
or U14498 (N_14498,N_14017,N_14107);
nand U14499 (N_14499,N_14232,N_14186);
and U14500 (N_14500,N_14370,N_14356);
or U14501 (N_14501,N_14255,N_14353);
nand U14502 (N_14502,N_14482,N_14374);
and U14503 (N_14503,N_14418,N_14253);
or U14504 (N_14504,N_14360,N_14382);
or U14505 (N_14505,N_14389,N_14423);
nand U14506 (N_14506,N_14419,N_14409);
or U14507 (N_14507,N_14266,N_14471);
xnor U14508 (N_14508,N_14256,N_14422);
nor U14509 (N_14509,N_14348,N_14481);
nand U14510 (N_14510,N_14317,N_14289);
xor U14511 (N_14511,N_14478,N_14371);
or U14512 (N_14512,N_14341,N_14414);
nand U14513 (N_14513,N_14495,N_14456);
and U14514 (N_14514,N_14251,N_14438);
or U14515 (N_14515,N_14489,N_14428);
nor U14516 (N_14516,N_14391,N_14402);
and U14517 (N_14517,N_14291,N_14430);
and U14518 (N_14518,N_14375,N_14257);
nand U14519 (N_14519,N_14448,N_14497);
nand U14520 (N_14520,N_14315,N_14258);
and U14521 (N_14521,N_14318,N_14493);
and U14522 (N_14522,N_14339,N_14297);
and U14523 (N_14523,N_14275,N_14465);
or U14524 (N_14524,N_14477,N_14436);
and U14525 (N_14525,N_14343,N_14377);
nand U14526 (N_14526,N_14264,N_14321);
and U14527 (N_14527,N_14250,N_14499);
nor U14528 (N_14528,N_14399,N_14309);
or U14529 (N_14529,N_14474,N_14486);
or U14530 (N_14530,N_14384,N_14447);
and U14531 (N_14531,N_14342,N_14420);
and U14532 (N_14532,N_14269,N_14329);
and U14533 (N_14533,N_14451,N_14293);
and U14534 (N_14534,N_14398,N_14458);
nand U14535 (N_14535,N_14330,N_14312);
and U14536 (N_14536,N_14473,N_14431);
or U14537 (N_14537,N_14461,N_14305);
nand U14538 (N_14538,N_14437,N_14443);
and U14539 (N_14539,N_14441,N_14401);
nand U14540 (N_14540,N_14310,N_14386);
and U14541 (N_14541,N_14316,N_14280);
nand U14542 (N_14542,N_14369,N_14426);
nor U14543 (N_14543,N_14262,N_14453);
nand U14544 (N_14544,N_14252,N_14279);
or U14545 (N_14545,N_14479,N_14427);
and U14546 (N_14546,N_14333,N_14492);
and U14547 (N_14547,N_14494,N_14350);
and U14548 (N_14548,N_14281,N_14366);
or U14549 (N_14549,N_14332,N_14496);
and U14550 (N_14550,N_14404,N_14285);
nand U14551 (N_14551,N_14484,N_14302);
and U14552 (N_14552,N_14439,N_14480);
nand U14553 (N_14553,N_14292,N_14372);
nand U14554 (N_14554,N_14299,N_14307);
or U14555 (N_14555,N_14467,N_14286);
nand U14556 (N_14556,N_14425,N_14429);
nand U14557 (N_14557,N_14271,N_14290);
and U14558 (N_14558,N_14254,N_14335);
and U14559 (N_14559,N_14485,N_14282);
nor U14560 (N_14560,N_14328,N_14294);
nand U14561 (N_14561,N_14381,N_14403);
nand U14562 (N_14562,N_14476,N_14354);
nor U14563 (N_14563,N_14413,N_14488);
nor U14564 (N_14564,N_14452,N_14411);
nor U14565 (N_14565,N_14393,N_14337);
or U14566 (N_14566,N_14498,N_14278);
nand U14567 (N_14567,N_14388,N_14346);
nand U14568 (N_14568,N_14440,N_14490);
nand U14569 (N_14569,N_14487,N_14373);
nor U14570 (N_14570,N_14324,N_14340);
nand U14571 (N_14571,N_14390,N_14455);
and U14572 (N_14572,N_14379,N_14460);
and U14573 (N_14573,N_14338,N_14412);
xnor U14574 (N_14574,N_14415,N_14394);
or U14575 (N_14575,N_14334,N_14259);
or U14576 (N_14576,N_14378,N_14367);
or U14577 (N_14577,N_14470,N_14416);
or U14578 (N_14578,N_14311,N_14261);
nor U14579 (N_14579,N_14450,N_14433);
or U14580 (N_14580,N_14263,N_14469);
or U14581 (N_14581,N_14344,N_14365);
nand U14582 (N_14582,N_14323,N_14421);
and U14583 (N_14583,N_14385,N_14319);
nor U14584 (N_14584,N_14444,N_14395);
or U14585 (N_14585,N_14359,N_14368);
nand U14586 (N_14586,N_14442,N_14272);
nand U14587 (N_14587,N_14265,N_14468);
nor U14588 (N_14588,N_14424,N_14417);
nor U14589 (N_14589,N_14407,N_14376);
and U14590 (N_14590,N_14273,N_14462);
xnor U14591 (N_14591,N_14432,N_14464);
or U14592 (N_14592,N_14288,N_14313);
nor U14593 (N_14593,N_14397,N_14274);
nand U14594 (N_14594,N_14459,N_14466);
and U14595 (N_14595,N_14295,N_14301);
and U14596 (N_14596,N_14277,N_14320);
and U14597 (N_14597,N_14408,N_14383);
and U14598 (N_14598,N_14362,N_14349);
nor U14599 (N_14599,N_14364,N_14276);
and U14600 (N_14600,N_14325,N_14267);
nor U14601 (N_14601,N_14435,N_14352);
nand U14602 (N_14602,N_14306,N_14457);
or U14603 (N_14603,N_14405,N_14284);
or U14604 (N_14604,N_14314,N_14434);
or U14605 (N_14605,N_14303,N_14351);
or U14606 (N_14606,N_14283,N_14300);
nand U14607 (N_14607,N_14445,N_14410);
nand U14608 (N_14608,N_14406,N_14472);
and U14609 (N_14609,N_14268,N_14347);
nand U14610 (N_14610,N_14326,N_14483);
xor U14611 (N_14611,N_14331,N_14400);
nand U14612 (N_14612,N_14358,N_14308);
nor U14613 (N_14613,N_14363,N_14449);
or U14614 (N_14614,N_14260,N_14287);
or U14615 (N_14615,N_14392,N_14345);
nor U14616 (N_14616,N_14298,N_14380);
nor U14617 (N_14617,N_14454,N_14475);
nor U14618 (N_14618,N_14446,N_14491);
nand U14619 (N_14619,N_14463,N_14357);
and U14620 (N_14620,N_14327,N_14322);
nor U14621 (N_14621,N_14355,N_14387);
nand U14622 (N_14622,N_14396,N_14296);
nand U14623 (N_14623,N_14336,N_14361);
nand U14624 (N_14624,N_14270,N_14304);
and U14625 (N_14625,N_14404,N_14337);
nand U14626 (N_14626,N_14258,N_14338);
nand U14627 (N_14627,N_14312,N_14372);
xor U14628 (N_14628,N_14364,N_14297);
nand U14629 (N_14629,N_14462,N_14309);
nand U14630 (N_14630,N_14426,N_14455);
or U14631 (N_14631,N_14296,N_14410);
nor U14632 (N_14632,N_14414,N_14340);
and U14633 (N_14633,N_14339,N_14450);
nand U14634 (N_14634,N_14465,N_14311);
nor U14635 (N_14635,N_14428,N_14466);
nor U14636 (N_14636,N_14353,N_14392);
or U14637 (N_14637,N_14466,N_14286);
nand U14638 (N_14638,N_14409,N_14330);
nand U14639 (N_14639,N_14277,N_14474);
nor U14640 (N_14640,N_14252,N_14463);
nand U14641 (N_14641,N_14251,N_14259);
nand U14642 (N_14642,N_14441,N_14455);
nor U14643 (N_14643,N_14279,N_14406);
nor U14644 (N_14644,N_14255,N_14486);
nand U14645 (N_14645,N_14433,N_14345);
or U14646 (N_14646,N_14355,N_14415);
and U14647 (N_14647,N_14313,N_14417);
and U14648 (N_14648,N_14405,N_14268);
nor U14649 (N_14649,N_14390,N_14395);
nand U14650 (N_14650,N_14495,N_14275);
nor U14651 (N_14651,N_14382,N_14497);
nand U14652 (N_14652,N_14416,N_14436);
or U14653 (N_14653,N_14283,N_14281);
nand U14654 (N_14654,N_14436,N_14297);
or U14655 (N_14655,N_14307,N_14366);
nor U14656 (N_14656,N_14395,N_14251);
nor U14657 (N_14657,N_14315,N_14262);
and U14658 (N_14658,N_14383,N_14332);
nor U14659 (N_14659,N_14426,N_14393);
and U14660 (N_14660,N_14261,N_14432);
and U14661 (N_14661,N_14346,N_14485);
nor U14662 (N_14662,N_14323,N_14355);
or U14663 (N_14663,N_14381,N_14278);
nand U14664 (N_14664,N_14445,N_14481);
and U14665 (N_14665,N_14383,N_14354);
and U14666 (N_14666,N_14474,N_14310);
and U14667 (N_14667,N_14338,N_14377);
nor U14668 (N_14668,N_14284,N_14423);
nor U14669 (N_14669,N_14478,N_14463);
or U14670 (N_14670,N_14481,N_14474);
nand U14671 (N_14671,N_14322,N_14461);
and U14672 (N_14672,N_14351,N_14265);
and U14673 (N_14673,N_14379,N_14466);
nor U14674 (N_14674,N_14383,N_14392);
and U14675 (N_14675,N_14279,N_14388);
nor U14676 (N_14676,N_14440,N_14381);
or U14677 (N_14677,N_14485,N_14318);
and U14678 (N_14678,N_14408,N_14371);
nand U14679 (N_14679,N_14492,N_14462);
and U14680 (N_14680,N_14260,N_14366);
or U14681 (N_14681,N_14471,N_14454);
or U14682 (N_14682,N_14351,N_14492);
or U14683 (N_14683,N_14450,N_14400);
nor U14684 (N_14684,N_14406,N_14300);
and U14685 (N_14685,N_14465,N_14285);
and U14686 (N_14686,N_14494,N_14434);
nand U14687 (N_14687,N_14314,N_14432);
nor U14688 (N_14688,N_14402,N_14300);
or U14689 (N_14689,N_14445,N_14289);
and U14690 (N_14690,N_14392,N_14430);
and U14691 (N_14691,N_14349,N_14466);
nor U14692 (N_14692,N_14409,N_14311);
or U14693 (N_14693,N_14426,N_14321);
and U14694 (N_14694,N_14491,N_14258);
and U14695 (N_14695,N_14456,N_14296);
or U14696 (N_14696,N_14379,N_14332);
or U14697 (N_14697,N_14489,N_14273);
or U14698 (N_14698,N_14351,N_14456);
and U14699 (N_14699,N_14353,N_14363);
and U14700 (N_14700,N_14346,N_14405);
or U14701 (N_14701,N_14253,N_14455);
nor U14702 (N_14702,N_14332,N_14394);
nor U14703 (N_14703,N_14357,N_14301);
and U14704 (N_14704,N_14360,N_14326);
nor U14705 (N_14705,N_14498,N_14477);
and U14706 (N_14706,N_14317,N_14334);
nor U14707 (N_14707,N_14289,N_14447);
nor U14708 (N_14708,N_14321,N_14499);
nor U14709 (N_14709,N_14375,N_14412);
and U14710 (N_14710,N_14328,N_14256);
or U14711 (N_14711,N_14479,N_14407);
and U14712 (N_14712,N_14358,N_14301);
nand U14713 (N_14713,N_14447,N_14339);
nand U14714 (N_14714,N_14484,N_14276);
or U14715 (N_14715,N_14372,N_14478);
or U14716 (N_14716,N_14479,N_14349);
and U14717 (N_14717,N_14406,N_14477);
and U14718 (N_14718,N_14373,N_14451);
nor U14719 (N_14719,N_14394,N_14302);
nand U14720 (N_14720,N_14454,N_14446);
and U14721 (N_14721,N_14379,N_14371);
nor U14722 (N_14722,N_14273,N_14366);
nand U14723 (N_14723,N_14375,N_14275);
and U14724 (N_14724,N_14418,N_14470);
nand U14725 (N_14725,N_14321,N_14317);
and U14726 (N_14726,N_14380,N_14451);
or U14727 (N_14727,N_14437,N_14389);
or U14728 (N_14728,N_14407,N_14482);
or U14729 (N_14729,N_14456,N_14395);
nand U14730 (N_14730,N_14315,N_14386);
or U14731 (N_14731,N_14263,N_14471);
nand U14732 (N_14732,N_14265,N_14394);
nand U14733 (N_14733,N_14291,N_14296);
or U14734 (N_14734,N_14266,N_14319);
and U14735 (N_14735,N_14363,N_14393);
and U14736 (N_14736,N_14292,N_14270);
nand U14737 (N_14737,N_14409,N_14447);
nand U14738 (N_14738,N_14250,N_14463);
or U14739 (N_14739,N_14470,N_14369);
nand U14740 (N_14740,N_14484,N_14299);
and U14741 (N_14741,N_14305,N_14331);
nor U14742 (N_14742,N_14479,N_14255);
or U14743 (N_14743,N_14276,N_14342);
nand U14744 (N_14744,N_14499,N_14352);
and U14745 (N_14745,N_14410,N_14426);
and U14746 (N_14746,N_14346,N_14496);
nor U14747 (N_14747,N_14313,N_14293);
nand U14748 (N_14748,N_14281,N_14453);
xnor U14749 (N_14749,N_14432,N_14398);
nor U14750 (N_14750,N_14662,N_14588);
nand U14751 (N_14751,N_14728,N_14580);
or U14752 (N_14752,N_14640,N_14736);
nor U14753 (N_14753,N_14561,N_14743);
nand U14754 (N_14754,N_14586,N_14725);
nand U14755 (N_14755,N_14641,N_14516);
xor U14756 (N_14756,N_14678,N_14585);
nor U14757 (N_14757,N_14649,N_14650);
and U14758 (N_14758,N_14537,N_14731);
nand U14759 (N_14759,N_14611,N_14621);
nor U14760 (N_14760,N_14705,N_14620);
and U14761 (N_14761,N_14735,N_14553);
and U14762 (N_14762,N_14646,N_14651);
nor U14763 (N_14763,N_14509,N_14505);
nor U14764 (N_14764,N_14571,N_14665);
and U14765 (N_14765,N_14700,N_14689);
or U14766 (N_14766,N_14520,N_14528);
nor U14767 (N_14767,N_14696,N_14666);
or U14768 (N_14768,N_14738,N_14744);
nor U14769 (N_14769,N_14562,N_14721);
or U14770 (N_14770,N_14637,N_14622);
or U14771 (N_14771,N_14625,N_14590);
or U14772 (N_14772,N_14681,N_14507);
nand U14773 (N_14773,N_14519,N_14693);
nor U14774 (N_14774,N_14600,N_14533);
and U14775 (N_14775,N_14708,N_14713);
nor U14776 (N_14776,N_14655,N_14638);
and U14777 (N_14777,N_14690,N_14603);
and U14778 (N_14778,N_14703,N_14527);
and U14779 (N_14779,N_14615,N_14591);
nand U14780 (N_14780,N_14543,N_14523);
nand U14781 (N_14781,N_14673,N_14630);
or U14782 (N_14782,N_14601,N_14563);
or U14783 (N_14783,N_14677,N_14557);
and U14784 (N_14784,N_14566,N_14732);
nand U14785 (N_14785,N_14579,N_14565);
nand U14786 (N_14786,N_14574,N_14572);
nor U14787 (N_14787,N_14577,N_14532);
nand U14788 (N_14788,N_14617,N_14530);
or U14789 (N_14789,N_14501,N_14560);
and U14790 (N_14790,N_14647,N_14682);
or U14791 (N_14791,N_14718,N_14619);
and U14792 (N_14792,N_14540,N_14547);
or U14793 (N_14793,N_14670,N_14564);
or U14794 (N_14794,N_14614,N_14748);
and U14795 (N_14795,N_14653,N_14531);
nand U14796 (N_14796,N_14500,N_14687);
and U14797 (N_14797,N_14645,N_14659);
nor U14798 (N_14798,N_14524,N_14550);
nand U14799 (N_14799,N_14582,N_14522);
or U14800 (N_14800,N_14511,N_14657);
and U14801 (N_14801,N_14644,N_14701);
or U14802 (N_14802,N_14639,N_14602);
nor U14803 (N_14803,N_14660,N_14631);
nand U14804 (N_14804,N_14658,N_14747);
nand U14805 (N_14805,N_14628,N_14538);
nand U14806 (N_14806,N_14612,N_14722);
and U14807 (N_14807,N_14584,N_14711);
and U14808 (N_14808,N_14556,N_14656);
or U14809 (N_14809,N_14545,N_14707);
nand U14810 (N_14810,N_14552,N_14740);
or U14811 (N_14811,N_14594,N_14683);
nor U14812 (N_14812,N_14695,N_14559);
or U14813 (N_14813,N_14742,N_14636);
or U14814 (N_14814,N_14723,N_14605);
nand U14815 (N_14815,N_14684,N_14536);
nor U14816 (N_14816,N_14717,N_14739);
nor U14817 (N_14817,N_14529,N_14569);
nand U14818 (N_14818,N_14633,N_14643);
xor U14819 (N_14819,N_14654,N_14675);
and U14820 (N_14820,N_14679,N_14508);
nor U14821 (N_14821,N_14724,N_14733);
nor U14822 (N_14822,N_14589,N_14672);
nor U14823 (N_14823,N_14555,N_14558);
and U14824 (N_14824,N_14570,N_14661);
or U14825 (N_14825,N_14737,N_14704);
nor U14826 (N_14826,N_14608,N_14518);
nor U14827 (N_14827,N_14746,N_14710);
nand U14828 (N_14828,N_14686,N_14549);
and U14829 (N_14829,N_14749,N_14674);
nor U14830 (N_14830,N_14715,N_14664);
or U14831 (N_14831,N_14583,N_14613);
nand U14832 (N_14832,N_14702,N_14669);
and U14833 (N_14833,N_14521,N_14635);
or U14834 (N_14834,N_14726,N_14729);
nand U14835 (N_14835,N_14627,N_14576);
nand U14836 (N_14836,N_14629,N_14539);
or U14837 (N_14837,N_14512,N_14648);
nand U14838 (N_14838,N_14607,N_14592);
and U14839 (N_14839,N_14598,N_14551);
nor U14840 (N_14840,N_14541,N_14618);
and U14841 (N_14841,N_14623,N_14513);
nor U14842 (N_14842,N_14548,N_14534);
nor U14843 (N_14843,N_14730,N_14642);
nor U14844 (N_14844,N_14734,N_14604);
or U14845 (N_14845,N_14680,N_14581);
or U14846 (N_14846,N_14609,N_14544);
nor U14847 (N_14847,N_14593,N_14510);
or U14848 (N_14848,N_14634,N_14663);
and U14849 (N_14849,N_14504,N_14578);
nor U14850 (N_14850,N_14667,N_14624);
and U14851 (N_14851,N_14567,N_14698);
or U14852 (N_14852,N_14692,N_14716);
nor U14853 (N_14853,N_14503,N_14587);
and U14854 (N_14854,N_14719,N_14616);
and U14855 (N_14855,N_14688,N_14514);
nand U14856 (N_14856,N_14517,N_14626);
nor U14857 (N_14857,N_14546,N_14694);
and U14858 (N_14858,N_14697,N_14535);
nand U14859 (N_14859,N_14573,N_14597);
and U14860 (N_14860,N_14709,N_14526);
nand U14861 (N_14861,N_14610,N_14632);
xor U14862 (N_14862,N_14525,N_14652);
nor U14863 (N_14863,N_14502,N_14599);
nand U14864 (N_14864,N_14676,N_14699);
nor U14865 (N_14865,N_14595,N_14691);
xnor U14866 (N_14866,N_14596,N_14706);
and U14867 (N_14867,N_14712,N_14714);
nor U14868 (N_14868,N_14554,N_14727);
or U14869 (N_14869,N_14685,N_14542);
xnor U14870 (N_14870,N_14606,N_14741);
nor U14871 (N_14871,N_14720,N_14515);
nor U14872 (N_14872,N_14668,N_14506);
and U14873 (N_14873,N_14568,N_14671);
nor U14874 (N_14874,N_14575,N_14745);
nand U14875 (N_14875,N_14735,N_14500);
and U14876 (N_14876,N_14707,N_14711);
and U14877 (N_14877,N_14641,N_14511);
or U14878 (N_14878,N_14719,N_14665);
nor U14879 (N_14879,N_14636,N_14687);
nand U14880 (N_14880,N_14543,N_14584);
nand U14881 (N_14881,N_14618,N_14744);
nor U14882 (N_14882,N_14517,N_14636);
or U14883 (N_14883,N_14517,N_14692);
xnor U14884 (N_14884,N_14558,N_14665);
and U14885 (N_14885,N_14649,N_14691);
and U14886 (N_14886,N_14526,N_14594);
nand U14887 (N_14887,N_14559,N_14507);
nand U14888 (N_14888,N_14548,N_14651);
nor U14889 (N_14889,N_14604,N_14560);
nor U14890 (N_14890,N_14574,N_14744);
nand U14891 (N_14891,N_14724,N_14696);
or U14892 (N_14892,N_14743,N_14622);
and U14893 (N_14893,N_14522,N_14668);
or U14894 (N_14894,N_14608,N_14601);
and U14895 (N_14895,N_14720,N_14524);
nand U14896 (N_14896,N_14502,N_14679);
and U14897 (N_14897,N_14728,N_14628);
or U14898 (N_14898,N_14696,N_14647);
or U14899 (N_14899,N_14738,N_14661);
and U14900 (N_14900,N_14531,N_14515);
nand U14901 (N_14901,N_14647,N_14550);
xor U14902 (N_14902,N_14515,N_14707);
xor U14903 (N_14903,N_14734,N_14699);
and U14904 (N_14904,N_14537,N_14657);
nand U14905 (N_14905,N_14685,N_14575);
nor U14906 (N_14906,N_14522,N_14502);
nor U14907 (N_14907,N_14500,N_14663);
or U14908 (N_14908,N_14625,N_14704);
xnor U14909 (N_14909,N_14614,N_14715);
nand U14910 (N_14910,N_14638,N_14733);
nor U14911 (N_14911,N_14517,N_14572);
and U14912 (N_14912,N_14729,N_14668);
or U14913 (N_14913,N_14683,N_14612);
nand U14914 (N_14914,N_14644,N_14543);
and U14915 (N_14915,N_14574,N_14560);
nor U14916 (N_14916,N_14638,N_14512);
nand U14917 (N_14917,N_14578,N_14562);
nand U14918 (N_14918,N_14503,N_14688);
and U14919 (N_14919,N_14518,N_14670);
nor U14920 (N_14920,N_14646,N_14548);
and U14921 (N_14921,N_14680,N_14614);
nand U14922 (N_14922,N_14521,N_14709);
and U14923 (N_14923,N_14713,N_14685);
nor U14924 (N_14924,N_14560,N_14686);
or U14925 (N_14925,N_14718,N_14633);
or U14926 (N_14926,N_14667,N_14682);
or U14927 (N_14927,N_14715,N_14557);
and U14928 (N_14928,N_14629,N_14721);
and U14929 (N_14929,N_14659,N_14573);
nor U14930 (N_14930,N_14661,N_14656);
nand U14931 (N_14931,N_14695,N_14711);
or U14932 (N_14932,N_14700,N_14693);
nor U14933 (N_14933,N_14558,N_14694);
and U14934 (N_14934,N_14638,N_14550);
nor U14935 (N_14935,N_14599,N_14710);
nor U14936 (N_14936,N_14548,N_14538);
nor U14937 (N_14937,N_14638,N_14615);
or U14938 (N_14938,N_14708,N_14677);
or U14939 (N_14939,N_14709,N_14729);
or U14940 (N_14940,N_14626,N_14513);
and U14941 (N_14941,N_14742,N_14709);
or U14942 (N_14942,N_14584,N_14519);
nand U14943 (N_14943,N_14638,N_14668);
nor U14944 (N_14944,N_14648,N_14588);
nor U14945 (N_14945,N_14697,N_14618);
and U14946 (N_14946,N_14553,N_14741);
nor U14947 (N_14947,N_14643,N_14664);
nand U14948 (N_14948,N_14684,N_14516);
and U14949 (N_14949,N_14688,N_14745);
nand U14950 (N_14950,N_14545,N_14731);
nor U14951 (N_14951,N_14735,N_14572);
or U14952 (N_14952,N_14544,N_14700);
nand U14953 (N_14953,N_14686,N_14744);
nand U14954 (N_14954,N_14528,N_14666);
and U14955 (N_14955,N_14566,N_14545);
nand U14956 (N_14956,N_14675,N_14668);
or U14957 (N_14957,N_14518,N_14725);
and U14958 (N_14958,N_14560,N_14625);
and U14959 (N_14959,N_14687,N_14664);
and U14960 (N_14960,N_14576,N_14748);
nor U14961 (N_14961,N_14583,N_14551);
nand U14962 (N_14962,N_14676,N_14571);
or U14963 (N_14963,N_14720,N_14564);
and U14964 (N_14964,N_14588,N_14522);
and U14965 (N_14965,N_14523,N_14626);
nand U14966 (N_14966,N_14736,N_14625);
and U14967 (N_14967,N_14524,N_14626);
nor U14968 (N_14968,N_14574,N_14737);
nor U14969 (N_14969,N_14666,N_14734);
nor U14970 (N_14970,N_14595,N_14514);
and U14971 (N_14971,N_14589,N_14520);
or U14972 (N_14972,N_14507,N_14702);
nor U14973 (N_14973,N_14670,N_14572);
nand U14974 (N_14974,N_14718,N_14549);
nor U14975 (N_14975,N_14646,N_14715);
or U14976 (N_14976,N_14594,N_14726);
and U14977 (N_14977,N_14731,N_14521);
or U14978 (N_14978,N_14662,N_14697);
or U14979 (N_14979,N_14647,N_14515);
and U14980 (N_14980,N_14732,N_14744);
and U14981 (N_14981,N_14557,N_14638);
and U14982 (N_14982,N_14535,N_14522);
nand U14983 (N_14983,N_14622,N_14725);
nor U14984 (N_14984,N_14553,N_14687);
nor U14985 (N_14985,N_14675,N_14571);
and U14986 (N_14986,N_14735,N_14658);
nand U14987 (N_14987,N_14653,N_14520);
or U14988 (N_14988,N_14597,N_14517);
or U14989 (N_14989,N_14619,N_14578);
or U14990 (N_14990,N_14646,N_14692);
nor U14991 (N_14991,N_14514,N_14695);
or U14992 (N_14992,N_14741,N_14546);
nor U14993 (N_14993,N_14698,N_14738);
nor U14994 (N_14994,N_14666,N_14634);
and U14995 (N_14995,N_14712,N_14624);
and U14996 (N_14996,N_14741,N_14521);
and U14997 (N_14997,N_14726,N_14558);
nand U14998 (N_14998,N_14564,N_14551);
and U14999 (N_14999,N_14557,N_14569);
nor U15000 (N_15000,N_14959,N_14996);
nor U15001 (N_15001,N_14914,N_14890);
nand U15002 (N_15002,N_14971,N_14800);
and U15003 (N_15003,N_14829,N_14979);
nor U15004 (N_15004,N_14757,N_14750);
nand U15005 (N_15005,N_14774,N_14934);
and U15006 (N_15006,N_14963,N_14886);
nand U15007 (N_15007,N_14933,N_14962);
nor U15008 (N_15008,N_14941,N_14834);
and U15009 (N_15009,N_14916,N_14789);
or U15010 (N_15010,N_14773,N_14901);
nand U15011 (N_15011,N_14831,N_14997);
xnor U15012 (N_15012,N_14777,N_14876);
or U15013 (N_15013,N_14906,N_14751);
and U15014 (N_15014,N_14824,N_14781);
or U15015 (N_15015,N_14938,N_14864);
nand U15016 (N_15016,N_14851,N_14999);
and U15017 (N_15017,N_14797,N_14947);
or U15018 (N_15018,N_14993,N_14818);
or U15019 (N_15019,N_14989,N_14983);
nand U15020 (N_15020,N_14986,N_14813);
nor U15021 (N_15021,N_14785,N_14994);
and U15022 (N_15022,N_14949,N_14759);
or U15023 (N_15023,N_14764,N_14907);
nor U15024 (N_15024,N_14809,N_14771);
nand U15025 (N_15025,N_14856,N_14839);
nand U15026 (N_15026,N_14844,N_14988);
nand U15027 (N_15027,N_14958,N_14793);
and U15028 (N_15028,N_14827,N_14841);
or U15029 (N_15029,N_14828,N_14919);
or U15030 (N_15030,N_14806,N_14882);
or U15031 (N_15031,N_14946,N_14917);
or U15032 (N_15032,N_14815,N_14816);
and U15033 (N_15033,N_14861,N_14762);
nand U15034 (N_15034,N_14953,N_14823);
and U15035 (N_15035,N_14926,N_14970);
and U15036 (N_15036,N_14910,N_14951);
nor U15037 (N_15037,N_14950,N_14790);
or U15038 (N_15038,N_14980,N_14837);
xor U15039 (N_15039,N_14911,N_14863);
and U15040 (N_15040,N_14812,N_14865);
and U15041 (N_15041,N_14881,N_14819);
nand U15042 (N_15042,N_14767,N_14794);
nand U15043 (N_15043,N_14768,N_14904);
and U15044 (N_15044,N_14991,N_14898);
nor U15045 (N_15045,N_14817,N_14981);
nand U15046 (N_15046,N_14803,N_14939);
or U15047 (N_15047,N_14845,N_14798);
nor U15048 (N_15048,N_14918,N_14935);
and U15049 (N_15049,N_14955,N_14804);
or U15050 (N_15050,N_14987,N_14968);
nand U15051 (N_15051,N_14811,N_14927);
and U15052 (N_15052,N_14975,N_14753);
nor U15053 (N_15053,N_14969,N_14884);
nor U15054 (N_15054,N_14874,N_14776);
or U15055 (N_15055,N_14807,N_14954);
nor U15056 (N_15056,N_14780,N_14943);
nand U15057 (N_15057,N_14887,N_14899);
xnor U15058 (N_15058,N_14932,N_14859);
nand U15059 (N_15059,N_14972,N_14867);
and U15060 (N_15060,N_14799,N_14847);
or U15061 (N_15061,N_14769,N_14929);
or U15062 (N_15062,N_14838,N_14843);
and U15063 (N_15063,N_14905,N_14973);
nand U15064 (N_15064,N_14995,N_14833);
or U15065 (N_15065,N_14755,N_14871);
or U15066 (N_15066,N_14866,N_14956);
or U15067 (N_15067,N_14897,N_14879);
nand U15068 (N_15068,N_14840,N_14858);
or U15069 (N_15069,N_14852,N_14822);
nand U15070 (N_15070,N_14931,N_14937);
nand U15071 (N_15071,N_14802,N_14779);
or U15072 (N_15072,N_14870,N_14909);
nor U15073 (N_15073,N_14786,N_14920);
nor U15074 (N_15074,N_14810,N_14922);
or U15075 (N_15075,N_14808,N_14795);
nor U15076 (N_15076,N_14900,N_14960);
or U15077 (N_15077,N_14763,N_14862);
or U15078 (N_15078,N_14825,N_14945);
and U15079 (N_15079,N_14814,N_14891);
nand U15080 (N_15080,N_14940,N_14872);
and U15081 (N_15081,N_14896,N_14869);
nand U15082 (N_15082,N_14835,N_14878);
nand U15083 (N_15083,N_14791,N_14842);
or U15084 (N_15084,N_14885,N_14784);
nor U15085 (N_15085,N_14990,N_14912);
nand U15086 (N_15086,N_14801,N_14977);
or U15087 (N_15087,N_14942,N_14855);
nand U15088 (N_15088,N_14752,N_14849);
nand U15089 (N_15089,N_14846,N_14913);
nand U15090 (N_15090,N_14782,N_14923);
nor U15091 (N_15091,N_14895,N_14765);
and U15092 (N_15092,N_14894,N_14772);
and U15093 (N_15093,N_14985,N_14915);
and U15094 (N_15094,N_14761,N_14830);
nor U15095 (N_15095,N_14787,N_14944);
nor U15096 (N_15096,N_14775,N_14967);
and U15097 (N_15097,N_14948,N_14778);
nand U15098 (N_15098,N_14902,N_14875);
nand U15099 (N_15099,N_14873,N_14850);
nand U15100 (N_15100,N_14889,N_14982);
and U15101 (N_15101,N_14820,N_14853);
and U15102 (N_15102,N_14832,N_14966);
nor U15103 (N_15103,N_14925,N_14908);
nor U15104 (N_15104,N_14783,N_14756);
nor U15105 (N_15105,N_14998,N_14854);
or U15106 (N_15106,N_14760,N_14826);
or U15107 (N_15107,N_14883,N_14992);
nand U15108 (N_15108,N_14952,N_14796);
and U15109 (N_15109,N_14857,N_14821);
nor U15110 (N_15110,N_14921,N_14766);
nor U15111 (N_15111,N_14930,N_14877);
nand U15112 (N_15112,N_14957,N_14893);
nor U15113 (N_15113,N_14924,N_14792);
and U15114 (N_15114,N_14848,N_14936);
and U15115 (N_15115,N_14974,N_14860);
or U15116 (N_15116,N_14961,N_14880);
or U15117 (N_15117,N_14888,N_14984);
nand U15118 (N_15118,N_14836,N_14788);
and U15119 (N_15119,N_14978,N_14976);
nor U15120 (N_15120,N_14892,N_14928);
and U15121 (N_15121,N_14754,N_14903);
and U15122 (N_15122,N_14758,N_14964);
or U15123 (N_15123,N_14965,N_14868);
nor U15124 (N_15124,N_14805,N_14770);
or U15125 (N_15125,N_14818,N_14962);
nand U15126 (N_15126,N_14876,N_14970);
and U15127 (N_15127,N_14760,N_14979);
nor U15128 (N_15128,N_14765,N_14853);
or U15129 (N_15129,N_14852,N_14775);
or U15130 (N_15130,N_14991,N_14784);
nor U15131 (N_15131,N_14820,N_14979);
nor U15132 (N_15132,N_14875,N_14960);
nor U15133 (N_15133,N_14800,N_14903);
and U15134 (N_15134,N_14817,N_14802);
or U15135 (N_15135,N_14982,N_14772);
and U15136 (N_15136,N_14867,N_14994);
and U15137 (N_15137,N_14827,N_14850);
or U15138 (N_15138,N_14814,N_14871);
or U15139 (N_15139,N_14895,N_14914);
and U15140 (N_15140,N_14862,N_14869);
or U15141 (N_15141,N_14903,N_14815);
nor U15142 (N_15142,N_14796,N_14787);
nor U15143 (N_15143,N_14796,N_14776);
nor U15144 (N_15144,N_14888,N_14858);
nor U15145 (N_15145,N_14759,N_14849);
nor U15146 (N_15146,N_14986,N_14934);
nand U15147 (N_15147,N_14930,N_14993);
nand U15148 (N_15148,N_14824,N_14750);
or U15149 (N_15149,N_14901,N_14984);
nor U15150 (N_15150,N_14997,N_14870);
nor U15151 (N_15151,N_14986,N_14900);
nor U15152 (N_15152,N_14883,N_14840);
and U15153 (N_15153,N_14752,N_14836);
or U15154 (N_15154,N_14916,N_14836);
nor U15155 (N_15155,N_14823,N_14835);
nor U15156 (N_15156,N_14774,N_14887);
nor U15157 (N_15157,N_14873,N_14761);
or U15158 (N_15158,N_14852,N_14910);
nand U15159 (N_15159,N_14795,N_14959);
nor U15160 (N_15160,N_14953,N_14970);
nor U15161 (N_15161,N_14788,N_14829);
or U15162 (N_15162,N_14972,N_14991);
nand U15163 (N_15163,N_14923,N_14798);
or U15164 (N_15164,N_14886,N_14879);
and U15165 (N_15165,N_14990,N_14928);
nor U15166 (N_15166,N_14851,N_14903);
nand U15167 (N_15167,N_14876,N_14857);
and U15168 (N_15168,N_14766,N_14956);
or U15169 (N_15169,N_14908,N_14794);
nor U15170 (N_15170,N_14850,N_14846);
and U15171 (N_15171,N_14958,N_14858);
and U15172 (N_15172,N_14801,N_14942);
and U15173 (N_15173,N_14871,N_14807);
and U15174 (N_15174,N_14999,N_14888);
and U15175 (N_15175,N_14998,N_14755);
and U15176 (N_15176,N_14871,N_14942);
and U15177 (N_15177,N_14750,N_14859);
and U15178 (N_15178,N_14932,N_14757);
or U15179 (N_15179,N_14981,N_14791);
nand U15180 (N_15180,N_14941,N_14881);
nand U15181 (N_15181,N_14821,N_14817);
and U15182 (N_15182,N_14854,N_14994);
nor U15183 (N_15183,N_14845,N_14769);
nand U15184 (N_15184,N_14932,N_14782);
nor U15185 (N_15185,N_14794,N_14953);
and U15186 (N_15186,N_14836,N_14994);
nand U15187 (N_15187,N_14930,N_14846);
or U15188 (N_15188,N_14858,N_14767);
nor U15189 (N_15189,N_14934,N_14782);
or U15190 (N_15190,N_14998,N_14781);
and U15191 (N_15191,N_14817,N_14904);
and U15192 (N_15192,N_14983,N_14946);
or U15193 (N_15193,N_14875,N_14903);
nor U15194 (N_15194,N_14993,N_14821);
nor U15195 (N_15195,N_14930,N_14823);
or U15196 (N_15196,N_14795,N_14942);
nand U15197 (N_15197,N_14770,N_14750);
nor U15198 (N_15198,N_14944,N_14925);
nor U15199 (N_15199,N_14764,N_14983);
or U15200 (N_15200,N_14966,N_14940);
nand U15201 (N_15201,N_14935,N_14963);
nand U15202 (N_15202,N_14969,N_14752);
nor U15203 (N_15203,N_14801,N_14789);
nor U15204 (N_15204,N_14869,N_14904);
nand U15205 (N_15205,N_14858,N_14999);
nand U15206 (N_15206,N_14751,N_14919);
nor U15207 (N_15207,N_14955,N_14900);
or U15208 (N_15208,N_14783,N_14934);
or U15209 (N_15209,N_14835,N_14896);
or U15210 (N_15210,N_14792,N_14982);
nor U15211 (N_15211,N_14806,N_14942);
and U15212 (N_15212,N_14848,N_14842);
and U15213 (N_15213,N_14797,N_14896);
and U15214 (N_15214,N_14921,N_14895);
and U15215 (N_15215,N_14772,N_14769);
or U15216 (N_15216,N_14973,N_14982);
nor U15217 (N_15217,N_14834,N_14958);
and U15218 (N_15218,N_14965,N_14776);
nor U15219 (N_15219,N_14876,N_14923);
nor U15220 (N_15220,N_14837,N_14756);
xnor U15221 (N_15221,N_14880,N_14888);
nor U15222 (N_15222,N_14766,N_14852);
or U15223 (N_15223,N_14776,N_14958);
nor U15224 (N_15224,N_14758,N_14904);
nor U15225 (N_15225,N_14832,N_14909);
and U15226 (N_15226,N_14993,N_14777);
or U15227 (N_15227,N_14752,N_14920);
nor U15228 (N_15228,N_14874,N_14965);
nand U15229 (N_15229,N_14848,N_14952);
nand U15230 (N_15230,N_14849,N_14787);
and U15231 (N_15231,N_14924,N_14908);
nor U15232 (N_15232,N_14925,N_14840);
nand U15233 (N_15233,N_14764,N_14759);
nor U15234 (N_15234,N_14751,N_14868);
and U15235 (N_15235,N_14789,N_14962);
nand U15236 (N_15236,N_14789,N_14815);
nand U15237 (N_15237,N_14921,N_14960);
or U15238 (N_15238,N_14879,N_14775);
nand U15239 (N_15239,N_14809,N_14859);
nor U15240 (N_15240,N_14968,N_14846);
nor U15241 (N_15241,N_14757,N_14936);
and U15242 (N_15242,N_14981,N_14849);
or U15243 (N_15243,N_14990,N_14919);
nor U15244 (N_15244,N_14960,N_14772);
nand U15245 (N_15245,N_14816,N_14925);
or U15246 (N_15246,N_14872,N_14885);
nand U15247 (N_15247,N_14810,N_14797);
nor U15248 (N_15248,N_14870,N_14754);
or U15249 (N_15249,N_14962,N_14804);
nand U15250 (N_15250,N_15232,N_15098);
and U15251 (N_15251,N_15087,N_15074);
or U15252 (N_15252,N_15249,N_15099);
nand U15253 (N_15253,N_15169,N_15130);
or U15254 (N_15254,N_15094,N_15159);
nor U15255 (N_15255,N_15201,N_15015);
nor U15256 (N_15256,N_15102,N_15118);
and U15257 (N_15257,N_15004,N_15078);
nor U15258 (N_15258,N_15104,N_15097);
nor U15259 (N_15259,N_15075,N_15008);
nand U15260 (N_15260,N_15124,N_15196);
and U15261 (N_15261,N_15095,N_15014);
nor U15262 (N_15262,N_15171,N_15138);
and U15263 (N_15263,N_15212,N_15068);
and U15264 (N_15264,N_15059,N_15139);
and U15265 (N_15265,N_15009,N_15243);
nor U15266 (N_15266,N_15076,N_15117);
nor U15267 (N_15267,N_15029,N_15000);
and U15268 (N_15268,N_15142,N_15048);
xnor U15269 (N_15269,N_15018,N_15120);
nand U15270 (N_15270,N_15032,N_15235);
and U15271 (N_15271,N_15016,N_15054);
nand U15272 (N_15272,N_15181,N_15127);
and U15273 (N_15273,N_15046,N_15161);
and U15274 (N_15274,N_15101,N_15012);
or U15275 (N_15275,N_15246,N_15100);
or U15276 (N_15276,N_15093,N_15019);
and U15277 (N_15277,N_15050,N_15038);
nand U15278 (N_15278,N_15224,N_15121);
and U15279 (N_15279,N_15233,N_15092);
nand U15280 (N_15280,N_15239,N_15109);
and U15281 (N_15281,N_15144,N_15136);
and U15282 (N_15282,N_15119,N_15112);
nor U15283 (N_15283,N_15024,N_15215);
or U15284 (N_15284,N_15220,N_15174);
or U15285 (N_15285,N_15203,N_15190);
and U15286 (N_15286,N_15085,N_15107);
and U15287 (N_15287,N_15185,N_15194);
nor U15288 (N_15288,N_15184,N_15156);
or U15289 (N_15289,N_15066,N_15027);
and U15290 (N_15290,N_15129,N_15137);
and U15291 (N_15291,N_15089,N_15219);
nand U15292 (N_15292,N_15060,N_15134);
nor U15293 (N_15293,N_15053,N_15162);
nor U15294 (N_15294,N_15153,N_15044);
or U15295 (N_15295,N_15062,N_15141);
nand U15296 (N_15296,N_15163,N_15225);
nand U15297 (N_15297,N_15216,N_15182);
nand U15298 (N_15298,N_15001,N_15248);
or U15299 (N_15299,N_15151,N_15072);
nand U15300 (N_15300,N_15126,N_15023);
nand U15301 (N_15301,N_15133,N_15170);
or U15302 (N_15302,N_15007,N_15135);
nand U15303 (N_15303,N_15025,N_15140);
nand U15304 (N_15304,N_15228,N_15242);
and U15305 (N_15305,N_15017,N_15166);
and U15306 (N_15306,N_15180,N_15222);
or U15307 (N_15307,N_15035,N_15067);
and U15308 (N_15308,N_15218,N_15186);
and U15309 (N_15309,N_15205,N_15211);
nor U15310 (N_15310,N_15083,N_15217);
and U15311 (N_15311,N_15021,N_15005);
or U15312 (N_15312,N_15192,N_15195);
nor U15313 (N_15313,N_15096,N_15150);
nor U15314 (N_15314,N_15110,N_15040);
or U15315 (N_15315,N_15208,N_15036);
nor U15316 (N_15316,N_15070,N_15176);
nand U15317 (N_15317,N_15223,N_15193);
or U15318 (N_15318,N_15073,N_15206);
and U15319 (N_15319,N_15152,N_15145);
nand U15320 (N_15320,N_15081,N_15241);
nand U15321 (N_15321,N_15006,N_15034);
or U15322 (N_15322,N_15230,N_15202);
and U15323 (N_15323,N_15113,N_15231);
nor U15324 (N_15324,N_15188,N_15227);
nor U15325 (N_15325,N_15221,N_15013);
or U15326 (N_15326,N_15091,N_15172);
or U15327 (N_15327,N_15031,N_15160);
and U15328 (N_15328,N_15103,N_15238);
nand U15329 (N_15329,N_15234,N_15049);
or U15330 (N_15330,N_15041,N_15183);
or U15331 (N_15331,N_15158,N_15236);
and U15332 (N_15332,N_15200,N_15042);
nor U15333 (N_15333,N_15058,N_15123);
and U15334 (N_15334,N_15199,N_15088);
or U15335 (N_15335,N_15164,N_15011);
nor U15336 (N_15336,N_15077,N_15177);
and U15337 (N_15337,N_15131,N_15079);
and U15338 (N_15338,N_15064,N_15115);
nor U15339 (N_15339,N_15132,N_15002);
and U15340 (N_15340,N_15111,N_15213);
nor U15341 (N_15341,N_15240,N_15244);
nand U15342 (N_15342,N_15214,N_15116);
and U15343 (N_15343,N_15179,N_15149);
or U15344 (N_15344,N_15010,N_15122);
or U15345 (N_15345,N_15055,N_15178);
nor U15346 (N_15346,N_15028,N_15045);
and U15347 (N_15347,N_15090,N_15069);
nor U15348 (N_15348,N_15051,N_15056);
nor U15349 (N_15349,N_15039,N_15229);
nor U15350 (N_15350,N_15147,N_15168);
and U15351 (N_15351,N_15080,N_15128);
and U15352 (N_15352,N_15189,N_15237);
nand U15353 (N_15353,N_15226,N_15084);
and U15354 (N_15354,N_15197,N_15148);
and U15355 (N_15355,N_15052,N_15175);
nor U15356 (N_15356,N_15154,N_15198);
nand U15357 (N_15357,N_15026,N_15071);
nor U15358 (N_15358,N_15207,N_15105);
or U15359 (N_15359,N_15204,N_15143);
and U15360 (N_15360,N_15245,N_15157);
nand U15361 (N_15361,N_15209,N_15106);
and U15362 (N_15362,N_15003,N_15173);
nor U15363 (N_15363,N_15030,N_15247);
or U15364 (N_15364,N_15061,N_15086);
nand U15365 (N_15365,N_15082,N_15125);
nand U15366 (N_15366,N_15191,N_15165);
nor U15367 (N_15367,N_15146,N_15057);
nand U15368 (N_15368,N_15108,N_15047);
nand U15369 (N_15369,N_15020,N_15114);
nand U15370 (N_15370,N_15043,N_15167);
and U15371 (N_15371,N_15033,N_15155);
nor U15372 (N_15372,N_15065,N_15187);
or U15373 (N_15373,N_15210,N_15022);
nand U15374 (N_15374,N_15063,N_15037);
nor U15375 (N_15375,N_15213,N_15019);
and U15376 (N_15376,N_15226,N_15140);
nor U15377 (N_15377,N_15247,N_15241);
nor U15378 (N_15378,N_15188,N_15197);
and U15379 (N_15379,N_15136,N_15200);
nor U15380 (N_15380,N_15212,N_15040);
nor U15381 (N_15381,N_15089,N_15232);
or U15382 (N_15382,N_15028,N_15203);
or U15383 (N_15383,N_15143,N_15066);
nor U15384 (N_15384,N_15029,N_15211);
nor U15385 (N_15385,N_15059,N_15144);
nand U15386 (N_15386,N_15188,N_15038);
nor U15387 (N_15387,N_15122,N_15058);
nor U15388 (N_15388,N_15007,N_15097);
xor U15389 (N_15389,N_15194,N_15133);
nor U15390 (N_15390,N_15246,N_15136);
nand U15391 (N_15391,N_15013,N_15156);
nand U15392 (N_15392,N_15004,N_15248);
nor U15393 (N_15393,N_15095,N_15078);
or U15394 (N_15394,N_15082,N_15032);
nand U15395 (N_15395,N_15225,N_15024);
nor U15396 (N_15396,N_15154,N_15219);
nand U15397 (N_15397,N_15022,N_15164);
nor U15398 (N_15398,N_15052,N_15111);
and U15399 (N_15399,N_15123,N_15014);
nor U15400 (N_15400,N_15152,N_15161);
nor U15401 (N_15401,N_15216,N_15040);
nand U15402 (N_15402,N_15153,N_15045);
and U15403 (N_15403,N_15152,N_15096);
and U15404 (N_15404,N_15137,N_15061);
xnor U15405 (N_15405,N_15206,N_15225);
nand U15406 (N_15406,N_15192,N_15157);
or U15407 (N_15407,N_15059,N_15056);
and U15408 (N_15408,N_15034,N_15095);
and U15409 (N_15409,N_15043,N_15228);
nand U15410 (N_15410,N_15083,N_15121);
and U15411 (N_15411,N_15090,N_15056);
nor U15412 (N_15412,N_15040,N_15197);
nor U15413 (N_15413,N_15237,N_15074);
nor U15414 (N_15414,N_15120,N_15203);
or U15415 (N_15415,N_15133,N_15106);
nand U15416 (N_15416,N_15115,N_15214);
or U15417 (N_15417,N_15200,N_15086);
and U15418 (N_15418,N_15148,N_15055);
or U15419 (N_15419,N_15071,N_15177);
or U15420 (N_15420,N_15039,N_15018);
nand U15421 (N_15421,N_15190,N_15094);
nand U15422 (N_15422,N_15145,N_15157);
nand U15423 (N_15423,N_15047,N_15016);
and U15424 (N_15424,N_15169,N_15133);
or U15425 (N_15425,N_15024,N_15197);
nand U15426 (N_15426,N_15138,N_15053);
nand U15427 (N_15427,N_15189,N_15210);
nand U15428 (N_15428,N_15016,N_15029);
or U15429 (N_15429,N_15021,N_15226);
or U15430 (N_15430,N_15131,N_15244);
or U15431 (N_15431,N_15193,N_15206);
nor U15432 (N_15432,N_15138,N_15134);
and U15433 (N_15433,N_15235,N_15123);
nand U15434 (N_15434,N_15076,N_15140);
nand U15435 (N_15435,N_15236,N_15013);
nand U15436 (N_15436,N_15043,N_15096);
nor U15437 (N_15437,N_15238,N_15017);
nand U15438 (N_15438,N_15229,N_15153);
or U15439 (N_15439,N_15055,N_15102);
or U15440 (N_15440,N_15218,N_15107);
nor U15441 (N_15441,N_15186,N_15190);
nand U15442 (N_15442,N_15107,N_15040);
nor U15443 (N_15443,N_15079,N_15116);
nand U15444 (N_15444,N_15233,N_15073);
and U15445 (N_15445,N_15173,N_15071);
nor U15446 (N_15446,N_15099,N_15244);
and U15447 (N_15447,N_15019,N_15237);
and U15448 (N_15448,N_15184,N_15226);
nand U15449 (N_15449,N_15225,N_15066);
or U15450 (N_15450,N_15177,N_15195);
or U15451 (N_15451,N_15117,N_15186);
and U15452 (N_15452,N_15014,N_15212);
and U15453 (N_15453,N_15210,N_15114);
or U15454 (N_15454,N_15045,N_15186);
nor U15455 (N_15455,N_15222,N_15061);
nor U15456 (N_15456,N_15060,N_15074);
nor U15457 (N_15457,N_15145,N_15099);
or U15458 (N_15458,N_15167,N_15053);
nor U15459 (N_15459,N_15117,N_15212);
or U15460 (N_15460,N_15069,N_15068);
xnor U15461 (N_15461,N_15056,N_15085);
nor U15462 (N_15462,N_15130,N_15097);
and U15463 (N_15463,N_15215,N_15202);
nor U15464 (N_15464,N_15053,N_15214);
or U15465 (N_15465,N_15133,N_15069);
nor U15466 (N_15466,N_15099,N_15204);
or U15467 (N_15467,N_15093,N_15040);
or U15468 (N_15468,N_15002,N_15130);
and U15469 (N_15469,N_15160,N_15145);
or U15470 (N_15470,N_15069,N_15239);
or U15471 (N_15471,N_15143,N_15130);
or U15472 (N_15472,N_15224,N_15102);
nand U15473 (N_15473,N_15001,N_15242);
nand U15474 (N_15474,N_15087,N_15130);
nand U15475 (N_15475,N_15055,N_15002);
nand U15476 (N_15476,N_15209,N_15006);
nand U15477 (N_15477,N_15022,N_15046);
or U15478 (N_15478,N_15090,N_15087);
nand U15479 (N_15479,N_15184,N_15056);
nand U15480 (N_15480,N_15096,N_15186);
nor U15481 (N_15481,N_15097,N_15032);
nor U15482 (N_15482,N_15050,N_15047);
nor U15483 (N_15483,N_15088,N_15195);
xor U15484 (N_15484,N_15015,N_15092);
and U15485 (N_15485,N_15114,N_15179);
or U15486 (N_15486,N_15064,N_15081);
nor U15487 (N_15487,N_15137,N_15026);
nor U15488 (N_15488,N_15177,N_15203);
and U15489 (N_15489,N_15046,N_15060);
and U15490 (N_15490,N_15225,N_15001);
nand U15491 (N_15491,N_15072,N_15103);
nor U15492 (N_15492,N_15069,N_15171);
or U15493 (N_15493,N_15196,N_15158);
nand U15494 (N_15494,N_15205,N_15235);
and U15495 (N_15495,N_15189,N_15033);
nand U15496 (N_15496,N_15141,N_15065);
nand U15497 (N_15497,N_15063,N_15065);
nor U15498 (N_15498,N_15044,N_15203);
or U15499 (N_15499,N_15122,N_15203);
and U15500 (N_15500,N_15472,N_15401);
nand U15501 (N_15501,N_15400,N_15427);
nor U15502 (N_15502,N_15359,N_15302);
and U15503 (N_15503,N_15489,N_15366);
or U15504 (N_15504,N_15375,N_15266);
nor U15505 (N_15505,N_15442,N_15311);
and U15506 (N_15506,N_15468,N_15297);
nand U15507 (N_15507,N_15345,N_15484);
and U15508 (N_15508,N_15316,N_15323);
and U15509 (N_15509,N_15336,N_15291);
nor U15510 (N_15510,N_15327,N_15313);
nor U15511 (N_15511,N_15305,N_15340);
nand U15512 (N_15512,N_15329,N_15378);
or U15513 (N_15513,N_15478,N_15462);
xnor U15514 (N_15514,N_15449,N_15274);
nor U15515 (N_15515,N_15318,N_15490);
and U15516 (N_15516,N_15360,N_15333);
nor U15517 (N_15517,N_15446,N_15381);
or U15518 (N_15518,N_15420,N_15289);
nor U15519 (N_15519,N_15288,N_15404);
nand U15520 (N_15520,N_15447,N_15418);
or U15521 (N_15521,N_15352,N_15441);
nand U15522 (N_15522,N_15388,N_15259);
and U15523 (N_15523,N_15453,N_15379);
and U15524 (N_15524,N_15406,N_15324);
nor U15525 (N_15525,N_15393,N_15399);
nand U15526 (N_15526,N_15486,N_15416);
and U15527 (N_15527,N_15306,N_15424);
and U15528 (N_15528,N_15402,N_15439);
nand U15529 (N_15529,N_15264,N_15372);
nand U15530 (N_15530,N_15321,N_15389);
and U15531 (N_15531,N_15475,N_15312);
and U15532 (N_15532,N_15304,N_15296);
and U15533 (N_15533,N_15431,N_15354);
or U15534 (N_15534,N_15386,N_15250);
nand U15535 (N_15535,N_15347,N_15328);
and U15536 (N_15536,N_15254,N_15283);
nand U15537 (N_15537,N_15367,N_15303);
and U15538 (N_15538,N_15383,N_15314);
nand U15539 (N_15539,N_15493,N_15298);
and U15540 (N_15540,N_15255,N_15355);
and U15541 (N_15541,N_15317,N_15451);
or U15542 (N_15542,N_15405,N_15445);
nand U15543 (N_15543,N_15448,N_15271);
nand U15544 (N_15544,N_15309,N_15498);
nor U15545 (N_15545,N_15377,N_15396);
nor U15546 (N_15546,N_15275,N_15260);
nor U15547 (N_15547,N_15488,N_15350);
nand U15548 (N_15548,N_15301,N_15487);
nand U15549 (N_15549,N_15335,N_15422);
nor U15550 (N_15550,N_15410,N_15343);
and U15551 (N_15551,N_15494,N_15346);
or U15552 (N_15552,N_15425,N_15411);
or U15553 (N_15553,N_15262,N_15270);
and U15554 (N_15554,N_15390,N_15339);
xor U15555 (N_15555,N_15459,N_15483);
and U15556 (N_15556,N_15436,N_15479);
nand U15557 (N_15557,N_15429,N_15307);
or U15558 (N_15558,N_15257,N_15435);
or U15559 (N_15559,N_15369,N_15368);
nand U15560 (N_15560,N_15403,N_15286);
nand U15561 (N_15561,N_15437,N_15408);
nor U15562 (N_15562,N_15457,N_15480);
and U15563 (N_15563,N_15438,N_15481);
nand U15564 (N_15564,N_15330,N_15466);
nand U15565 (N_15565,N_15473,N_15251);
nand U15566 (N_15566,N_15474,N_15491);
and U15567 (N_15567,N_15285,N_15461);
or U15568 (N_15568,N_15421,N_15348);
nand U15569 (N_15569,N_15256,N_15332);
and U15570 (N_15570,N_15353,N_15281);
nor U15571 (N_15571,N_15471,N_15452);
and U15572 (N_15572,N_15279,N_15428);
nand U15573 (N_15573,N_15342,N_15278);
nor U15574 (N_15574,N_15430,N_15252);
nand U15575 (N_15575,N_15398,N_15423);
or U15576 (N_15576,N_15391,N_15385);
nand U15577 (N_15577,N_15337,N_15365);
and U15578 (N_15578,N_15485,N_15432);
nand U15579 (N_15579,N_15287,N_15392);
nor U15580 (N_15580,N_15443,N_15356);
and U15581 (N_15581,N_15415,N_15394);
nand U15582 (N_15582,N_15300,N_15362);
and U15583 (N_15583,N_15496,N_15361);
or U15584 (N_15584,N_15450,N_15290);
nor U15585 (N_15585,N_15349,N_15334);
nor U15586 (N_15586,N_15276,N_15499);
and U15587 (N_15587,N_15456,N_15284);
nand U15588 (N_15588,N_15477,N_15414);
and U15589 (N_15589,N_15320,N_15364);
nor U15590 (N_15590,N_15294,N_15497);
and U15591 (N_15591,N_15444,N_15269);
and U15592 (N_15592,N_15413,N_15326);
nand U15593 (N_15593,N_15338,N_15370);
nor U15594 (N_15594,N_15322,N_15409);
or U15595 (N_15595,N_15407,N_15351);
or U15596 (N_15596,N_15267,N_15458);
or U15597 (N_15597,N_15253,N_15341);
nand U15598 (N_15598,N_15412,N_15299);
or U15599 (N_15599,N_15272,N_15469);
or U15600 (N_15600,N_15268,N_15292);
nor U15601 (N_15601,N_15482,N_15273);
nand U15602 (N_15602,N_15467,N_15454);
or U15603 (N_15603,N_15476,N_15325);
nor U15604 (N_15604,N_15387,N_15295);
nand U15605 (N_15605,N_15258,N_15265);
and U15606 (N_15606,N_15380,N_15344);
and U15607 (N_15607,N_15470,N_15280);
and U15608 (N_15608,N_15426,N_15277);
or U15609 (N_15609,N_15373,N_15417);
nor U15610 (N_15610,N_15495,N_15263);
and U15611 (N_15611,N_15382,N_15374);
nor U15612 (N_15612,N_15363,N_15308);
nor U15613 (N_15613,N_15358,N_15465);
or U15614 (N_15614,N_15319,N_15440);
nand U15615 (N_15615,N_15384,N_15460);
and U15616 (N_15616,N_15397,N_15395);
or U15617 (N_15617,N_15464,N_15357);
nand U15618 (N_15618,N_15376,N_15282);
nand U15619 (N_15619,N_15315,N_15419);
nor U15620 (N_15620,N_15463,N_15331);
nand U15621 (N_15621,N_15492,N_15261);
nand U15622 (N_15622,N_15434,N_15310);
and U15623 (N_15623,N_15433,N_15293);
or U15624 (N_15624,N_15455,N_15371);
and U15625 (N_15625,N_15379,N_15419);
and U15626 (N_15626,N_15336,N_15363);
nand U15627 (N_15627,N_15283,N_15494);
nor U15628 (N_15628,N_15469,N_15490);
nand U15629 (N_15629,N_15291,N_15421);
nor U15630 (N_15630,N_15354,N_15425);
nor U15631 (N_15631,N_15288,N_15381);
nor U15632 (N_15632,N_15476,N_15323);
or U15633 (N_15633,N_15293,N_15408);
and U15634 (N_15634,N_15434,N_15395);
nand U15635 (N_15635,N_15433,N_15426);
and U15636 (N_15636,N_15394,N_15398);
nor U15637 (N_15637,N_15421,N_15436);
and U15638 (N_15638,N_15375,N_15466);
nor U15639 (N_15639,N_15345,N_15378);
or U15640 (N_15640,N_15419,N_15278);
and U15641 (N_15641,N_15349,N_15319);
and U15642 (N_15642,N_15259,N_15375);
and U15643 (N_15643,N_15372,N_15341);
or U15644 (N_15644,N_15391,N_15266);
or U15645 (N_15645,N_15367,N_15341);
or U15646 (N_15646,N_15284,N_15323);
nand U15647 (N_15647,N_15268,N_15262);
nand U15648 (N_15648,N_15356,N_15347);
nor U15649 (N_15649,N_15409,N_15492);
nor U15650 (N_15650,N_15472,N_15469);
or U15651 (N_15651,N_15443,N_15361);
or U15652 (N_15652,N_15332,N_15499);
and U15653 (N_15653,N_15273,N_15484);
nor U15654 (N_15654,N_15255,N_15433);
and U15655 (N_15655,N_15441,N_15296);
or U15656 (N_15656,N_15445,N_15409);
and U15657 (N_15657,N_15319,N_15326);
nor U15658 (N_15658,N_15373,N_15295);
nand U15659 (N_15659,N_15436,N_15341);
nor U15660 (N_15660,N_15486,N_15268);
and U15661 (N_15661,N_15251,N_15408);
or U15662 (N_15662,N_15303,N_15488);
and U15663 (N_15663,N_15291,N_15364);
nor U15664 (N_15664,N_15346,N_15307);
nand U15665 (N_15665,N_15256,N_15364);
nand U15666 (N_15666,N_15332,N_15485);
and U15667 (N_15667,N_15310,N_15301);
nor U15668 (N_15668,N_15458,N_15337);
nand U15669 (N_15669,N_15490,N_15409);
or U15670 (N_15670,N_15328,N_15412);
and U15671 (N_15671,N_15277,N_15366);
and U15672 (N_15672,N_15316,N_15309);
nor U15673 (N_15673,N_15316,N_15413);
nor U15674 (N_15674,N_15376,N_15491);
and U15675 (N_15675,N_15395,N_15333);
or U15676 (N_15676,N_15417,N_15443);
and U15677 (N_15677,N_15460,N_15451);
nand U15678 (N_15678,N_15431,N_15320);
and U15679 (N_15679,N_15278,N_15270);
nand U15680 (N_15680,N_15329,N_15270);
nand U15681 (N_15681,N_15361,N_15403);
nor U15682 (N_15682,N_15486,N_15335);
or U15683 (N_15683,N_15370,N_15481);
and U15684 (N_15684,N_15428,N_15444);
nand U15685 (N_15685,N_15471,N_15433);
and U15686 (N_15686,N_15342,N_15250);
or U15687 (N_15687,N_15269,N_15380);
nand U15688 (N_15688,N_15313,N_15334);
and U15689 (N_15689,N_15338,N_15323);
and U15690 (N_15690,N_15467,N_15257);
and U15691 (N_15691,N_15309,N_15360);
or U15692 (N_15692,N_15289,N_15470);
nand U15693 (N_15693,N_15386,N_15251);
nor U15694 (N_15694,N_15343,N_15328);
or U15695 (N_15695,N_15417,N_15418);
or U15696 (N_15696,N_15335,N_15375);
or U15697 (N_15697,N_15431,N_15429);
nand U15698 (N_15698,N_15435,N_15488);
and U15699 (N_15699,N_15299,N_15250);
and U15700 (N_15700,N_15396,N_15491);
nor U15701 (N_15701,N_15359,N_15477);
and U15702 (N_15702,N_15268,N_15273);
nor U15703 (N_15703,N_15354,N_15406);
nor U15704 (N_15704,N_15444,N_15291);
nand U15705 (N_15705,N_15254,N_15380);
or U15706 (N_15706,N_15481,N_15285);
nand U15707 (N_15707,N_15487,N_15356);
or U15708 (N_15708,N_15312,N_15282);
or U15709 (N_15709,N_15359,N_15409);
or U15710 (N_15710,N_15324,N_15263);
and U15711 (N_15711,N_15495,N_15360);
or U15712 (N_15712,N_15418,N_15283);
or U15713 (N_15713,N_15324,N_15332);
and U15714 (N_15714,N_15276,N_15263);
nor U15715 (N_15715,N_15360,N_15411);
and U15716 (N_15716,N_15299,N_15417);
nor U15717 (N_15717,N_15351,N_15299);
or U15718 (N_15718,N_15406,N_15337);
nor U15719 (N_15719,N_15421,N_15374);
nor U15720 (N_15720,N_15284,N_15259);
or U15721 (N_15721,N_15492,N_15380);
xnor U15722 (N_15722,N_15337,N_15387);
or U15723 (N_15723,N_15413,N_15401);
and U15724 (N_15724,N_15340,N_15457);
nor U15725 (N_15725,N_15460,N_15461);
nand U15726 (N_15726,N_15335,N_15460);
nand U15727 (N_15727,N_15466,N_15448);
or U15728 (N_15728,N_15406,N_15461);
and U15729 (N_15729,N_15293,N_15262);
nor U15730 (N_15730,N_15271,N_15279);
or U15731 (N_15731,N_15452,N_15272);
or U15732 (N_15732,N_15325,N_15444);
nor U15733 (N_15733,N_15251,N_15448);
or U15734 (N_15734,N_15321,N_15292);
nor U15735 (N_15735,N_15290,N_15387);
or U15736 (N_15736,N_15445,N_15487);
nand U15737 (N_15737,N_15392,N_15250);
or U15738 (N_15738,N_15322,N_15300);
nor U15739 (N_15739,N_15306,N_15375);
nand U15740 (N_15740,N_15282,N_15423);
and U15741 (N_15741,N_15253,N_15452);
nand U15742 (N_15742,N_15387,N_15340);
nand U15743 (N_15743,N_15388,N_15350);
nor U15744 (N_15744,N_15374,N_15256);
nand U15745 (N_15745,N_15337,N_15250);
xnor U15746 (N_15746,N_15318,N_15393);
nor U15747 (N_15747,N_15262,N_15429);
and U15748 (N_15748,N_15388,N_15416);
and U15749 (N_15749,N_15259,N_15322);
or U15750 (N_15750,N_15581,N_15653);
and U15751 (N_15751,N_15659,N_15744);
nor U15752 (N_15752,N_15688,N_15730);
and U15753 (N_15753,N_15611,N_15605);
and U15754 (N_15754,N_15643,N_15531);
nand U15755 (N_15755,N_15544,N_15584);
and U15756 (N_15756,N_15525,N_15576);
or U15757 (N_15757,N_15704,N_15500);
and U15758 (N_15758,N_15747,N_15748);
and U15759 (N_15759,N_15509,N_15600);
or U15760 (N_15760,N_15523,N_15626);
nor U15761 (N_15761,N_15502,N_15732);
or U15762 (N_15762,N_15604,N_15568);
nand U15763 (N_15763,N_15705,N_15519);
nor U15764 (N_15764,N_15521,N_15571);
and U15765 (N_15765,N_15725,N_15634);
nor U15766 (N_15766,N_15669,N_15516);
nor U15767 (N_15767,N_15654,N_15520);
nand U15768 (N_15768,N_15529,N_15570);
and U15769 (N_15769,N_15560,N_15559);
nor U15770 (N_15770,N_15577,N_15713);
nand U15771 (N_15771,N_15565,N_15590);
nand U15772 (N_15772,N_15681,N_15506);
nand U15773 (N_15773,N_15627,N_15679);
nor U15774 (N_15774,N_15698,N_15632);
nor U15775 (N_15775,N_15629,N_15670);
nor U15776 (N_15776,N_15682,N_15586);
nor U15777 (N_15777,N_15539,N_15623);
or U15778 (N_15778,N_15512,N_15716);
or U15779 (N_15779,N_15518,N_15655);
nor U15780 (N_15780,N_15625,N_15697);
and U15781 (N_15781,N_15552,N_15667);
nand U15782 (N_15782,N_15622,N_15660);
or U15783 (N_15783,N_15657,N_15551);
and U15784 (N_15784,N_15609,N_15646);
nand U15785 (N_15785,N_15612,N_15537);
nor U15786 (N_15786,N_15595,N_15515);
nor U15787 (N_15787,N_15592,N_15596);
xnor U15788 (N_15788,N_15566,N_15749);
nand U15789 (N_15789,N_15714,N_15666);
and U15790 (N_15790,N_15610,N_15556);
nor U15791 (N_15791,N_15532,N_15517);
nor U15792 (N_15792,N_15553,N_15648);
or U15793 (N_15793,N_15637,N_15583);
nor U15794 (N_15794,N_15664,N_15734);
nor U15795 (N_15795,N_15696,N_15633);
nor U15796 (N_15796,N_15618,N_15613);
xnor U15797 (N_15797,N_15687,N_15593);
and U15798 (N_15798,N_15547,N_15673);
or U15799 (N_15799,N_15724,N_15630);
and U15800 (N_15800,N_15603,N_15614);
nor U15801 (N_15801,N_15639,N_15642);
and U15802 (N_15802,N_15700,N_15574);
nand U15803 (N_15803,N_15522,N_15636);
nand U15804 (N_15804,N_15645,N_15501);
nor U15805 (N_15805,N_15615,N_15649);
or U15806 (N_15806,N_15672,N_15675);
or U15807 (N_15807,N_15695,N_15647);
nand U15808 (N_15808,N_15685,N_15699);
and U15809 (N_15809,N_15567,N_15662);
and U15810 (N_15810,N_15710,N_15683);
nor U15811 (N_15811,N_15534,N_15686);
nor U15812 (N_15812,N_15737,N_15510);
and U15813 (N_15813,N_15694,N_15651);
nand U15814 (N_15814,N_15526,N_15650);
nand U15815 (N_15815,N_15527,N_15591);
and U15816 (N_15816,N_15652,N_15735);
nor U15817 (N_15817,N_15594,N_15663);
or U15818 (N_15818,N_15671,N_15569);
and U15819 (N_15819,N_15739,N_15691);
and U15820 (N_15820,N_15508,N_15720);
or U15821 (N_15821,N_15578,N_15674);
nor U15822 (N_15822,N_15729,N_15541);
and U15823 (N_15823,N_15665,N_15740);
nor U15824 (N_15824,N_15514,N_15719);
nand U15825 (N_15825,N_15545,N_15535);
and U15826 (N_15826,N_15606,N_15741);
or U15827 (N_15827,N_15558,N_15661);
and U15828 (N_15828,N_15589,N_15538);
nor U15829 (N_15829,N_15706,N_15728);
and U15830 (N_15830,N_15738,N_15548);
and U15831 (N_15831,N_15621,N_15597);
nor U15832 (N_15832,N_15717,N_15693);
or U15833 (N_15833,N_15587,N_15533);
nor U15834 (N_15834,N_15546,N_15680);
nand U15835 (N_15835,N_15746,N_15689);
nor U15836 (N_15836,N_15736,N_15715);
or U15837 (N_15837,N_15635,N_15550);
nor U15838 (N_15838,N_15555,N_15709);
nor U15839 (N_15839,N_15608,N_15563);
and U15840 (N_15840,N_15677,N_15513);
nor U15841 (N_15841,N_15742,N_15638);
nor U15842 (N_15842,N_15658,N_15505);
and U15843 (N_15843,N_15701,N_15524);
nor U15844 (N_15844,N_15598,N_15644);
nand U15845 (N_15845,N_15540,N_15549);
nand U15846 (N_15846,N_15631,N_15619);
and U15847 (N_15847,N_15718,N_15543);
nor U15848 (N_15848,N_15640,N_15712);
and U15849 (N_15849,N_15572,N_15743);
and U15850 (N_15850,N_15726,N_15708);
and U15851 (N_15851,N_15733,N_15711);
or U15852 (N_15852,N_15504,N_15684);
or U15853 (N_15853,N_15582,N_15690);
and U15854 (N_15854,N_15562,N_15692);
nand U15855 (N_15855,N_15580,N_15617);
nand U15856 (N_15856,N_15745,N_15601);
nand U15857 (N_15857,N_15707,N_15641);
nand U15858 (N_15858,N_15573,N_15678);
or U15859 (N_15859,N_15702,N_15511);
nor U15860 (N_15860,N_15575,N_15624);
and U15861 (N_15861,N_15607,N_15628);
nor U15862 (N_15862,N_15620,N_15721);
nand U15863 (N_15863,N_15676,N_15561);
xor U15864 (N_15864,N_15585,N_15727);
nor U15865 (N_15865,N_15731,N_15536);
nand U15866 (N_15866,N_15579,N_15530);
or U15867 (N_15867,N_15557,N_15507);
nor U15868 (N_15868,N_15722,N_15599);
or U15869 (N_15869,N_15668,N_15588);
nand U15870 (N_15870,N_15723,N_15602);
or U15871 (N_15871,N_15503,N_15703);
nor U15872 (N_15872,N_15554,N_15564);
nor U15873 (N_15873,N_15616,N_15542);
and U15874 (N_15874,N_15656,N_15528);
nor U15875 (N_15875,N_15605,N_15507);
nor U15876 (N_15876,N_15614,N_15628);
nand U15877 (N_15877,N_15711,N_15704);
nor U15878 (N_15878,N_15502,N_15554);
nand U15879 (N_15879,N_15692,N_15575);
xnor U15880 (N_15880,N_15606,N_15684);
and U15881 (N_15881,N_15744,N_15738);
or U15882 (N_15882,N_15558,N_15731);
or U15883 (N_15883,N_15582,N_15558);
nand U15884 (N_15884,N_15671,N_15659);
and U15885 (N_15885,N_15589,N_15621);
or U15886 (N_15886,N_15557,N_15717);
or U15887 (N_15887,N_15636,N_15529);
and U15888 (N_15888,N_15734,N_15745);
nor U15889 (N_15889,N_15712,N_15672);
nor U15890 (N_15890,N_15604,N_15677);
or U15891 (N_15891,N_15504,N_15557);
nand U15892 (N_15892,N_15553,N_15658);
nor U15893 (N_15893,N_15512,N_15601);
or U15894 (N_15894,N_15731,N_15664);
nand U15895 (N_15895,N_15574,N_15569);
or U15896 (N_15896,N_15592,N_15580);
and U15897 (N_15897,N_15620,N_15678);
nor U15898 (N_15898,N_15578,N_15569);
and U15899 (N_15899,N_15647,N_15634);
or U15900 (N_15900,N_15623,N_15725);
nand U15901 (N_15901,N_15546,N_15528);
nor U15902 (N_15902,N_15560,N_15529);
nand U15903 (N_15903,N_15583,N_15580);
nor U15904 (N_15904,N_15640,N_15520);
or U15905 (N_15905,N_15563,N_15735);
nand U15906 (N_15906,N_15530,N_15549);
or U15907 (N_15907,N_15550,N_15672);
nand U15908 (N_15908,N_15551,N_15600);
or U15909 (N_15909,N_15585,N_15525);
nand U15910 (N_15910,N_15662,N_15512);
nand U15911 (N_15911,N_15528,N_15561);
or U15912 (N_15912,N_15575,N_15538);
nor U15913 (N_15913,N_15594,N_15629);
or U15914 (N_15914,N_15740,N_15598);
nand U15915 (N_15915,N_15598,N_15691);
or U15916 (N_15916,N_15541,N_15717);
nor U15917 (N_15917,N_15564,N_15570);
or U15918 (N_15918,N_15636,N_15554);
nand U15919 (N_15919,N_15607,N_15604);
or U15920 (N_15920,N_15615,N_15735);
nand U15921 (N_15921,N_15713,N_15637);
or U15922 (N_15922,N_15626,N_15556);
nand U15923 (N_15923,N_15737,N_15720);
nand U15924 (N_15924,N_15537,N_15728);
or U15925 (N_15925,N_15650,N_15700);
nor U15926 (N_15926,N_15623,N_15518);
nand U15927 (N_15927,N_15607,N_15570);
or U15928 (N_15928,N_15711,N_15715);
nor U15929 (N_15929,N_15745,N_15700);
nand U15930 (N_15930,N_15518,N_15735);
nor U15931 (N_15931,N_15635,N_15698);
nand U15932 (N_15932,N_15743,N_15563);
nor U15933 (N_15933,N_15629,N_15707);
or U15934 (N_15934,N_15608,N_15558);
nand U15935 (N_15935,N_15631,N_15680);
and U15936 (N_15936,N_15543,N_15582);
and U15937 (N_15937,N_15644,N_15625);
or U15938 (N_15938,N_15561,N_15549);
or U15939 (N_15939,N_15571,N_15589);
nand U15940 (N_15940,N_15584,N_15645);
and U15941 (N_15941,N_15578,N_15749);
nand U15942 (N_15942,N_15537,N_15693);
nor U15943 (N_15943,N_15719,N_15700);
and U15944 (N_15944,N_15715,N_15633);
nor U15945 (N_15945,N_15577,N_15515);
and U15946 (N_15946,N_15747,N_15693);
nand U15947 (N_15947,N_15628,N_15659);
or U15948 (N_15948,N_15656,N_15722);
nand U15949 (N_15949,N_15599,N_15732);
and U15950 (N_15950,N_15634,N_15652);
or U15951 (N_15951,N_15717,N_15661);
nor U15952 (N_15952,N_15515,N_15624);
or U15953 (N_15953,N_15586,N_15518);
nand U15954 (N_15954,N_15643,N_15745);
nor U15955 (N_15955,N_15638,N_15549);
or U15956 (N_15956,N_15618,N_15684);
and U15957 (N_15957,N_15622,N_15700);
nand U15958 (N_15958,N_15605,N_15716);
or U15959 (N_15959,N_15734,N_15507);
and U15960 (N_15960,N_15607,N_15552);
nand U15961 (N_15961,N_15660,N_15530);
or U15962 (N_15962,N_15683,N_15637);
or U15963 (N_15963,N_15567,N_15747);
and U15964 (N_15964,N_15739,N_15743);
nor U15965 (N_15965,N_15719,N_15729);
and U15966 (N_15966,N_15586,N_15669);
and U15967 (N_15967,N_15500,N_15535);
nand U15968 (N_15968,N_15639,N_15624);
or U15969 (N_15969,N_15632,N_15736);
and U15970 (N_15970,N_15553,N_15591);
or U15971 (N_15971,N_15531,N_15652);
nand U15972 (N_15972,N_15594,N_15725);
nand U15973 (N_15973,N_15560,N_15679);
nand U15974 (N_15974,N_15688,N_15749);
or U15975 (N_15975,N_15505,N_15733);
nand U15976 (N_15976,N_15576,N_15578);
and U15977 (N_15977,N_15640,N_15603);
or U15978 (N_15978,N_15719,N_15624);
nor U15979 (N_15979,N_15553,N_15631);
and U15980 (N_15980,N_15612,N_15679);
nor U15981 (N_15981,N_15668,N_15638);
and U15982 (N_15982,N_15658,N_15689);
nor U15983 (N_15983,N_15515,N_15616);
xnor U15984 (N_15984,N_15588,N_15548);
and U15985 (N_15985,N_15543,N_15516);
nand U15986 (N_15986,N_15666,N_15622);
and U15987 (N_15987,N_15728,N_15667);
nor U15988 (N_15988,N_15624,N_15507);
nand U15989 (N_15989,N_15706,N_15732);
nand U15990 (N_15990,N_15565,N_15725);
or U15991 (N_15991,N_15506,N_15710);
and U15992 (N_15992,N_15533,N_15677);
and U15993 (N_15993,N_15719,N_15710);
nor U15994 (N_15994,N_15627,N_15565);
and U15995 (N_15995,N_15605,N_15624);
or U15996 (N_15996,N_15630,N_15729);
nor U15997 (N_15997,N_15666,N_15551);
nand U15998 (N_15998,N_15522,N_15729);
or U15999 (N_15999,N_15713,N_15732);
nand U16000 (N_16000,N_15808,N_15960);
or U16001 (N_16001,N_15804,N_15967);
nand U16002 (N_16002,N_15957,N_15920);
nor U16003 (N_16003,N_15823,N_15821);
and U16004 (N_16004,N_15914,N_15871);
or U16005 (N_16005,N_15828,N_15803);
and U16006 (N_16006,N_15831,N_15991);
or U16007 (N_16007,N_15979,N_15773);
or U16008 (N_16008,N_15964,N_15981);
and U16009 (N_16009,N_15854,N_15815);
and U16010 (N_16010,N_15949,N_15926);
nand U16011 (N_16011,N_15917,N_15867);
nor U16012 (N_16012,N_15761,N_15904);
and U16013 (N_16013,N_15848,N_15857);
nand U16014 (N_16014,N_15900,N_15916);
nand U16015 (N_16015,N_15787,N_15897);
and U16016 (N_16016,N_15983,N_15886);
and U16017 (N_16017,N_15930,N_15918);
or U16018 (N_16018,N_15766,N_15919);
nor U16019 (N_16019,N_15910,N_15890);
nor U16020 (N_16020,N_15998,N_15781);
nor U16021 (N_16021,N_15801,N_15866);
or U16022 (N_16022,N_15999,N_15845);
or U16023 (N_16023,N_15770,N_15977);
or U16024 (N_16024,N_15868,N_15806);
and U16025 (N_16025,N_15870,N_15956);
nor U16026 (N_16026,N_15975,N_15984);
nand U16027 (N_16027,N_15946,N_15836);
nand U16028 (N_16028,N_15753,N_15938);
nand U16029 (N_16029,N_15997,N_15853);
or U16030 (N_16030,N_15833,N_15811);
nor U16031 (N_16031,N_15896,N_15909);
nand U16032 (N_16032,N_15860,N_15915);
or U16033 (N_16033,N_15779,N_15951);
or U16034 (N_16034,N_15783,N_15762);
nand U16035 (N_16035,N_15832,N_15769);
or U16036 (N_16036,N_15844,N_15954);
nor U16037 (N_16037,N_15767,N_15934);
nor U16038 (N_16038,N_15862,N_15978);
xor U16039 (N_16039,N_15851,N_15782);
and U16040 (N_16040,N_15986,N_15928);
nor U16041 (N_16041,N_15841,N_15990);
nor U16042 (N_16042,N_15942,N_15838);
or U16043 (N_16043,N_15872,N_15879);
nor U16044 (N_16044,N_15789,N_15813);
nand U16045 (N_16045,N_15825,N_15941);
and U16046 (N_16046,N_15849,N_15893);
or U16047 (N_16047,N_15864,N_15876);
nand U16048 (N_16048,N_15971,N_15797);
nand U16049 (N_16049,N_15795,N_15810);
nand U16050 (N_16050,N_15932,N_15798);
nor U16051 (N_16051,N_15760,N_15993);
nor U16052 (N_16052,N_15976,N_15807);
and U16053 (N_16053,N_15752,N_15935);
and U16054 (N_16054,N_15814,N_15847);
nand U16055 (N_16055,N_15875,N_15771);
and U16056 (N_16056,N_15908,N_15843);
nand U16057 (N_16057,N_15889,N_15772);
nand U16058 (N_16058,N_15765,N_15863);
and U16059 (N_16059,N_15835,N_15922);
or U16060 (N_16060,N_15989,N_15995);
nand U16061 (N_16061,N_15817,N_15775);
and U16062 (N_16062,N_15774,N_15883);
nor U16063 (N_16063,N_15888,N_15834);
and U16064 (N_16064,N_15905,N_15757);
nand U16065 (N_16065,N_15891,N_15840);
nand U16066 (N_16066,N_15961,N_15982);
nand U16067 (N_16067,N_15895,N_15856);
and U16068 (N_16068,N_15755,N_15837);
xnor U16069 (N_16069,N_15933,N_15786);
nor U16070 (N_16070,N_15923,N_15820);
or U16071 (N_16071,N_15792,N_15974);
nand U16072 (N_16072,N_15793,N_15763);
or U16073 (N_16073,N_15819,N_15968);
nand U16074 (N_16074,N_15899,N_15987);
and U16075 (N_16075,N_15855,N_15903);
or U16076 (N_16076,N_15858,N_15940);
or U16077 (N_16077,N_15816,N_15812);
nand U16078 (N_16078,N_15962,N_15965);
and U16079 (N_16079,N_15958,N_15759);
and U16080 (N_16080,N_15796,N_15892);
nand U16081 (N_16081,N_15902,N_15826);
and U16082 (N_16082,N_15877,N_15906);
nand U16083 (N_16083,N_15913,N_15805);
or U16084 (N_16084,N_15980,N_15996);
nand U16085 (N_16085,N_15830,N_15839);
and U16086 (N_16086,N_15788,N_15970);
and U16087 (N_16087,N_15887,N_15850);
or U16088 (N_16088,N_15756,N_15952);
or U16089 (N_16089,N_15776,N_15794);
or U16090 (N_16090,N_15822,N_15754);
nand U16091 (N_16091,N_15925,N_15921);
nor U16092 (N_16092,N_15790,N_15994);
or U16093 (N_16093,N_15947,N_15829);
or U16094 (N_16094,N_15800,N_15791);
or U16095 (N_16095,N_15901,N_15939);
nor U16096 (N_16096,N_15865,N_15907);
nand U16097 (N_16097,N_15972,N_15818);
and U16098 (N_16098,N_15936,N_15912);
nor U16099 (N_16099,N_15885,N_15751);
nand U16100 (N_16100,N_15846,N_15880);
nand U16101 (N_16101,N_15898,N_15882);
nand U16102 (N_16102,N_15861,N_15944);
nor U16103 (N_16103,N_15852,N_15943);
and U16104 (N_16104,N_15924,N_15780);
nand U16105 (N_16105,N_15869,N_15784);
and U16106 (N_16106,N_15824,N_15778);
and U16107 (N_16107,N_15881,N_15955);
and U16108 (N_16108,N_15929,N_15950);
nor U16109 (N_16109,N_15963,N_15948);
nand U16110 (N_16110,N_15842,N_15873);
or U16111 (N_16111,N_15966,N_15809);
nor U16112 (N_16112,N_15827,N_15988);
nor U16113 (N_16113,N_15750,N_15785);
and U16114 (N_16114,N_15764,N_15768);
nor U16115 (N_16115,N_15945,N_15959);
and U16116 (N_16116,N_15874,N_15802);
and U16117 (N_16117,N_15969,N_15878);
or U16118 (N_16118,N_15992,N_15777);
and U16119 (N_16119,N_15799,N_15758);
nand U16120 (N_16120,N_15859,N_15973);
and U16121 (N_16121,N_15884,N_15911);
nor U16122 (N_16122,N_15927,N_15953);
and U16123 (N_16123,N_15894,N_15931);
and U16124 (N_16124,N_15985,N_15937);
nor U16125 (N_16125,N_15787,N_15964);
nor U16126 (N_16126,N_15984,N_15955);
nor U16127 (N_16127,N_15893,N_15757);
and U16128 (N_16128,N_15771,N_15893);
or U16129 (N_16129,N_15928,N_15848);
nand U16130 (N_16130,N_15947,N_15850);
or U16131 (N_16131,N_15819,N_15915);
nand U16132 (N_16132,N_15862,N_15754);
or U16133 (N_16133,N_15922,N_15846);
and U16134 (N_16134,N_15946,N_15791);
nor U16135 (N_16135,N_15967,N_15773);
nand U16136 (N_16136,N_15936,N_15822);
or U16137 (N_16137,N_15814,N_15934);
or U16138 (N_16138,N_15814,N_15920);
nand U16139 (N_16139,N_15890,N_15921);
nor U16140 (N_16140,N_15826,N_15800);
or U16141 (N_16141,N_15954,N_15760);
nor U16142 (N_16142,N_15763,N_15883);
or U16143 (N_16143,N_15830,N_15825);
nand U16144 (N_16144,N_15997,N_15976);
and U16145 (N_16145,N_15908,N_15983);
and U16146 (N_16146,N_15826,N_15973);
nor U16147 (N_16147,N_15866,N_15770);
nor U16148 (N_16148,N_15766,N_15905);
nor U16149 (N_16149,N_15952,N_15789);
and U16150 (N_16150,N_15834,N_15943);
and U16151 (N_16151,N_15926,N_15852);
nor U16152 (N_16152,N_15836,N_15977);
or U16153 (N_16153,N_15957,N_15788);
nand U16154 (N_16154,N_15881,N_15886);
nor U16155 (N_16155,N_15991,N_15985);
nor U16156 (N_16156,N_15951,N_15983);
nor U16157 (N_16157,N_15830,N_15884);
nand U16158 (N_16158,N_15774,N_15750);
nand U16159 (N_16159,N_15773,N_15836);
nor U16160 (N_16160,N_15879,N_15798);
nor U16161 (N_16161,N_15797,N_15893);
and U16162 (N_16162,N_15929,N_15969);
and U16163 (N_16163,N_15990,N_15896);
or U16164 (N_16164,N_15895,N_15833);
and U16165 (N_16165,N_15856,N_15806);
and U16166 (N_16166,N_15793,N_15977);
and U16167 (N_16167,N_15987,N_15970);
nand U16168 (N_16168,N_15835,N_15879);
or U16169 (N_16169,N_15967,N_15839);
or U16170 (N_16170,N_15967,N_15913);
or U16171 (N_16171,N_15878,N_15887);
and U16172 (N_16172,N_15827,N_15899);
nor U16173 (N_16173,N_15787,N_15905);
and U16174 (N_16174,N_15798,N_15838);
nor U16175 (N_16175,N_15897,N_15915);
nand U16176 (N_16176,N_15992,N_15764);
nor U16177 (N_16177,N_15973,N_15947);
or U16178 (N_16178,N_15882,N_15843);
nor U16179 (N_16179,N_15787,N_15840);
or U16180 (N_16180,N_15757,N_15811);
nor U16181 (N_16181,N_15862,N_15933);
nand U16182 (N_16182,N_15958,N_15807);
nor U16183 (N_16183,N_15974,N_15833);
nand U16184 (N_16184,N_15906,N_15829);
and U16185 (N_16185,N_15880,N_15940);
nor U16186 (N_16186,N_15986,N_15796);
or U16187 (N_16187,N_15975,N_15970);
nor U16188 (N_16188,N_15782,N_15822);
and U16189 (N_16189,N_15966,N_15753);
or U16190 (N_16190,N_15871,N_15775);
and U16191 (N_16191,N_15779,N_15833);
and U16192 (N_16192,N_15897,N_15760);
or U16193 (N_16193,N_15886,N_15844);
nor U16194 (N_16194,N_15999,N_15906);
or U16195 (N_16195,N_15934,N_15899);
nand U16196 (N_16196,N_15750,N_15861);
nand U16197 (N_16197,N_15803,N_15829);
and U16198 (N_16198,N_15997,N_15883);
or U16199 (N_16199,N_15752,N_15816);
and U16200 (N_16200,N_15877,N_15787);
and U16201 (N_16201,N_15928,N_15910);
or U16202 (N_16202,N_15967,N_15950);
nand U16203 (N_16203,N_15999,N_15947);
nor U16204 (N_16204,N_15796,N_15847);
nand U16205 (N_16205,N_15970,N_15763);
nor U16206 (N_16206,N_15952,N_15876);
nor U16207 (N_16207,N_15951,N_15988);
nand U16208 (N_16208,N_15816,N_15926);
nand U16209 (N_16209,N_15773,N_15841);
or U16210 (N_16210,N_15844,N_15947);
and U16211 (N_16211,N_15911,N_15788);
nor U16212 (N_16212,N_15850,N_15840);
nor U16213 (N_16213,N_15998,N_15795);
or U16214 (N_16214,N_15877,N_15997);
nor U16215 (N_16215,N_15963,N_15789);
nand U16216 (N_16216,N_15987,N_15890);
nand U16217 (N_16217,N_15903,N_15861);
nand U16218 (N_16218,N_15939,N_15978);
nand U16219 (N_16219,N_15869,N_15974);
nand U16220 (N_16220,N_15992,N_15963);
or U16221 (N_16221,N_15758,N_15764);
or U16222 (N_16222,N_15769,N_15959);
and U16223 (N_16223,N_15965,N_15809);
nand U16224 (N_16224,N_15878,N_15954);
nor U16225 (N_16225,N_15787,N_15774);
or U16226 (N_16226,N_15801,N_15985);
and U16227 (N_16227,N_15758,N_15920);
nand U16228 (N_16228,N_15941,N_15832);
or U16229 (N_16229,N_15762,N_15844);
nor U16230 (N_16230,N_15796,N_15808);
or U16231 (N_16231,N_15863,N_15771);
nand U16232 (N_16232,N_15988,N_15754);
or U16233 (N_16233,N_15909,N_15956);
and U16234 (N_16234,N_15967,N_15929);
nand U16235 (N_16235,N_15767,N_15926);
or U16236 (N_16236,N_15935,N_15892);
nand U16237 (N_16237,N_15864,N_15855);
nand U16238 (N_16238,N_15915,N_15958);
and U16239 (N_16239,N_15959,N_15937);
or U16240 (N_16240,N_15802,N_15758);
nor U16241 (N_16241,N_15907,N_15817);
nand U16242 (N_16242,N_15957,N_15774);
nand U16243 (N_16243,N_15995,N_15802);
nor U16244 (N_16244,N_15945,N_15987);
nand U16245 (N_16245,N_15891,N_15792);
or U16246 (N_16246,N_15752,N_15810);
and U16247 (N_16247,N_15853,N_15756);
and U16248 (N_16248,N_15909,N_15823);
nand U16249 (N_16249,N_15822,N_15801);
nor U16250 (N_16250,N_16117,N_16056);
and U16251 (N_16251,N_16200,N_16193);
nor U16252 (N_16252,N_16137,N_16051);
and U16253 (N_16253,N_16140,N_16170);
nor U16254 (N_16254,N_16009,N_16243);
nor U16255 (N_16255,N_16171,N_16155);
nand U16256 (N_16256,N_16135,N_16153);
nor U16257 (N_16257,N_16145,N_16008);
nor U16258 (N_16258,N_16142,N_16149);
or U16259 (N_16259,N_16078,N_16159);
and U16260 (N_16260,N_16132,N_16129);
and U16261 (N_16261,N_16107,N_16032);
or U16262 (N_16262,N_16033,N_16245);
and U16263 (N_16263,N_16123,N_16229);
and U16264 (N_16264,N_16094,N_16190);
nand U16265 (N_16265,N_16133,N_16103);
nor U16266 (N_16266,N_16226,N_16023);
nor U16267 (N_16267,N_16077,N_16037);
nand U16268 (N_16268,N_16172,N_16246);
and U16269 (N_16269,N_16227,N_16043);
nor U16270 (N_16270,N_16167,N_16218);
nand U16271 (N_16271,N_16191,N_16030);
and U16272 (N_16272,N_16166,N_16247);
nand U16273 (N_16273,N_16144,N_16128);
and U16274 (N_16274,N_16174,N_16138);
nor U16275 (N_16275,N_16163,N_16053);
nor U16276 (N_16276,N_16114,N_16101);
or U16277 (N_16277,N_16160,N_16189);
nor U16278 (N_16278,N_16064,N_16217);
and U16279 (N_16279,N_16231,N_16048);
nor U16280 (N_16280,N_16093,N_16236);
nand U16281 (N_16281,N_16084,N_16109);
nand U16282 (N_16282,N_16062,N_16196);
nand U16283 (N_16283,N_16080,N_16203);
and U16284 (N_16284,N_16201,N_16146);
and U16285 (N_16285,N_16112,N_16039);
nor U16286 (N_16286,N_16106,N_16016);
nor U16287 (N_16287,N_16169,N_16111);
nand U16288 (N_16288,N_16097,N_16240);
and U16289 (N_16289,N_16015,N_16177);
or U16290 (N_16290,N_16225,N_16082);
or U16291 (N_16291,N_16143,N_16052);
nor U16292 (N_16292,N_16206,N_16061);
or U16293 (N_16293,N_16134,N_16024);
nor U16294 (N_16294,N_16184,N_16042);
nand U16295 (N_16295,N_16074,N_16073);
or U16296 (N_16296,N_16248,N_16086);
or U16297 (N_16297,N_16154,N_16083);
or U16298 (N_16298,N_16207,N_16130);
or U16299 (N_16299,N_16025,N_16194);
or U16300 (N_16300,N_16228,N_16105);
nand U16301 (N_16301,N_16058,N_16014);
nor U16302 (N_16302,N_16199,N_16162);
nor U16303 (N_16303,N_16010,N_16113);
or U16304 (N_16304,N_16156,N_16244);
or U16305 (N_16305,N_16183,N_16221);
or U16306 (N_16306,N_16022,N_16213);
or U16307 (N_16307,N_16067,N_16099);
nand U16308 (N_16308,N_16238,N_16029);
or U16309 (N_16309,N_16168,N_16224);
nor U16310 (N_16310,N_16012,N_16188);
or U16311 (N_16311,N_16057,N_16066);
nor U16312 (N_16312,N_16136,N_16076);
nand U16313 (N_16313,N_16204,N_16141);
or U16314 (N_16314,N_16027,N_16045);
or U16315 (N_16315,N_16116,N_16187);
or U16316 (N_16316,N_16148,N_16070);
and U16317 (N_16317,N_16049,N_16063);
and U16318 (N_16318,N_16215,N_16095);
nand U16319 (N_16319,N_16069,N_16002);
or U16320 (N_16320,N_16216,N_16087);
or U16321 (N_16321,N_16249,N_16195);
and U16322 (N_16322,N_16055,N_16031);
nor U16323 (N_16323,N_16054,N_16036);
nand U16324 (N_16324,N_16180,N_16220);
or U16325 (N_16325,N_16185,N_16071);
nand U16326 (N_16326,N_16192,N_16085);
nor U16327 (N_16327,N_16173,N_16234);
nand U16328 (N_16328,N_16041,N_16013);
nor U16329 (N_16329,N_16122,N_16232);
and U16330 (N_16330,N_16222,N_16088);
and U16331 (N_16331,N_16241,N_16219);
nor U16332 (N_16332,N_16235,N_16242);
nand U16333 (N_16333,N_16131,N_16115);
nor U16334 (N_16334,N_16006,N_16104);
or U16335 (N_16335,N_16011,N_16021);
nand U16336 (N_16336,N_16124,N_16157);
nand U16337 (N_16337,N_16050,N_16119);
or U16338 (N_16338,N_16120,N_16026);
nor U16339 (N_16339,N_16202,N_16158);
or U16340 (N_16340,N_16000,N_16072);
nand U16341 (N_16341,N_16210,N_16019);
nand U16342 (N_16342,N_16127,N_16118);
nor U16343 (N_16343,N_16017,N_16059);
nand U16344 (N_16344,N_16100,N_16164);
and U16345 (N_16345,N_16020,N_16239);
and U16346 (N_16346,N_16147,N_16223);
nand U16347 (N_16347,N_16209,N_16197);
or U16348 (N_16348,N_16001,N_16108);
and U16349 (N_16349,N_16208,N_16178);
and U16350 (N_16350,N_16181,N_16151);
and U16351 (N_16351,N_16046,N_16179);
and U16352 (N_16352,N_16007,N_16150);
and U16353 (N_16353,N_16040,N_16152);
or U16354 (N_16354,N_16186,N_16237);
and U16355 (N_16355,N_16003,N_16211);
or U16356 (N_16356,N_16092,N_16176);
or U16357 (N_16357,N_16102,N_16165);
or U16358 (N_16358,N_16125,N_16233);
and U16359 (N_16359,N_16081,N_16126);
and U16360 (N_16360,N_16175,N_16047);
nor U16361 (N_16361,N_16161,N_16090);
nand U16362 (N_16362,N_16205,N_16075);
nor U16363 (N_16363,N_16121,N_16018);
nand U16364 (N_16364,N_16230,N_16198);
nor U16365 (N_16365,N_16098,N_16035);
nand U16366 (N_16366,N_16214,N_16065);
nor U16367 (N_16367,N_16004,N_16038);
nor U16368 (N_16368,N_16068,N_16182);
nor U16369 (N_16369,N_16060,N_16212);
and U16370 (N_16370,N_16034,N_16079);
and U16371 (N_16371,N_16139,N_16028);
nand U16372 (N_16372,N_16044,N_16110);
nor U16373 (N_16373,N_16005,N_16091);
or U16374 (N_16374,N_16089,N_16096);
and U16375 (N_16375,N_16229,N_16140);
or U16376 (N_16376,N_16175,N_16022);
nand U16377 (N_16377,N_16015,N_16169);
or U16378 (N_16378,N_16043,N_16204);
or U16379 (N_16379,N_16070,N_16206);
nor U16380 (N_16380,N_16190,N_16145);
nor U16381 (N_16381,N_16035,N_16166);
nand U16382 (N_16382,N_16122,N_16156);
xor U16383 (N_16383,N_16027,N_16005);
nand U16384 (N_16384,N_16148,N_16063);
nor U16385 (N_16385,N_16142,N_16187);
and U16386 (N_16386,N_16244,N_16168);
nor U16387 (N_16387,N_16240,N_16214);
nor U16388 (N_16388,N_16006,N_16168);
nand U16389 (N_16389,N_16072,N_16248);
nor U16390 (N_16390,N_16086,N_16203);
nor U16391 (N_16391,N_16226,N_16200);
nand U16392 (N_16392,N_16017,N_16218);
nor U16393 (N_16393,N_16064,N_16224);
and U16394 (N_16394,N_16093,N_16066);
and U16395 (N_16395,N_16124,N_16029);
and U16396 (N_16396,N_16238,N_16128);
nor U16397 (N_16397,N_16104,N_16147);
or U16398 (N_16398,N_16167,N_16207);
and U16399 (N_16399,N_16229,N_16058);
and U16400 (N_16400,N_16100,N_16065);
and U16401 (N_16401,N_16097,N_16223);
nand U16402 (N_16402,N_16161,N_16152);
or U16403 (N_16403,N_16203,N_16196);
or U16404 (N_16404,N_16018,N_16117);
or U16405 (N_16405,N_16048,N_16059);
and U16406 (N_16406,N_16177,N_16187);
nand U16407 (N_16407,N_16193,N_16209);
or U16408 (N_16408,N_16045,N_16203);
and U16409 (N_16409,N_16089,N_16162);
nor U16410 (N_16410,N_16049,N_16107);
or U16411 (N_16411,N_16114,N_16200);
nand U16412 (N_16412,N_16068,N_16127);
or U16413 (N_16413,N_16221,N_16242);
and U16414 (N_16414,N_16103,N_16138);
nand U16415 (N_16415,N_16042,N_16044);
nand U16416 (N_16416,N_16063,N_16096);
and U16417 (N_16417,N_16233,N_16146);
and U16418 (N_16418,N_16004,N_16205);
nand U16419 (N_16419,N_16057,N_16070);
and U16420 (N_16420,N_16218,N_16203);
nand U16421 (N_16421,N_16022,N_16043);
nor U16422 (N_16422,N_16242,N_16126);
and U16423 (N_16423,N_16003,N_16239);
nand U16424 (N_16424,N_16164,N_16129);
or U16425 (N_16425,N_16124,N_16056);
or U16426 (N_16426,N_16016,N_16000);
and U16427 (N_16427,N_16203,N_16109);
and U16428 (N_16428,N_16201,N_16207);
nand U16429 (N_16429,N_16141,N_16201);
or U16430 (N_16430,N_16249,N_16236);
nor U16431 (N_16431,N_16021,N_16004);
or U16432 (N_16432,N_16060,N_16247);
or U16433 (N_16433,N_16187,N_16205);
nand U16434 (N_16434,N_16024,N_16043);
or U16435 (N_16435,N_16010,N_16212);
nand U16436 (N_16436,N_16021,N_16040);
and U16437 (N_16437,N_16118,N_16207);
or U16438 (N_16438,N_16062,N_16113);
nor U16439 (N_16439,N_16061,N_16052);
and U16440 (N_16440,N_16217,N_16014);
and U16441 (N_16441,N_16063,N_16117);
xnor U16442 (N_16442,N_16154,N_16199);
nor U16443 (N_16443,N_16075,N_16226);
or U16444 (N_16444,N_16199,N_16107);
nand U16445 (N_16445,N_16208,N_16168);
or U16446 (N_16446,N_16127,N_16097);
nor U16447 (N_16447,N_16174,N_16228);
xnor U16448 (N_16448,N_16215,N_16193);
nor U16449 (N_16449,N_16217,N_16112);
or U16450 (N_16450,N_16215,N_16223);
nand U16451 (N_16451,N_16232,N_16076);
nor U16452 (N_16452,N_16162,N_16004);
or U16453 (N_16453,N_16180,N_16107);
xnor U16454 (N_16454,N_16116,N_16093);
and U16455 (N_16455,N_16115,N_16054);
and U16456 (N_16456,N_16031,N_16174);
or U16457 (N_16457,N_16037,N_16019);
and U16458 (N_16458,N_16129,N_16223);
xor U16459 (N_16459,N_16037,N_16204);
xnor U16460 (N_16460,N_16247,N_16104);
nor U16461 (N_16461,N_16101,N_16218);
and U16462 (N_16462,N_16001,N_16231);
and U16463 (N_16463,N_16169,N_16070);
nor U16464 (N_16464,N_16159,N_16166);
and U16465 (N_16465,N_16103,N_16130);
or U16466 (N_16466,N_16217,N_16201);
and U16467 (N_16467,N_16025,N_16154);
or U16468 (N_16468,N_16179,N_16217);
nand U16469 (N_16469,N_16056,N_16179);
and U16470 (N_16470,N_16203,N_16244);
and U16471 (N_16471,N_16017,N_16070);
nor U16472 (N_16472,N_16103,N_16248);
and U16473 (N_16473,N_16038,N_16019);
nand U16474 (N_16474,N_16069,N_16242);
nand U16475 (N_16475,N_16220,N_16006);
nand U16476 (N_16476,N_16123,N_16019);
and U16477 (N_16477,N_16171,N_16090);
and U16478 (N_16478,N_16023,N_16186);
xor U16479 (N_16479,N_16128,N_16235);
nor U16480 (N_16480,N_16101,N_16056);
and U16481 (N_16481,N_16183,N_16099);
nor U16482 (N_16482,N_16233,N_16029);
nand U16483 (N_16483,N_16049,N_16219);
and U16484 (N_16484,N_16026,N_16158);
nand U16485 (N_16485,N_16100,N_16234);
or U16486 (N_16486,N_16236,N_16036);
or U16487 (N_16487,N_16105,N_16136);
and U16488 (N_16488,N_16127,N_16086);
and U16489 (N_16489,N_16111,N_16068);
nor U16490 (N_16490,N_16051,N_16080);
and U16491 (N_16491,N_16135,N_16058);
or U16492 (N_16492,N_16070,N_16078);
or U16493 (N_16493,N_16134,N_16246);
nor U16494 (N_16494,N_16008,N_16082);
nor U16495 (N_16495,N_16055,N_16077);
nor U16496 (N_16496,N_16093,N_16175);
or U16497 (N_16497,N_16173,N_16171);
nor U16498 (N_16498,N_16200,N_16132);
and U16499 (N_16499,N_16142,N_16239);
or U16500 (N_16500,N_16313,N_16391);
nand U16501 (N_16501,N_16264,N_16452);
and U16502 (N_16502,N_16483,N_16438);
nand U16503 (N_16503,N_16300,N_16304);
nor U16504 (N_16504,N_16322,N_16494);
nand U16505 (N_16505,N_16498,N_16403);
and U16506 (N_16506,N_16473,N_16426);
or U16507 (N_16507,N_16307,N_16318);
nand U16508 (N_16508,N_16436,N_16326);
nand U16509 (N_16509,N_16456,N_16309);
nor U16510 (N_16510,N_16476,N_16298);
or U16511 (N_16511,N_16332,N_16464);
and U16512 (N_16512,N_16336,N_16489);
and U16513 (N_16513,N_16497,N_16370);
nand U16514 (N_16514,N_16375,N_16358);
nor U16515 (N_16515,N_16422,N_16439);
or U16516 (N_16516,N_16339,N_16496);
nor U16517 (N_16517,N_16351,N_16435);
nor U16518 (N_16518,N_16257,N_16325);
and U16519 (N_16519,N_16287,N_16294);
nor U16520 (N_16520,N_16386,N_16285);
nor U16521 (N_16521,N_16335,N_16470);
and U16522 (N_16522,N_16493,N_16341);
nand U16523 (N_16523,N_16297,N_16319);
or U16524 (N_16524,N_16434,N_16327);
and U16525 (N_16525,N_16475,N_16295);
and U16526 (N_16526,N_16468,N_16357);
and U16527 (N_16527,N_16479,N_16273);
nand U16528 (N_16528,N_16306,N_16372);
or U16529 (N_16529,N_16381,N_16465);
nor U16530 (N_16530,N_16344,N_16281);
or U16531 (N_16531,N_16413,N_16412);
nor U16532 (N_16532,N_16286,N_16352);
or U16533 (N_16533,N_16474,N_16384);
nor U16534 (N_16534,N_16356,N_16459);
nand U16535 (N_16535,N_16291,N_16427);
nand U16536 (N_16536,N_16308,N_16329);
or U16537 (N_16537,N_16311,N_16333);
or U16538 (N_16538,N_16283,N_16280);
and U16539 (N_16539,N_16272,N_16274);
nand U16540 (N_16540,N_16383,N_16278);
nor U16541 (N_16541,N_16312,N_16380);
nand U16542 (N_16542,N_16440,N_16321);
and U16543 (N_16543,N_16261,N_16362);
nand U16544 (N_16544,N_16346,N_16293);
or U16545 (N_16545,N_16446,N_16367);
and U16546 (N_16546,N_16348,N_16394);
or U16547 (N_16547,N_16451,N_16414);
or U16548 (N_16548,N_16487,N_16328);
and U16549 (N_16549,N_16392,N_16491);
or U16550 (N_16550,N_16292,N_16419);
or U16551 (N_16551,N_16461,N_16482);
and U16552 (N_16552,N_16423,N_16431);
nand U16553 (N_16553,N_16404,N_16396);
nand U16554 (N_16554,N_16428,N_16277);
and U16555 (N_16555,N_16365,N_16447);
nor U16556 (N_16556,N_16266,N_16499);
nand U16557 (N_16557,N_16323,N_16421);
nand U16558 (N_16558,N_16441,N_16387);
and U16559 (N_16559,N_16405,N_16402);
nand U16560 (N_16560,N_16444,N_16296);
nand U16561 (N_16561,N_16276,N_16409);
nor U16562 (N_16562,N_16455,N_16466);
or U16563 (N_16563,N_16477,N_16364);
xnor U16564 (N_16564,N_16343,N_16418);
xnor U16565 (N_16565,N_16393,N_16347);
or U16566 (N_16566,N_16263,N_16400);
and U16567 (N_16567,N_16432,N_16262);
nand U16568 (N_16568,N_16288,N_16317);
nor U16569 (N_16569,N_16401,N_16271);
and U16570 (N_16570,N_16349,N_16254);
nand U16571 (N_16571,N_16495,N_16429);
and U16572 (N_16572,N_16270,N_16361);
and U16573 (N_16573,N_16299,N_16467);
or U16574 (N_16574,N_16484,N_16469);
and U16575 (N_16575,N_16315,N_16488);
and U16576 (N_16576,N_16450,N_16269);
and U16577 (N_16577,N_16345,N_16268);
nand U16578 (N_16578,N_16279,N_16478);
nand U16579 (N_16579,N_16267,N_16282);
nand U16580 (N_16580,N_16457,N_16472);
nand U16581 (N_16581,N_16453,N_16250);
or U16582 (N_16582,N_16331,N_16260);
nand U16583 (N_16583,N_16442,N_16486);
nand U16584 (N_16584,N_16363,N_16355);
and U16585 (N_16585,N_16310,N_16462);
nor U16586 (N_16586,N_16395,N_16373);
or U16587 (N_16587,N_16303,N_16360);
and U16588 (N_16588,N_16256,N_16354);
nand U16589 (N_16589,N_16259,N_16424);
nor U16590 (N_16590,N_16338,N_16397);
and U16591 (N_16591,N_16284,N_16492);
nor U16592 (N_16592,N_16342,N_16289);
and U16593 (N_16593,N_16337,N_16471);
and U16594 (N_16594,N_16371,N_16454);
or U16595 (N_16595,N_16406,N_16350);
and U16596 (N_16596,N_16377,N_16265);
nor U16597 (N_16597,N_16382,N_16340);
nand U16598 (N_16598,N_16252,N_16445);
xnor U16599 (N_16599,N_16407,N_16378);
nor U16600 (N_16600,N_16388,N_16458);
and U16601 (N_16601,N_16334,N_16425);
and U16602 (N_16602,N_16390,N_16314);
nand U16603 (N_16603,N_16430,N_16253);
nand U16604 (N_16604,N_16290,N_16369);
nand U16605 (N_16605,N_16316,N_16376);
or U16606 (N_16606,N_16353,N_16389);
or U16607 (N_16607,N_16330,N_16411);
nor U16608 (N_16608,N_16408,N_16255);
or U16609 (N_16609,N_16368,N_16379);
and U16610 (N_16610,N_16448,N_16443);
or U16611 (N_16611,N_16480,N_16251);
nor U16612 (N_16612,N_16359,N_16415);
or U16613 (N_16613,N_16301,N_16420);
and U16614 (N_16614,N_16305,N_16410);
or U16615 (N_16615,N_16433,N_16324);
or U16616 (N_16616,N_16374,N_16366);
nor U16617 (N_16617,N_16463,N_16416);
or U16618 (N_16618,N_16481,N_16449);
nand U16619 (N_16619,N_16275,N_16490);
nand U16620 (N_16620,N_16385,N_16258);
or U16621 (N_16621,N_16460,N_16417);
nand U16622 (N_16622,N_16485,N_16320);
nor U16623 (N_16623,N_16302,N_16398);
nor U16624 (N_16624,N_16399,N_16437);
and U16625 (N_16625,N_16470,N_16350);
or U16626 (N_16626,N_16276,N_16327);
and U16627 (N_16627,N_16437,N_16357);
and U16628 (N_16628,N_16273,N_16445);
nand U16629 (N_16629,N_16395,N_16325);
and U16630 (N_16630,N_16489,N_16299);
nand U16631 (N_16631,N_16282,N_16262);
nor U16632 (N_16632,N_16286,N_16365);
and U16633 (N_16633,N_16456,N_16432);
and U16634 (N_16634,N_16497,N_16273);
or U16635 (N_16635,N_16360,N_16423);
nand U16636 (N_16636,N_16331,N_16251);
or U16637 (N_16637,N_16384,N_16303);
nand U16638 (N_16638,N_16463,N_16438);
nor U16639 (N_16639,N_16460,N_16311);
nand U16640 (N_16640,N_16431,N_16482);
and U16641 (N_16641,N_16312,N_16447);
and U16642 (N_16642,N_16321,N_16330);
nor U16643 (N_16643,N_16315,N_16314);
or U16644 (N_16644,N_16269,N_16437);
nor U16645 (N_16645,N_16377,N_16327);
nand U16646 (N_16646,N_16292,N_16338);
nor U16647 (N_16647,N_16302,N_16418);
or U16648 (N_16648,N_16473,N_16452);
or U16649 (N_16649,N_16298,N_16477);
nor U16650 (N_16650,N_16311,N_16455);
nor U16651 (N_16651,N_16256,N_16447);
or U16652 (N_16652,N_16320,N_16300);
nand U16653 (N_16653,N_16341,N_16281);
or U16654 (N_16654,N_16311,N_16322);
nand U16655 (N_16655,N_16477,N_16403);
nand U16656 (N_16656,N_16250,N_16386);
and U16657 (N_16657,N_16458,N_16367);
nand U16658 (N_16658,N_16359,N_16476);
or U16659 (N_16659,N_16335,N_16368);
or U16660 (N_16660,N_16472,N_16257);
nor U16661 (N_16661,N_16407,N_16477);
and U16662 (N_16662,N_16471,N_16329);
nor U16663 (N_16663,N_16356,N_16304);
and U16664 (N_16664,N_16409,N_16463);
nor U16665 (N_16665,N_16476,N_16469);
or U16666 (N_16666,N_16411,N_16486);
nor U16667 (N_16667,N_16279,N_16283);
nor U16668 (N_16668,N_16299,N_16355);
nor U16669 (N_16669,N_16279,N_16463);
nand U16670 (N_16670,N_16372,N_16300);
or U16671 (N_16671,N_16437,N_16471);
xnor U16672 (N_16672,N_16404,N_16358);
nand U16673 (N_16673,N_16400,N_16314);
nor U16674 (N_16674,N_16441,N_16313);
nor U16675 (N_16675,N_16355,N_16430);
nand U16676 (N_16676,N_16381,N_16428);
or U16677 (N_16677,N_16433,N_16482);
nand U16678 (N_16678,N_16382,N_16413);
or U16679 (N_16679,N_16297,N_16490);
or U16680 (N_16680,N_16431,N_16252);
or U16681 (N_16681,N_16304,N_16345);
nor U16682 (N_16682,N_16269,N_16315);
nand U16683 (N_16683,N_16424,N_16282);
or U16684 (N_16684,N_16317,N_16320);
or U16685 (N_16685,N_16393,N_16488);
and U16686 (N_16686,N_16380,N_16444);
nand U16687 (N_16687,N_16387,N_16356);
nor U16688 (N_16688,N_16420,N_16399);
nand U16689 (N_16689,N_16433,N_16460);
nand U16690 (N_16690,N_16485,N_16431);
or U16691 (N_16691,N_16409,N_16356);
nand U16692 (N_16692,N_16275,N_16322);
or U16693 (N_16693,N_16479,N_16266);
nand U16694 (N_16694,N_16260,N_16278);
nor U16695 (N_16695,N_16255,N_16484);
nand U16696 (N_16696,N_16488,N_16462);
nand U16697 (N_16697,N_16289,N_16499);
nor U16698 (N_16698,N_16412,N_16422);
nand U16699 (N_16699,N_16419,N_16386);
nor U16700 (N_16700,N_16324,N_16473);
nor U16701 (N_16701,N_16435,N_16326);
or U16702 (N_16702,N_16375,N_16433);
nor U16703 (N_16703,N_16360,N_16430);
or U16704 (N_16704,N_16363,N_16264);
or U16705 (N_16705,N_16345,N_16466);
and U16706 (N_16706,N_16293,N_16343);
or U16707 (N_16707,N_16381,N_16302);
and U16708 (N_16708,N_16311,N_16268);
and U16709 (N_16709,N_16366,N_16365);
or U16710 (N_16710,N_16455,N_16360);
nor U16711 (N_16711,N_16482,N_16465);
nor U16712 (N_16712,N_16441,N_16412);
or U16713 (N_16713,N_16425,N_16280);
nor U16714 (N_16714,N_16319,N_16381);
or U16715 (N_16715,N_16431,N_16348);
nor U16716 (N_16716,N_16269,N_16422);
or U16717 (N_16717,N_16297,N_16405);
nand U16718 (N_16718,N_16408,N_16440);
nor U16719 (N_16719,N_16436,N_16442);
and U16720 (N_16720,N_16491,N_16270);
and U16721 (N_16721,N_16321,N_16264);
nand U16722 (N_16722,N_16403,N_16431);
and U16723 (N_16723,N_16439,N_16330);
and U16724 (N_16724,N_16292,N_16255);
or U16725 (N_16725,N_16493,N_16266);
nand U16726 (N_16726,N_16294,N_16322);
and U16727 (N_16727,N_16398,N_16360);
and U16728 (N_16728,N_16440,N_16300);
or U16729 (N_16729,N_16327,N_16355);
or U16730 (N_16730,N_16403,N_16379);
and U16731 (N_16731,N_16481,N_16306);
or U16732 (N_16732,N_16481,N_16421);
and U16733 (N_16733,N_16429,N_16271);
or U16734 (N_16734,N_16349,N_16408);
nand U16735 (N_16735,N_16255,N_16318);
nor U16736 (N_16736,N_16427,N_16406);
nand U16737 (N_16737,N_16306,N_16478);
nand U16738 (N_16738,N_16359,N_16327);
nor U16739 (N_16739,N_16470,N_16288);
and U16740 (N_16740,N_16438,N_16300);
nand U16741 (N_16741,N_16415,N_16266);
nand U16742 (N_16742,N_16339,N_16449);
and U16743 (N_16743,N_16266,N_16400);
or U16744 (N_16744,N_16333,N_16430);
nand U16745 (N_16745,N_16418,N_16308);
and U16746 (N_16746,N_16350,N_16410);
nor U16747 (N_16747,N_16342,N_16467);
nor U16748 (N_16748,N_16286,N_16298);
nor U16749 (N_16749,N_16439,N_16364);
and U16750 (N_16750,N_16600,N_16599);
and U16751 (N_16751,N_16547,N_16597);
nor U16752 (N_16752,N_16728,N_16591);
nor U16753 (N_16753,N_16543,N_16735);
nor U16754 (N_16754,N_16635,N_16640);
or U16755 (N_16755,N_16573,N_16738);
nand U16756 (N_16756,N_16690,N_16523);
and U16757 (N_16757,N_16682,N_16525);
xnor U16758 (N_16758,N_16616,N_16664);
or U16759 (N_16759,N_16535,N_16565);
and U16760 (N_16760,N_16702,N_16617);
nand U16761 (N_16761,N_16744,N_16716);
or U16762 (N_16762,N_16522,N_16549);
nor U16763 (N_16763,N_16646,N_16688);
and U16764 (N_16764,N_16604,N_16677);
or U16765 (N_16765,N_16579,N_16590);
or U16766 (N_16766,N_16671,N_16595);
or U16767 (N_16767,N_16727,N_16734);
and U16768 (N_16768,N_16540,N_16627);
nand U16769 (N_16769,N_16584,N_16655);
and U16770 (N_16770,N_16569,N_16504);
xor U16771 (N_16771,N_16634,N_16544);
and U16772 (N_16772,N_16647,N_16656);
or U16773 (N_16773,N_16726,N_16680);
or U16774 (N_16774,N_16662,N_16737);
and U16775 (N_16775,N_16675,N_16511);
nor U16776 (N_16776,N_16562,N_16648);
and U16777 (N_16777,N_16629,N_16636);
nor U16778 (N_16778,N_16620,N_16577);
and U16779 (N_16779,N_16564,N_16615);
nand U16780 (N_16780,N_16623,N_16739);
and U16781 (N_16781,N_16588,N_16524);
nor U16782 (N_16782,N_16505,N_16742);
or U16783 (N_16783,N_16566,N_16575);
or U16784 (N_16784,N_16678,N_16542);
nor U16785 (N_16785,N_16691,N_16657);
nand U16786 (N_16786,N_16710,N_16606);
or U16787 (N_16787,N_16673,N_16619);
and U16788 (N_16788,N_16707,N_16663);
nor U16789 (N_16789,N_16724,N_16696);
nand U16790 (N_16790,N_16510,N_16743);
nand U16791 (N_16791,N_16731,N_16500);
nand U16792 (N_16792,N_16512,N_16693);
and U16793 (N_16793,N_16557,N_16704);
or U16794 (N_16794,N_16695,N_16637);
nand U16795 (N_16795,N_16578,N_16503);
nand U16796 (N_16796,N_16709,N_16536);
nor U16797 (N_16797,N_16558,N_16713);
nand U16798 (N_16798,N_16592,N_16618);
or U16799 (N_16799,N_16674,N_16596);
nand U16800 (N_16800,N_16659,N_16633);
and U16801 (N_16801,N_16715,N_16686);
and U16802 (N_16802,N_16506,N_16586);
and U16803 (N_16803,N_16749,N_16683);
nor U16804 (N_16804,N_16720,N_16718);
and U16805 (N_16805,N_16725,N_16703);
nand U16806 (N_16806,N_16626,N_16694);
nor U16807 (N_16807,N_16545,N_16745);
nand U16808 (N_16808,N_16526,N_16551);
and U16809 (N_16809,N_16651,N_16642);
nor U16810 (N_16810,N_16550,N_16507);
nand U16811 (N_16811,N_16747,N_16585);
and U16812 (N_16812,N_16661,N_16653);
or U16813 (N_16813,N_16692,N_16654);
nand U16814 (N_16814,N_16560,N_16607);
or U16815 (N_16815,N_16652,N_16721);
nand U16816 (N_16816,N_16666,N_16598);
or U16817 (N_16817,N_16705,N_16697);
or U16818 (N_16818,N_16563,N_16676);
or U16819 (N_16819,N_16576,N_16589);
nor U16820 (N_16820,N_16644,N_16553);
and U16821 (N_16821,N_16687,N_16555);
nand U16822 (N_16822,N_16541,N_16571);
nand U16823 (N_16823,N_16520,N_16670);
nand U16824 (N_16824,N_16527,N_16699);
nand U16825 (N_16825,N_16538,N_16612);
nand U16826 (N_16826,N_16548,N_16645);
or U16827 (N_16827,N_16632,N_16614);
nor U16828 (N_16828,N_16712,N_16667);
nand U16829 (N_16829,N_16554,N_16570);
and U16830 (N_16830,N_16723,N_16568);
nor U16831 (N_16831,N_16746,N_16574);
nand U16832 (N_16832,N_16665,N_16643);
or U16833 (N_16833,N_16602,N_16698);
and U16834 (N_16834,N_16650,N_16701);
or U16835 (N_16835,N_16719,N_16605);
or U16836 (N_16836,N_16609,N_16509);
or U16837 (N_16837,N_16649,N_16518);
or U16838 (N_16838,N_16639,N_16711);
nor U16839 (N_16839,N_16580,N_16740);
and U16840 (N_16840,N_16529,N_16729);
and U16841 (N_16841,N_16593,N_16641);
nand U16842 (N_16842,N_16733,N_16628);
or U16843 (N_16843,N_16722,N_16519);
nand U16844 (N_16844,N_16736,N_16537);
nor U16845 (N_16845,N_16530,N_16748);
nor U16846 (N_16846,N_16689,N_16610);
nand U16847 (N_16847,N_16594,N_16658);
or U16848 (N_16848,N_16681,N_16521);
or U16849 (N_16849,N_16621,N_16700);
nor U16850 (N_16850,N_16546,N_16531);
nand U16851 (N_16851,N_16515,N_16501);
nand U16852 (N_16852,N_16638,N_16502);
and U16853 (N_16853,N_16708,N_16679);
and U16854 (N_16854,N_16532,N_16567);
or U16855 (N_16855,N_16508,N_16660);
nor U16856 (N_16856,N_16516,N_16706);
nor U16857 (N_16857,N_16730,N_16669);
and U16858 (N_16858,N_16533,N_16539);
and U16859 (N_16859,N_16741,N_16517);
nor U16860 (N_16860,N_16611,N_16556);
or U16861 (N_16861,N_16717,N_16534);
or U16862 (N_16862,N_16685,N_16514);
nor U16863 (N_16863,N_16672,N_16601);
and U16864 (N_16864,N_16668,N_16714);
and U16865 (N_16865,N_16622,N_16513);
and U16866 (N_16866,N_16528,N_16630);
nor U16867 (N_16867,N_16684,N_16608);
and U16868 (N_16868,N_16572,N_16583);
and U16869 (N_16869,N_16624,N_16631);
and U16870 (N_16870,N_16603,N_16613);
or U16871 (N_16871,N_16552,N_16587);
or U16872 (N_16872,N_16732,N_16581);
nor U16873 (N_16873,N_16559,N_16582);
or U16874 (N_16874,N_16561,N_16625);
and U16875 (N_16875,N_16635,N_16717);
nor U16876 (N_16876,N_16716,N_16522);
or U16877 (N_16877,N_16510,N_16533);
nand U16878 (N_16878,N_16597,N_16672);
or U16879 (N_16879,N_16536,N_16659);
or U16880 (N_16880,N_16720,N_16604);
or U16881 (N_16881,N_16720,N_16539);
nand U16882 (N_16882,N_16533,N_16528);
and U16883 (N_16883,N_16639,N_16726);
or U16884 (N_16884,N_16706,N_16742);
nor U16885 (N_16885,N_16589,N_16582);
nor U16886 (N_16886,N_16733,N_16549);
nand U16887 (N_16887,N_16508,N_16737);
nor U16888 (N_16888,N_16559,N_16558);
and U16889 (N_16889,N_16561,N_16551);
nor U16890 (N_16890,N_16523,N_16694);
nor U16891 (N_16891,N_16641,N_16678);
and U16892 (N_16892,N_16735,N_16556);
nor U16893 (N_16893,N_16664,N_16572);
nor U16894 (N_16894,N_16585,N_16654);
nor U16895 (N_16895,N_16570,N_16640);
or U16896 (N_16896,N_16647,N_16663);
and U16897 (N_16897,N_16696,N_16579);
nand U16898 (N_16898,N_16744,N_16502);
nor U16899 (N_16899,N_16565,N_16610);
nor U16900 (N_16900,N_16564,N_16681);
or U16901 (N_16901,N_16688,N_16503);
and U16902 (N_16902,N_16572,N_16609);
or U16903 (N_16903,N_16570,N_16622);
or U16904 (N_16904,N_16606,N_16608);
nand U16905 (N_16905,N_16603,N_16611);
nand U16906 (N_16906,N_16560,N_16660);
or U16907 (N_16907,N_16667,N_16703);
nor U16908 (N_16908,N_16568,N_16521);
nand U16909 (N_16909,N_16686,N_16698);
nor U16910 (N_16910,N_16682,N_16640);
or U16911 (N_16911,N_16530,N_16608);
nand U16912 (N_16912,N_16716,N_16502);
nor U16913 (N_16913,N_16550,N_16627);
nor U16914 (N_16914,N_16518,N_16718);
and U16915 (N_16915,N_16679,N_16565);
and U16916 (N_16916,N_16563,N_16516);
nor U16917 (N_16917,N_16702,N_16640);
nor U16918 (N_16918,N_16745,N_16657);
or U16919 (N_16919,N_16625,N_16667);
or U16920 (N_16920,N_16629,N_16562);
nor U16921 (N_16921,N_16645,N_16631);
xor U16922 (N_16922,N_16706,N_16586);
or U16923 (N_16923,N_16621,N_16696);
or U16924 (N_16924,N_16607,N_16519);
or U16925 (N_16925,N_16541,N_16733);
nand U16926 (N_16926,N_16747,N_16665);
nand U16927 (N_16927,N_16555,N_16707);
nand U16928 (N_16928,N_16505,N_16570);
and U16929 (N_16929,N_16617,N_16525);
nand U16930 (N_16930,N_16650,N_16520);
nand U16931 (N_16931,N_16678,N_16633);
nor U16932 (N_16932,N_16549,N_16740);
xor U16933 (N_16933,N_16607,N_16532);
and U16934 (N_16934,N_16746,N_16534);
and U16935 (N_16935,N_16730,N_16531);
nand U16936 (N_16936,N_16725,N_16564);
nor U16937 (N_16937,N_16662,N_16578);
nand U16938 (N_16938,N_16726,N_16538);
nand U16939 (N_16939,N_16675,N_16645);
nor U16940 (N_16940,N_16594,N_16532);
or U16941 (N_16941,N_16713,N_16613);
or U16942 (N_16942,N_16706,N_16669);
nand U16943 (N_16943,N_16594,N_16564);
xor U16944 (N_16944,N_16696,N_16663);
nor U16945 (N_16945,N_16671,N_16639);
or U16946 (N_16946,N_16631,N_16542);
and U16947 (N_16947,N_16566,N_16685);
or U16948 (N_16948,N_16601,N_16545);
and U16949 (N_16949,N_16664,N_16722);
nand U16950 (N_16950,N_16736,N_16552);
nor U16951 (N_16951,N_16684,N_16618);
nor U16952 (N_16952,N_16522,N_16564);
nor U16953 (N_16953,N_16718,N_16514);
nor U16954 (N_16954,N_16626,N_16622);
and U16955 (N_16955,N_16511,N_16593);
nor U16956 (N_16956,N_16682,N_16747);
nand U16957 (N_16957,N_16567,N_16563);
and U16958 (N_16958,N_16740,N_16675);
or U16959 (N_16959,N_16555,N_16510);
or U16960 (N_16960,N_16515,N_16709);
or U16961 (N_16961,N_16698,N_16661);
and U16962 (N_16962,N_16530,N_16516);
nand U16963 (N_16963,N_16729,N_16672);
or U16964 (N_16964,N_16739,N_16556);
or U16965 (N_16965,N_16630,N_16522);
nand U16966 (N_16966,N_16514,N_16731);
nor U16967 (N_16967,N_16726,N_16586);
and U16968 (N_16968,N_16680,N_16710);
or U16969 (N_16969,N_16567,N_16611);
and U16970 (N_16970,N_16714,N_16525);
and U16971 (N_16971,N_16711,N_16624);
and U16972 (N_16972,N_16679,N_16587);
nor U16973 (N_16973,N_16525,N_16580);
and U16974 (N_16974,N_16731,N_16675);
and U16975 (N_16975,N_16634,N_16622);
nand U16976 (N_16976,N_16628,N_16676);
and U16977 (N_16977,N_16715,N_16664);
and U16978 (N_16978,N_16560,N_16624);
and U16979 (N_16979,N_16737,N_16721);
nand U16980 (N_16980,N_16628,N_16746);
nor U16981 (N_16981,N_16743,N_16745);
nand U16982 (N_16982,N_16509,N_16526);
and U16983 (N_16983,N_16582,N_16526);
nand U16984 (N_16984,N_16609,N_16623);
or U16985 (N_16985,N_16692,N_16741);
or U16986 (N_16986,N_16746,N_16632);
xor U16987 (N_16987,N_16504,N_16575);
or U16988 (N_16988,N_16673,N_16514);
nand U16989 (N_16989,N_16657,N_16664);
and U16990 (N_16990,N_16598,N_16602);
nand U16991 (N_16991,N_16549,N_16524);
nand U16992 (N_16992,N_16720,N_16730);
and U16993 (N_16993,N_16671,N_16733);
nor U16994 (N_16994,N_16688,N_16599);
nor U16995 (N_16995,N_16741,N_16524);
or U16996 (N_16996,N_16638,N_16690);
nor U16997 (N_16997,N_16533,N_16523);
nor U16998 (N_16998,N_16709,N_16632);
nand U16999 (N_16999,N_16573,N_16672);
or U17000 (N_17000,N_16863,N_16753);
nand U17001 (N_17001,N_16781,N_16893);
nand U17002 (N_17002,N_16920,N_16898);
nand U17003 (N_17003,N_16813,N_16976);
nand U17004 (N_17004,N_16862,N_16832);
or U17005 (N_17005,N_16861,N_16992);
nand U17006 (N_17006,N_16933,N_16883);
or U17007 (N_17007,N_16908,N_16944);
and U17008 (N_17008,N_16957,N_16991);
nor U17009 (N_17009,N_16972,N_16897);
and U17010 (N_17010,N_16939,N_16970);
or U17011 (N_17011,N_16826,N_16942);
nand U17012 (N_17012,N_16765,N_16916);
nand U17013 (N_17013,N_16874,N_16837);
or U17014 (N_17014,N_16949,N_16987);
nand U17015 (N_17015,N_16922,N_16932);
nand U17016 (N_17016,N_16806,N_16946);
nand U17017 (N_17017,N_16770,N_16919);
or U17018 (N_17018,N_16845,N_16959);
nand U17019 (N_17019,N_16854,N_16857);
nand U17020 (N_17020,N_16924,N_16860);
nand U17021 (N_17021,N_16888,N_16761);
or U17022 (N_17022,N_16941,N_16938);
nand U17023 (N_17023,N_16958,N_16852);
or U17024 (N_17024,N_16925,N_16929);
or U17025 (N_17025,N_16973,N_16772);
nor U17026 (N_17026,N_16954,N_16935);
nor U17027 (N_17027,N_16780,N_16760);
nor U17028 (N_17028,N_16870,N_16759);
or U17029 (N_17029,N_16989,N_16782);
or U17030 (N_17030,N_16799,N_16814);
or U17031 (N_17031,N_16762,N_16768);
or U17032 (N_17032,N_16786,N_16867);
and U17033 (N_17033,N_16827,N_16803);
nand U17034 (N_17034,N_16856,N_16966);
nor U17035 (N_17035,N_16890,N_16902);
nand U17036 (N_17036,N_16978,N_16828);
or U17037 (N_17037,N_16912,N_16968);
or U17038 (N_17038,N_16937,N_16879);
or U17039 (N_17039,N_16891,N_16940);
and U17040 (N_17040,N_16997,N_16994);
or U17041 (N_17041,N_16817,N_16905);
nand U17042 (N_17042,N_16953,N_16836);
and U17043 (N_17043,N_16947,N_16766);
nand U17044 (N_17044,N_16843,N_16907);
or U17045 (N_17045,N_16797,N_16808);
or U17046 (N_17046,N_16903,N_16921);
or U17047 (N_17047,N_16774,N_16985);
nor U17048 (N_17048,N_16988,N_16869);
and U17049 (N_17049,N_16993,N_16951);
nor U17050 (N_17050,N_16792,N_16775);
nor U17051 (N_17051,N_16923,N_16784);
or U17052 (N_17052,N_16796,N_16871);
nor U17053 (N_17053,N_16811,N_16794);
and U17054 (N_17054,N_16915,N_16795);
nor U17055 (N_17055,N_16977,N_16804);
nor U17056 (N_17056,N_16850,N_16855);
and U17057 (N_17057,N_16763,N_16886);
or U17058 (N_17058,N_16969,N_16787);
and U17059 (N_17059,N_16788,N_16834);
or U17060 (N_17060,N_16980,N_16877);
or U17061 (N_17061,N_16841,N_16918);
xor U17062 (N_17062,N_16764,N_16962);
and U17063 (N_17063,N_16830,N_16881);
nor U17064 (N_17064,N_16805,N_16816);
nand U17065 (N_17065,N_16838,N_16777);
nor U17066 (N_17066,N_16892,N_16823);
and U17067 (N_17067,N_16931,N_16757);
nand U17068 (N_17068,N_16943,N_16767);
and U17069 (N_17069,N_16906,N_16866);
or U17070 (N_17070,N_16983,N_16773);
and U17071 (N_17071,N_16831,N_16900);
or U17072 (N_17072,N_16961,N_16865);
and U17073 (N_17073,N_16776,N_16779);
or U17074 (N_17074,N_16926,N_16960);
nor U17075 (N_17075,N_16955,N_16878);
or U17076 (N_17076,N_16801,N_16825);
nor U17077 (N_17077,N_16755,N_16842);
nor U17078 (N_17078,N_16996,N_16858);
and U17079 (N_17079,N_16818,N_16810);
nand U17080 (N_17080,N_16887,N_16839);
nor U17081 (N_17081,N_16821,N_16868);
or U17082 (N_17082,N_16778,N_16798);
and U17083 (N_17083,N_16844,N_16956);
nor U17084 (N_17084,N_16975,N_16802);
or U17085 (N_17085,N_16945,N_16896);
nor U17086 (N_17086,N_16927,N_16979);
nand U17087 (N_17087,N_16952,N_16791);
or U17088 (N_17088,N_16930,N_16771);
or U17089 (N_17089,N_16769,N_16965);
and U17090 (N_17090,N_16750,N_16833);
and U17091 (N_17091,N_16789,N_16934);
and U17092 (N_17092,N_16793,N_16872);
nand U17093 (N_17093,N_16849,N_16884);
nor U17094 (N_17094,N_16785,N_16964);
nand U17095 (N_17095,N_16812,N_16851);
or U17096 (N_17096,N_16809,N_16936);
and U17097 (N_17097,N_16752,N_16822);
nor U17098 (N_17098,N_16901,N_16974);
or U17099 (N_17099,N_16853,N_16971);
nor U17100 (N_17100,N_16998,N_16894);
and U17101 (N_17101,N_16914,N_16899);
and U17102 (N_17102,N_16756,N_16783);
nand U17103 (N_17103,N_16859,N_16895);
or U17104 (N_17104,N_16950,N_16758);
nor U17105 (N_17105,N_16751,N_16882);
nand U17106 (N_17106,N_16981,N_16848);
and U17107 (N_17107,N_16819,N_16790);
or U17108 (N_17108,N_16889,N_16846);
nor U17109 (N_17109,N_16986,N_16995);
nand U17110 (N_17110,N_16873,N_16829);
nor U17111 (N_17111,N_16815,N_16820);
xor U17112 (N_17112,N_16913,N_16967);
nor U17113 (N_17113,N_16885,N_16875);
and U17114 (N_17114,N_16835,N_16963);
nand U17115 (N_17115,N_16876,N_16990);
and U17116 (N_17116,N_16917,N_16864);
or U17117 (N_17117,N_16904,N_16824);
nor U17118 (N_17118,N_16910,N_16800);
and U17119 (N_17119,N_16847,N_16948);
or U17120 (N_17120,N_16909,N_16840);
and U17121 (N_17121,N_16880,N_16982);
nor U17122 (N_17122,N_16984,N_16807);
and U17123 (N_17123,N_16999,N_16754);
nor U17124 (N_17124,N_16928,N_16911);
nand U17125 (N_17125,N_16804,N_16814);
nor U17126 (N_17126,N_16855,N_16780);
or U17127 (N_17127,N_16808,N_16771);
xnor U17128 (N_17128,N_16981,N_16911);
nand U17129 (N_17129,N_16938,N_16846);
or U17130 (N_17130,N_16904,N_16870);
nor U17131 (N_17131,N_16863,N_16875);
and U17132 (N_17132,N_16991,N_16992);
and U17133 (N_17133,N_16761,N_16982);
nand U17134 (N_17134,N_16888,N_16829);
nor U17135 (N_17135,N_16763,N_16927);
nand U17136 (N_17136,N_16963,N_16883);
or U17137 (N_17137,N_16955,N_16755);
and U17138 (N_17138,N_16938,N_16928);
nor U17139 (N_17139,N_16930,N_16880);
nor U17140 (N_17140,N_16807,N_16938);
nand U17141 (N_17141,N_16942,N_16992);
or U17142 (N_17142,N_16931,N_16942);
and U17143 (N_17143,N_16926,N_16794);
nand U17144 (N_17144,N_16927,N_16793);
nor U17145 (N_17145,N_16925,N_16924);
and U17146 (N_17146,N_16760,N_16931);
nor U17147 (N_17147,N_16882,N_16915);
nand U17148 (N_17148,N_16778,N_16824);
nand U17149 (N_17149,N_16758,N_16949);
and U17150 (N_17150,N_16754,N_16822);
or U17151 (N_17151,N_16894,N_16828);
or U17152 (N_17152,N_16817,N_16819);
nor U17153 (N_17153,N_16804,N_16951);
nand U17154 (N_17154,N_16901,N_16886);
and U17155 (N_17155,N_16973,N_16841);
nor U17156 (N_17156,N_16999,N_16829);
or U17157 (N_17157,N_16756,N_16944);
nand U17158 (N_17158,N_16807,N_16829);
nor U17159 (N_17159,N_16840,N_16854);
or U17160 (N_17160,N_16876,N_16793);
and U17161 (N_17161,N_16834,N_16862);
and U17162 (N_17162,N_16897,N_16756);
nor U17163 (N_17163,N_16906,N_16831);
nor U17164 (N_17164,N_16791,N_16753);
or U17165 (N_17165,N_16931,N_16970);
nor U17166 (N_17166,N_16786,N_16989);
nand U17167 (N_17167,N_16835,N_16822);
nor U17168 (N_17168,N_16879,N_16841);
nand U17169 (N_17169,N_16878,N_16991);
nand U17170 (N_17170,N_16870,N_16763);
nor U17171 (N_17171,N_16883,N_16869);
xor U17172 (N_17172,N_16965,N_16941);
nand U17173 (N_17173,N_16907,N_16882);
nand U17174 (N_17174,N_16903,N_16994);
or U17175 (N_17175,N_16840,N_16790);
nor U17176 (N_17176,N_16938,N_16756);
nand U17177 (N_17177,N_16971,N_16877);
or U17178 (N_17178,N_16849,N_16883);
or U17179 (N_17179,N_16967,N_16903);
and U17180 (N_17180,N_16970,N_16875);
nor U17181 (N_17181,N_16970,N_16880);
xor U17182 (N_17182,N_16919,N_16833);
and U17183 (N_17183,N_16948,N_16762);
nor U17184 (N_17184,N_16986,N_16829);
nor U17185 (N_17185,N_16947,N_16883);
nor U17186 (N_17186,N_16953,N_16900);
nand U17187 (N_17187,N_16905,N_16763);
nor U17188 (N_17188,N_16781,N_16810);
nand U17189 (N_17189,N_16917,N_16938);
nor U17190 (N_17190,N_16876,N_16808);
and U17191 (N_17191,N_16947,N_16782);
nand U17192 (N_17192,N_16966,N_16822);
nor U17193 (N_17193,N_16893,N_16902);
and U17194 (N_17194,N_16928,N_16808);
or U17195 (N_17195,N_16809,N_16993);
nand U17196 (N_17196,N_16967,N_16897);
or U17197 (N_17197,N_16785,N_16997);
nand U17198 (N_17198,N_16774,N_16809);
and U17199 (N_17199,N_16845,N_16756);
and U17200 (N_17200,N_16754,N_16824);
or U17201 (N_17201,N_16898,N_16783);
nor U17202 (N_17202,N_16941,N_16961);
nor U17203 (N_17203,N_16796,N_16754);
nand U17204 (N_17204,N_16968,N_16819);
nand U17205 (N_17205,N_16779,N_16853);
or U17206 (N_17206,N_16870,N_16857);
or U17207 (N_17207,N_16812,N_16960);
nor U17208 (N_17208,N_16846,N_16810);
nor U17209 (N_17209,N_16824,N_16781);
nor U17210 (N_17210,N_16862,N_16854);
and U17211 (N_17211,N_16878,N_16826);
or U17212 (N_17212,N_16884,N_16883);
or U17213 (N_17213,N_16811,N_16901);
and U17214 (N_17214,N_16852,N_16924);
and U17215 (N_17215,N_16808,N_16892);
or U17216 (N_17216,N_16982,N_16910);
and U17217 (N_17217,N_16982,N_16752);
or U17218 (N_17218,N_16820,N_16960);
nor U17219 (N_17219,N_16795,N_16868);
or U17220 (N_17220,N_16899,N_16955);
and U17221 (N_17221,N_16784,N_16922);
nor U17222 (N_17222,N_16914,N_16757);
nand U17223 (N_17223,N_16836,N_16944);
or U17224 (N_17224,N_16989,N_16820);
and U17225 (N_17225,N_16858,N_16755);
or U17226 (N_17226,N_16844,N_16873);
and U17227 (N_17227,N_16802,N_16833);
or U17228 (N_17228,N_16981,N_16798);
nor U17229 (N_17229,N_16817,N_16868);
nand U17230 (N_17230,N_16992,N_16837);
nor U17231 (N_17231,N_16864,N_16942);
or U17232 (N_17232,N_16814,N_16850);
nor U17233 (N_17233,N_16858,N_16910);
nand U17234 (N_17234,N_16839,N_16993);
or U17235 (N_17235,N_16818,N_16813);
nand U17236 (N_17236,N_16893,N_16833);
and U17237 (N_17237,N_16999,N_16980);
nor U17238 (N_17238,N_16942,N_16796);
nand U17239 (N_17239,N_16958,N_16879);
or U17240 (N_17240,N_16980,N_16928);
nor U17241 (N_17241,N_16809,N_16951);
nor U17242 (N_17242,N_16845,N_16996);
nand U17243 (N_17243,N_16940,N_16794);
nor U17244 (N_17244,N_16821,N_16870);
nand U17245 (N_17245,N_16755,N_16904);
or U17246 (N_17246,N_16934,N_16970);
or U17247 (N_17247,N_16760,N_16762);
and U17248 (N_17248,N_16761,N_16834);
nor U17249 (N_17249,N_16973,N_16797);
and U17250 (N_17250,N_17054,N_17123);
and U17251 (N_17251,N_17209,N_17215);
xor U17252 (N_17252,N_17078,N_17226);
or U17253 (N_17253,N_17018,N_17122);
nand U17254 (N_17254,N_17156,N_17224);
nand U17255 (N_17255,N_17165,N_17099);
nand U17256 (N_17256,N_17004,N_17195);
or U17257 (N_17257,N_17241,N_17221);
nand U17258 (N_17258,N_17100,N_17025);
nor U17259 (N_17259,N_17112,N_17184);
nand U17260 (N_17260,N_17111,N_17017);
nor U17261 (N_17261,N_17177,N_17074);
or U17262 (N_17262,N_17031,N_17124);
nand U17263 (N_17263,N_17013,N_17058);
or U17264 (N_17264,N_17213,N_17023);
nor U17265 (N_17265,N_17164,N_17007);
or U17266 (N_17266,N_17069,N_17231);
or U17267 (N_17267,N_17180,N_17237);
nand U17268 (N_17268,N_17079,N_17240);
or U17269 (N_17269,N_17137,N_17169);
or U17270 (N_17270,N_17066,N_17245);
or U17271 (N_17271,N_17027,N_17068);
or U17272 (N_17272,N_17026,N_17201);
nor U17273 (N_17273,N_17159,N_17009);
or U17274 (N_17274,N_17202,N_17194);
nand U17275 (N_17275,N_17121,N_17060);
or U17276 (N_17276,N_17236,N_17085);
nor U17277 (N_17277,N_17091,N_17010);
or U17278 (N_17278,N_17171,N_17002);
and U17279 (N_17279,N_17126,N_17132);
nand U17280 (N_17280,N_17063,N_17077);
or U17281 (N_17281,N_17097,N_17062);
nand U17282 (N_17282,N_17189,N_17248);
and U17283 (N_17283,N_17044,N_17016);
nor U17284 (N_17284,N_17092,N_17153);
or U17285 (N_17285,N_17155,N_17046);
or U17286 (N_17286,N_17141,N_17030);
nor U17287 (N_17287,N_17244,N_17093);
nor U17288 (N_17288,N_17197,N_17140);
or U17289 (N_17289,N_17117,N_17131);
and U17290 (N_17290,N_17029,N_17076);
and U17291 (N_17291,N_17130,N_17113);
nor U17292 (N_17292,N_17035,N_17109);
and U17293 (N_17293,N_17219,N_17056);
nand U17294 (N_17294,N_17229,N_17191);
nand U17295 (N_17295,N_17014,N_17214);
and U17296 (N_17296,N_17083,N_17116);
nand U17297 (N_17297,N_17034,N_17175);
and U17298 (N_17298,N_17082,N_17086);
nor U17299 (N_17299,N_17089,N_17235);
nand U17300 (N_17300,N_17115,N_17243);
nor U17301 (N_17301,N_17228,N_17182);
and U17302 (N_17302,N_17151,N_17238);
nor U17303 (N_17303,N_17040,N_17098);
and U17304 (N_17304,N_17166,N_17206);
nand U17305 (N_17305,N_17188,N_17216);
and U17306 (N_17306,N_17059,N_17106);
nand U17307 (N_17307,N_17144,N_17105);
nand U17308 (N_17308,N_17170,N_17203);
nand U17309 (N_17309,N_17249,N_17028);
or U17310 (N_17310,N_17208,N_17102);
xor U17311 (N_17311,N_17168,N_17220);
nor U17312 (N_17312,N_17185,N_17139);
nor U17313 (N_17313,N_17176,N_17071);
nand U17314 (N_17314,N_17133,N_17227);
and U17315 (N_17315,N_17101,N_17087);
nor U17316 (N_17316,N_17125,N_17043);
nor U17317 (N_17317,N_17088,N_17006);
or U17318 (N_17318,N_17193,N_17104);
nor U17319 (N_17319,N_17190,N_17142);
and U17320 (N_17320,N_17246,N_17212);
and U17321 (N_17321,N_17084,N_17048);
and U17322 (N_17322,N_17003,N_17128);
or U17323 (N_17323,N_17008,N_17036);
nand U17324 (N_17324,N_17021,N_17108);
nor U17325 (N_17325,N_17095,N_17136);
and U17326 (N_17326,N_17234,N_17223);
or U17327 (N_17327,N_17158,N_17075);
nand U17328 (N_17328,N_17051,N_17199);
nor U17329 (N_17329,N_17163,N_17019);
nor U17330 (N_17330,N_17129,N_17233);
nor U17331 (N_17331,N_17135,N_17055);
nand U17332 (N_17332,N_17174,N_17011);
or U17333 (N_17333,N_17012,N_17001);
or U17334 (N_17334,N_17147,N_17187);
nand U17335 (N_17335,N_17005,N_17196);
nor U17336 (N_17336,N_17067,N_17207);
nor U17337 (N_17337,N_17127,N_17038);
nor U17338 (N_17338,N_17161,N_17070);
nand U17339 (N_17339,N_17167,N_17049);
and U17340 (N_17340,N_17232,N_17081);
nand U17341 (N_17341,N_17042,N_17096);
or U17342 (N_17342,N_17178,N_17000);
nand U17343 (N_17343,N_17107,N_17211);
or U17344 (N_17344,N_17179,N_17150);
nand U17345 (N_17345,N_17103,N_17032);
and U17346 (N_17346,N_17080,N_17204);
nor U17347 (N_17347,N_17037,N_17045);
and U17348 (N_17348,N_17181,N_17218);
nor U17349 (N_17349,N_17015,N_17242);
and U17350 (N_17350,N_17053,N_17145);
or U17351 (N_17351,N_17198,N_17065);
or U17352 (N_17352,N_17192,N_17222);
nor U17353 (N_17353,N_17064,N_17173);
or U17354 (N_17354,N_17118,N_17039);
and U17355 (N_17355,N_17057,N_17183);
nand U17356 (N_17356,N_17210,N_17033);
or U17357 (N_17357,N_17114,N_17172);
or U17358 (N_17358,N_17072,N_17146);
nand U17359 (N_17359,N_17138,N_17247);
or U17360 (N_17360,N_17050,N_17022);
and U17361 (N_17361,N_17225,N_17061);
nand U17362 (N_17362,N_17217,N_17073);
nand U17363 (N_17363,N_17160,N_17047);
xnor U17364 (N_17364,N_17143,N_17119);
nor U17365 (N_17365,N_17024,N_17149);
or U17366 (N_17366,N_17154,N_17157);
and U17367 (N_17367,N_17052,N_17162);
and U17368 (N_17368,N_17134,N_17148);
or U17369 (N_17369,N_17020,N_17200);
nand U17370 (N_17370,N_17205,N_17041);
and U17371 (N_17371,N_17120,N_17230);
xor U17372 (N_17372,N_17094,N_17152);
and U17373 (N_17373,N_17110,N_17239);
nand U17374 (N_17374,N_17090,N_17186);
nor U17375 (N_17375,N_17140,N_17206);
nand U17376 (N_17376,N_17223,N_17086);
nor U17377 (N_17377,N_17164,N_17128);
or U17378 (N_17378,N_17170,N_17204);
or U17379 (N_17379,N_17102,N_17213);
and U17380 (N_17380,N_17182,N_17152);
nand U17381 (N_17381,N_17047,N_17244);
nor U17382 (N_17382,N_17025,N_17179);
or U17383 (N_17383,N_17142,N_17235);
or U17384 (N_17384,N_17013,N_17008);
or U17385 (N_17385,N_17215,N_17152);
or U17386 (N_17386,N_17086,N_17088);
nand U17387 (N_17387,N_17004,N_17196);
or U17388 (N_17388,N_17148,N_17204);
nor U17389 (N_17389,N_17132,N_17232);
nand U17390 (N_17390,N_17150,N_17094);
nand U17391 (N_17391,N_17209,N_17231);
nand U17392 (N_17392,N_17247,N_17199);
or U17393 (N_17393,N_17119,N_17043);
nor U17394 (N_17394,N_17028,N_17045);
or U17395 (N_17395,N_17220,N_17166);
nand U17396 (N_17396,N_17112,N_17088);
and U17397 (N_17397,N_17207,N_17127);
nor U17398 (N_17398,N_17099,N_17061);
or U17399 (N_17399,N_17236,N_17024);
or U17400 (N_17400,N_17009,N_17086);
and U17401 (N_17401,N_17142,N_17157);
or U17402 (N_17402,N_17180,N_17225);
nand U17403 (N_17403,N_17230,N_17172);
and U17404 (N_17404,N_17129,N_17133);
nor U17405 (N_17405,N_17184,N_17132);
nand U17406 (N_17406,N_17072,N_17012);
or U17407 (N_17407,N_17016,N_17058);
or U17408 (N_17408,N_17170,N_17118);
nand U17409 (N_17409,N_17198,N_17157);
nand U17410 (N_17410,N_17078,N_17029);
or U17411 (N_17411,N_17156,N_17171);
nor U17412 (N_17412,N_17033,N_17061);
nand U17413 (N_17413,N_17080,N_17167);
nor U17414 (N_17414,N_17185,N_17199);
and U17415 (N_17415,N_17190,N_17028);
nor U17416 (N_17416,N_17008,N_17144);
nand U17417 (N_17417,N_17156,N_17020);
nor U17418 (N_17418,N_17075,N_17081);
nand U17419 (N_17419,N_17091,N_17006);
nor U17420 (N_17420,N_17066,N_17232);
and U17421 (N_17421,N_17073,N_17064);
or U17422 (N_17422,N_17201,N_17179);
nor U17423 (N_17423,N_17103,N_17238);
nand U17424 (N_17424,N_17183,N_17215);
nand U17425 (N_17425,N_17183,N_17156);
nor U17426 (N_17426,N_17121,N_17072);
and U17427 (N_17427,N_17008,N_17137);
or U17428 (N_17428,N_17096,N_17053);
or U17429 (N_17429,N_17094,N_17182);
and U17430 (N_17430,N_17203,N_17035);
and U17431 (N_17431,N_17075,N_17230);
or U17432 (N_17432,N_17081,N_17003);
nor U17433 (N_17433,N_17136,N_17063);
nor U17434 (N_17434,N_17024,N_17084);
nand U17435 (N_17435,N_17172,N_17166);
or U17436 (N_17436,N_17073,N_17238);
nor U17437 (N_17437,N_17012,N_17165);
nand U17438 (N_17438,N_17143,N_17173);
nand U17439 (N_17439,N_17138,N_17197);
and U17440 (N_17440,N_17002,N_17113);
nor U17441 (N_17441,N_17207,N_17154);
nor U17442 (N_17442,N_17009,N_17174);
and U17443 (N_17443,N_17057,N_17120);
nand U17444 (N_17444,N_17045,N_17042);
and U17445 (N_17445,N_17085,N_17152);
nor U17446 (N_17446,N_17071,N_17243);
or U17447 (N_17447,N_17191,N_17216);
or U17448 (N_17448,N_17074,N_17239);
nor U17449 (N_17449,N_17112,N_17191);
nand U17450 (N_17450,N_17133,N_17184);
nor U17451 (N_17451,N_17239,N_17246);
nand U17452 (N_17452,N_17204,N_17056);
nand U17453 (N_17453,N_17026,N_17180);
or U17454 (N_17454,N_17034,N_17244);
xnor U17455 (N_17455,N_17213,N_17179);
nor U17456 (N_17456,N_17114,N_17185);
nand U17457 (N_17457,N_17003,N_17069);
and U17458 (N_17458,N_17115,N_17055);
nand U17459 (N_17459,N_17240,N_17243);
nand U17460 (N_17460,N_17170,N_17187);
or U17461 (N_17461,N_17238,N_17236);
nor U17462 (N_17462,N_17026,N_17110);
nor U17463 (N_17463,N_17174,N_17034);
nand U17464 (N_17464,N_17127,N_17031);
nor U17465 (N_17465,N_17065,N_17144);
and U17466 (N_17466,N_17036,N_17147);
xnor U17467 (N_17467,N_17187,N_17117);
nand U17468 (N_17468,N_17214,N_17192);
and U17469 (N_17469,N_17208,N_17221);
and U17470 (N_17470,N_17070,N_17038);
nand U17471 (N_17471,N_17236,N_17122);
nand U17472 (N_17472,N_17025,N_17018);
and U17473 (N_17473,N_17115,N_17155);
and U17474 (N_17474,N_17150,N_17067);
or U17475 (N_17475,N_17122,N_17098);
or U17476 (N_17476,N_17233,N_17206);
or U17477 (N_17477,N_17229,N_17091);
and U17478 (N_17478,N_17128,N_17113);
nor U17479 (N_17479,N_17042,N_17181);
and U17480 (N_17480,N_17140,N_17042);
nor U17481 (N_17481,N_17099,N_17038);
and U17482 (N_17482,N_17027,N_17004);
and U17483 (N_17483,N_17008,N_17071);
or U17484 (N_17484,N_17230,N_17198);
nand U17485 (N_17485,N_17093,N_17064);
nand U17486 (N_17486,N_17074,N_17200);
or U17487 (N_17487,N_17153,N_17169);
nor U17488 (N_17488,N_17152,N_17055);
or U17489 (N_17489,N_17126,N_17216);
nand U17490 (N_17490,N_17200,N_17214);
and U17491 (N_17491,N_17199,N_17049);
nand U17492 (N_17492,N_17068,N_17203);
nand U17493 (N_17493,N_17175,N_17134);
nand U17494 (N_17494,N_17181,N_17073);
nor U17495 (N_17495,N_17081,N_17098);
and U17496 (N_17496,N_17040,N_17016);
nor U17497 (N_17497,N_17174,N_17242);
nand U17498 (N_17498,N_17058,N_17208);
or U17499 (N_17499,N_17126,N_17154);
nand U17500 (N_17500,N_17361,N_17297);
nor U17501 (N_17501,N_17258,N_17444);
nor U17502 (N_17502,N_17296,N_17446);
and U17503 (N_17503,N_17450,N_17354);
or U17504 (N_17504,N_17334,N_17323);
and U17505 (N_17505,N_17307,N_17417);
nor U17506 (N_17506,N_17443,N_17329);
nor U17507 (N_17507,N_17411,N_17377);
nand U17508 (N_17508,N_17440,N_17295);
and U17509 (N_17509,N_17474,N_17403);
or U17510 (N_17510,N_17415,N_17331);
and U17511 (N_17511,N_17363,N_17448);
nand U17512 (N_17512,N_17313,N_17314);
and U17513 (N_17513,N_17370,N_17442);
and U17514 (N_17514,N_17283,N_17321);
or U17515 (N_17515,N_17461,N_17410);
and U17516 (N_17516,N_17468,N_17469);
or U17517 (N_17517,N_17421,N_17281);
and U17518 (N_17518,N_17357,N_17375);
nor U17519 (N_17519,N_17330,N_17325);
or U17520 (N_17520,N_17385,N_17301);
or U17521 (N_17521,N_17259,N_17310);
nor U17522 (N_17522,N_17378,N_17466);
nand U17523 (N_17523,N_17473,N_17482);
nor U17524 (N_17524,N_17389,N_17436);
or U17525 (N_17525,N_17472,N_17419);
or U17526 (N_17526,N_17449,N_17479);
and U17527 (N_17527,N_17272,N_17496);
nor U17528 (N_17528,N_17251,N_17464);
and U17529 (N_17529,N_17445,N_17367);
nand U17530 (N_17530,N_17453,N_17480);
xnor U17531 (N_17531,N_17342,N_17276);
nor U17532 (N_17532,N_17348,N_17260);
and U17533 (N_17533,N_17397,N_17412);
nand U17534 (N_17534,N_17339,N_17418);
and U17535 (N_17535,N_17358,N_17265);
or U17536 (N_17536,N_17499,N_17343);
or U17537 (N_17537,N_17253,N_17327);
and U17538 (N_17538,N_17484,N_17485);
nor U17539 (N_17539,N_17455,N_17393);
or U17540 (N_17540,N_17289,N_17438);
nand U17541 (N_17541,N_17381,N_17275);
or U17542 (N_17542,N_17288,N_17369);
or U17543 (N_17543,N_17332,N_17463);
nand U17544 (N_17544,N_17390,N_17405);
nand U17545 (N_17545,N_17382,N_17439);
or U17546 (N_17546,N_17372,N_17497);
nand U17547 (N_17547,N_17300,N_17432);
nand U17548 (N_17548,N_17498,N_17399);
nand U17549 (N_17549,N_17284,N_17293);
or U17550 (N_17550,N_17366,N_17317);
or U17551 (N_17551,N_17287,N_17319);
and U17552 (N_17552,N_17355,N_17413);
and U17553 (N_17553,N_17488,N_17353);
nor U17554 (N_17554,N_17487,N_17430);
or U17555 (N_17555,N_17494,N_17359);
nand U17556 (N_17556,N_17458,N_17368);
nor U17557 (N_17557,N_17280,N_17262);
nand U17558 (N_17558,N_17392,N_17282);
nor U17559 (N_17559,N_17263,N_17414);
nand U17560 (N_17560,N_17404,N_17407);
nand U17561 (N_17561,N_17252,N_17447);
and U17562 (N_17562,N_17303,N_17335);
nand U17563 (N_17563,N_17470,N_17338);
or U17564 (N_17564,N_17386,N_17427);
xnor U17565 (N_17565,N_17315,N_17416);
or U17566 (N_17566,N_17264,N_17356);
nor U17567 (N_17567,N_17268,N_17424);
nand U17568 (N_17568,N_17478,N_17437);
nor U17569 (N_17569,N_17400,N_17328);
or U17570 (N_17570,N_17364,N_17391);
nand U17571 (N_17571,N_17360,N_17476);
or U17572 (N_17572,N_17341,N_17306);
or U17573 (N_17573,N_17406,N_17379);
nand U17574 (N_17574,N_17495,N_17493);
nand U17575 (N_17575,N_17285,N_17322);
nor U17576 (N_17576,N_17344,N_17333);
and U17577 (N_17577,N_17398,N_17302);
nor U17578 (N_17578,N_17336,N_17428);
and U17579 (N_17579,N_17490,N_17489);
and U17580 (N_17580,N_17324,N_17471);
and U17581 (N_17581,N_17380,N_17483);
and U17582 (N_17582,N_17435,N_17475);
nor U17583 (N_17583,N_17441,N_17434);
and U17584 (N_17584,N_17451,N_17365);
or U17585 (N_17585,N_17273,N_17349);
nor U17586 (N_17586,N_17373,N_17290);
nor U17587 (N_17587,N_17374,N_17388);
and U17588 (N_17588,N_17409,N_17340);
or U17589 (N_17589,N_17278,N_17316);
nor U17590 (N_17590,N_17477,N_17267);
or U17591 (N_17591,N_17250,N_17426);
and U17592 (N_17592,N_17255,N_17350);
nor U17593 (N_17593,N_17491,N_17429);
xor U17594 (N_17594,N_17457,N_17486);
nor U17595 (N_17595,N_17311,N_17257);
nor U17596 (N_17596,N_17371,N_17459);
nor U17597 (N_17597,N_17384,N_17320);
nand U17598 (N_17598,N_17396,N_17423);
and U17599 (N_17599,N_17376,N_17347);
or U17600 (N_17600,N_17422,N_17420);
or U17601 (N_17601,N_17452,N_17394);
and U17602 (N_17602,N_17465,N_17454);
and U17603 (N_17603,N_17462,N_17298);
and U17604 (N_17604,N_17346,N_17299);
nand U17605 (N_17605,N_17304,N_17308);
or U17606 (N_17606,N_17395,N_17362);
and U17607 (N_17607,N_17277,N_17305);
or U17608 (N_17608,N_17279,N_17312);
nor U17609 (N_17609,N_17269,N_17309);
nor U17610 (N_17610,N_17286,N_17351);
nand U17611 (N_17611,N_17274,N_17433);
and U17612 (N_17612,N_17256,N_17318);
nand U17613 (N_17613,N_17270,N_17383);
and U17614 (N_17614,N_17408,N_17456);
and U17615 (N_17615,N_17387,N_17254);
and U17616 (N_17616,N_17292,N_17401);
nor U17617 (N_17617,N_17492,N_17266);
and U17618 (N_17618,N_17352,N_17337);
nor U17619 (N_17619,N_17460,N_17467);
nor U17620 (N_17620,N_17345,N_17261);
and U17621 (N_17621,N_17294,N_17481);
and U17622 (N_17622,N_17431,N_17402);
nand U17623 (N_17623,N_17425,N_17326);
nor U17624 (N_17624,N_17291,N_17271);
and U17625 (N_17625,N_17417,N_17314);
nand U17626 (N_17626,N_17295,N_17446);
nor U17627 (N_17627,N_17461,N_17296);
or U17628 (N_17628,N_17316,N_17256);
nand U17629 (N_17629,N_17376,N_17429);
nor U17630 (N_17630,N_17474,N_17268);
nand U17631 (N_17631,N_17250,N_17466);
and U17632 (N_17632,N_17479,N_17265);
and U17633 (N_17633,N_17405,N_17456);
nand U17634 (N_17634,N_17423,N_17482);
nand U17635 (N_17635,N_17396,N_17409);
nor U17636 (N_17636,N_17253,N_17458);
or U17637 (N_17637,N_17304,N_17339);
and U17638 (N_17638,N_17257,N_17378);
nand U17639 (N_17639,N_17409,N_17270);
and U17640 (N_17640,N_17489,N_17317);
nand U17641 (N_17641,N_17251,N_17491);
and U17642 (N_17642,N_17478,N_17449);
and U17643 (N_17643,N_17439,N_17297);
nand U17644 (N_17644,N_17498,N_17490);
nand U17645 (N_17645,N_17432,N_17390);
and U17646 (N_17646,N_17401,N_17489);
and U17647 (N_17647,N_17318,N_17409);
or U17648 (N_17648,N_17295,N_17351);
and U17649 (N_17649,N_17465,N_17382);
and U17650 (N_17650,N_17481,N_17344);
nand U17651 (N_17651,N_17321,N_17386);
or U17652 (N_17652,N_17292,N_17317);
and U17653 (N_17653,N_17307,N_17339);
nor U17654 (N_17654,N_17363,N_17475);
nor U17655 (N_17655,N_17470,N_17253);
or U17656 (N_17656,N_17315,N_17440);
nor U17657 (N_17657,N_17387,N_17319);
or U17658 (N_17658,N_17473,N_17262);
nand U17659 (N_17659,N_17325,N_17380);
nor U17660 (N_17660,N_17498,N_17328);
or U17661 (N_17661,N_17286,N_17400);
nor U17662 (N_17662,N_17271,N_17452);
and U17663 (N_17663,N_17329,N_17346);
nand U17664 (N_17664,N_17304,N_17385);
nor U17665 (N_17665,N_17295,N_17252);
xnor U17666 (N_17666,N_17320,N_17366);
nand U17667 (N_17667,N_17385,N_17498);
xor U17668 (N_17668,N_17423,N_17364);
or U17669 (N_17669,N_17466,N_17343);
and U17670 (N_17670,N_17324,N_17423);
and U17671 (N_17671,N_17442,N_17452);
nor U17672 (N_17672,N_17272,N_17311);
nand U17673 (N_17673,N_17284,N_17359);
nor U17674 (N_17674,N_17313,N_17275);
nand U17675 (N_17675,N_17315,N_17265);
and U17676 (N_17676,N_17454,N_17340);
nor U17677 (N_17677,N_17369,N_17437);
and U17678 (N_17678,N_17388,N_17308);
or U17679 (N_17679,N_17410,N_17442);
nand U17680 (N_17680,N_17262,N_17444);
nor U17681 (N_17681,N_17309,N_17294);
and U17682 (N_17682,N_17325,N_17407);
nor U17683 (N_17683,N_17383,N_17435);
nor U17684 (N_17684,N_17320,N_17371);
nand U17685 (N_17685,N_17351,N_17293);
nor U17686 (N_17686,N_17464,N_17303);
and U17687 (N_17687,N_17304,N_17487);
or U17688 (N_17688,N_17453,N_17256);
and U17689 (N_17689,N_17432,N_17448);
nand U17690 (N_17690,N_17374,N_17417);
and U17691 (N_17691,N_17409,N_17401);
or U17692 (N_17692,N_17436,N_17335);
or U17693 (N_17693,N_17391,N_17354);
nand U17694 (N_17694,N_17390,N_17356);
nor U17695 (N_17695,N_17356,N_17405);
nor U17696 (N_17696,N_17402,N_17286);
or U17697 (N_17697,N_17447,N_17310);
nand U17698 (N_17698,N_17481,N_17497);
or U17699 (N_17699,N_17316,N_17339);
or U17700 (N_17700,N_17440,N_17479);
nor U17701 (N_17701,N_17435,N_17472);
and U17702 (N_17702,N_17335,N_17393);
nor U17703 (N_17703,N_17387,N_17312);
or U17704 (N_17704,N_17310,N_17353);
nor U17705 (N_17705,N_17438,N_17376);
or U17706 (N_17706,N_17336,N_17446);
or U17707 (N_17707,N_17263,N_17409);
nor U17708 (N_17708,N_17272,N_17373);
or U17709 (N_17709,N_17282,N_17498);
nor U17710 (N_17710,N_17459,N_17342);
or U17711 (N_17711,N_17314,N_17321);
nor U17712 (N_17712,N_17264,N_17475);
or U17713 (N_17713,N_17281,N_17479);
and U17714 (N_17714,N_17261,N_17272);
nand U17715 (N_17715,N_17433,N_17376);
and U17716 (N_17716,N_17488,N_17336);
nor U17717 (N_17717,N_17370,N_17381);
xor U17718 (N_17718,N_17406,N_17330);
and U17719 (N_17719,N_17484,N_17257);
or U17720 (N_17720,N_17291,N_17261);
nand U17721 (N_17721,N_17346,N_17306);
nand U17722 (N_17722,N_17430,N_17434);
or U17723 (N_17723,N_17300,N_17344);
and U17724 (N_17724,N_17463,N_17313);
and U17725 (N_17725,N_17309,N_17453);
and U17726 (N_17726,N_17276,N_17499);
and U17727 (N_17727,N_17496,N_17256);
nand U17728 (N_17728,N_17373,N_17390);
and U17729 (N_17729,N_17499,N_17398);
or U17730 (N_17730,N_17360,N_17387);
and U17731 (N_17731,N_17329,N_17316);
or U17732 (N_17732,N_17416,N_17374);
and U17733 (N_17733,N_17284,N_17344);
nor U17734 (N_17734,N_17480,N_17442);
nor U17735 (N_17735,N_17464,N_17438);
nand U17736 (N_17736,N_17266,N_17332);
nand U17737 (N_17737,N_17350,N_17319);
nor U17738 (N_17738,N_17453,N_17400);
nand U17739 (N_17739,N_17274,N_17481);
or U17740 (N_17740,N_17316,N_17412);
nor U17741 (N_17741,N_17422,N_17365);
nor U17742 (N_17742,N_17427,N_17265);
nor U17743 (N_17743,N_17295,N_17271);
nor U17744 (N_17744,N_17353,N_17364);
nor U17745 (N_17745,N_17273,N_17347);
and U17746 (N_17746,N_17434,N_17397);
and U17747 (N_17747,N_17393,N_17279);
nand U17748 (N_17748,N_17483,N_17442);
and U17749 (N_17749,N_17469,N_17348);
nand U17750 (N_17750,N_17729,N_17727);
nor U17751 (N_17751,N_17582,N_17731);
and U17752 (N_17752,N_17535,N_17632);
nand U17753 (N_17753,N_17741,N_17611);
or U17754 (N_17754,N_17606,N_17531);
nand U17755 (N_17755,N_17537,N_17613);
nand U17756 (N_17756,N_17501,N_17629);
or U17757 (N_17757,N_17721,N_17726);
nand U17758 (N_17758,N_17500,N_17623);
or U17759 (N_17759,N_17749,N_17539);
nand U17760 (N_17760,N_17710,N_17697);
or U17761 (N_17761,N_17585,N_17738);
and U17762 (N_17762,N_17664,N_17517);
and U17763 (N_17763,N_17686,N_17590);
or U17764 (N_17764,N_17707,N_17593);
nor U17765 (N_17765,N_17547,N_17554);
nand U17766 (N_17766,N_17696,N_17739);
nand U17767 (N_17767,N_17532,N_17695);
nor U17768 (N_17768,N_17734,N_17534);
nand U17769 (N_17769,N_17600,N_17676);
nor U17770 (N_17770,N_17617,N_17518);
or U17771 (N_17771,N_17528,N_17591);
nor U17772 (N_17772,N_17589,N_17708);
or U17773 (N_17773,N_17608,N_17634);
nor U17774 (N_17774,N_17574,N_17704);
or U17775 (N_17775,N_17730,N_17713);
nand U17776 (N_17776,N_17723,N_17644);
nor U17777 (N_17777,N_17667,N_17712);
or U17778 (N_17778,N_17627,N_17706);
or U17779 (N_17779,N_17735,N_17603);
or U17780 (N_17780,N_17688,N_17596);
and U17781 (N_17781,N_17551,N_17659);
nor U17782 (N_17782,N_17636,N_17669);
nor U17783 (N_17783,N_17587,N_17642);
and U17784 (N_17784,N_17693,N_17553);
and U17785 (N_17785,N_17510,N_17631);
nor U17786 (N_17786,N_17665,N_17692);
xor U17787 (N_17787,N_17579,N_17572);
nor U17788 (N_17788,N_17702,N_17538);
and U17789 (N_17789,N_17575,N_17542);
nand U17790 (N_17790,N_17577,N_17679);
nand U17791 (N_17791,N_17717,N_17647);
nand U17792 (N_17792,N_17610,N_17663);
nor U17793 (N_17793,N_17609,N_17640);
or U17794 (N_17794,N_17545,N_17645);
or U17795 (N_17795,N_17732,N_17655);
nand U17796 (N_17796,N_17622,N_17715);
nor U17797 (N_17797,N_17556,N_17728);
nand U17798 (N_17798,N_17555,N_17653);
and U17799 (N_17799,N_17615,N_17525);
nor U17800 (N_17800,N_17526,N_17527);
nand U17801 (N_17801,N_17737,N_17700);
nand U17802 (N_17802,N_17658,N_17598);
or U17803 (N_17803,N_17549,N_17683);
nor U17804 (N_17804,N_17509,N_17540);
nor U17805 (N_17805,N_17505,N_17616);
or U17806 (N_17806,N_17668,N_17530);
nor U17807 (N_17807,N_17671,N_17543);
nand U17808 (N_17808,N_17744,N_17557);
or U17809 (N_17809,N_17568,N_17638);
or U17810 (N_17810,N_17595,N_17529);
nor U17811 (N_17811,N_17705,N_17566);
nor U17812 (N_17812,N_17628,N_17504);
or U17813 (N_17813,N_17607,N_17701);
and U17814 (N_17814,N_17612,N_17652);
nor U17815 (N_17815,N_17562,N_17633);
and U17816 (N_17816,N_17586,N_17619);
or U17817 (N_17817,N_17580,N_17604);
or U17818 (N_17818,N_17520,N_17550);
nor U17819 (N_17819,N_17649,N_17524);
and U17820 (N_17820,N_17719,N_17662);
nor U17821 (N_17821,N_17743,N_17694);
and U17822 (N_17822,N_17724,N_17541);
and U17823 (N_17823,N_17747,N_17681);
nand U17824 (N_17824,N_17523,N_17578);
nor U17825 (N_17825,N_17521,N_17740);
nand U17826 (N_17826,N_17650,N_17565);
nand U17827 (N_17827,N_17621,N_17718);
or U17828 (N_17828,N_17716,N_17677);
and U17829 (N_17829,N_17513,N_17745);
nand U17830 (N_17830,N_17552,N_17588);
nand U17831 (N_17831,N_17736,N_17670);
and U17832 (N_17832,N_17584,N_17507);
nand U17833 (N_17833,N_17639,N_17635);
or U17834 (N_17834,N_17680,N_17561);
nor U17835 (N_17835,N_17515,N_17742);
or U17836 (N_17836,N_17625,N_17714);
or U17837 (N_17837,N_17602,N_17559);
nor U17838 (N_17838,N_17657,N_17672);
nand U17839 (N_17839,N_17514,N_17624);
nor U17840 (N_17840,N_17516,N_17626);
and U17841 (N_17841,N_17682,N_17690);
or U17842 (N_17842,N_17605,N_17569);
nand U17843 (N_17843,N_17678,N_17666);
or U17844 (N_17844,N_17648,N_17583);
or U17845 (N_17845,N_17601,N_17685);
nor U17846 (N_17846,N_17506,N_17558);
or U17847 (N_17847,N_17502,N_17560);
nand U17848 (N_17848,N_17675,N_17673);
nor U17849 (N_17849,N_17709,N_17703);
nand U17850 (N_17850,N_17564,N_17711);
or U17851 (N_17851,N_17536,N_17630);
nand U17852 (N_17852,N_17687,N_17641);
nand U17853 (N_17853,N_17620,N_17508);
nand U17854 (N_17854,N_17643,N_17571);
nor U17855 (N_17855,N_17684,N_17592);
nor U17856 (N_17856,N_17614,N_17522);
and U17857 (N_17857,N_17699,N_17573);
and U17858 (N_17858,N_17722,N_17691);
nor U17859 (N_17859,N_17567,N_17599);
nor U17860 (N_17860,N_17544,N_17674);
nor U17861 (N_17861,N_17748,N_17511);
nor U17862 (N_17862,N_17533,N_17594);
nand U17863 (N_17863,N_17661,N_17576);
xor U17864 (N_17864,N_17698,N_17503);
nor U17865 (N_17865,N_17651,N_17637);
and U17866 (N_17866,N_17570,N_17563);
nor U17867 (N_17867,N_17646,N_17548);
xor U17868 (N_17868,N_17660,N_17720);
nand U17869 (N_17869,N_17581,N_17597);
and U17870 (N_17870,N_17519,N_17512);
nor U17871 (N_17871,N_17689,N_17546);
and U17872 (N_17872,N_17654,N_17733);
nand U17873 (N_17873,N_17746,N_17618);
nor U17874 (N_17874,N_17656,N_17725);
or U17875 (N_17875,N_17689,N_17549);
or U17876 (N_17876,N_17685,N_17749);
nor U17877 (N_17877,N_17563,N_17705);
and U17878 (N_17878,N_17671,N_17680);
or U17879 (N_17879,N_17641,N_17642);
xnor U17880 (N_17880,N_17722,N_17628);
nand U17881 (N_17881,N_17611,N_17553);
or U17882 (N_17882,N_17562,N_17579);
and U17883 (N_17883,N_17510,N_17536);
nand U17884 (N_17884,N_17585,N_17568);
xor U17885 (N_17885,N_17640,N_17610);
and U17886 (N_17886,N_17643,N_17599);
nor U17887 (N_17887,N_17661,N_17582);
and U17888 (N_17888,N_17721,N_17677);
nand U17889 (N_17889,N_17696,N_17510);
or U17890 (N_17890,N_17559,N_17694);
nor U17891 (N_17891,N_17636,N_17688);
or U17892 (N_17892,N_17749,N_17548);
and U17893 (N_17893,N_17578,N_17547);
and U17894 (N_17894,N_17730,N_17606);
or U17895 (N_17895,N_17657,N_17569);
nand U17896 (N_17896,N_17714,N_17530);
xnor U17897 (N_17897,N_17573,N_17643);
nand U17898 (N_17898,N_17582,N_17565);
and U17899 (N_17899,N_17734,N_17566);
nor U17900 (N_17900,N_17519,N_17698);
nor U17901 (N_17901,N_17625,N_17697);
or U17902 (N_17902,N_17740,N_17641);
nor U17903 (N_17903,N_17552,N_17645);
nand U17904 (N_17904,N_17585,N_17515);
and U17905 (N_17905,N_17550,N_17710);
or U17906 (N_17906,N_17663,N_17525);
or U17907 (N_17907,N_17525,N_17560);
and U17908 (N_17908,N_17648,N_17568);
nor U17909 (N_17909,N_17503,N_17513);
and U17910 (N_17910,N_17644,N_17635);
nand U17911 (N_17911,N_17597,N_17572);
or U17912 (N_17912,N_17540,N_17727);
and U17913 (N_17913,N_17704,N_17627);
nor U17914 (N_17914,N_17626,N_17598);
nor U17915 (N_17915,N_17505,N_17537);
and U17916 (N_17916,N_17736,N_17716);
and U17917 (N_17917,N_17644,N_17558);
nor U17918 (N_17918,N_17734,N_17560);
nand U17919 (N_17919,N_17597,N_17741);
nor U17920 (N_17920,N_17668,N_17555);
or U17921 (N_17921,N_17662,N_17619);
or U17922 (N_17922,N_17625,N_17597);
nor U17923 (N_17923,N_17512,N_17590);
nand U17924 (N_17924,N_17548,N_17526);
and U17925 (N_17925,N_17705,N_17604);
nor U17926 (N_17926,N_17714,N_17604);
and U17927 (N_17927,N_17546,N_17748);
nor U17928 (N_17928,N_17614,N_17537);
nand U17929 (N_17929,N_17531,N_17743);
and U17930 (N_17930,N_17623,N_17610);
nand U17931 (N_17931,N_17578,N_17519);
nor U17932 (N_17932,N_17556,N_17664);
nor U17933 (N_17933,N_17531,N_17747);
nand U17934 (N_17934,N_17587,N_17577);
and U17935 (N_17935,N_17657,N_17598);
nand U17936 (N_17936,N_17729,N_17560);
nor U17937 (N_17937,N_17672,N_17555);
nor U17938 (N_17938,N_17649,N_17725);
and U17939 (N_17939,N_17529,N_17696);
nand U17940 (N_17940,N_17625,N_17569);
and U17941 (N_17941,N_17549,N_17571);
and U17942 (N_17942,N_17721,N_17667);
nor U17943 (N_17943,N_17726,N_17624);
and U17944 (N_17944,N_17525,N_17700);
nor U17945 (N_17945,N_17637,N_17742);
or U17946 (N_17946,N_17530,N_17570);
nor U17947 (N_17947,N_17634,N_17590);
nor U17948 (N_17948,N_17558,N_17694);
nand U17949 (N_17949,N_17557,N_17539);
and U17950 (N_17950,N_17622,N_17602);
nor U17951 (N_17951,N_17638,N_17567);
or U17952 (N_17952,N_17675,N_17705);
nand U17953 (N_17953,N_17578,N_17657);
nor U17954 (N_17954,N_17705,N_17629);
or U17955 (N_17955,N_17625,N_17512);
nor U17956 (N_17956,N_17622,N_17547);
nor U17957 (N_17957,N_17650,N_17713);
nand U17958 (N_17958,N_17503,N_17669);
or U17959 (N_17959,N_17505,N_17615);
and U17960 (N_17960,N_17730,N_17545);
or U17961 (N_17961,N_17645,N_17553);
nor U17962 (N_17962,N_17734,N_17510);
nand U17963 (N_17963,N_17589,N_17699);
or U17964 (N_17964,N_17664,N_17631);
nand U17965 (N_17965,N_17543,N_17624);
nor U17966 (N_17966,N_17653,N_17693);
and U17967 (N_17967,N_17683,N_17739);
nor U17968 (N_17968,N_17618,N_17513);
or U17969 (N_17969,N_17568,N_17744);
nand U17970 (N_17970,N_17635,N_17660);
nand U17971 (N_17971,N_17689,N_17732);
nor U17972 (N_17972,N_17577,N_17655);
nor U17973 (N_17973,N_17631,N_17722);
or U17974 (N_17974,N_17570,N_17500);
and U17975 (N_17975,N_17500,N_17586);
nand U17976 (N_17976,N_17627,N_17679);
nand U17977 (N_17977,N_17605,N_17636);
and U17978 (N_17978,N_17544,N_17607);
nand U17979 (N_17979,N_17683,N_17681);
nor U17980 (N_17980,N_17722,N_17626);
nor U17981 (N_17981,N_17673,N_17649);
nor U17982 (N_17982,N_17684,N_17563);
and U17983 (N_17983,N_17667,N_17602);
and U17984 (N_17984,N_17719,N_17709);
nor U17985 (N_17985,N_17602,N_17556);
and U17986 (N_17986,N_17504,N_17678);
and U17987 (N_17987,N_17558,N_17675);
or U17988 (N_17988,N_17688,N_17599);
and U17989 (N_17989,N_17704,N_17549);
or U17990 (N_17990,N_17535,N_17595);
or U17991 (N_17991,N_17719,N_17547);
nand U17992 (N_17992,N_17568,N_17701);
nand U17993 (N_17993,N_17608,N_17746);
or U17994 (N_17994,N_17526,N_17505);
and U17995 (N_17995,N_17746,N_17633);
or U17996 (N_17996,N_17681,N_17529);
nor U17997 (N_17997,N_17649,N_17654);
and U17998 (N_17998,N_17594,N_17741);
or U17999 (N_17999,N_17627,N_17541);
or U18000 (N_18000,N_17980,N_17926);
nor U18001 (N_18001,N_17757,N_17835);
or U18002 (N_18002,N_17849,N_17953);
nand U18003 (N_18003,N_17852,N_17839);
or U18004 (N_18004,N_17791,N_17847);
nor U18005 (N_18005,N_17924,N_17758);
nor U18006 (N_18006,N_17827,N_17845);
or U18007 (N_18007,N_17884,N_17761);
nand U18008 (N_18008,N_17778,N_17957);
or U18009 (N_18009,N_17865,N_17972);
or U18010 (N_18010,N_17862,N_17906);
or U18011 (N_18011,N_17796,N_17755);
and U18012 (N_18012,N_17918,N_17903);
or U18013 (N_18013,N_17809,N_17867);
nor U18014 (N_18014,N_17797,N_17858);
and U18015 (N_18015,N_17876,N_17989);
and U18016 (N_18016,N_17805,N_17956);
nand U18017 (N_18017,N_17991,N_17985);
or U18018 (N_18018,N_17823,N_17922);
nand U18019 (N_18019,N_17764,N_17850);
and U18020 (N_18020,N_17766,N_17885);
nor U18021 (N_18021,N_17997,N_17949);
nand U18022 (N_18022,N_17759,N_17792);
and U18023 (N_18023,N_17774,N_17816);
and U18024 (N_18024,N_17905,N_17881);
and U18025 (N_18025,N_17769,N_17784);
or U18026 (N_18026,N_17841,N_17939);
nand U18027 (N_18027,N_17978,N_17836);
and U18028 (N_18028,N_17790,N_17781);
and U18029 (N_18029,N_17783,N_17954);
nand U18030 (N_18030,N_17808,N_17994);
and U18031 (N_18031,N_17813,N_17822);
nand U18032 (N_18032,N_17894,N_17833);
or U18033 (N_18033,N_17904,N_17892);
and U18034 (N_18034,N_17752,N_17819);
or U18035 (N_18035,N_17751,N_17834);
and U18036 (N_18036,N_17853,N_17967);
and U18037 (N_18037,N_17767,N_17898);
nor U18038 (N_18038,N_17795,N_17793);
nor U18039 (N_18039,N_17820,N_17756);
nand U18040 (N_18040,N_17986,N_17958);
or U18041 (N_18041,N_17840,N_17825);
or U18042 (N_18042,N_17977,N_17896);
nor U18043 (N_18043,N_17941,N_17832);
nor U18044 (N_18044,N_17889,N_17928);
and U18045 (N_18045,N_17855,N_17866);
nand U18046 (N_18046,N_17908,N_17937);
nor U18047 (N_18047,N_17948,N_17945);
or U18048 (N_18048,N_17762,N_17899);
or U18049 (N_18049,N_17984,N_17966);
and U18050 (N_18050,N_17817,N_17775);
and U18051 (N_18051,N_17914,N_17801);
nor U18052 (N_18052,N_17963,N_17981);
and U18053 (N_18053,N_17982,N_17869);
and U18054 (N_18054,N_17846,N_17814);
and U18055 (N_18055,N_17848,N_17938);
or U18056 (N_18056,N_17917,N_17976);
nand U18057 (N_18057,N_17975,N_17871);
nand U18058 (N_18058,N_17780,N_17870);
or U18059 (N_18059,N_17999,N_17973);
and U18060 (N_18060,N_17987,N_17887);
nand U18061 (N_18061,N_17873,N_17910);
nor U18062 (N_18062,N_17970,N_17893);
and U18063 (N_18063,N_17803,N_17806);
and U18064 (N_18064,N_17799,N_17824);
nand U18065 (N_18065,N_17837,N_17815);
nand U18066 (N_18066,N_17923,N_17777);
or U18067 (N_18067,N_17979,N_17830);
nand U18068 (N_18068,N_17988,N_17911);
or U18069 (N_18069,N_17753,N_17787);
and U18070 (N_18070,N_17912,N_17961);
nand U18071 (N_18071,N_17786,N_17990);
or U18072 (N_18072,N_17875,N_17965);
or U18073 (N_18073,N_17838,N_17765);
nor U18074 (N_18074,N_17831,N_17807);
nand U18075 (N_18075,N_17851,N_17951);
nand U18076 (N_18076,N_17854,N_17878);
nor U18077 (N_18077,N_17992,N_17930);
or U18078 (N_18078,N_17915,N_17901);
nor U18079 (N_18079,N_17935,N_17864);
nand U18080 (N_18080,N_17828,N_17868);
and U18081 (N_18081,N_17785,N_17789);
or U18082 (N_18082,N_17857,N_17770);
and U18083 (N_18083,N_17750,N_17993);
nand U18084 (N_18084,N_17932,N_17771);
nor U18085 (N_18085,N_17995,N_17947);
nand U18086 (N_18086,N_17944,N_17907);
or U18087 (N_18087,N_17931,N_17810);
nor U18088 (N_18088,N_17843,N_17955);
nand U18089 (N_18089,N_17925,N_17863);
nand U18090 (N_18090,N_17936,N_17798);
and U18091 (N_18091,N_17902,N_17888);
and U18092 (N_18092,N_17818,N_17996);
nand U18093 (N_18093,N_17952,N_17920);
nand U18094 (N_18094,N_17804,N_17763);
or U18095 (N_18095,N_17960,N_17971);
nor U18096 (N_18096,N_17964,N_17895);
or U18097 (N_18097,N_17859,N_17794);
or U18098 (N_18098,N_17890,N_17933);
or U18099 (N_18099,N_17942,N_17940);
nand U18100 (N_18100,N_17998,N_17877);
nand U18101 (N_18101,N_17844,N_17909);
and U18102 (N_18102,N_17934,N_17882);
nand U18103 (N_18103,N_17768,N_17913);
or U18104 (N_18104,N_17929,N_17821);
nand U18105 (N_18105,N_17826,N_17812);
and U18106 (N_18106,N_17874,N_17842);
and U18107 (N_18107,N_17879,N_17860);
nor U18108 (N_18108,N_17927,N_17946);
or U18109 (N_18109,N_17919,N_17891);
nor U18110 (N_18110,N_17897,N_17760);
nand U18111 (N_18111,N_17782,N_17779);
nand U18112 (N_18112,N_17983,N_17916);
nor U18113 (N_18113,N_17883,N_17811);
or U18114 (N_18114,N_17754,N_17776);
and U18115 (N_18115,N_17900,N_17950);
or U18116 (N_18116,N_17968,N_17943);
nand U18117 (N_18117,N_17772,N_17921);
nor U18118 (N_18118,N_17962,N_17872);
nor U18119 (N_18119,N_17829,N_17974);
nand U18120 (N_18120,N_17969,N_17788);
nor U18121 (N_18121,N_17880,N_17861);
nand U18122 (N_18122,N_17886,N_17802);
and U18123 (N_18123,N_17856,N_17959);
and U18124 (N_18124,N_17800,N_17773);
or U18125 (N_18125,N_17889,N_17791);
nand U18126 (N_18126,N_17909,N_17894);
and U18127 (N_18127,N_17797,N_17991);
nor U18128 (N_18128,N_17797,N_17986);
or U18129 (N_18129,N_17864,N_17874);
nand U18130 (N_18130,N_17914,N_17850);
nor U18131 (N_18131,N_17967,N_17891);
or U18132 (N_18132,N_17833,N_17814);
nor U18133 (N_18133,N_17836,N_17778);
and U18134 (N_18134,N_17902,N_17965);
and U18135 (N_18135,N_17953,N_17885);
and U18136 (N_18136,N_17883,N_17755);
nand U18137 (N_18137,N_17891,N_17925);
nand U18138 (N_18138,N_17955,N_17846);
nand U18139 (N_18139,N_17926,N_17989);
and U18140 (N_18140,N_17925,N_17869);
and U18141 (N_18141,N_17927,N_17919);
or U18142 (N_18142,N_17893,N_17833);
and U18143 (N_18143,N_17905,N_17879);
nand U18144 (N_18144,N_17958,N_17944);
or U18145 (N_18145,N_17954,N_17795);
nand U18146 (N_18146,N_17823,N_17804);
or U18147 (N_18147,N_17937,N_17960);
nand U18148 (N_18148,N_17880,N_17982);
nand U18149 (N_18149,N_17963,N_17858);
nand U18150 (N_18150,N_17787,N_17964);
nand U18151 (N_18151,N_17761,N_17780);
nor U18152 (N_18152,N_17798,N_17882);
nand U18153 (N_18153,N_17876,N_17823);
nand U18154 (N_18154,N_17802,N_17900);
nor U18155 (N_18155,N_17841,N_17825);
and U18156 (N_18156,N_17830,N_17928);
nand U18157 (N_18157,N_17835,N_17808);
nor U18158 (N_18158,N_17847,N_17994);
and U18159 (N_18159,N_17967,N_17939);
nand U18160 (N_18160,N_17909,N_17999);
or U18161 (N_18161,N_17782,N_17764);
or U18162 (N_18162,N_17888,N_17807);
nor U18163 (N_18163,N_17998,N_17944);
nor U18164 (N_18164,N_17999,N_17990);
or U18165 (N_18165,N_17961,N_17913);
or U18166 (N_18166,N_17865,N_17850);
or U18167 (N_18167,N_17948,N_17895);
and U18168 (N_18168,N_17862,N_17962);
and U18169 (N_18169,N_17892,N_17924);
nand U18170 (N_18170,N_17970,N_17830);
and U18171 (N_18171,N_17977,N_17995);
and U18172 (N_18172,N_17786,N_17851);
or U18173 (N_18173,N_17813,N_17817);
and U18174 (N_18174,N_17775,N_17786);
nand U18175 (N_18175,N_17773,N_17786);
or U18176 (N_18176,N_17936,N_17988);
or U18177 (N_18177,N_17827,N_17929);
or U18178 (N_18178,N_17897,N_17813);
xnor U18179 (N_18179,N_17780,N_17833);
or U18180 (N_18180,N_17895,N_17780);
or U18181 (N_18181,N_17812,N_17800);
nor U18182 (N_18182,N_17793,N_17825);
or U18183 (N_18183,N_17840,N_17893);
and U18184 (N_18184,N_17775,N_17997);
and U18185 (N_18185,N_17880,N_17826);
or U18186 (N_18186,N_17844,N_17952);
or U18187 (N_18187,N_17934,N_17876);
nor U18188 (N_18188,N_17790,N_17951);
or U18189 (N_18189,N_17872,N_17782);
nor U18190 (N_18190,N_17832,N_17917);
nand U18191 (N_18191,N_17993,N_17815);
and U18192 (N_18192,N_17839,N_17763);
and U18193 (N_18193,N_17841,N_17983);
and U18194 (N_18194,N_17990,N_17836);
nor U18195 (N_18195,N_17878,N_17817);
or U18196 (N_18196,N_17965,N_17821);
and U18197 (N_18197,N_17799,N_17798);
nand U18198 (N_18198,N_17848,N_17879);
nor U18199 (N_18199,N_17871,N_17890);
nand U18200 (N_18200,N_17956,N_17907);
or U18201 (N_18201,N_17914,N_17976);
and U18202 (N_18202,N_17952,N_17983);
or U18203 (N_18203,N_17928,N_17762);
nand U18204 (N_18204,N_17847,N_17936);
or U18205 (N_18205,N_17902,N_17825);
nand U18206 (N_18206,N_17988,N_17945);
or U18207 (N_18207,N_17833,N_17956);
nor U18208 (N_18208,N_17830,N_17905);
and U18209 (N_18209,N_17961,N_17795);
or U18210 (N_18210,N_17971,N_17918);
nand U18211 (N_18211,N_17888,N_17926);
and U18212 (N_18212,N_17981,N_17851);
nor U18213 (N_18213,N_17809,N_17903);
or U18214 (N_18214,N_17888,N_17972);
or U18215 (N_18215,N_17859,N_17934);
and U18216 (N_18216,N_17880,N_17936);
nand U18217 (N_18217,N_17822,N_17777);
or U18218 (N_18218,N_17910,N_17844);
and U18219 (N_18219,N_17989,N_17964);
nand U18220 (N_18220,N_17785,N_17786);
or U18221 (N_18221,N_17838,N_17850);
and U18222 (N_18222,N_17941,N_17919);
and U18223 (N_18223,N_17944,N_17896);
nor U18224 (N_18224,N_17831,N_17784);
nand U18225 (N_18225,N_17781,N_17773);
or U18226 (N_18226,N_17903,N_17997);
and U18227 (N_18227,N_17999,N_17984);
and U18228 (N_18228,N_17844,N_17785);
nand U18229 (N_18229,N_17825,N_17976);
and U18230 (N_18230,N_17779,N_17775);
and U18231 (N_18231,N_17773,N_17904);
and U18232 (N_18232,N_17826,N_17972);
nand U18233 (N_18233,N_17755,N_17811);
nor U18234 (N_18234,N_17828,N_17920);
nor U18235 (N_18235,N_17981,N_17926);
nor U18236 (N_18236,N_17903,N_17864);
or U18237 (N_18237,N_17914,N_17768);
nand U18238 (N_18238,N_17786,N_17772);
nand U18239 (N_18239,N_17914,N_17922);
and U18240 (N_18240,N_17887,N_17934);
nor U18241 (N_18241,N_17969,N_17973);
nor U18242 (N_18242,N_17998,N_17978);
nor U18243 (N_18243,N_17810,N_17852);
or U18244 (N_18244,N_17785,N_17846);
and U18245 (N_18245,N_17948,N_17763);
nor U18246 (N_18246,N_17833,N_17877);
or U18247 (N_18247,N_17963,N_17909);
and U18248 (N_18248,N_17831,N_17930);
or U18249 (N_18249,N_17904,N_17941);
nand U18250 (N_18250,N_18165,N_18173);
nand U18251 (N_18251,N_18241,N_18153);
nand U18252 (N_18252,N_18175,N_18086);
nor U18253 (N_18253,N_18215,N_18189);
nand U18254 (N_18254,N_18155,N_18043);
or U18255 (N_18255,N_18085,N_18192);
nand U18256 (N_18256,N_18007,N_18091);
nand U18257 (N_18257,N_18196,N_18166);
and U18258 (N_18258,N_18191,N_18233);
and U18259 (N_18259,N_18186,N_18059);
and U18260 (N_18260,N_18193,N_18117);
nor U18261 (N_18261,N_18230,N_18225);
nor U18262 (N_18262,N_18167,N_18018);
or U18263 (N_18263,N_18066,N_18161);
or U18264 (N_18264,N_18087,N_18111);
or U18265 (N_18265,N_18152,N_18096);
nor U18266 (N_18266,N_18122,N_18061);
nand U18267 (N_18267,N_18011,N_18158);
or U18268 (N_18268,N_18185,N_18072);
nor U18269 (N_18269,N_18075,N_18058);
or U18270 (N_18270,N_18099,N_18204);
nor U18271 (N_18271,N_18130,N_18178);
nor U18272 (N_18272,N_18201,N_18008);
and U18273 (N_18273,N_18208,N_18194);
nand U18274 (N_18274,N_18013,N_18235);
nor U18275 (N_18275,N_18198,N_18097);
and U18276 (N_18276,N_18114,N_18054);
or U18277 (N_18277,N_18027,N_18071);
and U18278 (N_18278,N_18041,N_18084);
nand U18279 (N_18279,N_18223,N_18222);
nor U18280 (N_18280,N_18141,N_18090);
and U18281 (N_18281,N_18074,N_18213);
or U18282 (N_18282,N_18184,N_18249);
or U18283 (N_18283,N_18144,N_18216);
or U18284 (N_18284,N_18202,N_18199);
or U18285 (N_18285,N_18020,N_18197);
or U18286 (N_18286,N_18177,N_18209);
and U18287 (N_18287,N_18247,N_18021);
nor U18288 (N_18288,N_18147,N_18169);
and U18289 (N_18289,N_18139,N_18120);
or U18290 (N_18290,N_18172,N_18137);
and U18291 (N_18291,N_18163,N_18132);
nor U18292 (N_18292,N_18181,N_18125);
nor U18293 (N_18293,N_18053,N_18157);
nor U18294 (N_18294,N_18131,N_18069);
and U18295 (N_18295,N_18047,N_18179);
or U18296 (N_18296,N_18035,N_18073);
and U18297 (N_18297,N_18156,N_18055);
nand U18298 (N_18298,N_18228,N_18102);
or U18299 (N_18299,N_18109,N_18226);
or U18300 (N_18300,N_18042,N_18010);
and U18301 (N_18301,N_18118,N_18077);
and U18302 (N_18302,N_18174,N_18040);
nand U18303 (N_18303,N_18134,N_18078);
nor U18304 (N_18304,N_18115,N_18211);
or U18305 (N_18305,N_18231,N_18049);
or U18306 (N_18306,N_18187,N_18088);
and U18307 (N_18307,N_18064,N_18103);
or U18308 (N_18308,N_18105,N_18092);
and U18309 (N_18309,N_18128,N_18151);
or U18310 (N_18310,N_18146,N_18205);
nand U18311 (N_18311,N_18026,N_18126);
nand U18312 (N_18312,N_18033,N_18224);
and U18313 (N_18313,N_18210,N_18002);
nor U18314 (N_18314,N_18127,N_18094);
nor U18315 (N_18315,N_18229,N_18168);
nand U18316 (N_18316,N_18046,N_18029);
or U18317 (N_18317,N_18037,N_18065);
nor U18318 (N_18318,N_18060,N_18217);
nor U18319 (N_18319,N_18098,N_18136);
nand U18320 (N_18320,N_18052,N_18039);
nand U18321 (N_18321,N_18237,N_18028);
or U18322 (N_18322,N_18232,N_18057);
nand U18323 (N_18323,N_18110,N_18032);
xor U18324 (N_18324,N_18017,N_18234);
nor U18325 (N_18325,N_18206,N_18089);
nor U18326 (N_18326,N_18081,N_18142);
or U18327 (N_18327,N_18243,N_18143);
or U18328 (N_18328,N_18000,N_18214);
and U18329 (N_18329,N_18176,N_18219);
and U18330 (N_18330,N_18148,N_18082);
nand U18331 (N_18331,N_18068,N_18221);
and U18332 (N_18332,N_18154,N_18116);
nand U18333 (N_18333,N_18006,N_18095);
nor U18334 (N_18334,N_18145,N_18030);
or U18335 (N_18335,N_18200,N_18004);
or U18336 (N_18336,N_18036,N_18083);
nand U18337 (N_18337,N_18014,N_18104);
nand U18338 (N_18338,N_18124,N_18170);
and U18339 (N_18339,N_18079,N_18121);
and U18340 (N_18340,N_18108,N_18164);
nor U18341 (N_18341,N_18016,N_18015);
nand U18342 (N_18342,N_18149,N_18019);
nand U18343 (N_18343,N_18113,N_18248);
nand U18344 (N_18344,N_18044,N_18080);
nand U18345 (N_18345,N_18159,N_18062);
and U18346 (N_18346,N_18107,N_18203);
and U18347 (N_18347,N_18245,N_18180);
nor U18348 (N_18348,N_18022,N_18050);
nand U18349 (N_18349,N_18093,N_18038);
and U18350 (N_18350,N_18025,N_18024);
nor U18351 (N_18351,N_18182,N_18100);
nand U18352 (N_18352,N_18140,N_18171);
and U18353 (N_18353,N_18045,N_18063);
and U18354 (N_18354,N_18001,N_18012);
or U18355 (N_18355,N_18138,N_18218);
or U18356 (N_18356,N_18129,N_18244);
and U18357 (N_18357,N_18227,N_18112);
nand U18358 (N_18358,N_18067,N_18003);
and U18359 (N_18359,N_18236,N_18188);
nor U18360 (N_18360,N_18135,N_18239);
nand U18361 (N_18361,N_18031,N_18190);
or U18362 (N_18362,N_18123,N_18240);
nor U18363 (N_18363,N_18195,N_18238);
or U18364 (N_18364,N_18023,N_18220);
nor U18365 (N_18365,N_18051,N_18246);
or U18366 (N_18366,N_18207,N_18242);
and U18367 (N_18367,N_18150,N_18162);
and U18368 (N_18368,N_18133,N_18160);
nand U18369 (N_18369,N_18183,N_18212);
and U18370 (N_18370,N_18005,N_18056);
and U18371 (N_18371,N_18009,N_18119);
or U18372 (N_18372,N_18048,N_18070);
and U18373 (N_18373,N_18106,N_18101);
or U18374 (N_18374,N_18034,N_18076);
nor U18375 (N_18375,N_18034,N_18025);
and U18376 (N_18376,N_18188,N_18159);
and U18377 (N_18377,N_18078,N_18003);
or U18378 (N_18378,N_18091,N_18201);
or U18379 (N_18379,N_18120,N_18068);
nor U18380 (N_18380,N_18086,N_18212);
nand U18381 (N_18381,N_18229,N_18203);
nor U18382 (N_18382,N_18030,N_18024);
or U18383 (N_18383,N_18113,N_18229);
nor U18384 (N_18384,N_18182,N_18158);
and U18385 (N_18385,N_18128,N_18017);
nor U18386 (N_18386,N_18246,N_18178);
or U18387 (N_18387,N_18198,N_18192);
or U18388 (N_18388,N_18036,N_18225);
nand U18389 (N_18389,N_18133,N_18242);
nor U18390 (N_18390,N_18169,N_18092);
nor U18391 (N_18391,N_18191,N_18187);
or U18392 (N_18392,N_18116,N_18136);
nand U18393 (N_18393,N_18069,N_18165);
nand U18394 (N_18394,N_18238,N_18242);
or U18395 (N_18395,N_18132,N_18037);
nor U18396 (N_18396,N_18044,N_18201);
or U18397 (N_18397,N_18083,N_18201);
and U18398 (N_18398,N_18029,N_18226);
nand U18399 (N_18399,N_18050,N_18104);
nor U18400 (N_18400,N_18065,N_18094);
or U18401 (N_18401,N_18047,N_18245);
and U18402 (N_18402,N_18156,N_18149);
and U18403 (N_18403,N_18237,N_18174);
and U18404 (N_18404,N_18138,N_18174);
nor U18405 (N_18405,N_18006,N_18181);
nor U18406 (N_18406,N_18235,N_18147);
and U18407 (N_18407,N_18006,N_18096);
or U18408 (N_18408,N_18078,N_18175);
and U18409 (N_18409,N_18075,N_18062);
and U18410 (N_18410,N_18191,N_18156);
or U18411 (N_18411,N_18138,N_18124);
or U18412 (N_18412,N_18010,N_18022);
and U18413 (N_18413,N_18081,N_18242);
and U18414 (N_18414,N_18072,N_18219);
or U18415 (N_18415,N_18121,N_18170);
or U18416 (N_18416,N_18149,N_18008);
nor U18417 (N_18417,N_18150,N_18187);
nand U18418 (N_18418,N_18212,N_18218);
and U18419 (N_18419,N_18164,N_18220);
nor U18420 (N_18420,N_18120,N_18005);
or U18421 (N_18421,N_18230,N_18146);
nand U18422 (N_18422,N_18207,N_18008);
and U18423 (N_18423,N_18232,N_18185);
and U18424 (N_18424,N_18230,N_18015);
nor U18425 (N_18425,N_18006,N_18221);
nand U18426 (N_18426,N_18155,N_18075);
and U18427 (N_18427,N_18066,N_18128);
or U18428 (N_18428,N_18064,N_18193);
or U18429 (N_18429,N_18042,N_18065);
xor U18430 (N_18430,N_18075,N_18034);
nand U18431 (N_18431,N_18206,N_18043);
or U18432 (N_18432,N_18165,N_18105);
nor U18433 (N_18433,N_18109,N_18242);
or U18434 (N_18434,N_18133,N_18067);
nand U18435 (N_18435,N_18214,N_18229);
nand U18436 (N_18436,N_18222,N_18111);
nand U18437 (N_18437,N_18100,N_18051);
and U18438 (N_18438,N_18168,N_18132);
nor U18439 (N_18439,N_18009,N_18046);
nand U18440 (N_18440,N_18182,N_18070);
nand U18441 (N_18441,N_18055,N_18179);
nor U18442 (N_18442,N_18025,N_18120);
and U18443 (N_18443,N_18098,N_18021);
or U18444 (N_18444,N_18140,N_18236);
or U18445 (N_18445,N_18059,N_18106);
and U18446 (N_18446,N_18204,N_18145);
nor U18447 (N_18447,N_18016,N_18043);
nand U18448 (N_18448,N_18228,N_18043);
nor U18449 (N_18449,N_18034,N_18072);
nor U18450 (N_18450,N_18093,N_18072);
or U18451 (N_18451,N_18034,N_18013);
or U18452 (N_18452,N_18234,N_18054);
or U18453 (N_18453,N_18102,N_18056);
or U18454 (N_18454,N_18082,N_18169);
nand U18455 (N_18455,N_18218,N_18249);
nand U18456 (N_18456,N_18073,N_18070);
nand U18457 (N_18457,N_18062,N_18136);
and U18458 (N_18458,N_18119,N_18142);
nor U18459 (N_18459,N_18085,N_18028);
and U18460 (N_18460,N_18221,N_18084);
or U18461 (N_18461,N_18012,N_18162);
nand U18462 (N_18462,N_18078,N_18085);
nand U18463 (N_18463,N_18135,N_18081);
nor U18464 (N_18464,N_18130,N_18138);
nand U18465 (N_18465,N_18234,N_18158);
or U18466 (N_18466,N_18054,N_18076);
or U18467 (N_18467,N_18175,N_18242);
nand U18468 (N_18468,N_18082,N_18159);
nand U18469 (N_18469,N_18076,N_18152);
nor U18470 (N_18470,N_18044,N_18234);
or U18471 (N_18471,N_18121,N_18187);
and U18472 (N_18472,N_18093,N_18145);
nor U18473 (N_18473,N_18056,N_18160);
nand U18474 (N_18474,N_18237,N_18166);
and U18475 (N_18475,N_18047,N_18099);
nand U18476 (N_18476,N_18175,N_18178);
nor U18477 (N_18477,N_18078,N_18034);
and U18478 (N_18478,N_18208,N_18024);
nand U18479 (N_18479,N_18185,N_18039);
nand U18480 (N_18480,N_18038,N_18143);
or U18481 (N_18481,N_18170,N_18036);
and U18482 (N_18482,N_18095,N_18163);
nand U18483 (N_18483,N_18190,N_18123);
xnor U18484 (N_18484,N_18200,N_18014);
and U18485 (N_18485,N_18198,N_18071);
nor U18486 (N_18486,N_18010,N_18137);
nor U18487 (N_18487,N_18148,N_18142);
nand U18488 (N_18488,N_18057,N_18215);
or U18489 (N_18489,N_18202,N_18005);
nand U18490 (N_18490,N_18172,N_18100);
nor U18491 (N_18491,N_18204,N_18146);
nor U18492 (N_18492,N_18248,N_18071);
and U18493 (N_18493,N_18085,N_18157);
nand U18494 (N_18494,N_18224,N_18211);
nand U18495 (N_18495,N_18059,N_18009);
and U18496 (N_18496,N_18051,N_18027);
and U18497 (N_18497,N_18201,N_18185);
or U18498 (N_18498,N_18204,N_18025);
or U18499 (N_18499,N_18025,N_18038);
nor U18500 (N_18500,N_18315,N_18441);
nand U18501 (N_18501,N_18496,N_18335);
and U18502 (N_18502,N_18381,N_18261);
nor U18503 (N_18503,N_18397,N_18330);
and U18504 (N_18504,N_18311,N_18491);
nor U18505 (N_18505,N_18332,N_18388);
nor U18506 (N_18506,N_18300,N_18375);
and U18507 (N_18507,N_18259,N_18385);
nand U18508 (N_18508,N_18394,N_18482);
nor U18509 (N_18509,N_18477,N_18488);
nand U18510 (N_18510,N_18449,N_18304);
and U18511 (N_18511,N_18478,N_18379);
nor U18512 (N_18512,N_18461,N_18498);
or U18513 (N_18513,N_18352,N_18299);
nand U18514 (N_18514,N_18278,N_18293);
nand U18515 (N_18515,N_18272,N_18402);
and U18516 (N_18516,N_18319,N_18426);
or U18517 (N_18517,N_18418,N_18376);
or U18518 (N_18518,N_18339,N_18427);
and U18519 (N_18519,N_18382,N_18398);
nand U18520 (N_18520,N_18267,N_18337);
or U18521 (N_18521,N_18322,N_18432);
or U18522 (N_18522,N_18495,N_18333);
and U18523 (N_18523,N_18362,N_18283);
or U18524 (N_18524,N_18301,N_18443);
nand U18525 (N_18525,N_18312,N_18253);
and U18526 (N_18526,N_18371,N_18479);
or U18527 (N_18527,N_18326,N_18417);
nor U18528 (N_18528,N_18303,N_18308);
and U18529 (N_18529,N_18442,N_18314);
nand U18530 (N_18530,N_18399,N_18468);
nor U18531 (N_18531,N_18462,N_18367);
nand U18532 (N_18532,N_18378,N_18305);
nor U18533 (N_18533,N_18291,N_18493);
nand U18534 (N_18534,N_18490,N_18374);
nand U18535 (N_18535,N_18438,N_18358);
or U18536 (N_18536,N_18483,N_18457);
nand U18537 (N_18537,N_18345,N_18331);
or U18538 (N_18538,N_18373,N_18282);
or U18539 (N_18539,N_18392,N_18324);
and U18540 (N_18540,N_18349,N_18307);
and U18541 (N_18541,N_18284,N_18342);
nor U18542 (N_18542,N_18419,N_18444);
or U18543 (N_18543,N_18411,N_18464);
or U18544 (N_18544,N_18273,N_18383);
nor U18545 (N_18545,N_18325,N_18369);
nand U18546 (N_18546,N_18439,N_18310);
and U18547 (N_18547,N_18252,N_18404);
and U18548 (N_18548,N_18389,N_18408);
and U18549 (N_18549,N_18487,N_18455);
or U18550 (N_18550,N_18452,N_18463);
or U18551 (N_18551,N_18258,N_18348);
or U18552 (N_18552,N_18396,N_18285);
and U18553 (N_18553,N_18356,N_18412);
or U18554 (N_18554,N_18409,N_18341);
and U18555 (N_18555,N_18336,N_18391);
nor U18556 (N_18556,N_18360,N_18355);
and U18557 (N_18557,N_18363,N_18286);
nor U18558 (N_18558,N_18485,N_18431);
or U18559 (N_18559,N_18289,N_18370);
or U18560 (N_18560,N_18338,N_18380);
and U18561 (N_18561,N_18274,N_18433);
nor U18562 (N_18562,N_18474,N_18472);
nand U18563 (N_18563,N_18421,N_18250);
nand U18564 (N_18564,N_18458,N_18263);
or U18565 (N_18565,N_18280,N_18422);
or U18566 (N_18566,N_18451,N_18275);
or U18567 (N_18567,N_18271,N_18364);
and U18568 (N_18568,N_18497,N_18454);
or U18569 (N_18569,N_18499,N_18296);
and U18570 (N_18570,N_18302,N_18269);
nand U18571 (N_18571,N_18266,N_18410);
nor U18572 (N_18572,N_18328,N_18471);
nand U18573 (N_18573,N_18453,N_18476);
nand U18574 (N_18574,N_18347,N_18297);
nor U18575 (N_18575,N_18288,N_18424);
and U18576 (N_18576,N_18340,N_18323);
nor U18577 (N_18577,N_18416,N_18413);
nand U18578 (N_18578,N_18465,N_18460);
nor U18579 (N_18579,N_18366,N_18405);
nand U18580 (N_18580,N_18268,N_18334);
or U18581 (N_18581,N_18287,N_18407);
nand U18582 (N_18582,N_18456,N_18329);
or U18583 (N_18583,N_18447,N_18436);
nor U18584 (N_18584,N_18459,N_18466);
or U18585 (N_18585,N_18480,N_18346);
and U18586 (N_18586,N_18414,N_18327);
or U18587 (N_18587,N_18470,N_18377);
nor U18588 (N_18588,N_18486,N_18313);
nand U18589 (N_18589,N_18429,N_18415);
nor U18590 (N_18590,N_18393,N_18386);
nor U18591 (N_18591,N_18469,N_18309);
or U18592 (N_18592,N_18489,N_18292);
and U18593 (N_18593,N_18401,N_18368);
nand U18594 (N_18594,N_18384,N_18492);
nand U18595 (N_18595,N_18318,N_18264);
nor U18596 (N_18596,N_18260,N_18387);
or U18597 (N_18597,N_18255,N_18425);
nand U18598 (N_18598,N_18279,N_18484);
or U18599 (N_18599,N_18434,N_18359);
and U18600 (N_18600,N_18467,N_18350);
nor U18601 (N_18601,N_18357,N_18400);
or U18602 (N_18602,N_18262,N_18361);
nor U18603 (N_18603,N_18372,N_18440);
or U18604 (N_18604,N_18277,N_18306);
or U18605 (N_18605,N_18270,N_18430);
or U18606 (N_18606,N_18256,N_18450);
nor U18607 (N_18607,N_18281,N_18365);
or U18608 (N_18608,N_18276,N_18354);
and U18609 (N_18609,N_18298,N_18475);
nand U18610 (N_18610,N_18316,N_18294);
nand U18611 (N_18611,N_18320,N_18351);
nand U18612 (N_18612,N_18428,N_18445);
and U18613 (N_18613,N_18317,N_18353);
nand U18614 (N_18614,N_18295,N_18265);
nand U18615 (N_18615,N_18420,N_18403);
nor U18616 (N_18616,N_18448,N_18254);
and U18617 (N_18617,N_18435,N_18251);
nand U18618 (N_18618,N_18257,N_18406);
or U18619 (N_18619,N_18321,N_18290);
nor U18620 (N_18620,N_18343,N_18437);
or U18621 (N_18621,N_18446,N_18390);
or U18622 (N_18622,N_18481,N_18494);
nor U18623 (N_18623,N_18344,N_18395);
nand U18624 (N_18624,N_18473,N_18423);
nor U18625 (N_18625,N_18426,N_18361);
nand U18626 (N_18626,N_18337,N_18276);
nor U18627 (N_18627,N_18363,N_18375);
nand U18628 (N_18628,N_18336,N_18372);
or U18629 (N_18629,N_18417,N_18399);
or U18630 (N_18630,N_18442,N_18285);
and U18631 (N_18631,N_18484,N_18285);
and U18632 (N_18632,N_18353,N_18373);
nor U18633 (N_18633,N_18413,N_18386);
nand U18634 (N_18634,N_18346,N_18492);
and U18635 (N_18635,N_18458,N_18486);
nand U18636 (N_18636,N_18365,N_18347);
nand U18637 (N_18637,N_18415,N_18499);
nand U18638 (N_18638,N_18481,N_18286);
nor U18639 (N_18639,N_18477,N_18400);
and U18640 (N_18640,N_18378,N_18291);
nor U18641 (N_18641,N_18459,N_18419);
nand U18642 (N_18642,N_18365,N_18395);
and U18643 (N_18643,N_18474,N_18485);
and U18644 (N_18644,N_18338,N_18289);
nor U18645 (N_18645,N_18265,N_18401);
nand U18646 (N_18646,N_18302,N_18336);
and U18647 (N_18647,N_18489,N_18325);
and U18648 (N_18648,N_18352,N_18401);
nand U18649 (N_18649,N_18449,N_18409);
nor U18650 (N_18650,N_18466,N_18333);
nand U18651 (N_18651,N_18369,N_18450);
or U18652 (N_18652,N_18264,N_18335);
nand U18653 (N_18653,N_18420,N_18417);
and U18654 (N_18654,N_18354,N_18310);
nand U18655 (N_18655,N_18250,N_18431);
nand U18656 (N_18656,N_18263,N_18431);
and U18657 (N_18657,N_18482,N_18339);
nor U18658 (N_18658,N_18335,N_18415);
or U18659 (N_18659,N_18377,N_18417);
or U18660 (N_18660,N_18433,N_18323);
or U18661 (N_18661,N_18377,N_18487);
or U18662 (N_18662,N_18486,N_18390);
and U18663 (N_18663,N_18309,N_18400);
nor U18664 (N_18664,N_18347,N_18323);
or U18665 (N_18665,N_18270,N_18366);
or U18666 (N_18666,N_18432,N_18343);
and U18667 (N_18667,N_18264,N_18479);
or U18668 (N_18668,N_18377,N_18293);
or U18669 (N_18669,N_18398,N_18484);
nand U18670 (N_18670,N_18423,N_18499);
and U18671 (N_18671,N_18495,N_18317);
or U18672 (N_18672,N_18448,N_18403);
nand U18673 (N_18673,N_18336,N_18272);
nor U18674 (N_18674,N_18370,N_18255);
or U18675 (N_18675,N_18430,N_18260);
and U18676 (N_18676,N_18251,N_18436);
nand U18677 (N_18677,N_18285,N_18358);
or U18678 (N_18678,N_18400,N_18436);
and U18679 (N_18679,N_18252,N_18484);
and U18680 (N_18680,N_18325,N_18294);
nor U18681 (N_18681,N_18441,N_18403);
nand U18682 (N_18682,N_18363,N_18330);
nand U18683 (N_18683,N_18423,N_18433);
nand U18684 (N_18684,N_18339,N_18323);
nor U18685 (N_18685,N_18322,N_18254);
nand U18686 (N_18686,N_18357,N_18479);
and U18687 (N_18687,N_18265,N_18398);
and U18688 (N_18688,N_18476,N_18285);
and U18689 (N_18689,N_18430,N_18428);
nand U18690 (N_18690,N_18399,N_18315);
and U18691 (N_18691,N_18480,N_18385);
nor U18692 (N_18692,N_18365,N_18372);
or U18693 (N_18693,N_18435,N_18266);
nand U18694 (N_18694,N_18438,N_18483);
nor U18695 (N_18695,N_18471,N_18433);
nand U18696 (N_18696,N_18356,N_18381);
and U18697 (N_18697,N_18383,N_18289);
and U18698 (N_18698,N_18254,N_18308);
nor U18699 (N_18699,N_18391,N_18459);
or U18700 (N_18700,N_18335,N_18408);
or U18701 (N_18701,N_18435,N_18338);
or U18702 (N_18702,N_18499,N_18276);
nor U18703 (N_18703,N_18363,N_18435);
and U18704 (N_18704,N_18258,N_18265);
nor U18705 (N_18705,N_18496,N_18375);
and U18706 (N_18706,N_18250,N_18305);
nor U18707 (N_18707,N_18375,N_18302);
nor U18708 (N_18708,N_18346,N_18289);
nand U18709 (N_18709,N_18277,N_18251);
or U18710 (N_18710,N_18297,N_18365);
and U18711 (N_18711,N_18406,N_18467);
nand U18712 (N_18712,N_18320,N_18477);
and U18713 (N_18713,N_18386,N_18258);
and U18714 (N_18714,N_18323,N_18370);
and U18715 (N_18715,N_18490,N_18304);
and U18716 (N_18716,N_18274,N_18329);
nor U18717 (N_18717,N_18486,N_18475);
nor U18718 (N_18718,N_18294,N_18323);
nor U18719 (N_18719,N_18472,N_18499);
nor U18720 (N_18720,N_18391,N_18348);
nand U18721 (N_18721,N_18396,N_18321);
or U18722 (N_18722,N_18328,N_18377);
nor U18723 (N_18723,N_18483,N_18439);
and U18724 (N_18724,N_18339,N_18425);
or U18725 (N_18725,N_18373,N_18313);
nand U18726 (N_18726,N_18390,N_18346);
and U18727 (N_18727,N_18322,N_18302);
nand U18728 (N_18728,N_18258,N_18497);
or U18729 (N_18729,N_18291,N_18332);
or U18730 (N_18730,N_18475,N_18450);
nor U18731 (N_18731,N_18329,N_18375);
nand U18732 (N_18732,N_18374,N_18353);
or U18733 (N_18733,N_18436,N_18459);
nor U18734 (N_18734,N_18341,N_18362);
nand U18735 (N_18735,N_18471,N_18495);
nor U18736 (N_18736,N_18259,N_18287);
nand U18737 (N_18737,N_18409,N_18348);
nand U18738 (N_18738,N_18307,N_18250);
xor U18739 (N_18739,N_18321,N_18278);
or U18740 (N_18740,N_18340,N_18250);
nand U18741 (N_18741,N_18453,N_18333);
and U18742 (N_18742,N_18352,N_18434);
and U18743 (N_18743,N_18491,N_18408);
nand U18744 (N_18744,N_18301,N_18354);
or U18745 (N_18745,N_18489,N_18428);
or U18746 (N_18746,N_18305,N_18394);
nand U18747 (N_18747,N_18322,N_18419);
and U18748 (N_18748,N_18388,N_18470);
nor U18749 (N_18749,N_18301,N_18333);
or U18750 (N_18750,N_18530,N_18620);
and U18751 (N_18751,N_18586,N_18612);
nor U18752 (N_18752,N_18602,N_18642);
nor U18753 (N_18753,N_18673,N_18617);
and U18754 (N_18754,N_18600,N_18544);
or U18755 (N_18755,N_18513,N_18564);
nand U18756 (N_18756,N_18587,N_18703);
or U18757 (N_18757,N_18524,N_18581);
nand U18758 (N_18758,N_18724,N_18690);
and U18759 (N_18759,N_18740,N_18507);
and U18760 (N_18760,N_18658,N_18652);
and U18761 (N_18761,N_18582,N_18662);
or U18762 (N_18762,N_18668,N_18599);
nand U18763 (N_18763,N_18726,N_18661);
and U18764 (N_18764,N_18552,N_18626);
and U18765 (N_18765,N_18710,N_18613);
nor U18766 (N_18766,N_18667,N_18562);
nor U18767 (N_18767,N_18611,N_18705);
or U18768 (N_18768,N_18670,N_18715);
or U18769 (N_18769,N_18547,N_18588);
or U18770 (N_18770,N_18559,N_18545);
nand U18771 (N_18771,N_18601,N_18747);
and U18772 (N_18772,N_18614,N_18538);
nand U18773 (N_18773,N_18645,N_18646);
and U18774 (N_18774,N_18501,N_18505);
nor U18775 (N_18775,N_18723,N_18503);
nand U18776 (N_18776,N_18688,N_18536);
nor U18777 (N_18777,N_18636,N_18727);
nand U18778 (N_18778,N_18725,N_18654);
nand U18779 (N_18779,N_18603,N_18627);
nor U18780 (N_18780,N_18735,N_18714);
nor U18781 (N_18781,N_18734,N_18696);
and U18782 (N_18782,N_18584,N_18707);
nand U18783 (N_18783,N_18693,N_18580);
nor U18784 (N_18784,N_18623,N_18593);
nor U18785 (N_18785,N_18649,N_18655);
and U18786 (N_18786,N_18618,N_18730);
nor U18787 (N_18787,N_18567,N_18633);
and U18788 (N_18788,N_18685,N_18678);
or U18789 (N_18789,N_18569,N_18589);
nand U18790 (N_18790,N_18517,N_18519);
nand U18791 (N_18791,N_18669,N_18577);
nor U18792 (N_18792,N_18526,N_18640);
and U18793 (N_18793,N_18651,N_18641);
nor U18794 (N_18794,N_18698,N_18644);
and U18795 (N_18795,N_18543,N_18558);
nor U18796 (N_18796,N_18539,N_18656);
or U18797 (N_18797,N_18728,N_18622);
or U18798 (N_18798,N_18598,N_18729);
nor U18799 (N_18799,N_18571,N_18718);
nand U18800 (N_18800,N_18548,N_18663);
nand U18801 (N_18801,N_18540,N_18709);
nand U18802 (N_18802,N_18511,N_18664);
or U18803 (N_18803,N_18731,N_18606);
and U18804 (N_18804,N_18504,N_18686);
or U18805 (N_18805,N_18736,N_18681);
or U18806 (N_18806,N_18522,N_18509);
nand U18807 (N_18807,N_18637,N_18512);
and U18808 (N_18808,N_18579,N_18721);
nand U18809 (N_18809,N_18672,N_18717);
or U18810 (N_18810,N_18716,N_18563);
nor U18811 (N_18811,N_18719,N_18702);
nand U18812 (N_18812,N_18518,N_18533);
nor U18813 (N_18813,N_18738,N_18607);
nor U18814 (N_18814,N_18619,N_18549);
or U18815 (N_18815,N_18572,N_18625);
and U18816 (N_18816,N_18525,N_18647);
nand U18817 (N_18817,N_18746,N_18510);
nand U18818 (N_18818,N_18534,N_18523);
nor U18819 (N_18819,N_18722,N_18632);
and U18820 (N_18820,N_18706,N_18745);
and U18821 (N_18821,N_18712,N_18648);
nand U18822 (N_18822,N_18554,N_18737);
nor U18823 (N_18823,N_18680,N_18605);
nor U18824 (N_18824,N_18527,N_18568);
or U18825 (N_18825,N_18508,N_18550);
nand U18826 (N_18826,N_18643,N_18628);
and U18827 (N_18827,N_18596,N_18675);
nor U18828 (N_18828,N_18674,N_18555);
or U18829 (N_18829,N_18621,N_18635);
nand U18830 (N_18830,N_18660,N_18700);
nor U18831 (N_18831,N_18741,N_18701);
and U18832 (N_18832,N_18535,N_18575);
or U18833 (N_18833,N_18608,N_18708);
and U18834 (N_18834,N_18665,N_18520);
or U18835 (N_18835,N_18687,N_18748);
and U18836 (N_18836,N_18565,N_18506);
nor U18837 (N_18837,N_18689,N_18743);
nor U18838 (N_18838,N_18624,N_18553);
or U18839 (N_18839,N_18590,N_18542);
or U18840 (N_18840,N_18629,N_18594);
nor U18841 (N_18841,N_18576,N_18695);
and U18842 (N_18842,N_18691,N_18585);
nand U18843 (N_18843,N_18566,N_18657);
or U18844 (N_18844,N_18749,N_18733);
xnor U18845 (N_18845,N_18631,N_18529);
xor U18846 (N_18846,N_18583,N_18595);
or U18847 (N_18847,N_18546,N_18720);
or U18848 (N_18848,N_18638,N_18556);
nor U18849 (N_18849,N_18615,N_18732);
and U18850 (N_18850,N_18516,N_18694);
and U18851 (N_18851,N_18653,N_18573);
and U18852 (N_18852,N_18528,N_18532);
nand U18853 (N_18853,N_18630,N_18610);
and U18854 (N_18854,N_18521,N_18502);
nand U18855 (N_18855,N_18541,N_18591);
and U18856 (N_18856,N_18604,N_18574);
nor U18857 (N_18857,N_18692,N_18561);
or U18858 (N_18858,N_18666,N_18739);
and U18859 (N_18859,N_18634,N_18704);
nand U18860 (N_18860,N_18713,N_18515);
and U18861 (N_18861,N_18650,N_18671);
nand U18862 (N_18862,N_18682,N_18570);
and U18863 (N_18863,N_18578,N_18742);
or U18864 (N_18864,N_18697,N_18744);
nand U18865 (N_18865,N_18699,N_18500);
nand U18866 (N_18866,N_18609,N_18531);
nor U18867 (N_18867,N_18560,N_18639);
nand U18868 (N_18868,N_18537,N_18557);
nand U18869 (N_18869,N_18616,N_18514);
nand U18870 (N_18870,N_18659,N_18683);
nor U18871 (N_18871,N_18676,N_18597);
xnor U18872 (N_18872,N_18684,N_18551);
nor U18873 (N_18873,N_18677,N_18592);
and U18874 (N_18874,N_18711,N_18679);
nor U18875 (N_18875,N_18626,N_18631);
or U18876 (N_18876,N_18744,N_18676);
nor U18877 (N_18877,N_18621,N_18604);
or U18878 (N_18878,N_18512,N_18568);
nor U18879 (N_18879,N_18572,N_18535);
nand U18880 (N_18880,N_18686,N_18554);
nand U18881 (N_18881,N_18724,N_18716);
or U18882 (N_18882,N_18545,N_18636);
nor U18883 (N_18883,N_18646,N_18725);
and U18884 (N_18884,N_18550,N_18547);
or U18885 (N_18885,N_18716,N_18675);
or U18886 (N_18886,N_18512,N_18739);
and U18887 (N_18887,N_18553,N_18536);
nand U18888 (N_18888,N_18521,N_18622);
nand U18889 (N_18889,N_18578,N_18571);
nor U18890 (N_18890,N_18736,N_18588);
nor U18891 (N_18891,N_18678,N_18723);
or U18892 (N_18892,N_18583,N_18616);
and U18893 (N_18893,N_18600,N_18681);
and U18894 (N_18894,N_18672,N_18563);
and U18895 (N_18895,N_18642,N_18624);
nand U18896 (N_18896,N_18697,N_18681);
nor U18897 (N_18897,N_18657,N_18711);
or U18898 (N_18898,N_18717,N_18686);
and U18899 (N_18899,N_18556,N_18702);
and U18900 (N_18900,N_18546,N_18738);
nand U18901 (N_18901,N_18509,N_18734);
or U18902 (N_18902,N_18519,N_18691);
and U18903 (N_18903,N_18553,N_18745);
nand U18904 (N_18904,N_18716,N_18633);
nand U18905 (N_18905,N_18653,N_18537);
and U18906 (N_18906,N_18738,N_18625);
nand U18907 (N_18907,N_18631,N_18639);
nor U18908 (N_18908,N_18561,N_18529);
or U18909 (N_18909,N_18556,N_18617);
or U18910 (N_18910,N_18612,N_18524);
and U18911 (N_18911,N_18618,N_18667);
nor U18912 (N_18912,N_18691,N_18681);
nand U18913 (N_18913,N_18574,N_18533);
xnor U18914 (N_18914,N_18734,N_18516);
and U18915 (N_18915,N_18582,N_18708);
nor U18916 (N_18916,N_18716,N_18729);
nor U18917 (N_18917,N_18652,N_18662);
and U18918 (N_18918,N_18529,N_18709);
and U18919 (N_18919,N_18584,N_18666);
and U18920 (N_18920,N_18636,N_18666);
and U18921 (N_18921,N_18673,N_18583);
nor U18922 (N_18922,N_18599,N_18501);
or U18923 (N_18923,N_18559,N_18729);
nor U18924 (N_18924,N_18573,N_18670);
and U18925 (N_18925,N_18551,N_18584);
and U18926 (N_18926,N_18715,N_18637);
and U18927 (N_18927,N_18578,N_18729);
and U18928 (N_18928,N_18735,N_18549);
nand U18929 (N_18929,N_18664,N_18567);
or U18930 (N_18930,N_18610,N_18736);
xnor U18931 (N_18931,N_18548,N_18710);
nand U18932 (N_18932,N_18646,N_18640);
or U18933 (N_18933,N_18515,N_18610);
or U18934 (N_18934,N_18523,N_18696);
or U18935 (N_18935,N_18714,N_18666);
nor U18936 (N_18936,N_18536,N_18515);
nor U18937 (N_18937,N_18542,N_18586);
or U18938 (N_18938,N_18683,N_18512);
nand U18939 (N_18939,N_18736,N_18694);
and U18940 (N_18940,N_18698,N_18596);
nor U18941 (N_18941,N_18555,N_18517);
or U18942 (N_18942,N_18580,N_18601);
and U18943 (N_18943,N_18509,N_18593);
and U18944 (N_18944,N_18545,N_18663);
nand U18945 (N_18945,N_18587,N_18532);
nand U18946 (N_18946,N_18616,N_18675);
or U18947 (N_18947,N_18574,N_18709);
and U18948 (N_18948,N_18617,N_18701);
nor U18949 (N_18949,N_18598,N_18743);
and U18950 (N_18950,N_18655,N_18714);
or U18951 (N_18951,N_18528,N_18728);
nand U18952 (N_18952,N_18584,N_18746);
nand U18953 (N_18953,N_18556,N_18633);
and U18954 (N_18954,N_18685,N_18593);
nor U18955 (N_18955,N_18606,N_18514);
or U18956 (N_18956,N_18553,N_18718);
nand U18957 (N_18957,N_18519,N_18614);
and U18958 (N_18958,N_18620,N_18615);
nor U18959 (N_18959,N_18737,N_18555);
nor U18960 (N_18960,N_18636,N_18619);
or U18961 (N_18961,N_18551,N_18635);
and U18962 (N_18962,N_18626,N_18566);
nand U18963 (N_18963,N_18513,N_18576);
nand U18964 (N_18964,N_18704,N_18601);
nor U18965 (N_18965,N_18709,N_18713);
or U18966 (N_18966,N_18658,N_18684);
nor U18967 (N_18967,N_18622,N_18645);
and U18968 (N_18968,N_18685,N_18563);
nor U18969 (N_18969,N_18631,N_18693);
or U18970 (N_18970,N_18528,N_18663);
nand U18971 (N_18971,N_18698,N_18686);
or U18972 (N_18972,N_18523,N_18706);
or U18973 (N_18973,N_18697,N_18623);
and U18974 (N_18974,N_18675,N_18728);
and U18975 (N_18975,N_18693,N_18709);
and U18976 (N_18976,N_18683,N_18654);
nand U18977 (N_18977,N_18574,N_18524);
and U18978 (N_18978,N_18588,N_18510);
nand U18979 (N_18979,N_18683,N_18510);
or U18980 (N_18980,N_18533,N_18677);
and U18981 (N_18981,N_18657,N_18522);
or U18982 (N_18982,N_18588,N_18717);
nand U18983 (N_18983,N_18612,N_18672);
nor U18984 (N_18984,N_18674,N_18642);
or U18985 (N_18985,N_18621,N_18676);
or U18986 (N_18986,N_18632,N_18700);
or U18987 (N_18987,N_18550,N_18654);
and U18988 (N_18988,N_18666,N_18608);
nand U18989 (N_18989,N_18504,N_18690);
nor U18990 (N_18990,N_18583,N_18721);
nand U18991 (N_18991,N_18664,N_18601);
and U18992 (N_18992,N_18521,N_18689);
or U18993 (N_18993,N_18609,N_18559);
or U18994 (N_18994,N_18663,N_18500);
xnor U18995 (N_18995,N_18629,N_18680);
nor U18996 (N_18996,N_18535,N_18733);
nand U18997 (N_18997,N_18515,N_18640);
and U18998 (N_18998,N_18717,N_18532);
and U18999 (N_18999,N_18706,N_18511);
or U19000 (N_19000,N_18966,N_18957);
and U19001 (N_19001,N_18760,N_18936);
xnor U19002 (N_19002,N_18789,N_18889);
and U19003 (N_19003,N_18925,N_18846);
nand U19004 (N_19004,N_18807,N_18849);
or U19005 (N_19005,N_18833,N_18796);
or U19006 (N_19006,N_18848,N_18751);
nor U19007 (N_19007,N_18867,N_18941);
or U19008 (N_19008,N_18905,N_18840);
or U19009 (N_19009,N_18860,N_18928);
and U19010 (N_19010,N_18894,N_18971);
or U19011 (N_19011,N_18825,N_18933);
nor U19012 (N_19012,N_18935,N_18986);
or U19013 (N_19013,N_18870,N_18998);
nor U19014 (N_19014,N_18864,N_18979);
and U19015 (N_19015,N_18818,N_18927);
nor U19016 (N_19016,N_18801,N_18806);
nor U19017 (N_19017,N_18978,N_18918);
nand U19018 (N_19018,N_18926,N_18775);
or U19019 (N_19019,N_18809,N_18902);
or U19020 (N_19020,N_18761,N_18871);
and U19021 (N_19021,N_18805,N_18960);
nor U19022 (N_19022,N_18920,N_18874);
nor U19023 (N_19023,N_18947,N_18800);
nand U19024 (N_19024,N_18802,N_18850);
or U19025 (N_19025,N_18768,N_18837);
nand U19026 (N_19026,N_18755,N_18845);
and U19027 (N_19027,N_18811,N_18777);
and U19028 (N_19028,N_18814,N_18753);
and U19029 (N_19029,N_18816,N_18876);
nor U19030 (N_19030,N_18922,N_18788);
or U19031 (N_19031,N_18949,N_18891);
nor U19032 (N_19032,N_18803,N_18893);
nand U19033 (N_19033,N_18985,N_18899);
nand U19034 (N_19034,N_18993,N_18968);
or U19035 (N_19035,N_18924,N_18886);
and U19036 (N_19036,N_18790,N_18911);
nor U19037 (N_19037,N_18835,N_18829);
nor U19038 (N_19038,N_18766,N_18884);
and U19039 (N_19039,N_18955,N_18838);
nor U19040 (N_19040,N_18784,N_18964);
nand U19041 (N_19041,N_18956,N_18822);
or U19042 (N_19042,N_18999,N_18878);
and U19043 (N_19043,N_18916,N_18832);
and U19044 (N_19044,N_18872,N_18974);
nand U19045 (N_19045,N_18810,N_18900);
or U19046 (N_19046,N_18912,N_18930);
nor U19047 (N_19047,N_18754,N_18821);
xor U19048 (N_19048,N_18799,N_18977);
or U19049 (N_19049,N_18831,N_18785);
or U19050 (N_19050,N_18923,N_18750);
nand U19051 (N_19051,N_18781,N_18853);
nand U19052 (N_19052,N_18885,N_18862);
and U19053 (N_19053,N_18765,N_18782);
nor U19054 (N_19054,N_18815,N_18813);
or U19055 (N_19055,N_18762,N_18909);
or U19056 (N_19056,N_18990,N_18841);
nor U19057 (N_19057,N_18827,N_18908);
nand U19058 (N_19058,N_18826,N_18939);
and U19059 (N_19059,N_18887,N_18839);
or U19060 (N_19060,N_18759,N_18919);
or U19061 (N_19061,N_18980,N_18959);
and U19062 (N_19062,N_18921,N_18836);
or U19063 (N_19063,N_18858,N_18962);
nor U19064 (N_19064,N_18896,N_18975);
nor U19065 (N_19065,N_18953,N_18972);
or U19066 (N_19066,N_18812,N_18793);
or U19067 (N_19067,N_18963,N_18830);
nand U19068 (N_19068,N_18844,N_18906);
or U19069 (N_19069,N_18779,N_18770);
nor U19070 (N_19070,N_18847,N_18932);
nor U19071 (N_19071,N_18890,N_18951);
or U19072 (N_19072,N_18969,N_18792);
and U19073 (N_19073,N_18786,N_18954);
nor U19074 (N_19074,N_18958,N_18989);
or U19075 (N_19075,N_18897,N_18945);
nor U19076 (N_19076,N_18970,N_18942);
or U19077 (N_19077,N_18764,N_18776);
nor U19078 (N_19078,N_18791,N_18861);
or U19079 (N_19079,N_18863,N_18946);
nand U19080 (N_19080,N_18882,N_18973);
xor U19081 (N_19081,N_18987,N_18778);
nand U19082 (N_19082,N_18904,N_18903);
and U19083 (N_19083,N_18859,N_18914);
nor U19084 (N_19084,N_18854,N_18895);
nor U19085 (N_19085,N_18856,N_18877);
or U19086 (N_19086,N_18868,N_18931);
or U19087 (N_19087,N_18820,N_18915);
and U19088 (N_19088,N_18881,N_18892);
and U19089 (N_19089,N_18984,N_18866);
or U19090 (N_19090,N_18869,N_18937);
or U19091 (N_19091,N_18763,N_18898);
nand U19092 (N_19092,N_18828,N_18907);
nor U19093 (N_19093,N_18819,N_18769);
or U19094 (N_19094,N_18780,N_18995);
nand U19095 (N_19095,N_18929,N_18804);
or U19096 (N_19096,N_18773,N_18879);
nor U19097 (N_19097,N_18997,N_18943);
and U19098 (N_19098,N_18823,N_18875);
and U19099 (N_19099,N_18852,N_18824);
nor U19100 (N_19100,N_18988,N_18940);
nand U19101 (N_19101,N_18851,N_18880);
and U19102 (N_19102,N_18797,N_18913);
or U19103 (N_19103,N_18873,N_18767);
nand U19104 (N_19104,N_18967,N_18772);
and U19105 (N_19105,N_18817,N_18783);
or U19106 (N_19106,N_18794,N_18865);
nor U19107 (N_19107,N_18976,N_18994);
nor U19108 (N_19108,N_18910,N_18883);
nor U19109 (N_19109,N_18934,N_18774);
nand U19110 (N_19110,N_18888,N_18901);
and U19111 (N_19111,N_18983,N_18996);
nor U19112 (N_19112,N_18834,N_18948);
or U19113 (N_19113,N_18950,N_18991);
nor U19114 (N_19114,N_18771,N_18752);
nor U19115 (N_19115,N_18842,N_18756);
or U19116 (N_19116,N_18757,N_18961);
or U19117 (N_19117,N_18843,N_18944);
nand U19118 (N_19118,N_18855,N_18857);
or U19119 (N_19119,N_18917,N_18758);
nand U19120 (N_19120,N_18981,N_18965);
nand U19121 (N_19121,N_18798,N_18938);
and U19122 (N_19122,N_18795,N_18992);
nand U19123 (N_19123,N_18808,N_18982);
and U19124 (N_19124,N_18952,N_18787);
and U19125 (N_19125,N_18869,N_18987);
and U19126 (N_19126,N_18958,N_18916);
and U19127 (N_19127,N_18878,N_18920);
or U19128 (N_19128,N_18965,N_18764);
nand U19129 (N_19129,N_18905,N_18812);
nor U19130 (N_19130,N_18851,N_18927);
nor U19131 (N_19131,N_18934,N_18895);
nor U19132 (N_19132,N_18836,N_18761);
or U19133 (N_19133,N_18834,N_18827);
nand U19134 (N_19134,N_18814,N_18971);
or U19135 (N_19135,N_18985,N_18816);
nand U19136 (N_19136,N_18953,N_18909);
nor U19137 (N_19137,N_18903,N_18969);
nor U19138 (N_19138,N_18750,N_18854);
or U19139 (N_19139,N_18949,N_18838);
nand U19140 (N_19140,N_18904,N_18974);
or U19141 (N_19141,N_18945,N_18784);
and U19142 (N_19142,N_18829,N_18764);
and U19143 (N_19143,N_18884,N_18921);
nor U19144 (N_19144,N_18994,N_18764);
nor U19145 (N_19145,N_18877,N_18781);
nor U19146 (N_19146,N_18764,N_18926);
and U19147 (N_19147,N_18943,N_18867);
nand U19148 (N_19148,N_18851,N_18900);
or U19149 (N_19149,N_18754,N_18984);
or U19150 (N_19150,N_18875,N_18947);
and U19151 (N_19151,N_18902,N_18833);
and U19152 (N_19152,N_18999,N_18759);
nor U19153 (N_19153,N_18911,N_18822);
nand U19154 (N_19154,N_18949,N_18983);
nor U19155 (N_19155,N_18842,N_18982);
nand U19156 (N_19156,N_18916,N_18787);
or U19157 (N_19157,N_18998,N_18753);
and U19158 (N_19158,N_18902,N_18800);
or U19159 (N_19159,N_18994,N_18964);
nor U19160 (N_19160,N_18898,N_18766);
or U19161 (N_19161,N_18857,N_18776);
nor U19162 (N_19162,N_18866,N_18897);
nor U19163 (N_19163,N_18970,N_18943);
and U19164 (N_19164,N_18860,N_18873);
nand U19165 (N_19165,N_18911,N_18756);
and U19166 (N_19166,N_18782,N_18868);
and U19167 (N_19167,N_18997,N_18892);
nand U19168 (N_19168,N_18793,N_18750);
and U19169 (N_19169,N_18759,N_18765);
nor U19170 (N_19170,N_18809,N_18804);
or U19171 (N_19171,N_18994,N_18885);
nand U19172 (N_19172,N_18881,N_18770);
or U19173 (N_19173,N_18761,N_18954);
nand U19174 (N_19174,N_18935,N_18889);
nand U19175 (N_19175,N_18931,N_18877);
or U19176 (N_19176,N_18941,N_18841);
and U19177 (N_19177,N_18963,N_18890);
or U19178 (N_19178,N_18912,N_18941);
or U19179 (N_19179,N_18971,N_18898);
or U19180 (N_19180,N_18864,N_18808);
nor U19181 (N_19181,N_18992,N_18813);
nand U19182 (N_19182,N_18804,N_18767);
and U19183 (N_19183,N_18817,N_18752);
nand U19184 (N_19184,N_18908,N_18959);
or U19185 (N_19185,N_18886,N_18875);
nor U19186 (N_19186,N_18786,N_18756);
nand U19187 (N_19187,N_18812,N_18768);
nand U19188 (N_19188,N_18772,N_18961);
nor U19189 (N_19189,N_18831,N_18901);
or U19190 (N_19190,N_18801,N_18924);
and U19191 (N_19191,N_18854,N_18932);
nor U19192 (N_19192,N_18780,N_18861);
or U19193 (N_19193,N_18838,N_18911);
and U19194 (N_19194,N_18833,N_18857);
nor U19195 (N_19195,N_18867,N_18875);
nor U19196 (N_19196,N_18774,N_18796);
nand U19197 (N_19197,N_18877,N_18770);
or U19198 (N_19198,N_18835,N_18973);
or U19199 (N_19199,N_18825,N_18787);
nor U19200 (N_19200,N_18893,N_18949);
nor U19201 (N_19201,N_18829,N_18766);
nand U19202 (N_19202,N_18888,N_18999);
or U19203 (N_19203,N_18943,N_18941);
or U19204 (N_19204,N_18912,N_18886);
or U19205 (N_19205,N_18998,N_18960);
nand U19206 (N_19206,N_18828,N_18806);
and U19207 (N_19207,N_18808,N_18983);
nor U19208 (N_19208,N_18864,N_18759);
or U19209 (N_19209,N_18909,N_18949);
and U19210 (N_19210,N_18767,N_18868);
nor U19211 (N_19211,N_18824,N_18969);
nand U19212 (N_19212,N_18907,N_18950);
nand U19213 (N_19213,N_18886,N_18871);
and U19214 (N_19214,N_18830,N_18991);
or U19215 (N_19215,N_18944,N_18966);
nand U19216 (N_19216,N_18933,N_18819);
and U19217 (N_19217,N_18886,N_18806);
nand U19218 (N_19218,N_18956,N_18838);
or U19219 (N_19219,N_18998,N_18795);
nand U19220 (N_19220,N_18884,N_18772);
or U19221 (N_19221,N_18995,N_18931);
or U19222 (N_19222,N_18869,N_18825);
and U19223 (N_19223,N_18837,N_18926);
nand U19224 (N_19224,N_18991,N_18840);
or U19225 (N_19225,N_18774,N_18825);
and U19226 (N_19226,N_18978,N_18763);
nand U19227 (N_19227,N_18889,N_18775);
nand U19228 (N_19228,N_18971,N_18951);
and U19229 (N_19229,N_18990,N_18957);
or U19230 (N_19230,N_18885,N_18818);
nor U19231 (N_19231,N_18801,N_18825);
nor U19232 (N_19232,N_18923,N_18896);
and U19233 (N_19233,N_18841,N_18818);
nor U19234 (N_19234,N_18971,N_18796);
nor U19235 (N_19235,N_18896,N_18870);
and U19236 (N_19236,N_18911,N_18860);
and U19237 (N_19237,N_18820,N_18902);
and U19238 (N_19238,N_18804,N_18920);
and U19239 (N_19239,N_18779,N_18952);
and U19240 (N_19240,N_18895,N_18976);
nor U19241 (N_19241,N_18941,N_18984);
nor U19242 (N_19242,N_18962,N_18850);
nand U19243 (N_19243,N_18877,N_18903);
and U19244 (N_19244,N_18850,N_18896);
and U19245 (N_19245,N_18932,N_18819);
or U19246 (N_19246,N_18784,N_18814);
and U19247 (N_19247,N_18898,N_18940);
nor U19248 (N_19248,N_18971,N_18986);
nand U19249 (N_19249,N_18800,N_18873);
nor U19250 (N_19250,N_19229,N_19180);
nand U19251 (N_19251,N_19101,N_19235);
and U19252 (N_19252,N_19013,N_19084);
and U19253 (N_19253,N_19223,N_19042);
and U19254 (N_19254,N_19183,N_19190);
or U19255 (N_19255,N_19028,N_19140);
nand U19256 (N_19256,N_19018,N_19054);
nor U19257 (N_19257,N_19160,N_19127);
or U19258 (N_19258,N_19184,N_19204);
and U19259 (N_19259,N_19202,N_19166);
nand U19260 (N_19260,N_19164,N_19114);
nor U19261 (N_19261,N_19194,N_19039);
nand U19262 (N_19262,N_19199,N_19002);
nand U19263 (N_19263,N_19227,N_19069);
or U19264 (N_19264,N_19167,N_19044);
or U19265 (N_19265,N_19175,N_19065);
and U19266 (N_19266,N_19106,N_19237);
or U19267 (N_19267,N_19100,N_19049);
and U19268 (N_19268,N_19245,N_19003);
and U19269 (N_19269,N_19083,N_19016);
nor U19270 (N_19270,N_19056,N_19105);
or U19271 (N_19271,N_19045,N_19179);
or U19272 (N_19272,N_19185,N_19080);
and U19273 (N_19273,N_19230,N_19189);
and U19274 (N_19274,N_19144,N_19210);
nor U19275 (N_19275,N_19170,N_19171);
or U19276 (N_19276,N_19238,N_19024);
nand U19277 (N_19277,N_19051,N_19121);
nand U19278 (N_19278,N_19010,N_19151);
or U19279 (N_19279,N_19012,N_19147);
nand U19280 (N_19280,N_19111,N_19015);
nor U19281 (N_19281,N_19120,N_19064);
nor U19282 (N_19282,N_19200,N_19131);
and U19283 (N_19283,N_19040,N_19108);
nand U19284 (N_19284,N_19244,N_19109);
nor U19285 (N_19285,N_19213,N_19197);
or U19286 (N_19286,N_19247,N_19152);
or U19287 (N_19287,N_19103,N_19061);
nor U19288 (N_19288,N_19236,N_19022);
or U19289 (N_19289,N_19163,N_19222);
or U19290 (N_19290,N_19225,N_19186);
nor U19291 (N_19291,N_19123,N_19034);
nand U19292 (N_19292,N_19192,N_19021);
nor U19293 (N_19293,N_19033,N_19072);
nand U19294 (N_19294,N_19214,N_19132);
nor U19295 (N_19295,N_19067,N_19232);
and U19296 (N_19296,N_19217,N_19137);
nand U19297 (N_19297,N_19154,N_19208);
nor U19298 (N_19298,N_19090,N_19148);
or U19299 (N_19299,N_19099,N_19193);
nor U19300 (N_19300,N_19095,N_19143);
nor U19301 (N_19301,N_19240,N_19188);
and U19302 (N_19302,N_19115,N_19216);
and U19303 (N_19303,N_19068,N_19187);
or U19304 (N_19304,N_19070,N_19094);
nor U19305 (N_19305,N_19119,N_19239);
and U19306 (N_19306,N_19159,N_19135);
nor U19307 (N_19307,N_19001,N_19116);
or U19308 (N_19308,N_19058,N_19117);
nand U19309 (N_19309,N_19146,N_19243);
nor U19310 (N_19310,N_19077,N_19172);
nand U19311 (N_19311,N_19052,N_19066);
nand U19312 (N_19312,N_19139,N_19027);
nand U19313 (N_19313,N_19161,N_19141);
and U19314 (N_19314,N_19129,N_19124);
nor U19315 (N_19315,N_19032,N_19110);
and U19316 (N_19316,N_19122,N_19218);
nand U19317 (N_19317,N_19165,N_19221);
nand U19318 (N_19318,N_19036,N_19014);
and U19319 (N_19319,N_19182,N_19037);
nor U19320 (N_19320,N_19025,N_19233);
nor U19321 (N_19321,N_19191,N_19102);
nand U19322 (N_19322,N_19075,N_19162);
nand U19323 (N_19323,N_19053,N_19228);
nand U19324 (N_19324,N_19063,N_19050);
nor U19325 (N_19325,N_19041,N_19035);
nor U19326 (N_19326,N_19215,N_19008);
or U19327 (N_19327,N_19181,N_19136);
or U19328 (N_19328,N_19219,N_19207);
or U19329 (N_19329,N_19005,N_19195);
or U19330 (N_19330,N_19157,N_19011);
nand U19331 (N_19331,N_19085,N_19071);
or U19332 (N_19332,N_19093,N_19059);
or U19333 (N_19333,N_19031,N_19060);
and U19334 (N_19334,N_19019,N_19241);
and U19335 (N_19335,N_19125,N_19091);
nor U19336 (N_19336,N_19089,N_19209);
and U19337 (N_19337,N_19074,N_19020);
nor U19338 (N_19338,N_19096,N_19087);
nand U19339 (N_19339,N_19178,N_19082);
and U19340 (N_19340,N_19150,N_19174);
nor U19341 (N_19341,N_19098,N_19038);
nand U19342 (N_19342,N_19249,N_19062);
nand U19343 (N_19343,N_19023,N_19113);
nand U19344 (N_19344,N_19134,N_19006);
nor U19345 (N_19345,N_19234,N_19176);
xor U19346 (N_19346,N_19198,N_19029);
nand U19347 (N_19347,N_19224,N_19104);
nand U19348 (N_19348,N_19128,N_19242);
and U19349 (N_19349,N_19142,N_19212);
and U19350 (N_19350,N_19126,N_19088);
or U19351 (N_19351,N_19205,N_19158);
nor U19352 (N_19352,N_19226,N_19133);
nor U19353 (N_19353,N_19047,N_19076);
and U19354 (N_19354,N_19118,N_19138);
nand U19355 (N_19355,N_19048,N_19009);
nand U19356 (N_19356,N_19086,N_19173);
nand U19357 (N_19357,N_19155,N_19026);
nor U19358 (N_19358,N_19248,N_19145);
and U19359 (N_19359,N_19004,N_19078);
and U19360 (N_19360,N_19156,N_19220);
nor U19361 (N_19361,N_19203,N_19112);
or U19362 (N_19362,N_19246,N_19057);
nor U19363 (N_19363,N_19097,N_19149);
nand U19364 (N_19364,N_19030,N_19092);
and U19365 (N_19365,N_19231,N_19017);
or U19366 (N_19366,N_19046,N_19079);
nand U19367 (N_19367,N_19073,N_19201);
nor U19368 (N_19368,N_19169,N_19211);
or U19369 (N_19369,N_19168,N_19000);
nand U19370 (N_19370,N_19196,N_19007);
or U19371 (N_19371,N_19130,N_19107);
nor U19372 (N_19372,N_19081,N_19206);
nor U19373 (N_19373,N_19055,N_19043);
nor U19374 (N_19374,N_19153,N_19177);
nor U19375 (N_19375,N_19135,N_19169);
xnor U19376 (N_19376,N_19175,N_19001);
nand U19377 (N_19377,N_19221,N_19139);
and U19378 (N_19378,N_19061,N_19005);
and U19379 (N_19379,N_19164,N_19137);
nor U19380 (N_19380,N_19060,N_19114);
and U19381 (N_19381,N_19158,N_19105);
or U19382 (N_19382,N_19039,N_19131);
nor U19383 (N_19383,N_19195,N_19033);
and U19384 (N_19384,N_19110,N_19195);
or U19385 (N_19385,N_19082,N_19135);
and U19386 (N_19386,N_19067,N_19154);
nand U19387 (N_19387,N_19021,N_19098);
nand U19388 (N_19388,N_19086,N_19098);
and U19389 (N_19389,N_19225,N_19066);
or U19390 (N_19390,N_19241,N_19026);
or U19391 (N_19391,N_19144,N_19167);
nor U19392 (N_19392,N_19096,N_19236);
nor U19393 (N_19393,N_19174,N_19054);
nand U19394 (N_19394,N_19156,N_19168);
nand U19395 (N_19395,N_19131,N_19183);
nand U19396 (N_19396,N_19101,N_19118);
nand U19397 (N_19397,N_19201,N_19225);
nand U19398 (N_19398,N_19216,N_19186);
xor U19399 (N_19399,N_19081,N_19029);
or U19400 (N_19400,N_19019,N_19215);
or U19401 (N_19401,N_19062,N_19034);
and U19402 (N_19402,N_19233,N_19208);
or U19403 (N_19403,N_19135,N_19103);
nor U19404 (N_19404,N_19054,N_19218);
nor U19405 (N_19405,N_19141,N_19078);
and U19406 (N_19406,N_19158,N_19018);
nor U19407 (N_19407,N_19033,N_19144);
nand U19408 (N_19408,N_19065,N_19063);
or U19409 (N_19409,N_19132,N_19162);
and U19410 (N_19410,N_19103,N_19028);
or U19411 (N_19411,N_19075,N_19206);
or U19412 (N_19412,N_19043,N_19034);
nand U19413 (N_19413,N_19099,N_19066);
nand U19414 (N_19414,N_19197,N_19004);
nor U19415 (N_19415,N_19049,N_19147);
or U19416 (N_19416,N_19218,N_19106);
and U19417 (N_19417,N_19015,N_19204);
nand U19418 (N_19418,N_19212,N_19111);
nor U19419 (N_19419,N_19192,N_19115);
and U19420 (N_19420,N_19151,N_19246);
nor U19421 (N_19421,N_19245,N_19172);
nor U19422 (N_19422,N_19062,N_19133);
nor U19423 (N_19423,N_19212,N_19084);
nand U19424 (N_19424,N_19126,N_19157);
and U19425 (N_19425,N_19036,N_19015);
nand U19426 (N_19426,N_19085,N_19114);
nor U19427 (N_19427,N_19115,N_19102);
or U19428 (N_19428,N_19072,N_19139);
or U19429 (N_19429,N_19107,N_19214);
nand U19430 (N_19430,N_19165,N_19105);
or U19431 (N_19431,N_19216,N_19241);
nand U19432 (N_19432,N_19158,N_19000);
nor U19433 (N_19433,N_19000,N_19132);
nor U19434 (N_19434,N_19102,N_19011);
and U19435 (N_19435,N_19053,N_19137);
nand U19436 (N_19436,N_19136,N_19089);
or U19437 (N_19437,N_19175,N_19152);
or U19438 (N_19438,N_19092,N_19099);
nand U19439 (N_19439,N_19047,N_19234);
and U19440 (N_19440,N_19119,N_19196);
and U19441 (N_19441,N_19176,N_19206);
or U19442 (N_19442,N_19048,N_19113);
or U19443 (N_19443,N_19050,N_19008);
nor U19444 (N_19444,N_19114,N_19172);
nor U19445 (N_19445,N_19249,N_19012);
xnor U19446 (N_19446,N_19238,N_19244);
or U19447 (N_19447,N_19121,N_19118);
and U19448 (N_19448,N_19178,N_19008);
nand U19449 (N_19449,N_19078,N_19216);
nand U19450 (N_19450,N_19087,N_19240);
nor U19451 (N_19451,N_19144,N_19056);
or U19452 (N_19452,N_19028,N_19136);
and U19453 (N_19453,N_19107,N_19211);
and U19454 (N_19454,N_19180,N_19021);
nand U19455 (N_19455,N_19076,N_19023);
and U19456 (N_19456,N_19142,N_19241);
and U19457 (N_19457,N_19079,N_19142);
and U19458 (N_19458,N_19217,N_19094);
nand U19459 (N_19459,N_19216,N_19246);
nor U19460 (N_19460,N_19019,N_19196);
and U19461 (N_19461,N_19091,N_19026);
xnor U19462 (N_19462,N_19124,N_19195);
and U19463 (N_19463,N_19059,N_19079);
nor U19464 (N_19464,N_19048,N_19071);
or U19465 (N_19465,N_19043,N_19201);
and U19466 (N_19466,N_19057,N_19053);
nor U19467 (N_19467,N_19173,N_19217);
nor U19468 (N_19468,N_19135,N_19186);
and U19469 (N_19469,N_19011,N_19034);
or U19470 (N_19470,N_19232,N_19094);
nor U19471 (N_19471,N_19089,N_19056);
or U19472 (N_19472,N_19185,N_19019);
or U19473 (N_19473,N_19112,N_19029);
or U19474 (N_19474,N_19143,N_19010);
and U19475 (N_19475,N_19248,N_19131);
and U19476 (N_19476,N_19150,N_19136);
nand U19477 (N_19477,N_19061,N_19117);
and U19478 (N_19478,N_19083,N_19091);
nor U19479 (N_19479,N_19111,N_19167);
nand U19480 (N_19480,N_19175,N_19168);
nor U19481 (N_19481,N_19068,N_19230);
and U19482 (N_19482,N_19149,N_19020);
or U19483 (N_19483,N_19118,N_19152);
and U19484 (N_19484,N_19035,N_19121);
and U19485 (N_19485,N_19044,N_19139);
and U19486 (N_19486,N_19138,N_19119);
and U19487 (N_19487,N_19080,N_19221);
and U19488 (N_19488,N_19117,N_19067);
and U19489 (N_19489,N_19055,N_19050);
nor U19490 (N_19490,N_19184,N_19169);
nor U19491 (N_19491,N_19240,N_19212);
or U19492 (N_19492,N_19019,N_19179);
or U19493 (N_19493,N_19166,N_19066);
and U19494 (N_19494,N_19041,N_19012);
or U19495 (N_19495,N_19068,N_19150);
or U19496 (N_19496,N_19182,N_19013);
or U19497 (N_19497,N_19145,N_19234);
nand U19498 (N_19498,N_19107,N_19035);
nand U19499 (N_19499,N_19073,N_19044);
or U19500 (N_19500,N_19340,N_19396);
nand U19501 (N_19501,N_19439,N_19425);
and U19502 (N_19502,N_19298,N_19277);
or U19503 (N_19503,N_19359,N_19457);
nand U19504 (N_19504,N_19366,N_19361);
nand U19505 (N_19505,N_19479,N_19471);
nand U19506 (N_19506,N_19349,N_19290);
or U19507 (N_19507,N_19369,N_19323);
or U19508 (N_19508,N_19266,N_19311);
nor U19509 (N_19509,N_19318,N_19449);
or U19510 (N_19510,N_19496,N_19360);
or U19511 (N_19511,N_19453,N_19443);
nand U19512 (N_19512,N_19476,N_19417);
nor U19513 (N_19513,N_19406,N_19351);
and U19514 (N_19514,N_19285,N_19488);
nor U19515 (N_19515,N_19489,N_19296);
nor U19516 (N_19516,N_19348,N_19353);
and U19517 (N_19517,N_19459,N_19436);
and U19518 (N_19518,N_19268,N_19368);
nand U19519 (N_19519,N_19448,N_19293);
and U19520 (N_19520,N_19251,N_19344);
nor U19521 (N_19521,N_19402,N_19352);
and U19522 (N_19522,N_19398,N_19421);
and U19523 (N_19523,N_19338,N_19445);
or U19524 (N_19524,N_19335,N_19450);
nand U19525 (N_19525,N_19393,N_19464);
nand U19526 (N_19526,N_19495,N_19317);
nor U19527 (N_19527,N_19250,N_19434);
nand U19528 (N_19528,N_19265,N_19438);
nor U19529 (N_19529,N_19283,N_19383);
and U19530 (N_19530,N_19331,N_19334);
and U19531 (N_19531,N_19339,N_19392);
or U19532 (N_19532,N_19423,N_19465);
or U19533 (N_19533,N_19345,N_19269);
or U19534 (N_19534,N_19254,N_19253);
and U19535 (N_19535,N_19259,N_19374);
nor U19536 (N_19536,N_19286,N_19400);
nor U19537 (N_19537,N_19395,N_19307);
nor U19538 (N_19538,N_19433,N_19258);
nor U19539 (N_19539,N_19410,N_19305);
and U19540 (N_19540,N_19316,N_19312);
nand U19541 (N_19541,N_19274,N_19446);
or U19542 (N_19542,N_19327,N_19412);
and U19543 (N_19543,N_19407,N_19405);
and U19544 (N_19544,N_19456,N_19263);
and U19545 (N_19545,N_19382,N_19288);
and U19546 (N_19546,N_19363,N_19435);
and U19547 (N_19547,N_19376,N_19300);
nor U19548 (N_19548,N_19420,N_19431);
and U19549 (N_19549,N_19452,N_19291);
or U19550 (N_19550,N_19267,N_19493);
and U19551 (N_19551,N_19252,N_19264);
and U19552 (N_19552,N_19299,N_19272);
nor U19553 (N_19553,N_19454,N_19362);
and U19554 (N_19554,N_19306,N_19325);
xnor U19555 (N_19555,N_19409,N_19469);
nand U19556 (N_19556,N_19364,N_19429);
and U19557 (N_19557,N_19278,N_19365);
nand U19558 (N_19558,N_19473,N_19371);
nand U19559 (N_19559,N_19416,N_19329);
nand U19560 (N_19560,N_19458,N_19411);
xnor U19561 (N_19561,N_19481,N_19455);
nand U19562 (N_19562,N_19432,N_19480);
nand U19563 (N_19563,N_19463,N_19372);
nand U19564 (N_19564,N_19320,N_19355);
and U19565 (N_19565,N_19482,N_19381);
and U19566 (N_19566,N_19295,N_19273);
or U19567 (N_19567,N_19377,N_19346);
or U19568 (N_19568,N_19328,N_19403);
and U19569 (N_19569,N_19271,N_19387);
or U19570 (N_19570,N_19260,N_19297);
nor U19571 (N_19571,N_19483,N_19379);
and U19572 (N_19572,N_19484,N_19408);
nor U19573 (N_19573,N_19342,N_19442);
nor U19574 (N_19574,N_19444,N_19310);
and U19575 (N_19575,N_19289,N_19462);
or U19576 (N_19576,N_19422,N_19401);
or U19577 (N_19577,N_19428,N_19279);
nand U19578 (N_19578,N_19261,N_19385);
or U19579 (N_19579,N_19497,N_19414);
nor U19580 (N_19580,N_19324,N_19294);
and U19581 (N_19581,N_19380,N_19315);
nor U19582 (N_19582,N_19321,N_19451);
or U19583 (N_19583,N_19499,N_19337);
or U19584 (N_19584,N_19378,N_19468);
nand U19585 (N_19585,N_19322,N_19319);
nor U19586 (N_19586,N_19257,N_19472);
and U19587 (N_19587,N_19301,N_19326);
or U19588 (N_19588,N_19440,N_19491);
nor U19589 (N_19589,N_19437,N_19354);
or U19590 (N_19590,N_19292,N_19478);
nor U19591 (N_19591,N_19370,N_19492);
and U19592 (N_19592,N_19313,N_19494);
nor U19593 (N_19593,N_19276,N_19341);
nor U19594 (N_19594,N_19397,N_19486);
or U19595 (N_19595,N_19389,N_19375);
or U19596 (N_19596,N_19343,N_19302);
or U19597 (N_19597,N_19373,N_19388);
and U19598 (N_19598,N_19485,N_19447);
nor U19599 (N_19599,N_19282,N_19308);
and U19600 (N_19600,N_19430,N_19303);
or U19601 (N_19601,N_19270,N_19415);
nand U19602 (N_19602,N_19424,N_19404);
nor U19603 (N_19603,N_19426,N_19441);
and U19604 (N_19604,N_19390,N_19427);
nand U19605 (N_19605,N_19418,N_19280);
nor U19606 (N_19606,N_19498,N_19461);
nor U19607 (N_19607,N_19314,N_19332);
nand U19608 (N_19608,N_19367,N_19466);
nand U19609 (N_19609,N_19487,N_19474);
nand U19610 (N_19610,N_19336,N_19399);
and U19611 (N_19611,N_19287,N_19255);
and U19612 (N_19612,N_19309,N_19460);
nor U19613 (N_19613,N_19330,N_19281);
or U19614 (N_19614,N_19413,N_19347);
or U19615 (N_19615,N_19490,N_19284);
or U19616 (N_19616,N_19384,N_19357);
or U19617 (N_19617,N_19333,N_19475);
and U19618 (N_19618,N_19419,N_19391);
or U19619 (N_19619,N_19477,N_19356);
or U19620 (N_19620,N_19350,N_19386);
nand U19621 (N_19621,N_19304,N_19256);
nand U19622 (N_19622,N_19467,N_19470);
and U19623 (N_19623,N_19275,N_19358);
and U19624 (N_19624,N_19394,N_19262);
or U19625 (N_19625,N_19271,N_19395);
nand U19626 (N_19626,N_19432,N_19360);
nor U19627 (N_19627,N_19493,N_19381);
or U19628 (N_19628,N_19339,N_19419);
and U19629 (N_19629,N_19261,N_19390);
and U19630 (N_19630,N_19462,N_19251);
or U19631 (N_19631,N_19410,N_19472);
nor U19632 (N_19632,N_19311,N_19443);
nor U19633 (N_19633,N_19361,N_19419);
nor U19634 (N_19634,N_19481,N_19287);
and U19635 (N_19635,N_19480,N_19274);
and U19636 (N_19636,N_19347,N_19378);
nor U19637 (N_19637,N_19335,N_19266);
and U19638 (N_19638,N_19422,N_19491);
nor U19639 (N_19639,N_19380,N_19469);
or U19640 (N_19640,N_19473,N_19453);
or U19641 (N_19641,N_19499,N_19454);
nand U19642 (N_19642,N_19492,N_19402);
or U19643 (N_19643,N_19407,N_19421);
and U19644 (N_19644,N_19384,N_19342);
nand U19645 (N_19645,N_19429,N_19346);
and U19646 (N_19646,N_19485,N_19345);
and U19647 (N_19647,N_19274,N_19385);
nor U19648 (N_19648,N_19328,N_19293);
nand U19649 (N_19649,N_19288,N_19319);
nor U19650 (N_19650,N_19415,N_19357);
and U19651 (N_19651,N_19360,N_19393);
or U19652 (N_19652,N_19364,N_19478);
nand U19653 (N_19653,N_19398,N_19382);
nand U19654 (N_19654,N_19274,N_19497);
and U19655 (N_19655,N_19344,N_19372);
or U19656 (N_19656,N_19455,N_19447);
nor U19657 (N_19657,N_19464,N_19349);
or U19658 (N_19658,N_19330,N_19475);
and U19659 (N_19659,N_19271,N_19258);
and U19660 (N_19660,N_19349,N_19410);
or U19661 (N_19661,N_19283,N_19411);
nor U19662 (N_19662,N_19406,N_19344);
and U19663 (N_19663,N_19365,N_19498);
nor U19664 (N_19664,N_19459,N_19371);
and U19665 (N_19665,N_19401,N_19427);
nor U19666 (N_19666,N_19343,N_19497);
or U19667 (N_19667,N_19289,N_19357);
nand U19668 (N_19668,N_19360,N_19385);
or U19669 (N_19669,N_19320,N_19440);
or U19670 (N_19670,N_19454,N_19300);
nor U19671 (N_19671,N_19323,N_19358);
and U19672 (N_19672,N_19494,N_19291);
nor U19673 (N_19673,N_19354,N_19269);
and U19674 (N_19674,N_19393,N_19254);
or U19675 (N_19675,N_19274,N_19357);
nor U19676 (N_19676,N_19276,N_19480);
and U19677 (N_19677,N_19287,N_19263);
nand U19678 (N_19678,N_19281,N_19417);
nor U19679 (N_19679,N_19325,N_19350);
and U19680 (N_19680,N_19446,N_19344);
nor U19681 (N_19681,N_19281,N_19448);
or U19682 (N_19682,N_19269,N_19291);
xnor U19683 (N_19683,N_19283,N_19250);
or U19684 (N_19684,N_19337,N_19370);
nor U19685 (N_19685,N_19451,N_19460);
and U19686 (N_19686,N_19455,N_19317);
and U19687 (N_19687,N_19327,N_19422);
or U19688 (N_19688,N_19475,N_19366);
nor U19689 (N_19689,N_19421,N_19488);
nor U19690 (N_19690,N_19416,N_19372);
nor U19691 (N_19691,N_19298,N_19380);
nand U19692 (N_19692,N_19322,N_19405);
nor U19693 (N_19693,N_19423,N_19367);
nand U19694 (N_19694,N_19414,N_19314);
or U19695 (N_19695,N_19317,N_19348);
and U19696 (N_19696,N_19257,N_19326);
nor U19697 (N_19697,N_19376,N_19326);
and U19698 (N_19698,N_19442,N_19291);
nor U19699 (N_19699,N_19497,N_19474);
nor U19700 (N_19700,N_19379,N_19255);
or U19701 (N_19701,N_19417,N_19382);
nand U19702 (N_19702,N_19383,N_19279);
and U19703 (N_19703,N_19306,N_19356);
nand U19704 (N_19704,N_19397,N_19291);
nand U19705 (N_19705,N_19498,N_19438);
and U19706 (N_19706,N_19445,N_19323);
nand U19707 (N_19707,N_19322,N_19352);
or U19708 (N_19708,N_19362,N_19466);
nor U19709 (N_19709,N_19325,N_19452);
nor U19710 (N_19710,N_19384,N_19317);
xnor U19711 (N_19711,N_19422,N_19404);
nor U19712 (N_19712,N_19259,N_19471);
and U19713 (N_19713,N_19438,N_19372);
nor U19714 (N_19714,N_19376,N_19299);
nand U19715 (N_19715,N_19274,N_19295);
nand U19716 (N_19716,N_19290,N_19435);
nand U19717 (N_19717,N_19264,N_19425);
nor U19718 (N_19718,N_19277,N_19394);
or U19719 (N_19719,N_19426,N_19366);
nand U19720 (N_19720,N_19255,N_19328);
and U19721 (N_19721,N_19412,N_19376);
and U19722 (N_19722,N_19362,N_19288);
nand U19723 (N_19723,N_19279,N_19482);
or U19724 (N_19724,N_19482,N_19479);
or U19725 (N_19725,N_19270,N_19459);
and U19726 (N_19726,N_19474,N_19459);
nand U19727 (N_19727,N_19341,N_19402);
and U19728 (N_19728,N_19456,N_19369);
and U19729 (N_19729,N_19385,N_19465);
nand U19730 (N_19730,N_19280,N_19444);
and U19731 (N_19731,N_19469,N_19395);
nor U19732 (N_19732,N_19328,N_19332);
and U19733 (N_19733,N_19466,N_19313);
nand U19734 (N_19734,N_19389,N_19252);
and U19735 (N_19735,N_19472,N_19467);
nor U19736 (N_19736,N_19388,N_19381);
nand U19737 (N_19737,N_19351,N_19462);
nor U19738 (N_19738,N_19325,N_19336);
or U19739 (N_19739,N_19272,N_19472);
nor U19740 (N_19740,N_19258,N_19461);
and U19741 (N_19741,N_19348,N_19261);
nand U19742 (N_19742,N_19258,N_19482);
or U19743 (N_19743,N_19274,N_19270);
nor U19744 (N_19744,N_19376,N_19342);
or U19745 (N_19745,N_19289,N_19465);
nor U19746 (N_19746,N_19386,N_19348);
or U19747 (N_19747,N_19401,N_19482);
and U19748 (N_19748,N_19465,N_19362);
nor U19749 (N_19749,N_19271,N_19400);
or U19750 (N_19750,N_19598,N_19633);
and U19751 (N_19751,N_19560,N_19626);
nand U19752 (N_19752,N_19713,N_19570);
nor U19753 (N_19753,N_19660,N_19621);
nand U19754 (N_19754,N_19706,N_19641);
nor U19755 (N_19755,N_19721,N_19656);
nand U19756 (N_19756,N_19515,N_19675);
nor U19757 (N_19757,N_19666,N_19501);
nor U19758 (N_19758,N_19748,N_19541);
nor U19759 (N_19759,N_19720,N_19636);
or U19760 (N_19760,N_19712,N_19571);
nand U19761 (N_19761,N_19627,N_19655);
nand U19762 (N_19762,N_19503,N_19579);
nand U19763 (N_19763,N_19601,N_19595);
or U19764 (N_19764,N_19698,N_19645);
nand U19765 (N_19765,N_19550,N_19718);
nand U19766 (N_19766,N_19743,N_19745);
nand U19767 (N_19767,N_19527,N_19671);
nor U19768 (N_19768,N_19646,N_19679);
nor U19769 (N_19769,N_19735,N_19584);
nand U19770 (N_19770,N_19510,N_19522);
nor U19771 (N_19771,N_19676,N_19524);
and U19772 (N_19772,N_19557,N_19723);
nand U19773 (N_19773,N_19521,N_19622);
or U19774 (N_19774,N_19613,N_19523);
or U19775 (N_19775,N_19661,N_19744);
nand U19776 (N_19776,N_19518,N_19673);
nor U19777 (N_19777,N_19746,N_19556);
nor U19778 (N_19778,N_19709,N_19725);
or U19779 (N_19779,N_19504,N_19545);
or U19780 (N_19780,N_19564,N_19596);
or U19781 (N_19781,N_19617,N_19525);
nor U19782 (N_19782,N_19719,N_19586);
or U19783 (N_19783,N_19508,N_19726);
and U19784 (N_19784,N_19511,N_19705);
nor U19785 (N_19785,N_19701,N_19702);
and U19786 (N_19786,N_19734,N_19670);
and U19787 (N_19787,N_19659,N_19509);
or U19788 (N_19788,N_19517,N_19665);
and U19789 (N_19789,N_19519,N_19620);
nand U19790 (N_19790,N_19590,N_19730);
nor U19791 (N_19791,N_19559,N_19500);
nor U19792 (N_19792,N_19604,N_19609);
nor U19793 (N_19793,N_19737,N_19612);
nor U19794 (N_19794,N_19693,N_19543);
nand U19795 (N_19795,N_19635,N_19736);
nand U19796 (N_19796,N_19710,N_19724);
and U19797 (N_19797,N_19630,N_19513);
or U19798 (N_19798,N_19614,N_19669);
and U19799 (N_19799,N_19667,N_19644);
and U19800 (N_19800,N_19534,N_19749);
or U19801 (N_19801,N_19615,N_19638);
nand U19802 (N_19802,N_19547,N_19649);
and U19803 (N_19803,N_19647,N_19592);
and U19804 (N_19804,N_19682,N_19632);
or U19805 (N_19805,N_19618,N_19568);
nor U19806 (N_19806,N_19738,N_19722);
nand U19807 (N_19807,N_19600,N_19603);
and U19808 (N_19808,N_19537,N_19739);
and U19809 (N_19809,N_19551,N_19565);
and U19810 (N_19810,N_19689,N_19623);
nand U19811 (N_19811,N_19505,N_19587);
nand U19812 (N_19812,N_19740,N_19628);
nand U19813 (N_19813,N_19696,N_19573);
nand U19814 (N_19814,N_19697,N_19566);
nor U19815 (N_19815,N_19715,N_19686);
and U19816 (N_19816,N_19528,N_19678);
or U19817 (N_19817,N_19652,N_19514);
nand U19818 (N_19818,N_19576,N_19585);
or U19819 (N_19819,N_19681,N_19529);
or U19820 (N_19820,N_19574,N_19555);
nand U19821 (N_19821,N_19677,N_19602);
or U19822 (N_19822,N_19512,N_19688);
nand U19823 (N_19823,N_19594,N_19629);
or U19824 (N_19824,N_19731,N_19732);
nor U19825 (N_19825,N_19599,N_19728);
nor U19826 (N_19826,N_19544,N_19711);
nor U19827 (N_19827,N_19563,N_19577);
or U19828 (N_19828,N_19692,N_19733);
nor U19829 (N_19829,N_19593,N_19658);
nand U19830 (N_19830,N_19639,N_19704);
nor U19831 (N_19831,N_19554,N_19664);
nand U19832 (N_19832,N_19727,N_19502);
and U19833 (N_19833,N_19624,N_19703);
or U19834 (N_19834,N_19606,N_19625);
nor U19835 (N_19835,N_19680,N_19663);
nor U19836 (N_19836,N_19516,N_19668);
nor U19837 (N_19837,N_19631,N_19538);
or U19838 (N_19838,N_19605,N_19540);
nand U19839 (N_19839,N_19552,N_19526);
nand U19840 (N_19840,N_19648,N_19691);
nand U19841 (N_19841,N_19684,N_19674);
nand U19842 (N_19842,N_19690,N_19533);
or U19843 (N_19843,N_19610,N_19597);
nand U19844 (N_19844,N_19536,N_19687);
nor U19845 (N_19845,N_19707,N_19507);
or U19846 (N_19846,N_19531,N_19716);
and U19847 (N_19847,N_19542,N_19549);
or U19848 (N_19848,N_19562,N_19535);
and U19849 (N_19849,N_19672,N_19608);
or U19850 (N_19850,N_19654,N_19685);
and U19851 (N_19851,N_19683,N_19619);
or U19852 (N_19852,N_19583,N_19506);
nor U19853 (N_19853,N_19561,N_19657);
nand U19854 (N_19854,N_19548,N_19589);
nand U19855 (N_19855,N_19651,N_19575);
or U19856 (N_19856,N_19642,N_19582);
nand U19857 (N_19857,N_19634,N_19567);
nor U19858 (N_19858,N_19714,N_19742);
nor U19859 (N_19859,N_19580,N_19611);
nand U19860 (N_19860,N_19581,N_19578);
nand U19861 (N_19861,N_19694,N_19569);
nand U19862 (N_19862,N_19532,N_19700);
nand U19863 (N_19863,N_19558,N_19616);
nor U19864 (N_19864,N_19643,N_19572);
nand U19865 (N_19865,N_19729,N_19653);
or U19866 (N_19866,N_19708,N_19588);
xor U19867 (N_19867,N_19747,N_19695);
or U19868 (N_19868,N_19640,N_19539);
nor U19869 (N_19869,N_19520,N_19699);
nand U19870 (N_19870,N_19637,N_19662);
or U19871 (N_19871,N_19546,N_19717);
nand U19872 (N_19872,N_19553,N_19741);
or U19873 (N_19873,N_19607,N_19650);
nor U19874 (N_19874,N_19530,N_19591);
and U19875 (N_19875,N_19733,N_19746);
and U19876 (N_19876,N_19638,N_19719);
nor U19877 (N_19877,N_19610,N_19550);
nor U19878 (N_19878,N_19711,N_19652);
nand U19879 (N_19879,N_19708,N_19620);
nor U19880 (N_19880,N_19594,N_19687);
and U19881 (N_19881,N_19665,N_19522);
nand U19882 (N_19882,N_19667,N_19614);
and U19883 (N_19883,N_19570,N_19715);
or U19884 (N_19884,N_19697,N_19620);
or U19885 (N_19885,N_19531,N_19693);
and U19886 (N_19886,N_19578,N_19739);
nor U19887 (N_19887,N_19584,N_19510);
and U19888 (N_19888,N_19636,N_19598);
or U19889 (N_19889,N_19540,N_19583);
or U19890 (N_19890,N_19723,N_19700);
and U19891 (N_19891,N_19732,N_19505);
or U19892 (N_19892,N_19552,N_19536);
and U19893 (N_19893,N_19564,N_19722);
nor U19894 (N_19894,N_19558,N_19660);
or U19895 (N_19895,N_19545,N_19634);
nand U19896 (N_19896,N_19586,N_19654);
or U19897 (N_19897,N_19704,N_19594);
and U19898 (N_19898,N_19651,N_19652);
nor U19899 (N_19899,N_19658,N_19657);
and U19900 (N_19900,N_19588,N_19613);
nand U19901 (N_19901,N_19612,N_19662);
or U19902 (N_19902,N_19713,N_19611);
or U19903 (N_19903,N_19712,N_19686);
and U19904 (N_19904,N_19672,N_19617);
and U19905 (N_19905,N_19748,N_19539);
or U19906 (N_19906,N_19563,N_19690);
nand U19907 (N_19907,N_19594,N_19729);
and U19908 (N_19908,N_19588,N_19653);
and U19909 (N_19909,N_19630,N_19715);
or U19910 (N_19910,N_19609,N_19522);
or U19911 (N_19911,N_19529,N_19574);
or U19912 (N_19912,N_19743,N_19593);
nor U19913 (N_19913,N_19718,N_19505);
or U19914 (N_19914,N_19510,N_19518);
nor U19915 (N_19915,N_19512,N_19617);
nand U19916 (N_19916,N_19621,N_19525);
and U19917 (N_19917,N_19674,N_19515);
or U19918 (N_19918,N_19743,N_19575);
nand U19919 (N_19919,N_19686,N_19504);
nand U19920 (N_19920,N_19573,N_19516);
and U19921 (N_19921,N_19668,N_19587);
and U19922 (N_19922,N_19637,N_19547);
or U19923 (N_19923,N_19640,N_19694);
or U19924 (N_19924,N_19728,N_19685);
nand U19925 (N_19925,N_19533,N_19581);
nand U19926 (N_19926,N_19609,N_19737);
nand U19927 (N_19927,N_19620,N_19675);
and U19928 (N_19928,N_19514,N_19740);
nand U19929 (N_19929,N_19608,N_19557);
or U19930 (N_19930,N_19649,N_19575);
nor U19931 (N_19931,N_19639,N_19636);
nand U19932 (N_19932,N_19597,N_19612);
nand U19933 (N_19933,N_19654,N_19557);
nand U19934 (N_19934,N_19583,N_19684);
nand U19935 (N_19935,N_19604,N_19513);
nor U19936 (N_19936,N_19646,N_19576);
nand U19937 (N_19937,N_19742,N_19662);
nand U19938 (N_19938,N_19613,N_19745);
xnor U19939 (N_19939,N_19738,N_19733);
and U19940 (N_19940,N_19603,N_19577);
nand U19941 (N_19941,N_19649,N_19670);
or U19942 (N_19942,N_19710,N_19664);
or U19943 (N_19943,N_19677,N_19605);
nand U19944 (N_19944,N_19698,N_19719);
and U19945 (N_19945,N_19543,N_19630);
nor U19946 (N_19946,N_19615,N_19541);
and U19947 (N_19947,N_19659,N_19610);
nand U19948 (N_19948,N_19542,N_19624);
or U19949 (N_19949,N_19698,N_19557);
or U19950 (N_19950,N_19648,N_19655);
and U19951 (N_19951,N_19632,N_19593);
and U19952 (N_19952,N_19562,N_19680);
nor U19953 (N_19953,N_19682,N_19629);
nand U19954 (N_19954,N_19691,N_19737);
and U19955 (N_19955,N_19584,N_19722);
or U19956 (N_19956,N_19739,N_19723);
and U19957 (N_19957,N_19638,N_19669);
and U19958 (N_19958,N_19635,N_19644);
nand U19959 (N_19959,N_19562,N_19665);
and U19960 (N_19960,N_19680,N_19732);
nor U19961 (N_19961,N_19566,N_19729);
and U19962 (N_19962,N_19524,N_19677);
nor U19963 (N_19963,N_19740,N_19676);
or U19964 (N_19964,N_19693,N_19666);
or U19965 (N_19965,N_19674,N_19724);
and U19966 (N_19966,N_19500,N_19715);
nand U19967 (N_19967,N_19585,N_19746);
or U19968 (N_19968,N_19629,N_19650);
nor U19969 (N_19969,N_19530,N_19547);
and U19970 (N_19970,N_19576,N_19745);
or U19971 (N_19971,N_19610,N_19726);
nand U19972 (N_19972,N_19737,N_19731);
or U19973 (N_19973,N_19516,N_19515);
nand U19974 (N_19974,N_19735,N_19576);
or U19975 (N_19975,N_19726,N_19564);
and U19976 (N_19976,N_19729,N_19604);
nor U19977 (N_19977,N_19609,N_19521);
nand U19978 (N_19978,N_19500,N_19644);
or U19979 (N_19979,N_19575,N_19525);
and U19980 (N_19980,N_19615,N_19746);
or U19981 (N_19981,N_19657,N_19563);
nor U19982 (N_19982,N_19592,N_19653);
or U19983 (N_19983,N_19617,N_19628);
nor U19984 (N_19984,N_19706,N_19599);
nand U19985 (N_19985,N_19737,N_19522);
nor U19986 (N_19986,N_19531,N_19715);
or U19987 (N_19987,N_19614,N_19689);
or U19988 (N_19988,N_19709,N_19647);
or U19989 (N_19989,N_19667,N_19725);
nand U19990 (N_19990,N_19515,N_19534);
xor U19991 (N_19991,N_19501,N_19560);
or U19992 (N_19992,N_19523,N_19524);
nor U19993 (N_19993,N_19741,N_19599);
and U19994 (N_19994,N_19666,N_19555);
nor U19995 (N_19995,N_19617,N_19571);
nand U19996 (N_19996,N_19605,N_19505);
and U19997 (N_19997,N_19531,N_19625);
xor U19998 (N_19998,N_19536,N_19647);
nor U19999 (N_19999,N_19739,N_19548);
nand U20000 (N_20000,N_19838,N_19930);
or U20001 (N_20001,N_19886,N_19985);
nor U20002 (N_20002,N_19891,N_19879);
nor U20003 (N_20003,N_19860,N_19785);
nand U20004 (N_20004,N_19874,N_19866);
and U20005 (N_20005,N_19793,N_19924);
or U20006 (N_20006,N_19913,N_19825);
and U20007 (N_20007,N_19798,N_19871);
nand U20008 (N_20008,N_19966,N_19971);
nor U20009 (N_20009,N_19997,N_19963);
and U20010 (N_20010,N_19750,N_19852);
nand U20011 (N_20011,N_19814,N_19956);
and U20012 (N_20012,N_19780,N_19868);
nor U20013 (N_20013,N_19911,N_19802);
nand U20014 (N_20014,N_19948,N_19964);
and U20015 (N_20015,N_19828,N_19884);
and U20016 (N_20016,N_19861,N_19847);
or U20017 (N_20017,N_19781,N_19987);
xor U20018 (N_20018,N_19915,N_19899);
nand U20019 (N_20019,N_19933,N_19901);
nand U20020 (N_20020,N_19876,N_19819);
nand U20021 (N_20021,N_19863,N_19962);
or U20022 (N_20022,N_19976,N_19960);
nor U20023 (N_20023,N_19822,N_19751);
nand U20024 (N_20024,N_19829,N_19921);
and U20025 (N_20025,N_19978,N_19936);
nand U20026 (N_20026,N_19902,N_19790);
or U20027 (N_20027,N_19881,N_19835);
nor U20028 (N_20028,N_19854,N_19760);
and U20029 (N_20029,N_19767,N_19801);
xor U20030 (N_20030,N_19920,N_19875);
nand U20031 (N_20031,N_19817,N_19859);
and U20032 (N_20032,N_19955,N_19942);
nor U20033 (N_20033,N_19969,N_19952);
and U20034 (N_20034,N_19990,N_19912);
or U20035 (N_20035,N_19797,N_19914);
and U20036 (N_20036,N_19944,N_19792);
nor U20037 (N_20037,N_19853,N_19977);
nor U20038 (N_20038,N_19938,N_19771);
or U20039 (N_20039,N_19768,N_19851);
nand U20040 (N_20040,N_19959,N_19783);
nor U20041 (N_20041,N_19919,N_19928);
and U20042 (N_20042,N_19756,N_19775);
nor U20043 (N_20043,N_19947,N_19981);
nor U20044 (N_20044,N_19968,N_19848);
and U20045 (N_20045,N_19776,N_19823);
and U20046 (N_20046,N_19856,N_19800);
and U20047 (N_20047,N_19777,N_19791);
nor U20048 (N_20048,N_19937,N_19932);
and U20049 (N_20049,N_19984,N_19845);
nor U20050 (N_20050,N_19880,N_19784);
nor U20051 (N_20051,N_19870,N_19894);
nor U20052 (N_20052,N_19909,N_19773);
or U20053 (N_20053,N_19973,N_19951);
or U20054 (N_20054,N_19795,N_19809);
nor U20055 (N_20055,N_19935,N_19883);
nand U20056 (N_20056,N_19769,N_19831);
or U20057 (N_20057,N_19830,N_19862);
nor U20058 (N_20058,N_19806,N_19839);
nor U20059 (N_20059,N_19836,N_19910);
nand U20060 (N_20060,N_19872,N_19762);
and U20061 (N_20061,N_19855,N_19957);
nand U20062 (N_20062,N_19753,N_19953);
nand U20063 (N_20063,N_19820,N_19869);
nand U20064 (N_20064,N_19898,N_19908);
or U20065 (N_20065,N_19815,N_19844);
and U20066 (N_20066,N_19788,N_19810);
nand U20067 (N_20067,N_19755,N_19865);
and U20068 (N_20068,N_19807,N_19922);
and U20069 (N_20069,N_19885,N_19877);
or U20070 (N_20070,N_19940,N_19967);
or U20071 (N_20071,N_19989,N_19918);
nor U20072 (N_20072,N_19794,N_19905);
and U20073 (N_20073,N_19778,N_19980);
nor U20074 (N_20074,N_19782,N_19988);
nor U20075 (N_20075,N_19974,N_19816);
or U20076 (N_20076,N_19850,N_19811);
nor U20077 (N_20077,N_19934,N_19796);
or U20078 (N_20078,N_19846,N_19943);
nor U20079 (N_20079,N_19900,N_19907);
or U20080 (N_20080,N_19925,N_19995);
and U20081 (N_20081,N_19896,N_19906);
nand U20082 (N_20082,N_19849,N_19808);
nand U20083 (N_20083,N_19897,N_19895);
and U20084 (N_20084,N_19917,N_19824);
or U20085 (N_20085,N_19818,N_19758);
nor U20086 (N_20086,N_19950,N_19982);
nor U20087 (N_20087,N_19949,N_19946);
or U20088 (N_20088,N_19993,N_19764);
or U20089 (N_20089,N_19770,N_19821);
and U20090 (N_20090,N_19941,N_19961);
and U20091 (N_20091,N_19787,N_19858);
or U20092 (N_20092,N_19834,N_19892);
or U20093 (N_20093,N_19752,N_19867);
or U20094 (N_20094,N_19903,N_19888);
nand U20095 (N_20095,N_19893,N_19887);
or U20096 (N_20096,N_19843,N_19999);
nor U20097 (N_20097,N_19970,N_19842);
nor U20098 (N_20098,N_19972,N_19983);
nand U20099 (N_20099,N_19841,N_19904);
nand U20100 (N_20100,N_19805,N_19786);
nor U20101 (N_20101,N_19890,N_19763);
and U20102 (N_20102,N_19864,N_19926);
nor U20103 (N_20103,N_19878,N_19833);
and U20104 (N_20104,N_19931,N_19799);
and U20105 (N_20105,N_19772,N_19827);
and U20106 (N_20106,N_19826,N_19992);
nand U20107 (N_20107,N_19857,N_19837);
nand U20108 (N_20108,N_19998,N_19916);
or U20109 (N_20109,N_19804,N_19975);
nor U20110 (N_20110,N_19832,N_19803);
nand U20111 (N_20111,N_19929,N_19939);
nand U20112 (N_20112,N_19927,N_19986);
nand U20113 (N_20113,N_19757,N_19954);
and U20114 (N_20114,N_19761,N_19754);
or U20115 (N_20115,N_19774,N_19889);
nand U20116 (N_20116,N_19979,N_19812);
nor U20117 (N_20117,N_19840,N_19965);
and U20118 (N_20118,N_19766,N_19996);
nor U20119 (N_20119,N_19759,N_19991);
and U20120 (N_20120,N_19923,N_19789);
and U20121 (N_20121,N_19873,N_19779);
nor U20122 (N_20122,N_19958,N_19882);
nor U20123 (N_20123,N_19765,N_19945);
nand U20124 (N_20124,N_19813,N_19994);
or U20125 (N_20125,N_19841,N_19957);
nor U20126 (N_20126,N_19811,N_19777);
and U20127 (N_20127,N_19927,N_19930);
nor U20128 (N_20128,N_19946,N_19772);
nor U20129 (N_20129,N_19794,N_19785);
or U20130 (N_20130,N_19980,N_19767);
nor U20131 (N_20131,N_19824,N_19989);
nor U20132 (N_20132,N_19972,N_19958);
or U20133 (N_20133,N_19832,N_19807);
or U20134 (N_20134,N_19849,N_19817);
or U20135 (N_20135,N_19932,N_19854);
nor U20136 (N_20136,N_19830,N_19857);
and U20137 (N_20137,N_19973,N_19800);
and U20138 (N_20138,N_19826,N_19871);
nor U20139 (N_20139,N_19919,N_19965);
nand U20140 (N_20140,N_19763,N_19971);
or U20141 (N_20141,N_19885,N_19996);
or U20142 (N_20142,N_19778,N_19865);
or U20143 (N_20143,N_19830,N_19979);
or U20144 (N_20144,N_19983,N_19804);
and U20145 (N_20145,N_19923,N_19802);
and U20146 (N_20146,N_19768,N_19904);
xor U20147 (N_20147,N_19823,N_19986);
nor U20148 (N_20148,N_19831,N_19943);
nor U20149 (N_20149,N_19760,N_19940);
and U20150 (N_20150,N_19765,N_19750);
nand U20151 (N_20151,N_19855,N_19975);
or U20152 (N_20152,N_19940,N_19898);
nand U20153 (N_20153,N_19840,N_19767);
nor U20154 (N_20154,N_19764,N_19955);
and U20155 (N_20155,N_19781,N_19970);
nand U20156 (N_20156,N_19937,N_19901);
nor U20157 (N_20157,N_19914,N_19824);
and U20158 (N_20158,N_19901,N_19979);
nand U20159 (N_20159,N_19891,N_19845);
nand U20160 (N_20160,N_19818,N_19868);
nor U20161 (N_20161,N_19943,N_19991);
nand U20162 (N_20162,N_19999,N_19781);
and U20163 (N_20163,N_19997,N_19857);
or U20164 (N_20164,N_19861,N_19990);
nor U20165 (N_20165,N_19931,N_19906);
and U20166 (N_20166,N_19955,N_19919);
or U20167 (N_20167,N_19948,N_19876);
or U20168 (N_20168,N_19988,N_19999);
and U20169 (N_20169,N_19798,N_19982);
nor U20170 (N_20170,N_19751,N_19936);
nor U20171 (N_20171,N_19838,N_19962);
nand U20172 (N_20172,N_19824,N_19780);
nand U20173 (N_20173,N_19977,N_19835);
and U20174 (N_20174,N_19873,N_19776);
xnor U20175 (N_20175,N_19784,N_19860);
xor U20176 (N_20176,N_19818,N_19776);
or U20177 (N_20177,N_19912,N_19833);
xnor U20178 (N_20178,N_19781,N_19788);
nand U20179 (N_20179,N_19760,N_19927);
or U20180 (N_20180,N_19960,N_19977);
nand U20181 (N_20181,N_19839,N_19857);
nand U20182 (N_20182,N_19768,N_19796);
nand U20183 (N_20183,N_19895,N_19964);
nor U20184 (N_20184,N_19949,N_19842);
nor U20185 (N_20185,N_19937,N_19849);
or U20186 (N_20186,N_19772,N_19826);
and U20187 (N_20187,N_19874,N_19924);
or U20188 (N_20188,N_19855,N_19832);
nand U20189 (N_20189,N_19777,N_19993);
nand U20190 (N_20190,N_19984,N_19755);
and U20191 (N_20191,N_19843,N_19798);
or U20192 (N_20192,N_19851,N_19849);
nand U20193 (N_20193,N_19884,N_19914);
and U20194 (N_20194,N_19937,N_19813);
nand U20195 (N_20195,N_19864,N_19928);
or U20196 (N_20196,N_19886,N_19989);
or U20197 (N_20197,N_19906,N_19886);
or U20198 (N_20198,N_19827,N_19879);
nor U20199 (N_20199,N_19860,N_19870);
nor U20200 (N_20200,N_19936,N_19790);
and U20201 (N_20201,N_19785,N_19955);
or U20202 (N_20202,N_19971,N_19838);
nand U20203 (N_20203,N_19996,N_19974);
nor U20204 (N_20204,N_19904,N_19903);
nand U20205 (N_20205,N_19880,N_19937);
and U20206 (N_20206,N_19778,N_19983);
and U20207 (N_20207,N_19965,N_19949);
and U20208 (N_20208,N_19856,N_19812);
nand U20209 (N_20209,N_19898,N_19770);
nor U20210 (N_20210,N_19918,N_19928);
or U20211 (N_20211,N_19887,N_19945);
or U20212 (N_20212,N_19805,N_19897);
or U20213 (N_20213,N_19935,N_19901);
or U20214 (N_20214,N_19837,N_19912);
nand U20215 (N_20215,N_19826,N_19762);
nand U20216 (N_20216,N_19872,N_19873);
and U20217 (N_20217,N_19815,N_19872);
nor U20218 (N_20218,N_19944,N_19764);
nand U20219 (N_20219,N_19867,N_19799);
or U20220 (N_20220,N_19943,N_19916);
nor U20221 (N_20221,N_19979,N_19986);
nand U20222 (N_20222,N_19833,N_19889);
or U20223 (N_20223,N_19869,N_19922);
nor U20224 (N_20224,N_19833,N_19916);
nor U20225 (N_20225,N_19798,N_19779);
nand U20226 (N_20226,N_19973,N_19888);
nand U20227 (N_20227,N_19899,N_19963);
or U20228 (N_20228,N_19897,N_19788);
nor U20229 (N_20229,N_19949,N_19862);
and U20230 (N_20230,N_19777,N_19770);
and U20231 (N_20231,N_19909,N_19817);
nand U20232 (N_20232,N_19850,N_19757);
nand U20233 (N_20233,N_19841,N_19839);
and U20234 (N_20234,N_19850,N_19986);
or U20235 (N_20235,N_19868,N_19907);
nand U20236 (N_20236,N_19825,N_19927);
or U20237 (N_20237,N_19988,N_19792);
and U20238 (N_20238,N_19828,N_19996);
and U20239 (N_20239,N_19760,N_19845);
and U20240 (N_20240,N_19835,N_19933);
nand U20241 (N_20241,N_19828,N_19881);
nand U20242 (N_20242,N_19978,N_19895);
nor U20243 (N_20243,N_19826,N_19874);
nor U20244 (N_20244,N_19959,N_19876);
or U20245 (N_20245,N_19806,N_19879);
xnor U20246 (N_20246,N_19917,N_19940);
nand U20247 (N_20247,N_19964,N_19886);
nor U20248 (N_20248,N_19887,N_19787);
nand U20249 (N_20249,N_19869,N_19843);
or U20250 (N_20250,N_20182,N_20129);
and U20251 (N_20251,N_20221,N_20151);
nor U20252 (N_20252,N_20010,N_20077);
and U20253 (N_20253,N_20229,N_20216);
nand U20254 (N_20254,N_20237,N_20206);
and U20255 (N_20255,N_20018,N_20139);
nand U20256 (N_20256,N_20224,N_20164);
nand U20257 (N_20257,N_20191,N_20054);
or U20258 (N_20258,N_20176,N_20154);
or U20259 (N_20259,N_20080,N_20050);
nand U20260 (N_20260,N_20005,N_20003);
and U20261 (N_20261,N_20170,N_20214);
or U20262 (N_20262,N_20231,N_20060);
nor U20263 (N_20263,N_20022,N_20245);
nand U20264 (N_20264,N_20135,N_20081);
nor U20265 (N_20265,N_20033,N_20131);
nand U20266 (N_20266,N_20194,N_20123);
nand U20267 (N_20267,N_20052,N_20101);
and U20268 (N_20268,N_20041,N_20169);
nand U20269 (N_20269,N_20161,N_20198);
nand U20270 (N_20270,N_20115,N_20248);
nand U20271 (N_20271,N_20099,N_20104);
or U20272 (N_20272,N_20053,N_20177);
nor U20273 (N_20273,N_20044,N_20166);
or U20274 (N_20274,N_20049,N_20227);
nor U20275 (N_20275,N_20056,N_20094);
nand U20276 (N_20276,N_20186,N_20168);
and U20277 (N_20277,N_20174,N_20090);
or U20278 (N_20278,N_20061,N_20238);
nor U20279 (N_20279,N_20069,N_20037);
nor U20280 (N_20280,N_20178,N_20163);
nor U20281 (N_20281,N_20014,N_20149);
and U20282 (N_20282,N_20035,N_20147);
nand U20283 (N_20283,N_20046,N_20109);
nand U20284 (N_20284,N_20218,N_20140);
nor U20285 (N_20285,N_20235,N_20097);
nor U20286 (N_20286,N_20153,N_20181);
or U20287 (N_20287,N_20084,N_20193);
nand U20288 (N_20288,N_20088,N_20212);
nand U20289 (N_20289,N_20152,N_20211);
and U20290 (N_20290,N_20171,N_20236);
nor U20291 (N_20291,N_20209,N_20007);
nor U20292 (N_20292,N_20015,N_20102);
and U20293 (N_20293,N_20136,N_20145);
nor U20294 (N_20294,N_20200,N_20133);
nor U20295 (N_20295,N_20043,N_20141);
nand U20296 (N_20296,N_20073,N_20100);
nand U20297 (N_20297,N_20012,N_20172);
nor U20298 (N_20298,N_20042,N_20219);
nand U20299 (N_20299,N_20086,N_20112);
or U20300 (N_20300,N_20091,N_20239);
and U20301 (N_20301,N_20114,N_20000);
or U20302 (N_20302,N_20232,N_20160);
and U20303 (N_20303,N_20197,N_20165);
or U20304 (N_20304,N_20247,N_20184);
or U20305 (N_20305,N_20233,N_20026);
and U20306 (N_20306,N_20064,N_20024);
nor U20307 (N_20307,N_20029,N_20196);
nand U20308 (N_20308,N_20220,N_20120);
or U20309 (N_20309,N_20116,N_20199);
and U20310 (N_20310,N_20208,N_20040);
nor U20311 (N_20311,N_20021,N_20180);
nand U20312 (N_20312,N_20002,N_20070);
nand U20313 (N_20313,N_20083,N_20051);
nand U20314 (N_20314,N_20106,N_20078);
or U20315 (N_20315,N_20144,N_20118);
nor U20316 (N_20316,N_20074,N_20187);
nand U20317 (N_20317,N_20119,N_20110);
and U20318 (N_20318,N_20215,N_20242);
nand U20319 (N_20319,N_20016,N_20201);
or U20320 (N_20320,N_20210,N_20143);
and U20321 (N_20321,N_20146,N_20167);
and U20322 (N_20322,N_20020,N_20223);
and U20323 (N_20323,N_20013,N_20008);
and U20324 (N_20324,N_20138,N_20059);
nor U20325 (N_20325,N_20028,N_20096);
nand U20326 (N_20326,N_20103,N_20023);
or U20327 (N_20327,N_20063,N_20241);
or U20328 (N_20328,N_20189,N_20132);
nor U20329 (N_20329,N_20039,N_20019);
nor U20330 (N_20330,N_20017,N_20038);
and U20331 (N_20331,N_20148,N_20113);
nor U20332 (N_20332,N_20072,N_20156);
nor U20333 (N_20333,N_20213,N_20031);
and U20334 (N_20334,N_20195,N_20190);
or U20335 (N_20335,N_20157,N_20062);
nand U20336 (N_20336,N_20142,N_20107);
nor U20337 (N_20337,N_20048,N_20082);
xnor U20338 (N_20338,N_20126,N_20202);
or U20339 (N_20339,N_20246,N_20068);
and U20340 (N_20340,N_20205,N_20192);
and U20341 (N_20341,N_20032,N_20226);
and U20342 (N_20342,N_20240,N_20111);
nor U20343 (N_20343,N_20127,N_20225);
and U20344 (N_20344,N_20159,N_20222);
nand U20345 (N_20345,N_20004,N_20089);
or U20346 (N_20346,N_20066,N_20030);
and U20347 (N_20347,N_20117,N_20175);
nand U20348 (N_20348,N_20230,N_20057);
nand U20349 (N_20349,N_20155,N_20093);
or U20350 (N_20350,N_20085,N_20036);
nand U20351 (N_20351,N_20158,N_20121);
nand U20352 (N_20352,N_20034,N_20025);
nand U20353 (N_20353,N_20228,N_20130);
nand U20354 (N_20354,N_20150,N_20011);
nand U20355 (N_20355,N_20217,N_20162);
nand U20356 (N_20356,N_20058,N_20179);
nor U20357 (N_20357,N_20045,N_20108);
and U20358 (N_20358,N_20128,N_20087);
and U20359 (N_20359,N_20009,N_20067);
nand U20360 (N_20360,N_20001,N_20185);
or U20361 (N_20361,N_20098,N_20075);
nor U20362 (N_20362,N_20125,N_20065);
nor U20363 (N_20363,N_20234,N_20183);
or U20364 (N_20364,N_20071,N_20124);
and U20365 (N_20365,N_20095,N_20173);
nor U20366 (N_20366,N_20244,N_20207);
nand U20367 (N_20367,N_20092,N_20134);
or U20368 (N_20368,N_20027,N_20243);
and U20369 (N_20369,N_20122,N_20203);
nand U20370 (N_20370,N_20055,N_20047);
nand U20371 (N_20371,N_20204,N_20188);
and U20372 (N_20372,N_20249,N_20006);
or U20373 (N_20373,N_20137,N_20079);
or U20374 (N_20374,N_20105,N_20076);
and U20375 (N_20375,N_20029,N_20220);
nand U20376 (N_20376,N_20156,N_20041);
or U20377 (N_20377,N_20236,N_20005);
nor U20378 (N_20378,N_20097,N_20201);
or U20379 (N_20379,N_20009,N_20111);
nor U20380 (N_20380,N_20065,N_20202);
nand U20381 (N_20381,N_20142,N_20055);
or U20382 (N_20382,N_20078,N_20151);
and U20383 (N_20383,N_20127,N_20222);
nand U20384 (N_20384,N_20113,N_20242);
and U20385 (N_20385,N_20078,N_20100);
nand U20386 (N_20386,N_20150,N_20246);
nor U20387 (N_20387,N_20140,N_20000);
nor U20388 (N_20388,N_20163,N_20079);
or U20389 (N_20389,N_20239,N_20092);
or U20390 (N_20390,N_20183,N_20094);
xnor U20391 (N_20391,N_20105,N_20233);
nor U20392 (N_20392,N_20074,N_20189);
nand U20393 (N_20393,N_20163,N_20116);
or U20394 (N_20394,N_20070,N_20149);
and U20395 (N_20395,N_20215,N_20218);
nor U20396 (N_20396,N_20039,N_20034);
nand U20397 (N_20397,N_20102,N_20082);
nand U20398 (N_20398,N_20033,N_20172);
or U20399 (N_20399,N_20029,N_20225);
nor U20400 (N_20400,N_20220,N_20231);
nor U20401 (N_20401,N_20200,N_20130);
or U20402 (N_20402,N_20001,N_20019);
nor U20403 (N_20403,N_20049,N_20246);
nand U20404 (N_20404,N_20121,N_20008);
nor U20405 (N_20405,N_20148,N_20025);
and U20406 (N_20406,N_20161,N_20061);
nand U20407 (N_20407,N_20081,N_20141);
nand U20408 (N_20408,N_20011,N_20116);
or U20409 (N_20409,N_20109,N_20099);
nor U20410 (N_20410,N_20042,N_20176);
and U20411 (N_20411,N_20071,N_20002);
and U20412 (N_20412,N_20123,N_20122);
or U20413 (N_20413,N_20026,N_20137);
and U20414 (N_20414,N_20207,N_20194);
and U20415 (N_20415,N_20224,N_20248);
nor U20416 (N_20416,N_20099,N_20001);
or U20417 (N_20417,N_20151,N_20234);
or U20418 (N_20418,N_20151,N_20071);
nand U20419 (N_20419,N_20044,N_20178);
nor U20420 (N_20420,N_20139,N_20091);
nor U20421 (N_20421,N_20090,N_20088);
and U20422 (N_20422,N_20103,N_20136);
and U20423 (N_20423,N_20219,N_20203);
nor U20424 (N_20424,N_20200,N_20153);
nor U20425 (N_20425,N_20078,N_20072);
nor U20426 (N_20426,N_20110,N_20240);
nor U20427 (N_20427,N_20168,N_20092);
or U20428 (N_20428,N_20116,N_20210);
nor U20429 (N_20429,N_20121,N_20043);
nor U20430 (N_20430,N_20172,N_20206);
and U20431 (N_20431,N_20245,N_20186);
or U20432 (N_20432,N_20020,N_20141);
nor U20433 (N_20433,N_20051,N_20150);
and U20434 (N_20434,N_20079,N_20034);
and U20435 (N_20435,N_20215,N_20237);
and U20436 (N_20436,N_20132,N_20175);
or U20437 (N_20437,N_20161,N_20047);
nor U20438 (N_20438,N_20215,N_20049);
or U20439 (N_20439,N_20074,N_20218);
and U20440 (N_20440,N_20162,N_20070);
or U20441 (N_20441,N_20249,N_20038);
nor U20442 (N_20442,N_20024,N_20109);
nor U20443 (N_20443,N_20018,N_20085);
and U20444 (N_20444,N_20092,N_20034);
and U20445 (N_20445,N_20147,N_20125);
nand U20446 (N_20446,N_20107,N_20191);
and U20447 (N_20447,N_20158,N_20162);
nor U20448 (N_20448,N_20043,N_20184);
and U20449 (N_20449,N_20006,N_20155);
or U20450 (N_20450,N_20127,N_20004);
and U20451 (N_20451,N_20241,N_20179);
nor U20452 (N_20452,N_20191,N_20189);
nor U20453 (N_20453,N_20044,N_20084);
and U20454 (N_20454,N_20038,N_20016);
and U20455 (N_20455,N_20215,N_20090);
and U20456 (N_20456,N_20228,N_20019);
nor U20457 (N_20457,N_20037,N_20181);
or U20458 (N_20458,N_20064,N_20074);
nor U20459 (N_20459,N_20154,N_20053);
or U20460 (N_20460,N_20174,N_20168);
nand U20461 (N_20461,N_20087,N_20002);
or U20462 (N_20462,N_20096,N_20071);
and U20463 (N_20463,N_20238,N_20173);
nor U20464 (N_20464,N_20174,N_20037);
and U20465 (N_20465,N_20206,N_20238);
or U20466 (N_20466,N_20139,N_20033);
xnor U20467 (N_20467,N_20137,N_20213);
or U20468 (N_20468,N_20004,N_20126);
nor U20469 (N_20469,N_20064,N_20098);
and U20470 (N_20470,N_20113,N_20003);
nor U20471 (N_20471,N_20234,N_20094);
and U20472 (N_20472,N_20036,N_20242);
nor U20473 (N_20473,N_20121,N_20159);
nand U20474 (N_20474,N_20197,N_20208);
and U20475 (N_20475,N_20115,N_20151);
or U20476 (N_20476,N_20202,N_20109);
or U20477 (N_20477,N_20018,N_20095);
and U20478 (N_20478,N_20004,N_20002);
and U20479 (N_20479,N_20169,N_20023);
and U20480 (N_20480,N_20156,N_20048);
and U20481 (N_20481,N_20024,N_20077);
nand U20482 (N_20482,N_20138,N_20033);
or U20483 (N_20483,N_20143,N_20174);
and U20484 (N_20484,N_20033,N_20185);
nor U20485 (N_20485,N_20222,N_20058);
and U20486 (N_20486,N_20235,N_20020);
nand U20487 (N_20487,N_20221,N_20013);
or U20488 (N_20488,N_20069,N_20115);
nand U20489 (N_20489,N_20089,N_20061);
and U20490 (N_20490,N_20003,N_20051);
nor U20491 (N_20491,N_20192,N_20050);
or U20492 (N_20492,N_20091,N_20071);
nand U20493 (N_20493,N_20175,N_20231);
or U20494 (N_20494,N_20078,N_20016);
or U20495 (N_20495,N_20180,N_20025);
and U20496 (N_20496,N_20151,N_20100);
and U20497 (N_20497,N_20236,N_20168);
nand U20498 (N_20498,N_20115,N_20243);
or U20499 (N_20499,N_20050,N_20029);
or U20500 (N_20500,N_20448,N_20413);
xnor U20501 (N_20501,N_20287,N_20252);
and U20502 (N_20502,N_20317,N_20495);
or U20503 (N_20503,N_20302,N_20262);
nor U20504 (N_20504,N_20292,N_20488);
nand U20505 (N_20505,N_20473,N_20293);
or U20506 (N_20506,N_20264,N_20390);
or U20507 (N_20507,N_20394,N_20297);
and U20508 (N_20508,N_20340,N_20274);
nand U20509 (N_20509,N_20385,N_20463);
and U20510 (N_20510,N_20343,N_20439);
and U20511 (N_20511,N_20377,N_20408);
or U20512 (N_20512,N_20373,N_20357);
nand U20513 (N_20513,N_20458,N_20254);
nor U20514 (N_20514,N_20266,N_20371);
and U20515 (N_20515,N_20349,N_20367);
and U20516 (N_20516,N_20376,N_20393);
nor U20517 (N_20517,N_20299,N_20291);
xnor U20518 (N_20518,N_20354,N_20263);
and U20519 (N_20519,N_20432,N_20479);
nor U20520 (N_20520,N_20335,N_20279);
or U20521 (N_20521,N_20267,N_20350);
or U20522 (N_20522,N_20417,N_20484);
nand U20523 (N_20523,N_20325,N_20273);
nor U20524 (N_20524,N_20490,N_20326);
and U20525 (N_20525,N_20375,N_20486);
nand U20526 (N_20526,N_20482,N_20380);
and U20527 (N_20527,N_20301,N_20277);
or U20528 (N_20528,N_20281,N_20269);
and U20529 (N_20529,N_20427,N_20493);
nand U20530 (N_20530,N_20285,N_20461);
or U20531 (N_20531,N_20494,N_20328);
or U20532 (N_20532,N_20419,N_20289);
nor U20533 (N_20533,N_20497,N_20383);
or U20534 (N_20534,N_20369,N_20341);
and U20535 (N_20535,N_20405,N_20446);
or U20536 (N_20536,N_20378,N_20467);
or U20537 (N_20537,N_20403,N_20499);
nor U20538 (N_20538,N_20401,N_20331);
and U20539 (N_20539,N_20434,N_20351);
nor U20540 (N_20540,N_20455,N_20443);
or U20541 (N_20541,N_20409,N_20352);
nand U20542 (N_20542,N_20290,N_20339);
nor U20543 (N_20543,N_20337,N_20433);
or U20544 (N_20544,N_20253,N_20276);
nor U20545 (N_20545,N_20363,N_20338);
or U20546 (N_20546,N_20321,N_20355);
nor U20547 (N_20547,N_20307,N_20345);
nand U20548 (N_20548,N_20300,N_20422);
nor U20549 (N_20549,N_20392,N_20360);
or U20550 (N_20550,N_20358,N_20362);
or U20551 (N_20551,N_20415,N_20283);
nor U20552 (N_20552,N_20381,N_20462);
and U20553 (N_20553,N_20284,N_20323);
and U20554 (N_20554,N_20332,N_20318);
nand U20555 (N_20555,N_20436,N_20478);
nand U20556 (N_20556,N_20327,N_20399);
or U20557 (N_20557,N_20344,N_20426);
nor U20558 (N_20558,N_20372,N_20465);
or U20559 (N_20559,N_20334,N_20464);
or U20560 (N_20560,N_20275,N_20388);
or U20561 (N_20561,N_20305,N_20472);
nor U20562 (N_20562,N_20389,N_20485);
nor U20563 (N_20563,N_20286,N_20410);
nand U20564 (N_20564,N_20402,N_20368);
nor U20565 (N_20565,N_20260,N_20476);
and U20566 (N_20566,N_20329,N_20498);
nand U20567 (N_20567,N_20456,N_20333);
and U20568 (N_20568,N_20404,N_20310);
nor U20569 (N_20569,N_20441,N_20431);
or U20570 (N_20570,N_20353,N_20312);
nor U20571 (N_20571,N_20255,N_20480);
nor U20572 (N_20572,N_20425,N_20356);
or U20573 (N_20573,N_20492,N_20481);
or U20574 (N_20574,N_20469,N_20280);
or U20575 (N_20575,N_20282,N_20272);
or U20576 (N_20576,N_20347,N_20454);
nand U20577 (N_20577,N_20396,N_20459);
nand U20578 (N_20578,N_20346,N_20361);
or U20579 (N_20579,N_20270,N_20364);
or U20580 (N_20580,N_20430,N_20314);
nand U20581 (N_20581,N_20421,N_20444);
nor U20582 (N_20582,N_20295,N_20489);
or U20583 (N_20583,N_20429,N_20397);
nor U20584 (N_20584,N_20437,N_20445);
nand U20585 (N_20585,N_20496,N_20453);
nand U20586 (N_20586,N_20251,N_20250);
or U20587 (N_20587,N_20424,N_20450);
or U20588 (N_20588,N_20370,N_20483);
or U20589 (N_20589,N_20395,N_20420);
or U20590 (N_20590,N_20412,N_20451);
or U20591 (N_20591,N_20468,N_20296);
nand U20592 (N_20592,N_20406,N_20442);
nand U20593 (N_20593,N_20475,N_20259);
or U20594 (N_20594,N_20379,N_20382);
or U20595 (N_20595,N_20306,N_20257);
nand U20596 (N_20596,N_20278,N_20391);
or U20597 (N_20597,N_20342,N_20400);
nor U20598 (N_20598,N_20319,N_20311);
nand U20599 (N_20599,N_20265,N_20271);
and U20600 (N_20600,N_20366,N_20298);
or U20601 (N_20601,N_20470,N_20438);
nor U20602 (N_20602,N_20309,N_20303);
and U20603 (N_20603,N_20418,N_20374);
and U20604 (N_20604,N_20474,N_20449);
or U20605 (N_20605,N_20471,N_20457);
nor U20606 (N_20606,N_20313,N_20466);
nand U20607 (N_20607,N_20435,N_20304);
or U20608 (N_20608,N_20411,N_20386);
or U20609 (N_20609,N_20407,N_20330);
nand U20610 (N_20610,N_20387,N_20315);
nand U20611 (N_20611,N_20428,N_20316);
or U20612 (N_20612,N_20261,N_20487);
nand U20613 (N_20613,N_20322,N_20256);
nor U20614 (N_20614,N_20336,N_20440);
or U20615 (N_20615,N_20452,N_20477);
nor U20616 (N_20616,N_20320,N_20324);
and U20617 (N_20617,N_20308,N_20268);
nor U20618 (N_20618,N_20348,N_20447);
or U20619 (N_20619,N_20414,N_20460);
nor U20620 (N_20620,N_20416,N_20384);
or U20621 (N_20621,N_20398,N_20365);
nand U20622 (N_20622,N_20491,N_20359);
nand U20623 (N_20623,N_20294,N_20423);
nand U20624 (N_20624,N_20258,N_20288);
xor U20625 (N_20625,N_20463,N_20256);
or U20626 (N_20626,N_20445,N_20460);
nor U20627 (N_20627,N_20427,N_20385);
xor U20628 (N_20628,N_20251,N_20495);
nand U20629 (N_20629,N_20272,N_20430);
nor U20630 (N_20630,N_20353,N_20442);
nand U20631 (N_20631,N_20468,N_20297);
and U20632 (N_20632,N_20415,N_20254);
nand U20633 (N_20633,N_20291,N_20315);
or U20634 (N_20634,N_20289,N_20276);
nor U20635 (N_20635,N_20348,N_20252);
and U20636 (N_20636,N_20353,N_20324);
nor U20637 (N_20637,N_20464,N_20406);
or U20638 (N_20638,N_20470,N_20493);
nor U20639 (N_20639,N_20496,N_20374);
and U20640 (N_20640,N_20415,N_20473);
and U20641 (N_20641,N_20441,N_20410);
and U20642 (N_20642,N_20285,N_20488);
and U20643 (N_20643,N_20312,N_20446);
nor U20644 (N_20644,N_20266,N_20280);
xnor U20645 (N_20645,N_20470,N_20439);
and U20646 (N_20646,N_20495,N_20270);
nand U20647 (N_20647,N_20456,N_20486);
or U20648 (N_20648,N_20424,N_20478);
nand U20649 (N_20649,N_20254,N_20409);
or U20650 (N_20650,N_20425,N_20348);
nand U20651 (N_20651,N_20263,N_20421);
nor U20652 (N_20652,N_20280,N_20394);
and U20653 (N_20653,N_20307,N_20319);
nand U20654 (N_20654,N_20476,N_20343);
nor U20655 (N_20655,N_20355,N_20258);
or U20656 (N_20656,N_20436,N_20453);
nor U20657 (N_20657,N_20250,N_20377);
and U20658 (N_20658,N_20359,N_20315);
or U20659 (N_20659,N_20262,N_20274);
nor U20660 (N_20660,N_20250,N_20422);
nand U20661 (N_20661,N_20446,N_20266);
nand U20662 (N_20662,N_20273,N_20277);
or U20663 (N_20663,N_20381,N_20383);
nand U20664 (N_20664,N_20390,N_20251);
nand U20665 (N_20665,N_20353,N_20345);
nor U20666 (N_20666,N_20330,N_20338);
or U20667 (N_20667,N_20304,N_20254);
or U20668 (N_20668,N_20419,N_20324);
nand U20669 (N_20669,N_20470,N_20311);
and U20670 (N_20670,N_20335,N_20492);
or U20671 (N_20671,N_20285,N_20485);
or U20672 (N_20672,N_20402,N_20473);
and U20673 (N_20673,N_20447,N_20290);
and U20674 (N_20674,N_20496,N_20293);
nor U20675 (N_20675,N_20341,N_20483);
nor U20676 (N_20676,N_20339,N_20457);
nor U20677 (N_20677,N_20466,N_20257);
or U20678 (N_20678,N_20284,N_20257);
and U20679 (N_20679,N_20419,N_20427);
or U20680 (N_20680,N_20442,N_20378);
or U20681 (N_20681,N_20463,N_20383);
and U20682 (N_20682,N_20398,N_20499);
nand U20683 (N_20683,N_20369,N_20264);
and U20684 (N_20684,N_20449,N_20423);
or U20685 (N_20685,N_20313,N_20250);
nand U20686 (N_20686,N_20447,N_20441);
nor U20687 (N_20687,N_20303,N_20473);
or U20688 (N_20688,N_20489,N_20442);
and U20689 (N_20689,N_20297,N_20303);
nand U20690 (N_20690,N_20483,N_20332);
nand U20691 (N_20691,N_20427,N_20338);
nor U20692 (N_20692,N_20337,N_20374);
or U20693 (N_20693,N_20304,N_20408);
nor U20694 (N_20694,N_20311,N_20349);
and U20695 (N_20695,N_20489,N_20356);
nand U20696 (N_20696,N_20429,N_20305);
or U20697 (N_20697,N_20356,N_20331);
nand U20698 (N_20698,N_20438,N_20257);
nor U20699 (N_20699,N_20352,N_20443);
nor U20700 (N_20700,N_20373,N_20465);
nor U20701 (N_20701,N_20408,N_20493);
nor U20702 (N_20702,N_20282,N_20269);
or U20703 (N_20703,N_20497,N_20498);
or U20704 (N_20704,N_20425,N_20476);
nor U20705 (N_20705,N_20302,N_20273);
nand U20706 (N_20706,N_20254,N_20298);
and U20707 (N_20707,N_20260,N_20251);
and U20708 (N_20708,N_20302,N_20360);
nand U20709 (N_20709,N_20403,N_20324);
nor U20710 (N_20710,N_20461,N_20259);
nand U20711 (N_20711,N_20407,N_20309);
nand U20712 (N_20712,N_20436,N_20373);
or U20713 (N_20713,N_20381,N_20496);
and U20714 (N_20714,N_20489,N_20388);
and U20715 (N_20715,N_20280,N_20483);
and U20716 (N_20716,N_20309,N_20251);
nand U20717 (N_20717,N_20453,N_20478);
and U20718 (N_20718,N_20398,N_20296);
nor U20719 (N_20719,N_20472,N_20357);
and U20720 (N_20720,N_20281,N_20277);
and U20721 (N_20721,N_20375,N_20277);
and U20722 (N_20722,N_20283,N_20277);
or U20723 (N_20723,N_20312,N_20391);
nor U20724 (N_20724,N_20374,N_20388);
nand U20725 (N_20725,N_20376,N_20395);
and U20726 (N_20726,N_20463,N_20488);
or U20727 (N_20727,N_20491,N_20345);
and U20728 (N_20728,N_20328,N_20287);
nand U20729 (N_20729,N_20298,N_20439);
or U20730 (N_20730,N_20277,N_20261);
nand U20731 (N_20731,N_20345,N_20405);
or U20732 (N_20732,N_20422,N_20384);
nand U20733 (N_20733,N_20490,N_20311);
or U20734 (N_20734,N_20435,N_20334);
nand U20735 (N_20735,N_20480,N_20436);
nor U20736 (N_20736,N_20290,N_20430);
nor U20737 (N_20737,N_20325,N_20338);
and U20738 (N_20738,N_20366,N_20275);
or U20739 (N_20739,N_20431,N_20429);
or U20740 (N_20740,N_20480,N_20334);
or U20741 (N_20741,N_20402,N_20288);
nand U20742 (N_20742,N_20294,N_20298);
nor U20743 (N_20743,N_20336,N_20479);
or U20744 (N_20744,N_20284,N_20390);
nand U20745 (N_20745,N_20388,N_20471);
nand U20746 (N_20746,N_20299,N_20439);
nor U20747 (N_20747,N_20395,N_20379);
nor U20748 (N_20748,N_20421,N_20362);
and U20749 (N_20749,N_20358,N_20336);
nand U20750 (N_20750,N_20742,N_20642);
or U20751 (N_20751,N_20622,N_20703);
and U20752 (N_20752,N_20508,N_20712);
and U20753 (N_20753,N_20546,N_20530);
nand U20754 (N_20754,N_20547,N_20625);
nor U20755 (N_20755,N_20554,N_20549);
and U20756 (N_20756,N_20569,N_20671);
and U20757 (N_20757,N_20567,N_20641);
nand U20758 (N_20758,N_20689,N_20679);
nand U20759 (N_20759,N_20714,N_20531);
nor U20760 (N_20760,N_20706,N_20621);
or U20761 (N_20761,N_20705,N_20609);
nand U20762 (N_20762,N_20558,N_20574);
and U20763 (N_20763,N_20675,N_20638);
or U20764 (N_20764,N_20583,N_20709);
or U20765 (N_20765,N_20749,N_20582);
and U20766 (N_20766,N_20686,N_20618);
or U20767 (N_20767,N_20735,N_20544);
nand U20768 (N_20768,N_20692,N_20639);
and U20769 (N_20769,N_20654,N_20718);
xnor U20770 (N_20770,N_20635,N_20651);
nand U20771 (N_20771,N_20726,N_20652);
and U20772 (N_20772,N_20595,N_20680);
and U20773 (N_20773,N_20528,N_20690);
and U20774 (N_20774,N_20503,N_20676);
nand U20775 (N_20775,N_20616,N_20725);
nor U20776 (N_20776,N_20716,N_20673);
or U20777 (N_20777,N_20516,N_20632);
nor U20778 (N_20778,N_20555,N_20536);
nand U20779 (N_20779,N_20643,N_20729);
nand U20780 (N_20780,N_20747,N_20738);
and U20781 (N_20781,N_20532,N_20501);
or U20782 (N_20782,N_20707,N_20548);
or U20783 (N_20783,N_20637,N_20540);
nand U20784 (N_20784,N_20698,N_20667);
or U20785 (N_20785,N_20745,N_20545);
nand U20786 (N_20786,N_20629,N_20526);
nor U20787 (N_20787,N_20513,N_20507);
nor U20788 (N_20788,N_20724,N_20727);
nor U20789 (N_20789,N_20552,N_20674);
nand U20790 (N_20790,N_20636,N_20500);
nor U20791 (N_20791,N_20693,N_20715);
or U20792 (N_20792,N_20743,N_20597);
nor U20793 (N_20793,N_20587,N_20506);
or U20794 (N_20794,N_20559,N_20653);
and U20795 (N_20795,N_20575,N_20691);
and U20796 (N_20796,N_20541,N_20662);
nand U20797 (N_20797,N_20576,N_20614);
or U20798 (N_20798,N_20739,N_20746);
and U20799 (N_20799,N_20599,N_20626);
and U20800 (N_20800,N_20631,N_20646);
nor U20801 (N_20801,N_20624,N_20577);
and U20802 (N_20802,N_20593,N_20570);
or U20803 (N_20803,N_20634,N_20700);
nor U20804 (N_20804,N_20717,N_20606);
or U20805 (N_20805,N_20610,N_20556);
nor U20806 (N_20806,N_20564,N_20603);
nand U20807 (N_20807,N_20578,N_20605);
and U20808 (N_20808,N_20627,N_20568);
nor U20809 (N_20809,N_20537,N_20645);
nor U20810 (N_20810,N_20542,N_20668);
or U20811 (N_20811,N_20663,N_20522);
nand U20812 (N_20812,N_20719,N_20511);
nor U20813 (N_20813,N_20509,N_20648);
nor U20814 (N_20814,N_20563,N_20685);
nand U20815 (N_20815,N_20551,N_20505);
or U20816 (N_20816,N_20702,N_20615);
nand U20817 (N_20817,N_20658,N_20670);
nand U20818 (N_20818,N_20561,N_20590);
nand U20819 (N_20819,N_20594,N_20666);
and U20820 (N_20820,N_20699,N_20741);
nor U20821 (N_20821,N_20527,N_20688);
nand U20822 (N_20822,N_20677,N_20617);
and U20823 (N_20823,N_20650,N_20521);
and U20824 (N_20824,N_20557,N_20630);
xor U20825 (N_20825,N_20713,N_20697);
nor U20826 (N_20826,N_20602,N_20589);
nand U20827 (N_20827,N_20592,N_20598);
nor U20828 (N_20828,N_20601,N_20612);
and U20829 (N_20829,N_20591,N_20730);
and U20830 (N_20830,N_20720,N_20684);
and U20831 (N_20831,N_20734,N_20647);
nand U20832 (N_20832,N_20525,N_20687);
nor U20833 (N_20833,N_20571,N_20728);
or U20834 (N_20834,N_20669,N_20731);
or U20835 (N_20835,N_20607,N_20533);
nor U20836 (N_20836,N_20623,N_20504);
nand U20837 (N_20837,N_20672,N_20732);
and U20838 (N_20838,N_20748,N_20694);
nor U20839 (N_20839,N_20562,N_20560);
nor U20840 (N_20840,N_20538,N_20619);
or U20841 (N_20841,N_20737,N_20512);
nor U20842 (N_20842,N_20581,N_20529);
or U20843 (N_20843,N_20661,N_20701);
nand U20844 (N_20844,N_20539,N_20704);
or U20845 (N_20845,N_20584,N_20519);
or U20846 (N_20846,N_20600,N_20620);
nand U20847 (N_20847,N_20604,N_20644);
or U20848 (N_20848,N_20611,N_20524);
nand U20849 (N_20849,N_20740,N_20565);
or U20850 (N_20850,N_20534,N_20640);
or U20851 (N_20851,N_20520,N_20553);
nor U20852 (N_20852,N_20733,N_20683);
or U20853 (N_20853,N_20566,N_20543);
nand U20854 (N_20854,N_20696,N_20678);
and U20855 (N_20855,N_20723,N_20514);
nor U20856 (N_20856,N_20596,N_20517);
or U20857 (N_20857,N_20711,N_20585);
nor U20858 (N_20858,N_20510,N_20608);
nand U20859 (N_20859,N_20515,N_20657);
and U20860 (N_20860,N_20682,N_20695);
and U20861 (N_20861,N_20660,N_20744);
nand U20862 (N_20862,N_20710,N_20580);
nor U20863 (N_20863,N_20633,N_20681);
nor U20864 (N_20864,N_20572,N_20588);
nor U20865 (N_20865,N_20722,N_20535);
nand U20866 (N_20866,N_20573,N_20628);
and U20867 (N_20867,N_20518,N_20664);
xor U20868 (N_20868,N_20708,N_20502);
or U20869 (N_20869,N_20659,N_20579);
or U20870 (N_20870,N_20613,N_20550);
nand U20871 (N_20871,N_20649,N_20523);
nand U20872 (N_20872,N_20721,N_20736);
nand U20873 (N_20873,N_20655,N_20656);
or U20874 (N_20874,N_20586,N_20665);
nand U20875 (N_20875,N_20517,N_20633);
nor U20876 (N_20876,N_20543,N_20695);
and U20877 (N_20877,N_20690,N_20733);
nand U20878 (N_20878,N_20513,N_20699);
nand U20879 (N_20879,N_20702,N_20621);
and U20880 (N_20880,N_20703,N_20585);
and U20881 (N_20881,N_20675,N_20503);
nor U20882 (N_20882,N_20651,N_20733);
nor U20883 (N_20883,N_20719,N_20557);
nand U20884 (N_20884,N_20614,N_20639);
or U20885 (N_20885,N_20699,N_20728);
or U20886 (N_20886,N_20615,N_20689);
or U20887 (N_20887,N_20558,N_20611);
and U20888 (N_20888,N_20736,N_20747);
nand U20889 (N_20889,N_20550,N_20600);
nor U20890 (N_20890,N_20684,N_20591);
nor U20891 (N_20891,N_20575,N_20703);
or U20892 (N_20892,N_20678,N_20627);
nand U20893 (N_20893,N_20521,N_20614);
nand U20894 (N_20894,N_20570,N_20702);
nand U20895 (N_20895,N_20703,N_20640);
nand U20896 (N_20896,N_20549,N_20556);
nor U20897 (N_20897,N_20571,N_20563);
and U20898 (N_20898,N_20559,N_20749);
and U20899 (N_20899,N_20663,N_20530);
nand U20900 (N_20900,N_20625,N_20679);
nand U20901 (N_20901,N_20524,N_20712);
nor U20902 (N_20902,N_20558,N_20517);
nand U20903 (N_20903,N_20615,N_20671);
or U20904 (N_20904,N_20689,N_20672);
nor U20905 (N_20905,N_20502,N_20532);
nand U20906 (N_20906,N_20528,N_20556);
nand U20907 (N_20907,N_20549,N_20500);
nand U20908 (N_20908,N_20682,N_20704);
and U20909 (N_20909,N_20644,N_20745);
nor U20910 (N_20910,N_20747,N_20670);
nand U20911 (N_20911,N_20689,N_20700);
nand U20912 (N_20912,N_20664,N_20532);
xor U20913 (N_20913,N_20545,N_20633);
or U20914 (N_20914,N_20709,N_20658);
xor U20915 (N_20915,N_20697,N_20554);
or U20916 (N_20916,N_20524,N_20674);
and U20917 (N_20917,N_20715,N_20531);
and U20918 (N_20918,N_20580,N_20612);
or U20919 (N_20919,N_20637,N_20682);
and U20920 (N_20920,N_20655,N_20732);
nand U20921 (N_20921,N_20534,N_20517);
nand U20922 (N_20922,N_20646,N_20543);
and U20923 (N_20923,N_20503,N_20659);
nor U20924 (N_20924,N_20622,N_20689);
nand U20925 (N_20925,N_20626,N_20560);
or U20926 (N_20926,N_20552,N_20745);
and U20927 (N_20927,N_20690,N_20517);
and U20928 (N_20928,N_20700,N_20545);
and U20929 (N_20929,N_20741,N_20553);
and U20930 (N_20930,N_20578,N_20521);
nand U20931 (N_20931,N_20709,N_20531);
nor U20932 (N_20932,N_20587,N_20637);
xor U20933 (N_20933,N_20704,N_20626);
nor U20934 (N_20934,N_20743,N_20564);
nand U20935 (N_20935,N_20535,N_20665);
and U20936 (N_20936,N_20729,N_20565);
or U20937 (N_20937,N_20738,N_20748);
nor U20938 (N_20938,N_20676,N_20510);
nor U20939 (N_20939,N_20616,N_20655);
or U20940 (N_20940,N_20541,N_20597);
and U20941 (N_20941,N_20692,N_20525);
nand U20942 (N_20942,N_20666,N_20749);
nor U20943 (N_20943,N_20680,N_20735);
or U20944 (N_20944,N_20540,N_20582);
nand U20945 (N_20945,N_20616,N_20659);
nor U20946 (N_20946,N_20509,N_20556);
nand U20947 (N_20947,N_20534,N_20740);
or U20948 (N_20948,N_20511,N_20634);
nor U20949 (N_20949,N_20707,N_20738);
or U20950 (N_20950,N_20628,N_20632);
nand U20951 (N_20951,N_20520,N_20565);
nand U20952 (N_20952,N_20553,N_20697);
or U20953 (N_20953,N_20693,N_20563);
and U20954 (N_20954,N_20650,N_20615);
or U20955 (N_20955,N_20555,N_20651);
nand U20956 (N_20956,N_20737,N_20520);
and U20957 (N_20957,N_20545,N_20585);
and U20958 (N_20958,N_20587,N_20676);
or U20959 (N_20959,N_20517,N_20617);
nand U20960 (N_20960,N_20545,N_20570);
or U20961 (N_20961,N_20523,N_20589);
and U20962 (N_20962,N_20739,N_20641);
nor U20963 (N_20963,N_20545,N_20602);
nor U20964 (N_20964,N_20715,N_20642);
nand U20965 (N_20965,N_20634,N_20718);
nor U20966 (N_20966,N_20563,N_20560);
or U20967 (N_20967,N_20704,N_20625);
nor U20968 (N_20968,N_20515,N_20588);
nor U20969 (N_20969,N_20629,N_20690);
and U20970 (N_20970,N_20680,N_20504);
and U20971 (N_20971,N_20683,N_20712);
or U20972 (N_20972,N_20550,N_20673);
nand U20973 (N_20973,N_20677,N_20666);
and U20974 (N_20974,N_20580,N_20648);
nor U20975 (N_20975,N_20680,N_20742);
or U20976 (N_20976,N_20541,N_20585);
or U20977 (N_20977,N_20540,N_20565);
nand U20978 (N_20978,N_20651,N_20625);
nor U20979 (N_20979,N_20587,N_20639);
nor U20980 (N_20980,N_20747,N_20682);
and U20981 (N_20981,N_20661,N_20674);
and U20982 (N_20982,N_20636,N_20521);
nor U20983 (N_20983,N_20684,N_20608);
and U20984 (N_20984,N_20720,N_20524);
nand U20985 (N_20985,N_20624,N_20718);
or U20986 (N_20986,N_20589,N_20522);
nand U20987 (N_20987,N_20739,N_20678);
nor U20988 (N_20988,N_20717,N_20639);
and U20989 (N_20989,N_20626,N_20719);
nand U20990 (N_20990,N_20640,N_20667);
nand U20991 (N_20991,N_20631,N_20517);
nand U20992 (N_20992,N_20549,N_20645);
nor U20993 (N_20993,N_20512,N_20597);
nor U20994 (N_20994,N_20619,N_20573);
nand U20995 (N_20995,N_20506,N_20613);
or U20996 (N_20996,N_20703,N_20687);
or U20997 (N_20997,N_20502,N_20514);
nor U20998 (N_20998,N_20688,N_20702);
or U20999 (N_20999,N_20722,N_20542);
and U21000 (N_21000,N_20767,N_20975);
or U21001 (N_21001,N_20854,N_20903);
nand U21002 (N_21002,N_20887,N_20984);
or U21003 (N_21003,N_20750,N_20789);
nand U21004 (N_21004,N_20781,N_20818);
nor U21005 (N_21005,N_20960,N_20798);
nor U21006 (N_21006,N_20764,N_20782);
nor U21007 (N_21007,N_20950,N_20753);
and U21008 (N_21008,N_20925,N_20996);
and U21009 (N_21009,N_20986,N_20904);
and U21010 (N_21010,N_20922,N_20963);
and U21011 (N_21011,N_20916,N_20858);
and U21012 (N_21012,N_20876,N_20882);
nor U21013 (N_21013,N_20968,N_20843);
nand U21014 (N_21014,N_20787,N_20779);
nor U21015 (N_21015,N_20971,N_20848);
or U21016 (N_21016,N_20997,N_20805);
nor U21017 (N_21017,N_20969,N_20861);
nand U21018 (N_21018,N_20771,N_20883);
or U21019 (N_21019,N_20754,N_20994);
nor U21020 (N_21020,N_20772,N_20927);
and U21021 (N_21021,N_20948,N_20900);
nand U21022 (N_21022,N_20838,N_20826);
nand U21023 (N_21023,N_20845,N_20766);
and U21024 (N_21024,N_20831,N_20769);
nor U21025 (N_21025,N_20979,N_20906);
and U21026 (N_21026,N_20919,N_20983);
or U21027 (N_21027,N_20911,N_20929);
nand U21028 (N_21028,N_20801,N_20758);
nor U21029 (N_21029,N_20774,N_20988);
and U21030 (N_21030,N_20846,N_20952);
nor U21031 (N_21031,N_20870,N_20913);
and U21032 (N_21032,N_20940,N_20851);
nand U21033 (N_21033,N_20866,N_20755);
and U21034 (N_21034,N_20867,N_20822);
or U21035 (N_21035,N_20943,N_20933);
nor U21036 (N_21036,N_20809,N_20751);
or U21037 (N_21037,N_20918,N_20966);
and U21038 (N_21038,N_20856,N_20784);
nor U21039 (N_21039,N_20930,N_20797);
and U21040 (N_21040,N_20901,N_20990);
nor U21041 (N_21041,N_20978,N_20862);
nand U21042 (N_21042,N_20821,N_20874);
and U21043 (N_21043,N_20756,N_20850);
nand U21044 (N_21044,N_20880,N_20871);
and U21045 (N_21045,N_20985,N_20763);
and U21046 (N_21046,N_20820,N_20967);
and U21047 (N_21047,N_20965,N_20895);
nor U21048 (N_21048,N_20891,N_20802);
and U21049 (N_21049,N_20863,N_20780);
nand U21050 (N_21050,N_20869,N_20855);
nor U21051 (N_21051,N_20910,N_20860);
nor U21052 (N_21052,N_20907,N_20795);
nor U21053 (N_21053,N_20872,N_20897);
and U21054 (N_21054,N_20998,N_20973);
or U21055 (N_21055,N_20878,N_20808);
or U21056 (N_21056,N_20972,N_20834);
and U21057 (N_21057,N_20841,N_20977);
nor U21058 (N_21058,N_20892,N_20951);
nand U21059 (N_21059,N_20823,N_20945);
nand U21060 (N_21060,N_20859,N_20964);
or U21061 (N_21061,N_20926,N_20825);
nor U21062 (N_21062,N_20937,N_20885);
nor U21063 (N_21063,N_20877,N_20803);
nand U21064 (N_21064,N_20777,N_20909);
nand U21065 (N_21065,N_20835,N_20836);
and U21066 (N_21066,N_20778,N_20917);
nand U21067 (N_21067,N_20840,N_20768);
and U21068 (N_21068,N_20824,N_20944);
nor U21069 (N_21069,N_20844,N_20786);
nor U21070 (N_21070,N_20793,N_20810);
and U21071 (N_21071,N_20816,N_20959);
nor U21072 (N_21072,N_20961,N_20899);
or U21073 (N_21073,N_20773,N_20814);
nor U21074 (N_21074,N_20800,N_20832);
nor U21075 (N_21075,N_20954,N_20757);
nor U21076 (N_21076,N_20941,N_20938);
or U21077 (N_21077,N_20982,N_20837);
and U21078 (N_21078,N_20981,N_20776);
and U21079 (N_21079,N_20953,N_20886);
nand U21080 (N_21080,N_20760,N_20970);
and U21081 (N_21081,N_20830,N_20939);
or U21082 (N_21082,N_20962,N_20914);
or U21083 (N_21083,N_20864,N_20879);
or U21084 (N_21084,N_20934,N_20991);
nand U21085 (N_21085,N_20912,N_20752);
and U21086 (N_21086,N_20857,N_20765);
nand U21087 (N_21087,N_20759,N_20842);
and U21088 (N_21088,N_20819,N_20935);
or U21089 (N_21089,N_20908,N_20770);
nand U21090 (N_21090,N_20839,N_20799);
or U21091 (N_21091,N_20889,N_20807);
and U21092 (N_21092,N_20888,N_20949);
and U21093 (N_21093,N_20788,N_20898);
nand U21094 (N_21094,N_20833,N_20804);
nor U21095 (N_21095,N_20813,N_20920);
and U21096 (N_21096,N_20868,N_20956);
or U21097 (N_21097,N_20884,N_20791);
nor U21098 (N_21098,N_20931,N_20811);
and U21099 (N_21099,N_20915,N_20995);
nand U21100 (N_21100,N_20894,N_20974);
and U21101 (N_21101,N_20924,N_20955);
nor U21102 (N_21102,N_20783,N_20828);
or U21103 (N_21103,N_20928,N_20853);
and U21104 (N_21104,N_20827,N_20881);
or U21105 (N_21105,N_20806,N_20976);
or U21106 (N_21106,N_20921,N_20932);
and U21107 (N_21107,N_20829,N_20902);
and U21108 (N_21108,N_20989,N_20957);
or U21109 (N_21109,N_20796,N_20815);
nor U21110 (N_21110,N_20812,N_20923);
nand U21111 (N_21111,N_20992,N_20905);
and U21112 (N_21112,N_20785,N_20847);
xor U21113 (N_21113,N_20958,N_20794);
or U21114 (N_21114,N_20987,N_20936);
and U21115 (N_21115,N_20946,N_20775);
and U21116 (N_21116,N_20792,N_20942);
xor U21117 (N_21117,N_20875,N_20790);
nor U21118 (N_21118,N_20896,N_20817);
or U21119 (N_21119,N_20865,N_20873);
and U21120 (N_21120,N_20980,N_20762);
or U21121 (N_21121,N_20893,N_20890);
or U21122 (N_21122,N_20993,N_20761);
nor U21123 (N_21123,N_20849,N_20999);
nor U21124 (N_21124,N_20852,N_20947);
and U21125 (N_21125,N_20817,N_20813);
nand U21126 (N_21126,N_20986,N_20866);
nor U21127 (N_21127,N_20775,N_20962);
and U21128 (N_21128,N_20877,N_20935);
and U21129 (N_21129,N_20952,N_20752);
nand U21130 (N_21130,N_20817,N_20951);
or U21131 (N_21131,N_20968,N_20877);
and U21132 (N_21132,N_20762,N_20934);
or U21133 (N_21133,N_20776,N_20858);
or U21134 (N_21134,N_20768,N_20927);
nor U21135 (N_21135,N_20865,N_20764);
nand U21136 (N_21136,N_20869,N_20980);
and U21137 (N_21137,N_20994,N_20898);
nor U21138 (N_21138,N_20984,N_20895);
or U21139 (N_21139,N_20781,N_20789);
nor U21140 (N_21140,N_20887,N_20803);
or U21141 (N_21141,N_20797,N_20947);
and U21142 (N_21142,N_20994,N_20959);
nor U21143 (N_21143,N_20751,N_20808);
nor U21144 (N_21144,N_20816,N_20836);
nand U21145 (N_21145,N_20762,N_20937);
nor U21146 (N_21146,N_20907,N_20936);
nor U21147 (N_21147,N_20787,N_20999);
nor U21148 (N_21148,N_20871,N_20901);
and U21149 (N_21149,N_20762,N_20948);
and U21150 (N_21150,N_20944,N_20941);
nand U21151 (N_21151,N_20848,N_20950);
nor U21152 (N_21152,N_20781,N_20928);
nand U21153 (N_21153,N_20810,N_20970);
or U21154 (N_21154,N_20968,N_20862);
or U21155 (N_21155,N_20965,N_20819);
nor U21156 (N_21156,N_20979,N_20812);
and U21157 (N_21157,N_20840,N_20995);
or U21158 (N_21158,N_20983,N_20757);
or U21159 (N_21159,N_20771,N_20913);
or U21160 (N_21160,N_20918,N_20980);
nor U21161 (N_21161,N_20766,N_20970);
nor U21162 (N_21162,N_20835,N_20857);
or U21163 (N_21163,N_20956,N_20936);
nor U21164 (N_21164,N_20823,N_20802);
nand U21165 (N_21165,N_20978,N_20865);
and U21166 (N_21166,N_20987,N_20991);
nor U21167 (N_21167,N_20920,N_20781);
nand U21168 (N_21168,N_20930,N_20808);
or U21169 (N_21169,N_20954,N_20958);
or U21170 (N_21170,N_20869,N_20958);
or U21171 (N_21171,N_20907,N_20837);
nand U21172 (N_21172,N_20917,N_20811);
and U21173 (N_21173,N_20918,N_20976);
nor U21174 (N_21174,N_20920,N_20940);
nor U21175 (N_21175,N_20990,N_20865);
or U21176 (N_21176,N_20990,N_20995);
nand U21177 (N_21177,N_20857,N_20788);
nor U21178 (N_21178,N_20921,N_20954);
or U21179 (N_21179,N_20872,N_20798);
nand U21180 (N_21180,N_20853,N_20757);
or U21181 (N_21181,N_20952,N_20837);
and U21182 (N_21182,N_20814,N_20962);
or U21183 (N_21183,N_20985,N_20757);
nor U21184 (N_21184,N_20897,N_20962);
or U21185 (N_21185,N_20755,N_20803);
and U21186 (N_21186,N_20929,N_20913);
nand U21187 (N_21187,N_20823,N_20967);
or U21188 (N_21188,N_20765,N_20811);
xnor U21189 (N_21189,N_20772,N_20974);
nand U21190 (N_21190,N_20988,N_20864);
and U21191 (N_21191,N_20750,N_20792);
nand U21192 (N_21192,N_20938,N_20930);
nand U21193 (N_21193,N_20798,N_20799);
nor U21194 (N_21194,N_20815,N_20897);
and U21195 (N_21195,N_20865,N_20864);
nand U21196 (N_21196,N_20808,N_20950);
and U21197 (N_21197,N_20790,N_20954);
nor U21198 (N_21198,N_20943,N_20863);
nand U21199 (N_21199,N_20788,N_20843);
or U21200 (N_21200,N_20825,N_20982);
or U21201 (N_21201,N_20988,N_20907);
nor U21202 (N_21202,N_20837,N_20814);
nand U21203 (N_21203,N_20969,N_20957);
or U21204 (N_21204,N_20805,N_20803);
or U21205 (N_21205,N_20856,N_20818);
nand U21206 (N_21206,N_20802,N_20779);
nor U21207 (N_21207,N_20798,N_20967);
nand U21208 (N_21208,N_20832,N_20936);
or U21209 (N_21209,N_20856,N_20844);
or U21210 (N_21210,N_20919,N_20992);
nand U21211 (N_21211,N_20861,N_20977);
nor U21212 (N_21212,N_20983,N_20960);
and U21213 (N_21213,N_20822,N_20884);
nand U21214 (N_21214,N_20852,N_20898);
and U21215 (N_21215,N_20823,N_20822);
and U21216 (N_21216,N_20899,N_20780);
nor U21217 (N_21217,N_20918,N_20834);
nor U21218 (N_21218,N_20988,N_20760);
nor U21219 (N_21219,N_20998,N_20901);
xnor U21220 (N_21220,N_20834,N_20957);
nor U21221 (N_21221,N_20840,N_20850);
nand U21222 (N_21222,N_20987,N_20912);
and U21223 (N_21223,N_20898,N_20906);
nor U21224 (N_21224,N_20915,N_20825);
or U21225 (N_21225,N_20993,N_20943);
or U21226 (N_21226,N_20835,N_20952);
nor U21227 (N_21227,N_20911,N_20970);
nand U21228 (N_21228,N_20845,N_20984);
and U21229 (N_21229,N_20915,N_20798);
or U21230 (N_21230,N_20959,N_20810);
and U21231 (N_21231,N_20878,N_20830);
nor U21232 (N_21232,N_20824,N_20937);
nor U21233 (N_21233,N_20752,N_20753);
nor U21234 (N_21234,N_20756,N_20771);
and U21235 (N_21235,N_20894,N_20889);
or U21236 (N_21236,N_20854,N_20835);
or U21237 (N_21237,N_20960,N_20889);
and U21238 (N_21238,N_20764,N_20772);
and U21239 (N_21239,N_20846,N_20886);
nor U21240 (N_21240,N_20752,N_20755);
and U21241 (N_21241,N_20895,N_20958);
nor U21242 (N_21242,N_20859,N_20959);
or U21243 (N_21243,N_20972,N_20796);
nor U21244 (N_21244,N_20835,N_20868);
nand U21245 (N_21245,N_20996,N_20829);
nor U21246 (N_21246,N_20805,N_20792);
and U21247 (N_21247,N_20952,N_20782);
or U21248 (N_21248,N_20846,N_20934);
and U21249 (N_21249,N_20889,N_20976);
nand U21250 (N_21250,N_21102,N_21033);
nand U21251 (N_21251,N_21009,N_21079);
nor U21252 (N_21252,N_21249,N_21001);
or U21253 (N_21253,N_21062,N_21141);
or U21254 (N_21254,N_21220,N_21107);
and U21255 (N_21255,N_21061,N_21140);
or U21256 (N_21256,N_21166,N_21074);
nand U21257 (N_21257,N_21188,N_21086);
nor U21258 (N_21258,N_21103,N_21064);
nor U21259 (N_21259,N_21087,N_21017);
nand U21260 (N_21260,N_21012,N_21067);
or U21261 (N_21261,N_21145,N_21022);
and U21262 (N_21262,N_21124,N_21100);
nand U21263 (N_21263,N_21010,N_21076);
nor U21264 (N_21264,N_21167,N_21117);
and U21265 (N_21265,N_21023,N_21218);
and U21266 (N_21266,N_21097,N_21189);
or U21267 (N_21267,N_21197,N_21057);
or U21268 (N_21268,N_21131,N_21169);
nand U21269 (N_21269,N_21090,N_21049);
or U21270 (N_21270,N_21186,N_21201);
or U21271 (N_21271,N_21066,N_21094);
nor U21272 (N_21272,N_21025,N_21164);
nor U21273 (N_21273,N_21165,N_21198);
nand U21274 (N_21274,N_21109,N_21154);
and U21275 (N_21275,N_21194,N_21006);
or U21276 (N_21276,N_21146,N_21065);
or U21277 (N_21277,N_21014,N_21002);
or U21278 (N_21278,N_21055,N_21228);
and U21279 (N_21279,N_21245,N_21044);
and U21280 (N_21280,N_21138,N_21068);
nand U21281 (N_21281,N_21199,N_21207);
nor U21282 (N_21282,N_21230,N_21018);
nor U21283 (N_21283,N_21120,N_21248);
and U21284 (N_21284,N_21106,N_21227);
nor U21285 (N_21285,N_21004,N_21225);
nor U21286 (N_21286,N_21026,N_21091);
nor U21287 (N_21287,N_21233,N_21213);
or U21288 (N_21288,N_21125,N_21187);
and U21289 (N_21289,N_21095,N_21035);
nand U21290 (N_21290,N_21132,N_21144);
or U21291 (N_21291,N_21204,N_21029);
nor U21292 (N_21292,N_21147,N_21093);
and U21293 (N_21293,N_21172,N_21115);
and U21294 (N_21294,N_21151,N_21092);
nand U21295 (N_21295,N_21148,N_21110);
nand U21296 (N_21296,N_21142,N_21008);
nand U21297 (N_21297,N_21206,N_21239);
and U21298 (N_21298,N_21114,N_21080);
or U21299 (N_21299,N_21098,N_21123);
or U21300 (N_21300,N_21101,N_21081);
nor U21301 (N_21301,N_21217,N_21232);
or U21302 (N_21302,N_21021,N_21112);
nand U21303 (N_21303,N_21036,N_21136);
and U21304 (N_21304,N_21129,N_21168);
or U21305 (N_21305,N_21040,N_21237);
and U21306 (N_21306,N_21089,N_21244);
nand U21307 (N_21307,N_21236,N_21143);
or U21308 (N_21308,N_21139,N_21046);
or U21309 (N_21309,N_21108,N_21174);
or U21310 (N_21310,N_21192,N_21212);
or U21311 (N_21311,N_21039,N_21134);
nor U21312 (N_21312,N_21191,N_21231);
and U21313 (N_21313,N_21111,N_21041);
or U21314 (N_21314,N_21122,N_21105);
or U21315 (N_21315,N_21128,N_21203);
and U21316 (N_21316,N_21032,N_21047);
and U21317 (N_21317,N_21037,N_21241);
or U21318 (N_21318,N_21177,N_21162);
nand U21319 (N_21319,N_21156,N_21137);
and U21320 (N_21320,N_21229,N_21003);
nor U21321 (N_21321,N_21159,N_21030);
nand U21322 (N_21322,N_21069,N_21027);
nand U21323 (N_21323,N_21020,N_21000);
nand U21324 (N_21324,N_21222,N_21171);
or U21325 (N_21325,N_21082,N_21173);
and U21326 (N_21326,N_21011,N_21034);
and U21327 (N_21327,N_21059,N_21083);
or U21328 (N_21328,N_21121,N_21056);
nor U21329 (N_21329,N_21084,N_21242);
or U21330 (N_21330,N_21053,N_21214);
nor U21331 (N_21331,N_21050,N_21208);
or U21332 (N_21332,N_21119,N_21005);
nand U21333 (N_21333,N_21163,N_21113);
and U21334 (N_21334,N_21135,N_21216);
and U21335 (N_21335,N_21054,N_21099);
nand U21336 (N_21336,N_21221,N_21118);
nor U21337 (N_21337,N_21038,N_21190);
nor U21338 (N_21338,N_21060,N_21007);
nand U21339 (N_21339,N_21150,N_21104);
nor U21340 (N_21340,N_21031,N_21149);
nor U21341 (N_21341,N_21161,N_21200);
nand U21342 (N_21342,N_21077,N_21016);
and U21343 (N_21343,N_21158,N_21210);
and U21344 (N_21344,N_21176,N_21179);
nand U21345 (N_21345,N_21127,N_21235);
and U21346 (N_21346,N_21178,N_21058);
nand U21347 (N_21347,N_21075,N_21015);
or U21348 (N_21348,N_21073,N_21205);
and U21349 (N_21349,N_21185,N_21045);
and U21350 (N_21350,N_21063,N_21219);
nor U21351 (N_21351,N_21234,N_21211);
or U21352 (N_21352,N_21133,N_21052);
or U21353 (N_21353,N_21152,N_21019);
or U21354 (N_21354,N_21160,N_21195);
or U21355 (N_21355,N_21088,N_21238);
or U21356 (N_21356,N_21196,N_21202);
or U21357 (N_21357,N_21013,N_21184);
or U21358 (N_21358,N_21078,N_21070);
or U21359 (N_21359,N_21024,N_21240);
and U21360 (N_21360,N_21243,N_21223);
nor U21361 (N_21361,N_21048,N_21130);
nand U21362 (N_21362,N_21155,N_21180);
nor U21363 (N_21363,N_21072,N_21182);
xnor U21364 (N_21364,N_21181,N_21193);
xor U21365 (N_21365,N_21175,N_21247);
nand U21366 (N_21366,N_21153,N_21215);
or U21367 (N_21367,N_21126,N_21085);
or U21368 (N_21368,N_21043,N_21051);
or U21369 (N_21369,N_21209,N_21183);
or U21370 (N_21370,N_21246,N_21116);
nand U21371 (N_21371,N_21157,N_21096);
and U21372 (N_21372,N_21042,N_21226);
nand U21373 (N_21373,N_21028,N_21071);
or U21374 (N_21374,N_21224,N_21170);
or U21375 (N_21375,N_21235,N_21209);
nand U21376 (N_21376,N_21070,N_21010);
nand U21377 (N_21377,N_21050,N_21019);
and U21378 (N_21378,N_21182,N_21056);
or U21379 (N_21379,N_21205,N_21102);
nand U21380 (N_21380,N_21140,N_21034);
nor U21381 (N_21381,N_21137,N_21169);
and U21382 (N_21382,N_21027,N_21046);
nand U21383 (N_21383,N_21054,N_21021);
or U21384 (N_21384,N_21121,N_21045);
nand U21385 (N_21385,N_21047,N_21201);
and U21386 (N_21386,N_21084,N_21105);
or U21387 (N_21387,N_21217,N_21040);
nand U21388 (N_21388,N_21142,N_21183);
nand U21389 (N_21389,N_21030,N_21172);
nand U21390 (N_21390,N_21247,N_21144);
nand U21391 (N_21391,N_21029,N_21019);
nor U21392 (N_21392,N_21242,N_21220);
or U21393 (N_21393,N_21040,N_21176);
nor U21394 (N_21394,N_21231,N_21065);
nand U21395 (N_21395,N_21023,N_21139);
nor U21396 (N_21396,N_21111,N_21201);
nor U21397 (N_21397,N_21084,N_21077);
nor U21398 (N_21398,N_21018,N_21209);
nand U21399 (N_21399,N_21131,N_21179);
nand U21400 (N_21400,N_21003,N_21246);
nand U21401 (N_21401,N_21199,N_21031);
nand U21402 (N_21402,N_21141,N_21026);
and U21403 (N_21403,N_21182,N_21171);
or U21404 (N_21404,N_21074,N_21196);
nor U21405 (N_21405,N_21102,N_21234);
nor U21406 (N_21406,N_21118,N_21115);
and U21407 (N_21407,N_21022,N_21157);
nand U21408 (N_21408,N_21007,N_21100);
nand U21409 (N_21409,N_21195,N_21043);
and U21410 (N_21410,N_21155,N_21111);
and U21411 (N_21411,N_21091,N_21082);
or U21412 (N_21412,N_21114,N_21157);
and U21413 (N_21413,N_21029,N_21082);
or U21414 (N_21414,N_21189,N_21010);
or U21415 (N_21415,N_21172,N_21147);
nand U21416 (N_21416,N_21179,N_21148);
and U21417 (N_21417,N_21225,N_21068);
and U21418 (N_21418,N_21029,N_21203);
nand U21419 (N_21419,N_21034,N_21062);
nand U21420 (N_21420,N_21035,N_21040);
or U21421 (N_21421,N_21097,N_21147);
nor U21422 (N_21422,N_21105,N_21039);
or U21423 (N_21423,N_21179,N_21096);
nand U21424 (N_21424,N_21083,N_21020);
or U21425 (N_21425,N_21028,N_21039);
nand U21426 (N_21426,N_21163,N_21195);
nor U21427 (N_21427,N_21179,N_21086);
and U21428 (N_21428,N_21186,N_21207);
and U21429 (N_21429,N_21053,N_21078);
and U21430 (N_21430,N_21210,N_21025);
or U21431 (N_21431,N_21134,N_21032);
nand U21432 (N_21432,N_21192,N_21097);
nor U21433 (N_21433,N_21216,N_21001);
nor U21434 (N_21434,N_21087,N_21096);
nand U21435 (N_21435,N_21133,N_21097);
nand U21436 (N_21436,N_21021,N_21148);
nor U21437 (N_21437,N_21011,N_21013);
nand U21438 (N_21438,N_21199,N_21019);
or U21439 (N_21439,N_21091,N_21036);
and U21440 (N_21440,N_21021,N_21022);
nor U21441 (N_21441,N_21022,N_21163);
nand U21442 (N_21442,N_21179,N_21055);
or U21443 (N_21443,N_21197,N_21129);
nand U21444 (N_21444,N_21028,N_21198);
xor U21445 (N_21445,N_21022,N_21189);
nor U21446 (N_21446,N_21239,N_21010);
and U21447 (N_21447,N_21222,N_21150);
nand U21448 (N_21448,N_21149,N_21132);
or U21449 (N_21449,N_21018,N_21109);
nand U21450 (N_21450,N_21219,N_21004);
and U21451 (N_21451,N_21165,N_21225);
or U21452 (N_21452,N_21141,N_21031);
xor U21453 (N_21453,N_21123,N_21243);
or U21454 (N_21454,N_21234,N_21004);
or U21455 (N_21455,N_21043,N_21203);
nor U21456 (N_21456,N_21142,N_21126);
nand U21457 (N_21457,N_21240,N_21133);
nand U21458 (N_21458,N_21075,N_21110);
and U21459 (N_21459,N_21211,N_21158);
nor U21460 (N_21460,N_21182,N_21031);
and U21461 (N_21461,N_21048,N_21193);
nor U21462 (N_21462,N_21206,N_21120);
nor U21463 (N_21463,N_21032,N_21013);
nor U21464 (N_21464,N_21045,N_21198);
and U21465 (N_21465,N_21191,N_21072);
or U21466 (N_21466,N_21020,N_21018);
nor U21467 (N_21467,N_21042,N_21097);
or U21468 (N_21468,N_21033,N_21012);
nor U21469 (N_21469,N_21167,N_21190);
or U21470 (N_21470,N_21041,N_21006);
nor U21471 (N_21471,N_21005,N_21104);
or U21472 (N_21472,N_21073,N_21133);
or U21473 (N_21473,N_21154,N_21133);
nand U21474 (N_21474,N_21117,N_21033);
nand U21475 (N_21475,N_21140,N_21046);
or U21476 (N_21476,N_21025,N_21064);
nor U21477 (N_21477,N_21115,N_21084);
nand U21478 (N_21478,N_21145,N_21134);
and U21479 (N_21479,N_21210,N_21160);
and U21480 (N_21480,N_21121,N_21010);
nand U21481 (N_21481,N_21024,N_21104);
nand U21482 (N_21482,N_21177,N_21070);
and U21483 (N_21483,N_21054,N_21174);
or U21484 (N_21484,N_21216,N_21239);
or U21485 (N_21485,N_21136,N_21122);
and U21486 (N_21486,N_21138,N_21045);
nor U21487 (N_21487,N_21087,N_21064);
and U21488 (N_21488,N_21227,N_21080);
or U21489 (N_21489,N_21134,N_21113);
and U21490 (N_21490,N_21178,N_21003);
or U21491 (N_21491,N_21246,N_21062);
nor U21492 (N_21492,N_21178,N_21240);
nand U21493 (N_21493,N_21037,N_21205);
nor U21494 (N_21494,N_21047,N_21249);
nor U21495 (N_21495,N_21027,N_21206);
or U21496 (N_21496,N_21099,N_21124);
and U21497 (N_21497,N_21074,N_21089);
and U21498 (N_21498,N_21247,N_21199);
nand U21499 (N_21499,N_21205,N_21086);
or U21500 (N_21500,N_21486,N_21282);
xnor U21501 (N_21501,N_21459,N_21386);
and U21502 (N_21502,N_21340,N_21287);
and U21503 (N_21503,N_21328,N_21451);
nor U21504 (N_21504,N_21312,N_21415);
nor U21505 (N_21505,N_21498,N_21339);
nand U21506 (N_21506,N_21338,N_21349);
nand U21507 (N_21507,N_21447,N_21381);
nor U21508 (N_21508,N_21416,N_21412);
and U21509 (N_21509,N_21280,N_21315);
nor U21510 (N_21510,N_21421,N_21460);
nor U21511 (N_21511,N_21275,N_21495);
nor U21512 (N_21512,N_21331,N_21329);
and U21513 (N_21513,N_21389,N_21347);
and U21514 (N_21514,N_21298,N_21255);
xnor U21515 (N_21515,N_21292,N_21343);
and U21516 (N_21516,N_21403,N_21448);
or U21517 (N_21517,N_21436,N_21390);
nor U21518 (N_21518,N_21363,N_21470);
nand U21519 (N_21519,N_21336,N_21377);
nor U21520 (N_21520,N_21308,N_21469);
nor U21521 (N_21521,N_21466,N_21424);
and U21522 (N_21522,N_21361,N_21324);
and U21523 (N_21523,N_21290,N_21409);
nand U21524 (N_21524,N_21283,N_21482);
or U21525 (N_21525,N_21358,N_21410);
and U21526 (N_21526,N_21422,N_21462);
nor U21527 (N_21527,N_21395,N_21333);
and U21528 (N_21528,N_21446,N_21406);
nor U21529 (N_21529,N_21429,N_21352);
and U21530 (N_21530,N_21369,N_21260);
nor U21531 (N_21531,N_21267,N_21440);
nor U21532 (N_21532,N_21357,N_21285);
nand U21533 (N_21533,N_21423,N_21301);
xnor U21534 (N_21534,N_21305,N_21316);
and U21535 (N_21535,N_21350,N_21437);
or U21536 (N_21536,N_21334,N_21491);
nand U21537 (N_21537,N_21360,N_21456);
nor U21538 (N_21538,N_21380,N_21262);
or U21539 (N_21539,N_21346,N_21345);
and U21540 (N_21540,N_21319,N_21259);
or U21541 (N_21541,N_21373,N_21256);
nor U21542 (N_21542,N_21487,N_21480);
nand U21543 (N_21543,N_21253,N_21356);
nor U21544 (N_21544,N_21266,N_21318);
or U21545 (N_21545,N_21393,N_21281);
or U21546 (N_21546,N_21370,N_21310);
nor U21547 (N_21547,N_21457,N_21418);
xnor U21548 (N_21548,N_21304,N_21427);
or U21549 (N_21549,N_21320,N_21379);
nand U21550 (N_21550,N_21453,N_21289);
and U21551 (N_21551,N_21264,N_21426);
and U21552 (N_21552,N_21367,N_21279);
nand U21553 (N_21553,N_21420,N_21384);
nand U21554 (N_21554,N_21365,N_21351);
or U21555 (N_21555,N_21394,N_21483);
and U21556 (N_21556,N_21408,N_21332);
or U21557 (N_21557,N_21385,N_21317);
nor U21558 (N_21558,N_21321,N_21295);
nor U21559 (N_21559,N_21404,N_21261);
nor U21560 (N_21560,N_21489,N_21414);
and U21561 (N_21561,N_21330,N_21323);
nand U21562 (N_21562,N_21327,N_21477);
nor U21563 (N_21563,N_21311,N_21382);
or U21564 (N_21564,N_21461,N_21433);
and U21565 (N_21565,N_21258,N_21467);
nand U21566 (N_21566,N_21326,N_21428);
and U21567 (N_21567,N_21374,N_21413);
nand U21568 (N_21568,N_21419,N_21371);
and U21569 (N_21569,N_21454,N_21263);
nand U21570 (N_21570,N_21432,N_21344);
or U21571 (N_21571,N_21376,N_21274);
and U21572 (N_21572,N_21368,N_21271);
and U21573 (N_21573,N_21400,N_21322);
and U21574 (N_21574,N_21388,N_21354);
and U21575 (N_21575,N_21391,N_21257);
or U21576 (N_21576,N_21284,N_21299);
nor U21577 (N_21577,N_21435,N_21364);
nand U21578 (N_21578,N_21383,N_21300);
and U21579 (N_21579,N_21399,N_21476);
nand U21580 (N_21580,N_21337,N_21397);
nor U21581 (N_21581,N_21484,N_21309);
nand U21582 (N_21582,N_21473,N_21431);
and U21583 (N_21583,N_21341,N_21288);
and U21584 (N_21584,N_21492,N_21475);
nor U21585 (N_21585,N_21313,N_21471);
nand U21586 (N_21586,N_21254,N_21335);
nor U21587 (N_21587,N_21425,N_21272);
and U21588 (N_21588,N_21439,N_21252);
nand U21589 (N_21589,N_21375,N_21302);
nand U21590 (N_21590,N_21401,N_21297);
nor U21591 (N_21591,N_21478,N_21499);
nor U21592 (N_21592,N_21496,N_21441);
or U21593 (N_21593,N_21296,N_21303);
nand U21594 (N_21594,N_21455,N_21407);
nand U21595 (N_21595,N_21430,N_21493);
nand U21596 (N_21596,N_21325,N_21474);
and U21597 (N_21597,N_21268,N_21291);
nor U21598 (N_21598,N_21494,N_21396);
nand U21599 (N_21599,N_21438,N_21434);
and U21600 (N_21600,N_21355,N_21402);
nand U21601 (N_21601,N_21278,N_21468);
and U21602 (N_21602,N_21444,N_21306);
or U21603 (N_21603,N_21270,N_21276);
and U21604 (N_21604,N_21443,N_21464);
nand U21605 (N_21605,N_21465,N_21342);
or U21606 (N_21606,N_21314,N_21265);
nor U21607 (N_21607,N_21449,N_21307);
or U21608 (N_21608,N_21411,N_21445);
and U21609 (N_21609,N_21458,N_21250);
nand U21610 (N_21610,N_21359,N_21348);
nand U21611 (N_21611,N_21452,N_21366);
xor U21612 (N_21612,N_21481,N_21392);
and U21613 (N_21613,N_21251,N_21472);
nor U21614 (N_21614,N_21417,N_21362);
nand U21615 (N_21615,N_21479,N_21273);
nor U21616 (N_21616,N_21463,N_21353);
and U21617 (N_21617,N_21294,N_21405);
nor U21618 (N_21618,N_21286,N_21497);
or U21619 (N_21619,N_21442,N_21378);
or U21620 (N_21620,N_21269,N_21485);
nand U21621 (N_21621,N_21450,N_21488);
and U21622 (N_21622,N_21372,N_21293);
nor U21623 (N_21623,N_21387,N_21277);
or U21624 (N_21624,N_21398,N_21490);
or U21625 (N_21625,N_21441,N_21343);
nor U21626 (N_21626,N_21400,N_21440);
nand U21627 (N_21627,N_21292,N_21379);
or U21628 (N_21628,N_21496,N_21483);
and U21629 (N_21629,N_21433,N_21370);
nor U21630 (N_21630,N_21479,N_21423);
and U21631 (N_21631,N_21398,N_21295);
nand U21632 (N_21632,N_21400,N_21394);
and U21633 (N_21633,N_21424,N_21253);
or U21634 (N_21634,N_21396,N_21271);
nand U21635 (N_21635,N_21338,N_21469);
or U21636 (N_21636,N_21347,N_21413);
or U21637 (N_21637,N_21370,N_21333);
or U21638 (N_21638,N_21305,N_21404);
nor U21639 (N_21639,N_21311,N_21491);
nor U21640 (N_21640,N_21309,N_21409);
or U21641 (N_21641,N_21481,N_21463);
or U21642 (N_21642,N_21385,N_21402);
nor U21643 (N_21643,N_21363,N_21487);
and U21644 (N_21644,N_21250,N_21279);
or U21645 (N_21645,N_21275,N_21470);
nand U21646 (N_21646,N_21422,N_21467);
nor U21647 (N_21647,N_21431,N_21373);
nor U21648 (N_21648,N_21475,N_21267);
and U21649 (N_21649,N_21385,N_21434);
nor U21650 (N_21650,N_21324,N_21284);
nor U21651 (N_21651,N_21282,N_21492);
nand U21652 (N_21652,N_21491,N_21374);
or U21653 (N_21653,N_21485,N_21340);
nand U21654 (N_21654,N_21474,N_21307);
nor U21655 (N_21655,N_21272,N_21284);
nor U21656 (N_21656,N_21279,N_21267);
nand U21657 (N_21657,N_21492,N_21388);
nand U21658 (N_21658,N_21376,N_21424);
nor U21659 (N_21659,N_21484,N_21374);
nor U21660 (N_21660,N_21343,N_21275);
nand U21661 (N_21661,N_21359,N_21408);
or U21662 (N_21662,N_21394,N_21424);
and U21663 (N_21663,N_21258,N_21429);
nor U21664 (N_21664,N_21354,N_21360);
and U21665 (N_21665,N_21475,N_21349);
and U21666 (N_21666,N_21425,N_21350);
or U21667 (N_21667,N_21388,N_21380);
or U21668 (N_21668,N_21374,N_21319);
nor U21669 (N_21669,N_21358,N_21277);
and U21670 (N_21670,N_21476,N_21466);
nand U21671 (N_21671,N_21361,N_21496);
and U21672 (N_21672,N_21351,N_21379);
or U21673 (N_21673,N_21295,N_21277);
nand U21674 (N_21674,N_21250,N_21432);
nand U21675 (N_21675,N_21292,N_21398);
or U21676 (N_21676,N_21314,N_21251);
nor U21677 (N_21677,N_21433,N_21478);
or U21678 (N_21678,N_21381,N_21426);
or U21679 (N_21679,N_21365,N_21264);
or U21680 (N_21680,N_21419,N_21452);
or U21681 (N_21681,N_21453,N_21397);
nand U21682 (N_21682,N_21458,N_21413);
and U21683 (N_21683,N_21332,N_21302);
or U21684 (N_21684,N_21405,N_21451);
or U21685 (N_21685,N_21470,N_21495);
and U21686 (N_21686,N_21418,N_21421);
and U21687 (N_21687,N_21375,N_21279);
nor U21688 (N_21688,N_21305,N_21262);
and U21689 (N_21689,N_21425,N_21472);
xor U21690 (N_21690,N_21417,N_21382);
or U21691 (N_21691,N_21367,N_21282);
and U21692 (N_21692,N_21348,N_21394);
nand U21693 (N_21693,N_21469,N_21370);
or U21694 (N_21694,N_21368,N_21381);
or U21695 (N_21695,N_21457,N_21437);
nor U21696 (N_21696,N_21420,N_21289);
nor U21697 (N_21697,N_21412,N_21315);
and U21698 (N_21698,N_21315,N_21284);
or U21699 (N_21699,N_21431,N_21336);
nor U21700 (N_21700,N_21401,N_21444);
and U21701 (N_21701,N_21281,N_21352);
nand U21702 (N_21702,N_21346,N_21471);
or U21703 (N_21703,N_21487,N_21428);
or U21704 (N_21704,N_21345,N_21286);
and U21705 (N_21705,N_21351,N_21349);
or U21706 (N_21706,N_21397,N_21322);
nor U21707 (N_21707,N_21414,N_21324);
nor U21708 (N_21708,N_21341,N_21393);
and U21709 (N_21709,N_21434,N_21498);
and U21710 (N_21710,N_21391,N_21447);
or U21711 (N_21711,N_21395,N_21358);
or U21712 (N_21712,N_21290,N_21259);
or U21713 (N_21713,N_21360,N_21369);
and U21714 (N_21714,N_21256,N_21303);
nand U21715 (N_21715,N_21400,N_21480);
nor U21716 (N_21716,N_21329,N_21460);
nor U21717 (N_21717,N_21261,N_21285);
nor U21718 (N_21718,N_21304,N_21435);
or U21719 (N_21719,N_21379,N_21483);
and U21720 (N_21720,N_21355,N_21283);
or U21721 (N_21721,N_21330,N_21341);
nand U21722 (N_21722,N_21440,N_21446);
and U21723 (N_21723,N_21375,N_21264);
and U21724 (N_21724,N_21310,N_21420);
nor U21725 (N_21725,N_21331,N_21361);
nand U21726 (N_21726,N_21444,N_21446);
and U21727 (N_21727,N_21424,N_21347);
and U21728 (N_21728,N_21284,N_21399);
and U21729 (N_21729,N_21262,N_21329);
nand U21730 (N_21730,N_21477,N_21325);
or U21731 (N_21731,N_21415,N_21343);
or U21732 (N_21732,N_21349,N_21353);
or U21733 (N_21733,N_21344,N_21375);
and U21734 (N_21734,N_21468,N_21459);
nor U21735 (N_21735,N_21353,N_21409);
nor U21736 (N_21736,N_21484,N_21495);
and U21737 (N_21737,N_21452,N_21290);
nand U21738 (N_21738,N_21298,N_21270);
nor U21739 (N_21739,N_21359,N_21278);
nand U21740 (N_21740,N_21414,N_21317);
and U21741 (N_21741,N_21339,N_21316);
nor U21742 (N_21742,N_21384,N_21255);
or U21743 (N_21743,N_21429,N_21403);
and U21744 (N_21744,N_21301,N_21390);
nor U21745 (N_21745,N_21357,N_21418);
or U21746 (N_21746,N_21414,N_21366);
nor U21747 (N_21747,N_21461,N_21377);
or U21748 (N_21748,N_21307,N_21264);
and U21749 (N_21749,N_21405,N_21446);
or U21750 (N_21750,N_21747,N_21678);
or U21751 (N_21751,N_21510,N_21583);
and U21752 (N_21752,N_21502,N_21738);
nor U21753 (N_21753,N_21689,N_21721);
and U21754 (N_21754,N_21637,N_21607);
and U21755 (N_21755,N_21735,N_21642);
nor U21756 (N_21756,N_21509,N_21670);
nand U21757 (N_21757,N_21596,N_21739);
or U21758 (N_21758,N_21620,N_21711);
and U21759 (N_21759,N_21547,N_21654);
nand U21760 (N_21760,N_21538,N_21543);
or U21761 (N_21761,N_21588,N_21591);
or U21762 (N_21762,N_21699,N_21665);
nor U21763 (N_21763,N_21575,N_21663);
nand U21764 (N_21764,N_21651,N_21594);
nand U21765 (N_21765,N_21707,N_21730);
nor U21766 (N_21766,N_21659,N_21568);
or U21767 (N_21767,N_21694,N_21649);
nor U21768 (N_21768,N_21504,N_21683);
and U21769 (N_21769,N_21718,N_21710);
and U21770 (N_21770,N_21644,N_21597);
or U21771 (N_21771,N_21517,N_21657);
nor U21772 (N_21772,N_21746,N_21674);
or U21773 (N_21773,N_21723,N_21539);
nand U21774 (N_21774,N_21586,N_21668);
nand U21775 (N_21775,N_21622,N_21650);
nor U21776 (N_21776,N_21574,N_21701);
and U21777 (N_21777,N_21673,N_21567);
nor U21778 (N_21778,N_21636,N_21566);
and U21779 (N_21779,N_21676,N_21605);
nor U21780 (N_21780,N_21514,N_21703);
nand U21781 (N_21781,N_21634,N_21688);
nor U21782 (N_21782,N_21684,N_21530);
or U21783 (N_21783,N_21598,N_21506);
and U21784 (N_21784,N_21742,N_21616);
or U21785 (N_21785,N_21508,N_21612);
nor U21786 (N_21786,N_21719,N_21615);
and U21787 (N_21787,N_21545,N_21706);
nand U21788 (N_21788,N_21600,N_21534);
and U21789 (N_21789,N_21695,N_21685);
nor U21790 (N_21790,N_21628,N_21696);
and U21791 (N_21791,N_21589,N_21648);
nor U21792 (N_21792,N_21516,N_21512);
and U21793 (N_21793,N_21617,N_21572);
nand U21794 (N_21794,N_21669,N_21546);
nor U21795 (N_21795,N_21520,N_21613);
nand U21796 (N_21796,N_21737,N_21677);
nand U21797 (N_21797,N_21700,N_21667);
and U21798 (N_21798,N_21533,N_21681);
and U21799 (N_21799,N_21671,N_21716);
nand U21800 (N_21800,N_21554,N_21741);
and U21801 (N_21801,N_21528,N_21560);
nand U21802 (N_21802,N_21578,N_21705);
and U21803 (N_21803,N_21527,N_21563);
or U21804 (N_21804,N_21725,N_21585);
and U21805 (N_21805,N_21631,N_21590);
nand U21806 (N_21806,N_21748,N_21724);
or U21807 (N_21807,N_21714,N_21555);
or U21808 (N_21808,N_21736,N_21556);
and U21809 (N_21809,N_21536,N_21732);
nor U21810 (N_21810,N_21561,N_21624);
nor U21811 (N_21811,N_21623,N_21733);
or U21812 (N_21812,N_21698,N_21690);
nor U21813 (N_21813,N_21569,N_21522);
xnor U21814 (N_21814,N_21728,N_21708);
nand U21815 (N_21815,N_21614,N_21571);
nor U21816 (N_21816,N_21603,N_21525);
nand U21817 (N_21817,N_21715,N_21749);
xor U21818 (N_21818,N_21601,N_21658);
or U21819 (N_21819,N_21579,N_21515);
and U21820 (N_21820,N_21519,N_21672);
nor U21821 (N_21821,N_21505,N_21626);
nor U21822 (N_21822,N_21645,N_21576);
nand U21823 (N_21823,N_21661,N_21544);
or U21824 (N_21824,N_21702,N_21584);
nor U21825 (N_21825,N_21581,N_21662);
and U21826 (N_21826,N_21744,N_21604);
nand U21827 (N_21827,N_21666,N_21635);
and U21828 (N_21828,N_21608,N_21712);
or U21829 (N_21829,N_21686,N_21557);
nand U21830 (N_21830,N_21691,N_21729);
and U21831 (N_21831,N_21619,N_21646);
or U21832 (N_21832,N_21565,N_21523);
nor U21833 (N_21833,N_21518,N_21580);
xor U21834 (N_21834,N_21592,N_21629);
nor U21835 (N_21835,N_21679,N_21611);
or U21836 (N_21836,N_21656,N_21507);
nand U21837 (N_21837,N_21664,N_21549);
or U21838 (N_21838,N_21550,N_21660);
xnor U21839 (N_21839,N_21731,N_21529);
nor U21840 (N_21840,N_21501,N_21675);
or U21841 (N_21841,N_21693,N_21599);
nand U21842 (N_21842,N_21524,N_21734);
or U21843 (N_21843,N_21602,N_21652);
and U21844 (N_21844,N_21521,N_21541);
nand U21845 (N_21845,N_21542,N_21513);
or U21846 (N_21846,N_21717,N_21641);
nor U21847 (N_21847,N_21627,N_21593);
nor U21848 (N_21848,N_21595,N_21639);
or U21849 (N_21849,N_21720,N_21535);
nor U21850 (N_21850,N_21537,N_21552);
xor U21851 (N_21851,N_21532,N_21638);
or U21852 (N_21852,N_21562,N_21697);
nor U21853 (N_21853,N_21726,N_21621);
or U21854 (N_21854,N_21680,N_21573);
nor U21855 (N_21855,N_21609,N_21618);
nor U21856 (N_21856,N_21587,N_21606);
nand U21857 (N_21857,N_21540,N_21643);
nand U21858 (N_21858,N_21511,N_21500);
nor U21859 (N_21859,N_21727,N_21553);
and U21860 (N_21860,N_21577,N_21655);
nand U21861 (N_21861,N_21558,N_21526);
or U21862 (N_21862,N_21503,N_21709);
nand U21863 (N_21863,N_21704,N_21740);
and U21864 (N_21864,N_21713,N_21625);
or U21865 (N_21865,N_21632,N_21531);
nand U21866 (N_21866,N_21610,N_21745);
nand U21867 (N_21867,N_21722,N_21548);
nand U21868 (N_21868,N_21582,N_21692);
nor U21869 (N_21869,N_21570,N_21633);
nand U21870 (N_21870,N_21564,N_21653);
nand U21871 (N_21871,N_21630,N_21640);
nor U21872 (N_21872,N_21551,N_21559);
and U21873 (N_21873,N_21682,N_21647);
nand U21874 (N_21874,N_21743,N_21687);
or U21875 (N_21875,N_21688,N_21534);
nand U21876 (N_21876,N_21676,N_21626);
or U21877 (N_21877,N_21740,N_21609);
or U21878 (N_21878,N_21697,N_21513);
or U21879 (N_21879,N_21683,N_21715);
nor U21880 (N_21880,N_21661,N_21749);
and U21881 (N_21881,N_21580,N_21601);
or U21882 (N_21882,N_21652,N_21512);
nand U21883 (N_21883,N_21544,N_21568);
nor U21884 (N_21884,N_21523,N_21603);
nor U21885 (N_21885,N_21653,N_21703);
and U21886 (N_21886,N_21635,N_21742);
and U21887 (N_21887,N_21592,N_21677);
nor U21888 (N_21888,N_21749,N_21581);
nor U21889 (N_21889,N_21552,N_21555);
and U21890 (N_21890,N_21552,N_21663);
and U21891 (N_21891,N_21689,N_21533);
or U21892 (N_21892,N_21523,N_21633);
xnor U21893 (N_21893,N_21628,N_21675);
or U21894 (N_21894,N_21622,N_21530);
nor U21895 (N_21895,N_21608,N_21672);
and U21896 (N_21896,N_21636,N_21715);
and U21897 (N_21897,N_21572,N_21660);
or U21898 (N_21898,N_21624,N_21573);
and U21899 (N_21899,N_21700,N_21726);
nand U21900 (N_21900,N_21748,N_21532);
nand U21901 (N_21901,N_21642,N_21502);
or U21902 (N_21902,N_21583,N_21595);
or U21903 (N_21903,N_21532,N_21609);
nand U21904 (N_21904,N_21647,N_21658);
or U21905 (N_21905,N_21732,N_21516);
nor U21906 (N_21906,N_21726,N_21598);
or U21907 (N_21907,N_21681,N_21731);
or U21908 (N_21908,N_21587,N_21588);
nor U21909 (N_21909,N_21620,N_21653);
nand U21910 (N_21910,N_21726,N_21652);
and U21911 (N_21911,N_21649,N_21511);
and U21912 (N_21912,N_21740,N_21566);
nand U21913 (N_21913,N_21523,N_21503);
or U21914 (N_21914,N_21735,N_21584);
or U21915 (N_21915,N_21725,N_21688);
and U21916 (N_21916,N_21649,N_21544);
nor U21917 (N_21917,N_21602,N_21576);
nand U21918 (N_21918,N_21610,N_21615);
or U21919 (N_21919,N_21625,N_21565);
and U21920 (N_21920,N_21583,N_21615);
nand U21921 (N_21921,N_21720,N_21570);
or U21922 (N_21922,N_21749,N_21731);
or U21923 (N_21923,N_21590,N_21646);
and U21924 (N_21924,N_21592,N_21602);
nand U21925 (N_21925,N_21614,N_21509);
nor U21926 (N_21926,N_21690,N_21667);
or U21927 (N_21927,N_21696,N_21735);
nor U21928 (N_21928,N_21604,N_21535);
nand U21929 (N_21929,N_21525,N_21660);
nand U21930 (N_21930,N_21611,N_21571);
nor U21931 (N_21931,N_21746,N_21510);
nor U21932 (N_21932,N_21525,N_21527);
nor U21933 (N_21933,N_21502,N_21650);
nor U21934 (N_21934,N_21519,N_21622);
and U21935 (N_21935,N_21510,N_21630);
nor U21936 (N_21936,N_21605,N_21653);
and U21937 (N_21937,N_21522,N_21591);
nand U21938 (N_21938,N_21534,N_21663);
and U21939 (N_21939,N_21513,N_21516);
and U21940 (N_21940,N_21714,N_21533);
nand U21941 (N_21941,N_21725,N_21650);
and U21942 (N_21942,N_21552,N_21548);
nand U21943 (N_21943,N_21519,N_21529);
nor U21944 (N_21944,N_21578,N_21742);
or U21945 (N_21945,N_21596,N_21627);
and U21946 (N_21946,N_21580,N_21598);
nor U21947 (N_21947,N_21702,N_21510);
and U21948 (N_21948,N_21553,N_21638);
nor U21949 (N_21949,N_21705,N_21589);
nor U21950 (N_21950,N_21696,N_21639);
nand U21951 (N_21951,N_21513,N_21636);
or U21952 (N_21952,N_21641,N_21671);
and U21953 (N_21953,N_21692,N_21691);
and U21954 (N_21954,N_21695,N_21586);
and U21955 (N_21955,N_21649,N_21705);
or U21956 (N_21956,N_21634,N_21670);
and U21957 (N_21957,N_21534,N_21721);
nor U21958 (N_21958,N_21635,N_21537);
and U21959 (N_21959,N_21619,N_21513);
nor U21960 (N_21960,N_21742,N_21590);
nand U21961 (N_21961,N_21686,N_21714);
nand U21962 (N_21962,N_21709,N_21663);
and U21963 (N_21963,N_21659,N_21717);
nor U21964 (N_21964,N_21574,N_21576);
nor U21965 (N_21965,N_21721,N_21676);
nand U21966 (N_21966,N_21535,N_21710);
or U21967 (N_21967,N_21562,N_21503);
nor U21968 (N_21968,N_21661,N_21715);
nor U21969 (N_21969,N_21521,N_21675);
nand U21970 (N_21970,N_21697,N_21579);
and U21971 (N_21971,N_21718,N_21605);
nor U21972 (N_21972,N_21692,N_21503);
and U21973 (N_21973,N_21746,N_21665);
or U21974 (N_21974,N_21623,N_21742);
or U21975 (N_21975,N_21636,N_21556);
and U21976 (N_21976,N_21530,N_21657);
and U21977 (N_21977,N_21541,N_21734);
or U21978 (N_21978,N_21698,N_21625);
nand U21979 (N_21979,N_21657,N_21535);
nor U21980 (N_21980,N_21531,N_21519);
nand U21981 (N_21981,N_21648,N_21603);
nor U21982 (N_21982,N_21625,N_21634);
nor U21983 (N_21983,N_21743,N_21536);
or U21984 (N_21984,N_21726,N_21563);
nand U21985 (N_21985,N_21559,N_21524);
nor U21986 (N_21986,N_21687,N_21737);
nand U21987 (N_21987,N_21508,N_21539);
nor U21988 (N_21988,N_21585,N_21532);
or U21989 (N_21989,N_21676,N_21515);
and U21990 (N_21990,N_21730,N_21565);
and U21991 (N_21991,N_21667,N_21727);
and U21992 (N_21992,N_21644,N_21593);
and U21993 (N_21993,N_21613,N_21553);
nor U21994 (N_21994,N_21652,N_21735);
or U21995 (N_21995,N_21650,N_21617);
and U21996 (N_21996,N_21525,N_21720);
nor U21997 (N_21997,N_21719,N_21597);
nand U21998 (N_21998,N_21725,N_21601);
nand U21999 (N_21999,N_21517,N_21669);
nor U22000 (N_22000,N_21970,N_21947);
or U22001 (N_22001,N_21792,N_21773);
and U22002 (N_22002,N_21956,N_21924);
and U22003 (N_22003,N_21759,N_21819);
or U22004 (N_22004,N_21876,N_21920);
nor U22005 (N_22005,N_21941,N_21841);
or U22006 (N_22006,N_21969,N_21968);
nand U22007 (N_22007,N_21880,N_21774);
or U22008 (N_22008,N_21788,N_21828);
nand U22009 (N_22009,N_21755,N_21972);
or U22010 (N_22010,N_21952,N_21764);
and U22011 (N_22011,N_21845,N_21900);
or U22012 (N_22012,N_21894,N_21959);
or U22013 (N_22013,N_21975,N_21884);
and U22014 (N_22014,N_21929,N_21987);
nor U22015 (N_22015,N_21800,N_21766);
nand U22016 (N_22016,N_21901,N_21862);
or U22017 (N_22017,N_21937,N_21855);
or U22018 (N_22018,N_21878,N_21754);
nor U22019 (N_22019,N_21958,N_21799);
nand U22020 (N_22020,N_21820,N_21810);
nor U22021 (N_22021,N_21981,N_21818);
nor U22022 (N_22022,N_21778,N_21756);
and U22023 (N_22023,N_21775,N_21921);
and U22024 (N_22024,N_21886,N_21791);
nor U22025 (N_22025,N_21860,N_21893);
nand U22026 (N_22026,N_21814,N_21967);
nor U22027 (N_22027,N_21837,N_21945);
nand U22028 (N_22028,N_21783,N_21846);
and U22029 (N_22029,N_21848,N_21892);
or U22030 (N_22030,N_21903,N_21888);
or U22031 (N_22031,N_21808,N_21962);
and U22032 (N_22032,N_21809,N_21827);
and U22033 (N_22033,N_21912,N_21861);
or U22034 (N_22034,N_21785,N_21798);
and U22035 (N_22035,N_21789,N_21939);
nand U22036 (N_22036,N_21770,N_21872);
nand U22037 (N_22037,N_21781,N_21832);
nor U22038 (N_22038,N_21935,N_21866);
nand U22039 (N_22039,N_21913,N_21856);
or U22040 (N_22040,N_21768,N_21990);
nor U22041 (N_22041,N_21836,N_21905);
nand U22042 (N_22042,N_21867,N_21907);
nor U22043 (N_22043,N_21964,N_21854);
and U22044 (N_22044,N_21923,N_21853);
nor U22045 (N_22045,N_21915,N_21927);
or U22046 (N_22046,N_21925,N_21869);
nand U22047 (N_22047,N_21833,N_21896);
nor U22048 (N_22048,N_21991,N_21851);
and U22049 (N_22049,N_21988,N_21843);
or U22050 (N_22050,N_21950,N_21931);
nand U22051 (N_22051,N_21859,N_21909);
nand U22052 (N_22052,N_21976,N_21993);
nand U22053 (N_22053,N_21813,N_21839);
or U22054 (N_22054,N_21954,N_21812);
and U22055 (N_22055,N_21961,N_21895);
or U22056 (N_22056,N_21807,N_21918);
nor U22057 (N_22057,N_21890,N_21863);
nand U22058 (N_22058,N_21877,N_21752);
or U22059 (N_22059,N_21994,N_21995);
nor U22060 (N_22060,N_21948,N_21889);
and U22061 (N_22061,N_21771,N_21883);
or U22062 (N_22062,N_21762,N_21999);
nor U22063 (N_22063,N_21955,N_21760);
or U22064 (N_22064,N_21917,N_21758);
or U22065 (N_22065,N_21902,N_21757);
and U22066 (N_22066,N_21897,N_21767);
or U22067 (N_22067,N_21934,N_21782);
nand U22068 (N_22068,N_21787,N_21780);
and U22069 (N_22069,N_21986,N_21858);
nand U22070 (N_22070,N_21891,N_21944);
nor U22071 (N_22071,N_21942,N_21777);
or U22072 (N_22072,N_21911,N_21761);
and U22073 (N_22073,N_21849,N_21802);
and U22074 (N_22074,N_21772,N_21831);
nor U22075 (N_22075,N_21879,N_21885);
or U22076 (N_22076,N_21838,N_21795);
or U22077 (N_22077,N_21823,N_21984);
and U22078 (N_22078,N_21992,N_21974);
nand U22079 (N_22079,N_21870,N_21864);
nor U22080 (N_22080,N_21973,N_21805);
nor U22081 (N_22081,N_21763,N_21835);
and U22082 (N_22082,N_21834,N_21936);
or U22083 (N_22083,N_21922,N_21830);
nand U22084 (N_22084,N_21978,N_21857);
and U22085 (N_22085,N_21804,N_21998);
nor U22086 (N_22086,N_21906,N_21882);
nand U22087 (N_22087,N_21914,N_21957);
and U22088 (N_22088,N_21908,N_21904);
or U22089 (N_22089,N_21997,N_21801);
nand U22090 (N_22090,N_21815,N_21868);
nor U22091 (N_22091,N_21769,N_21806);
or U22092 (N_22092,N_21951,N_21874);
and U22093 (N_22093,N_21817,N_21946);
or U22094 (N_22094,N_21811,N_21933);
or U22095 (N_22095,N_21982,N_21928);
nor U22096 (N_22096,N_21985,N_21847);
nor U22097 (N_22097,N_21963,N_21793);
nor U22098 (N_22098,N_21751,N_21794);
nand U22099 (N_22099,N_21949,N_21887);
nor U22100 (N_22100,N_21797,N_21824);
and U22101 (N_22101,N_21786,N_21871);
nor U22102 (N_22102,N_21996,N_21926);
and U22103 (N_22103,N_21776,N_21852);
and U22104 (N_22104,N_21796,N_21980);
or U22105 (N_22105,N_21919,N_21932);
or U22106 (N_22106,N_21881,N_21873);
or U22107 (N_22107,N_21753,N_21790);
and U22108 (N_22108,N_21979,N_21750);
and U22109 (N_22109,N_21765,N_21816);
nor U22110 (N_22110,N_21938,N_21898);
and U22111 (N_22111,N_21875,N_21865);
nand U22112 (N_22112,N_21953,N_21784);
nor U22113 (N_22113,N_21826,N_21977);
and U22114 (N_22114,N_21930,N_21822);
or U22115 (N_22115,N_21971,N_21910);
or U22116 (N_22116,N_21989,N_21844);
and U22117 (N_22117,N_21821,N_21965);
or U22118 (N_22118,N_21960,N_21829);
nor U22119 (N_22119,N_21899,N_21803);
xnor U22120 (N_22120,N_21850,N_21983);
nand U22121 (N_22121,N_21943,N_21916);
and U22122 (N_22122,N_21779,N_21842);
or U22123 (N_22123,N_21825,N_21840);
nor U22124 (N_22124,N_21940,N_21966);
and U22125 (N_22125,N_21903,N_21784);
or U22126 (N_22126,N_21984,N_21991);
or U22127 (N_22127,N_21857,N_21886);
nand U22128 (N_22128,N_21941,N_21907);
nand U22129 (N_22129,N_21965,N_21872);
nor U22130 (N_22130,N_21978,N_21828);
nand U22131 (N_22131,N_21949,N_21919);
and U22132 (N_22132,N_21973,N_21783);
nor U22133 (N_22133,N_21898,N_21869);
nor U22134 (N_22134,N_21861,N_21785);
and U22135 (N_22135,N_21868,N_21800);
nand U22136 (N_22136,N_21914,N_21834);
nor U22137 (N_22137,N_21788,N_21997);
or U22138 (N_22138,N_21928,N_21962);
nand U22139 (N_22139,N_21767,N_21860);
nand U22140 (N_22140,N_21826,N_21769);
nand U22141 (N_22141,N_21878,N_21800);
xor U22142 (N_22142,N_21843,N_21879);
and U22143 (N_22143,N_21898,N_21774);
nor U22144 (N_22144,N_21993,N_21956);
xor U22145 (N_22145,N_21810,N_21933);
or U22146 (N_22146,N_21981,N_21942);
nor U22147 (N_22147,N_21786,N_21887);
and U22148 (N_22148,N_21877,N_21763);
and U22149 (N_22149,N_21884,N_21971);
nor U22150 (N_22150,N_21989,N_21767);
nor U22151 (N_22151,N_21770,N_21885);
nor U22152 (N_22152,N_21891,N_21825);
or U22153 (N_22153,N_21905,N_21782);
or U22154 (N_22154,N_21922,N_21829);
nand U22155 (N_22155,N_21876,N_21902);
nor U22156 (N_22156,N_21970,N_21827);
or U22157 (N_22157,N_21968,N_21903);
and U22158 (N_22158,N_21776,N_21884);
nand U22159 (N_22159,N_21982,N_21841);
and U22160 (N_22160,N_21861,N_21982);
and U22161 (N_22161,N_21818,N_21996);
and U22162 (N_22162,N_21913,N_21932);
and U22163 (N_22163,N_21765,N_21962);
nor U22164 (N_22164,N_21910,N_21887);
nand U22165 (N_22165,N_21858,N_21894);
nand U22166 (N_22166,N_21768,N_21819);
nor U22167 (N_22167,N_21919,N_21903);
and U22168 (N_22168,N_21937,N_21801);
and U22169 (N_22169,N_21823,N_21779);
and U22170 (N_22170,N_21786,N_21866);
and U22171 (N_22171,N_21839,N_21952);
and U22172 (N_22172,N_21822,N_21866);
nand U22173 (N_22173,N_21796,N_21820);
and U22174 (N_22174,N_21908,N_21765);
and U22175 (N_22175,N_21932,N_21958);
or U22176 (N_22176,N_21998,N_21820);
and U22177 (N_22177,N_21765,N_21978);
nor U22178 (N_22178,N_21930,N_21818);
nor U22179 (N_22179,N_21842,N_21763);
nand U22180 (N_22180,N_21873,N_21941);
nand U22181 (N_22181,N_21768,N_21760);
nand U22182 (N_22182,N_21945,N_21825);
nand U22183 (N_22183,N_21947,N_21800);
or U22184 (N_22184,N_21878,N_21923);
nor U22185 (N_22185,N_21848,N_21768);
nor U22186 (N_22186,N_21938,N_21765);
and U22187 (N_22187,N_21987,N_21784);
nand U22188 (N_22188,N_21987,N_21867);
or U22189 (N_22189,N_21981,N_21823);
and U22190 (N_22190,N_21867,N_21768);
nand U22191 (N_22191,N_21815,N_21877);
nand U22192 (N_22192,N_21928,N_21915);
and U22193 (N_22193,N_21837,N_21896);
and U22194 (N_22194,N_21941,N_21829);
nor U22195 (N_22195,N_21977,N_21841);
and U22196 (N_22196,N_21933,N_21792);
and U22197 (N_22197,N_21898,N_21756);
or U22198 (N_22198,N_21939,N_21988);
nor U22199 (N_22199,N_21790,N_21886);
or U22200 (N_22200,N_21850,N_21765);
nor U22201 (N_22201,N_21874,N_21771);
nand U22202 (N_22202,N_21850,N_21787);
nor U22203 (N_22203,N_21997,N_21987);
nand U22204 (N_22204,N_21888,N_21972);
nand U22205 (N_22205,N_21762,N_21803);
or U22206 (N_22206,N_21855,N_21812);
and U22207 (N_22207,N_21897,N_21878);
nor U22208 (N_22208,N_21907,N_21856);
nand U22209 (N_22209,N_21773,N_21882);
nand U22210 (N_22210,N_21897,N_21794);
and U22211 (N_22211,N_21769,N_21816);
or U22212 (N_22212,N_21880,N_21893);
nor U22213 (N_22213,N_21968,N_21795);
or U22214 (N_22214,N_21922,N_21834);
or U22215 (N_22215,N_21864,N_21838);
nand U22216 (N_22216,N_21900,N_21908);
nand U22217 (N_22217,N_21812,N_21815);
nor U22218 (N_22218,N_21792,N_21769);
nor U22219 (N_22219,N_21864,N_21753);
nand U22220 (N_22220,N_21858,N_21969);
xnor U22221 (N_22221,N_21854,N_21821);
and U22222 (N_22222,N_21940,N_21884);
and U22223 (N_22223,N_21785,N_21796);
nand U22224 (N_22224,N_21861,N_21990);
nand U22225 (N_22225,N_21799,N_21918);
or U22226 (N_22226,N_21879,N_21765);
nand U22227 (N_22227,N_21886,N_21793);
nand U22228 (N_22228,N_21943,N_21965);
and U22229 (N_22229,N_21833,N_21878);
or U22230 (N_22230,N_21962,N_21986);
nand U22231 (N_22231,N_21989,N_21818);
nor U22232 (N_22232,N_21788,N_21947);
nand U22233 (N_22233,N_21835,N_21955);
and U22234 (N_22234,N_21779,N_21792);
and U22235 (N_22235,N_21958,N_21888);
or U22236 (N_22236,N_21972,N_21981);
or U22237 (N_22237,N_21799,N_21959);
or U22238 (N_22238,N_21887,N_21799);
or U22239 (N_22239,N_21779,N_21829);
or U22240 (N_22240,N_21967,N_21795);
nor U22241 (N_22241,N_21752,N_21952);
nor U22242 (N_22242,N_21886,N_21788);
and U22243 (N_22243,N_21885,N_21952);
nor U22244 (N_22244,N_21912,N_21786);
nor U22245 (N_22245,N_21894,N_21768);
or U22246 (N_22246,N_21779,N_21899);
and U22247 (N_22247,N_21960,N_21979);
and U22248 (N_22248,N_21879,N_21996);
nand U22249 (N_22249,N_21848,N_21959);
or U22250 (N_22250,N_22164,N_22154);
nand U22251 (N_22251,N_22069,N_22249);
and U22252 (N_22252,N_22059,N_22063);
nand U22253 (N_22253,N_22028,N_22090);
and U22254 (N_22254,N_22165,N_22212);
nor U22255 (N_22255,N_22171,N_22104);
or U22256 (N_22256,N_22129,N_22246);
nor U22257 (N_22257,N_22117,N_22032);
and U22258 (N_22258,N_22210,N_22177);
or U22259 (N_22259,N_22141,N_22087);
nand U22260 (N_22260,N_22030,N_22079);
and U22261 (N_22261,N_22189,N_22005);
and U22262 (N_22262,N_22179,N_22060);
or U22263 (N_22263,N_22245,N_22144);
or U22264 (N_22264,N_22248,N_22176);
or U22265 (N_22265,N_22233,N_22197);
nor U22266 (N_22266,N_22035,N_22068);
or U22267 (N_22267,N_22206,N_22088);
and U22268 (N_22268,N_22053,N_22092);
nand U22269 (N_22269,N_22225,N_22103);
or U22270 (N_22270,N_22124,N_22222);
and U22271 (N_22271,N_22123,N_22198);
or U22272 (N_22272,N_22047,N_22058);
and U22273 (N_22273,N_22169,N_22247);
and U22274 (N_22274,N_22099,N_22007);
nor U22275 (N_22275,N_22105,N_22094);
or U22276 (N_22276,N_22037,N_22242);
nor U22277 (N_22277,N_22076,N_22102);
or U22278 (N_22278,N_22056,N_22220);
or U22279 (N_22279,N_22033,N_22082);
nor U22280 (N_22280,N_22119,N_22193);
and U22281 (N_22281,N_22025,N_22050);
or U22282 (N_22282,N_22042,N_22113);
or U22283 (N_22283,N_22041,N_22009);
nand U22284 (N_22284,N_22024,N_22133);
nand U22285 (N_22285,N_22150,N_22223);
or U22286 (N_22286,N_22192,N_22040);
and U22287 (N_22287,N_22095,N_22004);
nand U22288 (N_22288,N_22071,N_22039);
or U22289 (N_22289,N_22203,N_22089);
and U22290 (N_22290,N_22204,N_22235);
nor U22291 (N_22291,N_22110,N_22074);
or U22292 (N_22292,N_22085,N_22116);
nand U22293 (N_22293,N_22243,N_22158);
nor U22294 (N_22294,N_22013,N_22127);
nand U22295 (N_22295,N_22010,N_22178);
nor U22296 (N_22296,N_22021,N_22145);
and U22297 (N_22297,N_22211,N_22077);
or U22298 (N_22298,N_22240,N_22136);
or U22299 (N_22299,N_22126,N_22143);
or U22300 (N_22300,N_22062,N_22147);
xor U22301 (N_22301,N_22016,N_22208);
nor U22302 (N_22302,N_22006,N_22221);
and U22303 (N_22303,N_22148,N_22234);
and U22304 (N_22304,N_22218,N_22086);
and U22305 (N_22305,N_22084,N_22167);
nor U22306 (N_22306,N_22049,N_22029);
and U22307 (N_22307,N_22114,N_22201);
and U22308 (N_22308,N_22231,N_22186);
or U22309 (N_22309,N_22140,N_22236);
and U22310 (N_22310,N_22217,N_22188);
and U22311 (N_22311,N_22151,N_22051);
nor U22312 (N_22312,N_22230,N_22213);
nor U22313 (N_22313,N_22057,N_22239);
nand U22314 (N_22314,N_22142,N_22020);
nand U22315 (N_22315,N_22215,N_22160);
and U22316 (N_22316,N_22112,N_22111);
or U22317 (N_22317,N_22080,N_22012);
or U22318 (N_22318,N_22159,N_22115);
nor U22319 (N_22319,N_22044,N_22043);
nor U22320 (N_22320,N_22138,N_22139);
nand U22321 (N_22321,N_22034,N_22216);
or U22322 (N_22322,N_22070,N_22132);
or U22323 (N_22323,N_22023,N_22214);
nand U22324 (N_22324,N_22135,N_22199);
or U22325 (N_22325,N_22194,N_22001);
nand U22326 (N_22326,N_22002,N_22081);
nor U22327 (N_22327,N_22046,N_22128);
and U22328 (N_22328,N_22134,N_22196);
nor U22329 (N_22329,N_22232,N_22026);
or U22330 (N_22330,N_22219,N_22075);
and U22331 (N_22331,N_22054,N_22064);
nor U22332 (N_22332,N_22195,N_22008);
nor U22333 (N_22333,N_22022,N_22120);
and U22334 (N_22334,N_22187,N_22066);
and U22335 (N_22335,N_22118,N_22055);
nor U22336 (N_22336,N_22202,N_22162);
nand U22337 (N_22337,N_22163,N_22183);
nand U22338 (N_22338,N_22172,N_22153);
and U22339 (N_22339,N_22067,N_22241);
or U22340 (N_22340,N_22036,N_22238);
nand U22341 (N_22341,N_22149,N_22166);
nor U22342 (N_22342,N_22122,N_22237);
and U22343 (N_22343,N_22106,N_22107);
nor U22344 (N_22344,N_22000,N_22018);
or U22345 (N_22345,N_22011,N_22228);
nor U22346 (N_22346,N_22181,N_22027);
nand U22347 (N_22347,N_22146,N_22096);
nor U22348 (N_22348,N_22207,N_22173);
nor U22349 (N_22349,N_22014,N_22038);
and U22350 (N_22350,N_22155,N_22168);
nand U22351 (N_22351,N_22078,N_22061);
nor U22352 (N_22352,N_22048,N_22065);
nand U22353 (N_22353,N_22152,N_22161);
or U22354 (N_22354,N_22100,N_22244);
nand U22355 (N_22355,N_22180,N_22015);
nor U22356 (N_22356,N_22200,N_22184);
and U22357 (N_22357,N_22073,N_22229);
nor U22358 (N_22358,N_22174,N_22108);
and U22359 (N_22359,N_22072,N_22101);
nand U22360 (N_22360,N_22083,N_22205);
or U22361 (N_22361,N_22045,N_22224);
nand U22362 (N_22362,N_22031,N_22190);
or U22363 (N_22363,N_22017,N_22182);
nor U22364 (N_22364,N_22209,N_22097);
nor U22365 (N_22365,N_22003,N_22052);
or U22366 (N_22366,N_22226,N_22130);
nand U22367 (N_22367,N_22098,N_22175);
nor U22368 (N_22368,N_22191,N_22019);
nor U22369 (N_22369,N_22131,N_22227);
or U22370 (N_22370,N_22125,N_22121);
or U22371 (N_22371,N_22185,N_22091);
and U22372 (N_22372,N_22157,N_22109);
and U22373 (N_22373,N_22137,N_22156);
and U22374 (N_22374,N_22093,N_22170);
nor U22375 (N_22375,N_22120,N_22021);
and U22376 (N_22376,N_22241,N_22072);
nor U22377 (N_22377,N_22058,N_22012);
and U22378 (N_22378,N_22049,N_22105);
and U22379 (N_22379,N_22046,N_22026);
or U22380 (N_22380,N_22182,N_22124);
nand U22381 (N_22381,N_22049,N_22180);
and U22382 (N_22382,N_22237,N_22025);
nor U22383 (N_22383,N_22145,N_22089);
nor U22384 (N_22384,N_22009,N_22107);
nor U22385 (N_22385,N_22171,N_22112);
nand U22386 (N_22386,N_22236,N_22219);
nand U22387 (N_22387,N_22114,N_22124);
or U22388 (N_22388,N_22222,N_22041);
nand U22389 (N_22389,N_22072,N_22164);
nand U22390 (N_22390,N_22218,N_22095);
or U22391 (N_22391,N_22022,N_22198);
nand U22392 (N_22392,N_22118,N_22085);
and U22393 (N_22393,N_22028,N_22136);
nand U22394 (N_22394,N_22245,N_22101);
nor U22395 (N_22395,N_22105,N_22006);
nor U22396 (N_22396,N_22221,N_22208);
or U22397 (N_22397,N_22106,N_22138);
and U22398 (N_22398,N_22200,N_22033);
nand U22399 (N_22399,N_22022,N_22065);
nor U22400 (N_22400,N_22131,N_22171);
or U22401 (N_22401,N_22208,N_22005);
and U22402 (N_22402,N_22101,N_22096);
nor U22403 (N_22403,N_22131,N_22052);
nor U22404 (N_22404,N_22083,N_22125);
nand U22405 (N_22405,N_22136,N_22171);
and U22406 (N_22406,N_22126,N_22009);
nand U22407 (N_22407,N_22072,N_22243);
and U22408 (N_22408,N_22042,N_22097);
nor U22409 (N_22409,N_22001,N_22094);
nand U22410 (N_22410,N_22169,N_22064);
nor U22411 (N_22411,N_22006,N_22204);
nor U22412 (N_22412,N_22057,N_22204);
or U22413 (N_22413,N_22069,N_22106);
or U22414 (N_22414,N_22049,N_22185);
nor U22415 (N_22415,N_22052,N_22139);
nor U22416 (N_22416,N_22217,N_22227);
nand U22417 (N_22417,N_22172,N_22079);
or U22418 (N_22418,N_22076,N_22031);
and U22419 (N_22419,N_22123,N_22103);
or U22420 (N_22420,N_22174,N_22161);
or U22421 (N_22421,N_22104,N_22205);
or U22422 (N_22422,N_22067,N_22151);
nor U22423 (N_22423,N_22116,N_22005);
nor U22424 (N_22424,N_22215,N_22093);
nand U22425 (N_22425,N_22037,N_22000);
or U22426 (N_22426,N_22194,N_22098);
or U22427 (N_22427,N_22211,N_22198);
or U22428 (N_22428,N_22117,N_22148);
or U22429 (N_22429,N_22051,N_22136);
or U22430 (N_22430,N_22085,N_22208);
nor U22431 (N_22431,N_22240,N_22092);
and U22432 (N_22432,N_22226,N_22092);
xnor U22433 (N_22433,N_22119,N_22059);
and U22434 (N_22434,N_22108,N_22039);
nor U22435 (N_22435,N_22130,N_22118);
or U22436 (N_22436,N_22080,N_22164);
nand U22437 (N_22437,N_22180,N_22057);
or U22438 (N_22438,N_22180,N_22029);
nor U22439 (N_22439,N_22127,N_22103);
or U22440 (N_22440,N_22239,N_22217);
and U22441 (N_22441,N_22198,N_22133);
or U22442 (N_22442,N_22174,N_22195);
or U22443 (N_22443,N_22088,N_22022);
and U22444 (N_22444,N_22092,N_22198);
or U22445 (N_22445,N_22144,N_22140);
or U22446 (N_22446,N_22246,N_22143);
nor U22447 (N_22447,N_22003,N_22095);
or U22448 (N_22448,N_22181,N_22023);
and U22449 (N_22449,N_22146,N_22076);
nand U22450 (N_22450,N_22030,N_22152);
or U22451 (N_22451,N_22181,N_22235);
or U22452 (N_22452,N_22211,N_22249);
or U22453 (N_22453,N_22068,N_22071);
nand U22454 (N_22454,N_22213,N_22040);
or U22455 (N_22455,N_22168,N_22058);
nand U22456 (N_22456,N_22049,N_22205);
or U22457 (N_22457,N_22116,N_22191);
nand U22458 (N_22458,N_22194,N_22085);
or U22459 (N_22459,N_22143,N_22132);
or U22460 (N_22460,N_22210,N_22042);
or U22461 (N_22461,N_22080,N_22121);
and U22462 (N_22462,N_22205,N_22059);
nor U22463 (N_22463,N_22100,N_22217);
nand U22464 (N_22464,N_22200,N_22027);
nor U22465 (N_22465,N_22168,N_22025);
or U22466 (N_22466,N_22237,N_22247);
or U22467 (N_22467,N_22009,N_22246);
nor U22468 (N_22468,N_22171,N_22140);
nand U22469 (N_22469,N_22196,N_22067);
nand U22470 (N_22470,N_22202,N_22078);
nand U22471 (N_22471,N_22123,N_22134);
nor U22472 (N_22472,N_22072,N_22153);
nand U22473 (N_22473,N_22188,N_22007);
nand U22474 (N_22474,N_22131,N_22069);
nand U22475 (N_22475,N_22042,N_22194);
nor U22476 (N_22476,N_22200,N_22199);
nand U22477 (N_22477,N_22234,N_22199);
nor U22478 (N_22478,N_22092,N_22178);
and U22479 (N_22479,N_22137,N_22146);
or U22480 (N_22480,N_22198,N_22013);
and U22481 (N_22481,N_22102,N_22239);
nor U22482 (N_22482,N_22217,N_22249);
and U22483 (N_22483,N_22065,N_22075);
and U22484 (N_22484,N_22031,N_22211);
and U22485 (N_22485,N_22035,N_22124);
nor U22486 (N_22486,N_22126,N_22108);
or U22487 (N_22487,N_22245,N_22200);
and U22488 (N_22488,N_22047,N_22024);
nor U22489 (N_22489,N_22088,N_22124);
and U22490 (N_22490,N_22022,N_22053);
or U22491 (N_22491,N_22030,N_22049);
and U22492 (N_22492,N_22073,N_22061);
nand U22493 (N_22493,N_22094,N_22240);
nand U22494 (N_22494,N_22029,N_22168);
or U22495 (N_22495,N_22009,N_22185);
nand U22496 (N_22496,N_22164,N_22167);
or U22497 (N_22497,N_22153,N_22219);
or U22498 (N_22498,N_22130,N_22027);
or U22499 (N_22499,N_22095,N_22207);
or U22500 (N_22500,N_22432,N_22405);
nand U22501 (N_22501,N_22366,N_22499);
nor U22502 (N_22502,N_22253,N_22357);
nor U22503 (N_22503,N_22483,N_22462);
and U22504 (N_22504,N_22303,N_22350);
or U22505 (N_22505,N_22380,N_22400);
or U22506 (N_22506,N_22266,N_22375);
nor U22507 (N_22507,N_22480,N_22419);
nand U22508 (N_22508,N_22442,N_22361);
and U22509 (N_22509,N_22343,N_22374);
nand U22510 (N_22510,N_22311,N_22440);
and U22511 (N_22511,N_22482,N_22300);
nand U22512 (N_22512,N_22356,N_22466);
or U22513 (N_22513,N_22265,N_22276);
and U22514 (N_22514,N_22398,N_22360);
or U22515 (N_22515,N_22306,N_22488);
or U22516 (N_22516,N_22365,N_22332);
nor U22517 (N_22517,N_22349,N_22444);
nor U22518 (N_22518,N_22368,N_22302);
or U22519 (N_22519,N_22386,N_22289);
and U22520 (N_22520,N_22438,N_22463);
nor U22521 (N_22521,N_22330,N_22478);
nand U22522 (N_22522,N_22290,N_22342);
nand U22523 (N_22523,N_22448,N_22433);
nor U22524 (N_22524,N_22335,N_22313);
nor U22525 (N_22525,N_22337,N_22327);
nand U22526 (N_22526,N_22468,N_22291);
and U22527 (N_22527,N_22404,N_22315);
nand U22528 (N_22528,N_22331,N_22270);
or U22529 (N_22529,N_22317,N_22464);
nor U22530 (N_22530,N_22422,N_22436);
nand U22531 (N_22531,N_22322,N_22394);
or U22532 (N_22532,N_22373,N_22370);
nor U22533 (N_22533,N_22431,N_22257);
nor U22534 (N_22534,N_22428,N_22274);
or U22535 (N_22535,N_22498,N_22258);
or U22536 (N_22536,N_22399,N_22369);
nor U22537 (N_22537,N_22473,N_22434);
and U22538 (N_22538,N_22487,N_22465);
and U22539 (N_22539,N_22409,N_22421);
or U22540 (N_22540,N_22391,N_22486);
nand U22541 (N_22541,N_22389,N_22408);
or U22542 (N_22542,N_22351,N_22268);
or U22543 (N_22543,N_22286,N_22344);
and U22544 (N_22544,N_22275,N_22471);
nor U22545 (N_22545,N_22447,N_22340);
nand U22546 (N_22546,N_22424,N_22390);
and U22547 (N_22547,N_22251,N_22445);
and U22548 (N_22548,N_22309,N_22407);
nand U22549 (N_22549,N_22272,N_22314);
nor U22550 (N_22550,N_22381,N_22295);
nor U22551 (N_22551,N_22437,N_22446);
nor U22552 (N_22552,N_22296,N_22481);
nor U22553 (N_22553,N_22493,N_22496);
nor U22554 (N_22554,N_22283,N_22441);
nor U22555 (N_22555,N_22382,N_22469);
and U22556 (N_22556,N_22297,N_22352);
or U22557 (N_22557,N_22417,N_22321);
and U22558 (N_22558,N_22395,N_22287);
and U22559 (N_22559,N_22485,N_22363);
nand U22560 (N_22560,N_22401,N_22397);
nor U22561 (N_22561,N_22310,N_22308);
and U22562 (N_22562,N_22454,N_22304);
nor U22563 (N_22563,N_22282,N_22293);
nand U22564 (N_22564,N_22477,N_22443);
nor U22565 (N_22565,N_22489,N_22474);
nand U22566 (N_22566,N_22279,N_22455);
nor U22567 (N_22567,N_22467,N_22346);
and U22568 (N_22568,N_22354,N_22336);
and U22569 (N_22569,N_22425,N_22423);
nor U22570 (N_22570,N_22353,N_22288);
and U22571 (N_22571,N_22457,N_22415);
nand U22572 (N_22572,N_22472,N_22367);
and U22573 (N_22573,N_22345,N_22377);
nand U22574 (N_22574,N_22362,N_22470);
nand U22575 (N_22575,N_22262,N_22359);
nand U22576 (N_22576,N_22403,N_22338);
or U22577 (N_22577,N_22255,N_22497);
nor U22578 (N_22578,N_22261,N_22326);
and U22579 (N_22579,N_22319,N_22298);
nand U22580 (N_22580,N_22430,N_22324);
and U22581 (N_22581,N_22435,N_22396);
and U22582 (N_22582,N_22284,N_22411);
nand U22583 (N_22583,N_22260,N_22263);
nor U22584 (N_22584,N_22292,N_22294);
or U22585 (N_22585,N_22460,N_22267);
nor U22586 (N_22586,N_22372,N_22339);
or U22587 (N_22587,N_22256,N_22393);
nand U22588 (N_22588,N_22416,N_22459);
nand U22589 (N_22589,N_22250,N_22334);
nor U22590 (N_22590,N_22439,N_22252);
and U22591 (N_22591,N_22280,N_22476);
nand U22592 (N_22592,N_22376,N_22452);
nand U22593 (N_22593,N_22413,N_22301);
nand U22594 (N_22594,N_22278,N_22458);
nor U22595 (N_22595,N_22358,N_22410);
nand U22596 (N_22596,N_22273,N_22412);
or U22597 (N_22597,N_22347,N_22371);
or U22598 (N_22598,N_22449,N_22341);
nand U22599 (N_22599,N_22318,N_22254);
and U22600 (N_22600,N_22348,N_22325);
nor U22601 (N_22601,N_22406,N_22323);
nand U22602 (N_22602,N_22385,N_22379);
and U22603 (N_22603,N_22383,N_22420);
nor U22604 (N_22604,N_22299,N_22484);
and U22605 (N_22605,N_22264,N_22378);
nand U22606 (N_22606,N_22491,N_22414);
and U22607 (N_22607,N_22418,N_22388);
nor U22608 (N_22608,N_22328,N_22492);
nor U22609 (N_22609,N_22312,N_22320);
or U22610 (N_22610,N_22402,N_22333);
nand U22611 (N_22611,N_22456,N_22461);
or U22612 (N_22612,N_22285,N_22429);
nand U22613 (N_22613,N_22387,N_22269);
nand U22614 (N_22614,N_22479,N_22490);
and U22615 (N_22615,N_22450,N_22307);
and U22616 (N_22616,N_22364,N_22277);
or U22617 (N_22617,N_22427,N_22426);
or U22618 (N_22618,N_22281,N_22305);
or U22619 (N_22619,N_22475,N_22316);
nand U22620 (N_22620,N_22384,N_22453);
nand U22621 (N_22621,N_22495,N_22392);
or U22622 (N_22622,N_22329,N_22259);
or U22623 (N_22623,N_22451,N_22355);
nor U22624 (N_22624,N_22494,N_22271);
and U22625 (N_22625,N_22464,N_22250);
nand U22626 (N_22626,N_22464,N_22442);
and U22627 (N_22627,N_22337,N_22370);
nand U22628 (N_22628,N_22375,N_22260);
nor U22629 (N_22629,N_22430,N_22468);
and U22630 (N_22630,N_22469,N_22349);
or U22631 (N_22631,N_22275,N_22384);
and U22632 (N_22632,N_22414,N_22487);
and U22633 (N_22633,N_22362,N_22319);
or U22634 (N_22634,N_22450,N_22424);
or U22635 (N_22635,N_22495,N_22375);
nand U22636 (N_22636,N_22427,N_22408);
or U22637 (N_22637,N_22261,N_22430);
nand U22638 (N_22638,N_22484,N_22280);
and U22639 (N_22639,N_22266,N_22429);
nor U22640 (N_22640,N_22264,N_22470);
and U22641 (N_22641,N_22354,N_22480);
and U22642 (N_22642,N_22340,N_22391);
or U22643 (N_22643,N_22371,N_22426);
and U22644 (N_22644,N_22408,N_22267);
nand U22645 (N_22645,N_22425,N_22321);
and U22646 (N_22646,N_22413,N_22419);
or U22647 (N_22647,N_22439,N_22296);
nor U22648 (N_22648,N_22273,N_22345);
and U22649 (N_22649,N_22432,N_22372);
or U22650 (N_22650,N_22426,N_22380);
nor U22651 (N_22651,N_22444,N_22498);
nor U22652 (N_22652,N_22464,N_22462);
and U22653 (N_22653,N_22454,N_22298);
nor U22654 (N_22654,N_22292,N_22466);
nand U22655 (N_22655,N_22288,N_22380);
nand U22656 (N_22656,N_22273,N_22477);
nor U22657 (N_22657,N_22497,N_22257);
nor U22658 (N_22658,N_22343,N_22320);
nand U22659 (N_22659,N_22408,N_22402);
nand U22660 (N_22660,N_22354,N_22482);
nand U22661 (N_22661,N_22250,N_22423);
nor U22662 (N_22662,N_22412,N_22369);
and U22663 (N_22663,N_22386,N_22366);
nor U22664 (N_22664,N_22481,N_22337);
nor U22665 (N_22665,N_22440,N_22309);
nor U22666 (N_22666,N_22324,N_22432);
or U22667 (N_22667,N_22453,N_22259);
nand U22668 (N_22668,N_22391,N_22435);
nor U22669 (N_22669,N_22469,N_22449);
nand U22670 (N_22670,N_22375,N_22374);
or U22671 (N_22671,N_22306,N_22455);
nand U22672 (N_22672,N_22429,N_22442);
nor U22673 (N_22673,N_22286,N_22340);
nand U22674 (N_22674,N_22491,N_22388);
nand U22675 (N_22675,N_22283,N_22483);
nand U22676 (N_22676,N_22437,N_22252);
nor U22677 (N_22677,N_22493,N_22373);
or U22678 (N_22678,N_22420,N_22446);
nand U22679 (N_22679,N_22297,N_22345);
or U22680 (N_22680,N_22426,N_22484);
and U22681 (N_22681,N_22382,N_22383);
nand U22682 (N_22682,N_22354,N_22359);
or U22683 (N_22683,N_22405,N_22394);
and U22684 (N_22684,N_22418,N_22372);
nand U22685 (N_22685,N_22352,N_22361);
or U22686 (N_22686,N_22474,N_22352);
and U22687 (N_22687,N_22449,N_22299);
or U22688 (N_22688,N_22320,N_22382);
and U22689 (N_22689,N_22358,N_22257);
and U22690 (N_22690,N_22453,N_22422);
and U22691 (N_22691,N_22436,N_22388);
or U22692 (N_22692,N_22280,N_22434);
nor U22693 (N_22693,N_22490,N_22435);
or U22694 (N_22694,N_22283,N_22278);
or U22695 (N_22695,N_22289,N_22340);
or U22696 (N_22696,N_22482,N_22438);
nand U22697 (N_22697,N_22472,N_22404);
nand U22698 (N_22698,N_22472,N_22421);
or U22699 (N_22699,N_22353,N_22476);
and U22700 (N_22700,N_22286,N_22463);
nor U22701 (N_22701,N_22399,N_22386);
and U22702 (N_22702,N_22363,N_22452);
or U22703 (N_22703,N_22407,N_22375);
or U22704 (N_22704,N_22269,N_22431);
or U22705 (N_22705,N_22294,N_22489);
and U22706 (N_22706,N_22313,N_22258);
or U22707 (N_22707,N_22286,N_22456);
and U22708 (N_22708,N_22451,N_22320);
or U22709 (N_22709,N_22310,N_22399);
nor U22710 (N_22710,N_22385,N_22389);
nand U22711 (N_22711,N_22462,N_22434);
xor U22712 (N_22712,N_22477,N_22478);
nand U22713 (N_22713,N_22486,N_22286);
or U22714 (N_22714,N_22457,N_22350);
nor U22715 (N_22715,N_22330,N_22460);
or U22716 (N_22716,N_22374,N_22290);
nor U22717 (N_22717,N_22435,N_22346);
and U22718 (N_22718,N_22380,N_22378);
or U22719 (N_22719,N_22365,N_22385);
nand U22720 (N_22720,N_22460,N_22282);
and U22721 (N_22721,N_22442,N_22333);
or U22722 (N_22722,N_22339,N_22251);
or U22723 (N_22723,N_22265,N_22316);
and U22724 (N_22724,N_22336,N_22469);
nor U22725 (N_22725,N_22424,N_22498);
nand U22726 (N_22726,N_22414,N_22347);
nand U22727 (N_22727,N_22347,N_22344);
nor U22728 (N_22728,N_22276,N_22394);
nand U22729 (N_22729,N_22342,N_22397);
or U22730 (N_22730,N_22480,N_22320);
and U22731 (N_22731,N_22454,N_22315);
nand U22732 (N_22732,N_22402,N_22492);
and U22733 (N_22733,N_22267,N_22252);
nand U22734 (N_22734,N_22483,N_22312);
nor U22735 (N_22735,N_22389,N_22287);
or U22736 (N_22736,N_22436,N_22345);
or U22737 (N_22737,N_22480,N_22326);
nand U22738 (N_22738,N_22338,N_22251);
or U22739 (N_22739,N_22267,N_22393);
nand U22740 (N_22740,N_22449,N_22442);
nand U22741 (N_22741,N_22293,N_22331);
or U22742 (N_22742,N_22255,N_22250);
nor U22743 (N_22743,N_22331,N_22327);
and U22744 (N_22744,N_22448,N_22314);
or U22745 (N_22745,N_22444,N_22280);
or U22746 (N_22746,N_22480,N_22437);
nand U22747 (N_22747,N_22331,N_22360);
nand U22748 (N_22748,N_22412,N_22443);
nand U22749 (N_22749,N_22400,N_22309);
or U22750 (N_22750,N_22584,N_22574);
and U22751 (N_22751,N_22604,N_22729);
nand U22752 (N_22752,N_22718,N_22674);
or U22753 (N_22753,N_22601,N_22596);
or U22754 (N_22754,N_22611,N_22665);
nand U22755 (N_22755,N_22614,N_22739);
nand U22756 (N_22756,N_22548,N_22624);
nor U22757 (N_22757,N_22555,N_22513);
nand U22758 (N_22758,N_22605,N_22618);
nand U22759 (N_22759,N_22667,N_22664);
nor U22760 (N_22760,N_22632,N_22704);
or U22761 (N_22761,N_22675,N_22515);
nand U22762 (N_22762,N_22510,N_22528);
or U22763 (N_22763,N_22737,N_22659);
nor U22764 (N_22764,N_22657,N_22625);
nand U22765 (N_22765,N_22736,N_22606);
or U22766 (N_22766,N_22685,N_22690);
or U22767 (N_22767,N_22655,N_22587);
nor U22768 (N_22768,N_22658,N_22546);
or U22769 (N_22769,N_22620,N_22529);
or U22770 (N_22770,N_22539,N_22749);
nor U22771 (N_22771,N_22720,N_22716);
or U22772 (N_22772,N_22557,N_22568);
nor U22773 (N_22773,N_22647,N_22609);
nor U22774 (N_22774,N_22600,N_22560);
nor U22775 (N_22775,N_22563,N_22644);
or U22776 (N_22776,N_22676,N_22705);
and U22777 (N_22777,N_22504,N_22530);
nor U22778 (N_22778,N_22503,N_22554);
nor U22779 (N_22779,N_22662,N_22575);
or U22780 (N_22780,N_22559,N_22651);
and U22781 (N_22781,N_22520,N_22589);
nor U22782 (N_22782,N_22607,N_22516);
nand U22783 (N_22783,N_22580,N_22523);
nand U22784 (N_22784,N_22715,N_22613);
and U22785 (N_22785,N_22687,N_22512);
nand U22786 (N_22786,N_22509,N_22506);
nor U22787 (N_22787,N_22550,N_22610);
nor U22788 (N_22788,N_22725,N_22670);
or U22789 (N_22789,N_22514,N_22558);
nor U22790 (N_22790,N_22538,N_22719);
or U22791 (N_22791,N_22707,N_22653);
or U22792 (N_22792,N_22572,N_22570);
nor U22793 (N_22793,N_22518,N_22608);
nor U22794 (N_22794,N_22733,N_22746);
nor U22795 (N_22795,N_22660,N_22534);
nand U22796 (N_22796,N_22717,N_22508);
nor U22797 (N_22797,N_22745,N_22527);
and U22798 (N_22798,N_22661,N_22710);
nor U22799 (N_22799,N_22623,N_22627);
or U22800 (N_22800,N_22723,N_22597);
and U22801 (N_22801,N_22693,N_22650);
or U22802 (N_22802,N_22590,N_22556);
or U22803 (N_22803,N_22615,N_22566);
or U22804 (N_22804,N_22540,N_22639);
nand U22805 (N_22805,N_22629,N_22592);
or U22806 (N_22806,N_22748,N_22544);
nor U22807 (N_22807,N_22581,N_22689);
and U22808 (N_22808,N_22669,N_22680);
nor U22809 (N_22809,N_22635,N_22543);
and U22810 (N_22810,N_22549,N_22722);
nor U22811 (N_22811,N_22649,N_22526);
and U22812 (N_22812,N_22691,N_22619);
nand U22813 (N_22813,N_22697,N_22634);
nor U22814 (N_22814,N_22631,N_22582);
and U22815 (N_22815,N_22700,N_22652);
and U22816 (N_22816,N_22542,N_22740);
and U22817 (N_22817,N_22640,N_22501);
nand U22818 (N_22818,N_22714,N_22517);
nand U22819 (N_22819,N_22552,N_22636);
and U22820 (N_22820,N_22709,N_22594);
nand U22821 (N_22821,N_22562,N_22599);
and U22822 (N_22822,N_22583,N_22547);
nand U22823 (N_22823,N_22648,N_22525);
or U22824 (N_22824,N_22521,N_22698);
and U22825 (N_22825,N_22500,N_22735);
nor U22826 (N_22826,N_22626,N_22708);
and U22827 (N_22827,N_22679,N_22683);
nand U22828 (N_22828,N_22533,N_22701);
nor U22829 (N_22829,N_22622,N_22673);
or U22830 (N_22830,N_22569,N_22642);
and U22831 (N_22831,N_22688,N_22564);
xor U22832 (N_22832,N_22612,N_22541);
and U22833 (N_22833,N_22595,N_22668);
or U22834 (N_22834,N_22643,N_22703);
nand U22835 (N_22835,N_22522,N_22593);
nor U22836 (N_22836,N_22507,N_22532);
and U22837 (N_22837,N_22565,N_22617);
and U22838 (N_22838,N_22677,N_22699);
nand U22839 (N_22839,N_22633,N_22535);
nand U22840 (N_22840,N_22684,N_22567);
nor U22841 (N_22841,N_22505,N_22603);
and U22842 (N_22842,N_22553,N_22654);
nand U22843 (N_22843,N_22598,N_22731);
xor U22844 (N_22844,N_22578,N_22637);
and U22845 (N_22845,N_22645,N_22721);
nand U22846 (N_22846,N_22616,N_22702);
nor U22847 (N_22847,N_22656,N_22638);
nand U22848 (N_22848,N_22681,N_22672);
and U22849 (N_22849,N_22628,N_22686);
nand U22850 (N_22850,N_22711,N_22511);
nand U22851 (N_22851,N_22730,N_22577);
and U22852 (N_22852,N_22696,N_22573);
xor U22853 (N_22853,N_22663,N_22727);
nor U22854 (N_22854,N_22712,N_22666);
and U22855 (N_22855,N_22646,N_22744);
and U22856 (N_22856,N_22561,N_22706);
and U22857 (N_22857,N_22728,N_22678);
or U22858 (N_22858,N_22531,N_22741);
nand U22859 (N_22859,N_22537,N_22588);
nor U22860 (N_22860,N_22630,N_22591);
or U22861 (N_22861,N_22545,N_22519);
nand U22862 (N_22862,N_22524,N_22621);
nand U22863 (N_22863,N_22585,N_22692);
nand U22864 (N_22864,N_22641,N_22586);
nor U22865 (N_22865,N_22502,N_22576);
nor U22866 (N_22866,N_22536,N_22747);
nor U22867 (N_22867,N_22551,N_22671);
nor U22868 (N_22868,N_22682,N_22742);
nand U22869 (N_22869,N_22579,N_22732);
or U22870 (N_22870,N_22734,N_22571);
and U22871 (N_22871,N_22695,N_22602);
or U22872 (N_22872,N_22713,N_22726);
nand U22873 (N_22873,N_22738,N_22743);
nand U22874 (N_22874,N_22694,N_22724);
nand U22875 (N_22875,N_22585,N_22531);
or U22876 (N_22876,N_22742,N_22688);
nor U22877 (N_22877,N_22678,N_22687);
nor U22878 (N_22878,N_22682,N_22561);
or U22879 (N_22879,N_22697,N_22642);
nand U22880 (N_22880,N_22725,N_22550);
or U22881 (N_22881,N_22700,N_22732);
nand U22882 (N_22882,N_22608,N_22649);
and U22883 (N_22883,N_22664,N_22572);
nor U22884 (N_22884,N_22686,N_22670);
nor U22885 (N_22885,N_22699,N_22653);
and U22886 (N_22886,N_22737,N_22517);
nand U22887 (N_22887,N_22721,N_22725);
nand U22888 (N_22888,N_22534,N_22716);
or U22889 (N_22889,N_22653,N_22708);
nor U22890 (N_22890,N_22629,N_22727);
nand U22891 (N_22891,N_22651,N_22620);
and U22892 (N_22892,N_22563,N_22585);
or U22893 (N_22893,N_22738,N_22650);
or U22894 (N_22894,N_22664,N_22596);
xor U22895 (N_22895,N_22595,N_22698);
nand U22896 (N_22896,N_22650,N_22551);
nand U22897 (N_22897,N_22607,N_22604);
nor U22898 (N_22898,N_22628,N_22597);
or U22899 (N_22899,N_22608,N_22718);
or U22900 (N_22900,N_22672,N_22687);
or U22901 (N_22901,N_22654,N_22675);
nor U22902 (N_22902,N_22693,N_22677);
and U22903 (N_22903,N_22644,N_22688);
or U22904 (N_22904,N_22611,N_22624);
or U22905 (N_22905,N_22697,N_22735);
and U22906 (N_22906,N_22694,N_22608);
or U22907 (N_22907,N_22587,N_22588);
and U22908 (N_22908,N_22721,N_22677);
nand U22909 (N_22909,N_22514,N_22741);
and U22910 (N_22910,N_22521,N_22744);
or U22911 (N_22911,N_22604,N_22615);
and U22912 (N_22912,N_22561,N_22667);
nor U22913 (N_22913,N_22691,N_22554);
nand U22914 (N_22914,N_22618,N_22650);
nand U22915 (N_22915,N_22697,N_22689);
or U22916 (N_22916,N_22540,N_22580);
nor U22917 (N_22917,N_22549,N_22610);
nor U22918 (N_22918,N_22726,N_22746);
and U22919 (N_22919,N_22705,N_22516);
and U22920 (N_22920,N_22689,N_22588);
nor U22921 (N_22921,N_22563,N_22652);
and U22922 (N_22922,N_22629,N_22648);
and U22923 (N_22923,N_22682,N_22598);
and U22924 (N_22924,N_22552,N_22695);
nand U22925 (N_22925,N_22636,N_22602);
and U22926 (N_22926,N_22529,N_22611);
nor U22927 (N_22927,N_22521,N_22719);
or U22928 (N_22928,N_22669,N_22591);
nor U22929 (N_22929,N_22703,N_22561);
and U22930 (N_22930,N_22731,N_22623);
and U22931 (N_22931,N_22698,N_22527);
nor U22932 (N_22932,N_22643,N_22531);
or U22933 (N_22933,N_22720,N_22551);
nor U22934 (N_22934,N_22747,N_22681);
nand U22935 (N_22935,N_22687,N_22574);
and U22936 (N_22936,N_22611,N_22677);
or U22937 (N_22937,N_22734,N_22744);
nor U22938 (N_22938,N_22562,N_22572);
or U22939 (N_22939,N_22748,N_22525);
or U22940 (N_22940,N_22610,N_22656);
and U22941 (N_22941,N_22721,N_22607);
nand U22942 (N_22942,N_22717,N_22528);
or U22943 (N_22943,N_22686,N_22642);
or U22944 (N_22944,N_22527,N_22657);
nor U22945 (N_22945,N_22624,N_22534);
and U22946 (N_22946,N_22601,N_22666);
and U22947 (N_22947,N_22706,N_22587);
or U22948 (N_22948,N_22644,N_22542);
and U22949 (N_22949,N_22710,N_22600);
nand U22950 (N_22950,N_22675,N_22596);
nor U22951 (N_22951,N_22574,N_22507);
or U22952 (N_22952,N_22597,N_22502);
or U22953 (N_22953,N_22512,N_22590);
and U22954 (N_22954,N_22533,N_22669);
and U22955 (N_22955,N_22641,N_22746);
and U22956 (N_22956,N_22550,N_22650);
nand U22957 (N_22957,N_22696,N_22742);
nor U22958 (N_22958,N_22591,N_22523);
and U22959 (N_22959,N_22687,N_22747);
nand U22960 (N_22960,N_22615,N_22514);
nor U22961 (N_22961,N_22601,N_22679);
or U22962 (N_22962,N_22720,N_22574);
or U22963 (N_22963,N_22581,N_22578);
nand U22964 (N_22964,N_22589,N_22618);
or U22965 (N_22965,N_22613,N_22568);
nand U22966 (N_22966,N_22744,N_22635);
and U22967 (N_22967,N_22701,N_22522);
or U22968 (N_22968,N_22692,N_22648);
nor U22969 (N_22969,N_22559,N_22703);
and U22970 (N_22970,N_22568,N_22541);
or U22971 (N_22971,N_22616,N_22733);
or U22972 (N_22972,N_22593,N_22585);
nor U22973 (N_22973,N_22709,N_22602);
or U22974 (N_22974,N_22715,N_22668);
or U22975 (N_22975,N_22541,N_22531);
or U22976 (N_22976,N_22618,N_22508);
and U22977 (N_22977,N_22675,N_22512);
nor U22978 (N_22978,N_22545,N_22735);
and U22979 (N_22979,N_22609,N_22539);
xnor U22980 (N_22980,N_22664,N_22539);
nand U22981 (N_22981,N_22674,N_22549);
nand U22982 (N_22982,N_22626,N_22649);
and U22983 (N_22983,N_22525,N_22615);
and U22984 (N_22984,N_22721,N_22589);
or U22985 (N_22985,N_22672,N_22533);
and U22986 (N_22986,N_22642,N_22606);
nand U22987 (N_22987,N_22518,N_22631);
nor U22988 (N_22988,N_22664,N_22634);
and U22989 (N_22989,N_22609,N_22564);
nor U22990 (N_22990,N_22662,N_22680);
and U22991 (N_22991,N_22504,N_22614);
or U22992 (N_22992,N_22749,N_22525);
and U22993 (N_22993,N_22585,N_22654);
and U22994 (N_22994,N_22733,N_22716);
nor U22995 (N_22995,N_22704,N_22691);
and U22996 (N_22996,N_22684,N_22710);
and U22997 (N_22997,N_22682,N_22563);
and U22998 (N_22998,N_22517,N_22732);
and U22999 (N_22999,N_22623,N_22682);
nand U23000 (N_23000,N_22796,N_22919);
or U23001 (N_23001,N_22899,N_22798);
nor U23002 (N_23002,N_22876,N_22957);
or U23003 (N_23003,N_22766,N_22981);
and U23004 (N_23004,N_22922,N_22974);
nor U23005 (N_23005,N_22832,N_22801);
nor U23006 (N_23006,N_22911,N_22964);
or U23007 (N_23007,N_22794,N_22849);
nor U23008 (N_23008,N_22753,N_22847);
nand U23009 (N_23009,N_22912,N_22888);
nand U23010 (N_23010,N_22809,N_22978);
and U23011 (N_23011,N_22928,N_22987);
and U23012 (N_23012,N_22971,N_22800);
nor U23013 (N_23013,N_22767,N_22810);
nand U23014 (N_23014,N_22945,N_22902);
nor U23015 (N_23015,N_22841,N_22967);
or U23016 (N_23016,N_22958,N_22782);
nand U23017 (N_23017,N_22940,N_22965);
and U23018 (N_23018,N_22952,N_22771);
and U23019 (N_23019,N_22861,N_22938);
and U23020 (N_23020,N_22909,N_22779);
and U23021 (N_23021,N_22828,N_22860);
or U23022 (N_23022,N_22975,N_22830);
or U23023 (N_23023,N_22880,N_22781);
nor U23024 (N_23024,N_22803,N_22890);
nand U23025 (N_23025,N_22769,N_22775);
or U23026 (N_23026,N_22825,N_22807);
nand U23027 (N_23027,N_22959,N_22823);
nand U23028 (N_23028,N_22813,N_22770);
or U23029 (N_23029,N_22793,N_22929);
and U23030 (N_23030,N_22961,N_22976);
or U23031 (N_23031,N_22821,N_22894);
and U23032 (N_23032,N_22937,N_22996);
nor U23033 (N_23033,N_22903,N_22916);
and U23034 (N_23034,N_22924,N_22984);
nor U23035 (N_23035,N_22994,N_22776);
nor U23036 (N_23036,N_22802,N_22754);
or U23037 (N_23037,N_22925,N_22921);
and U23038 (N_23038,N_22804,N_22914);
and U23039 (N_23039,N_22787,N_22907);
nor U23040 (N_23040,N_22791,N_22881);
and U23041 (N_23041,N_22837,N_22756);
or U23042 (N_23042,N_22820,N_22953);
and U23043 (N_23043,N_22969,N_22943);
and U23044 (N_23044,N_22785,N_22883);
nor U23045 (N_23045,N_22864,N_22910);
or U23046 (N_23046,N_22752,N_22946);
and U23047 (N_23047,N_22757,N_22777);
nand U23048 (N_23048,N_22973,N_22962);
or U23049 (N_23049,N_22778,N_22855);
and U23050 (N_23050,N_22970,N_22838);
and U23051 (N_23051,N_22873,N_22942);
nor U23052 (N_23052,N_22759,N_22853);
and U23053 (N_23053,N_22901,N_22980);
or U23054 (N_23054,N_22790,N_22886);
and U23055 (N_23055,N_22963,N_22816);
and U23056 (N_23056,N_22815,N_22833);
nor U23057 (N_23057,N_22991,N_22908);
nor U23058 (N_23058,N_22751,N_22898);
nand U23059 (N_23059,N_22818,N_22986);
or U23060 (N_23060,N_22765,N_22863);
nor U23061 (N_23061,N_22896,N_22805);
nor U23062 (N_23062,N_22842,N_22939);
nor U23063 (N_23063,N_22934,N_22764);
nand U23064 (N_23064,N_22789,N_22835);
and U23065 (N_23065,N_22871,N_22915);
nand U23066 (N_23066,N_22755,N_22993);
nand U23067 (N_23067,N_22941,N_22786);
nor U23068 (N_23068,N_22836,N_22761);
nor U23069 (N_23069,N_22808,N_22913);
nand U23070 (N_23070,N_22892,N_22875);
nand U23071 (N_23071,N_22867,N_22762);
and U23072 (N_23072,N_22799,N_22960);
nand U23073 (N_23073,N_22877,N_22859);
nor U23074 (N_23074,N_22992,N_22997);
nand U23075 (N_23075,N_22850,N_22819);
nand U23076 (N_23076,N_22868,N_22750);
or U23077 (N_23077,N_22848,N_22917);
or U23078 (N_23078,N_22931,N_22900);
or U23079 (N_23079,N_22872,N_22874);
or U23080 (N_23080,N_22988,N_22840);
nand U23081 (N_23081,N_22936,N_22889);
nor U23082 (N_23082,N_22930,N_22893);
nor U23083 (N_23083,N_22846,N_22814);
nor U23084 (N_23084,N_22956,N_22783);
nand U23085 (N_23085,N_22862,N_22950);
nand U23086 (N_23086,N_22839,N_22772);
nor U23087 (N_23087,N_22904,N_22845);
or U23088 (N_23088,N_22985,N_22990);
or U23089 (N_23089,N_22951,N_22812);
and U23090 (N_23090,N_22944,N_22829);
or U23091 (N_23091,N_22884,N_22932);
nor U23092 (N_23092,N_22858,N_22966);
nor U23093 (N_23093,N_22995,N_22948);
and U23094 (N_23094,N_22857,N_22852);
nor U23095 (N_23095,N_22768,N_22891);
nor U23096 (N_23096,N_22773,N_22882);
nor U23097 (N_23097,N_22935,N_22999);
and U23098 (N_23098,N_22954,N_22879);
nand U23099 (N_23099,N_22983,N_22895);
or U23100 (N_23100,N_22824,N_22949);
nand U23101 (N_23101,N_22806,N_22885);
and U23102 (N_23102,N_22968,N_22826);
and U23103 (N_23103,N_22977,N_22982);
or U23104 (N_23104,N_22933,N_22920);
nand U23105 (N_23105,N_22788,N_22865);
or U23106 (N_23106,N_22760,N_22831);
nor U23107 (N_23107,N_22887,N_22763);
or U23108 (N_23108,N_22972,N_22827);
nand U23109 (N_23109,N_22784,N_22795);
or U23110 (N_23110,N_22905,N_22955);
and U23111 (N_23111,N_22797,N_22947);
nand U23112 (N_23112,N_22780,N_22926);
nor U23113 (N_23113,N_22927,N_22989);
or U23114 (N_23114,N_22869,N_22878);
or U23115 (N_23115,N_22897,N_22998);
and U23116 (N_23116,N_22822,N_22843);
or U23117 (N_23117,N_22866,N_22979);
xnor U23118 (N_23118,N_22792,N_22774);
nand U23119 (N_23119,N_22851,N_22811);
or U23120 (N_23120,N_22870,N_22906);
and U23121 (N_23121,N_22923,N_22844);
nand U23122 (N_23122,N_22856,N_22834);
and U23123 (N_23123,N_22817,N_22758);
or U23124 (N_23124,N_22918,N_22854);
and U23125 (N_23125,N_22955,N_22867);
and U23126 (N_23126,N_22995,N_22902);
or U23127 (N_23127,N_22800,N_22754);
and U23128 (N_23128,N_22902,N_22752);
and U23129 (N_23129,N_22760,N_22835);
nand U23130 (N_23130,N_22984,N_22967);
and U23131 (N_23131,N_22795,N_22781);
and U23132 (N_23132,N_22988,N_22784);
nor U23133 (N_23133,N_22898,N_22805);
nand U23134 (N_23134,N_22843,N_22948);
or U23135 (N_23135,N_22906,N_22856);
and U23136 (N_23136,N_22823,N_22885);
or U23137 (N_23137,N_22861,N_22892);
or U23138 (N_23138,N_22995,N_22851);
or U23139 (N_23139,N_22920,N_22946);
and U23140 (N_23140,N_22866,N_22943);
nand U23141 (N_23141,N_22983,N_22785);
or U23142 (N_23142,N_22773,N_22932);
or U23143 (N_23143,N_22943,N_22974);
nand U23144 (N_23144,N_22760,N_22813);
nand U23145 (N_23145,N_22997,N_22804);
nor U23146 (N_23146,N_22833,N_22907);
and U23147 (N_23147,N_22775,N_22865);
or U23148 (N_23148,N_22822,N_22828);
or U23149 (N_23149,N_22985,N_22886);
or U23150 (N_23150,N_22851,N_22915);
or U23151 (N_23151,N_22826,N_22963);
nand U23152 (N_23152,N_22810,N_22919);
or U23153 (N_23153,N_22835,N_22957);
and U23154 (N_23154,N_22769,N_22897);
nand U23155 (N_23155,N_22847,N_22808);
nand U23156 (N_23156,N_22894,N_22772);
and U23157 (N_23157,N_22989,N_22909);
nor U23158 (N_23158,N_22792,N_22886);
and U23159 (N_23159,N_22987,N_22802);
nand U23160 (N_23160,N_22765,N_22983);
nand U23161 (N_23161,N_22801,N_22939);
or U23162 (N_23162,N_22755,N_22852);
nand U23163 (N_23163,N_22825,N_22838);
nand U23164 (N_23164,N_22892,N_22930);
or U23165 (N_23165,N_22992,N_22773);
nor U23166 (N_23166,N_22915,N_22772);
and U23167 (N_23167,N_22967,N_22904);
nand U23168 (N_23168,N_22948,N_22860);
nand U23169 (N_23169,N_22939,N_22935);
nand U23170 (N_23170,N_22974,N_22986);
nand U23171 (N_23171,N_22881,N_22864);
nand U23172 (N_23172,N_22791,N_22868);
xor U23173 (N_23173,N_22913,N_22893);
nor U23174 (N_23174,N_22798,N_22955);
and U23175 (N_23175,N_22773,N_22797);
nor U23176 (N_23176,N_22823,N_22917);
or U23177 (N_23177,N_22990,N_22896);
or U23178 (N_23178,N_22906,N_22787);
and U23179 (N_23179,N_22987,N_22848);
nor U23180 (N_23180,N_22921,N_22895);
nor U23181 (N_23181,N_22901,N_22770);
and U23182 (N_23182,N_22757,N_22862);
and U23183 (N_23183,N_22864,N_22926);
nand U23184 (N_23184,N_22852,N_22787);
nor U23185 (N_23185,N_22831,N_22836);
and U23186 (N_23186,N_22767,N_22920);
nand U23187 (N_23187,N_22809,N_22893);
nand U23188 (N_23188,N_22901,N_22803);
nor U23189 (N_23189,N_22799,N_22948);
and U23190 (N_23190,N_22875,N_22960);
and U23191 (N_23191,N_22933,N_22811);
or U23192 (N_23192,N_22866,N_22829);
nand U23193 (N_23193,N_22901,N_22927);
nor U23194 (N_23194,N_22775,N_22762);
and U23195 (N_23195,N_22838,N_22815);
nor U23196 (N_23196,N_22785,N_22967);
nor U23197 (N_23197,N_22975,N_22958);
nor U23198 (N_23198,N_22911,N_22918);
or U23199 (N_23199,N_22949,N_22864);
and U23200 (N_23200,N_22916,N_22987);
nor U23201 (N_23201,N_22768,N_22919);
or U23202 (N_23202,N_22957,N_22988);
and U23203 (N_23203,N_22868,N_22919);
nand U23204 (N_23204,N_22874,N_22949);
nand U23205 (N_23205,N_22911,N_22794);
and U23206 (N_23206,N_22776,N_22842);
nor U23207 (N_23207,N_22868,N_22963);
nor U23208 (N_23208,N_22858,N_22964);
nor U23209 (N_23209,N_22902,N_22926);
nor U23210 (N_23210,N_22750,N_22814);
nand U23211 (N_23211,N_22896,N_22983);
nand U23212 (N_23212,N_22812,N_22865);
nand U23213 (N_23213,N_22922,N_22899);
and U23214 (N_23214,N_22922,N_22935);
and U23215 (N_23215,N_22768,N_22774);
nand U23216 (N_23216,N_22955,N_22978);
nor U23217 (N_23217,N_22890,N_22857);
or U23218 (N_23218,N_22952,N_22989);
nand U23219 (N_23219,N_22959,N_22795);
and U23220 (N_23220,N_22827,N_22930);
and U23221 (N_23221,N_22809,N_22939);
or U23222 (N_23222,N_22801,N_22761);
xor U23223 (N_23223,N_22756,N_22790);
nand U23224 (N_23224,N_22910,N_22922);
or U23225 (N_23225,N_22847,N_22966);
nor U23226 (N_23226,N_22987,N_22965);
nand U23227 (N_23227,N_22756,N_22872);
nand U23228 (N_23228,N_22967,N_22868);
nor U23229 (N_23229,N_22788,N_22880);
nor U23230 (N_23230,N_22842,N_22855);
nand U23231 (N_23231,N_22750,N_22834);
nor U23232 (N_23232,N_22862,N_22934);
nor U23233 (N_23233,N_22802,N_22969);
and U23234 (N_23234,N_22772,N_22795);
nor U23235 (N_23235,N_22909,N_22997);
nand U23236 (N_23236,N_22779,N_22953);
or U23237 (N_23237,N_22975,N_22781);
nand U23238 (N_23238,N_22807,N_22875);
or U23239 (N_23239,N_22913,N_22977);
and U23240 (N_23240,N_22996,N_22902);
nor U23241 (N_23241,N_22910,N_22952);
and U23242 (N_23242,N_22899,N_22797);
nor U23243 (N_23243,N_22951,N_22752);
and U23244 (N_23244,N_22894,N_22789);
nand U23245 (N_23245,N_22999,N_22964);
nor U23246 (N_23246,N_22861,N_22932);
and U23247 (N_23247,N_22764,N_22970);
or U23248 (N_23248,N_22767,N_22971);
nor U23249 (N_23249,N_22794,N_22786);
nand U23250 (N_23250,N_23186,N_23113);
and U23251 (N_23251,N_23036,N_23061);
or U23252 (N_23252,N_23229,N_23143);
nand U23253 (N_23253,N_23006,N_23232);
and U23254 (N_23254,N_23074,N_23086);
or U23255 (N_23255,N_23050,N_23035);
nand U23256 (N_23256,N_23028,N_23091);
and U23257 (N_23257,N_23058,N_23238);
nor U23258 (N_23258,N_23168,N_23083);
nor U23259 (N_23259,N_23048,N_23125);
or U23260 (N_23260,N_23241,N_23248);
nand U23261 (N_23261,N_23191,N_23000);
and U23262 (N_23262,N_23246,N_23226);
nor U23263 (N_23263,N_23115,N_23208);
nor U23264 (N_23264,N_23129,N_23233);
nor U23265 (N_23265,N_23249,N_23069);
and U23266 (N_23266,N_23009,N_23105);
nor U23267 (N_23267,N_23221,N_23173);
and U23268 (N_23268,N_23158,N_23088);
nand U23269 (N_23269,N_23064,N_23022);
nand U23270 (N_23270,N_23066,N_23167);
and U23271 (N_23271,N_23040,N_23203);
nand U23272 (N_23272,N_23179,N_23101);
and U23273 (N_23273,N_23080,N_23166);
nor U23274 (N_23274,N_23193,N_23150);
nor U23275 (N_23275,N_23020,N_23135);
and U23276 (N_23276,N_23044,N_23140);
nor U23277 (N_23277,N_23122,N_23062);
or U23278 (N_23278,N_23037,N_23205);
nor U23279 (N_23279,N_23038,N_23100);
or U23280 (N_23280,N_23130,N_23170);
and U23281 (N_23281,N_23021,N_23239);
or U23282 (N_23282,N_23180,N_23075);
nand U23283 (N_23283,N_23121,N_23185);
or U23284 (N_23284,N_23025,N_23056);
and U23285 (N_23285,N_23133,N_23141);
or U23286 (N_23286,N_23215,N_23218);
or U23287 (N_23287,N_23123,N_23007);
xnor U23288 (N_23288,N_23161,N_23010);
or U23289 (N_23289,N_23003,N_23071);
or U23290 (N_23290,N_23078,N_23070);
nor U23291 (N_23291,N_23176,N_23102);
nor U23292 (N_23292,N_23231,N_23013);
nand U23293 (N_23293,N_23174,N_23089);
nor U23294 (N_23294,N_23195,N_23212);
nor U23295 (N_23295,N_23116,N_23054);
nand U23296 (N_23296,N_23156,N_23237);
nand U23297 (N_23297,N_23151,N_23137);
or U23298 (N_23298,N_23154,N_23242);
nor U23299 (N_23299,N_23094,N_23159);
nor U23300 (N_23300,N_23128,N_23029);
or U23301 (N_23301,N_23181,N_23096);
or U23302 (N_23302,N_23107,N_23019);
and U23303 (N_23303,N_23085,N_23207);
and U23304 (N_23304,N_23202,N_23063);
and U23305 (N_23305,N_23136,N_23126);
and U23306 (N_23306,N_23030,N_23024);
or U23307 (N_23307,N_23228,N_23244);
and U23308 (N_23308,N_23211,N_23124);
and U23309 (N_23309,N_23104,N_23082);
nor U23310 (N_23310,N_23027,N_23077);
nor U23311 (N_23311,N_23081,N_23095);
and U23312 (N_23312,N_23189,N_23068);
nor U23313 (N_23313,N_23204,N_23031);
nor U23314 (N_23314,N_23149,N_23008);
nor U23315 (N_23315,N_23165,N_23178);
nand U23316 (N_23316,N_23132,N_23002);
nand U23317 (N_23317,N_23192,N_23162);
or U23318 (N_23318,N_23134,N_23004);
or U23319 (N_23319,N_23046,N_23067);
nand U23320 (N_23320,N_23073,N_23087);
or U23321 (N_23321,N_23214,N_23099);
and U23322 (N_23322,N_23005,N_23160);
or U23323 (N_23323,N_23043,N_23112);
or U23324 (N_23324,N_23245,N_23222);
nand U23325 (N_23325,N_23045,N_23057);
or U23326 (N_23326,N_23240,N_23023);
xor U23327 (N_23327,N_23227,N_23164);
nor U23328 (N_23328,N_23190,N_23175);
and U23329 (N_23329,N_23197,N_23060);
nand U23330 (N_23330,N_23147,N_23033);
and U23331 (N_23331,N_23182,N_23117);
and U23332 (N_23332,N_23219,N_23011);
xor U23333 (N_23333,N_23097,N_23153);
nand U23334 (N_23334,N_23243,N_23213);
or U23335 (N_23335,N_23118,N_23001);
nand U23336 (N_23336,N_23157,N_23217);
or U23337 (N_23337,N_23016,N_23041);
or U23338 (N_23338,N_23236,N_23093);
nand U23339 (N_23339,N_23177,N_23216);
or U23340 (N_23340,N_23059,N_23032);
and U23341 (N_23341,N_23146,N_23187);
or U23342 (N_23342,N_23201,N_23014);
and U23343 (N_23343,N_23065,N_23017);
or U23344 (N_23344,N_23184,N_23224);
nor U23345 (N_23345,N_23034,N_23206);
nor U23346 (N_23346,N_23053,N_23051);
nor U23347 (N_23347,N_23090,N_23103);
nor U23348 (N_23348,N_23163,N_23171);
and U23349 (N_23349,N_23072,N_23199);
nand U23350 (N_23350,N_23230,N_23225);
and U23351 (N_23351,N_23110,N_23200);
nor U23352 (N_23352,N_23148,N_23049);
and U23353 (N_23353,N_23127,N_23194);
nand U23354 (N_23354,N_23052,N_23012);
and U23355 (N_23355,N_23018,N_23039);
and U23356 (N_23356,N_23138,N_23247);
and U23357 (N_23357,N_23209,N_23152);
nor U23358 (N_23358,N_23114,N_23098);
and U23359 (N_23359,N_23234,N_23108);
and U23360 (N_23360,N_23188,N_23144);
or U23361 (N_23361,N_23111,N_23015);
or U23362 (N_23362,N_23172,N_23047);
nand U23363 (N_23363,N_23142,N_23120);
xor U23364 (N_23364,N_23145,N_23026);
and U23365 (N_23365,N_23235,N_23131);
and U23366 (N_23366,N_23042,N_23106);
and U23367 (N_23367,N_23220,N_23092);
or U23368 (N_23368,N_23139,N_23198);
and U23369 (N_23369,N_23196,N_23076);
or U23370 (N_23370,N_23084,N_23155);
xor U23371 (N_23371,N_23079,N_23169);
and U23372 (N_23372,N_23055,N_23119);
nand U23373 (N_23373,N_23183,N_23223);
or U23374 (N_23374,N_23210,N_23109);
nand U23375 (N_23375,N_23117,N_23186);
nand U23376 (N_23376,N_23066,N_23135);
nor U23377 (N_23377,N_23154,N_23245);
nand U23378 (N_23378,N_23110,N_23160);
and U23379 (N_23379,N_23089,N_23066);
nand U23380 (N_23380,N_23212,N_23123);
or U23381 (N_23381,N_23057,N_23178);
nand U23382 (N_23382,N_23170,N_23152);
and U23383 (N_23383,N_23081,N_23038);
nand U23384 (N_23384,N_23085,N_23219);
and U23385 (N_23385,N_23099,N_23146);
nor U23386 (N_23386,N_23026,N_23113);
and U23387 (N_23387,N_23225,N_23163);
or U23388 (N_23388,N_23113,N_23204);
or U23389 (N_23389,N_23227,N_23157);
nor U23390 (N_23390,N_23215,N_23122);
and U23391 (N_23391,N_23164,N_23220);
nor U23392 (N_23392,N_23036,N_23063);
nor U23393 (N_23393,N_23061,N_23013);
and U23394 (N_23394,N_23056,N_23248);
or U23395 (N_23395,N_23183,N_23160);
nor U23396 (N_23396,N_23170,N_23225);
or U23397 (N_23397,N_23119,N_23048);
and U23398 (N_23398,N_23183,N_23054);
and U23399 (N_23399,N_23208,N_23214);
and U23400 (N_23400,N_23215,N_23131);
nand U23401 (N_23401,N_23223,N_23133);
or U23402 (N_23402,N_23152,N_23074);
and U23403 (N_23403,N_23137,N_23082);
and U23404 (N_23404,N_23031,N_23008);
nand U23405 (N_23405,N_23209,N_23229);
nand U23406 (N_23406,N_23163,N_23066);
or U23407 (N_23407,N_23165,N_23234);
and U23408 (N_23408,N_23085,N_23244);
nand U23409 (N_23409,N_23235,N_23249);
or U23410 (N_23410,N_23010,N_23047);
nor U23411 (N_23411,N_23226,N_23202);
or U23412 (N_23412,N_23021,N_23130);
nor U23413 (N_23413,N_23143,N_23030);
nor U23414 (N_23414,N_23060,N_23226);
or U23415 (N_23415,N_23202,N_23225);
nor U23416 (N_23416,N_23191,N_23165);
and U23417 (N_23417,N_23147,N_23183);
nor U23418 (N_23418,N_23138,N_23219);
nor U23419 (N_23419,N_23013,N_23217);
nand U23420 (N_23420,N_23010,N_23046);
and U23421 (N_23421,N_23160,N_23025);
and U23422 (N_23422,N_23091,N_23035);
or U23423 (N_23423,N_23193,N_23199);
nor U23424 (N_23424,N_23132,N_23074);
nor U23425 (N_23425,N_23222,N_23094);
nor U23426 (N_23426,N_23189,N_23055);
and U23427 (N_23427,N_23236,N_23068);
and U23428 (N_23428,N_23108,N_23102);
and U23429 (N_23429,N_23087,N_23232);
nand U23430 (N_23430,N_23082,N_23201);
and U23431 (N_23431,N_23105,N_23182);
and U23432 (N_23432,N_23123,N_23086);
nor U23433 (N_23433,N_23212,N_23114);
or U23434 (N_23434,N_23076,N_23118);
and U23435 (N_23435,N_23029,N_23106);
nor U23436 (N_23436,N_23177,N_23151);
nand U23437 (N_23437,N_23147,N_23016);
or U23438 (N_23438,N_23154,N_23143);
and U23439 (N_23439,N_23243,N_23128);
nand U23440 (N_23440,N_23073,N_23137);
nand U23441 (N_23441,N_23006,N_23125);
or U23442 (N_23442,N_23153,N_23172);
or U23443 (N_23443,N_23197,N_23122);
and U23444 (N_23444,N_23172,N_23208);
and U23445 (N_23445,N_23004,N_23239);
nor U23446 (N_23446,N_23138,N_23017);
and U23447 (N_23447,N_23188,N_23097);
and U23448 (N_23448,N_23129,N_23079);
or U23449 (N_23449,N_23200,N_23124);
nand U23450 (N_23450,N_23068,N_23181);
and U23451 (N_23451,N_23079,N_23140);
nand U23452 (N_23452,N_23071,N_23100);
or U23453 (N_23453,N_23168,N_23085);
nand U23454 (N_23454,N_23207,N_23241);
nor U23455 (N_23455,N_23239,N_23001);
or U23456 (N_23456,N_23148,N_23063);
and U23457 (N_23457,N_23141,N_23225);
nor U23458 (N_23458,N_23104,N_23063);
nor U23459 (N_23459,N_23209,N_23053);
or U23460 (N_23460,N_23014,N_23130);
nand U23461 (N_23461,N_23088,N_23226);
and U23462 (N_23462,N_23107,N_23237);
nor U23463 (N_23463,N_23195,N_23190);
and U23464 (N_23464,N_23195,N_23102);
or U23465 (N_23465,N_23002,N_23188);
and U23466 (N_23466,N_23150,N_23005);
and U23467 (N_23467,N_23080,N_23103);
or U23468 (N_23468,N_23203,N_23084);
nand U23469 (N_23469,N_23169,N_23107);
nor U23470 (N_23470,N_23020,N_23129);
or U23471 (N_23471,N_23073,N_23199);
nor U23472 (N_23472,N_23194,N_23202);
and U23473 (N_23473,N_23119,N_23141);
nor U23474 (N_23474,N_23099,N_23248);
nor U23475 (N_23475,N_23098,N_23125);
and U23476 (N_23476,N_23070,N_23148);
nand U23477 (N_23477,N_23183,N_23226);
nor U23478 (N_23478,N_23238,N_23191);
nor U23479 (N_23479,N_23162,N_23112);
and U23480 (N_23480,N_23149,N_23238);
and U23481 (N_23481,N_23127,N_23027);
nor U23482 (N_23482,N_23097,N_23092);
or U23483 (N_23483,N_23224,N_23028);
and U23484 (N_23484,N_23107,N_23208);
and U23485 (N_23485,N_23010,N_23243);
or U23486 (N_23486,N_23142,N_23062);
nor U23487 (N_23487,N_23101,N_23067);
or U23488 (N_23488,N_23068,N_23043);
or U23489 (N_23489,N_23166,N_23200);
or U23490 (N_23490,N_23160,N_23211);
or U23491 (N_23491,N_23165,N_23183);
nand U23492 (N_23492,N_23214,N_23051);
nand U23493 (N_23493,N_23051,N_23227);
and U23494 (N_23494,N_23056,N_23174);
nand U23495 (N_23495,N_23190,N_23205);
nor U23496 (N_23496,N_23211,N_23120);
nor U23497 (N_23497,N_23050,N_23242);
nand U23498 (N_23498,N_23201,N_23135);
and U23499 (N_23499,N_23139,N_23163);
or U23500 (N_23500,N_23475,N_23480);
or U23501 (N_23501,N_23365,N_23272);
and U23502 (N_23502,N_23273,N_23461);
nor U23503 (N_23503,N_23392,N_23363);
xor U23504 (N_23504,N_23263,N_23374);
or U23505 (N_23505,N_23487,N_23427);
and U23506 (N_23506,N_23446,N_23282);
and U23507 (N_23507,N_23373,N_23401);
nand U23508 (N_23508,N_23416,N_23357);
nand U23509 (N_23509,N_23448,N_23460);
nor U23510 (N_23510,N_23425,N_23330);
nor U23511 (N_23511,N_23256,N_23474);
or U23512 (N_23512,N_23421,N_23422);
nand U23513 (N_23513,N_23499,N_23364);
nand U23514 (N_23514,N_23488,N_23483);
or U23515 (N_23515,N_23320,N_23262);
nand U23516 (N_23516,N_23289,N_23294);
nor U23517 (N_23517,N_23361,N_23465);
and U23518 (N_23518,N_23325,N_23444);
and U23519 (N_23519,N_23291,N_23267);
nand U23520 (N_23520,N_23277,N_23476);
and U23521 (N_23521,N_23259,N_23455);
nand U23522 (N_23522,N_23381,N_23472);
nor U23523 (N_23523,N_23355,N_23441);
nand U23524 (N_23524,N_23454,N_23317);
or U23525 (N_23525,N_23390,N_23346);
and U23526 (N_23526,N_23301,N_23412);
nor U23527 (N_23527,N_23459,N_23307);
or U23528 (N_23528,N_23286,N_23351);
or U23529 (N_23529,N_23309,N_23481);
nor U23530 (N_23530,N_23395,N_23464);
nand U23531 (N_23531,N_23283,N_23251);
and U23532 (N_23532,N_23398,N_23322);
or U23533 (N_23533,N_23492,N_23431);
nor U23534 (N_23534,N_23397,N_23469);
nand U23535 (N_23535,N_23336,N_23407);
nand U23536 (N_23536,N_23255,N_23359);
or U23537 (N_23537,N_23348,N_23367);
or U23538 (N_23538,N_23389,N_23478);
nor U23539 (N_23539,N_23400,N_23497);
nor U23540 (N_23540,N_23369,N_23275);
nor U23541 (N_23541,N_23423,N_23331);
nand U23542 (N_23542,N_23344,N_23276);
and U23543 (N_23543,N_23388,N_23386);
and U23544 (N_23544,N_23442,N_23350);
and U23545 (N_23545,N_23493,N_23312);
nand U23546 (N_23546,N_23266,N_23477);
xnor U23547 (N_23547,N_23304,N_23436);
nor U23548 (N_23548,N_23462,N_23486);
nand U23549 (N_23549,N_23418,N_23471);
or U23550 (N_23550,N_23385,N_23470);
and U23551 (N_23551,N_23405,N_23450);
nor U23552 (N_23552,N_23298,N_23303);
or U23553 (N_23553,N_23437,N_23340);
or U23554 (N_23554,N_23335,N_23252);
and U23555 (N_23555,N_23278,N_23473);
nand U23556 (N_23556,N_23338,N_23482);
and U23557 (N_23557,N_23353,N_23314);
or U23558 (N_23558,N_23430,N_23453);
and U23559 (N_23559,N_23270,N_23377);
nand U23560 (N_23560,N_23253,N_23484);
and U23561 (N_23561,N_23250,N_23403);
nor U23562 (N_23562,N_23349,N_23417);
nand U23563 (N_23563,N_23467,N_23409);
and U23564 (N_23564,N_23347,N_23491);
and U23565 (N_23565,N_23438,N_23457);
xnor U23566 (N_23566,N_23447,N_23415);
nand U23567 (N_23567,N_23326,N_23410);
nor U23568 (N_23568,N_23274,N_23420);
and U23569 (N_23569,N_23396,N_23424);
and U23570 (N_23570,N_23305,N_23260);
nor U23571 (N_23571,N_23362,N_23290);
nand U23572 (N_23572,N_23280,N_23258);
nor U23573 (N_23573,N_23382,N_23439);
or U23574 (N_23574,N_23321,N_23341);
nand U23575 (N_23575,N_23287,N_23449);
and U23576 (N_23576,N_23296,N_23333);
nor U23577 (N_23577,N_23408,N_23302);
nand U23578 (N_23578,N_23337,N_23281);
nand U23579 (N_23579,N_23358,N_23434);
nand U23580 (N_23580,N_23490,N_23443);
nand U23581 (N_23581,N_23285,N_23261);
nor U23582 (N_23582,N_23458,N_23393);
nand U23583 (N_23583,N_23269,N_23495);
or U23584 (N_23584,N_23257,N_23310);
nor U23585 (N_23585,N_23391,N_23496);
and U23586 (N_23586,N_23383,N_23368);
nand U23587 (N_23587,N_23354,N_23297);
nand U23588 (N_23588,N_23380,N_23378);
nand U23589 (N_23589,N_23360,N_23288);
or U23590 (N_23590,N_23295,N_23414);
nand U23591 (N_23591,N_23494,N_23463);
or U23592 (N_23592,N_23432,N_23268);
nand U23593 (N_23593,N_23334,N_23399);
nand U23594 (N_23594,N_23329,N_23429);
and U23595 (N_23595,N_23313,N_23306);
and U23596 (N_23596,N_23327,N_23379);
and U23597 (N_23597,N_23370,N_23284);
nand U23598 (N_23598,N_23428,N_23387);
and U23599 (N_23599,N_23498,N_23406);
or U23600 (N_23600,N_23489,N_23384);
and U23601 (N_23601,N_23411,N_23339);
nor U23602 (N_23602,N_23332,N_23308);
or U23603 (N_23603,N_23375,N_23479);
and U23604 (N_23604,N_23323,N_23343);
nand U23605 (N_23605,N_23402,N_23394);
nand U23606 (N_23606,N_23316,N_23371);
and U23607 (N_23607,N_23254,N_23324);
nand U23608 (N_23608,N_23413,N_23419);
nand U23609 (N_23609,N_23319,N_23356);
and U23610 (N_23610,N_23445,N_23318);
and U23611 (N_23611,N_23404,N_23299);
and U23612 (N_23612,N_23279,N_23352);
nand U23613 (N_23613,N_23345,N_23264);
and U23614 (N_23614,N_23292,N_23435);
or U23615 (N_23615,N_23466,N_23485);
and U23616 (N_23616,N_23265,N_23328);
or U23617 (N_23617,N_23426,N_23271);
and U23618 (N_23618,N_23376,N_23452);
or U23619 (N_23619,N_23300,N_23440);
nor U23620 (N_23620,N_23372,N_23433);
and U23621 (N_23621,N_23311,N_23468);
or U23622 (N_23622,N_23293,N_23451);
and U23623 (N_23623,N_23342,N_23366);
or U23624 (N_23624,N_23456,N_23315);
or U23625 (N_23625,N_23489,N_23362);
and U23626 (N_23626,N_23384,N_23396);
and U23627 (N_23627,N_23335,N_23426);
nand U23628 (N_23628,N_23441,N_23351);
nor U23629 (N_23629,N_23311,N_23393);
and U23630 (N_23630,N_23384,N_23450);
or U23631 (N_23631,N_23264,N_23291);
nand U23632 (N_23632,N_23395,N_23456);
nor U23633 (N_23633,N_23314,N_23330);
nand U23634 (N_23634,N_23297,N_23434);
xnor U23635 (N_23635,N_23328,N_23363);
and U23636 (N_23636,N_23343,N_23429);
nand U23637 (N_23637,N_23290,N_23380);
or U23638 (N_23638,N_23480,N_23445);
nand U23639 (N_23639,N_23281,N_23319);
or U23640 (N_23640,N_23378,N_23466);
nor U23641 (N_23641,N_23489,N_23466);
nand U23642 (N_23642,N_23437,N_23406);
nor U23643 (N_23643,N_23310,N_23435);
nor U23644 (N_23644,N_23352,N_23288);
nor U23645 (N_23645,N_23255,N_23441);
and U23646 (N_23646,N_23487,N_23349);
or U23647 (N_23647,N_23261,N_23299);
and U23648 (N_23648,N_23251,N_23403);
and U23649 (N_23649,N_23442,N_23433);
nor U23650 (N_23650,N_23388,N_23438);
nand U23651 (N_23651,N_23341,N_23490);
nor U23652 (N_23652,N_23326,N_23254);
or U23653 (N_23653,N_23336,N_23283);
nor U23654 (N_23654,N_23327,N_23269);
and U23655 (N_23655,N_23418,N_23422);
and U23656 (N_23656,N_23298,N_23342);
nor U23657 (N_23657,N_23285,N_23483);
or U23658 (N_23658,N_23452,N_23441);
and U23659 (N_23659,N_23280,N_23361);
nand U23660 (N_23660,N_23334,N_23474);
nand U23661 (N_23661,N_23378,N_23464);
nand U23662 (N_23662,N_23483,N_23250);
nor U23663 (N_23663,N_23401,N_23308);
nor U23664 (N_23664,N_23359,N_23274);
and U23665 (N_23665,N_23433,N_23351);
nand U23666 (N_23666,N_23389,N_23469);
and U23667 (N_23667,N_23276,N_23419);
nor U23668 (N_23668,N_23349,N_23435);
and U23669 (N_23669,N_23359,N_23494);
nor U23670 (N_23670,N_23430,N_23497);
and U23671 (N_23671,N_23288,N_23346);
nand U23672 (N_23672,N_23351,N_23298);
nor U23673 (N_23673,N_23301,N_23318);
nand U23674 (N_23674,N_23264,N_23443);
nor U23675 (N_23675,N_23306,N_23412);
and U23676 (N_23676,N_23338,N_23494);
nor U23677 (N_23677,N_23410,N_23342);
nand U23678 (N_23678,N_23494,N_23266);
or U23679 (N_23679,N_23270,N_23359);
or U23680 (N_23680,N_23498,N_23429);
and U23681 (N_23681,N_23387,N_23250);
or U23682 (N_23682,N_23403,N_23372);
and U23683 (N_23683,N_23284,N_23309);
and U23684 (N_23684,N_23408,N_23259);
and U23685 (N_23685,N_23455,N_23349);
and U23686 (N_23686,N_23457,N_23255);
nor U23687 (N_23687,N_23298,N_23432);
or U23688 (N_23688,N_23444,N_23424);
nand U23689 (N_23689,N_23304,N_23448);
nand U23690 (N_23690,N_23385,N_23360);
nor U23691 (N_23691,N_23277,N_23424);
nor U23692 (N_23692,N_23252,N_23403);
or U23693 (N_23693,N_23369,N_23425);
nand U23694 (N_23694,N_23493,N_23456);
and U23695 (N_23695,N_23339,N_23330);
or U23696 (N_23696,N_23345,N_23321);
nand U23697 (N_23697,N_23296,N_23497);
nand U23698 (N_23698,N_23456,N_23482);
nand U23699 (N_23699,N_23268,N_23353);
and U23700 (N_23700,N_23448,N_23425);
and U23701 (N_23701,N_23274,N_23334);
or U23702 (N_23702,N_23411,N_23486);
nand U23703 (N_23703,N_23418,N_23465);
and U23704 (N_23704,N_23314,N_23324);
nor U23705 (N_23705,N_23377,N_23280);
nand U23706 (N_23706,N_23472,N_23453);
nand U23707 (N_23707,N_23257,N_23453);
or U23708 (N_23708,N_23394,N_23333);
nor U23709 (N_23709,N_23354,N_23269);
and U23710 (N_23710,N_23254,N_23468);
and U23711 (N_23711,N_23385,N_23486);
nor U23712 (N_23712,N_23477,N_23491);
or U23713 (N_23713,N_23358,N_23375);
xor U23714 (N_23714,N_23487,N_23335);
nor U23715 (N_23715,N_23447,N_23369);
and U23716 (N_23716,N_23264,N_23374);
nor U23717 (N_23717,N_23365,N_23258);
or U23718 (N_23718,N_23379,N_23318);
nor U23719 (N_23719,N_23427,N_23470);
nand U23720 (N_23720,N_23422,N_23321);
nand U23721 (N_23721,N_23446,N_23479);
nand U23722 (N_23722,N_23342,N_23433);
and U23723 (N_23723,N_23268,N_23369);
or U23724 (N_23724,N_23323,N_23413);
or U23725 (N_23725,N_23417,N_23289);
nand U23726 (N_23726,N_23260,N_23332);
and U23727 (N_23727,N_23360,N_23351);
nand U23728 (N_23728,N_23356,N_23257);
nor U23729 (N_23729,N_23477,N_23432);
or U23730 (N_23730,N_23373,N_23488);
and U23731 (N_23731,N_23392,N_23413);
nand U23732 (N_23732,N_23374,N_23472);
and U23733 (N_23733,N_23352,N_23401);
or U23734 (N_23734,N_23382,N_23359);
nor U23735 (N_23735,N_23291,N_23299);
or U23736 (N_23736,N_23273,N_23329);
nor U23737 (N_23737,N_23361,N_23366);
and U23738 (N_23738,N_23469,N_23412);
nor U23739 (N_23739,N_23252,N_23493);
and U23740 (N_23740,N_23322,N_23387);
nor U23741 (N_23741,N_23446,N_23256);
and U23742 (N_23742,N_23440,N_23276);
nor U23743 (N_23743,N_23288,N_23275);
and U23744 (N_23744,N_23349,N_23463);
nor U23745 (N_23745,N_23450,N_23372);
nand U23746 (N_23746,N_23292,N_23398);
or U23747 (N_23747,N_23424,N_23386);
nor U23748 (N_23748,N_23349,N_23471);
and U23749 (N_23749,N_23340,N_23301);
nand U23750 (N_23750,N_23597,N_23732);
and U23751 (N_23751,N_23506,N_23581);
and U23752 (N_23752,N_23706,N_23702);
nand U23753 (N_23753,N_23683,N_23502);
nor U23754 (N_23754,N_23690,N_23657);
nand U23755 (N_23755,N_23640,N_23611);
or U23756 (N_23756,N_23652,N_23691);
nand U23757 (N_23757,N_23517,N_23641);
nand U23758 (N_23758,N_23610,N_23513);
nor U23759 (N_23759,N_23730,N_23606);
nand U23760 (N_23760,N_23627,N_23547);
nor U23761 (N_23761,N_23615,N_23623);
nor U23762 (N_23762,N_23625,N_23736);
nor U23763 (N_23763,N_23514,N_23582);
and U23764 (N_23764,N_23621,N_23618);
or U23765 (N_23765,N_23599,N_23649);
nor U23766 (N_23766,N_23684,N_23583);
and U23767 (N_23767,N_23563,N_23558);
or U23768 (N_23768,N_23604,N_23670);
nand U23769 (N_23769,N_23532,N_23737);
or U23770 (N_23770,N_23723,N_23603);
nor U23771 (N_23771,N_23744,N_23573);
and U23772 (N_23772,N_23725,N_23645);
and U23773 (N_23773,N_23561,N_23629);
and U23774 (N_23774,N_23659,N_23646);
or U23775 (N_23775,N_23607,N_23704);
nor U23776 (N_23776,N_23734,N_23701);
xor U23777 (N_23777,N_23520,N_23524);
nand U23778 (N_23778,N_23556,N_23507);
and U23779 (N_23779,N_23743,N_23698);
nand U23780 (N_23780,N_23576,N_23711);
nor U23781 (N_23781,N_23686,N_23504);
and U23782 (N_23782,N_23579,N_23601);
and U23783 (N_23783,N_23523,N_23567);
nor U23784 (N_23784,N_23516,N_23585);
or U23785 (N_23785,N_23674,N_23669);
and U23786 (N_23786,N_23527,N_23663);
nor U23787 (N_23787,N_23637,N_23577);
nor U23788 (N_23788,N_23694,N_23594);
and U23789 (N_23789,N_23667,N_23555);
nand U23790 (N_23790,N_23554,N_23617);
nand U23791 (N_23791,N_23720,N_23589);
nor U23792 (N_23792,N_23682,N_23644);
and U23793 (N_23793,N_23528,N_23748);
nor U23794 (N_23794,N_23501,N_23505);
nor U23795 (N_23795,N_23697,N_23733);
nor U23796 (N_23796,N_23650,N_23651);
or U23797 (N_23797,N_23551,N_23560);
or U23798 (N_23798,N_23656,N_23677);
and U23799 (N_23799,N_23535,N_23544);
nand U23800 (N_23800,N_23526,N_23689);
or U23801 (N_23801,N_23512,N_23570);
nand U23802 (N_23802,N_23643,N_23562);
or U23803 (N_23803,N_23655,N_23692);
and U23804 (N_23804,N_23566,N_23537);
or U23805 (N_23805,N_23620,N_23543);
and U23806 (N_23806,N_23545,N_23548);
and U23807 (N_23807,N_23553,N_23742);
or U23808 (N_23808,N_23578,N_23633);
or U23809 (N_23809,N_23587,N_23634);
nand U23810 (N_23810,N_23534,N_23719);
or U23811 (N_23811,N_23636,N_23500);
nor U23812 (N_23812,N_23605,N_23679);
nor U23813 (N_23813,N_23609,N_23665);
and U23814 (N_23814,N_23724,N_23681);
nand U23815 (N_23815,N_23729,N_23590);
nor U23816 (N_23816,N_23635,N_23626);
nor U23817 (N_23817,N_23592,N_23530);
and U23818 (N_23818,N_23708,N_23735);
or U23819 (N_23819,N_23675,N_23559);
nand U23820 (N_23820,N_23531,N_23678);
or U23821 (N_23821,N_23664,N_23540);
nor U23822 (N_23822,N_23613,N_23666);
or U23823 (N_23823,N_23749,N_23614);
nand U23824 (N_23824,N_23747,N_23575);
nor U23825 (N_23825,N_23713,N_23549);
or U23826 (N_23826,N_23588,N_23638);
and U23827 (N_23827,N_23726,N_23728);
nor U23828 (N_23828,N_23718,N_23557);
or U23829 (N_23829,N_23624,N_23596);
nor U23830 (N_23830,N_23565,N_23612);
or U23831 (N_23831,N_23550,N_23569);
and U23832 (N_23832,N_23510,N_23519);
or U23833 (N_23833,N_23727,N_23685);
or U23834 (N_23834,N_23695,N_23673);
and U23835 (N_23835,N_23738,N_23705);
or U23836 (N_23836,N_23511,N_23741);
and U23837 (N_23837,N_23688,N_23658);
nor U23838 (N_23838,N_23538,N_23714);
nand U23839 (N_23839,N_23696,N_23630);
or U23840 (N_23840,N_23642,N_23568);
nor U23841 (N_23841,N_23740,N_23508);
nand U23842 (N_23842,N_23653,N_23687);
nand U23843 (N_23843,N_23648,N_23572);
and U23844 (N_23844,N_23522,N_23598);
nor U23845 (N_23845,N_23717,N_23552);
or U23846 (N_23846,N_23586,N_23710);
and U23847 (N_23847,N_23716,N_23739);
nand U23848 (N_23848,N_23647,N_23542);
nor U23849 (N_23849,N_23722,N_23518);
nand U23850 (N_23850,N_23662,N_23571);
nor U23851 (N_23851,N_23593,N_23721);
or U23852 (N_23852,N_23654,N_23616);
nor U23853 (N_23853,N_23541,N_23503);
nand U23854 (N_23854,N_23703,N_23745);
and U23855 (N_23855,N_23574,N_23546);
nor U23856 (N_23856,N_23515,N_23539);
and U23857 (N_23857,N_23693,N_23564);
or U23858 (N_23858,N_23672,N_23580);
or U23859 (N_23859,N_23536,N_23715);
nor U23860 (N_23860,N_23660,N_23584);
nor U23861 (N_23861,N_23608,N_23628);
or U23862 (N_23862,N_23631,N_23619);
or U23863 (N_23863,N_23700,N_23746);
nand U23864 (N_23864,N_23602,N_23529);
nand U23865 (N_23865,N_23680,N_23668);
nor U23866 (N_23866,N_23591,N_23521);
nand U23867 (N_23867,N_23509,N_23622);
or U23868 (N_23868,N_23712,N_23671);
xnor U23869 (N_23869,N_23533,N_23525);
and U23870 (N_23870,N_23595,N_23676);
and U23871 (N_23871,N_23707,N_23632);
nand U23872 (N_23872,N_23709,N_23639);
or U23873 (N_23873,N_23661,N_23699);
nand U23874 (N_23874,N_23600,N_23731);
or U23875 (N_23875,N_23535,N_23689);
nand U23876 (N_23876,N_23621,N_23722);
nor U23877 (N_23877,N_23593,N_23748);
or U23878 (N_23878,N_23606,N_23511);
nand U23879 (N_23879,N_23679,N_23531);
nor U23880 (N_23880,N_23724,N_23737);
or U23881 (N_23881,N_23556,N_23746);
or U23882 (N_23882,N_23729,N_23515);
nor U23883 (N_23883,N_23652,N_23649);
or U23884 (N_23884,N_23606,N_23717);
and U23885 (N_23885,N_23698,N_23577);
nor U23886 (N_23886,N_23541,N_23738);
and U23887 (N_23887,N_23662,N_23584);
nor U23888 (N_23888,N_23652,N_23505);
nand U23889 (N_23889,N_23741,N_23702);
or U23890 (N_23890,N_23534,N_23563);
and U23891 (N_23891,N_23504,N_23526);
and U23892 (N_23892,N_23721,N_23728);
nor U23893 (N_23893,N_23593,N_23604);
or U23894 (N_23894,N_23505,N_23508);
or U23895 (N_23895,N_23630,N_23520);
or U23896 (N_23896,N_23713,N_23507);
xor U23897 (N_23897,N_23517,N_23684);
nand U23898 (N_23898,N_23714,N_23518);
and U23899 (N_23899,N_23668,N_23585);
nor U23900 (N_23900,N_23621,N_23516);
nand U23901 (N_23901,N_23718,N_23612);
xor U23902 (N_23902,N_23550,N_23669);
or U23903 (N_23903,N_23618,N_23719);
and U23904 (N_23904,N_23564,N_23723);
nor U23905 (N_23905,N_23626,N_23588);
nand U23906 (N_23906,N_23585,N_23603);
nor U23907 (N_23907,N_23606,N_23532);
nand U23908 (N_23908,N_23656,N_23588);
nor U23909 (N_23909,N_23536,N_23739);
nand U23910 (N_23910,N_23512,N_23710);
nand U23911 (N_23911,N_23629,N_23625);
nor U23912 (N_23912,N_23663,N_23644);
nand U23913 (N_23913,N_23529,N_23690);
and U23914 (N_23914,N_23594,N_23539);
nor U23915 (N_23915,N_23528,N_23575);
nor U23916 (N_23916,N_23589,N_23607);
nor U23917 (N_23917,N_23615,N_23515);
or U23918 (N_23918,N_23607,N_23679);
or U23919 (N_23919,N_23612,N_23674);
nand U23920 (N_23920,N_23616,N_23552);
and U23921 (N_23921,N_23637,N_23642);
nand U23922 (N_23922,N_23532,N_23564);
xor U23923 (N_23923,N_23511,N_23708);
nor U23924 (N_23924,N_23599,N_23665);
and U23925 (N_23925,N_23620,N_23717);
and U23926 (N_23926,N_23548,N_23650);
nand U23927 (N_23927,N_23747,N_23701);
and U23928 (N_23928,N_23509,N_23585);
or U23929 (N_23929,N_23707,N_23602);
and U23930 (N_23930,N_23595,N_23562);
and U23931 (N_23931,N_23515,N_23736);
and U23932 (N_23932,N_23599,N_23660);
and U23933 (N_23933,N_23637,N_23691);
nand U23934 (N_23934,N_23746,N_23644);
nor U23935 (N_23935,N_23655,N_23582);
or U23936 (N_23936,N_23699,N_23593);
and U23937 (N_23937,N_23706,N_23648);
and U23938 (N_23938,N_23525,N_23731);
nor U23939 (N_23939,N_23571,N_23624);
nor U23940 (N_23940,N_23708,N_23643);
and U23941 (N_23941,N_23557,N_23560);
nand U23942 (N_23942,N_23629,N_23689);
or U23943 (N_23943,N_23698,N_23629);
or U23944 (N_23944,N_23535,N_23586);
nand U23945 (N_23945,N_23585,N_23639);
nor U23946 (N_23946,N_23670,N_23652);
nor U23947 (N_23947,N_23528,N_23718);
and U23948 (N_23948,N_23561,N_23601);
nor U23949 (N_23949,N_23647,N_23688);
nor U23950 (N_23950,N_23704,N_23560);
and U23951 (N_23951,N_23734,N_23662);
and U23952 (N_23952,N_23601,N_23590);
or U23953 (N_23953,N_23732,N_23632);
or U23954 (N_23954,N_23535,N_23631);
nor U23955 (N_23955,N_23584,N_23598);
nor U23956 (N_23956,N_23747,N_23622);
nor U23957 (N_23957,N_23638,N_23527);
nand U23958 (N_23958,N_23565,N_23588);
nor U23959 (N_23959,N_23536,N_23534);
nand U23960 (N_23960,N_23648,N_23512);
nor U23961 (N_23961,N_23675,N_23679);
nand U23962 (N_23962,N_23740,N_23644);
nor U23963 (N_23963,N_23554,N_23556);
and U23964 (N_23964,N_23668,N_23557);
or U23965 (N_23965,N_23734,N_23725);
and U23966 (N_23966,N_23700,N_23744);
and U23967 (N_23967,N_23614,N_23708);
nor U23968 (N_23968,N_23682,N_23602);
nor U23969 (N_23969,N_23546,N_23514);
nand U23970 (N_23970,N_23594,N_23561);
nand U23971 (N_23971,N_23748,N_23586);
nand U23972 (N_23972,N_23522,N_23585);
or U23973 (N_23973,N_23600,N_23547);
and U23974 (N_23974,N_23694,N_23558);
nor U23975 (N_23975,N_23549,N_23705);
and U23976 (N_23976,N_23695,N_23538);
or U23977 (N_23977,N_23507,N_23711);
nor U23978 (N_23978,N_23653,N_23641);
nor U23979 (N_23979,N_23720,N_23639);
nor U23980 (N_23980,N_23591,N_23653);
and U23981 (N_23981,N_23547,N_23633);
nor U23982 (N_23982,N_23560,N_23647);
or U23983 (N_23983,N_23503,N_23651);
nor U23984 (N_23984,N_23514,N_23501);
or U23985 (N_23985,N_23743,N_23582);
and U23986 (N_23986,N_23593,N_23525);
nor U23987 (N_23987,N_23679,N_23594);
and U23988 (N_23988,N_23693,N_23682);
nand U23989 (N_23989,N_23511,N_23598);
and U23990 (N_23990,N_23589,N_23547);
or U23991 (N_23991,N_23742,N_23671);
and U23992 (N_23992,N_23503,N_23736);
or U23993 (N_23993,N_23656,N_23560);
nor U23994 (N_23994,N_23713,N_23727);
or U23995 (N_23995,N_23592,N_23699);
or U23996 (N_23996,N_23508,N_23659);
or U23997 (N_23997,N_23500,N_23718);
nand U23998 (N_23998,N_23544,N_23550);
nand U23999 (N_23999,N_23567,N_23671);
or U24000 (N_24000,N_23836,N_23961);
nand U24001 (N_24001,N_23766,N_23849);
nand U24002 (N_24002,N_23998,N_23823);
or U24003 (N_24003,N_23866,N_23951);
nor U24004 (N_24004,N_23964,N_23832);
nand U24005 (N_24005,N_23820,N_23932);
nor U24006 (N_24006,N_23877,N_23883);
or U24007 (N_24007,N_23830,N_23908);
nand U24008 (N_24008,N_23799,N_23874);
or U24009 (N_24009,N_23843,N_23989);
or U24010 (N_24010,N_23914,N_23927);
nand U24011 (N_24011,N_23965,N_23751);
or U24012 (N_24012,N_23783,N_23835);
or U24013 (N_24013,N_23757,N_23827);
nand U24014 (N_24014,N_23829,N_23987);
nor U24015 (N_24015,N_23966,N_23769);
nor U24016 (N_24016,N_23910,N_23756);
nor U24017 (N_24017,N_23833,N_23778);
or U24018 (N_24018,N_23846,N_23784);
nand U24019 (N_24019,N_23958,N_23868);
and U24020 (N_24020,N_23930,N_23776);
or U24021 (N_24021,N_23812,N_23762);
nand U24022 (N_24022,N_23763,N_23881);
nand U24023 (N_24023,N_23894,N_23750);
and U24024 (N_24024,N_23978,N_23925);
or U24025 (N_24025,N_23774,N_23999);
nand U24026 (N_24026,N_23882,N_23809);
and U24027 (N_24027,N_23811,N_23771);
nor U24028 (N_24028,N_23963,N_23937);
and U24029 (N_24029,N_23879,N_23845);
or U24030 (N_24030,N_23921,N_23785);
and U24031 (N_24031,N_23847,N_23788);
and U24032 (N_24032,N_23918,N_23939);
nand U24033 (N_24033,N_23828,N_23772);
and U24034 (N_24034,N_23924,N_23856);
or U24035 (N_24035,N_23972,N_23878);
nand U24036 (N_24036,N_23888,N_23831);
or U24037 (N_24037,N_23895,N_23926);
and U24038 (N_24038,N_23848,N_23897);
or U24039 (N_24039,N_23933,N_23957);
or U24040 (N_24040,N_23754,N_23816);
or U24041 (N_24041,N_23791,N_23873);
nor U24042 (N_24042,N_23867,N_23983);
nand U24043 (N_24043,N_23802,N_23949);
xor U24044 (N_24044,N_23889,N_23807);
and U24045 (N_24045,N_23923,N_23969);
nor U24046 (N_24046,N_23870,N_23980);
or U24047 (N_24047,N_23904,N_23796);
nand U24048 (N_24048,N_23821,N_23858);
nand U24049 (N_24049,N_23981,N_23907);
or U24050 (N_24050,N_23946,N_23770);
or U24051 (N_24051,N_23786,N_23941);
or U24052 (N_24052,N_23797,N_23928);
or U24053 (N_24053,N_23765,N_23901);
or U24054 (N_24054,N_23935,N_23896);
nand U24055 (N_24055,N_23768,N_23872);
or U24056 (N_24056,N_23824,N_23875);
and U24057 (N_24057,N_23902,N_23837);
or U24058 (N_24058,N_23929,N_23956);
or U24059 (N_24059,N_23947,N_23962);
and U24060 (N_24060,N_23759,N_23819);
or U24061 (N_24061,N_23931,N_23840);
nand U24062 (N_24062,N_23953,N_23991);
nor U24063 (N_24063,N_23940,N_23884);
nor U24064 (N_24064,N_23764,N_23892);
nand U24065 (N_24065,N_23942,N_23880);
nand U24066 (N_24066,N_23793,N_23917);
nand U24067 (N_24067,N_23990,N_23822);
and U24068 (N_24068,N_23876,N_23862);
nor U24069 (N_24069,N_23973,N_23825);
nor U24070 (N_24070,N_23909,N_23944);
nor U24071 (N_24071,N_23915,N_23936);
and U24072 (N_24072,N_23752,N_23992);
nand U24073 (N_24073,N_23893,N_23852);
nand U24074 (N_24074,N_23865,N_23842);
nor U24075 (N_24075,N_23859,N_23971);
or U24076 (N_24076,N_23760,N_23808);
and U24077 (N_24077,N_23781,N_23975);
nor U24078 (N_24078,N_23945,N_23974);
nand U24079 (N_24079,N_23864,N_23985);
and U24080 (N_24080,N_23948,N_23773);
nand U24081 (N_24081,N_23789,N_23993);
or U24082 (N_24082,N_23861,N_23817);
and U24083 (N_24083,N_23818,N_23871);
or U24084 (N_24084,N_23790,N_23885);
nor U24085 (N_24085,N_23954,N_23857);
nor U24086 (N_24086,N_23813,N_23806);
nand U24087 (N_24087,N_23955,N_23995);
nand U24088 (N_24088,N_23805,N_23959);
and U24089 (N_24089,N_23869,N_23795);
xor U24090 (N_24090,N_23798,N_23887);
nor U24091 (N_24091,N_23792,N_23834);
nand U24092 (N_24092,N_23758,N_23986);
nand U24093 (N_24093,N_23952,N_23838);
or U24094 (N_24094,N_23779,N_23938);
or U24095 (N_24095,N_23815,N_23968);
nand U24096 (N_24096,N_23755,N_23800);
nand U24097 (N_24097,N_23943,N_23753);
or U24098 (N_24098,N_23960,N_23919);
or U24099 (N_24099,N_23782,N_23810);
nor U24100 (N_24100,N_23922,N_23841);
or U24101 (N_24101,N_23803,N_23997);
or U24102 (N_24102,N_23905,N_23787);
nand U24103 (N_24103,N_23826,N_23839);
nand U24104 (N_24104,N_23801,N_23898);
nor U24105 (N_24105,N_23934,N_23844);
nor U24106 (N_24106,N_23775,N_23886);
nand U24107 (N_24107,N_23851,N_23967);
and U24108 (N_24108,N_23913,N_23761);
or U24109 (N_24109,N_23970,N_23920);
or U24110 (N_24110,N_23891,N_23780);
nand U24111 (N_24111,N_23984,N_23863);
or U24112 (N_24112,N_23906,N_23850);
or U24113 (N_24113,N_23994,N_23777);
or U24114 (N_24114,N_23890,N_23976);
and U24115 (N_24115,N_23814,N_23899);
nor U24116 (N_24116,N_23911,N_23979);
or U24117 (N_24117,N_23900,N_23950);
or U24118 (N_24118,N_23916,N_23860);
nand U24119 (N_24119,N_23996,N_23912);
or U24120 (N_24120,N_23804,N_23988);
and U24121 (N_24121,N_23853,N_23854);
or U24122 (N_24122,N_23977,N_23903);
or U24123 (N_24123,N_23794,N_23982);
and U24124 (N_24124,N_23767,N_23855);
nor U24125 (N_24125,N_23793,N_23857);
or U24126 (N_24126,N_23754,N_23991);
or U24127 (N_24127,N_23759,N_23997);
nor U24128 (N_24128,N_23773,N_23895);
nor U24129 (N_24129,N_23884,N_23764);
nand U24130 (N_24130,N_23826,N_23798);
and U24131 (N_24131,N_23938,N_23862);
and U24132 (N_24132,N_23755,N_23829);
nor U24133 (N_24133,N_23977,N_23985);
or U24134 (N_24134,N_23777,N_23886);
nand U24135 (N_24135,N_23964,N_23802);
and U24136 (N_24136,N_23842,N_23969);
and U24137 (N_24137,N_23809,N_23783);
or U24138 (N_24138,N_23775,N_23998);
nor U24139 (N_24139,N_23989,N_23813);
nand U24140 (N_24140,N_23991,N_23786);
nand U24141 (N_24141,N_23933,N_23821);
xor U24142 (N_24142,N_23939,N_23820);
or U24143 (N_24143,N_23908,N_23885);
nand U24144 (N_24144,N_23956,N_23814);
nand U24145 (N_24145,N_23789,N_23871);
and U24146 (N_24146,N_23750,N_23819);
nor U24147 (N_24147,N_23862,N_23954);
or U24148 (N_24148,N_23930,N_23882);
and U24149 (N_24149,N_23983,N_23960);
nor U24150 (N_24150,N_23942,N_23906);
nor U24151 (N_24151,N_23781,N_23824);
and U24152 (N_24152,N_23843,N_23807);
nand U24153 (N_24153,N_23873,N_23995);
nor U24154 (N_24154,N_23980,N_23869);
and U24155 (N_24155,N_23986,N_23904);
or U24156 (N_24156,N_23853,N_23915);
xor U24157 (N_24157,N_23966,N_23869);
nand U24158 (N_24158,N_23980,N_23903);
and U24159 (N_24159,N_23790,N_23788);
or U24160 (N_24160,N_23776,N_23867);
and U24161 (N_24161,N_23808,N_23837);
nand U24162 (N_24162,N_23827,N_23794);
nand U24163 (N_24163,N_23961,N_23975);
and U24164 (N_24164,N_23972,N_23839);
or U24165 (N_24165,N_23750,N_23940);
nor U24166 (N_24166,N_23976,N_23977);
and U24167 (N_24167,N_23935,N_23868);
nor U24168 (N_24168,N_23928,N_23862);
nor U24169 (N_24169,N_23959,N_23789);
nor U24170 (N_24170,N_23777,N_23961);
and U24171 (N_24171,N_23752,N_23912);
nand U24172 (N_24172,N_23769,N_23773);
and U24173 (N_24173,N_23826,N_23922);
nand U24174 (N_24174,N_23847,N_23855);
and U24175 (N_24175,N_23756,N_23991);
and U24176 (N_24176,N_23790,N_23755);
or U24177 (N_24177,N_23921,N_23954);
xnor U24178 (N_24178,N_23821,N_23929);
or U24179 (N_24179,N_23869,N_23752);
nor U24180 (N_24180,N_23797,N_23794);
nand U24181 (N_24181,N_23889,N_23997);
nor U24182 (N_24182,N_23880,N_23809);
and U24183 (N_24183,N_23858,N_23792);
or U24184 (N_24184,N_23855,N_23969);
nor U24185 (N_24185,N_23990,N_23950);
and U24186 (N_24186,N_23978,N_23837);
or U24187 (N_24187,N_23757,N_23989);
and U24188 (N_24188,N_23834,N_23887);
or U24189 (N_24189,N_23866,N_23875);
nor U24190 (N_24190,N_23753,N_23896);
nand U24191 (N_24191,N_23761,N_23993);
and U24192 (N_24192,N_23997,N_23988);
nor U24193 (N_24193,N_23833,N_23840);
nor U24194 (N_24194,N_23797,N_23904);
nand U24195 (N_24195,N_23795,N_23872);
and U24196 (N_24196,N_23908,N_23842);
or U24197 (N_24197,N_23775,N_23779);
and U24198 (N_24198,N_23877,N_23993);
xor U24199 (N_24199,N_23897,N_23814);
or U24200 (N_24200,N_23812,N_23754);
nand U24201 (N_24201,N_23801,N_23904);
nand U24202 (N_24202,N_23886,N_23837);
or U24203 (N_24203,N_23816,N_23814);
nor U24204 (N_24204,N_23758,N_23948);
or U24205 (N_24205,N_23975,N_23778);
or U24206 (N_24206,N_23803,N_23893);
and U24207 (N_24207,N_23770,N_23758);
nand U24208 (N_24208,N_23897,N_23792);
or U24209 (N_24209,N_23776,N_23841);
nand U24210 (N_24210,N_23754,N_23908);
and U24211 (N_24211,N_23778,N_23899);
or U24212 (N_24212,N_23891,N_23974);
and U24213 (N_24213,N_23796,N_23895);
or U24214 (N_24214,N_23851,N_23997);
and U24215 (N_24215,N_23890,N_23979);
or U24216 (N_24216,N_23967,N_23798);
and U24217 (N_24217,N_23988,N_23768);
or U24218 (N_24218,N_23844,N_23978);
nor U24219 (N_24219,N_23953,N_23777);
and U24220 (N_24220,N_23765,N_23825);
nor U24221 (N_24221,N_23856,N_23932);
and U24222 (N_24222,N_23866,N_23854);
nand U24223 (N_24223,N_23771,N_23815);
or U24224 (N_24224,N_23775,N_23838);
and U24225 (N_24225,N_23815,N_23831);
nand U24226 (N_24226,N_23959,N_23996);
and U24227 (N_24227,N_23808,N_23963);
or U24228 (N_24228,N_23800,N_23777);
or U24229 (N_24229,N_23801,N_23833);
nand U24230 (N_24230,N_23858,N_23966);
nand U24231 (N_24231,N_23834,N_23799);
and U24232 (N_24232,N_23781,N_23940);
and U24233 (N_24233,N_23905,N_23826);
or U24234 (N_24234,N_23843,N_23793);
nor U24235 (N_24235,N_23825,N_23788);
nand U24236 (N_24236,N_23818,N_23791);
or U24237 (N_24237,N_23861,N_23847);
nor U24238 (N_24238,N_23959,N_23985);
nor U24239 (N_24239,N_23983,N_23874);
nand U24240 (N_24240,N_23968,N_23778);
nor U24241 (N_24241,N_23872,N_23983);
nor U24242 (N_24242,N_23945,N_23969);
and U24243 (N_24243,N_23801,N_23754);
and U24244 (N_24244,N_23951,N_23931);
nor U24245 (N_24245,N_23757,N_23868);
nand U24246 (N_24246,N_23937,N_23951);
nor U24247 (N_24247,N_23990,N_23995);
or U24248 (N_24248,N_23955,N_23968);
nand U24249 (N_24249,N_23955,N_23761);
nand U24250 (N_24250,N_24100,N_24126);
nand U24251 (N_24251,N_24074,N_24080);
nand U24252 (N_24252,N_24248,N_24067);
nor U24253 (N_24253,N_24240,N_24024);
nand U24254 (N_24254,N_24028,N_24189);
or U24255 (N_24255,N_24236,N_24219);
or U24256 (N_24256,N_24031,N_24002);
nand U24257 (N_24257,N_24192,N_24018);
or U24258 (N_24258,N_24165,N_24150);
and U24259 (N_24259,N_24110,N_24178);
nand U24260 (N_24260,N_24147,N_24224);
and U24261 (N_24261,N_24006,N_24191);
and U24262 (N_24262,N_24141,N_24013);
nor U24263 (N_24263,N_24144,N_24016);
and U24264 (N_24264,N_24133,N_24057);
or U24265 (N_24265,N_24123,N_24140);
nand U24266 (N_24266,N_24233,N_24156);
nand U24267 (N_24267,N_24217,N_24047);
or U24268 (N_24268,N_24188,N_24004);
and U24269 (N_24269,N_24201,N_24120);
or U24270 (N_24270,N_24174,N_24102);
and U24271 (N_24271,N_24075,N_24104);
or U24272 (N_24272,N_24220,N_24081);
or U24273 (N_24273,N_24161,N_24235);
nor U24274 (N_24274,N_24051,N_24181);
and U24275 (N_24275,N_24000,N_24227);
or U24276 (N_24276,N_24148,N_24089);
and U24277 (N_24277,N_24158,N_24135);
or U24278 (N_24278,N_24115,N_24244);
nor U24279 (N_24279,N_24033,N_24097);
nand U24280 (N_24280,N_24059,N_24096);
and U24281 (N_24281,N_24228,N_24182);
or U24282 (N_24282,N_24054,N_24014);
and U24283 (N_24283,N_24169,N_24106);
nand U24284 (N_24284,N_24091,N_24105);
nand U24285 (N_24285,N_24194,N_24122);
and U24286 (N_24286,N_24160,N_24037);
and U24287 (N_24287,N_24211,N_24232);
or U24288 (N_24288,N_24116,N_24168);
nand U24289 (N_24289,N_24060,N_24107);
nor U24290 (N_24290,N_24172,N_24086);
or U24291 (N_24291,N_24173,N_24242);
nor U24292 (N_24292,N_24114,N_24222);
nor U24293 (N_24293,N_24132,N_24163);
and U24294 (N_24294,N_24177,N_24125);
and U24295 (N_24295,N_24069,N_24052);
and U24296 (N_24296,N_24195,N_24185);
and U24297 (N_24297,N_24022,N_24078);
nor U24298 (N_24298,N_24076,N_24119);
nor U24299 (N_24299,N_24036,N_24111);
or U24300 (N_24300,N_24130,N_24246);
or U24301 (N_24301,N_24044,N_24193);
or U24302 (N_24302,N_24145,N_24001);
and U24303 (N_24303,N_24103,N_24070);
nand U24304 (N_24304,N_24046,N_24085);
nand U24305 (N_24305,N_24143,N_24127);
and U24306 (N_24306,N_24061,N_24179);
or U24307 (N_24307,N_24056,N_24093);
nor U24308 (N_24308,N_24108,N_24050);
nor U24309 (N_24309,N_24084,N_24011);
and U24310 (N_24310,N_24071,N_24058);
and U24311 (N_24311,N_24162,N_24212);
or U24312 (N_24312,N_24009,N_24041);
nor U24313 (N_24313,N_24138,N_24010);
and U24314 (N_24314,N_24208,N_24083);
or U24315 (N_24315,N_24077,N_24203);
nor U24316 (N_24316,N_24207,N_24053);
nand U24317 (N_24317,N_24021,N_24007);
and U24318 (N_24318,N_24237,N_24247);
or U24319 (N_24319,N_24038,N_24099);
and U24320 (N_24320,N_24230,N_24090);
or U24321 (N_24321,N_24205,N_24012);
or U24322 (N_24322,N_24095,N_24213);
and U24323 (N_24323,N_24063,N_24045);
nand U24324 (N_24324,N_24226,N_24048);
and U24325 (N_24325,N_24094,N_24197);
or U24326 (N_24326,N_24043,N_24055);
or U24327 (N_24327,N_24079,N_24129);
and U24328 (N_24328,N_24154,N_24015);
xor U24329 (N_24329,N_24131,N_24020);
nor U24330 (N_24330,N_24124,N_24121);
nor U24331 (N_24331,N_24152,N_24239);
nand U24332 (N_24332,N_24029,N_24101);
xnor U24333 (N_24333,N_24146,N_24068);
nor U24334 (N_24334,N_24249,N_24064);
and U24335 (N_24335,N_24164,N_24032);
nand U24336 (N_24336,N_24109,N_24087);
or U24337 (N_24337,N_24238,N_24034);
nand U24338 (N_24338,N_24196,N_24088);
or U24339 (N_24339,N_24128,N_24082);
nor U24340 (N_24340,N_24215,N_24072);
and U24341 (N_24341,N_24204,N_24118);
and U24342 (N_24342,N_24170,N_24030);
or U24343 (N_24343,N_24026,N_24035);
or U24344 (N_24344,N_24065,N_24008);
and U24345 (N_24345,N_24200,N_24223);
nand U24346 (N_24346,N_24202,N_24159);
and U24347 (N_24347,N_24042,N_24025);
or U24348 (N_24348,N_24184,N_24112);
or U24349 (N_24349,N_24183,N_24136);
and U24350 (N_24350,N_24005,N_24229);
and U24351 (N_24351,N_24199,N_24216);
or U24352 (N_24352,N_24003,N_24098);
and U24353 (N_24353,N_24231,N_24073);
or U24354 (N_24354,N_24151,N_24049);
and U24355 (N_24355,N_24198,N_24218);
and U24356 (N_24356,N_24190,N_24066);
or U24357 (N_24357,N_24062,N_24092);
or U24358 (N_24358,N_24241,N_24149);
nor U24359 (N_24359,N_24023,N_24019);
nand U24360 (N_24360,N_24243,N_24153);
nand U24361 (N_24361,N_24187,N_24027);
and U24362 (N_24362,N_24157,N_24155);
nand U24363 (N_24363,N_24040,N_24142);
or U24364 (N_24364,N_24117,N_24214);
and U24365 (N_24365,N_24221,N_24176);
nand U24366 (N_24366,N_24113,N_24017);
nand U24367 (N_24367,N_24167,N_24186);
and U24368 (N_24368,N_24166,N_24206);
or U24369 (N_24369,N_24209,N_24234);
or U24370 (N_24370,N_24137,N_24171);
nor U24371 (N_24371,N_24210,N_24180);
nand U24372 (N_24372,N_24139,N_24245);
nor U24373 (N_24373,N_24039,N_24175);
and U24374 (N_24374,N_24225,N_24134);
and U24375 (N_24375,N_24142,N_24189);
nand U24376 (N_24376,N_24186,N_24088);
nor U24377 (N_24377,N_24075,N_24182);
and U24378 (N_24378,N_24224,N_24140);
and U24379 (N_24379,N_24129,N_24218);
or U24380 (N_24380,N_24168,N_24143);
nor U24381 (N_24381,N_24064,N_24149);
or U24382 (N_24382,N_24062,N_24198);
nor U24383 (N_24383,N_24144,N_24209);
and U24384 (N_24384,N_24135,N_24209);
or U24385 (N_24385,N_24179,N_24088);
nor U24386 (N_24386,N_24238,N_24026);
and U24387 (N_24387,N_24220,N_24071);
and U24388 (N_24388,N_24036,N_24098);
nor U24389 (N_24389,N_24088,N_24004);
nand U24390 (N_24390,N_24172,N_24145);
or U24391 (N_24391,N_24000,N_24191);
nor U24392 (N_24392,N_24077,N_24078);
or U24393 (N_24393,N_24021,N_24115);
nor U24394 (N_24394,N_24117,N_24227);
and U24395 (N_24395,N_24027,N_24046);
and U24396 (N_24396,N_24116,N_24016);
or U24397 (N_24397,N_24014,N_24229);
nor U24398 (N_24398,N_24118,N_24224);
nand U24399 (N_24399,N_24183,N_24015);
nand U24400 (N_24400,N_24020,N_24245);
nand U24401 (N_24401,N_24089,N_24205);
nor U24402 (N_24402,N_24079,N_24190);
and U24403 (N_24403,N_24008,N_24134);
or U24404 (N_24404,N_24241,N_24145);
or U24405 (N_24405,N_24113,N_24185);
nor U24406 (N_24406,N_24118,N_24002);
and U24407 (N_24407,N_24204,N_24155);
and U24408 (N_24408,N_24203,N_24213);
nand U24409 (N_24409,N_24214,N_24015);
nor U24410 (N_24410,N_24173,N_24166);
and U24411 (N_24411,N_24157,N_24099);
or U24412 (N_24412,N_24242,N_24001);
or U24413 (N_24413,N_24042,N_24243);
nor U24414 (N_24414,N_24091,N_24134);
or U24415 (N_24415,N_24103,N_24089);
nor U24416 (N_24416,N_24077,N_24213);
and U24417 (N_24417,N_24135,N_24098);
or U24418 (N_24418,N_24242,N_24089);
nor U24419 (N_24419,N_24091,N_24138);
nand U24420 (N_24420,N_24028,N_24077);
nor U24421 (N_24421,N_24157,N_24076);
nor U24422 (N_24422,N_24021,N_24238);
and U24423 (N_24423,N_24180,N_24118);
nor U24424 (N_24424,N_24187,N_24190);
and U24425 (N_24425,N_24108,N_24246);
or U24426 (N_24426,N_24226,N_24133);
nor U24427 (N_24427,N_24086,N_24236);
or U24428 (N_24428,N_24044,N_24121);
nor U24429 (N_24429,N_24200,N_24061);
xor U24430 (N_24430,N_24184,N_24072);
nand U24431 (N_24431,N_24041,N_24044);
and U24432 (N_24432,N_24205,N_24041);
nor U24433 (N_24433,N_24159,N_24077);
and U24434 (N_24434,N_24026,N_24208);
nor U24435 (N_24435,N_24149,N_24063);
nor U24436 (N_24436,N_24036,N_24169);
or U24437 (N_24437,N_24106,N_24191);
nor U24438 (N_24438,N_24186,N_24099);
nor U24439 (N_24439,N_24161,N_24139);
or U24440 (N_24440,N_24174,N_24143);
and U24441 (N_24441,N_24142,N_24166);
nand U24442 (N_24442,N_24161,N_24176);
and U24443 (N_24443,N_24059,N_24141);
and U24444 (N_24444,N_24212,N_24157);
nand U24445 (N_24445,N_24051,N_24246);
nand U24446 (N_24446,N_24004,N_24010);
nor U24447 (N_24447,N_24144,N_24240);
or U24448 (N_24448,N_24136,N_24139);
nor U24449 (N_24449,N_24168,N_24056);
and U24450 (N_24450,N_24227,N_24160);
and U24451 (N_24451,N_24153,N_24127);
nor U24452 (N_24452,N_24208,N_24087);
nand U24453 (N_24453,N_24004,N_24092);
and U24454 (N_24454,N_24001,N_24240);
nor U24455 (N_24455,N_24031,N_24244);
or U24456 (N_24456,N_24101,N_24157);
or U24457 (N_24457,N_24127,N_24202);
nand U24458 (N_24458,N_24069,N_24161);
or U24459 (N_24459,N_24106,N_24001);
nand U24460 (N_24460,N_24061,N_24131);
nor U24461 (N_24461,N_24083,N_24134);
or U24462 (N_24462,N_24079,N_24051);
and U24463 (N_24463,N_24235,N_24017);
nand U24464 (N_24464,N_24086,N_24022);
nor U24465 (N_24465,N_24197,N_24167);
nand U24466 (N_24466,N_24241,N_24065);
nand U24467 (N_24467,N_24222,N_24178);
and U24468 (N_24468,N_24140,N_24025);
nand U24469 (N_24469,N_24031,N_24217);
or U24470 (N_24470,N_24036,N_24091);
nor U24471 (N_24471,N_24076,N_24060);
nor U24472 (N_24472,N_24008,N_24154);
nand U24473 (N_24473,N_24153,N_24103);
and U24474 (N_24474,N_24219,N_24127);
nand U24475 (N_24475,N_24100,N_24239);
nor U24476 (N_24476,N_24160,N_24214);
nor U24477 (N_24477,N_24151,N_24226);
or U24478 (N_24478,N_24053,N_24215);
nor U24479 (N_24479,N_24115,N_24222);
nand U24480 (N_24480,N_24083,N_24027);
or U24481 (N_24481,N_24137,N_24240);
or U24482 (N_24482,N_24098,N_24170);
and U24483 (N_24483,N_24111,N_24093);
and U24484 (N_24484,N_24167,N_24036);
and U24485 (N_24485,N_24117,N_24236);
nand U24486 (N_24486,N_24170,N_24074);
nand U24487 (N_24487,N_24094,N_24247);
nor U24488 (N_24488,N_24119,N_24106);
nor U24489 (N_24489,N_24109,N_24063);
and U24490 (N_24490,N_24180,N_24160);
or U24491 (N_24491,N_24031,N_24046);
nand U24492 (N_24492,N_24238,N_24014);
nor U24493 (N_24493,N_24049,N_24086);
nand U24494 (N_24494,N_24249,N_24076);
or U24495 (N_24495,N_24041,N_24242);
nor U24496 (N_24496,N_24126,N_24028);
or U24497 (N_24497,N_24118,N_24141);
nor U24498 (N_24498,N_24099,N_24152);
and U24499 (N_24499,N_24172,N_24162);
nand U24500 (N_24500,N_24460,N_24340);
or U24501 (N_24501,N_24353,N_24393);
and U24502 (N_24502,N_24292,N_24435);
or U24503 (N_24503,N_24333,N_24357);
or U24504 (N_24504,N_24411,N_24322);
or U24505 (N_24505,N_24402,N_24277);
nand U24506 (N_24506,N_24406,N_24485);
or U24507 (N_24507,N_24397,N_24455);
nor U24508 (N_24508,N_24434,N_24308);
and U24509 (N_24509,N_24414,N_24392);
nor U24510 (N_24510,N_24454,N_24334);
nand U24511 (N_24511,N_24264,N_24358);
or U24512 (N_24512,N_24461,N_24428);
nand U24513 (N_24513,N_24294,N_24363);
or U24514 (N_24514,N_24272,N_24463);
and U24515 (N_24515,N_24360,N_24429);
or U24516 (N_24516,N_24490,N_24419);
xor U24517 (N_24517,N_24315,N_24251);
nor U24518 (N_24518,N_24332,N_24499);
nor U24519 (N_24519,N_24316,N_24314);
nand U24520 (N_24520,N_24293,N_24327);
nor U24521 (N_24521,N_24346,N_24278);
and U24522 (N_24522,N_24412,N_24443);
or U24523 (N_24523,N_24386,N_24341);
nand U24524 (N_24524,N_24480,N_24469);
or U24525 (N_24525,N_24311,N_24389);
and U24526 (N_24526,N_24351,N_24288);
nand U24527 (N_24527,N_24262,N_24255);
nand U24528 (N_24528,N_24296,N_24440);
or U24529 (N_24529,N_24398,N_24487);
or U24530 (N_24530,N_24467,N_24457);
or U24531 (N_24531,N_24298,N_24422);
or U24532 (N_24532,N_24361,N_24410);
nand U24533 (N_24533,N_24374,N_24376);
nor U24534 (N_24534,N_24498,N_24491);
or U24535 (N_24535,N_24330,N_24381);
nand U24536 (N_24536,N_24415,N_24405);
or U24537 (N_24537,N_24365,N_24470);
nor U24538 (N_24538,N_24475,N_24369);
nand U24539 (N_24539,N_24441,N_24489);
nand U24540 (N_24540,N_24328,N_24399);
and U24541 (N_24541,N_24452,N_24382);
and U24542 (N_24542,N_24342,N_24312);
nor U24543 (N_24543,N_24418,N_24484);
nor U24544 (N_24544,N_24413,N_24466);
nand U24545 (N_24545,N_24305,N_24432);
nor U24546 (N_24546,N_24362,N_24323);
or U24547 (N_24547,N_24396,N_24430);
or U24548 (N_24548,N_24377,N_24338);
nand U24549 (N_24549,N_24453,N_24462);
nand U24550 (N_24550,N_24404,N_24364);
nor U24551 (N_24551,N_24492,N_24437);
nor U24552 (N_24552,N_24421,N_24426);
nor U24553 (N_24553,N_24252,N_24354);
or U24554 (N_24554,N_24335,N_24494);
and U24555 (N_24555,N_24408,N_24456);
nand U24556 (N_24556,N_24486,N_24446);
and U24557 (N_24557,N_24303,N_24263);
or U24558 (N_24558,N_24451,N_24458);
nor U24559 (N_24559,N_24331,N_24258);
nor U24560 (N_24560,N_24250,N_24481);
and U24561 (N_24561,N_24472,N_24395);
and U24562 (N_24562,N_24387,N_24479);
and U24563 (N_24563,N_24468,N_24326);
nor U24564 (N_24564,N_24299,N_24478);
and U24565 (N_24565,N_24266,N_24254);
nand U24566 (N_24566,N_24496,N_24319);
and U24567 (N_24567,N_24442,N_24465);
nor U24568 (N_24568,N_24269,N_24268);
nor U24569 (N_24569,N_24257,N_24459);
or U24570 (N_24570,N_24420,N_24276);
nand U24571 (N_24571,N_24444,N_24271);
and U24572 (N_24572,N_24388,N_24321);
or U24573 (N_24573,N_24380,N_24337);
or U24574 (N_24574,N_24253,N_24476);
nand U24575 (N_24575,N_24306,N_24345);
or U24576 (N_24576,N_24291,N_24400);
or U24577 (N_24577,N_24401,N_24290);
or U24578 (N_24578,N_24347,N_24301);
nand U24579 (N_24579,N_24371,N_24403);
and U24580 (N_24580,N_24273,N_24320);
and U24581 (N_24581,N_24495,N_24355);
or U24582 (N_24582,N_24416,N_24394);
nor U24583 (N_24583,N_24309,N_24493);
and U24584 (N_24584,N_24431,N_24307);
nor U24585 (N_24585,N_24438,N_24280);
or U24586 (N_24586,N_24448,N_24267);
and U24587 (N_24587,N_24433,N_24318);
nor U24588 (N_24588,N_24281,N_24447);
nand U24589 (N_24589,N_24259,N_24350);
and U24590 (N_24590,N_24317,N_24423);
and U24591 (N_24591,N_24283,N_24450);
nand U24592 (N_24592,N_24379,N_24297);
nand U24593 (N_24593,N_24343,N_24324);
and U24594 (N_24594,N_24424,N_24390);
nor U24595 (N_24595,N_24329,N_24336);
and U24596 (N_24596,N_24284,N_24449);
nor U24597 (N_24597,N_24310,N_24407);
or U24598 (N_24598,N_24482,N_24473);
and U24599 (N_24599,N_24425,N_24352);
and U24600 (N_24600,N_24367,N_24282);
and U24601 (N_24601,N_24391,N_24471);
nand U24602 (N_24602,N_24265,N_24445);
nand U24603 (N_24603,N_24295,N_24274);
and U24604 (N_24604,N_24409,N_24261);
nor U24605 (N_24605,N_24488,N_24373);
nand U24606 (N_24606,N_24287,N_24436);
or U24607 (N_24607,N_24464,N_24370);
nor U24608 (N_24608,N_24348,N_24325);
or U24609 (N_24609,N_24366,N_24417);
nor U24610 (N_24610,N_24286,N_24304);
nor U24611 (N_24611,N_24300,N_24439);
or U24612 (N_24612,N_24270,N_24356);
nand U24613 (N_24613,N_24427,N_24260);
or U24614 (N_24614,N_24289,N_24313);
nor U24615 (N_24615,N_24477,N_24368);
nand U24616 (N_24616,N_24275,N_24349);
nand U24617 (N_24617,N_24383,N_24339);
nor U24618 (N_24618,N_24344,N_24378);
and U24619 (N_24619,N_24474,N_24279);
nand U24620 (N_24620,N_24359,N_24285);
or U24621 (N_24621,N_24256,N_24384);
nor U24622 (N_24622,N_24385,N_24497);
nand U24623 (N_24623,N_24375,N_24372);
or U24624 (N_24624,N_24483,N_24302);
nor U24625 (N_24625,N_24461,N_24424);
nor U24626 (N_24626,N_24260,N_24382);
nor U24627 (N_24627,N_24441,N_24250);
or U24628 (N_24628,N_24410,N_24375);
nor U24629 (N_24629,N_24474,N_24467);
nand U24630 (N_24630,N_24384,N_24319);
nand U24631 (N_24631,N_24444,N_24339);
nand U24632 (N_24632,N_24468,N_24306);
and U24633 (N_24633,N_24373,N_24399);
nand U24634 (N_24634,N_24496,N_24392);
and U24635 (N_24635,N_24376,N_24425);
nand U24636 (N_24636,N_24262,N_24381);
and U24637 (N_24637,N_24476,N_24459);
nand U24638 (N_24638,N_24356,N_24391);
and U24639 (N_24639,N_24372,N_24456);
or U24640 (N_24640,N_24291,N_24371);
or U24641 (N_24641,N_24282,N_24269);
nor U24642 (N_24642,N_24328,N_24353);
or U24643 (N_24643,N_24360,N_24494);
and U24644 (N_24644,N_24398,N_24463);
and U24645 (N_24645,N_24258,N_24449);
xnor U24646 (N_24646,N_24380,N_24323);
and U24647 (N_24647,N_24304,N_24405);
nor U24648 (N_24648,N_24311,N_24285);
or U24649 (N_24649,N_24302,N_24337);
nor U24650 (N_24650,N_24441,N_24439);
nor U24651 (N_24651,N_24413,N_24397);
nand U24652 (N_24652,N_24478,N_24287);
nand U24653 (N_24653,N_24381,N_24439);
nand U24654 (N_24654,N_24403,N_24336);
nor U24655 (N_24655,N_24450,N_24293);
nand U24656 (N_24656,N_24330,N_24417);
and U24657 (N_24657,N_24365,N_24270);
xor U24658 (N_24658,N_24371,N_24411);
and U24659 (N_24659,N_24359,N_24447);
and U24660 (N_24660,N_24454,N_24250);
nand U24661 (N_24661,N_24329,N_24282);
nand U24662 (N_24662,N_24426,N_24468);
nor U24663 (N_24663,N_24400,N_24475);
or U24664 (N_24664,N_24491,N_24417);
and U24665 (N_24665,N_24284,N_24259);
or U24666 (N_24666,N_24493,N_24282);
or U24667 (N_24667,N_24465,N_24256);
nor U24668 (N_24668,N_24376,N_24369);
or U24669 (N_24669,N_24372,N_24379);
nor U24670 (N_24670,N_24491,N_24256);
or U24671 (N_24671,N_24272,N_24394);
nor U24672 (N_24672,N_24443,N_24327);
or U24673 (N_24673,N_24436,N_24298);
or U24674 (N_24674,N_24391,N_24372);
nor U24675 (N_24675,N_24335,N_24337);
nand U24676 (N_24676,N_24302,N_24277);
and U24677 (N_24677,N_24429,N_24269);
and U24678 (N_24678,N_24390,N_24296);
nand U24679 (N_24679,N_24322,N_24433);
nor U24680 (N_24680,N_24275,N_24421);
nand U24681 (N_24681,N_24311,N_24451);
nand U24682 (N_24682,N_24433,N_24389);
or U24683 (N_24683,N_24460,N_24448);
or U24684 (N_24684,N_24361,N_24411);
or U24685 (N_24685,N_24379,N_24465);
nand U24686 (N_24686,N_24354,N_24420);
nor U24687 (N_24687,N_24491,N_24291);
xor U24688 (N_24688,N_24316,N_24461);
nor U24689 (N_24689,N_24293,N_24267);
or U24690 (N_24690,N_24289,N_24470);
and U24691 (N_24691,N_24339,N_24334);
and U24692 (N_24692,N_24331,N_24476);
nor U24693 (N_24693,N_24270,N_24272);
nand U24694 (N_24694,N_24407,N_24481);
nand U24695 (N_24695,N_24320,N_24337);
or U24696 (N_24696,N_24360,N_24267);
or U24697 (N_24697,N_24290,N_24333);
or U24698 (N_24698,N_24484,N_24494);
nand U24699 (N_24699,N_24310,N_24482);
nor U24700 (N_24700,N_24310,N_24398);
nand U24701 (N_24701,N_24329,N_24328);
and U24702 (N_24702,N_24428,N_24427);
and U24703 (N_24703,N_24299,N_24464);
nor U24704 (N_24704,N_24275,N_24444);
nand U24705 (N_24705,N_24374,N_24385);
nor U24706 (N_24706,N_24396,N_24321);
or U24707 (N_24707,N_24421,N_24285);
nor U24708 (N_24708,N_24354,N_24427);
or U24709 (N_24709,N_24385,N_24489);
nor U24710 (N_24710,N_24489,N_24285);
or U24711 (N_24711,N_24255,N_24363);
or U24712 (N_24712,N_24432,N_24467);
nand U24713 (N_24713,N_24407,N_24328);
and U24714 (N_24714,N_24359,N_24376);
and U24715 (N_24715,N_24412,N_24490);
nand U24716 (N_24716,N_24337,N_24358);
nor U24717 (N_24717,N_24309,N_24474);
or U24718 (N_24718,N_24490,N_24497);
or U24719 (N_24719,N_24313,N_24459);
nand U24720 (N_24720,N_24254,N_24323);
nor U24721 (N_24721,N_24498,N_24471);
or U24722 (N_24722,N_24355,N_24359);
and U24723 (N_24723,N_24326,N_24441);
nor U24724 (N_24724,N_24477,N_24440);
and U24725 (N_24725,N_24492,N_24459);
and U24726 (N_24726,N_24307,N_24330);
and U24727 (N_24727,N_24256,N_24267);
and U24728 (N_24728,N_24476,N_24456);
or U24729 (N_24729,N_24340,N_24412);
or U24730 (N_24730,N_24317,N_24309);
nor U24731 (N_24731,N_24437,N_24351);
nand U24732 (N_24732,N_24444,N_24483);
nand U24733 (N_24733,N_24414,N_24252);
and U24734 (N_24734,N_24306,N_24254);
or U24735 (N_24735,N_24394,N_24424);
or U24736 (N_24736,N_24444,N_24476);
nor U24737 (N_24737,N_24364,N_24329);
and U24738 (N_24738,N_24416,N_24412);
and U24739 (N_24739,N_24328,N_24378);
nand U24740 (N_24740,N_24373,N_24351);
or U24741 (N_24741,N_24311,N_24268);
nand U24742 (N_24742,N_24277,N_24466);
and U24743 (N_24743,N_24483,N_24487);
nand U24744 (N_24744,N_24463,N_24410);
and U24745 (N_24745,N_24426,N_24325);
nor U24746 (N_24746,N_24277,N_24350);
nand U24747 (N_24747,N_24322,N_24388);
and U24748 (N_24748,N_24298,N_24346);
and U24749 (N_24749,N_24367,N_24469);
and U24750 (N_24750,N_24669,N_24556);
or U24751 (N_24751,N_24642,N_24675);
and U24752 (N_24752,N_24531,N_24581);
and U24753 (N_24753,N_24664,N_24717);
nor U24754 (N_24754,N_24706,N_24626);
or U24755 (N_24755,N_24627,N_24588);
nand U24756 (N_24756,N_24644,N_24598);
nor U24757 (N_24757,N_24557,N_24618);
xor U24758 (N_24758,N_24682,N_24502);
nand U24759 (N_24759,N_24635,N_24668);
or U24760 (N_24760,N_24736,N_24575);
nand U24761 (N_24761,N_24729,N_24580);
or U24762 (N_24762,N_24709,N_24564);
nor U24763 (N_24763,N_24689,N_24503);
nor U24764 (N_24764,N_24551,N_24552);
nand U24765 (N_24765,N_24590,N_24704);
nor U24766 (N_24766,N_24585,N_24624);
and U24767 (N_24767,N_24631,N_24587);
and U24768 (N_24768,N_24549,N_24607);
nor U24769 (N_24769,N_24544,N_24659);
and U24770 (N_24770,N_24534,N_24600);
or U24771 (N_24771,N_24604,N_24529);
or U24772 (N_24772,N_24539,N_24686);
nor U24773 (N_24773,N_24672,N_24712);
nand U24774 (N_24774,N_24540,N_24730);
or U24775 (N_24775,N_24743,N_24608);
and U24776 (N_24776,N_24514,N_24542);
or U24777 (N_24777,N_24578,N_24696);
nand U24778 (N_24778,N_24545,N_24654);
and U24779 (N_24779,N_24550,N_24603);
nand U24780 (N_24780,N_24582,N_24638);
or U24781 (N_24781,N_24700,N_24636);
nor U24782 (N_24782,N_24733,N_24667);
or U24783 (N_24783,N_24630,N_24525);
nor U24784 (N_24784,N_24538,N_24698);
or U24785 (N_24785,N_24732,N_24537);
nand U24786 (N_24786,N_24504,N_24524);
or U24787 (N_24787,N_24715,N_24719);
nor U24788 (N_24788,N_24740,N_24532);
nor U24789 (N_24789,N_24513,N_24708);
nor U24790 (N_24790,N_24727,N_24560);
and U24791 (N_24791,N_24593,N_24623);
and U24792 (N_24792,N_24597,N_24703);
nor U24793 (N_24793,N_24613,N_24634);
nand U24794 (N_24794,N_24579,N_24517);
or U24795 (N_24795,N_24574,N_24522);
nor U24796 (N_24796,N_24662,N_24749);
nor U24797 (N_24797,N_24620,N_24702);
nor U24798 (N_24798,N_24705,N_24652);
nand U24799 (N_24799,N_24650,N_24554);
nand U24800 (N_24800,N_24561,N_24562);
nor U24801 (N_24801,N_24619,N_24665);
and U24802 (N_24802,N_24713,N_24536);
or U24803 (N_24803,N_24515,N_24605);
or U24804 (N_24804,N_24610,N_24621);
nor U24805 (N_24805,N_24673,N_24596);
or U24806 (N_24806,N_24584,N_24663);
nand U24807 (N_24807,N_24691,N_24695);
and U24808 (N_24808,N_24523,N_24699);
nand U24809 (N_24809,N_24693,N_24723);
nor U24810 (N_24810,N_24547,N_24692);
and U24811 (N_24811,N_24647,N_24565);
and U24812 (N_24812,N_24566,N_24519);
and U24813 (N_24813,N_24521,N_24611);
nor U24814 (N_24814,N_24528,N_24701);
nand U24815 (N_24815,N_24602,N_24670);
nand U24816 (N_24816,N_24697,N_24601);
nand U24817 (N_24817,N_24666,N_24722);
and U24818 (N_24818,N_24671,N_24684);
xor U24819 (N_24819,N_24718,N_24726);
nor U24820 (N_24820,N_24609,N_24681);
nand U24821 (N_24821,N_24614,N_24592);
or U24822 (N_24822,N_24506,N_24563);
and U24823 (N_24823,N_24543,N_24643);
nor U24824 (N_24824,N_24559,N_24518);
nand U24825 (N_24825,N_24651,N_24530);
or U24826 (N_24826,N_24572,N_24594);
nor U24827 (N_24827,N_24688,N_24744);
nand U24828 (N_24828,N_24586,N_24512);
and U24829 (N_24829,N_24622,N_24520);
or U24830 (N_24830,N_24628,N_24555);
and U24831 (N_24831,N_24747,N_24678);
nand U24832 (N_24832,N_24548,N_24616);
or U24833 (N_24833,N_24655,N_24728);
nor U24834 (N_24834,N_24511,N_24646);
nor U24835 (N_24835,N_24735,N_24649);
and U24836 (N_24836,N_24558,N_24738);
nand U24837 (N_24837,N_24576,N_24516);
nand U24838 (N_24838,N_24734,N_24741);
nand U24839 (N_24839,N_24707,N_24546);
or U24840 (N_24840,N_24731,N_24617);
nor U24841 (N_24841,N_24660,N_24577);
or U24842 (N_24842,N_24658,N_24685);
or U24843 (N_24843,N_24510,N_24687);
nand U24844 (N_24844,N_24720,N_24508);
xnor U24845 (N_24845,N_24641,N_24739);
nor U24846 (N_24846,N_24721,N_24568);
nor U24847 (N_24847,N_24639,N_24637);
nand U24848 (N_24848,N_24674,N_24589);
and U24849 (N_24849,N_24745,N_24573);
nand U24850 (N_24850,N_24571,N_24742);
and U24851 (N_24851,N_24748,N_24711);
nor U24852 (N_24852,N_24680,N_24683);
and U24853 (N_24853,N_24612,N_24633);
and U24854 (N_24854,N_24676,N_24656);
or U24855 (N_24855,N_24541,N_24507);
nand U24856 (N_24856,N_24615,N_24710);
nor U24857 (N_24857,N_24567,N_24679);
or U24858 (N_24858,N_24533,N_24746);
nand U24859 (N_24859,N_24677,N_24535);
and U24860 (N_24860,N_24737,N_24509);
nand U24861 (N_24861,N_24553,N_24501);
and U24862 (N_24862,N_24694,N_24645);
nor U24863 (N_24863,N_24625,N_24725);
or U24864 (N_24864,N_24606,N_24599);
nor U24865 (N_24865,N_24724,N_24570);
or U24866 (N_24866,N_24648,N_24657);
nor U24867 (N_24867,N_24690,N_24569);
nor U24868 (N_24868,N_24661,N_24505);
or U24869 (N_24869,N_24640,N_24716);
xor U24870 (N_24870,N_24653,N_24595);
and U24871 (N_24871,N_24632,N_24591);
and U24872 (N_24872,N_24583,N_24527);
and U24873 (N_24873,N_24629,N_24500);
nor U24874 (N_24874,N_24714,N_24526);
and U24875 (N_24875,N_24585,N_24587);
nand U24876 (N_24876,N_24647,N_24557);
nand U24877 (N_24877,N_24571,N_24516);
nor U24878 (N_24878,N_24722,N_24571);
nand U24879 (N_24879,N_24640,N_24530);
nand U24880 (N_24880,N_24604,N_24543);
nor U24881 (N_24881,N_24645,N_24635);
or U24882 (N_24882,N_24585,N_24649);
or U24883 (N_24883,N_24618,N_24598);
nand U24884 (N_24884,N_24657,N_24609);
and U24885 (N_24885,N_24621,N_24624);
nand U24886 (N_24886,N_24701,N_24736);
nand U24887 (N_24887,N_24723,N_24549);
and U24888 (N_24888,N_24602,N_24611);
or U24889 (N_24889,N_24744,N_24602);
nand U24890 (N_24890,N_24504,N_24717);
nand U24891 (N_24891,N_24704,N_24571);
xnor U24892 (N_24892,N_24632,N_24561);
or U24893 (N_24893,N_24647,N_24507);
and U24894 (N_24894,N_24713,N_24690);
nand U24895 (N_24895,N_24523,N_24529);
and U24896 (N_24896,N_24726,N_24529);
or U24897 (N_24897,N_24535,N_24646);
nor U24898 (N_24898,N_24594,N_24558);
nand U24899 (N_24899,N_24735,N_24528);
or U24900 (N_24900,N_24623,N_24694);
xor U24901 (N_24901,N_24559,N_24706);
nand U24902 (N_24902,N_24723,N_24748);
and U24903 (N_24903,N_24666,N_24613);
xnor U24904 (N_24904,N_24610,N_24743);
nor U24905 (N_24905,N_24727,N_24551);
nor U24906 (N_24906,N_24557,N_24566);
or U24907 (N_24907,N_24633,N_24707);
nor U24908 (N_24908,N_24601,N_24558);
or U24909 (N_24909,N_24537,N_24545);
nand U24910 (N_24910,N_24647,N_24736);
or U24911 (N_24911,N_24540,N_24579);
nand U24912 (N_24912,N_24596,N_24651);
or U24913 (N_24913,N_24659,N_24504);
nor U24914 (N_24914,N_24584,N_24637);
nand U24915 (N_24915,N_24679,N_24682);
nor U24916 (N_24916,N_24640,N_24634);
nor U24917 (N_24917,N_24546,N_24714);
xnor U24918 (N_24918,N_24599,N_24557);
nor U24919 (N_24919,N_24571,N_24565);
nor U24920 (N_24920,N_24617,N_24583);
and U24921 (N_24921,N_24610,N_24501);
xnor U24922 (N_24922,N_24567,N_24569);
and U24923 (N_24923,N_24507,N_24699);
and U24924 (N_24924,N_24683,N_24699);
nor U24925 (N_24925,N_24747,N_24643);
or U24926 (N_24926,N_24576,N_24537);
and U24927 (N_24927,N_24729,N_24737);
or U24928 (N_24928,N_24549,N_24526);
and U24929 (N_24929,N_24681,N_24724);
and U24930 (N_24930,N_24635,N_24656);
and U24931 (N_24931,N_24507,N_24534);
nor U24932 (N_24932,N_24580,N_24585);
nand U24933 (N_24933,N_24572,N_24714);
and U24934 (N_24934,N_24709,N_24744);
or U24935 (N_24935,N_24533,N_24519);
nor U24936 (N_24936,N_24658,N_24672);
or U24937 (N_24937,N_24566,N_24562);
or U24938 (N_24938,N_24507,N_24674);
and U24939 (N_24939,N_24602,N_24604);
nand U24940 (N_24940,N_24703,N_24577);
nor U24941 (N_24941,N_24648,N_24525);
nor U24942 (N_24942,N_24605,N_24662);
nor U24943 (N_24943,N_24732,N_24544);
and U24944 (N_24944,N_24700,N_24546);
nor U24945 (N_24945,N_24663,N_24696);
nor U24946 (N_24946,N_24637,N_24504);
or U24947 (N_24947,N_24544,N_24627);
and U24948 (N_24948,N_24721,N_24563);
and U24949 (N_24949,N_24618,N_24590);
and U24950 (N_24950,N_24727,N_24510);
nand U24951 (N_24951,N_24512,N_24557);
nand U24952 (N_24952,N_24515,N_24544);
and U24953 (N_24953,N_24687,N_24566);
xor U24954 (N_24954,N_24626,N_24656);
and U24955 (N_24955,N_24652,N_24620);
nor U24956 (N_24956,N_24674,N_24590);
or U24957 (N_24957,N_24597,N_24620);
or U24958 (N_24958,N_24685,N_24561);
nand U24959 (N_24959,N_24592,N_24580);
and U24960 (N_24960,N_24545,N_24649);
nand U24961 (N_24961,N_24566,N_24505);
or U24962 (N_24962,N_24576,N_24731);
nor U24963 (N_24963,N_24588,N_24731);
and U24964 (N_24964,N_24580,N_24596);
and U24965 (N_24965,N_24694,N_24615);
nor U24966 (N_24966,N_24598,N_24626);
and U24967 (N_24967,N_24551,N_24745);
or U24968 (N_24968,N_24505,N_24620);
and U24969 (N_24969,N_24562,N_24588);
nand U24970 (N_24970,N_24638,N_24746);
nand U24971 (N_24971,N_24707,N_24593);
nand U24972 (N_24972,N_24625,N_24592);
and U24973 (N_24973,N_24608,N_24718);
and U24974 (N_24974,N_24646,N_24649);
and U24975 (N_24975,N_24670,N_24509);
nor U24976 (N_24976,N_24737,N_24646);
nor U24977 (N_24977,N_24538,N_24642);
nor U24978 (N_24978,N_24747,N_24625);
or U24979 (N_24979,N_24659,N_24505);
nor U24980 (N_24980,N_24629,N_24564);
nand U24981 (N_24981,N_24547,N_24512);
nand U24982 (N_24982,N_24589,N_24548);
nand U24983 (N_24983,N_24507,N_24598);
or U24984 (N_24984,N_24698,N_24593);
nand U24985 (N_24985,N_24738,N_24618);
nand U24986 (N_24986,N_24619,N_24650);
nor U24987 (N_24987,N_24567,N_24723);
nor U24988 (N_24988,N_24737,N_24684);
and U24989 (N_24989,N_24729,N_24681);
or U24990 (N_24990,N_24723,N_24515);
nand U24991 (N_24991,N_24528,N_24527);
nor U24992 (N_24992,N_24657,N_24747);
nor U24993 (N_24993,N_24730,N_24591);
and U24994 (N_24994,N_24620,N_24551);
nand U24995 (N_24995,N_24666,N_24703);
and U24996 (N_24996,N_24566,N_24713);
and U24997 (N_24997,N_24616,N_24529);
and U24998 (N_24998,N_24696,N_24568);
and U24999 (N_24999,N_24690,N_24623);
and UO_0 (O_0,N_24918,N_24852);
nand UO_1 (O_1,N_24983,N_24760);
or UO_2 (O_2,N_24772,N_24759);
or UO_3 (O_3,N_24997,N_24825);
nor UO_4 (O_4,N_24890,N_24930);
and UO_5 (O_5,N_24803,N_24783);
nand UO_6 (O_6,N_24875,N_24885);
and UO_7 (O_7,N_24887,N_24870);
nor UO_8 (O_8,N_24769,N_24859);
nor UO_9 (O_9,N_24917,N_24854);
nor UO_10 (O_10,N_24750,N_24906);
and UO_11 (O_11,N_24795,N_24903);
and UO_12 (O_12,N_24861,N_24856);
and UO_13 (O_13,N_24857,N_24848);
or UO_14 (O_14,N_24784,N_24786);
or UO_15 (O_15,N_24810,N_24976);
or UO_16 (O_16,N_24884,N_24782);
or UO_17 (O_17,N_24805,N_24931);
nand UO_18 (O_18,N_24863,N_24763);
and UO_19 (O_19,N_24921,N_24947);
nand UO_20 (O_20,N_24833,N_24912);
nor UO_21 (O_21,N_24876,N_24788);
or UO_22 (O_22,N_24847,N_24826);
nand UO_23 (O_23,N_24993,N_24896);
nor UO_24 (O_24,N_24928,N_24868);
nand UO_25 (O_25,N_24964,N_24967);
or UO_26 (O_26,N_24755,N_24820);
and UO_27 (O_27,N_24756,N_24821);
or UO_28 (O_28,N_24991,N_24837);
nand UO_29 (O_29,N_24956,N_24771);
nor UO_30 (O_30,N_24951,N_24839);
or UO_31 (O_31,N_24969,N_24984);
nand UO_32 (O_32,N_24879,N_24758);
and UO_33 (O_33,N_24781,N_24902);
nor UO_34 (O_34,N_24946,N_24933);
or UO_35 (O_35,N_24831,N_24836);
and UO_36 (O_36,N_24809,N_24910);
nor UO_37 (O_37,N_24777,N_24920);
nor UO_38 (O_38,N_24971,N_24923);
nand UO_39 (O_39,N_24874,N_24845);
or UO_40 (O_40,N_24934,N_24913);
or UO_41 (O_41,N_24904,N_24787);
nand UO_42 (O_42,N_24979,N_24855);
nand UO_43 (O_43,N_24998,N_24959);
nand UO_44 (O_44,N_24768,N_24916);
and UO_45 (O_45,N_24880,N_24774);
nor UO_46 (O_46,N_24754,N_24924);
nand UO_47 (O_47,N_24775,N_24966);
or UO_48 (O_48,N_24866,N_24909);
nor UO_49 (O_49,N_24864,N_24850);
or UO_50 (O_50,N_24941,N_24767);
or UO_51 (O_51,N_24865,N_24958);
or UO_52 (O_52,N_24927,N_24982);
and UO_53 (O_53,N_24962,N_24778);
and UO_54 (O_54,N_24765,N_24939);
and UO_55 (O_55,N_24994,N_24925);
and UO_56 (O_56,N_24897,N_24849);
or UO_57 (O_57,N_24869,N_24793);
or UO_58 (O_58,N_24840,N_24844);
nor UO_59 (O_59,N_24828,N_24996);
or UO_60 (O_60,N_24862,N_24761);
nand UO_61 (O_61,N_24842,N_24886);
and UO_62 (O_62,N_24851,N_24968);
and UO_63 (O_63,N_24999,N_24888);
and UO_64 (O_64,N_24955,N_24992);
xnor UO_65 (O_65,N_24948,N_24780);
nor UO_66 (O_66,N_24832,N_24792);
and UO_67 (O_67,N_24822,N_24881);
or UO_68 (O_68,N_24882,N_24853);
nor UO_69 (O_69,N_24977,N_24988);
nand UO_70 (O_70,N_24799,N_24929);
nor UO_71 (O_71,N_24892,N_24935);
or UO_72 (O_72,N_24807,N_24800);
or UO_73 (O_73,N_24814,N_24762);
nand UO_74 (O_74,N_24938,N_24907);
and UO_75 (O_75,N_24751,N_24773);
and UO_76 (O_76,N_24798,N_24891);
nand UO_77 (O_77,N_24950,N_24752);
and UO_78 (O_78,N_24899,N_24936);
nand UO_79 (O_79,N_24858,N_24894);
and UO_80 (O_80,N_24794,N_24804);
nand UO_81 (O_81,N_24974,N_24843);
or UO_82 (O_82,N_24957,N_24835);
nand UO_83 (O_83,N_24813,N_24900);
nor UO_84 (O_84,N_24915,N_24883);
xnor UO_85 (O_85,N_24944,N_24841);
and UO_86 (O_86,N_24908,N_24978);
nand UO_87 (O_87,N_24970,N_24986);
nand UO_88 (O_88,N_24953,N_24770);
and UO_89 (O_89,N_24785,N_24827);
nand UO_90 (O_90,N_24764,N_24817);
nand UO_91 (O_91,N_24872,N_24878);
nand UO_92 (O_92,N_24797,N_24949);
and UO_93 (O_93,N_24753,N_24816);
and UO_94 (O_94,N_24806,N_24942);
and UO_95 (O_95,N_24838,N_24873);
nor UO_96 (O_96,N_24802,N_24819);
and UO_97 (O_97,N_24973,N_24954);
nor UO_98 (O_98,N_24779,N_24945);
nand UO_99 (O_99,N_24889,N_24943);
nor UO_100 (O_100,N_24960,N_24877);
nand UO_101 (O_101,N_24989,N_24975);
or UO_102 (O_102,N_24815,N_24829);
or UO_103 (O_103,N_24985,N_24789);
and UO_104 (O_104,N_24914,N_24811);
or UO_105 (O_105,N_24871,N_24757);
nand UO_106 (O_106,N_24823,N_24846);
nor UO_107 (O_107,N_24972,N_24965);
or UO_108 (O_108,N_24952,N_24801);
nand UO_109 (O_109,N_24860,N_24961);
nor UO_110 (O_110,N_24919,N_24766);
or UO_111 (O_111,N_24867,N_24834);
and UO_112 (O_112,N_24791,N_24893);
nor UO_113 (O_113,N_24790,N_24812);
or UO_114 (O_114,N_24990,N_24922);
nand UO_115 (O_115,N_24830,N_24937);
and UO_116 (O_116,N_24995,N_24898);
nand UO_117 (O_117,N_24926,N_24905);
and UO_118 (O_118,N_24963,N_24940);
nor UO_119 (O_119,N_24980,N_24818);
and UO_120 (O_120,N_24981,N_24808);
nand UO_121 (O_121,N_24776,N_24895);
nand UO_122 (O_122,N_24987,N_24824);
nor UO_123 (O_123,N_24932,N_24796);
and UO_124 (O_124,N_24901,N_24911);
or UO_125 (O_125,N_24766,N_24900);
nor UO_126 (O_126,N_24858,N_24873);
nand UO_127 (O_127,N_24816,N_24860);
or UO_128 (O_128,N_24885,N_24999);
nor UO_129 (O_129,N_24943,N_24811);
nand UO_130 (O_130,N_24896,N_24903);
and UO_131 (O_131,N_24855,N_24753);
and UO_132 (O_132,N_24960,N_24857);
or UO_133 (O_133,N_24823,N_24880);
or UO_134 (O_134,N_24823,N_24803);
nor UO_135 (O_135,N_24793,N_24938);
and UO_136 (O_136,N_24989,N_24764);
nor UO_137 (O_137,N_24895,N_24881);
nor UO_138 (O_138,N_24972,N_24877);
or UO_139 (O_139,N_24900,N_24753);
nand UO_140 (O_140,N_24769,N_24864);
or UO_141 (O_141,N_24751,N_24767);
or UO_142 (O_142,N_24938,N_24919);
or UO_143 (O_143,N_24847,N_24898);
nor UO_144 (O_144,N_24966,N_24871);
nand UO_145 (O_145,N_24999,N_24891);
nand UO_146 (O_146,N_24855,N_24938);
nor UO_147 (O_147,N_24768,N_24854);
and UO_148 (O_148,N_24900,N_24855);
nor UO_149 (O_149,N_24991,N_24858);
nand UO_150 (O_150,N_24977,N_24779);
nor UO_151 (O_151,N_24969,N_24762);
nor UO_152 (O_152,N_24820,N_24885);
and UO_153 (O_153,N_24935,N_24757);
and UO_154 (O_154,N_24924,N_24843);
nor UO_155 (O_155,N_24787,N_24968);
nand UO_156 (O_156,N_24980,N_24991);
nand UO_157 (O_157,N_24829,N_24800);
and UO_158 (O_158,N_24875,N_24887);
and UO_159 (O_159,N_24911,N_24863);
nand UO_160 (O_160,N_24849,N_24887);
nand UO_161 (O_161,N_24900,N_24974);
and UO_162 (O_162,N_24751,N_24792);
nor UO_163 (O_163,N_24971,N_24769);
or UO_164 (O_164,N_24996,N_24988);
or UO_165 (O_165,N_24987,N_24882);
nand UO_166 (O_166,N_24785,N_24949);
nor UO_167 (O_167,N_24916,N_24817);
nand UO_168 (O_168,N_24964,N_24955);
nor UO_169 (O_169,N_24911,N_24970);
nor UO_170 (O_170,N_24907,N_24860);
nor UO_171 (O_171,N_24962,N_24851);
nor UO_172 (O_172,N_24999,N_24975);
nor UO_173 (O_173,N_24819,N_24932);
and UO_174 (O_174,N_24951,N_24958);
nor UO_175 (O_175,N_24881,N_24951);
and UO_176 (O_176,N_24772,N_24934);
or UO_177 (O_177,N_24786,N_24973);
nor UO_178 (O_178,N_24763,N_24892);
nand UO_179 (O_179,N_24856,N_24940);
nand UO_180 (O_180,N_24960,N_24829);
nand UO_181 (O_181,N_24864,N_24949);
nor UO_182 (O_182,N_24801,N_24881);
and UO_183 (O_183,N_24750,N_24958);
or UO_184 (O_184,N_24857,N_24751);
and UO_185 (O_185,N_24900,N_24910);
and UO_186 (O_186,N_24890,N_24957);
nor UO_187 (O_187,N_24875,N_24994);
nor UO_188 (O_188,N_24872,N_24917);
nand UO_189 (O_189,N_24843,N_24884);
or UO_190 (O_190,N_24803,N_24955);
or UO_191 (O_191,N_24804,N_24974);
nand UO_192 (O_192,N_24900,N_24809);
and UO_193 (O_193,N_24782,N_24936);
and UO_194 (O_194,N_24790,N_24847);
nand UO_195 (O_195,N_24879,N_24955);
nand UO_196 (O_196,N_24779,N_24967);
nor UO_197 (O_197,N_24996,N_24939);
nand UO_198 (O_198,N_24844,N_24972);
nand UO_199 (O_199,N_24849,N_24856);
and UO_200 (O_200,N_24828,N_24858);
or UO_201 (O_201,N_24914,N_24886);
or UO_202 (O_202,N_24937,N_24969);
nor UO_203 (O_203,N_24882,N_24886);
or UO_204 (O_204,N_24843,N_24815);
nand UO_205 (O_205,N_24930,N_24794);
nor UO_206 (O_206,N_24993,N_24891);
nand UO_207 (O_207,N_24866,N_24872);
or UO_208 (O_208,N_24801,N_24804);
nand UO_209 (O_209,N_24858,N_24882);
and UO_210 (O_210,N_24899,N_24839);
nand UO_211 (O_211,N_24751,N_24761);
or UO_212 (O_212,N_24892,N_24799);
nand UO_213 (O_213,N_24851,N_24958);
and UO_214 (O_214,N_24876,N_24750);
or UO_215 (O_215,N_24835,N_24869);
and UO_216 (O_216,N_24938,N_24828);
nand UO_217 (O_217,N_24851,N_24765);
and UO_218 (O_218,N_24907,N_24843);
nor UO_219 (O_219,N_24865,N_24892);
or UO_220 (O_220,N_24963,N_24966);
and UO_221 (O_221,N_24949,N_24771);
and UO_222 (O_222,N_24825,N_24867);
nand UO_223 (O_223,N_24952,N_24838);
nand UO_224 (O_224,N_24751,N_24903);
or UO_225 (O_225,N_24803,N_24940);
and UO_226 (O_226,N_24771,N_24765);
nor UO_227 (O_227,N_24991,N_24974);
xor UO_228 (O_228,N_24772,N_24971);
nand UO_229 (O_229,N_24979,N_24904);
nand UO_230 (O_230,N_24945,N_24772);
or UO_231 (O_231,N_24999,N_24991);
nand UO_232 (O_232,N_24889,N_24873);
nand UO_233 (O_233,N_24785,N_24757);
nand UO_234 (O_234,N_24797,N_24828);
and UO_235 (O_235,N_24983,N_24859);
and UO_236 (O_236,N_24907,N_24767);
nor UO_237 (O_237,N_24771,N_24933);
and UO_238 (O_238,N_24815,N_24784);
and UO_239 (O_239,N_24808,N_24906);
or UO_240 (O_240,N_24956,N_24777);
nand UO_241 (O_241,N_24865,N_24978);
nand UO_242 (O_242,N_24973,N_24869);
and UO_243 (O_243,N_24868,N_24846);
or UO_244 (O_244,N_24923,N_24777);
nand UO_245 (O_245,N_24944,N_24902);
and UO_246 (O_246,N_24783,N_24811);
nand UO_247 (O_247,N_24963,N_24895);
nor UO_248 (O_248,N_24934,N_24895);
or UO_249 (O_249,N_24777,N_24928);
nand UO_250 (O_250,N_24821,N_24970);
xor UO_251 (O_251,N_24891,N_24915);
and UO_252 (O_252,N_24977,N_24924);
nand UO_253 (O_253,N_24959,N_24900);
or UO_254 (O_254,N_24817,N_24863);
or UO_255 (O_255,N_24796,N_24948);
nor UO_256 (O_256,N_24936,N_24857);
and UO_257 (O_257,N_24811,N_24969);
and UO_258 (O_258,N_24941,N_24884);
or UO_259 (O_259,N_24886,N_24757);
or UO_260 (O_260,N_24959,N_24939);
nand UO_261 (O_261,N_24847,N_24837);
nor UO_262 (O_262,N_24865,N_24893);
nand UO_263 (O_263,N_24922,N_24778);
or UO_264 (O_264,N_24936,N_24795);
or UO_265 (O_265,N_24815,N_24789);
nor UO_266 (O_266,N_24958,N_24880);
or UO_267 (O_267,N_24793,N_24858);
nor UO_268 (O_268,N_24877,N_24908);
and UO_269 (O_269,N_24806,N_24811);
or UO_270 (O_270,N_24901,N_24837);
and UO_271 (O_271,N_24773,N_24888);
nand UO_272 (O_272,N_24858,N_24940);
or UO_273 (O_273,N_24997,N_24871);
or UO_274 (O_274,N_24985,N_24758);
nand UO_275 (O_275,N_24974,N_24751);
nor UO_276 (O_276,N_24943,N_24924);
or UO_277 (O_277,N_24891,N_24859);
nand UO_278 (O_278,N_24775,N_24827);
nor UO_279 (O_279,N_24907,N_24958);
or UO_280 (O_280,N_24829,N_24888);
or UO_281 (O_281,N_24750,N_24798);
nor UO_282 (O_282,N_24935,N_24954);
or UO_283 (O_283,N_24801,N_24904);
nor UO_284 (O_284,N_24928,N_24885);
nor UO_285 (O_285,N_24960,N_24818);
and UO_286 (O_286,N_24992,N_24813);
and UO_287 (O_287,N_24852,N_24945);
nor UO_288 (O_288,N_24920,N_24781);
and UO_289 (O_289,N_24920,N_24769);
nor UO_290 (O_290,N_24912,N_24952);
and UO_291 (O_291,N_24773,N_24850);
nand UO_292 (O_292,N_24855,N_24880);
and UO_293 (O_293,N_24978,N_24895);
or UO_294 (O_294,N_24878,N_24913);
and UO_295 (O_295,N_24906,N_24925);
nor UO_296 (O_296,N_24954,N_24887);
nand UO_297 (O_297,N_24903,N_24799);
or UO_298 (O_298,N_24812,N_24896);
nor UO_299 (O_299,N_24978,N_24993);
nand UO_300 (O_300,N_24878,N_24870);
or UO_301 (O_301,N_24788,N_24820);
and UO_302 (O_302,N_24874,N_24809);
nor UO_303 (O_303,N_24840,N_24936);
or UO_304 (O_304,N_24952,N_24984);
and UO_305 (O_305,N_24989,N_24941);
or UO_306 (O_306,N_24842,N_24780);
and UO_307 (O_307,N_24981,N_24829);
nor UO_308 (O_308,N_24808,N_24869);
nor UO_309 (O_309,N_24876,N_24977);
nand UO_310 (O_310,N_24836,N_24764);
or UO_311 (O_311,N_24827,N_24855);
or UO_312 (O_312,N_24790,N_24907);
or UO_313 (O_313,N_24829,N_24808);
or UO_314 (O_314,N_24794,N_24840);
and UO_315 (O_315,N_24835,N_24829);
nand UO_316 (O_316,N_24924,N_24898);
and UO_317 (O_317,N_24797,N_24961);
nor UO_318 (O_318,N_24816,N_24988);
nor UO_319 (O_319,N_24896,N_24830);
and UO_320 (O_320,N_24794,N_24830);
nand UO_321 (O_321,N_24759,N_24983);
or UO_322 (O_322,N_24946,N_24907);
xnor UO_323 (O_323,N_24879,N_24990);
and UO_324 (O_324,N_24975,N_24982);
nand UO_325 (O_325,N_24867,N_24934);
and UO_326 (O_326,N_24998,N_24948);
or UO_327 (O_327,N_24886,N_24798);
and UO_328 (O_328,N_24798,N_24795);
and UO_329 (O_329,N_24804,N_24904);
and UO_330 (O_330,N_24900,N_24759);
nor UO_331 (O_331,N_24788,N_24839);
or UO_332 (O_332,N_24817,N_24940);
or UO_333 (O_333,N_24821,N_24814);
nor UO_334 (O_334,N_24918,N_24913);
and UO_335 (O_335,N_24752,N_24802);
and UO_336 (O_336,N_24759,N_24897);
and UO_337 (O_337,N_24768,N_24998);
nand UO_338 (O_338,N_24803,N_24969);
or UO_339 (O_339,N_24978,N_24853);
nand UO_340 (O_340,N_24750,N_24779);
nor UO_341 (O_341,N_24865,N_24840);
nor UO_342 (O_342,N_24824,N_24755);
nor UO_343 (O_343,N_24955,N_24965);
nor UO_344 (O_344,N_24939,N_24775);
nor UO_345 (O_345,N_24970,N_24953);
or UO_346 (O_346,N_24798,N_24864);
nor UO_347 (O_347,N_24944,N_24766);
and UO_348 (O_348,N_24827,N_24824);
nand UO_349 (O_349,N_24855,N_24906);
and UO_350 (O_350,N_24874,N_24977);
and UO_351 (O_351,N_24901,N_24821);
nor UO_352 (O_352,N_24834,N_24849);
nor UO_353 (O_353,N_24837,N_24914);
and UO_354 (O_354,N_24837,N_24908);
nand UO_355 (O_355,N_24976,N_24894);
and UO_356 (O_356,N_24900,N_24784);
and UO_357 (O_357,N_24792,N_24919);
and UO_358 (O_358,N_24853,N_24810);
nor UO_359 (O_359,N_24923,N_24858);
or UO_360 (O_360,N_24805,N_24795);
nor UO_361 (O_361,N_24964,N_24809);
nor UO_362 (O_362,N_24871,N_24783);
nand UO_363 (O_363,N_24830,N_24915);
and UO_364 (O_364,N_24771,N_24857);
or UO_365 (O_365,N_24784,N_24874);
nand UO_366 (O_366,N_24987,N_24763);
nand UO_367 (O_367,N_24966,N_24774);
nand UO_368 (O_368,N_24769,N_24816);
nand UO_369 (O_369,N_24760,N_24832);
nor UO_370 (O_370,N_24778,N_24824);
nor UO_371 (O_371,N_24914,N_24763);
or UO_372 (O_372,N_24825,N_24849);
or UO_373 (O_373,N_24967,N_24765);
nor UO_374 (O_374,N_24958,N_24998);
xor UO_375 (O_375,N_24927,N_24816);
or UO_376 (O_376,N_24889,N_24907);
nor UO_377 (O_377,N_24933,N_24940);
nor UO_378 (O_378,N_24769,N_24918);
nand UO_379 (O_379,N_24922,N_24776);
nand UO_380 (O_380,N_24833,N_24808);
nand UO_381 (O_381,N_24937,N_24941);
or UO_382 (O_382,N_24984,N_24979);
xnor UO_383 (O_383,N_24863,N_24862);
and UO_384 (O_384,N_24985,N_24977);
nor UO_385 (O_385,N_24792,N_24999);
or UO_386 (O_386,N_24908,N_24881);
nor UO_387 (O_387,N_24831,N_24955);
nand UO_388 (O_388,N_24874,N_24783);
nor UO_389 (O_389,N_24973,N_24843);
and UO_390 (O_390,N_24960,N_24840);
and UO_391 (O_391,N_24982,N_24771);
nand UO_392 (O_392,N_24882,N_24915);
or UO_393 (O_393,N_24784,N_24881);
nor UO_394 (O_394,N_24915,N_24970);
and UO_395 (O_395,N_24869,N_24768);
or UO_396 (O_396,N_24835,N_24986);
and UO_397 (O_397,N_24778,N_24954);
or UO_398 (O_398,N_24906,N_24827);
nor UO_399 (O_399,N_24765,N_24900);
nand UO_400 (O_400,N_24904,N_24921);
nor UO_401 (O_401,N_24849,N_24799);
and UO_402 (O_402,N_24952,N_24812);
and UO_403 (O_403,N_24976,N_24783);
or UO_404 (O_404,N_24828,N_24982);
or UO_405 (O_405,N_24899,N_24807);
nor UO_406 (O_406,N_24849,N_24989);
or UO_407 (O_407,N_24830,N_24873);
and UO_408 (O_408,N_24949,N_24987);
and UO_409 (O_409,N_24997,N_24783);
and UO_410 (O_410,N_24909,N_24851);
and UO_411 (O_411,N_24847,N_24992);
nor UO_412 (O_412,N_24873,N_24992);
xor UO_413 (O_413,N_24847,N_24983);
nor UO_414 (O_414,N_24852,N_24815);
and UO_415 (O_415,N_24883,N_24953);
and UO_416 (O_416,N_24871,N_24822);
or UO_417 (O_417,N_24907,N_24984);
nand UO_418 (O_418,N_24770,N_24948);
nor UO_419 (O_419,N_24789,N_24791);
or UO_420 (O_420,N_24811,N_24814);
or UO_421 (O_421,N_24942,N_24771);
nor UO_422 (O_422,N_24815,N_24828);
xnor UO_423 (O_423,N_24799,N_24820);
and UO_424 (O_424,N_24803,N_24768);
nor UO_425 (O_425,N_24766,N_24818);
or UO_426 (O_426,N_24765,N_24872);
and UO_427 (O_427,N_24779,N_24974);
nor UO_428 (O_428,N_24823,N_24965);
and UO_429 (O_429,N_24885,N_24810);
or UO_430 (O_430,N_24770,N_24939);
nand UO_431 (O_431,N_24871,N_24933);
nor UO_432 (O_432,N_24992,N_24891);
or UO_433 (O_433,N_24773,N_24780);
nand UO_434 (O_434,N_24788,N_24949);
and UO_435 (O_435,N_24973,N_24761);
nand UO_436 (O_436,N_24965,N_24826);
nor UO_437 (O_437,N_24942,N_24820);
or UO_438 (O_438,N_24823,N_24887);
and UO_439 (O_439,N_24980,N_24939);
and UO_440 (O_440,N_24987,N_24753);
nor UO_441 (O_441,N_24797,N_24996);
nand UO_442 (O_442,N_24879,N_24766);
or UO_443 (O_443,N_24924,N_24923);
and UO_444 (O_444,N_24935,N_24870);
nor UO_445 (O_445,N_24847,N_24772);
nand UO_446 (O_446,N_24941,N_24902);
and UO_447 (O_447,N_24768,N_24908);
nand UO_448 (O_448,N_24833,N_24986);
and UO_449 (O_449,N_24965,N_24979);
and UO_450 (O_450,N_24965,N_24771);
or UO_451 (O_451,N_24832,N_24935);
or UO_452 (O_452,N_24796,N_24833);
and UO_453 (O_453,N_24974,N_24830);
or UO_454 (O_454,N_24902,N_24810);
and UO_455 (O_455,N_24765,N_24793);
or UO_456 (O_456,N_24911,N_24938);
nor UO_457 (O_457,N_24970,N_24958);
nor UO_458 (O_458,N_24883,N_24762);
nor UO_459 (O_459,N_24799,N_24990);
nand UO_460 (O_460,N_24839,N_24953);
nand UO_461 (O_461,N_24933,N_24961);
and UO_462 (O_462,N_24896,N_24818);
nor UO_463 (O_463,N_24810,N_24940);
or UO_464 (O_464,N_24843,N_24830);
xor UO_465 (O_465,N_24922,N_24840);
nor UO_466 (O_466,N_24869,N_24972);
nand UO_467 (O_467,N_24823,N_24872);
nand UO_468 (O_468,N_24917,N_24853);
nand UO_469 (O_469,N_24986,N_24947);
or UO_470 (O_470,N_24968,N_24806);
xor UO_471 (O_471,N_24847,N_24884);
and UO_472 (O_472,N_24953,N_24907);
nor UO_473 (O_473,N_24874,N_24776);
and UO_474 (O_474,N_24794,N_24940);
and UO_475 (O_475,N_24774,N_24861);
nand UO_476 (O_476,N_24951,N_24869);
nand UO_477 (O_477,N_24901,N_24985);
or UO_478 (O_478,N_24848,N_24976);
and UO_479 (O_479,N_24896,N_24990);
or UO_480 (O_480,N_24951,N_24791);
and UO_481 (O_481,N_24832,N_24874);
nor UO_482 (O_482,N_24852,N_24988);
and UO_483 (O_483,N_24775,N_24903);
or UO_484 (O_484,N_24792,N_24907);
nor UO_485 (O_485,N_24830,N_24763);
or UO_486 (O_486,N_24785,N_24765);
nor UO_487 (O_487,N_24989,N_24867);
nand UO_488 (O_488,N_24825,N_24752);
nand UO_489 (O_489,N_24823,N_24949);
and UO_490 (O_490,N_24834,N_24798);
nand UO_491 (O_491,N_24940,N_24772);
nor UO_492 (O_492,N_24826,N_24941);
and UO_493 (O_493,N_24833,N_24913);
nand UO_494 (O_494,N_24984,N_24862);
nor UO_495 (O_495,N_24902,N_24995);
or UO_496 (O_496,N_24793,N_24904);
nor UO_497 (O_497,N_24752,N_24828);
nand UO_498 (O_498,N_24755,N_24798);
or UO_499 (O_499,N_24823,N_24893);
or UO_500 (O_500,N_24844,N_24834);
or UO_501 (O_501,N_24803,N_24903);
and UO_502 (O_502,N_24937,N_24804);
or UO_503 (O_503,N_24886,N_24765);
nand UO_504 (O_504,N_24929,N_24775);
and UO_505 (O_505,N_24904,N_24757);
or UO_506 (O_506,N_24879,N_24936);
and UO_507 (O_507,N_24944,N_24818);
or UO_508 (O_508,N_24839,N_24757);
and UO_509 (O_509,N_24795,N_24775);
xor UO_510 (O_510,N_24787,N_24752);
nor UO_511 (O_511,N_24796,N_24935);
and UO_512 (O_512,N_24817,N_24829);
and UO_513 (O_513,N_24960,N_24967);
nor UO_514 (O_514,N_24827,N_24779);
nand UO_515 (O_515,N_24762,N_24811);
and UO_516 (O_516,N_24894,N_24837);
nand UO_517 (O_517,N_24834,N_24941);
nand UO_518 (O_518,N_24879,N_24960);
nand UO_519 (O_519,N_24922,N_24766);
or UO_520 (O_520,N_24757,N_24970);
or UO_521 (O_521,N_24797,N_24999);
and UO_522 (O_522,N_24856,N_24795);
nor UO_523 (O_523,N_24960,N_24802);
nor UO_524 (O_524,N_24874,N_24923);
nand UO_525 (O_525,N_24998,N_24861);
nor UO_526 (O_526,N_24856,N_24919);
nand UO_527 (O_527,N_24919,N_24964);
and UO_528 (O_528,N_24921,N_24945);
and UO_529 (O_529,N_24884,N_24772);
nor UO_530 (O_530,N_24889,N_24833);
nor UO_531 (O_531,N_24757,N_24975);
nand UO_532 (O_532,N_24927,N_24932);
or UO_533 (O_533,N_24895,N_24754);
nor UO_534 (O_534,N_24957,N_24761);
nand UO_535 (O_535,N_24766,N_24908);
or UO_536 (O_536,N_24800,N_24968);
nand UO_537 (O_537,N_24997,N_24852);
or UO_538 (O_538,N_24953,N_24898);
and UO_539 (O_539,N_24868,N_24995);
nor UO_540 (O_540,N_24914,N_24849);
or UO_541 (O_541,N_24997,N_24982);
nor UO_542 (O_542,N_24974,N_24858);
nand UO_543 (O_543,N_24843,N_24983);
or UO_544 (O_544,N_24944,N_24858);
nand UO_545 (O_545,N_24890,N_24904);
or UO_546 (O_546,N_24902,N_24853);
and UO_547 (O_547,N_24755,N_24924);
nor UO_548 (O_548,N_24912,N_24960);
nand UO_549 (O_549,N_24795,N_24905);
and UO_550 (O_550,N_24955,N_24793);
or UO_551 (O_551,N_24904,N_24846);
or UO_552 (O_552,N_24805,N_24878);
or UO_553 (O_553,N_24833,N_24863);
and UO_554 (O_554,N_24841,N_24978);
or UO_555 (O_555,N_24916,N_24753);
and UO_556 (O_556,N_24801,N_24778);
and UO_557 (O_557,N_24911,N_24881);
or UO_558 (O_558,N_24790,N_24958);
nand UO_559 (O_559,N_24890,N_24752);
nand UO_560 (O_560,N_24980,N_24843);
nand UO_561 (O_561,N_24952,N_24769);
or UO_562 (O_562,N_24962,N_24979);
nand UO_563 (O_563,N_24853,N_24875);
nand UO_564 (O_564,N_24848,N_24887);
and UO_565 (O_565,N_24908,N_24848);
nand UO_566 (O_566,N_24895,N_24924);
or UO_567 (O_567,N_24805,N_24989);
nand UO_568 (O_568,N_24856,N_24938);
nor UO_569 (O_569,N_24958,N_24954);
and UO_570 (O_570,N_24931,N_24905);
or UO_571 (O_571,N_24867,N_24927);
and UO_572 (O_572,N_24914,N_24956);
and UO_573 (O_573,N_24949,N_24940);
or UO_574 (O_574,N_24937,N_24791);
nand UO_575 (O_575,N_24874,N_24957);
and UO_576 (O_576,N_24794,N_24791);
or UO_577 (O_577,N_24823,N_24818);
or UO_578 (O_578,N_24792,N_24943);
nor UO_579 (O_579,N_24807,N_24818);
and UO_580 (O_580,N_24814,N_24906);
nor UO_581 (O_581,N_24862,N_24884);
and UO_582 (O_582,N_24950,N_24907);
nor UO_583 (O_583,N_24904,N_24880);
nor UO_584 (O_584,N_24902,N_24758);
or UO_585 (O_585,N_24806,N_24900);
or UO_586 (O_586,N_24844,N_24926);
and UO_587 (O_587,N_24819,N_24828);
or UO_588 (O_588,N_24771,N_24829);
nand UO_589 (O_589,N_24770,N_24970);
nor UO_590 (O_590,N_24794,N_24771);
and UO_591 (O_591,N_24784,N_24851);
or UO_592 (O_592,N_24869,N_24879);
or UO_593 (O_593,N_24835,N_24828);
nand UO_594 (O_594,N_24852,N_24881);
nand UO_595 (O_595,N_24950,N_24821);
nor UO_596 (O_596,N_24911,N_24940);
nand UO_597 (O_597,N_24837,N_24799);
nand UO_598 (O_598,N_24804,N_24771);
nand UO_599 (O_599,N_24999,N_24983);
nor UO_600 (O_600,N_24898,N_24883);
and UO_601 (O_601,N_24889,N_24818);
and UO_602 (O_602,N_24861,N_24947);
nand UO_603 (O_603,N_24976,N_24996);
or UO_604 (O_604,N_24787,N_24923);
or UO_605 (O_605,N_24966,N_24851);
nand UO_606 (O_606,N_24996,N_24863);
xnor UO_607 (O_607,N_24755,N_24807);
nor UO_608 (O_608,N_24754,N_24988);
nand UO_609 (O_609,N_24842,N_24914);
and UO_610 (O_610,N_24916,N_24773);
or UO_611 (O_611,N_24796,N_24933);
or UO_612 (O_612,N_24820,N_24981);
or UO_613 (O_613,N_24798,N_24822);
nor UO_614 (O_614,N_24793,N_24933);
nor UO_615 (O_615,N_24954,N_24761);
or UO_616 (O_616,N_24865,N_24798);
and UO_617 (O_617,N_24856,N_24928);
nor UO_618 (O_618,N_24984,N_24850);
and UO_619 (O_619,N_24956,N_24867);
nor UO_620 (O_620,N_24914,N_24786);
nand UO_621 (O_621,N_24884,N_24776);
or UO_622 (O_622,N_24845,N_24962);
nand UO_623 (O_623,N_24799,N_24930);
and UO_624 (O_624,N_24842,N_24990);
nor UO_625 (O_625,N_24987,N_24931);
and UO_626 (O_626,N_24808,N_24826);
nor UO_627 (O_627,N_24765,N_24820);
or UO_628 (O_628,N_24969,N_24781);
and UO_629 (O_629,N_24986,N_24781);
and UO_630 (O_630,N_24840,N_24898);
and UO_631 (O_631,N_24842,N_24844);
or UO_632 (O_632,N_24958,N_24971);
nor UO_633 (O_633,N_24767,N_24801);
xor UO_634 (O_634,N_24973,N_24916);
or UO_635 (O_635,N_24754,N_24792);
nand UO_636 (O_636,N_24841,N_24796);
or UO_637 (O_637,N_24931,N_24873);
and UO_638 (O_638,N_24841,N_24771);
nor UO_639 (O_639,N_24953,N_24798);
or UO_640 (O_640,N_24772,N_24781);
nor UO_641 (O_641,N_24944,N_24814);
and UO_642 (O_642,N_24947,N_24841);
or UO_643 (O_643,N_24959,N_24804);
and UO_644 (O_644,N_24843,N_24938);
and UO_645 (O_645,N_24975,N_24995);
nor UO_646 (O_646,N_24841,N_24787);
nor UO_647 (O_647,N_24957,N_24877);
or UO_648 (O_648,N_24865,N_24762);
nand UO_649 (O_649,N_24791,N_24897);
nor UO_650 (O_650,N_24860,N_24968);
nor UO_651 (O_651,N_24859,N_24883);
and UO_652 (O_652,N_24972,N_24806);
xor UO_653 (O_653,N_24753,N_24840);
nand UO_654 (O_654,N_24858,N_24877);
or UO_655 (O_655,N_24902,N_24901);
and UO_656 (O_656,N_24936,N_24760);
nor UO_657 (O_657,N_24940,N_24921);
or UO_658 (O_658,N_24966,N_24839);
nand UO_659 (O_659,N_24869,N_24983);
and UO_660 (O_660,N_24886,N_24766);
and UO_661 (O_661,N_24806,N_24931);
nand UO_662 (O_662,N_24904,N_24841);
nand UO_663 (O_663,N_24897,N_24845);
or UO_664 (O_664,N_24911,N_24861);
nand UO_665 (O_665,N_24766,N_24981);
and UO_666 (O_666,N_24859,N_24918);
nor UO_667 (O_667,N_24927,N_24975);
or UO_668 (O_668,N_24761,N_24968);
or UO_669 (O_669,N_24797,N_24947);
or UO_670 (O_670,N_24808,N_24949);
or UO_671 (O_671,N_24938,N_24751);
nand UO_672 (O_672,N_24844,N_24761);
or UO_673 (O_673,N_24929,N_24836);
and UO_674 (O_674,N_24929,N_24890);
or UO_675 (O_675,N_24915,N_24788);
and UO_676 (O_676,N_24951,N_24989);
nand UO_677 (O_677,N_24814,N_24842);
and UO_678 (O_678,N_24809,N_24946);
nor UO_679 (O_679,N_24802,N_24863);
and UO_680 (O_680,N_24816,N_24784);
or UO_681 (O_681,N_24925,N_24953);
or UO_682 (O_682,N_24893,N_24962);
and UO_683 (O_683,N_24893,N_24880);
and UO_684 (O_684,N_24765,N_24920);
nand UO_685 (O_685,N_24774,N_24849);
and UO_686 (O_686,N_24961,N_24846);
nor UO_687 (O_687,N_24997,N_24778);
nor UO_688 (O_688,N_24973,N_24941);
nor UO_689 (O_689,N_24905,N_24821);
and UO_690 (O_690,N_24922,N_24869);
nand UO_691 (O_691,N_24991,N_24853);
nand UO_692 (O_692,N_24869,N_24909);
and UO_693 (O_693,N_24897,N_24860);
nor UO_694 (O_694,N_24879,N_24863);
nand UO_695 (O_695,N_24958,N_24856);
nor UO_696 (O_696,N_24835,N_24961);
or UO_697 (O_697,N_24762,N_24758);
nor UO_698 (O_698,N_24759,N_24771);
nand UO_699 (O_699,N_24926,N_24895);
nand UO_700 (O_700,N_24807,N_24901);
nor UO_701 (O_701,N_24990,N_24871);
or UO_702 (O_702,N_24752,N_24788);
nor UO_703 (O_703,N_24971,N_24870);
and UO_704 (O_704,N_24864,N_24826);
nor UO_705 (O_705,N_24866,N_24751);
nor UO_706 (O_706,N_24969,N_24851);
or UO_707 (O_707,N_24818,N_24975);
nor UO_708 (O_708,N_24813,N_24847);
nand UO_709 (O_709,N_24988,N_24850);
and UO_710 (O_710,N_24862,N_24860);
and UO_711 (O_711,N_24948,N_24776);
nor UO_712 (O_712,N_24949,N_24762);
and UO_713 (O_713,N_24862,N_24875);
or UO_714 (O_714,N_24998,N_24855);
and UO_715 (O_715,N_24966,N_24902);
nand UO_716 (O_716,N_24943,N_24888);
nor UO_717 (O_717,N_24968,N_24886);
nor UO_718 (O_718,N_24854,N_24939);
nor UO_719 (O_719,N_24798,N_24959);
and UO_720 (O_720,N_24837,N_24993);
nor UO_721 (O_721,N_24868,N_24921);
nand UO_722 (O_722,N_24961,N_24885);
nor UO_723 (O_723,N_24828,N_24943);
nor UO_724 (O_724,N_24985,N_24893);
nand UO_725 (O_725,N_24768,N_24899);
nor UO_726 (O_726,N_24930,N_24956);
nand UO_727 (O_727,N_24909,N_24806);
and UO_728 (O_728,N_24872,N_24951);
nor UO_729 (O_729,N_24965,N_24929);
or UO_730 (O_730,N_24959,N_24805);
nand UO_731 (O_731,N_24924,N_24976);
nor UO_732 (O_732,N_24810,N_24982);
and UO_733 (O_733,N_24845,N_24923);
nor UO_734 (O_734,N_24769,N_24762);
and UO_735 (O_735,N_24874,N_24818);
nor UO_736 (O_736,N_24897,N_24865);
and UO_737 (O_737,N_24916,N_24955);
nand UO_738 (O_738,N_24926,N_24947);
nand UO_739 (O_739,N_24890,N_24999);
nor UO_740 (O_740,N_24885,N_24954);
nand UO_741 (O_741,N_24857,N_24961);
or UO_742 (O_742,N_24810,N_24825);
and UO_743 (O_743,N_24782,N_24772);
or UO_744 (O_744,N_24857,N_24879);
or UO_745 (O_745,N_24878,N_24967);
nor UO_746 (O_746,N_24890,N_24893);
or UO_747 (O_747,N_24809,N_24926);
nand UO_748 (O_748,N_24806,N_24861);
nor UO_749 (O_749,N_24780,N_24834);
and UO_750 (O_750,N_24823,N_24807);
and UO_751 (O_751,N_24877,N_24765);
and UO_752 (O_752,N_24854,N_24974);
or UO_753 (O_753,N_24804,N_24854);
or UO_754 (O_754,N_24980,N_24794);
nor UO_755 (O_755,N_24786,N_24840);
and UO_756 (O_756,N_24792,N_24942);
or UO_757 (O_757,N_24825,N_24850);
nor UO_758 (O_758,N_24757,N_24942);
nand UO_759 (O_759,N_24821,N_24947);
nor UO_760 (O_760,N_24872,N_24995);
nor UO_761 (O_761,N_24917,N_24989);
and UO_762 (O_762,N_24908,N_24898);
or UO_763 (O_763,N_24984,N_24908);
and UO_764 (O_764,N_24877,N_24851);
nand UO_765 (O_765,N_24835,N_24956);
nand UO_766 (O_766,N_24873,N_24952);
nor UO_767 (O_767,N_24921,N_24784);
nor UO_768 (O_768,N_24922,N_24802);
or UO_769 (O_769,N_24977,N_24775);
nand UO_770 (O_770,N_24814,N_24878);
nor UO_771 (O_771,N_24974,N_24820);
or UO_772 (O_772,N_24996,N_24814);
and UO_773 (O_773,N_24944,N_24982);
nand UO_774 (O_774,N_24752,N_24838);
and UO_775 (O_775,N_24982,N_24826);
nand UO_776 (O_776,N_24891,N_24767);
nor UO_777 (O_777,N_24837,N_24941);
or UO_778 (O_778,N_24942,N_24907);
or UO_779 (O_779,N_24807,N_24940);
or UO_780 (O_780,N_24988,N_24831);
and UO_781 (O_781,N_24905,N_24891);
nor UO_782 (O_782,N_24759,N_24963);
nor UO_783 (O_783,N_24897,N_24889);
and UO_784 (O_784,N_24777,N_24786);
or UO_785 (O_785,N_24983,N_24962);
nand UO_786 (O_786,N_24922,N_24883);
or UO_787 (O_787,N_24782,N_24818);
and UO_788 (O_788,N_24785,N_24817);
nand UO_789 (O_789,N_24899,N_24792);
nand UO_790 (O_790,N_24948,N_24930);
nor UO_791 (O_791,N_24877,N_24836);
and UO_792 (O_792,N_24917,N_24828);
nor UO_793 (O_793,N_24896,N_24858);
or UO_794 (O_794,N_24835,N_24921);
or UO_795 (O_795,N_24888,N_24819);
nor UO_796 (O_796,N_24935,N_24794);
nand UO_797 (O_797,N_24768,N_24985);
and UO_798 (O_798,N_24969,N_24896);
nor UO_799 (O_799,N_24923,N_24948);
or UO_800 (O_800,N_24898,N_24932);
nand UO_801 (O_801,N_24866,N_24936);
nor UO_802 (O_802,N_24951,N_24955);
and UO_803 (O_803,N_24971,N_24758);
and UO_804 (O_804,N_24773,N_24924);
nor UO_805 (O_805,N_24947,N_24886);
or UO_806 (O_806,N_24829,N_24961);
nor UO_807 (O_807,N_24995,N_24969);
nor UO_808 (O_808,N_24918,N_24843);
nor UO_809 (O_809,N_24777,N_24800);
and UO_810 (O_810,N_24851,N_24826);
nand UO_811 (O_811,N_24771,N_24880);
or UO_812 (O_812,N_24968,N_24985);
nand UO_813 (O_813,N_24855,N_24837);
and UO_814 (O_814,N_24798,N_24952);
nor UO_815 (O_815,N_24801,N_24902);
nor UO_816 (O_816,N_24947,N_24916);
nor UO_817 (O_817,N_24904,N_24878);
nor UO_818 (O_818,N_24752,N_24775);
and UO_819 (O_819,N_24985,N_24912);
nand UO_820 (O_820,N_24854,N_24888);
and UO_821 (O_821,N_24953,N_24911);
nor UO_822 (O_822,N_24771,N_24789);
nand UO_823 (O_823,N_24958,N_24939);
nor UO_824 (O_824,N_24957,N_24971);
and UO_825 (O_825,N_24996,N_24892);
or UO_826 (O_826,N_24810,N_24837);
nor UO_827 (O_827,N_24886,N_24825);
or UO_828 (O_828,N_24868,N_24775);
and UO_829 (O_829,N_24866,N_24911);
nor UO_830 (O_830,N_24897,N_24846);
or UO_831 (O_831,N_24813,N_24828);
nor UO_832 (O_832,N_24898,N_24965);
nand UO_833 (O_833,N_24997,N_24978);
nand UO_834 (O_834,N_24844,N_24768);
and UO_835 (O_835,N_24887,N_24986);
nor UO_836 (O_836,N_24992,N_24878);
nand UO_837 (O_837,N_24790,N_24937);
or UO_838 (O_838,N_24777,N_24957);
nor UO_839 (O_839,N_24753,N_24844);
nand UO_840 (O_840,N_24988,N_24843);
or UO_841 (O_841,N_24819,N_24991);
and UO_842 (O_842,N_24868,N_24797);
and UO_843 (O_843,N_24962,N_24814);
or UO_844 (O_844,N_24790,N_24777);
nand UO_845 (O_845,N_24935,N_24969);
or UO_846 (O_846,N_24969,N_24907);
or UO_847 (O_847,N_24941,N_24772);
nor UO_848 (O_848,N_24970,N_24975);
nor UO_849 (O_849,N_24783,N_24777);
and UO_850 (O_850,N_24847,N_24937);
and UO_851 (O_851,N_24974,N_24980);
or UO_852 (O_852,N_24998,N_24832);
or UO_853 (O_853,N_24990,N_24941);
nor UO_854 (O_854,N_24879,N_24969);
or UO_855 (O_855,N_24867,N_24884);
or UO_856 (O_856,N_24953,N_24995);
or UO_857 (O_857,N_24899,N_24868);
nor UO_858 (O_858,N_24971,N_24892);
nand UO_859 (O_859,N_24943,N_24773);
and UO_860 (O_860,N_24942,N_24909);
nor UO_861 (O_861,N_24785,N_24885);
nor UO_862 (O_862,N_24815,N_24778);
and UO_863 (O_863,N_24907,N_24968);
and UO_864 (O_864,N_24953,N_24958);
nand UO_865 (O_865,N_24827,N_24793);
and UO_866 (O_866,N_24774,N_24793);
and UO_867 (O_867,N_24766,N_24845);
nand UO_868 (O_868,N_24915,N_24906);
nor UO_869 (O_869,N_24979,N_24775);
nor UO_870 (O_870,N_24797,N_24950);
or UO_871 (O_871,N_24946,N_24797);
and UO_872 (O_872,N_24751,N_24971);
nor UO_873 (O_873,N_24881,N_24903);
nand UO_874 (O_874,N_24908,N_24889);
and UO_875 (O_875,N_24816,N_24859);
nor UO_876 (O_876,N_24769,N_24895);
nand UO_877 (O_877,N_24875,N_24977);
nand UO_878 (O_878,N_24952,N_24836);
nand UO_879 (O_879,N_24883,N_24941);
and UO_880 (O_880,N_24818,N_24970);
or UO_881 (O_881,N_24974,N_24990);
nand UO_882 (O_882,N_24949,N_24924);
or UO_883 (O_883,N_24965,N_24887);
nand UO_884 (O_884,N_24916,N_24849);
nand UO_885 (O_885,N_24761,N_24982);
nor UO_886 (O_886,N_24759,N_24895);
nand UO_887 (O_887,N_24914,N_24996);
and UO_888 (O_888,N_24976,N_24842);
or UO_889 (O_889,N_24983,N_24832);
or UO_890 (O_890,N_24775,N_24765);
nor UO_891 (O_891,N_24861,N_24858);
nor UO_892 (O_892,N_24862,N_24812);
nor UO_893 (O_893,N_24754,N_24941);
or UO_894 (O_894,N_24930,N_24825);
or UO_895 (O_895,N_24816,N_24856);
nor UO_896 (O_896,N_24796,N_24842);
nand UO_897 (O_897,N_24980,N_24852);
and UO_898 (O_898,N_24767,N_24993);
and UO_899 (O_899,N_24860,N_24820);
nor UO_900 (O_900,N_24824,N_24862);
nand UO_901 (O_901,N_24901,N_24841);
and UO_902 (O_902,N_24941,N_24957);
nand UO_903 (O_903,N_24870,N_24854);
and UO_904 (O_904,N_24876,N_24838);
nor UO_905 (O_905,N_24982,N_24790);
nand UO_906 (O_906,N_24931,N_24810);
nor UO_907 (O_907,N_24916,N_24928);
or UO_908 (O_908,N_24788,N_24810);
and UO_909 (O_909,N_24862,N_24757);
and UO_910 (O_910,N_24786,N_24986);
or UO_911 (O_911,N_24895,N_24809);
or UO_912 (O_912,N_24842,N_24957);
xor UO_913 (O_913,N_24829,N_24862);
or UO_914 (O_914,N_24771,N_24997);
nor UO_915 (O_915,N_24878,N_24959);
nor UO_916 (O_916,N_24908,N_24965);
nand UO_917 (O_917,N_24901,N_24816);
nand UO_918 (O_918,N_24847,N_24755);
nor UO_919 (O_919,N_24931,N_24922);
or UO_920 (O_920,N_24998,N_24826);
nand UO_921 (O_921,N_24782,N_24847);
or UO_922 (O_922,N_24909,N_24846);
and UO_923 (O_923,N_24880,N_24992);
nand UO_924 (O_924,N_24805,N_24830);
or UO_925 (O_925,N_24812,N_24844);
or UO_926 (O_926,N_24783,N_24875);
or UO_927 (O_927,N_24839,N_24821);
or UO_928 (O_928,N_24778,N_24886);
or UO_929 (O_929,N_24880,N_24918);
and UO_930 (O_930,N_24803,N_24830);
and UO_931 (O_931,N_24797,N_24777);
nand UO_932 (O_932,N_24888,N_24952);
nand UO_933 (O_933,N_24835,N_24892);
or UO_934 (O_934,N_24888,N_24750);
nor UO_935 (O_935,N_24855,N_24974);
and UO_936 (O_936,N_24971,N_24846);
or UO_937 (O_937,N_24817,N_24866);
nor UO_938 (O_938,N_24848,N_24753);
nor UO_939 (O_939,N_24805,N_24845);
and UO_940 (O_940,N_24909,N_24796);
nand UO_941 (O_941,N_24772,N_24998);
nand UO_942 (O_942,N_24850,N_24998);
nor UO_943 (O_943,N_24755,N_24881);
nand UO_944 (O_944,N_24828,N_24984);
nor UO_945 (O_945,N_24947,N_24824);
xnor UO_946 (O_946,N_24800,N_24948);
nand UO_947 (O_947,N_24867,N_24814);
and UO_948 (O_948,N_24943,N_24775);
nand UO_949 (O_949,N_24966,N_24911);
nor UO_950 (O_950,N_24994,N_24848);
or UO_951 (O_951,N_24986,N_24874);
and UO_952 (O_952,N_24987,N_24832);
nand UO_953 (O_953,N_24899,N_24924);
or UO_954 (O_954,N_24837,N_24891);
nand UO_955 (O_955,N_24951,N_24846);
or UO_956 (O_956,N_24850,N_24962);
nand UO_957 (O_957,N_24946,N_24936);
xnor UO_958 (O_958,N_24855,N_24842);
or UO_959 (O_959,N_24944,N_24882);
nor UO_960 (O_960,N_24971,N_24902);
and UO_961 (O_961,N_24751,N_24775);
or UO_962 (O_962,N_24890,N_24868);
nor UO_963 (O_963,N_24881,N_24884);
and UO_964 (O_964,N_24945,N_24885);
and UO_965 (O_965,N_24888,N_24758);
or UO_966 (O_966,N_24896,N_24857);
and UO_967 (O_967,N_24786,N_24769);
and UO_968 (O_968,N_24889,N_24979);
nand UO_969 (O_969,N_24970,N_24999);
and UO_970 (O_970,N_24871,N_24957);
or UO_971 (O_971,N_24967,N_24778);
and UO_972 (O_972,N_24777,N_24921);
nand UO_973 (O_973,N_24881,N_24821);
and UO_974 (O_974,N_24995,N_24876);
nor UO_975 (O_975,N_24902,N_24979);
and UO_976 (O_976,N_24835,N_24788);
and UO_977 (O_977,N_24793,N_24832);
or UO_978 (O_978,N_24770,N_24908);
nor UO_979 (O_979,N_24828,N_24822);
nand UO_980 (O_980,N_24990,N_24751);
xnor UO_981 (O_981,N_24915,N_24945);
or UO_982 (O_982,N_24986,N_24933);
nand UO_983 (O_983,N_24933,N_24931);
nor UO_984 (O_984,N_24890,N_24808);
or UO_985 (O_985,N_24889,N_24875);
nor UO_986 (O_986,N_24974,N_24923);
and UO_987 (O_987,N_24853,N_24756);
nand UO_988 (O_988,N_24929,N_24945);
or UO_989 (O_989,N_24975,N_24843);
nand UO_990 (O_990,N_24798,N_24871);
or UO_991 (O_991,N_24817,N_24773);
or UO_992 (O_992,N_24757,N_24775);
or UO_993 (O_993,N_24920,N_24846);
nor UO_994 (O_994,N_24994,N_24902);
nor UO_995 (O_995,N_24822,N_24961);
and UO_996 (O_996,N_24857,N_24892);
nand UO_997 (O_997,N_24806,N_24913);
and UO_998 (O_998,N_24891,N_24856);
nor UO_999 (O_999,N_24834,N_24908);
or UO_1000 (O_1000,N_24833,N_24972);
and UO_1001 (O_1001,N_24886,N_24988);
nor UO_1002 (O_1002,N_24864,N_24822);
and UO_1003 (O_1003,N_24754,N_24953);
nor UO_1004 (O_1004,N_24807,N_24975);
or UO_1005 (O_1005,N_24930,N_24834);
and UO_1006 (O_1006,N_24946,N_24803);
and UO_1007 (O_1007,N_24808,N_24791);
nand UO_1008 (O_1008,N_24814,N_24841);
and UO_1009 (O_1009,N_24777,N_24810);
nor UO_1010 (O_1010,N_24905,N_24938);
nor UO_1011 (O_1011,N_24832,N_24784);
nor UO_1012 (O_1012,N_24856,N_24967);
or UO_1013 (O_1013,N_24972,N_24835);
nor UO_1014 (O_1014,N_24772,N_24768);
and UO_1015 (O_1015,N_24951,N_24868);
nor UO_1016 (O_1016,N_24935,N_24976);
nand UO_1017 (O_1017,N_24796,N_24775);
and UO_1018 (O_1018,N_24784,N_24943);
or UO_1019 (O_1019,N_24853,N_24813);
or UO_1020 (O_1020,N_24945,N_24820);
and UO_1021 (O_1021,N_24909,N_24785);
and UO_1022 (O_1022,N_24945,N_24812);
or UO_1023 (O_1023,N_24893,N_24903);
nor UO_1024 (O_1024,N_24855,N_24821);
nor UO_1025 (O_1025,N_24867,N_24844);
nor UO_1026 (O_1026,N_24997,N_24780);
and UO_1027 (O_1027,N_24954,N_24922);
or UO_1028 (O_1028,N_24802,N_24987);
nand UO_1029 (O_1029,N_24839,N_24962);
and UO_1030 (O_1030,N_24842,N_24995);
nor UO_1031 (O_1031,N_24879,N_24827);
nor UO_1032 (O_1032,N_24774,N_24823);
nor UO_1033 (O_1033,N_24812,N_24869);
nor UO_1034 (O_1034,N_24995,N_24864);
or UO_1035 (O_1035,N_24793,N_24841);
and UO_1036 (O_1036,N_24997,N_24943);
nor UO_1037 (O_1037,N_24893,N_24858);
nor UO_1038 (O_1038,N_24823,N_24776);
nor UO_1039 (O_1039,N_24938,N_24864);
and UO_1040 (O_1040,N_24876,N_24948);
nand UO_1041 (O_1041,N_24873,N_24939);
or UO_1042 (O_1042,N_24805,N_24963);
and UO_1043 (O_1043,N_24912,N_24791);
and UO_1044 (O_1044,N_24871,N_24902);
or UO_1045 (O_1045,N_24914,N_24838);
or UO_1046 (O_1046,N_24780,N_24919);
nor UO_1047 (O_1047,N_24885,N_24769);
xor UO_1048 (O_1048,N_24932,N_24957);
nor UO_1049 (O_1049,N_24775,N_24832);
nor UO_1050 (O_1050,N_24976,N_24975);
nand UO_1051 (O_1051,N_24821,N_24915);
xnor UO_1052 (O_1052,N_24865,N_24968);
nor UO_1053 (O_1053,N_24827,N_24881);
nor UO_1054 (O_1054,N_24827,N_24849);
nor UO_1055 (O_1055,N_24935,N_24975);
and UO_1056 (O_1056,N_24833,N_24784);
nor UO_1057 (O_1057,N_24781,N_24823);
and UO_1058 (O_1058,N_24772,N_24963);
or UO_1059 (O_1059,N_24787,N_24932);
and UO_1060 (O_1060,N_24837,N_24900);
nand UO_1061 (O_1061,N_24943,N_24886);
xor UO_1062 (O_1062,N_24901,N_24942);
or UO_1063 (O_1063,N_24781,N_24921);
nor UO_1064 (O_1064,N_24807,N_24908);
nor UO_1065 (O_1065,N_24798,N_24954);
and UO_1066 (O_1066,N_24903,N_24911);
nand UO_1067 (O_1067,N_24834,N_24784);
nor UO_1068 (O_1068,N_24906,N_24920);
or UO_1069 (O_1069,N_24776,N_24810);
nand UO_1070 (O_1070,N_24831,N_24933);
nand UO_1071 (O_1071,N_24759,N_24782);
nand UO_1072 (O_1072,N_24890,N_24896);
nor UO_1073 (O_1073,N_24763,N_24887);
or UO_1074 (O_1074,N_24844,N_24783);
nand UO_1075 (O_1075,N_24894,N_24851);
nand UO_1076 (O_1076,N_24978,N_24888);
and UO_1077 (O_1077,N_24804,N_24950);
and UO_1078 (O_1078,N_24753,N_24979);
nand UO_1079 (O_1079,N_24865,N_24880);
or UO_1080 (O_1080,N_24835,N_24994);
and UO_1081 (O_1081,N_24969,N_24859);
nand UO_1082 (O_1082,N_24778,N_24823);
or UO_1083 (O_1083,N_24802,N_24883);
nand UO_1084 (O_1084,N_24795,N_24779);
and UO_1085 (O_1085,N_24895,N_24762);
or UO_1086 (O_1086,N_24969,N_24828);
nand UO_1087 (O_1087,N_24884,N_24822);
nand UO_1088 (O_1088,N_24954,N_24785);
or UO_1089 (O_1089,N_24902,N_24912);
nand UO_1090 (O_1090,N_24961,N_24759);
nand UO_1091 (O_1091,N_24962,N_24924);
or UO_1092 (O_1092,N_24784,N_24993);
or UO_1093 (O_1093,N_24855,N_24944);
or UO_1094 (O_1094,N_24778,N_24803);
nand UO_1095 (O_1095,N_24762,N_24823);
nand UO_1096 (O_1096,N_24887,N_24813);
nand UO_1097 (O_1097,N_24874,N_24960);
nor UO_1098 (O_1098,N_24902,N_24765);
and UO_1099 (O_1099,N_24933,N_24934);
or UO_1100 (O_1100,N_24763,N_24875);
nand UO_1101 (O_1101,N_24940,N_24758);
nand UO_1102 (O_1102,N_24800,N_24973);
or UO_1103 (O_1103,N_24757,N_24834);
nand UO_1104 (O_1104,N_24993,N_24883);
nand UO_1105 (O_1105,N_24989,N_24777);
or UO_1106 (O_1106,N_24912,N_24798);
and UO_1107 (O_1107,N_24913,N_24977);
nor UO_1108 (O_1108,N_24832,N_24927);
nand UO_1109 (O_1109,N_24867,N_24781);
nand UO_1110 (O_1110,N_24851,N_24847);
and UO_1111 (O_1111,N_24848,N_24971);
and UO_1112 (O_1112,N_24772,N_24974);
nor UO_1113 (O_1113,N_24792,N_24978);
nand UO_1114 (O_1114,N_24892,N_24842);
or UO_1115 (O_1115,N_24795,N_24846);
or UO_1116 (O_1116,N_24985,N_24861);
nand UO_1117 (O_1117,N_24933,N_24881);
or UO_1118 (O_1118,N_24875,N_24786);
nand UO_1119 (O_1119,N_24839,N_24825);
or UO_1120 (O_1120,N_24874,N_24863);
and UO_1121 (O_1121,N_24948,N_24758);
or UO_1122 (O_1122,N_24861,N_24833);
or UO_1123 (O_1123,N_24815,N_24888);
or UO_1124 (O_1124,N_24814,N_24860);
and UO_1125 (O_1125,N_24995,N_24800);
or UO_1126 (O_1126,N_24761,N_24938);
or UO_1127 (O_1127,N_24925,N_24846);
or UO_1128 (O_1128,N_24814,N_24988);
nor UO_1129 (O_1129,N_24917,N_24910);
and UO_1130 (O_1130,N_24761,N_24965);
and UO_1131 (O_1131,N_24809,N_24848);
and UO_1132 (O_1132,N_24983,N_24955);
xor UO_1133 (O_1133,N_24834,N_24988);
or UO_1134 (O_1134,N_24792,N_24827);
nand UO_1135 (O_1135,N_24791,N_24756);
and UO_1136 (O_1136,N_24936,N_24952);
nor UO_1137 (O_1137,N_24795,N_24926);
nand UO_1138 (O_1138,N_24877,N_24817);
and UO_1139 (O_1139,N_24959,N_24943);
or UO_1140 (O_1140,N_24807,N_24754);
nor UO_1141 (O_1141,N_24941,N_24872);
and UO_1142 (O_1142,N_24786,N_24802);
nand UO_1143 (O_1143,N_24945,N_24911);
or UO_1144 (O_1144,N_24893,N_24931);
nor UO_1145 (O_1145,N_24841,N_24795);
and UO_1146 (O_1146,N_24821,N_24806);
nand UO_1147 (O_1147,N_24790,N_24833);
or UO_1148 (O_1148,N_24757,N_24916);
or UO_1149 (O_1149,N_24836,N_24819);
or UO_1150 (O_1150,N_24802,N_24847);
nand UO_1151 (O_1151,N_24781,N_24972);
or UO_1152 (O_1152,N_24893,N_24936);
nor UO_1153 (O_1153,N_24758,N_24855);
nor UO_1154 (O_1154,N_24862,N_24971);
nor UO_1155 (O_1155,N_24858,N_24830);
nor UO_1156 (O_1156,N_24921,N_24908);
or UO_1157 (O_1157,N_24946,N_24938);
nand UO_1158 (O_1158,N_24968,N_24855);
nand UO_1159 (O_1159,N_24759,N_24872);
and UO_1160 (O_1160,N_24977,N_24851);
or UO_1161 (O_1161,N_24976,N_24886);
or UO_1162 (O_1162,N_24812,N_24820);
and UO_1163 (O_1163,N_24794,N_24895);
and UO_1164 (O_1164,N_24890,N_24806);
and UO_1165 (O_1165,N_24963,N_24892);
nand UO_1166 (O_1166,N_24956,N_24946);
or UO_1167 (O_1167,N_24992,N_24960);
nor UO_1168 (O_1168,N_24802,N_24871);
and UO_1169 (O_1169,N_24815,N_24876);
or UO_1170 (O_1170,N_24765,N_24828);
and UO_1171 (O_1171,N_24758,N_24837);
nand UO_1172 (O_1172,N_24934,N_24943);
or UO_1173 (O_1173,N_24922,N_24988);
or UO_1174 (O_1174,N_24833,N_24976);
nand UO_1175 (O_1175,N_24954,N_24828);
nand UO_1176 (O_1176,N_24845,N_24869);
nand UO_1177 (O_1177,N_24938,N_24970);
and UO_1178 (O_1178,N_24964,N_24917);
or UO_1179 (O_1179,N_24757,N_24928);
nor UO_1180 (O_1180,N_24948,N_24792);
and UO_1181 (O_1181,N_24807,N_24956);
and UO_1182 (O_1182,N_24868,N_24956);
or UO_1183 (O_1183,N_24785,N_24984);
or UO_1184 (O_1184,N_24886,N_24936);
or UO_1185 (O_1185,N_24808,N_24810);
nand UO_1186 (O_1186,N_24940,N_24765);
nand UO_1187 (O_1187,N_24778,N_24755);
nor UO_1188 (O_1188,N_24978,N_24766);
nor UO_1189 (O_1189,N_24946,N_24823);
and UO_1190 (O_1190,N_24864,N_24781);
or UO_1191 (O_1191,N_24936,N_24873);
or UO_1192 (O_1192,N_24875,N_24774);
or UO_1193 (O_1193,N_24992,N_24946);
and UO_1194 (O_1194,N_24777,N_24941);
and UO_1195 (O_1195,N_24832,N_24810);
or UO_1196 (O_1196,N_24880,N_24948);
nor UO_1197 (O_1197,N_24918,N_24865);
nor UO_1198 (O_1198,N_24799,N_24896);
nand UO_1199 (O_1199,N_24979,N_24795);
nor UO_1200 (O_1200,N_24978,N_24988);
or UO_1201 (O_1201,N_24942,N_24835);
or UO_1202 (O_1202,N_24840,N_24928);
nand UO_1203 (O_1203,N_24929,N_24794);
or UO_1204 (O_1204,N_24860,N_24836);
nand UO_1205 (O_1205,N_24932,N_24852);
nor UO_1206 (O_1206,N_24803,N_24985);
and UO_1207 (O_1207,N_24888,N_24986);
and UO_1208 (O_1208,N_24907,N_24839);
or UO_1209 (O_1209,N_24798,N_24866);
and UO_1210 (O_1210,N_24987,N_24819);
nor UO_1211 (O_1211,N_24836,N_24938);
or UO_1212 (O_1212,N_24785,N_24910);
and UO_1213 (O_1213,N_24806,N_24791);
nor UO_1214 (O_1214,N_24778,N_24788);
and UO_1215 (O_1215,N_24902,N_24924);
or UO_1216 (O_1216,N_24859,N_24955);
nand UO_1217 (O_1217,N_24918,N_24778);
or UO_1218 (O_1218,N_24833,N_24791);
nor UO_1219 (O_1219,N_24773,N_24988);
nor UO_1220 (O_1220,N_24806,N_24973);
or UO_1221 (O_1221,N_24956,N_24755);
or UO_1222 (O_1222,N_24946,N_24824);
nand UO_1223 (O_1223,N_24783,N_24847);
or UO_1224 (O_1224,N_24933,N_24957);
nor UO_1225 (O_1225,N_24914,N_24985);
and UO_1226 (O_1226,N_24919,N_24769);
or UO_1227 (O_1227,N_24896,N_24753);
and UO_1228 (O_1228,N_24850,N_24903);
and UO_1229 (O_1229,N_24822,N_24953);
nor UO_1230 (O_1230,N_24970,N_24794);
nor UO_1231 (O_1231,N_24780,N_24846);
and UO_1232 (O_1232,N_24951,N_24765);
and UO_1233 (O_1233,N_24763,N_24915);
nor UO_1234 (O_1234,N_24859,N_24907);
nor UO_1235 (O_1235,N_24831,N_24958);
nand UO_1236 (O_1236,N_24883,N_24867);
nor UO_1237 (O_1237,N_24839,N_24990);
or UO_1238 (O_1238,N_24866,N_24810);
or UO_1239 (O_1239,N_24835,N_24940);
nor UO_1240 (O_1240,N_24858,N_24885);
and UO_1241 (O_1241,N_24885,N_24880);
xnor UO_1242 (O_1242,N_24871,N_24876);
nor UO_1243 (O_1243,N_24794,N_24994);
nand UO_1244 (O_1244,N_24945,N_24984);
or UO_1245 (O_1245,N_24954,N_24987);
or UO_1246 (O_1246,N_24953,N_24824);
or UO_1247 (O_1247,N_24818,N_24916);
nand UO_1248 (O_1248,N_24793,N_24885);
nor UO_1249 (O_1249,N_24940,N_24967);
nor UO_1250 (O_1250,N_24908,N_24973);
nand UO_1251 (O_1251,N_24810,N_24887);
nor UO_1252 (O_1252,N_24879,N_24782);
nor UO_1253 (O_1253,N_24933,N_24873);
nand UO_1254 (O_1254,N_24957,N_24935);
nor UO_1255 (O_1255,N_24898,N_24911);
and UO_1256 (O_1256,N_24870,N_24957);
and UO_1257 (O_1257,N_24946,N_24795);
or UO_1258 (O_1258,N_24968,N_24887);
and UO_1259 (O_1259,N_24784,N_24911);
and UO_1260 (O_1260,N_24903,N_24858);
nor UO_1261 (O_1261,N_24972,N_24823);
and UO_1262 (O_1262,N_24817,N_24814);
nand UO_1263 (O_1263,N_24972,N_24790);
nor UO_1264 (O_1264,N_24941,N_24975);
nor UO_1265 (O_1265,N_24890,N_24794);
nor UO_1266 (O_1266,N_24990,N_24862);
or UO_1267 (O_1267,N_24923,N_24935);
nor UO_1268 (O_1268,N_24994,N_24960);
or UO_1269 (O_1269,N_24781,N_24787);
nor UO_1270 (O_1270,N_24956,N_24870);
nor UO_1271 (O_1271,N_24843,N_24899);
nand UO_1272 (O_1272,N_24790,N_24987);
nor UO_1273 (O_1273,N_24952,N_24785);
and UO_1274 (O_1274,N_24825,N_24913);
xor UO_1275 (O_1275,N_24756,N_24858);
nor UO_1276 (O_1276,N_24956,N_24816);
or UO_1277 (O_1277,N_24987,N_24750);
nor UO_1278 (O_1278,N_24752,N_24992);
nand UO_1279 (O_1279,N_24826,N_24953);
nor UO_1280 (O_1280,N_24807,N_24753);
or UO_1281 (O_1281,N_24986,N_24827);
nand UO_1282 (O_1282,N_24914,N_24833);
and UO_1283 (O_1283,N_24875,N_24936);
nor UO_1284 (O_1284,N_24912,N_24763);
nand UO_1285 (O_1285,N_24861,N_24936);
nand UO_1286 (O_1286,N_24798,N_24778);
nand UO_1287 (O_1287,N_24966,N_24752);
and UO_1288 (O_1288,N_24988,N_24971);
nand UO_1289 (O_1289,N_24751,N_24794);
nand UO_1290 (O_1290,N_24835,N_24923);
nand UO_1291 (O_1291,N_24788,N_24861);
or UO_1292 (O_1292,N_24980,N_24833);
nand UO_1293 (O_1293,N_24925,N_24859);
or UO_1294 (O_1294,N_24829,N_24993);
and UO_1295 (O_1295,N_24775,N_24974);
and UO_1296 (O_1296,N_24899,N_24828);
nor UO_1297 (O_1297,N_24807,N_24856);
nor UO_1298 (O_1298,N_24891,N_24904);
and UO_1299 (O_1299,N_24839,N_24797);
nand UO_1300 (O_1300,N_24952,N_24981);
nor UO_1301 (O_1301,N_24867,N_24924);
nor UO_1302 (O_1302,N_24857,N_24838);
nor UO_1303 (O_1303,N_24820,N_24862);
nand UO_1304 (O_1304,N_24816,N_24938);
nor UO_1305 (O_1305,N_24773,N_24976);
nor UO_1306 (O_1306,N_24965,N_24872);
nor UO_1307 (O_1307,N_24894,N_24809);
nand UO_1308 (O_1308,N_24997,N_24946);
nand UO_1309 (O_1309,N_24814,N_24946);
nor UO_1310 (O_1310,N_24943,N_24946);
nor UO_1311 (O_1311,N_24977,N_24939);
or UO_1312 (O_1312,N_24821,N_24777);
and UO_1313 (O_1313,N_24866,N_24764);
or UO_1314 (O_1314,N_24845,N_24816);
nand UO_1315 (O_1315,N_24926,N_24755);
nor UO_1316 (O_1316,N_24758,N_24922);
nand UO_1317 (O_1317,N_24856,N_24927);
and UO_1318 (O_1318,N_24812,N_24900);
nand UO_1319 (O_1319,N_24769,N_24802);
nand UO_1320 (O_1320,N_24826,N_24902);
nor UO_1321 (O_1321,N_24899,N_24992);
or UO_1322 (O_1322,N_24995,N_24770);
nor UO_1323 (O_1323,N_24828,N_24780);
nand UO_1324 (O_1324,N_24839,N_24823);
nand UO_1325 (O_1325,N_24879,N_24811);
nand UO_1326 (O_1326,N_24968,N_24767);
and UO_1327 (O_1327,N_24864,N_24796);
nor UO_1328 (O_1328,N_24907,N_24817);
or UO_1329 (O_1329,N_24769,N_24981);
or UO_1330 (O_1330,N_24970,N_24874);
nand UO_1331 (O_1331,N_24952,N_24916);
nor UO_1332 (O_1332,N_24965,N_24774);
or UO_1333 (O_1333,N_24757,N_24848);
nor UO_1334 (O_1334,N_24951,N_24816);
nor UO_1335 (O_1335,N_24769,N_24856);
nand UO_1336 (O_1336,N_24973,N_24887);
nand UO_1337 (O_1337,N_24886,N_24811);
nor UO_1338 (O_1338,N_24967,N_24761);
nor UO_1339 (O_1339,N_24901,N_24957);
or UO_1340 (O_1340,N_24852,N_24984);
or UO_1341 (O_1341,N_24841,N_24834);
or UO_1342 (O_1342,N_24925,N_24901);
nor UO_1343 (O_1343,N_24994,N_24946);
nand UO_1344 (O_1344,N_24943,N_24913);
or UO_1345 (O_1345,N_24940,N_24902);
and UO_1346 (O_1346,N_24921,N_24790);
and UO_1347 (O_1347,N_24848,N_24924);
nand UO_1348 (O_1348,N_24970,N_24764);
and UO_1349 (O_1349,N_24863,N_24993);
nand UO_1350 (O_1350,N_24896,N_24846);
or UO_1351 (O_1351,N_24966,N_24945);
or UO_1352 (O_1352,N_24886,N_24917);
nor UO_1353 (O_1353,N_24963,N_24869);
or UO_1354 (O_1354,N_24906,N_24962);
nor UO_1355 (O_1355,N_24970,N_24916);
or UO_1356 (O_1356,N_24913,N_24781);
nand UO_1357 (O_1357,N_24885,N_24930);
or UO_1358 (O_1358,N_24997,N_24932);
nand UO_1359 (O_1359,N_24928,N_24923);
nor UO_1360 (O_1360,N_24850,N_24926);
or UO_1361 (O_1361,N_24825,N_24887);
nor UO_1362 (O_1362,N_24910,N_24933);
nor UO_1363 (O_1363,N_24755,N_24999);
nand UO_1364 (O_1364,N_24935,N_24797);
nand UO_1365 (O_1365,N_24812,N_24860);
nand UO_1366 (O_1366,N_24963,N_24920);
or UO_1367 (O_1367,N_24948,N_24892);
nor UO_1368 (O_1368,N_24926,N_24995);
nor UO_1369 (O_1369,N_24909,N_24801);
and UO_1370 (O_1370,N_24789,N_24853);
nor UO_1371 (O_1371,N_24823,N_24917);
and UO_1372 (O_1372,N_24855,N_24775);
and UO_1373 (O_1373,N_24854,N_24822);
nor UO_1374 (O_1374,N_24899,N_24760);
or UO_1375 (O_1375,N_24771,N_24840);
or UO_1376 (O_1376,N_24879,N_24852);
or UO_1377 (O_1377,N_24818,N_24955);
and UO_1378 (O_1378,N_24825,N_24784);
and UO_1379 (O_1379,N_24853,N_24787);
nor UO_1380 (O_1380,N_24843,N_24765);
nor UO_1381 (O_1381,N_24925,N_24940);
or UO_1382 (O_1382,N_24877,N_24822);
or UO_1383 (O_1383,N_24945,N_24794);
nand UO_1384 (O_1384,N_24987,N_24923);
nor UO_1385 (O_1385,N_24828,N_24806);
nand UO_1386 (O_1386,N_24882,N_24911);
nor UO_1387 (O_1387,N_24892,N_24897);
or UO_1388 (O_1388,N_24845,N_24928);
nor UO_1389 (O_1389,N_24781,N_24766);
nor UO_1390 (O_1390,N_24939,N_24917);
or UO_1391 (O_1391,N_24914,N_24963);
nor UO_1392 (O_1392,N_24777,N_24874);
nor UO_1393 (O_1393,N_24767,N_24836);
nand UO_1394 (O_1394,N_24878,N_24788);
or UO_1395 (O_1395,N_24896,N_24894);
nand UO_1396 (O_1396,N_24779,N_24851);
nand UO_1397 (O_1397,N_24968,N_24853);
nand UO_1398 (O_1398,N_24912,N_24842);
and UO_1399 (O_1399,N_24899,N_24824);
nand UO_1400 (O_1400,N_24841,N_24994);
and UO_1401 (O_1401,N_24771,N_24937);
nand UO_1402 (O_1402,N_24800,N_24855);
and UO_1403 (O_1403,N_24937,N_24856);
nor UO_1404 (O_1404,N_24971,N_24891);
nand UO_1405 (O_1405,N_24799,N_24753);
or UO_1406 (O_1406,N_24865,N_24842);
and UO_1407 (O_1407,N_24852,N_24816);
nor UO_1408 (O_1408,N_24880,N_24860);
or UO_1409 (O_1409,N_24846,N_24931);
nor UO_1410 (O_1410,N_24776,N_24833);
or UO_1411 (O_1411,N_24857,N_24772);
nand UO_1412 (O_1412,N_24793,N_24881);
nand UO_1413 (O_1413,N_24825,N_24940);
and UO_1414 (O_1414,N_24986,N_24785);
nand UO_1415 (O_1415,N_24798,N_24806);
and UO_1416 (O_1416,N_24965,N_24808);
nand UO_1417 (O_1417,N_24921,N_24848);
nor UO_1418 (O_1418,N_24961,N_24818);
nand UO_1419 (O_1419,N_24913,N_24877);
nand UO_1420 (O_1420,N_24935,N_24980);
or UO_1421 (O_1421,N_24954,N_24776);
nand UO_1422 (O_1422,N_24797,N_24903);
and UO_1423 (O_1423,N_24874,N_24948);
nand UO_1424 (O_1424,N_24788,N_24847);
nor UO_1425 (O_1425,N_24982,N_24873);
and UO_1426 (O_1426,N_24978,N_24985);
nand UO_1427 (O_1427,N_24757,N_24963);
nor UO_1428 (O_1428,N_24877,N_24991);
nor UO_1429 (O_1429,N_24944,N_24845);
and UO_1430 (O_1430,N_24974,N_24913);
or UO_1431 (O_1431,N_24990,N_24905);
and UO_1432 (O_1432,N_24868,N_24982);
or UO_1433 (O_1433,N_24863,N_24780);
nand UO_1434 (O_1434,N_24888,N_24981);
or UO_1435 (O_1435,N_24770,N_24960);
and UO_1436 (O_1436,N_24753,N_24927);
nand UO_1437 (O_1437,N_24821,N_24876);
or UO_1438 (O_1438,N_24982,N_24918);
or UO_1439 (O_1439,N_24959,N_24974);
nand UO_1440 (O_1440,N_24974,N_24754);
and UO_1441 (O_1441,N_24822,N_24964);
nor UO_1442 (O_1442,N_24906,N_24765);
and UO_1443 (O_1443,N_24969,N_24829);
nor UO_1444 (O_1444,N_24775,N_24870);
or UO_1445 (O_1445,N_24805,N_24838);
or UO_1446 (O_1446,N_24969,N_24771);
xor UO_1447 (O_1447,N_24799,N_24868);
and UO_1448 (O_1448,N_24776,N_24907);
and UO_1449 (O_1449,N_24889,N_24851);
or UO_1450 (O_1450,N_24793,N_24845);
and UO_1451 (O_1451,N_24800,N_24993);
and UO_1452 (O_1452,N_24913,N_24896);
xor UO_1453 (O_1453,N_24785,N_24967);
nand UO_1454 (O_1454,N_24930,N_24779);
nand UO_1455 (O_1455,N_24901,N_24879);
nand UO_1456 (O_1456,N_24763,N_24820);
nand UO_1457 (O_1457,N_24842,N_24862);
or UO_1458 (O_1458,N_24939,N_24968);
nand UO_1459 (O_1459,N_24827,N_24991);
nand UO_1460 (O_1460,N_24769,N_24979);
nor UO_1461 (O_1461,N_24988,N_24956);
and UO_1462 (O_1462,N_24962,N_24967);
nor UO_1463 (O_1463,N_24799,N_24966);
nor UO_1464 (O_1464,N_24993,N_24773);
and UO_1465 (O_1465,N_24789,N_24781);
nor UO_1466 (O_1466,N_24998,N_24859);
nand UO_1467 (O_1467,N_24901,N_24820);
nand UO_1468 (O_1468,N_24873,N_24829);
nand UO_1469 (O_1469,N_24973,N_24893);
nor UO_1470 (O_1470,N_24983,N_24944);
or UO_1471 (O_1471,N_24988,N_24954);
and UO_1472 (O_1472,N_24984,N_24915);
and UO_1473 (O_1473,N_24899,N_24794);
and UO_1474 (O_1474,N_24774,N_24921);
and UO_1475 (O_1475,N_24914,N_24869);
nor UO_1476 (O_1476,N_24757,N_24869);
nor UO_1477 (O_1477,N_24903,N_24875);
nand UO_1478 (O_1478,N_24896,N_24775);
nand UO_1479 (O_1479,N_24997,N_24755);
nand UO_1480 (O_1480,N_24823,N_24822);
and UO_1481 (O_1481,N_24892,N_24891);
nand UO_1482 (O_1482,N_24985,N_24910);
nor UO_1483 (O_1483,N_24990,N_24910);
and UO_1484 (O_1484,N_24918,N_24891);
nand UO_1485 (O_1485,N_24888,N_24987);
nor UO_1486 (O_1486,N_24950,N_24796);
nor UO_1487 (O_1487,N_24824,N_24858);
nand UO_1488 (O_1488,N_24926,N_24780);
nand UO_1489 (O_1489,N_24781,N_24863);
or UO_1490 (O_1490,N_24922,N_24893);
nor UO_1491 (O_1491,N_24804,N_24922);
or UO_1492 (O_1492,N_24863,N_24991);
nand UO_1493 (O_1493,N_24814,N_24911);
nand UO_1494 (O_1494,N_24995,N_24933);
or UO_1495 (O_1495,N_24917,N_24950);
nor UO_1496 (O_1496,N_24908,N_24801);
nand UO_1497 (O_1497,N_24835,N_24906);
or UO_1498 (O_1498,N_24864,N_24805);
or UO_1499 (O_1499,N_24780,N_24794);
xor UO_1500 (O_1500,N_24891,N_24776);
nand UO_1501 (O_1501,N_24791,N_24790);
nor UO_1502 (O_1502,N_24787,N_24849);
nor UO_1503 (O_1503,N_24767,N_24945);
or UO_1504 (O_1504,N_24751,N_24917);
nand UO_1505 (O_1505,N_24994,N_24962);
nor UO_1506 (O_1506,N_24937,N_24921);
nor UO_1507 (O_1507,N_24864,N_24978);
or UO_1508 (O_1508,N_24881,N_24750);
and UO_1509 (O_1509,N_24982,N_24911);
nor UO_1510 (O_1510,N_24879,N_24897);
and UO_1511 (O_1511,N_24882,N_24857);
nor UO_1512 (O_1512,N_24968,N_24827);
and UO_1513 (O_1513,N_24874,N_24983);
or UO_1514 (O_1514,N_24898,N_24842);
and UO_1515 (O_1515,N_24756,N_24806);
nand UO_1516 (O_1516,N_24762,N_24959);
and UO_1517 (O_1517,N_24927,N_24780);
nand UO_1518 (O_1518,N_24972,N_24754);
nor UO_1519 (O_1519,N_24833,N_24917);
nor UO_1520 (O_1520,N_24795,N_24861);
nand UO_1521 (O_1521,N_24760,N_24852);
and UO_1522 (O_1522,N_24753,N_24936);
nor UO_1523 (O_1523,N_24961,N_24827);
or UO_1524 (O_1524,N_24966,N_24810);
or UO_1525 (O_1525,N_24889,N_24759);
or UO_1526 (O_1526,N_24761,N_24782);
or UO_1527 (O_1527,N_24778,N_24968);
and UO_1528 (O_1528,N_24758,N_24939);
nand UO_1529 (O_1529,N_24867,N_24869);
nand UO_1530 (O_1530,N_24767,N_24949);
and UO_1531 (O_1531,N_24870,N_24904);
or UO_1532 (O_1532,N_24786,N_24944);
and UO_1533 (O_1533,N_24924,N_24791);
nand UO_1534 (O_1534,N_24860,N_24769);
nand UO_1535 (O_1535,N_24875,N_24917);
nor UO_1536 (O_1536,N_24879,N_24945);
and UO_1537 (O_1537,N_24959,N_24932);
and UO_1538 (O_1538,N_24951,N_24931);
nor UO_1539 (O_1539,N_24776,N_24750);
and UO_1540 (O_1540,N_24766,N_24819);
and UO_1541 (O_1541,N_24868,N_24958);
nor UO_1542 (O_1542,N_24886,N_24895);
nor UO_1543 (O_1543,N_24900,N_24935);
nor UO_1544 (O_1544,N_24757,N_24905);
nand UO_1545 (O_1545,N_24815,N_24987);
or UO_1546 (O_1546,N_24825,N_24860);
nand UO_1547 (O_1547,N_24888,N_24794);
nor UO_1548 (O_1548,N_24838,N_24815);
or UO_1549 (O_1549,N_24819,N_24913);
nand UO_1550 (O_1550,N_24983,N_24958);
nand UO_1551 (O_1551,N_24970,N_24969);
and UO_1552 (O_1552,N_24759,N_24763);
nor UO_1553 (O_1553,N_24817,N_24889);
nand UO_1554 (O_1554,N_24956,N_24853);
nand UO_1555 (O_1555,N_24888,N_24836);
or UO_1556 (O_1556,N_24920,N_24806);
or UO_1557 (O_1557,N_24812,N_24819);
or UO_1558 (O_1558,N_24958,N_24871);
or UO_1559 (O_1559,N_24807,N_24923);
or UO_1560 (O_1560,N_24893,N_24970);
nor UO_1561 (O_1561,N_24822,N_24979);
nor UO_1562 (O_1562,N_24874,N_24808);
and UO_1563 (O_1563,N_24792,N_24911);
nand UO_1564 (O_1564,N_24805,N_24921);
and UO_1565 (O_1565,N_24822,N_24892);
and UO_1566 (O_1566,N_24979,N_24998);
nor UO_1567 (O_1567,N_24945,N_24765);
nor UO_1568 (O_1568,N_24922,N_24909);
or UO_1569 (O_1569,N_24846,N_24927);
and UO_1570 (O_1570,N_24855,N_24889);
or UO_1571 (O_1571,N_24978,N_24965);
nor UO_1572 (O_1572,N_24893,N_24781);
nor UO_1573 (O_1573,N_24823,N_24790);
and UO_1574 (O_1574,N_24918,N_24961);
nor UO_1575 (O_1575,N_24894,N_24971);
or UO_1576 (O_1576,N_24881,N_24899);
nand UO_1577 (O_1577,N_24942,N_24854);
and UO_1578 (O_1578,N_24803,N_24857);
nand UO_1579 (O_1579,N_24817,N_24884);
or UO_1580 (O_1580,N_24952,N_24991);
nor UO_1581 (O_1581,N_24981,N_24870);
nand UO_1582 (O_1582,N_24754,N_24902);
or UO_1583 (O_1583,N_24863,N_24844);
and UO_1584 (O_1584,N_24979,N_24802);
nor UO_1585 (O_1585,N_24923,N_24762);
nor UO_1586 (O_1586,N_24926,N_24972);
and UO_1587 (O_1587,N_24935,N_24843);
or UO_1588 (O_1588,N_24889,N_24990);
or UO_1589 (O_1589,N_24820,N_24907);
nand UO_1590 (O_1590,N_24798,N_24927);
nand UO_1591 (O_1591,N_24868,N_24776);
and UO_1592 (O_1592,N_24874,N_24779);
nor UO_1593 (O_1593,N_24841,N_24912);
nor UO_1594 (O_1594,N_24967,N_24991);
or UO_1595 (O_1595,N_24931,N_24838);
nor UO_1596 (O_1596,N_24800,N_24781);
or UO_1597 (O_1597,N_24980,N_24940);
xor UO_1598 (O_1598,N_24894,N_24838);
nand UO_1599 (O_1599,N_24930,N_24791);
nor UO_1600 (O_1600,N_24760,N_24861);
nor UO_1601 (O_1601,N_24887,N_24991);
or UO_1602 (O_1602,N_24781,N_24993);
or UO_1603 (O_1603,N_24899,N_24995);
nand UO_1604 (O_1604,N_24944,N_24967);
nand UO_1605 (O_1605,N_24795,N_24867);
nor UO_1606 (O_1606,N_24834,N_24795);
nand UO_1607 (O_1607,N_24919,N_24920);
and UO_1608 (O_1608,N_24836,N_24775);
nor UO_1609 (O_1609,N_24998,N_24925);
or UO_1610 (O_1610,N_24865,N_24916);
and UO_1611 (O_1611,N_24998,N_24950);
nand UO_1612 (O_1612,N_24869,N_24776);
or UO_1613 (O_1613,N_24840,N_24834);
or UO_1614 (O_1614,N_24934,N_24801);
nand UO_1615 (O_1615,N_24767,N_24879);
nand UO_1616 (O_1616,N_24955,N_24887);
or UO_1617 (O_1617,N_24912,N_24821);
nor UO_1618 (O_1618,N_24885,N_24953);
or UO_1619 (O_1619,N_24810,N_24911);
nor UO_1620 (O_1620,N_24791,N_24973);
xnor UO_1621 (O_1621,N_24831,N_24925);
nand UO_1622 (O_1622,N_24844,N_24943);
nor UO_1623 (O_1623,N_24866,N_24757);
or UO_1624 (O_1624,N_24884,N_24876);
or UO_1625 (O_1625,N_24856,N_24785);
nor UO_1626 (O_1626,N_24845,N_24976);
or UO_1627 (O_1627,N_24905,N_24954);
nor UO_1628 (O_1628,N_24874,N_24769);
or UO_1629 (O_1629,N_24909,N_24932);
or UO_1630 (O_1630,N_24923,N_24890);
and UO_1631 (O_1631,N_24778,N_24943);
nand UO_1632 (O_1632,N_24845,N_24950);
nand UO_1633 (O_1633,N_24989,N_24776);
nand UO_1634 (O_1634,N_24939,N_24960);
or UO_1635 (O_1635,N_24812,N_24991);
nand UO_1636 (O_1636,N_24813,N_24758);
and UO_1637 (O_1637,N_24763,N_24979);
nor UO_1638 (O_1638,N_24843,N_24768);
and UO_1639 (O_1639,N_24992,N_24832);
nor UO_1640 (O_1640,N_24904,N_24873);
and UO_1641 (O_1641,N_24791,N_24847);
nor UO_1642 (O_1642,N_24800,N_24805);
nor UO_1643 (O_1643,N_24962,N_24951);
nand UO_1644 (O_1644,N_24876,N_24978);
nand UO_1645 (O_1645,N_24968,N_24812);
nor UO_1646 (O_1646,N_24896,N_24984);
nor UO_1647 (O_1647,N_24889,N_24779);
nor UO_1648 (O_1648,N_24816,N_24846);
nand UO_1649 (O_1649,N_24907,N_24804);
or UO_1650 (O_1650,N_24955,N_24902);
and UO_1651 (O_1651,N_24955,N_24927);
or UO_1652 (O_1652,N_24777,N_24857);
or UO_1653 (O_1653,N_24933,N_24780);
or UO_1654 (O_1654,N_24865,N_24770);
nand UO_1655 (O_1655,N_24769,N_24990);
nor UO_1656 (O_1656,N_24854,N_24983);
nand UO_1657 (O_1657,N_24957,N_24880);
and UO_1658 (O_1658,N_24943,N_24980);
and UO_1659 (O_1659,N_24947,N_24806);
and UO_1660 (O_1660,N_24960,N_24811);
and UO_1661 (O_1661,N_24800,N_24825);
nand UO_1662 (O_1662,N_24754,N_24934);
or UO_1663 (O_1663,N_24896,N_24773);
and UO_1664 (O_1664,N_24775,N_24794);
or UO_1665 (O_1665,N_24912,N_24903);
and UO_1666 (O_1666,N_24764,N_24751);
or UO_1667 (O_1667,N_24797,N_24785);
or UO_1668 (O_1668,N_24925,N_24888);
nor UO_1669 (O_1669,N_24825,N_24921);
or UO_1670 (O_1670,N_24840,N_24964);
or UO_1671 (O_1671,N_24961,N_24841);
nand UO_1672 (O_1672,N_24849,N_24844);
or UO_1673 (O_1673,N_24893,N_24874);
nor UO_1674 (O_1674,N_24776,N_24979);
or UO_1675 (O_1675,N_24834,N_24958);
and UO_1676 (O_1676,N_24823,N_24993);
and UO_1677 (O_1677,N_24944,N_24838);
nor UO_1678 (O_1678,N_24808,N_24993);
and UO_1679 (O_1679,N_24858,N_24987);
nor UO_1680 (O_1680,N_24854,N_24997);
or UO_1681 (O_1681,N_24836,N_24960);
nor UO_1682 (O_1682,N_24980,N_24959);
and UO_1683 (O_1683,N_24844,N_24928);
or UO_1684 (O_1684,N_24769,N_24765);
or UO_1685 (O_1685,N_24901,N_24997);
nand UO_1686 (O_1686,N_24778,N_24780);
nor UO_1687 (O_1687,N_24822,N_24885);
or UO_1688 (O_1688,N_24817,N_24790);
nor UO_1689 (O_1689,N_24750,N_24823);
nand UO_1690 (O_1690,N_24831,N_24892);
nand UO_1691 (O_1691,N_24863,N_24931);
nand UO_1692 (O_1692,N_24786,N_24910);
nor UO_1693 (O_1693,N_24789,N_24776);
nand UO_1694 (O_1694,N_24842,N_24878);
or UO_1695 (O_1695,N_24838,N_24917);
or UO_1696 (O_1696,N_24992,N_24839);
or UO_1697 (O_1697,N_24853,N_24826);
nand UO_1698 (O_1698,N_24981,N_24893);
nor UO_1699 (O_1699,N_24940,N_24973);
or UO_1700 (O_1700,N_24974,N_24832);
nand UO_1701 (O_1701,N_24952,N_24965);
nor UO_1702 (O_1702,N_24869,N_24957);
or UO_1703 (O_1703,N_24948,N_24959);
nor UO_1704 (O_1704,N_24897,N_24970);
and UO_1705 (O_1705,N_24782,N_24765);
nor UO_1706 (O_1706,N_24768,N_24767);
nor UO_1707 (O_1707,N_24891,N_24921);
and UO_1708 (O_1708,N_24755,N_24832);
nand UO_1709 (O_1709,N_24772,N_24753);
and UO_1710 (O_1710,N_24873,N_24752);
or UO_1711 (O_1711,N_24801,N_24795);
nor UO_1712 (O_1712,N_24792,N_24906);
and UO_1713 (O_1713,N_24819,N_24929);
nor UO_1714 (O_1714,N_24896,N_24994);
nand UO_1715 (O_1715,N_24986,N_24826);
or UO_1716 (O_1716,N_24881,N_24963);
nand UO_1717 (O_1717,N_24930,N_24865);
and UO_1718 (O_1718,N_24770,N_24902);
and UO_1719 (O_1719,N_24785,N_24800);
nor UO_1720 (O_1720,N_24808,N_24954);
or UO_1721 (O_1721,N_24909,N_24808);
and UO_1722 (O_1722,N_24816,N_24923);
and UO_1723 (O_1723,N_24799,N_24988);
xor UO_1724 (O_1724,N_24819,N_24867);
or UO_1725 (O_1725,N_24874,N_24899);
and UO_1726 (O_1726,N_24800,N_24895);
and UO_1727 (O_1727,N_24927,N_24959);
nand UO_1728 (O_1728,N_24870,N_24823);
and UO_1729 (O_1729,N_24937,N_24931);
and UO_1730 (O_1730,N_24852,N_24869);
nand UO_1731 (O_1731,N_24898,N_24906);
or UO_1732 (O_1732,N_24874,N_24931);
or UO_1733 (O_1733,N_24820,N_24825);
nand UO_1734 (O_1734,N_24835,N_24968);
or UO_1735 (O_1735,N_24970,N_24813);
and UO_1736 (O_1736,N_24942,N_24760);
or UO_1737 (O_1737,N_24773,N_24779);
nor UO_1738 (O_1738,N_24903,N_24982);
or UO_1739 (O_1739,N_24988,N_24876);
or UO_1740 (O_1740,N_24878,N_24944);
nand UO_1741 (O_1741,N_24827,N_24786);
nand UO_1742 (O_1742,N_24970,N_24919);
nand UO_1743 (O_1743,N_24802,N_24929);
nand UO_1744 (O_1744,N_24894,N_24945);
and UO_1745 (O_1745,N_24857,N_24910);
and UO_1746 (O_1746,N_24771,N_24823);
and UO_1747 (O_1747,N_24901,N_24790);
or UO_1748 (O_1748,N_24916,N_24882);
nor UO_1749 (O_1749,N_24928,N_24830);
nand UO_1750 (O_1750,N_24967,N_24989);
and UO_1751 (O_1751,N_24920,N_24841);
nor UO_1752 (O_1752,N_24787,N_24921);
nor UO_1753 (O_1753,N_24980,N_24967);
nor UO_1754 (O_1754,N_24979,N_24892);
or UO_1755 (O_1755,N_24901,N_24952);
and UO_1756 (O_1756,N_24908,N_24958);
nand UO_1757 (O_1757,N_24894,N_24981);
nor UO_1758 (O_1758,N_24914,N_24831);
and UO_1759 (O_1759,N_24854,N_24785);
nand UO_1760 (O_1760,N_24990,N_24837);
or UO_1761 (O_1761,N_24965,N_24936);
or UO_1762 (O_1762,N_24887,N_24981);
or UO_1763 (O_1763,N_24851,N_24780);
and UO_1764 (O_1764,N_24994,N_24890);
nor UO_1765 (O_1765,N_24929,N_24760);
nor UO_1766 (O_1766,N_24850,N_24816);
xnor UO_1767 (O_1767,N_24837,N_24931);
or UO_1768 (O_1768,N_24986,N_24832);
or UO_1769 (O_1769,N_24768,N_24990);
or UO_1770 (O_1770,N_24959,N_24889);
and UO_1771 (O_1771,N_24970,N_24860);
nor UO_1772 (O_1772,N_24980,N_24906);
or UO_1773 (O_1773,N_24940,N_24852);
or UO_1774 (O_1774,N_24774,N_24931);
or UO_1775 (O_1775,N_24969,N_24832);
or UO_1776 (O_1776,N_24835,N_24843);
and UO_1777 (O_1777,N_24878,N_24917);
nor UO_1778 (O_1778,N_24789,N_24788);
and UO_1779 (O_1779,N_24894,N_24794);
nor UO_1780 (O_1780,N_24766,N_24924);
nor UO_1781 (O_1781,N_24955,N_24764);
nor UO_1782 (O_1782,N_24969,N_24936);
nand UO_1783 (O_1783,N_24910,N_24882);
and UO_1784 (O_1784,N_24851,N_24903);
and UO_1785 (O_1785,N_24764,N_24898);
and UO_1786 (O_1786,N_24873,N_24810);
nor UO_1787 (O_1787,N_24994,N_24873);
and UO_1788 (O_1788,N_24943,N_24818);
and UO_1789 (O_1789,N_24966,N_24974);
or UO_1790 (O_1790,N_24781,N_24948);
and UO_1791 (O_1791,N_24995,N_24959);
nor UO_1792 (O_1792,N_24957,N_24804);
or UO_1793 (O_1793,N_24776,N_24771);
xnor UO_1794 (O_1794,N_24756,N_24950);
nor UO_1795 (O_1795,N_24944,N_24938);
and UO_1796 (O_1796,N_24976,N_24909);
nand UO_1797 (O_1797,N_24894,N_24982);
nand UO_1798 (O_1798,N_24853,N_24969);
nand UO_1799 (O_1799,N_24767,N_24815);
or UO_1800 (O_1800,N_24932,N_24885);
xnor UO_1801 (O_1801,N_24791,N_24955);
or UO_1802 (O_1802,N_24907,N_24872);
nand UO_1803 (O_1803,N_24791,N_24830);
and UO_1804 (O_1804,N_24894,N_24958);
nor UO_1805 (O_1805,N_24810,N_24912);
nor UO_1806 (O_1806,N_24935,N_24936);
nand UO_1807 (O_1807,N_24861,N_24989);
and UO_1808 (O_1808,N_24939,N_24957);
nand UO_1809 (O_1809,N_24808,N_24908);
nand UO_1810 (O_1810,N_24754,N_24861);
xor UO_1811 (O_1811,N_24829,N_24853);
nor UO_1812 (O_1812,N_24863,N_24819);
and UO_1813 (O_1813,N_24791,N_24921);
nor UO_1814 (O_1814,N_24824,N_24817);
or UO_1815 (O_1815,N_24762,N_24773);
nor UO_1816 (O_1816,N_24967,N_24922);
nand UO_1817 (O_1817,N_24906,N_24917);
or UO_1818 (O_1818,N_24881,N_24803);
or UO_1819 (O_1819,N_24985,N_24882);
nand UO_1820 (O_1820,N_24945,N_24902);
nor UO_1821 (O_1821,N_24807,N_24840);
or UO_1822 (O_1822,N_24981,N_24796);
and UO_1823 (O_1823,N_24807,N_24904);
nand UO_1824 (O_1824,N_24801,N_24873);
or UO_1825 (O_1825,N_24933,N_24926);
nor UO_1826 (O_1826,N_24788,N_24866);
nand UO_1827 (O_1827,N_24832,N_24979);
nand UO_1828 (O_1828,N_24988,N_24776);
nand UO_1829 (O_1829,N_24837,N_24917);
nand UO_1830 (O_1830,N_24809,N_24930);
nand UO_1831 (O_1831,N_24843,N_24786);
nor UO_1832 (O_1832,N_24923,N_24982);
nand UO_1833 (O_1833,N_24928,N_24811);
or UO_1834 (O_1834,N_24785,N_24832);
nand UO_1835 (O_1835,N_24865,N_24862);
or UO_1836 (O_1836,N_24959,N_24753);
nand UO_1837 (O_1837,N_24885,N_24870);
and UO_1838 (O_1838,N_24968,N_24910);
or UO_1839 (O_1839,N_24900,N_24861);
or UO_1840 (O_1840,N_24949,N_24832);
or UO_1841 (O_1841,N_24800,N_24818);
or UO_1842 (O_1842,N_24839,N_24878);
and UO_1843 (O_1843,N_24929,N_24995);
nor UO_1844 (O_1844,N_24788,N_24905);
and UO_1845 (O_1845,N_24803,N_24947);
nor UO_1846 (O_1846,N_24868,N_24940);
nor UO_1847 (O_1847,N_24797,N_24919);
xnor UO_1848 (O_1848,N_24770,N_24947);
and UO_1849 (O_1849,N_24883,N_24995);
and UO_1850 (O_1850,N_24999,N_24894);
nand UO_1851 (O_1851,N_24844,N_24869);
and UO_1852 (O_1852,N_24933,N_24877);
nor UO_1853 (O_1853,N_24799,N_24818);
and UO_1854 (O_1854,N_24896,N_24978);
and UO_1855 (O_1855,N_24935,N_24752);
and UO_1856 (O_1856,N_24964,N_24985);
nor UO_1857 (O_1857,N_24812,N_24811);
nor UO_1858 (O_1858,N_24963,N_24847);
and UO_1859 (O_1859,N_24900,N_24934);
nand UO_1860 (O_1860,N_24781,N_24974);
nor UO_1861 (O_1861,N_24960,N_24786);
nand UO_1862 (O_1862,N_24910,N_24777);
nor UO_1863 (O_1863,N_24843,N_24991);
or UO_1864 (O_1864,N_24883,N_24943);
and UO_1865 (O_1865,N_24766,N_24761);
and UO_1866 (O_1866,N_24917,N_24919);
nand UO_1867 (O_1867,N_24785,N_24971);
or UO_1868 (O_1868,N_24798,N_24797);
nand UO_1869 (O_1869,N_24969,N_24973);
or UO_1870 (O_1870,N_24961,N_24922);
and UO_1871 (O_1871,N_24813,N_24911);
nor UO_1872 (O_1872,N_24780,N_24829);
or UO_1873 (O_1873,N_24995,N_24793);
or UO_1874 (O_1874,N_24797,N_24960);
and UO_1875 (O_1875,N_24985,N_24907);
or UO_1876 (O_1876,N_24791,N_24803);
and UO_1877 (O_1877,N_24934,N_24979);
and UO_1878 (O_1878,N_24994,N_24963);
nor UO_1879 (O_1879,N_24791,N_24991);
or UO_1880 (O_1880,N_24870,N_24925);
and UO_1881 (O_1881,N_24760,N_24979);
or UO_1882 (O_1882,N_24993,N_24768);
nand UO_1883 (O_1883,N_24813,N_24886);
and UO_1884 (O_1884,N_24953,N_24944);
nor UO_1885 (O_1885,N_24800,N_24838);
nand UO_1886 (O_1886,N_24833,N_24887);
nand UO_1887 (O_1887,N_24849,N_24870);
nor UO_1888 (O_1888,N_24865,N_24777);
or UO_1889 (O_1889,N_24896,N_24933);
nor UO_1890 (O_1890,N_24758,N_24969);
or UO_1891 (O_1891,N_24830,N_24904);
nor UO_1892 (O_1892,N_24895,N_24814);
xor UO_1893 (O_1893,N_24750,N_24794);
and UO_1894 (O_1894,N_24900,N_24933);
nor UO_1895 (O_1895,N_24920,N_24790);
and UO_1896 (O_1896,N_24926,N_24791);
nand UO_1897 (O_1897,N_24751,N_24782);
and UO_1898 (O_1898,N_24871,N_24853);
and UO_1899 (O_1899,N_24939,N_24901);
nor UO_1900 (O_1900,N_24938,N_24899);
and UO_1901 (O_1901,N_24954,N_24766);
or UO_1902 (O_1902,N_24835,N_24930);
nor UO_1903 (O_1903,N_24812,N_24792);
or UO_1904 (O_1904,N_24900,N_24901);
or UO_1905 (O_1905,N_24800,N_24915);
nor UO_1906 (O_1906,N_24782,N_24965);
or UO_1907 (O_1907,N_24906,N_24828);
and UO_1908 (O_1908,N_24932,N_24910);
nor UO_1909 (O_1909,N_24815,N_24775);
nor UO_1910 (O_1910,N_24917,N_24943);
or UO_1911 (O_1911,N_24798,N_24943);
and UO_1912 (O_1912,N_24974,N_24916);
and UO_1913 (O_1913,N_24950,N_24934);
nand UO_1914 (O_1914,N_24838,N_24992);
or UO_1915 (O_1915,N_24856,N_24775);
or UO_1916 (O_1916,N_24762,N_24934);
nand UO_1917 (O_1917,N_24985,N_24816);
and UO_1918 (O_1918,N_24789,N_24831);
or UO_1919 (O_1919,N_24772,N_24797);
nor UO_1920 (O_1920,N_24943,N_24925);
and UO_1921 (O_1921,N_24972,N_24957);
nor UO_1922 (O_1922,N_24967,N_24974);
and UO_1923 (O_1923,N_24999,N_24912);
nand UO_1924 (O_1924,N_24974,N_24972);
or UO_1925 (O_1925,N_24882,N_24881);
nand UO_1926 (O_1926,N_24853,N_24797);
nor UO_1927 (O_1927,N_24901,N_24994);
and UO_1928 (O_1928,N_24754,N_24970);
or UO_1929 (O_1929,N_24772,N_24846);
nand UO_1930 (O_1930,N_24880,N_24778);
nor UO_1931 (O_1931,N_24825,N_24938);
or UO_1932 (O_1932,N_24953,N_24843);
nor UO_1933 (O_1933,N_24800,N_24962);
or UO_1934 (O_1934,N_24920,N_24760);
nand UO_1935 (O_1935,N_24793,N_24868);
nor UO_1936 (O_1936,N_24920,N_24948);
nand UO_1937 (O_1937,N_24780,N_24818);
or UO_1938 (O_1938,N_24956,N_24872);
or UO_1939 (O_1939,N_24962,N_24981);
nand UO_1940 (O_1940,N_24853,N_24964);
or UO_1941 (O_1941,N_24955,N_24809);
or UO_1942 (O_1942,N_24987,N_24957);
nor UO_1943 (O_1943,N_24771,N_24787);
or UO_1944 (O_1944,N_24806,N_24773);
or UO_1945 (O_1945,N_24882,N_24959);
nand UO_1946 (O_1946,N_24780,N_24958);
or UO_1947 (O_1947,N_24955,N_24989);
and UO_1948 (O_1948,N_24889,N_24903);
and UO_1949 (O_1949,N_24968,N_24815);
nand UO_1950 (O_1950,N_24827,N_24870);
nand UO_1951 (O_1951,N_24850,N_24889);
or UO_1952 (O_1952,N_24774,N_24890);
or UO_1953 (O_1953,N_24989,N_24766);
nand UO_1954 (O_1954,N_24829,N_24785);
or UO_1955 (O_1955,N_24997,N_24926);
nand UO_1956 (O_1956,N_24762,N_24908);
and UO_1957 (O_1957,N_24947,N_24831);
nor UO_1958 (O_1958,N_24992,N_24965);
nand UO_1959 (O_1959,N_24907,N_24967);
or UO_1960 (O_1960,N_24923,N_24848);
and UO_1961 (O_1961,N_24969,N_24954);
or UO_1962 (O_1962,N_24899,N_24798);
or UO_1963 (O_1963,N_24934,N_24795);
nor UO_1964 (O_1964,N_24938,N_24915);
nand UO_1965 (O_1965,N_24927,N_24765);
and UO_1966 (O_1966,N_24927,N_24962);
nor UO_1967 (O_1967,N_24922,N_24754);
and UO_1968 (O_1968,N_24801,N_24799);
nor UO_1969 (O_1969,N_24762,N_24856);
nand UO_1970 (O_1970,N_24794,N_24916);
and UO_1971 (O_1971,N_24983,N_24919);
nand UO_1972 (O_1972,N_24858,N_24996);
nor UO_1973 (O_1973,N_24840,N_24992);
nand UO_1974 (O_1974,N_24926,N_24902);
nand UO_1975 (O_1975,N_24923,N_24771);
and UO_1976 (O_1976,N_24781,N_24843);
and UO_1977 (O_1977,N_24807,N_24996);
nand UO_1978 (O_1978,N_24966,N_24903);
or UO_1979 (O_1979,N_24839,N_24786);
nand UO_1980 (O_1980,N_24999,N_24979);
or UO_1981 (O_1981,N_24885,N_24808);
nand UO_1982 (O_1982,N_24936,N_24813);
or UO_1983 (O_1983,N_24774,N_24784);
nand UO_1984 (O_1984,N_24855,N_24795);
nand UO_1985 (O_1985,N_24910,N_24991);
or UO_1986 (O_1986,N_24903,N_24778);
nand UO_1987 (O_1987,N_24850,N_24867);
nand UO_1988 (O_1988,N_24925,N_24950);
and UO_1989 (O_1989,N_24854,N_24977);
nor UO_1990 (O_1990,N_24868,N_24981);
and UO_1991 (O_1991,N_24939,N_24949);
or UO_1992 (O_1992,N_24818,N_24995);
or UO_1993 (O_1993,N_24809,N_24925);
and UO_1994 (O_1994,N_24941,N_24985);
or UO_1995 (O_1995,N_24883,N_24908);
nand UO_1996 (O_1996,N_24778,N_24885);
and UO_1997 (O_1997,N_24860,N_24813);
nor UO_1998 (O_1998,N_24935,N_24829);
nand UO_1999 (O_1999,N_24756,N_24997);
nand UO_2000 (O_2000,N_24966,N_24763);
or UO_2001 (O_2001,N_24783,N_24925);
or UO_2002 (O_2002,N_24844,N_24881);
nor UO_2003 (O_2003,N_24967,N_24809);
and UO_2004 (O_2004,N_24826,N_24860);
nor UO_2005 (O_2005,N_24955,N_24821);
or UO_2006 (O_2006,N_24839,N_24760);
and UO_2007 (O_2007,N_24933,N_24976);
nor UO_2008 (O_2008,N_24985,N_24808);
nand UO_2009 (O_2009,N_24999,N_24781);
nand UO_2010 (O_2010,N_24882,N_24918);
nor UO_2011 (O_2011,N_24800,N_24782);
or UO_2012 (O_2012,N_24923,N_24842);
nand UO_2013 (O_2013,N_24967,N_24958);
or UO_2014 (O_2014,N_24934,N_24910);
or UO_2015 (O_2015,N_24830,N_24861);
or UO_2016 (O_2016,N_24966,N_24940);
nor UO_2017 (O_2017,N_24909,N_24782);
and UO_2018 (O_2018,N_24776,N_24751);
and UO_2019 (O_2019,N_24759,N_24869);
and UO_2020 (O_2020,N_24985,N_24898);
nand UO_2021 (O_2021,N_24845,N_24839);
or UO_2022 (O_2022,N_24889,N_24986);
or UO_2023 (O_2023,N_24923,N_24876);
nand UO_2024 (O_2024,N_24961,N_24836);
and UO_2025 (O_2025,N_24811,N_24937);
nor UO_2026 (O_2026,N_24777,N_24903);
nand UO_2027 (O_2027,N_24837,N_24964);
and UO_2028 (O_2028,N_24875,N_24926);
and UO_2029 (O_2029,N_24981,N_24814);
and UO_2030 (O_2030,N_24960,N_24754);
nand UO_2031 (O_2031,N_24843,N_24969);
and UO_2032 (O_2032,N_24854,N_24856);
or UO_2033 (O_2033,N_24877,N_24893);
nand UO_2034 (O_2034,N_24780,N_24874);
or UO_2035 (O_2035,N_24819,N_24814);
or UO_2036 (O_2036,N_24881,N_24965);
or UO_2037 (O_2037,N_24961,N_24863);
nand UO_2038 (O_2038,N_24921,N_24792);
and UO_2039 (O_2039,N_24860,N_24790);
and UO_2040 (O_2040,N_24836,N_24982);
nand UO_2041 (O_2041,N_24899,N_24879);
nor UO_2042 (O_2042,N_24795,N_24782);
nand UO_2043 (O_2043,N_24981,N_24892);
nand UO_2044 (O_2044,N_24978,N_24764);
and UO_2045 (O_2045,N_24959,N_24861);
nand UO_2046 (O_2046,N_24823,N_24789);
and UO_2047 (O_2047,N_24784,N_24969);
nand UO_2048 (O_2048,N_24849,N_24990);
nor UO_2049 (O_2049,N_24877,N_24995);
nor UO_2050 (O_2050,N_24875,N_24785);
and UO_2051 (O_2051,N_24993,N_24952);
nor UO_2052 (O_2052,N_24910,N_24843);
nand UO_2053 (O_2053,N_24793,N_24814);
nand UO_2054 (O_2054,N_24768,N_24962);
nand UO_2055 (O_2055,N_24931,N_24921);
or UO_2056 (O_2056,N_24843,N_24771);
nor UO_2057 (O_2057,N_24757,N_24751);
nand UO_2058 (O_2058,N_24813,N_24963);
nor UO_2059 (O_2059,N_24901,N_24873);
or UO_2060 (O_2060,N_24872,N_24779);
and UO_2061 (O_2061,N_24795,N_24887);
or UO_2062 (O_2062,N_24914,N_24947);
nand UO_2063 (O_2063,N_24860,N_24780);
xnor UO_2064 (O_2064,N_24853,N_24758);
nor UO_2065 (O_2065,N_24867,N_24804);
and UO_2066 (O_2066,N_24822,N_24760);
or UO_2067 (O_2067,N_24893,N_24928);
or UO_2068 (O_2068,N_24839,N_24919);
and UO_2069 (O_2069,N_24765,N_24885);
or UO_2070 (O_2070,N_24989,N_24826);
or UO_2071 (O_2071,N_24755,N_24890);
xnor UO_2072 (O_2072,N_24968,N_24764);
and UO_2073 (O_2073,N_24762,N_24820);
nor UO_2074 (O_2074,N_24798,N_24896);
or UO_2075 (O_2075,N_24911,N_24851);
or UO_2076 (O_2076,N_24850,N_24876);
and UO_2077 (O_2077,N_24949,N_24833);
nand UO_2078 (O_2078,N_24850,N_24942);
nand UO_2079 (O_2079,N_24839,N_24790);
and UO_2080 (O_2080,N_24969,N_24940);
nor UO_2081 (O_2081,N_24770,N_24915);
nor UO_2082 (O_2082,N_24923,N_24763);
or UO_2083 (O_2083,N_24827,N_24766);
or UO_2084 (O_2084,N_24771,N_24947);
and UO_2085 (O_2085,N_24930,N_24776);
or UO_2086 (O_2086,N_24810,N_24933);
nand UO_2087 (O_2087,N_24960,N_24903);
nor UO_2088 (O_2088,N_24882,N_24906);
nand UO_2089 (O_2089,N_24955,N_24807);
and UO_2090 (O_2090,N_24974,N_24911);
xnor UO_2091 (O_2091,N_24801,N_24890);
nor UO_2092 (O_2092,N_24980,N_24984);
nor UO_2093 (O_2093,N_24824,N_24761);
or UO_2094 (O_2094,N_24967,N_24896);
nand UO_2095 (O_2095,N_24959,N_24922);
nor UO_2096 (O_2096,N_24847,N_24938);
nand UO_2097 (O_2097,N_24839,N_24950);
and UO_2098 (O_2098,N_24798,N_24990);
or UO_2099 (O_2099,N_24846,N_24946);
nand UO_2100 (O_2100,N_24946,N_24973);
or UO_2101 (O_2101,N_24858,N_24892);
nor UO_2102 (O_2102,N_24906,N_24774);
or UO_2103 (O_2103,N_24753,N_24851);
or UO_2104 (O_2104,N_24780,N_24882);
nand UO_2105 (O_2105,N_24961,N_24806);
and UO_2106 (O_2106,N_24795,N_24944);
and UO_2107 (O_2107,N_24846,N_24875);
or UO_2108 (O_2108,N_24935,N_24926);
or UO_2109 (O_2109,N_24847,N_24916);
nand UO_2110 (O_2110,N_24882,N_24811);
or UO_2111 (O_2111,N_24946,N_24843);
and UO_2112 (O_2112,N_24908,N_24826);
or UO_2113 (O_2113,N_24912,N_24939);
or UO_2114 (O_2114,N_24969,N_24972);
nand UO_2115 (O_2115,N_24852,N_24971);
or UO_2116 (O_2116,N_24978,N_24957);
nor UO_2117 (O_2117,N_24754,N_24813);
nand UO_2118 (O_2118,N_24848,N_24898);
and UO_2119 (O_2119,N_24886,N_24884);
and UO_2120 (O_2120,N_24779,N_24842);
and UO_2121 (O_2121,N_24903,N_24832);
and UO_2122 (O_2122,N_24786,N_24824);
nand UO_2123 (O_2123,N_24882,N_24949);
nor UO_2124 (O_2124,N_24868,N_24941);
nand UO_2125 (O_2125,N_24828,N_24905);
or UO_2126 (O_2126,N_24866,N_24935);
nor UO_2127 (O_2127,N_24869,N_24807);
nor UO_2128 (O_2128,N_24875,N_24915);
nand UO_2129 (O_2129,N_24822,N_24755);
nor UO_2130 (O_2130,N_24877,N_24959);
nand UO_2131 (O_2131,N_24907,N_24992);
and UO_2132 (O_2132,N_24772,N_24935);
or UO_2133 (O_2133,N_24787,N_24910);
nor UO_2134 (O_2134,N_24767,N_24791);
or UO_2135 (O_2135,N_24853,N_24814);
and UO_2136 (O_2136,N_24878,N_24916);
nor UO_2137 (O_2137,N_24861,N_24903);
nand UO_2138 (O_2138,N_24954,N_24955);
nand UO_2139 (O_2139,N_24783,N_24936);
or UO_2140 (O_2140,N_24940,N_24887);
nand UO_2141 (O_2141,N_24754,N_24829);
or UO_2142 (O_2142,N_24808,N_24924);
and UO_2143 (O_2143,N_24754,N_24812);
or UO_2144 (O_2144,N_24879,N_24763);
or UO_2145 (O_2145,N_24869,N_24976);
nor UO_2146 (O_2146,N_24814,N_24785);
nor UO_2147 (O_2147,N_24996,N_24859);
nor UO_2148 (O_2148,N_24997,N_24821);
nand UO_2149 (O_2149,N_24786,N_24854);
and UO_2150 (O_2150,N_24916,N_24965);
nor UO_2151 (O_2151,N_24779,N_24759);
nand UO_2152 (O_2152,N_24769,N_24833);
and UO_2153 (O_2153,N_24956,N_24788);
nand UO_2154 (O_2154,N_24797,N_24967);
and UO_2155 (O_2155,N_24813,N_24885);
and UO_2156 (O_2156,N_24967,N_24859);
nand UO_2157 (O_2157,N_24833,N_24934);
nor UO_2158 (O_2158,N_24983,N_24784);
or UO_2159 (O_2159,N_24755,N_24792);
nor UO_2160 (O_2160,N_24808,N_24901);
nor UO_2161 (O_2161,N_24779,N_24891);
nand UO_2162 (O_2162,N_24920,N_24916);
or UO_2163 (O_2163,N_24894,N_24782);
nor UO_2164 (O_2164,N_24931,N_24967);
nor UO_2165 (O_2165,N_24985,N_24847);
nand UO_2166 (O_2166,N_24794,N_24803);
and UO_2167 (O_2167,N_24983,N_24762);
nand UO_2168 (O_2168,N_24914,N_24813);
nand UO_2169 (O_2169,N_24853,N_24751);
or UO_2170 (O_2170,N_24834,N_24876);
and UO_2171 (O_2171,N_24821,N_24910);
or UO_2172 (O_2172,N_24985,N_24777);
and UO_2173 (O_2173,N_24782,N_24919);
and UO_2174 (O_2174,N_24862,N_24818);
nor UO_2175 (O_2175,N_24934,N_24945);
and UO_2176 (O_2176,N_24830,N_24888);
nor UO_2177 (O_2177,N_24803,N_24923);
nor UO_2178 (O_2178,N_24798,N_24826);
or UO_2179 (O_2179,N_24962,N_24961);
and UO_2180 (O_2180,N_24826,N_24837);
or UO_2181 (O_2181,N_24829,N_24941);
or UO_2182 (O_2182,N_24983,N_24846);
and UO_2183 (O_2183,N_24984,N_24978);
nand UO_2184 (O_2184,N_24931,N_24798);
or UO_2185 (O_2185,N_24771,N_24802);
nand UO_2186 (O_2186,N_24873,N_24750);
nand UO_2187 (O_2187,N_24949,N_24974);
or UO_2188 (O_2188,N_24826,N_24802);
nand UO_2189 (O_2189,N_24779,N_24923);
and UO_2190 (O_2190,N_24908,N_24945);
nor UO_2191 (O_2191,N_24988,N_24854);
or UO_2192 (O_2192,N_24939,N_24806);
or UO_2193 (O_2193,N_24880,N_24869);
nand UO_2194 (O_2194,N_24954,N_24879);
or UO_2195 (O_2195,N_24951,N_24770);
or UO_2196 (O_2196,N_24805,N_24987);
and UO_2197 (O_2197,N_24914,N_24776);
nand UO_2198 (O_2198,N_24939,N_24850);
or UO_2199 (O_2199,N_24857,N_24821);
and UO_2200 (O_2200,N_24912,N_24834);
or UO_2201 (O_2201,N_24908,N_24903);
and UO_2202 (O_2202,N_24935,N_24977);
nand UO_2203 (O_2203,N_24883,N_24824);
nand UO_2204 (O_2204,N_24838,N_24933);
or UO_2205 (O_2205,N_24765,N_24806);
and UO_2206 (O_2206,N_24775,N_24930);
nor UO_2207 (O_2207,N_24933,N_24907);
or UO_2208 (O_2208,N_24889,N_24772);
or UO_2209 (O_2209,N_24754,N_24954);
and UO_2210 (O_2210,N_24908,N_24887);
nor UO_2211 (O_2211,N_24856,N_24847);
or UO_2212 (O_2212,N_24777,N_24846);
and UO_2213 (O_2213,N_24766,N_24839);
nor UO_2214 (O_2214,N_24813,N_24794);
and UO_2215 (O_2215,N_24910,N_24975);
or UO_2216 (O_2216,N_24905,N_24956);
and UO_2217 (O_2217,N_24792,N_24833);
or UO_2218 (O_2218,N_24823,N_24753);
or UO_2219 (O_2219,N_24861,N_24952);
and UO_2220 (O_2220,N_24999,N_24919);
nor UO_2221 (O_2221,N_24811,N_24922);
and UO_2222 (O_2222,N_24841,N_24862);
nand UO_2223 (O_2223,N_24920,N_24927);
and UO_2224 (O_2224,N_24761,N_24756);
nand UO_2225 (O_2225,N_24793,N_24783);
nor UO_2226 (O_2226,N_24799,N_24948);
nand UO_2227 (O_2227,N_24822,N_24880);
and UO_2228 (O_2228,N_24943,N_24759);
and UO_2229 (O_2229,N_24960,N_24881);
nand UO_2230 (O_2230,N_24843,N_24875);
nor UO_2231 (O_2231,N_24891,N_24994);
nand UO_2232 (O_2232,N_24852,N_24896);
nor UO_2233 (O_2233,N_24900,N_24930);
and UO_2234 (O_2234,N_24873,N_24869);
nand UO_2235 (O_2235,N_24894,N_24898);
nor UO_2236 (O_2236,N_24963,N_24852);
nor UO_2237 (O_2237,N_24926,N_24787);
or UO_2238 (O_2238,N_24933,N_24879);
or UO_2239 (O_2239,N_24860,N_24980);
nand UO_2240 (O_2240,N_24930,N_24846);
nor UO_2241 (O_2241,N_24822,N_24917);
and UO_2242 (O_2242,N_24819,N_24807);
nor UO_2243 (O_2243,N_24898,N_24884);
nor UO_2244 (O_2244,N_24784,N_24866);
nand UO_2245 (O_2245,N_24891,N_24803);
and UO_2246 (O_2246,N_24870,N_24795);
and UO_2247 (O_2247,N_24863,N_24926);
or UO_2248 (O_2248,N_24993,N_24843);
nand UO_2249 (O_2249,N_24844,N_24855);
or UO_2250 (O_2250,N_24823,N_24956);
nand UO_2251 (O_2251,N_24998,N_24750);
nand UO_2252 (O_2252,N_24923,N_24764);
nand UO_2253 (O_2253,N_24790,N_24875);
and UO_2254 (O_2254,N_24830,N_24881);
nor UO_2255 (O_2255,N_24750,N_24965);
and UO_2256 (O_2256,N_24976,N_24797);
nor UO_2257 (O_2257,N_24969,N_24927);
or UO_2258 (O_2258,N_24859,N_24904);
and UO_2259 (O_2259,N_24875,N_24809);
and UO_2260 (O_2260,N_24855,N_24934);
or UO_2261 (O_2261,N_24864,N_24806);
or UO_2262 (O_2262,N_24895,N_24790);
and UO_2263 (O_2263,N_24972,N_24941);
nand UO_2264 (O_2264,N_24953,N_24796);
and UO_2265 (O_2265,N_24949,N_24792);
nand UO_2266 (O_2266,N_24890,N_24943);
and UO_2267 (O_2267,N_24934,N_24798);
or UO_2268 (O_2268,N_24899,N_24867);
nand UO_2269 (O_2269,N_24989,N_24831);
nand UO_2270 (O_2270,N_24979,N_24971);
or UO_2271 (O_2271,N_24917,N_24932);
and UO_2272 (O_2272,N_24769,N_24923);
nor UO_2273 (O_2273,N_24773,N_24934);
nand UO_2274 (O_2274,N_24886,N_24861);
or UO_2275 (O_2275,N_24925,N_24889);
or UO_2276 (O_2276,N_24977,N_24767);
and UO_2277 (O_2277,N_24924,N_24866);
nand UO_2278 (O_2278,N_24892,N_24784);
nand UO_2279 (O_2279,N_24888,N_24768);
or UO_2280 (O_2280,N_24815,N_24995);
nor UO_2281 (O_2281,N_24903,N_24779);
or UO_2282 (O_2282,N_24841,N_24953);
or UO_2283 (O_2283,N_24987,N_24771);
and UO_2284 (O_2284,N_24866,N_24949);
nor UO_2285 (O_2285,N_24856,N_24872);
and UO_2286 (O_2286,N_24896,N_24983);
and UO_2287 (O_2287,N_24786,N_24856);
or UO_2288 (O_2288,N_24785,N_24893);
nand UO_2289 (O_2289,N_24921,N_24892);
and UO_2290 (O_2290,N_24778,N_24980);
or UO_2291 (O_2291,N_24975,N_24759);
and UO_2292 (O_2292,N_24813,N_24809);
nor UO_2293 (O_2293,N_24877,N_24931);
and UO_2294 (O_2294,N_24883,N_24874);
nand UO_2295 (O_2295,N_24980,N_24937);
or UO_2296 (O_2296,N_24756,N_24921);
and UO_2297 (O_2297,N_24973,N_24801);
and UO_2298 (O_2298,N_24891,N_24998);
nor UO_2299 (O_2299,N_24778,N_24964);
nand UO_2300 (O_2300,N_24993,N_24839);
or UO_2301 (O_2301,N_24870,N_24767);
nor UO_2302 (O_2302,N_24753,N_24908);
nor UO_2303 (O_2303,N_24817,N_24859);
nor UO_2304 (O_2304,N_24896,N_24960);
nor UO_2305 (O_2305,N_24858,N_24959);
or UO_2306 (O_2306,N_24777,N_24812);
xor UO_2307 (O_2307,N_24844,N_24968);
nor UO_2308 (O_2308,N_24795,N_24771);
or UO_2309 (O_2309,N_24821,N_24875);
and UO_2310 (O_2310,N_24991,N_24885);
or UO_2311 (O_2311,N_24819,N_24887);
nand UO_2312 (O_2312,N_24965,N_24906);
and UO_2313 (O_2313,N_24769,N_24774);
or UO_2314 (O_2314,N_24960,N_24937);
nor UO_2315 (O_2315,N_24852,N_24855);
nand UO_2316 (O_2316,N_24993,N_24755);
or UO_2317 (O_2317,N_24936,N_24987);
or UO_2318 (O_2318,N_24920,N_24827);
or UO_2319 (O_2319,N_24928,N_24941);
xor UO_2320 (O_2320,N_24791,N_24933);
nand UO_2321 (O_2321,N_24768,N_24760);
or UO_2322 (O_2322,N_24820,N_24890);
nand UO_2323 (O_2323,N_24774,N_24938);
nand UO_2324 (O_2324,N_24987,N_24883);
nor UO_2325 (O_2325,N_24803,N_24977);
nand UO_2326 (O_2326,N_24961,N_24899);
nor UO_2327 (O_2327,N_24811,N_24946);
nand UO_2328 (O_2328,N_24965,N_24937);
or UO_2329 (O_2329,N_24778,N_24847);
nand UO_2330 (O_2330,N_24992,N_24938);
nand UO_2331 (O_2331,N_24877,N_24910);
nand UO_2332 (O_2332,N_24977,N_24835);
nand UO_2333 (O_2333,N_24781,N_24750);
and UO_2334 (O_2334,N_24989,N_24970);
nor UO_2335 (O_2335,N_24838,N_24809);
nor UO_2336 (O_2336,N_24939,N_24913);
or UO_2337 (O_2337,N_24862,N_24805);
nand UO_2338 (O_2338,N_24781,N_24798);
nor UO_2339 (O_2339,N_24886,N_24869);
and UO_2340 (O_2340,N_24869,N_24796);
nand UO_2341 (O_2341,N_24921,N_24934);
and UO_2342 (O_2342,N_24960,N_24964);
or UO_2343 (O_2343,N_24938,N_24932);
nor UO_2344 (O_2344,N_24821,N_24945);
nand UO_2345 (O_2345,N_24977,N_24774);
or UO_2346 (O_2346,N_24824,N_24779);
or UO_2347 (O_2347,N_24852,N_24998);
and UO_2348 (O_2348,N_24756,N_24939);
nand UO_2349 (O_2349,N_24993,N_24797);
nand UO_2350 (O_2350,N_24787,N_24867);
nor UO_2351 (O_2351,N_24878,N_24905);
and UO_2352 (O_2352,N_24979,N_24951);
nor UO_2353 (O_2353,N_24855,N_24851);
nand UO_2354 (O_2354,N_24878,N_24811);
nand UO_2355 (O_2355,N_24770,N_24936);
and UO_2356 (O_2356,N_24792,N_24790);
nand UO_2357 (O_2357,N_24951,N_24974);
and UO_2358 (O_2358,N_24983,N_24971);
or UO_2359 (O_2359,N_24774,N_24883);
and UO_2360 (O_2360,N_24961,N_24983);
and UO_2361 (O_2361,N_24938,N_24951);
or UO_2362 (O_2362,N_24993,N_24987);
or UO_2363 (O_2363,N_24924,N_24758);
xor UO_2364 (O_2364,N_24878,N_24926);
and UO_2365 (O_2365,N_24883,N_24795);
nand UO_2366 (O_2366,N_24770,N_24871);
and UO_2367 (O_2367,N_24903,N_24975);
nand UO_2368 (O_2368,N_24755,N_24990);
nand UO_2369 (O_2369,N_24782,N_24803);
nor UO_2370 (O_2370,N_24830,N_24934);
nand UO_2371 (O_2371,N_24914,N_24808);
nand UO_2372 (O_2372,N_24771,N_24825);
or UO_2373 (O_2373,N_24795,N_24961);
and UO_2374 (O_2374,N_24980,N_24754);
nor UO_2375 (O_2375,N_24944,N_24762);
and UO_2376 (O_2376,N_24795,N_24876);
nand UO_2377 (O_2377,N_24839,N_24928);
nor UO_2378 (O_2378,N_24886,N_24932);
or UO_2379 (O_2379,N_24821,N_24911);
xor UO_2380 (O_2380,N_24809,N_24841);
nor UO_2381 (O_2381,N_24926,N_24909);
or UO_2382 (O_2382,N_24836,N_24874);
or UO_2383 (O_2383,N_24931,N_24984);
and UO_2384 (O_2384,N_24797,N_24882);
nand UO_2385 (O_2385,N_24777,N_24955);
nor UO_2386 (O_2386,N_24919,N_24931);
nand UO_2387 (O_2387,N_24934,N_24767);
or UO_2388 (O_2388,N_24842,N_24996);
and UO_2389 (O_2389,N_24997,N_24836);
or UO_2390 (O_2390,N_24947,N_24817);
or UO_2391 (O_2391,N_24872,N_24762);
nand UO_2392 (O_2392,N_24780,N_24962);
and UO_2393 (O_2393,N_24788,N_24815);
and UO_2394 (O_2394,N_24917,N_24975);
or UO_2395 (O_2395,N_24845,N_24808);
or UO_2396 (O_2396,N_24752,N_24907);
and UO_2397 (O_2397,N_24986,N_24914);
or UO_2398 (O_2398,N_24929,N_24788);
or UO_2399 (O_2399,N_24756,N_24757);
nand UO_2400 (O_2400,N_24959,N_24945);
and UO_2401 (O_2401,N_24933,N_24798);
or UO_2402 (O_2402,N_24939,N_24993);
nor UO_2403 (O_2403,N_24931,N_24960);
nor UO_2404 (O_2404,N_24897,N_24898);
nand UO_2405 (O_2405,N_24883,N_24957);
and UO_2406 (O_2406,N_24871,N_24807);
nor UO_2407 (O_2407,N_24893,N_24980);
and UO_2408 (O_2408,N_24919,N_24853);
and UO_2409 (O_2409,N_24845,N_24855);
and UO_2410 (O_2410,N_24751,N_24941);
nand UO_2411 (O_2411,N_24783,N_24751);
or UO_2412 (O_2412,N_24945,N_24960);
nand UO_2413 (O_2413,N_24812,N_24852);
nand UO_2414 (O_2414,N_24772,N_24806);
nor UO_2415 (O_2415,N_24759,N_24867);
and UO_2416 (O_2416,N_24754,N_24816);
or UO_2417 (O_2417,N_24984,N_24752);
nand UO_2418 (O_2418,N_24778,N_24804);
nor UO_2419 (O_2419,N_24856,N_24804);
and UO_2420 (O_2420,N_24862,N_24970);
nand UO_2421 (O_2421,N_24847,N_24940);
or UO_2422 (O_2422,N_24842,N_24970);
and UO_2423 (O_2423,N_24869,N_24981);
nor UO_2424 (O_2424,N_24973,N_24774);
or UO_2425 (O_2425,N_24931,N_24900);
and UO_2426 (O_2426,N_24878,N_24785);
and UO_2427 (O_2427,N_24779,N_24987);
and UO_2428 (O_2428,N_24916,N_24770);
nor UO_2429 (O_2429,N_24835,N_24798);
or UO_2430 (O_2430,N_24772,N_24836);
nor UO_2431 (O_2431,N_24886,N_24815);
nor UO_2432 (O_2432,N_24966,N_24972);
nor UO_2433 (O_2433,N_24923,N_24925);
nor UO_2434 (O_2434,N_24975,N_24951);
nor UO_2435 (O_2435,N_24782,N_24928);
or UO_2436 (O_2436,N_24781,N_24874);
and UO_2437 (O_2437,N_24854,N_24984);
and UO_2438 (O_2438,N_24972,N_24773);
nor UO_2439 (O_2439,N_24968,N_24789);
nand UO_2440 (O_2440,N_24863,N_24975);
nand UO_2441 (O_2441,N_24963,N_24975);
nor UO_2442 (O_2442,N_24952,N_24768);
or UO_2443 (O_2443,N_24832,N_24971);
and UO_2444 (O_2444,N_24757,N_24828);
and UO_2445 (O_2445,N_24882,N_24997);
and UO_2446 (O_2446,N_24782,N_24770);
and UO_2447 (O_2447,N_24775,N_24791);
nor UO_2448 (O_2448,N_24945,N_24951);
nand UO_2449 (O_2449,N_24976,N_24966);
nor UO_2450 (O_2450,N_24807,N_24928);
or UO_2451 (O_2451,N_24940,N_24872);
nor UO_2452 (O_2452,N_24943,N_24830);
nor UO_2453 (O_2453,N_24968,N_24796);
nor UO_2454 (O_2454,N_24995,N_24804);
xnor UO_2455 (O_2455,N_24865,N_24898);
or UO_2456 (O_2456,N_24874,N_24920);
or UO_2457 (O_2457,N_24837,N_24995);
and UO_2458 (O_2458,N_24852,N_24854);
nor UO_2459 (O_2459,N_24891,N_24863);
nor UO_2460 (O_2460,N_24831,N_24756);
nor UO_2461 (O_2461,N_24770,N_24832);
or UO_2462 (O_2462,N_24847,N_24868);
nor UO_2463 (O_2463,N_24946,N_24962);
nand UO_2464 (O_2464,N_24981,N_24855);
nand UO_2465 (O_2465,N_24964,N_24771);
and UO_2466 (O_2466,N_24755,N_24829);
xor UO_2467 (O_2467,N_24815,N_24947);
xnor UO_2468 (O_2468,N_24768,N_24886);
or UO_2469 (O_2469,N_24824,N_24787);
or UO_2470 (O_2470,N_24997,N_24972);
and UO_2471 (O_2471,N_24750,N_24905);
nand UO_2472 (O_2472,N_24759,N_24820);
nor UO_2473 (O_2473,N_24981,N_24933);
or UO_2474 (O_2474,N_24937,N_24818);
and UO_2475 (O_2475,N_24934,N_24756);
or UO_2476 (O_2476,N_24922,N_24970);
nand UO_2477 (O_2477,N_24849,N_24909);
or UO_2478 (O_2478,N_24854,N_24834);
and UO_2479 (O_2479,N_24794,N_24936);
or UO_2480 (O_2480,N_24860,N_24842);
or UO_2481 (O_2481,N_24950,N_24979);
and UO_2482 (O_2482,N_24778,N_24795);
or UO_2483 (O_2483,N_24904,N_24797);
and UO_2484 (O_2484,N_24950,N_24952);
and UO_2485 (O_2485,N_24807,N_24974);
nor UO_2486 (O_2486,N_24813,N_24961);
nand UO_2487 (O_2487,N_24853,N_24881);
or UO_2488 (O_2488,N_24984,N_24757);
nand UO_2489 (O_2489,N_24972,N_24923);
or UO_2490 (O_2490,N_24929,N_24913);
or UO_2491 (O_2491,N_24841,N_24759);
nand UO_2492 (O_2492,N_24974,N_24765);
nor UO_2493 (O_2493,N_24911,N_24776);
and UO_2494 (O_2494,N_24782,N_24949);
nand UO_2495 (O_2495,N_24861,N_24984);
or UO_2496 (O_2496,N_24991,N_24896);
or UO_2497 (O_2497,N_24766,N_24959);
nor UO_2498 (O_2498,N_24879,N_24989);
nand UO_2499 (O_2499,N_24988,N_24768);
and UO_2500 (O_2500,N_24795,N_24773);
or UO_2501 (O_2501,N_24949,N_24800);
nand UO_2502 (O_2502,N_24938,N_24763);
nor UO_2503 (O_2503,N_24998,N_24991);
or UO_2504 (O_2504,N_24914,N_24822);
or UO_2505 (O_2505,N_24837,N_24792);
nor UO_2506 (O_2506,N_24902,N_24807);
or UO_2507 (O_2507,N_24963,N_24839);
nor UO_2508 (O_2508,N_24885,N_24955);
nand UO_2509 (O_2509,N_24997,N_24803);
nor UO_2510 (O_2510,N_24809,N_24963);
nand UO_2511 (O_2511,N_24899,N_24942);
or UO_2512 (O_2512,N_24760,N_24994);
nor UO_2513 (O_2513,N_24922,N_24771);
nor UO_2514 (O_2514,N_24852,N_24837);
nand UO_2515 (O_2515,N_24899,N_24758);
or UO_2516 (O_2516,N_24753,N_24836);
nand UO_2517 (O_2517,N_24966,N_24803);
or UO_2518 (O_2518,N_24800,N_24870);
nand UO_2519 (O_2519,N_24830,N_24849);
nor UO_2520 (O_2520,N_24751,N_24752);
nor UO_2521 (O_2521,N_24917,N_24928);
and UO_2522 (O_2522,N_24923,N_24765);
nor UO_2523 (O_2523,N_24794,N_24861);
nor UO_2524 (O_2524,N_24794,N_24909);
nand UO_2525 (O_2525,N_24811,N_24985);
nand UO_2526 (O_2526,N_24908,N_24867);
and UO_2527 (O_2527,N_24895,N_24878);
nand UO_2528 (O_2528,N_24930,N_24770);
and UO_2529 (O_2529,N_24768,N_24960);
and UO_2530 (O_2530,N_24783,N_24807);
nor UO_2531 (O_2531,N_24925,N_24999);
xor UO_2532 (O_2532,N_24813,N_24969);
nand UO_2533 (O_2533,N_24774,N_24885);
nand UO_2534 (O_2534,N_24922,N_24850);
and UO_2535 (O_2535,N_24825,N_24908);
and UO_2536 (O_2536,N_24792,N_24784);
nand UO_2537 (O_2537,N_24958,N_24824);
and UO_2538 (O_2538,N_24961,N_24913);
and UO_2539 (O_2539,N_24764,N_24802);
nand UO_2540 (O_2540,N_24817,N_24970);
nand UO_2541 (O_2541,N_24850,N_24953);
or UO_2542 (O_2542,N_24989,N_24894);
or UO_2543 (O_2543,N_24876,N_24878);
or UO_2544 (O_2544,N_24991,N_24761);
nand UO_2545 (O_2545,N_24835,N_24902);
and UO_2546 (O_2546,N_24895,N_24780);
nor UO_2547 (O_2547,N_24801,N_24972);
or UO_2548 (O_2548,N_24821,N_24916);
or UO_2549 (O_2549,N_24832,N_24806);
and UO_2550 (O_2550,N_24869,N_24883);
or UO_2551 (O_2551,N_24902,N_24963);
and UO_2552 (O_2552,N_24844,N_24979);
and UO_2553 (O_2553,N_24796,N_24998);
or UO_2554 (O_2554,N_24792,N_24852);
and UO_2555 (O_2555,N_24900,N_24955);
nor UO_2556 (O_2556,N_24913,N_24834);
nor UO_2557 (O_2557,N_24955,N_24947);
nor UO_2558 (O_2558,N_24889,N_24882);
and UO_2559 (O_2559,N_24893,N_24996);
nor UO_2560 (O_2560,N_24765,N_24797);
or UO_2561 (O_2561,N_24780,N_24820);
nor UO_2562 (O_2562,N_24875,N_24973);
and UO_2563 (O_2563,N_24976,N_24956);
nor UO_2564 (O_2564,N_24937,N_24787);
nor UO_2565 (O_2565,N_24962,N_24892);
or UO_2566 (O_2566,N_24853,N_24883);
nand UO_2567 (O_2567,N_24762,N_24889);
or UO_2568 (O_2568,N_24919,N_24948);
nand UO_2569 (O_2569,N_24801,N_24866);
and UO_2570 (O_2570,N_24983,N_24942);
nor UO_2571 (O_2571,N_24924,N_24809);
and UO_2572 (O_2572,N_24956,N_24999);
nor UO_2573 (O_2573,N_24950,N_24755);
and UO_2574 (O_2574,N_24770,N_24751);
or UO_2575 (O_2575,N_24823,N_24999);
nand UO_2576 (O_2576,N_24921,N_24785);
or UO_2577 (O_2577,N_24905,N_24758);
nand UO_2578 (O_2578,N_24815,N_24975);
nor UO_2579 (O_2579,N_24846,N_24940);
and UO_2580 (O_2580,N_24803,N_24793);
nand UO_2581 (O_2581,N_24924,N_24817);
or UO_2582 (O_2582,N_24750,N_24974);
nand UO_2583 (O_2583,N_24932,N_24990);
nand UO_2584 (O_2584,N_24813,N_24787);
nand UO_2585 (O_2585,N_24822,N_24898);
nand UO_2586 (O_2586,N_24931,N_24757);
nor UO_2587 (O_2587,N_24972,N_24904);
and UO_2588 (O_2588,N_24895,N_24923);
nand UO_2589 (O_2589,N_24995,N_24786);
nor UO_2590 (O_2590,N_24840,N_24823);
nand UO_2591 (O_2591,N_24884,N_24829);
nor UO_2592 (O_2592,N_24997,N_24829);
nor UO_2593 (O_2593,N_24880,N_24945);
nor UO_2594 (O_2594,N_24827,N_24889);
and UO_2595 (O_2595,N_24902,N_24967);
and UO_2596 (O_2596,N_24928,N_24987);
nor UO_2597 (O_2597,N_24771,N_24973);
nor UO_2598 (O_2598,N_24932,N_24764);
or UO_2599 (O_2599,N_24911,N_24785);
nand UO_2600 (O_2600,N_24783,N_24880);
or UO_2601 (O_2601,N_24843,N_24822);
nand UO_2602 (O_2602,N_24942,N_24826);
nor UO_2603 (O_2603,N_24921,N_24845);
and UO_2604 (O_2604,N_24961,N_24910);
and UO_2605 (O_2605,N_24943,N_24900);
nand UO_2606 (O_2606,N_24913,N_24782);
and UO_2607 (O_2607,N_24947,N_24812);
or UO_2608 (O_2608,N_24951,N_24855);
or UO_2609 (O_2609,N_24917,N_24970);
or UO_2610 (O_2610,N_24839,N_24939);
and UO_2611 (O_2611,N_24831,N_24907);
xnor UO_2612 (O_2612,N_24787,N_24899);
or UO_2613 (O_2613,N_24927,N_24875);
or UO_2614 (O_2614,N_24988,N_24871);
and UO_2615 (O_2615,N_24975,N_24923);
nand UO_2616 (O_2616,N_24852,N_24872);
nor UO_2617 (O_2617,N_24775,N_24787);
and UO_2618 (O_2618,N_24949,N_24776);
and UO_2619 (O_2619,N_24899,N_24761);
nor UO_2620 (O_2620,N_24986,N_24989);
or UO_2621 (O_2621,N_24926,N_24946);
nand UO_2622 (O_2622,N_24976,N_24940);
or UO_2623 (O_2623,N_24835,N_24857);
nor UO_2624 (O_2624,N_24883,N_24878);
nor UO_2625 (O_2625,N_24869,N_24887);
and UO_2626 (O_2626,N_24883,N_24765);
and UO_2627 (O_2627,N_24779,N_24879);
and UO_2628 (O_2628,N_24765,N_24830);
or UO_2629 (O_2629,N_24937,N_24820);
or UO_2630 (O_2630,N_24905,N_24822);
nor UO_2631 (O_2631,N_24886,N_24876);
and UO_2632 (O_2632,N_24882,N_24763);
nand UO_2633 (O_2633,N_24884,N_24920);
and UO_2634 (O_2634,N_24971,N_24913);
nor UO_2635 (O_2635,N_24796,N_24910);
or UO_2636 (O_2636,N_24798,N_24851);
nor UO_2637 (O_2637,N_24772,N_24909);
nor UO_2638 (O_2638,N_24869,N_24829);
and UO_2639 (O_2639,N_24908,N_24816);
or UO_2640 (O_2640,N_24958,N_24919);
and UO_2641 (O_2641,N_24807,N_24849);
and UO_2642 (O_2642,N_24990,N_24867);
and UO_2643 (O_2643,N_24929,N_24847);
nand UO_2644 (O_2644,N_24913,N_24881);
nand UO_2645 (O_2645,N_24858,N_24876);
nand UO_2646 (O_2646,N_24792,N_24851);
nand UO_2647 (O_2647,N_24997,N_24811);
or UO_2648 (O_2648,N_24835,N_24804);
nand UO_2649 (O_2649,N_24753,N_24849);
and UO_2650 (O_2650,N_24886,N_24812);
nor UO_2651 (O_2651,N_24907,N_24803);
nand UO_2652 (O_2652,N_24927,N_24901);
nor UO_2653 (O_2653,N_24860,N_24898);
or UO_2654 (O_2654,N_24771,N_24931);
nor UO_2655 (O_2655,N_24859,N_24845);
and UO_2656 (O_2656,N_24807,N_24987);
nor UO_2657 (O_2657,N_24924,N_24834);
nor UO_2658 (O_2658,N_24975,N_24755);
nor UO_2659 (O_2659,N_24765,N_24957);
and UO_2660 (O_2660,N_24930,N_24990);
nand UO_2661 (O_2661,N_24903,N_24957);
and UO_2662 (O_2662,N_24816,N_24989);
nand UO_2663 (O_2663,N_24853,N_24840);
or UO_2664 (O_2664,N_24802,N_24966);
nand UO_2665 (O_2665,N_24783,N_24930);
or UO_2666 (O_2666,N_24837,N_24987);
nor UO_2667 (O_2667,N_24954,N_24978);
and UO_2668 (O_2668,N_24882,N_24872);
nand UO_2669 (O_2669,N_24830,N_24909);
or UO_2670 (O_2670,N_24870,N_24841);
nor UO_2671 (O_2671,N_24953,N_24927);
or UO_2672 (O_2672,N_24932,N_24971);
or UO_2673 (O_2673,N_24790,N_24976);
or UO_2674 (O_2674,N_24772,N_24862);
nor UO_2675 (O_2675,N_24874,N_24754);
nand UO_2676 (O_2676,N_24979,N_24982);
and UO_2677 (O_2677,N_24968,N_24917);
nand UO_2678 (O_2678,N_24763,N_24848);
and UO_2679 (O_2679,N_24769,N_24842);
and UO_2680 (O_2680,N_24885,N_24807);
and UO_2681 (O_2681,N_24907,N_24974);
nand UO_2682 (O_2682,N_24849,N_24832);
or UO_2683 (O_2683,N_24820,N_24940);
and UO_2684 (O_2684,N_24895,N_24887);
and UO_2685 (O_2685,N_24770,N_24918);
nor UO_2686 (O_2686,N_24801,N_24760);
or UO_2687 (O_2687,N_24764,N_24965);
or UO_2688 (O_2688,N_24820,N_24994);
nor UO_2689 (O_2689,N_24951,N_24971);
or UO_2690 (O_2690,N_24859,N_24872);
nor UO_2691 (O_2691,N_24820,N_24846);
nand UO_2692 (O_2692,N_24804,N_24853);
or UO_2693 (O_2693,N_24875,N_24959);
nand UO_2694 (O_2694,N_24861,N_24935);
nand UO_2695 (O_2695,N_24864,N_24838);
and UO_2696 (O_2696,N_24965,N_24805);
or UO_2697 (O_2697,N_24820,N_24992);
nand UO_2698 (O_2698,N_24822,N_24941);
nand UO_2699 (O_2699,N_24809,N_24941);
nor UO_2700 (O_2700,N_24990,N_24934);
and UO_2701 (O_2701,N_24891,N_24881);
or UO_2702 (O_2702,N_24936,N_24910);
and UO_2703 (O_2703,N_24947,N_24963);
nor UO_2704 (O_2704,N_24921,N_24779);
nor UO_2705 (O_2705,N_24912,N_24869);
nand UO_2706 (O_2706,N_24995,N_24982);
and UO_2707 (O_2707,N_24940,N_24865);
nand UO_2708 (O_2708,N_24962,N_24888);
nand UO_2709 (O_2709,N_24779,N_24866);
or UO_2710 (O_2710,N_24786,N_24938);
nand UO_2711 (O_2711,N_24762,N_24987);
nand UO_2712 (O_2712,N_24771,N_24894);
nand UO_2713 (O_2713,N_24972,N_24917);
nand UO_2714 (O_2714,N_24782,N_24920);
or UO_2715 (O_2715,N_24902,N_24752);
nand UO_2716 (O_2716,N_24773,N_24945);
or UO_2717 (O_2717,N_24779,N_24907);
nor UO_2718 (O_2718,N_24846,N_24864);
nand UO_2719 (O_2719,N_24951,N_24887);
nor UO_2720 (O_2720,N_24993,N_24886);
nand UO_2721 (O_2721,N_24862,N_24916);
nor UO_2722 (O_2722,N_24823,N_24862);
or UO_2723 (O_2723,N_24942,N_24989);
or UO_2724 (O_2724,N_24912,N_24752);
and UO_2725 (O_2725,N_24985,N_24822);
nand UO_2726 (O_2726,N_24950,N_24943);
and UO_2727 (O_2727,N_24955,N_24912);
nor UO_2728 (O_2728,N_24888,N_24991);
nor UO_2729 (O_2729,N_24832,N_24922);
nor UO_2730 (O_2730,N_24853,N_24816);
nand UO_2731 (O_2731,N_24932,N_24825);
or UO_2732 (O_2732,N_24919,N_24836);
nand UO_2733 (O_2733,N_24778,N_24783);
nand UO_2734 (O_2734,N_24801,N_24776);
nor UO_2735 (O_2735,N_24788,N_24942);
nor UO_2736 (O_2736,N_24776,N_24792);
xnor UO_2737 (O_2737,N_24964,N_24821);
or UO_2738 (O_2738,N_24930,N_24884);
nand UO_2739 (O_2739,N_24996,N_24969);
nand UO_2740 (O_2740,N_24814,N_24886);
nand UO_2741 (O_2741,N_24972,N_24765);
and UO_2742 (O_2742,N_24811,N_24785);
nor UO_2743 (O_2743,N_24762,N_24853);
and UO_2744 (O_2744,N_24759,N_24792);
or UO_2745 (O_2745,N_24871,N_24900);
and UO_2746 (O_2746,N_24781,N_24947);
and UO_2747 (O_2747,N_24845,N_24798);
and UO_2748 (O_2748,N_24862,N_24799);
and UO_2749 (O_2749,N_24852,N_24874);
or UO_2750 (O_2750,N_24975,N_24820);
nor UO_2751 (O_2751,N_24964,N_24970);
nor UO_2752 (O_2752,N_24970,N_24934);
and UO_2753 (O_2753,N_24841,N_24828);
nand UO_2754 (O_2754,N_24791,N_24816);
nor UO_2755 (O_2755,N_24991,N_24808);
and UO_2756 (O_2756,N_24960,N_24933);
nand UO_2757 (O_2757,N_24821,N_24946);
and UO_2758 (O_2758,N_24907,N_24884);
or UO_2759 (O_2759,N_24931,N_24988);
and UO_2760 (O_2760,N_24800,N_24844);
nand UO_2761 (O_2761,N_24809,N_24935);
or UO_2762 (O_2762,N_24958,N_24904);
or UO_2763 (O_2763,N_24870,N_24919);
and UO_2764 (O_2764,N_24986,N_24992);
or UO_2765 (O_2765,N_24829,N_24865);
nor UO_2766 (O_2766,N_24861,N_24937);
nor UO_2767 (O_2767,N_24782,N_24868);
or UO_2768 (O_2768,N_24994,N_24763);
or UO_2769 (O_2769,N_24914,N_24965);
and UO_2770 (O_2770,N_24842,N_24820);
or UO_2771 (O_2771,N_24957,N_24809);
or UO_2772 (O_2772,N_24891,N_24973);
nor UO_2773 (O_2773,N_24809,N_24944);
or UO_2774 (O_2774,N_24871,N_24943);
and UO_2775 (O_2775,N_24914,N_24826);
nand UO_2776 (O_2776,N_24980,N_24750);
nand UO_2777 (O_2777,N_24813,N_24869);
and UO_2778 (O_2778,N_24946,N_24765);
or UO_2779 (O_2779,N_24951,N_24803);
or UO_2780 (O_2780,N_24766,N_24928);
nand UO_2781 (O_2781,N_24990,N_24991);
and UO_2782 (O_2782,N_24841,N_24998);
nor UO_2783 (O_2783,N_24992,N_24968);
or UO_2784 (O_2784,N_24957,N_24928);
nand UO_2785 (O_2785,N_24785,N_24862);
and UO_2786 (O_2786,N_24825,N_24917);
nor UO_2787 (O_2787,N_24982,N_24850);
nand UO_2788 (O_2788,N_24926,N_24944);
and UO_2789 (O_2789,N_24830,N_24852);
nand UO_2790 (O_2790,N_24986,N_24842);
and UO_2791 (O_2791,N_24866,N_24840);
nand UO_2792 (O_2792,N_24895,N_24870);
nor UO_2793 (O_2793,N_24911,N_24873);
and UO_2794 (O_2794,N_24906,N_24979);
and UO_2795 (O_2795,N_24840,N_24772);
nor UO_2796 (O_2796,N_24821,N_24976);
nor UO_2797 (O_2797,N_24901,N_24976);
nand UO_2798 (O_2798,N_24984,N_24784);
nor UO_2799 (O_2799,N_24766,N_24915);
nand UO_2800 (O_2800,N_24892,N_24904);
nand UO_2801 (O_2801,N_24837,N_24811);
or UO_2802 (O_2802,N_24790,N_24990);
nand UO_2803 (O_2803,N_24872,N_24772);
nand UO_2804 (O_2804,N_24968,N_24879);
nor UO_2805 (O_2805,N_24815,N_24953);
nand UO_2806 (O_2806,N_24907,N_24954);
or UO_2807 (O_2807,N_24864,N_24899);
nand UO_2808 (O_2808,N_24877,N_24763);
and UO_2809 (O_2809,N_24772,N_24950);
nand UO_2810 (O_2810,N_24794,N_24832);
nor UO_2811 (O_2811,N_24891,N_24875);
nand UO_2812 (O_2812,N_24801,N_24790);
nand UO_2813 (O_2813,N_24954,N_24923);
nor UO_2814 (O_2814,N_24914,N_24829);
or UO_2815 (O_2815,N_24964,N_24841);
and UO_2816 (O_2816,N_24913,N_24917);
nor UO_2817 (O_2817,N_24782,N_24780);
nor UO_2818 (O_2818,N_24838,N_24779);
nand UO_2819 (O_2819,N_24858,N_24785);
or UO_2820 (O_2820,N_24902,N_24938);
nor UO_2821 (O_2821,N_24954,N_24772);
and UO_2822 (O_2822,N_24902,N_24929);
nand UO_2823 (O_2823,N_24876,N_24857);
nor UO_2824 (O_2824,N_24757,N_24899);
and UO_2825 (O_2825,N_24962,N_24842);
and UO_2826 (O_2826,N_24810,N_24794);
nor UO_2827 (O_2827,N_24846,N_24797);
and UO_2828 (O_2828,N_24912,N_24824);
nand UO_2829 (O_2829,N_24845,N_24978);
nor UO_2830 (O_2830,N_24823,N_24852);
nor UO_2831 (O_2831,N_24838,N_24764);
nand UO_2832 (O_2832,N_24989,N_24883);
nor UO_2833 (O_2833,N_24762,N_24792);
nand UO_2834 (O_2834,N_24846,N_24952);
nor UO_2835 (O_2835,N_24943,N_24891);
nand UO_2836 (O_2836,N_24755,N_24902);
and UO_2837 (O_2837,N_24958,N_24799);
or UO_2838 (O_2838,N_24903,N_24843);
and UO_2839 (O_2839,N_24989,N_24931);
nand UO_2840 (O_2840,N_24893,N_24813);
nand UO_2841 (O_2841,N_24823,N_24770);
nor UO_2842 (O_2842,N_24864,N_24786);
and UO_2843 (O_2843,N_24783,N_24795);
or UO_2844 (O_2844,N_24913,N_24849);
or UO_2845 (O_2845,N_24880,N_24924);
or UO_2846 (O_2846,N_24955,N_24778);
and UO_2847 (O_2847,N_24789,N_24978);
or UO_2848 (O_2848,N_24765,N_24921);
nand UO_2849 (O_2849,N_24874,N_24771);
nor UO_2850 (O_2850,N_24965,N_24817);
and UO_2851 (O_2851,N_24980,N_24877);
nand UO_2852 (O_2852,N_24752,N_24943);
nand UO_2853 (O_2853,N_24910,N_24835);
and UO_2854 (O_2854,N_24842,N_24961);
and UO_2855 (O_2855,N_24925,N_24838);
or UO_2856 (O_2856,N_24814,N_24812);
nor UO_2857 (O_2857,N_24807,N_24895);
or UO_2858 (O_2858,N_24821,N_24817);
or UO_2859 (O_2859,N_24901,N_24846);
or UO_2860 (O_2860,N_24806,N_24915);
and UO_2861 (O_2861,N_24942,N_24962);
nor UO_2862 (O_2862,N_24854,N_24827);
and UO_2863 (O_2863,N_24944,N_24843);
xor UO_2864 (O_2864,N_24964,N_24873);
and UO_2865 (O_2865,N_24848,N_24770);
nand UO_2866 (O_2866,N_24872,N_24768);
nand UO_2867 (O_2867,N_24891,N_24946);
and UO_2868 (O_2868,N_24972,N_24807);
or UO_2869 (O_2869,N_24833,N_24960);
or UO_2870 (O_2870,N_24818,N_24829);
or UO_2871 (O_2871,N_24880,N_24888);
or UO_2872 (O_2872,N_24976,N_24798);
and UO_2873 (O_2873,N_24916,N_24805);
xor UO_2874 (O_2874,N_24854,N_24832);
and UO_2875 (O_2875,N_24790,N_24754);
and UO_2876 (O_2876,N_24836,N_24965);
nand UO_2877 (O_2877,N_24843,N_24951);
nor UO_2878 (O_2878,N_24851,N_24810);
nor UO_2879 (O_2879,N_24761,N_24884);
or UO_2880 (O_2880,N_24826,N_24917);
or UO_2881 (O_2881,N_24914,N_24906);
nor UO_2882 (O_2882,N_24915,N_24868);
nand UO_2883 (O_2883,N_24906,N_24806);
nand UO_2884 (O_2884,N_24873,N_24977);
xor UO_2885 (O_2885,N_24759,N_24814);
nor UO_2886 (O_2886,N_24855,N_24962);
or UO_2887 (O_2887,N_24908,N_24950);
or UO_2888 (O_2888,N_24825,N_24922);
nor UO_2889 (O_2889,N_24839,N_24850);
or UO_2890 (O_2890,N_24819,N_24894);
or UO_2891 (O_2891,N_24981,N_24783);
or UO_2892 (O_2892,N_24792,N_24879);
and UO_2893 (O_2893,N_24872,N_24912);
nor UO_2894 (O_2894,N_24860,N_24810);
and UO_2895 (O_2895,N_24774,N_24945);
and UO_2896 (O_2896,N_24754,N_24758);
nor UO_2897 (O_2897,N_24903,N_24932);
or UO_2898 (O_2898,N_24903,N_24768);
nand UO_2899 (O_2899,N_24966,N_24792);
xnor UO_2900 (O_2900,N_24913,N_24941);
or UO_2901 (O_2901,N_24760,N_24857);
and UO_2902 (O_2902,N_24776,N_24827);
nand UO_2903 (O_2903,N_24907,N_24913);
nand UO_2904 (O_2904,N_24809,N_24980);
nand UO_2905 (O_2905,N_24945,N_24854);
and UO_2906 (O_2906,N_24947,N_24940);
and UO_2907 (O_2907,N_24844,N_24980);
nand UO_2908 (O_2908,N_24784,N_24961);
nor UO_2909 (O_2909,N_24856,N_24829);
nor UO_2910 (O_2910,N_24920,N_24840);
or UO_2911 (O_2911,N_24927,N_24993);
or UO_2912 (O_2912,N_24929,N_24761);
xor UO_2913 (O_2913,N_24973,N_24924);
nor UO_2914 (O_2914,N_24841,N_24801);
nand UO_2915 (O_2915,N_24964,N_24842);
nand UO_2916 (O_2916,N_24988,N_24912);
and UO_2917 (O_2917,N_24936,N_24954);
nor UO_2918 (O_2918,N_24794,N_24848);
or UO_2919 (O_2919,N_24755,N_24775);
or UO_2920 (O_2920,N_24906,N_24938);
or UO_2921 (O_2921,N_24784,N_24818);
nor UO_2922 (O_2922,N_24951,N_24760);
and UO_2923 (O_2923,N_24863,N_24914);
nor UO_2924 (O_2924,N_24973,N_24877);
nand UO_2925 (O_2925,N_24859,N_24828);
or UO_2926 (O_2926,N_24816,N_24943);
nand UO_2927 (O_2927,N_24891,N_24967);
nor UO_2928 (O_2928,N_24860,N_24933);
and UO_2929 (O_2929,N_24878,N_24820);
or UO_2930 (O_2930,N_24908,N_24781);
nor UO_2931 (O_2931,N_24963,N_24858);
and UO_2932 (O_2932,N_24851,N_24927);
and UO_2933 (O_2933,N_24914,N_24950);
nor UO_2934 (O_2934,N_24763,N_24768);
nor UO_2935 (O_2935,N_24950,N_24920);
nand UO_2936 (O_2936,N_24771,N_24809);
nand UO_2937 (O_2937,N_24851,N_24835);
or UO_2938 (O_2938,N_24899,N_24849);
or UO_2939 (O_2939,N_24829,N_24784);
and UO_2940 (O_2940,N_24987,N_24894);
nor UO_2941 (O_2941,N_24951,N_24928);
and UO_2942 (O_2942,N_24831,N_24883);
nor UO_2943 (O_2943,N_24951,N_24959);
or UO_2944 (O_2944,N_24945,N_24892);
nand UO_2945 (O_2945,N_24796,N_24870);
and UO_2946 (O_2946,N_24978,N_24844);
or UO_2947 (O_2947,N_24844,N_24945);
and UO_2948 (O_2948,N_24972,N_24758);
and UO_2949 (O_2949,N_24864,N_24828);
or UO_2950 (O_2950,N_24849,N_24792);
nor UO_2951 (O_2951,N_24966,N_24968);
nand UO_2952 (O_2952,N_24755,N_24846);
nand UO_2953 (O_2953,N_24755,N_24923);
or UO_2954 (O_2954,N_24757,N_24985);
nand UO_2955 (O_2955,N_24887,N_24933);
nor UO_2956 (O_2956,N_24818,N_24990);
or UO_2957 (O_2957,N_24950,N_24887);
or UO_2958 (O_2958,N_24950,N_24949);
and UO_2959 (O_2959,N_24965,N_24863);
nand UO_2960 (O_2960,N_24765,N_24854);
or UO_2961 (O_2961,N_24758,N_24870);
and UO_2962 (O_2962,N_24950,N_24838);
nand UO_2963 (O_2963,N_24934,N_24982);
or UO_2964 (O_2964,N_24961,N_24873);
nand UO_2965 (O_2965,N_24974,N_24940);
and UO_2966 (O_2966,N_24869,N_24767);
nand UO_2967 (O_2967,N_24904,N_24981);
or UO_2968 (O_2968,N_24804,N_24887);
and UO_2969 (O_2969,N_24776,N_24850);
and UO_2970 (O_2970,N_24956,N_24859);
or UO_2971 (O_2971,N_24982,N_24801);
nand UO_2972 (O_2972,N_24841,N_24955);
nor UO_2973 (O_2973,N_24982,N_24919);
nand UO_2974 (O_2974,N_24831,N_24880);
nor UO_2975 (O_2975,N_24928,N_24843);
nor UO_2976 (O_2976,N_24811,N_24877);
nand UO_2977 (O_2977,N_24965,N_24795);
or UO_2978 (O_2978,N_24951,N_24961);
nor UO_2979 (O_2979,N_24768,N_24969);
nor UO_2980 (O_2980,N_24756,N_24856);
or UO_2981 (O_2981,N_24922,N_24865);
or UO_2982 (O_2982,N_24971,N_24755);
nor UO_2983 (O_2983,N_24973,N_24939);
or UO_2984 (O_2984,N_24809,N_24876);
or UO_2985 (O_2985,N_24759,N_24908);
and UO_2986 (O_2986,N_24903,N_24870);
nor UO_2987 (O_2987,N_24788,N_24855);
nor UO_2988 (O_2988,N_24758,N_24789);
nand UO_2989 (O_2989,N_24919,N_24811);
and UO_2990 (O_2990,N_24810,N_24773);
nor UO_2991 (O_2991,N_24900,N_24756);
and UO_2992 (O_2992,N_24925,N_24986);
and UO_2993 (O_2993,N_24899,N_24809);
nand UO_2994 (O_2994,N_24979,N_24872);
nor UO_2995 (O_2995,N_24910,N_24898);
nor UO_2996 (O_2996,N_24772,N_24870);
and UO_2997 (O_2997,N_24885,N_24971);
xor UO_2998 (O_2998,N_24885,N_24886);
nand UO_2999 (O_2999,N_24947,N_24905);
endmodule