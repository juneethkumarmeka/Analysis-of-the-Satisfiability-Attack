module basic_750_5000_1000_25_levels_5xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
or U0 (N_0,In_430,In_244);
nor U1 (N_1,In_0,In_688);
and U2 (N_2,In_741,In_297);
or U3 (N_3,In_474,In_260);
and U4 (N_4,In_344,In_480);
nand U5 (N_5,In_740,In_34);
nand U6 (N_6,In_300,In_536);
and U7 (N_7,In_451,In_222);
and U8 (N_8,In_711,In_21);
and U9 (N_9,In_130,In_689);
and U10 (N_10,In_216,In_403);
and U11 (N_11,In_482,In_353);
or U12 (N_12,In_282,In_737);
or U13 (N_13,In_660,In_165);
nand U14 (N_14,In_155,In_184);
xnor U15 (N_15,In_89,In_32);
nor U16 (N_16,In_732,In_734);
and U17 (N_17,In_228,In_475);
xnor U18 (N_18,In_603,In_271);
and U19 (N_19,In_15,In_294);
and U20 (N_20,In_377,In_618);
nor U21 (N_21,In_20,In_70);
nand U22 (N_22,In_29,In_3);
nor U23 (N_23,In_638,In_63);
or U24 (N_24,In_658,In_628);
or U25 (N_25,In_731,In_133);
or U26 (N_26,In_419,In_635);
nand U27 (N_27,In_490,In_37);
or U28 (N_28,In_370,In_306);
xnor U29 (N_29,In_380,In_484);
nor U30 (N_30,In_97,In_22);
nand U31 (N_31,In_647,In_42);
or U32 (N_32,In_366,In_262);
nor U33 (N_33,In_568,In_322);
xnor U34 (N_34,In_295,In_50);
or U35 (N_35,In_381,In_162);
nor U36 (N_36,In_195,In_388);
nor U37 (N_37,In_429,In_398);
nor U38 (N_38,In_213,In_746);
and U39 (N_39,In_329,In_411);
and U40 (N_40,In_446,In_352);
and U41 (N_41,In_717,In_90);
or U42 (N_42,In_41,In_587);
and U43 (N_43,In_11,In_697);
nand U44 (N_44,In_609,In_449);
nand U45 (N_45,In_249,In_566);
nand U46 (N_46,In_85,In_55);
and U47 (N_47,In_721,In_495);
and U48 (N_48,In_576,In_525);
and U49 (N_49,In_650,In_747);
or U50 (N_50,In_448,In_535);
nor U51 (N_51,In_78,In_269);
and U52 (N_52,In_296,In_119);
nor U53 (N_53,In_293,In_643);
and U54 (N_54,In_567,In_48);
and U55 (N_55,In_283,In_542);
nand U56 (N_56,In_455,In_585);
nor U57 (N_57,In_151,In_725);
nor U58 (N_58,In_652,In_376);
nor U59 (N_59,In_524,In_290);
nand U60 (N_60,In_164,In_514);
nor U61 (N_61,In_51,In_40);
or U62 (N_62,In_371,In_2);
or U63 (N_63,In_407,In_553);
nand U64 (N_64,In_320,In_281);
nor U65 (N_65,In_272,In_503);
and U66 (N_66,In_251,In_13);
or U67 (N_67,In_708,In_664);
or U68 (N_68,In_496,In_189);
or U69 (N_69,In_248,In_175);
nor U70 (N_70,In_476,In_236);
nand U71 (N_71,In_325,In_68);
and U72 (N_72,In_543,In_274);
nand U73 (N_73,In_631,In_375);
or U74 (N_74,In_137,In_678);
and U75 (N_75,In_594,In_400);
or U76 (N_76,In_198,In_18);
nand U77 (N_77,In_98,In_44);
or U78 (N_78,In_642,In_280);
or U79 (N_79,In_373,In_277);
nor U80 (N_80,In_554,In_465);
nand U81 (N_81,In_6,In_147);
or U82 (N_82,In_634,In_359);
nor U83 (N_83,In_96,In_405);
or U84 (N_84,In_415,In_580);
and U85 (N_85,In_578,In_588);
and U86 (N_86,In_434,In_232);
or U87 (N_87,In_571,In_64);
and U88 (N_88,In_669,In_592);
and U89 (N_89,In_527,In_569);
xnor U90 (N_90,In_632,In_31);
xor U91 (N_91,In_605,In_74);
or U92 (N_92,In_76,In_606);
and U93 (N_93,In_614,In_245);
xnor U94 (N_94,In_414,In_683);
xnor U95 (N_95,In_461,In_109);
nand U96 (N_96,In_142,In_410);
xnor U97 (N_97,In_182,In_518);
or U98 (N_98,In_462,In_626);
or U99 (N_99,In_512,In_218);
nor U100 (N_100,In_431,In_701);
or U101 (N_101,In_75,In_181);
and U102 (N_102,In_268,In_661);
nor U103 (N_103,In_302,In_129);
nand U104 (N_104,In_674,In_387);
nand U105 (N_105,In_421,In_196);
nand U106 (N_106,In_104,In_315);
nor U107 (N_107,In_612,In_651);
nand U108 (N_108,In_648,In_341);
nand U109 (N_109,In_545,In_368);
xor U110 (N_110,In_197,In_87);
or U111 (N_111,In_173,In_289);
nand U112 (N_112,In_478,In_549);
and U113 (N_113,In_310,In_561);
or U114 (N_114,In_221,In_60);
xnor U115 (N_115,In_397,In_241);
or U116 (N_116,In_105,In_227);
nor U117 (N_117,In_102,In_305);
nand U118 (N_118,In_724,In_103);
nand U119 (N_119,In_59,In_176);
nand U120 (N_120,In_161,In_481);
and U121 (N_121,In_187,In_360);
nor U122 (N_122,In_573,In_7);
nand U123 (N_123,In_625,In_742);
and U124 (N_124,In_439,In_572);
or U125 (N_125,In_443,In_316);
xnor U126 (N_126,In_574,In_728);
nor U127 (N_127,In_676,In_629);
and U128 (N_128,In_125,In_16);
or U129 (N_129,In_672,In_623);
nor U130 (N_130,In_190,In_214);
nand U131 (N_131,In_358,In_257);
and U132 (N_132,In_179,In_158);
nand U133 (N_133,In_499,In_541);
and U134 (N_134,In_203,In_719);
or U135 (N_135,In_327,In_589);
nor U136 (N_136,In_205,In_408);
nand U137 (N_137,In_464,In_347);
nand U138 (N_138,In_229,In_687);
nor U139 (N_139,In_166,In_523);
and U140 (N_140,In_318,In_457);
and U141 (N_141,In_575,In_231);
nand U142 (N_142,In_486,In_428);
or U143 (N_143,In_167,In_77);
and U144 (N_144,In_420,In_171);
or U145 (N_145,In_492,In_186);
and U146 (N_146,In_695,In_286);
or U147 (N_147,In_345,In_440);
and U148 (N_148,In_264,In_378);
and U149 (N_149,In_738,In_406);
or U150 (N_150,In_662,In_533);
and U151 (N_151,In_616,In_510);
and U152 (N_152,In_655,In_361);
and U153 (N_153,In_132,In_255);
nand U154 (N_154,In_511,In_72);
or U155 (N_155,In_385,In_583);
or U156 (N_156,In_624,In_540);
and U157 (N_157,In_694,In_83);
nor U158 (N_158,In_394,In_256);
or U159 (N_159,In_491,In_644);
xnor U160 (N_160,In_143,In_226);
or U161 (N_161,In_577,In_659);
nand U162 (N_162,In_209,In_706);
or U163 (N_163,In_372,In_617);
xnor U164 (N_164,In_562,In_532);
nand U165 (N_165,In_704,In_513);
xnor U166 (N_166,In_416,In_471);
and U167 (N_167,In_299,In_160);
xor U168 (N_168,In_667,In_671);
nor U169 (N_169,In_699,In_364);
or U170 (N_170,In_346,In_93);
nand U171 (N_171,In_319,In_404);
and U172 (N_172,In_253,In_639);
xnor U173 (N_173,In_707,In_590);
nand U174 (N_174,In_714,In_23);
or U175 (N_175,In_680,In_646);
xor U176 (N_176,In_735,In_424);
nor U177 (N_177,In_5,In_350);
or U178 (N_178,In_39,In_450);
or U179 (N_179,In_409,In_399);
or U180 (N_180,In_479,In_30);
nand U181 (N_181,In_716,In_24);
nor U182 (N_182,In_62,In_489);
xnor U183 (N_183,In_131,In_237);
nor U184 (N_184,In_202,In_92);
and U185 (N_185,In_211,In_718);
or U186 (N_186,In_670,In_206);
nor U187 (N_187,In_28,In_52);
nor U188 (N_188,In_663,In_460);
nor U189 (N_189,In_627,In_733);
or U190 (N_190,In_331,In_555);
xnor U191 (N_191,In_247,In_235);
nor U192 (N_192,In_224,In_351);
nor U193 (N_193,In_138,In_116);
nor U194 (N_194,In_111,In_238);
or U195 (N_195,In_212,In_123);
nand U196 (N_196,In_355,In_303);
and U197 (N_197,In_516,In_526);
nand U198 (N_198,In_470,In_56);
or U199 (N_199,In_422,In_563);
nand U200 (N_200,N_101,N_197);
nor U201 (N_201,N_158,In_58);
and U202 (N_202,In_715,In_565);
nor U203 (N_203,In_487,N_44);
xor U204 (N_204,In_630,In_710);
or U205 (N_205,In_615,In_335);
and U206 (N_206,In_654,N_32);
or U207 (N_207,N_23,N_62);
nor U208 (N_208,In_192,N_121);
and U209 (N_209,In_640,N_184);
nand U210 (N_210,N_171,N_10);
or U211 (N_211,In_743,In_323);
or U212 (N_212,N_125,In_602);
or U213 (N_213,N_73,N_130);
and U214 (N_214,In_501,In_447);
nand U215 (N_215,In_657,In_508);
and U216 (N_216,In_180,In_517);
nor U217 (N_217,In_515,In_684);
or U218 (N_218,N_114,In_504);
or U219 (N_219,In_122,In_357);
and U220 (N_220,In_598,In_390);
nand U221 (N_221,N_119,In_270);
or U222 (N_222,In_520,N_98);
nor U223 (N_223,In_656,N_126);
nand U224 (N_224,In_432,In_183);
nor U225 (N_225,N_88,In_595);
nor U226 (N_226,In_284,N_19);
and U227 (N_227,N_38,In_621);
and U228 (N_228,In_149,In_9);
or U229 (N_229,N_156,In_472);
and U230 (N_230,In_273,N_22);
nand U231 (N_231,N_53,In_691);
or U232 (N_232,In_66,In_81);
nand U233 (N_233,In_392,N_8);
and U234 (N_234,In_442,In_321);
and U235 (N_235,N_34,N_166);
nor U236 (N_236,In_497,In_275);
nand U237 (N_237,N_111,N_24);
xor U238 (N_238,In_311,In_703);
nand U239 (N_239,In_54,N_96);
or U240 (N_240,In_210,In_312);
nand U241 (N_241,In_188,N_81);
nand U242 (N_242,In_534,N_31);
nand U243 (N_243,In_313,In_108);
nand U244 (N_244,In_584,In_739);
nand U245 (N_245,N_169,N_113);
and U246 (N_246,In_106,N_122);
and U247 (N_247,In_258,In_225);
nand U248 (N_248,In_134,In_47);
nand U249 (N_249,N_76,N_149);
nor U250 (N_250,In_170,In_367);
or U251 (N_251,N_71,N_164);
nand U252 (N_252,N_68,In_217);
and U253 (N_253,N_77,N_58);
or U254 (N_254,In_596,N_117);
and U255 (N_255,N_192,In_675);
and U256 (N_256,N_139,In_118);
and U257 (N_257,In_342,In_622);
or U258 (N_258,N_28,In_308);
and U259 (N_259,In_36,N_105);
xnor U260 (N_260,In_17,In_292);
or U261 (N_261,In_564,N_141);
or U262 (N_262,N_78,N_48);
or U263 (N_263,In_604,In_425);
nand U264 (N_264,In_494,In_653);
nand U265 (N_265,In_49,In_383);
nand U266 (N_266,N_40,In_88);
and U267 (N_267,In_682,In_417);
nor U268 (N_268,In_298,N_74);
or U269 (N_269,N_102,N_60);
nor U270 (N_270,In_80,In_485);
and U271 (N_271,In_339,In_552);
and U272 (N_272,In_426,In_250);
or U273 (N_273,In_278,In_259);
and U274 (N_274,N_135,N_93);
nand U275 (N_275,N_45,In_722);
or U276 (N_276,In_453,In_4);
nor U277 (N_277,In_110,In_150);
or U278 (N_278,In_727,In_500);
or U279 (N_279,In_379,N_146);
nor U280 (N_280,In_246,N_20);
nor U281 (N_281,N_51,In_698);
xor U282 (N_282,In_673,N_97);
or U283 (N_283,In_267,In_193);
or U284 (N_284,In_681,N_123);
or U285 (N_285,N_147,N_106);
nor U286 (N_286,In_94,In_666);
or U287 (N_287,N_116,N_17);
nand U288 (N_288,N_35,In_506);
and U289 (N_289,In_43,In_240);
or U290 (N_290,N_87,In_729);
nor U291 (N_291,N_167,N_191);
and U292 (N_292,In_522,N_120);
nor U293 (N_293,In_709,In_679);
or U294 (N_294,In_548,N_3);
and U295 (N_295,N_49,In_582);
nor U296 (N_296,N_150,N_7);
or U297 (N_297,In_121,N_85);
or U298 (N_298,N_170,In_692);
and U299 (N_299,N_61,In_649);
nand U300 (N_300,In_570,N_127);
nand U301 (N_301,In_384,N_155);
or U302 (N_302,N_15,N_79);
nor U303 (N_303,N_186,In_477);
or U304 (N_304,In_550,In_730);
nor U305 (N_305,In_597,In_117);
xnor U306 (N_306,In_433,In_276);
and U307 (N_307,N_174,N_140);
and U308 (N_308,In_745,N_134);
or U309 (N_309,N_178,In_113);
xor U310 (N_310,N_54,In_423);
xnor U311 (N_311,N_39,In_334);
and U312 (N_312,N_153,N_115);
xnor U313 (N_313,In_208,In_748);
xor U314 (N_314,N_65,N_132);
or U315 (N_315,In_168,In_362);
nand U316 (N_316,In_645,N_13);
nand U317 (N_317,In_374,In_601);
or U318 (N_318,In_291,In_530);
nand U319 (N_319,In_369,In_437);
or U320 (N_320,N_161,N_30);
nor U321 (N_321,N_70,N_138);
nor U322 (N_322,In_544,In_185);
and U323 (N_323,In_230,In_95);
nor U324 (N_324,In_744,N_108);
and U325 (N_325,In_100,N_162);
nor U326 (N_326,In_389,N_90);
nor U327 (N_327,In_194,In_613);
nor U328 (N_328,In_67,In_233);
or U329 (N_329,In_35,In_713);
and U330 (N_330,N_2,In_463);
or U331 (N_331,In_124,N_1);
xnor U332 (N_332,In_263,In_27);
and U333 (N_333,N_41,In_705);
and U334 (N_334,In_483,N_67);
and U335 (N_335,In_19,N_80);
or U336 (N_336,In_599,In_677);
nor U337 (N_337,N_188,In_586);
and U338 (N_338,In_159,In_396);
and U339 (N_339,N_152,N_50);
or U340 (N_340,In_69,In_363);
nor U341 (N_341,N_143,In_114);
and U342 (N_342,N_92,N_5);
nor U343 (N_343,In_469,In_135);
xnor U344 (N_344,N_100,In_330);
or U345 (N_345,In_45,N_42);
nor U346 (N_346,In_539,N_128);
and U347 (N_347,In_333,In_636);
nor U348 (N_348,N_64,In_99);
and U349 (N_349,In_473,N_185);
or U350 (N_350,In_309,In_157);
nor U351 (N_351,In_607,In_65);
and U352 (N_352,In_239,In_86);
nor U353 (N_353,N_94,In_393);
nand U354 (N_354,In_91,N_129);
nor U355 (N_355,In_12,N_173);
or U356 (N_356,N_0,In_152);
xor U357 (N_357,In_242,In_382);
nand U358 (N_358,In_467,In_163);
nand U359 (N_359,In_243,In_234);
nand U360 (N_360,N_118,In_207);
xnor U361 (N_361,N_72,N_18);
or U362 (N_362,In_509,In_120);
nand U363 (N_363,In_354,In_452);
xnor U364 (N_364,In_386,In_726);
or U365 (N_365,In_73,N_133);
nor U366 (N_366,N_55,In_71);
and U367 (N_367,In_438,N_187);
and U368 (N_368,N_33,N_63);
and U369 (N_369,In_493,In_8);
nor U370 (N_370,N_124,In_26);
or U371 (N_371,In_317,In_82);
xnor U372 (N_372,In_591,In_619);
nand U373 (N_373,In_145,In_547);
and U374 (N_374,In_712,In_172);
or U375 (N_375,N_47,In_140);
nand U376 (N_376,N_4,N_183);
or U377 (N_377,In_529,In_169);
nand U378 (N_378,N_46,In_337);
nand U379 (N_379,N_59,N_189);
nand U380 (N_380,N_11,In_454);
and U381 (N_381,N_82,In_459);
nor U382 (N_382,In_436,N_52);
nand U383 (N_383,In_338,N_195);
xnor U384 (N_384,N_145,N_6);
or U385 (N_385,In_191,In_201);
nor U386 (N_386,In_252,In_314);
nor U387 (N_387,In_488,In_200);
nand U388 (N_388,In_215,In_115);
or U389 (N_389,N_182,In_402);
nand U390 (N_390,In_307,In_127);
nand U391 (N_391,N_142,In_441);
nand U392 (N_392,N_179,In_418);
or U393 (N_393,In_519,In_136);
nor U394 (N_394,N_136,N_21);
xor U395 (N_395,N_194,In_693);
nand U396 (N_396,In_220,In_332);
nor U397 (N_397,N_157,N_16);
or U398 (N_398,In_556,N_27);
nor U399 (N_399,In_177,In_498);
or U400 (N_400,N_103,N_56);
xnor U401 (N_401,N_381,N_86);
nor U402 (N_402,N_159,N_305);
nor U403 (N_403,In_199,N_387);
xnor U404 (N_404,N_256,N_239);
or U405 (N_405,N_356,N_244);
nor U406 (N_406,N_272,N_190);
nor U407 (N_407,N_277,N_209);
nor U408 (N_408,N_237,N_361);
and U409 (N_409,N_375,N_91);
nand U410 (N_410,N_328,N_376);
nor U411 (N_411,In_61,N_388);
or U412 (N_412,N_254,N_260);
and U413 (N_413,In_139,In_466);
nor U414 (N_414,In_25,N_199);
nand U415 (N_415,N_255,N_95);
nor U416 (N_416,N_368,N_215);
or U417 (N_417,In_749,N_303);
or U418 (N_418,N_9,N_193);
nor U419 (N_419,N_234,In_304);
and U420 (N_420,N_261,N_320);
and U421 (N_421,N_296,N_112);
or U422 (N_422,In_608,N_395);
nand U423 (N_423,N_289,N_240);
nand U424 (N_424,N_219,In_458);
nand U425 (N_425,In_33,In_690);
nor U426 (N_426,N_264,N_306);
xnor U427 (N_427,In_1,N_351);
and U428 (N_428,N_270,N_390);
or U429 (N_429,N_276,N_357);
nand U430 (N_430,N_218,N_246);
nor U431 (N_431,N_338,N_373);
nor U432 (N_432,N_257,N_236);
or U433 (N_433,N_224,N_287);
or U434 (N_434,N_229,N_226);
and U435 (N_435,N_252,N_263);
and U436 (N_436,In_356,N_377);
or U437 (N_437,N_332,In_261);
nand U438 (N_438,In_219,N_216);
or U439 (N_439,N_269,N_144);
nor U440 (N_440,N_367,N_363);
or U441 (N_441,N_137,N_109);
nor U442 (N_442,N_366,N_107);
or U443 (N_443,In_254,N_278);
and U444 (N_444,In_620,N_172);
or U445 (N_445,N_175,In_340);
or U446 (N_446,In_156,N_342);
nor U447 (N_447,In_444,N_304);
or U448 (N_448,N_308,N_235);
and U449 (N_449,N_330,In_79);
nor U450 (N_450,N_223,N_371);
or U451 (N_451,In_328,N_352);
nand U452 (N_452,In_557,In_112);
and U453 (N_453,In_528,In_301);
nand U454 (N_454,N_231,N_313);
nor U455 (N_455,N_307,N_220);
xnor U456 (N_456,N_327,In_560);
and U457 (N_457,N_393,N_232);
or U458 (N_458,In_10,N_354);
and U459 (N_459,N_25,N_259);
nor U460 (N_460,N_201,In_287);
or U461 (N_461,In_736,N_383);
and U462 (N_462,N_253,N_394);
nand U463 (N_463,In_505,N_310);
xnor U464 (N_464,N_341,N_372);
and U465 (N_465,In_593,N_285);
or U466 (N_466,N_300,N_360);
nor U467 (N_467,N_359,N_322);
nor U468 (N_468,N_281,In_141);
and U469 (N_469,N_26,N_43);
nor U470 (N_470,N_154,N_200);
and U471 (N_471,In_696,In_413);
or U472 (N_472,N_248,N_347);
nor U473 (N_473,N_283,N_99);
nor U474 (N_474,N_37,N_241);
nand U475 (N_475,In_174,N_397);
nor U476 (N_476,N_317,N_294);
or U477 (N_477,In_531,N_384);
and U478 (N_478,N_316,N_181);
or U479 (N_479,N_318,N_299);
nor U480 (N_480,In_154,N_364);
nor U481 (N_481,N_233,In_558);
nand U482 (N_482,In_502,N_399);
nor U483 (N_483,In_324,N_104);
or U484 (N_484,N_160,N_398);
and U485 (N_485,N_279,N_392);
and U486 (N_486,N_290,In_101);
or U487 (N_487,In_107,In_611);
nor U488 (N_488,N_386,N_326);
nor U489 (N_489,N_271,N_315);
xnor U490 (N_490,In_468,N_291);
and U491 (N_491,In_204,N_83);
or U492 (N_492,N_280,In_288);
nor U493 (N_493,N_230,In_279);
nand U494 (N_494,N_222,In_46);
nand U495 (N_495,N_284,In_57);
nor U496 (N_496,N_66,N_148);
and U497 (N_497,N_228,In_395);
or U498 (N_498,N_391,N_331);
and U499 (N_499,N_309,N_214);
and U500 (N_500,In_685,N_225);
and U501 (N_501,N_221,N_337);
or U502 (N_502,N_266,N_345);
and U503 (N_503,N_319,In_600);
and U504 (N_504,N_324,In_579);
xor U505 (N_505,N_89,In_551);
nor U506 (N_506,N_274,In_637);
nor U507 (N_507,In_427,In_412);
xnor U508 (N_508,N_333,In_538);
or U509 (N_509,In_178,N_336);
or U510 (N_510,N_335,N_355);
and U511 (N_511,N_245,In_146);
and U512 (N_512,N_302,N_168);
nor U513 (N_513,N_12,In_391);
or U514 (N_514,In_559,N_348);
xnor U515 (N_515,N_349,N_379);
and U516 (N_516,In_343,N_288);
xor U517 (N_517,In_665,N_208);
nand U518 (N_518,In_285,In_266);
and U519 (N_519,N_374,In_53);
nor U520 (N_520,N_268,N_212);
nor U521 (N_521,N_389,N_227);
nand U522 (N_522,In_546,N_365);
nand U523 (N_523,N_370,N_84);
nor U524 (N_524,N_273,In_507);
nor U525 (N_525,In_435,N_110);
and U526 (N_526,N_211,N_380);
nand U527 (N_527,N_292,In_641);
or U528 (N_528,N_382,In_348);
or U529 (N_529,In_581,N_131);
and U530 (N_530,N_343,N_385);
nand U531 (N_531,N_75,N_265);
xnor U532 (N_532,N_314,N_282);
or U533 (N_533,N_262,N_242);
or U534 (N_534,In_128,N_340);
or U535 (N_535,N_286,N_210);
nand U536 (N_536,N_312,N_323);
and U537 (N_537,N_176,N_198);
xnor U538 (N_538,N_69,In_126);
nor U539 (N_539,N_151,In_144);
or U540 (N_540,In_148,N_258);
nand U541 (N_541,In_38,N_202);
xor U542 (N_542,N_350,N_369);
nor U543 (N_543,N_295,N_396);
or U544 (N_544,In_686,In_700);
xnor U545 (N_545,N_180,N_36);
or U546 (N_546,In_14,N_29);
nor U547 (N_547,N_301,N_196);
nand U548 (N_548,In_633,N_249);
nor U549 (N_549,In_702,N_329);
nor U550 (N_550,In_153,N_298);
and U551 (N_551,N_344,N_205);
and U552 (N_552,N_325,N_378);
or U553 (N_553,In_445,N_346);
or U554 (N_554,N_14,N_207);
or U555 (N_555,In_326,N_358);
nor U556 (N_556,In_265,N_217);
and U557 (N_557,In_537,In_223);
xor U558 (N_558,N_165,In_723);
and U559 (N_559,N_311,N_321);
nand U560 (N_560,N_251,N_206);
or U561 (N_561,N_250,N_293);
nand U562 (N_562,N_267,In_349);
nor U563 (N_563,In_668,N_204);
nand U564 (N_564,In_610,In_720);
or U565 (N_565,N_275,In_401);
nand U566 (N_566,N_243,N_203);
or U567 (N_567,In_521,N_213);
and U568 (N_568,N_238,N_177);
nand U569 (N_569,N_362,N_334);
and U570 (N_570,N_353,In_336);
or U571 (N_571,N_247,N_339);
and U572 (N_572,In_365,In_456);
nor U573 (N_573,N_297,N_163);
or U574 (N_574,In_84,N_57);
nand U575 (N_575,In_348,N_320);
nor U576 (N_576,N_376,N_393);
and U577 (N_577,N_329,N_308);
nand U578 (N_578,N_205,In_391);
and U579 (N_579,N_154,N_202);
nand U580 (N_580,N_325,N_217);
nor U581 (N_581,In_141,N_374);
nor U582 (N_582,N_66,In_84);
nand U583 (N_583,N_378,In_340);
nor U584 (N_584,In_444,In_144);
nor U585 (N_585,In_348,In_608);
nor U586 (N_586,N_84,In_46);
and U587 (N_587,N_237,In_156);
nand U588 (N_588,In_702,N_363);
and U589 (N_589,N_262,N_29);
nand U590 (N_590,In_301,In_723);
or U591 (N_591,N_148,N_328);
nand U592 (N_592,In_401,N_232);
nor U593 (N_593,N_237,N_151);
nor U594 (N_594,N_399,In_665);
or U595 (N_595,N_276,In_254);
or U596 (N_596,N_240,N_295);
and U597 (N_597,N_270,N_371);
or U598 (N_598,N_340,In_223);
and U599 (N_599,In_531,In_33);
nor U600 (N_600,N_500,N_553);
nor U601 (N_601,N_546,N_496);
xor U602 (N_602,N_490,N_503);
nor U603 (N_603,N_540,N_404);
nand U604 (N_604,N_545,N_477);
and U605 (N_605,N_463,N_589);
nor U606 (N_606,N_572,N_409);
nand U607 (N_607,N_515,N_487);
or U608 (N_608,N_510,N_554);
and U609 (N_609,N_587,N_439);
nand U610 (N_610,N_531,N_432);
and U611 (N_611,N_507,N_414);
or U612 (N_612,N_440,N_529);
or U613 (N_613,N_418,N_449);
and U614 (N_614,N_471,N_468);
and U615 (N_615,N_446,N_465);
or U616 (N_616,N_537,N_481);
nand U617 (N_617,N_528,N_522);
and U618 (N_618,N_413,N_588);
nand U619 (N_619,N_582,N_591);
and U620 (N_620,N_548,N_520);
or U621 (N_621,N_599,N_493);
or U622 (N_622,N_562,N_486);
nor U623 (N_623,N_473,N_451);
or U624 (N_624,N_556,N_488);
and U625 (N_625,N_502,N_571);
and U626 (N_626,N_469,N_585);
and U627 (N_627,N_586,N_530);
or U628 (N_628,N_420,N_443);
xor U629 (N_629,N_547,N_580);
nor U630 (N_630,N_434,N_506);
or U631 (N_631,N_564,N_457);
and U632 (N_632,N_593,N_576);
and U633 (N_633,N_596,N_517);
or U634 (N_634,N_430,N_544);
nor U635 (N_635,N_410,N_559);
and U636 (N_636,N_533,N_565);
or U637 (N_637,N_497,N_532);
nor U638 (N_638,N_460,N_513);
nor U639 (N_639,N_476,N_479);
nor U640 (N_640,N_498,N_508);
or U641 (N_641,N_595,N_436);
and U642 (N_642,N_470,N_442);
nand U643 (N_643,N_594,N_483);
or U644 (N_644,N_577,N_549);
or U645 (N_645,N_592,N_561);
xnor U646 (N_646,N_569,N_485);
or U647 (N_647,N_438,N_521);
or U648 (N_648,N_590,N_407);
and U649 (N_649,N_467,N_459);
xnor U650 (N_650,N_455,N_495);
nand U651 (N_651,N_570,N_504);
and U652 (N_652,N_519,N_447);
xnor U653 (N_653,N_558,N_478);
xor U654 (N_654,N_429,N_505);
xor U655 (N_655,N_482,N_421);
and U656 (N_656,N_491,N_405);
nor U657 (N_657,N_437,N_536);
and U658 (N_658,N_466,N_550);
nor U659 (N_659,N_567,N_575);
nor U660 (N_660,N_492,N_452);
xnor U661 (N_661,N_526,N_484);
nand U662 (N_662,N_597,N_480);
nand U663 (N_663,N_419,N_444);
xor U664 (N_664,N_448,N_598);
nand U665 (N_665,N_415,N_525);
nand U666 (N_666,N_475,N_541);
and U667 (N_667,N_450,N_535);
or U668 (N_668,N_583,N_401);
nor U669 (N_669,N_560,N_453);
nor U670 (N_670,N_555,N_524);
and U671 (N_671,N_581,N_514);
or U672 (N_672,N_563,N_584);
nand U673 (N_673,N_441,N_445);
or U674 (N_674,N_462,N_422);
nand U675 (N_675,N_400,N_557);
nor U676 (N_676,N_494,N_426);
nand U677 (N_677,N_534,N_464);
nor U678 (N_678,N_474,N_417);
xnor U679 (N_679,N_412,N_423);
or U680 (N_680,N_406,N_551);
nand U681 (N_681,N_472,N_552);
or U682 (N_682,N_489,N_425);
nor U683 (N_683,N_458,N_512);
nor U684 (N_684,N_431,N_454);
xnor U685 (N_685,N_566,N_427);
nor U686 (N_686,N_527,N_573);
or U687 (N_687,N_456,N_501);
and U688 (N_688,N_402,N_509);
nor U689 (N_689,N_435,N_416);
xor U690 (N_690,N_574,N_461);
nand U691 (N_691,N_516,N_543);
nand U692 (N_692,N_539,N_428);
nand U693 (N_693,N_424,N_518);
and U694 (N_694,N_499,N_411);
nor U695 (N_695,N_511,N_538);
nand U696 (N_696,N_542,N_408);
nand U697 (N_697,N_568,N_523);
or U698 (N_698,N_403,N_578);
nor U699 (N_699,N_433,N_579);
and U700 (N_700,N_467,N_550);
and U701 (N_701,N_453,N_564);
nor U702 (N_702,N_438,N_422);
xor U703 (N_703,N_501,N_475);
nor U704 (N_704,N_521,N_574);
nor U705 (N_705,N_445,N_555);
or U706 (N_706,N_470,N_559);
or U707 (N_707,N_456,N_582);
nand U708 (N_708,N_463,N_468);
nor U709 (N_709,N_461,N_400);
xor U710 (N_710,N_550,N_529);
nand U711 (N_711,N_417,N_575);
nor U712 (N_712,N_550,N_442);
nor U713 (N_713,N_543,N_525);
nand U714 (N_714,N_412,N_549);
nand U715 (N_715,N_508,N_544);
and U716 (N_716,N_464,N_437);
nand U717 (N_717,N_502,N_435);
and U718 (N_718,N_461,N_580);
nor U719 (N_719,N_454,N_472);
xnor U720 (N_720,N_432,N_446);
nor U721 (N_721,N_568,N_574);
or U722 (N_722,N_549,N_481);
nand U723 (N_723,N_518,N_538);
nand U724 (N_724,N_444,N_429);
nand U725 (N_725,N_588,N_479);
and U726 (N_726,N_540,N_416);
and U727 (N_727,N_467,N_533);
nor U728 (N_728,N_558,N_570);
nand U729 (N_729,N_509,N_549);
nand U730 (N_730,N_459,N_584);
nand U731 (N_731,N_559,N_482);
and U732 (N_732,N_453,N_553);
nor U733 (N_733,N_569,N_512);
or U734 (N_734,N_455,N_577);
nand U735 (N_735,N_458,N_443);
nand U736 (N_736,N_491,N_564);
nand U737 (N_737,N_472,N_521);
nor U738 (N_738,N_566,N_579);
and U739 (N_739,N_413,N_551);
and U740 (N_740,N_532,N_479);
nand U741 (N_741,N_590,N_452);
or U742 (N_742,N_402,N_598);
or U743 (N_743,N_409,N_505);
xor U744 (N_744,N_469,N_588);
nor U745 (N_745,N_438,N_490);
or U746 (N_746,N_504,N_530);
or U747 (N_747,N_409,N_427);
and U748 (N_748,N_489,N_577);
or U749 (N_749,N_457,N_525);
or U750 (N_750,N_409,N_598);
nor U751 (N_751,N_546,N_502);
nand U752 (N_752,N_460,N_591);
nor U753 (N_753,N_462,N_432);
and U754 (N_754,N_512,N_498);
xor U755 (N_755,N_550,N_423);
or U756 (N_756,N_527,N_463);
or U757 (N_757,N_538,N_408);
nand U758 (N_758,N_472,N_560);
nor U759 (N_759,N_564,N_581);
or U760 (N_760,N_416,N_425);
nor U761 (N_761,N_507,N_501);
and U762 (N_762,N_517,N_453);
nand U763 (N_763,N_520,N_536);
nor U764 (N_764,N_568,N_456);
xnor U765 (N_765,N_411,N_402);
nand U766 (N_766,N_578,N_469);
nand U767 (N_767,N_417,N_512);
and U768 (N_768,N_481,N_433);
nor U769 (N_769,N_409,N_420);
xor U770 (N_770,N_509,N_542);
xnor U771 (N_771,N_545,N_547);
and U772 (N_772,N_418,N_487);
and U773 (N_773,N_565,N_488);
nor U774 (N_774,N_588,N_530);
nand U775 (N_775,N_591,N_553);
and U776 (N_776,N_411,N_427);
nor U777 (N_777,N_423,N_564);
or U778 (N_778,N_519,N_457);
or U779 (N_779,N_476,N_407);
nor U780 (N_780,N_572,N_464);
xnor U781 (N_781,N_575,N_409);
nor U782 (N_782,N_426,N_531);
and U783 (N_783,N_501,N_537);
and U784 (N_784,N_424,N_419);
and U785 (N_785,N_465,N_544);
nor U786 (N_786,N_571,N_530);
xor U787 (N_787,N_487,N_520);
and U788 (N_788,N_526,N_400);
nand U789 (N_789,N_530,N_506);
or U790 (N_790,N_453,N_554);
or U791 (N_791,N_562,N_438);
or U792 (N_792,N_565,N_468);
nand U793 (N_793,N_509,N_404);
and U794 (N_794,N_479,N_570);
and U795 (N_795,N_590,N_416);
nand U796 (N_796,N_486,N_480);
nor U797 (N_797,N_494,N_459);
or U798 (N_798,N_456,N_468);
nand U799 (N_799,N_572,N_579);
nand U800 (N_800,N_611,N_615);
nor U801 (N_801,N_664,N_649);
nor U802 (N_802,N_776,N_788);
nand U803 (N_803,N_631,N_627);
nor U804 (N_804,N_687,N_797);
xor U805 (N_805,N_626,N_744);
and U806 (N_806,N_614,N_613);
and U807 (N_807,N_679,N_737);
or U808 (N_808,N_640,N_724);
nand U809 (N_809,N_714,N_655);
or U810 (N_810,N_644,N_790);
nand U811 (N_811,N_602,N_792);
nor U812 (N_812,N_796,N_641);
nor U813 (N_813,N_674,N_675);
nand U814 (N_814,N_717,N_771);
nand U815 (N_815,N_783,N_617);
and U816 (N_816,N_745,N_632);
or U817 (N_817,N_688,N_630);
or U818 (N_818,N_736,N_731);
nor U819 (N_819,N_622,N_703);
and U820 (N_820,N_657,N_713);
and U821 (N_821,N_633,N_734);
or U822 (N_822,N_682,N_693);
nor U823 (N_823,N_738,N_639);
nor U824 (N_824,N_642,N_695);
or U825 (N_825,N_667,N_718);
nand U826 (N_826,N_634,N_780);
nand U827 (N_827,N_681,N_707);
nor U828 (N_828,N_750,N_685);
nand U829 (N_829,N_747,N_710);
or U830 (N_830,N_794,N_658);
or U831 (N_831,N_648,N_786);
nand U832 (N_832,N_752,N_726);
nand U833 (N_833,N_689,N_694);
and U834 (N_834,N_765,N_696);
and U835 (N_835,N_720,N_697);
or U836 (N_836,N_704,N_635);
nand U837 (N_837,N_767,N_764);
nand U838 (N_838,N_663,N_773);
and U839 (N_839,N_768,N_661);
and U840 (N_840,N_690,N_761);
nor U841 (N_841,N_741,N_754);
or U842 (N_842,N_763,N_743);
or U843 (N_843,N_733,N_722);
nor U844 (N_844,N_723,N_643);
or U845 (N_845,N_730,N_612);
and U846 (N_846,N_715,N_691);
nand U847 (N_847,N_711,N_683);
nor U848 (N_848,N_636,N_610);
and U849 (N_849,N_719,N_660);
and U850 (N_850,N_784,N_787);
or U851 (N_851,N_653,N_621);
xnor U852 (N_852,N_753,N_620);
and U853 (N_853,N_791,N_705);
nand U854 (N_854,N_605,N_651);
and U855 (N_855,N_650,N_646);
and U856 (N_856,N_762,N_662);
nor U857 (N_857,N_680,N_647);
or U858 (N_858,N_729,N_686);
and U859 (N_859,N_795,N_725);
nor U860 (N_860,N_672,N_619);
nor U861 (N_861,N_669,N_656);
or U862 (N_862,N_668,N_769);
nor U863 (N_863,N_751,N_666);
or U864 (N_864,N_727,N_676);
or U865 (N_865,N_757,N_637);
and U866 (N_866,N_766,N_606);
and U867 (N_867,N_673,N_789);
nand U868 (N_868,N_645,N_735);
nand U869 (N_869,N_659,N_774);
nand U870 (N_870,N_748,N_770);
and U871 (N_871,N_625,N_624);
xnor U872 (N_872,N_758,N_712);
or U873 (N_873,N_609,N_742);
or U874 (N_874,N_706,N_785);
or U875 (N_875,N_670,N_708);
nand U876 (N_876,N_608,N_671);
nor U877 (N_877,N_755,N_778);
or U878 (N_878,N_775,N_604);
nor U879 (N_879,N_777,N_760);
nand U880 (N_880,N_793,N_749);
xor U881 (N_881,N_799,N_699);
nor U882 (N_882,N_603,N_652);
and U883 (N_883,N_772,N_702);
nand U884 (N_884,N_779,N_759);
nand U885 (N_885,N_798,N_623);
or U886 (N_886,N_746,N_756);
xnor U887 (N_887,N_739,N_684);
xor U888 (N_888,N_740,N_728);
xor U889 (N_889,N_628,N_692);
xor U890 (N_890,N_701,N_600);
nand U891 (N_891,N_654,N_629);
nor U892 (N_892,N_698,N_607);
xnor U893 (N_893,N_618,N_732);
nand U894 (N_894,N_616,N_677);
nand U895 (N_895,N_782,N_678);
nor U896 (N_896,N_665,N_638);
and U897 (N_897,N_601,N_781);
nand U898 (N_898,N_716,N_700);
nor U899 (N_899,N_721,N_709);
nand U900 (N_900,N_705,N_600);
nor U901 (N_901,N_667,N_648);
nor U902 (N_902,N_628,N_637);
nor U903 (N_903,N_632,N_797);
and U904 (N_904,N_601,N_611);
and U905 (N_905,N_660,N_680);
or U906 (N_906,N_729,N_664);
nor U907 (N_907,N_772,N_701);
and U908 (N_908,N_680,N_650);
nor U909 (N_909,N_695,N_630);
xnor U910 (N_910,N_689,N_786);
or U911 (N_911,N_661,N_655);
nand U912 (N_912,N_788,N_622);
or U913 (N_913,N_764,N_717);
or U914 (N_914,N_699,N_640);
or U915 (N_915,N_682,N_744);
nand U916 (N_916,N_648,N_761);
nand U917 (N_917,N_792,N_678);
nand U918 (N_918,N_641,N_798);
and U919 (N_919,N_790,N_712);
nor U920 (N_920,N_600,N_650);
nor U921 (N_921,N_699,N_674);
nand U922 (N_922,N_662,N_688);
xnor U923 (N_923,N_694,N_782);
nand U924 (N_924,N_786,N_700);
nor U925 (N_925,N_761,N_722);
xor U926 (N_926,N_760,N_654);
nor U927 (N_927,N_795,N_713);
xor U928 (N_928,N_765,N_642);
nor U929 (N_929,N_680,N_722);
xor U930 (N_930,N_744,N_646);
or U931 (N_931,N_699,N_660);
and U932 (N_932,N_664,N_717);
nand U933 (N_933,N_773,N_751);
and U934 (N_934,N_620,N_679);
and U935 (N_935,N_638,N_713);
xor U936 (N_936,N_693,N_672);
nand U937 (N_937,N_654,N_750);
nand U938 (N_938,N_604,N_614);
or U939 (N_939,N_703,N_696);
nor U940 (N_940,N_637,N_759);
nand U941 (N_941,N_635,N_642);
nor U942 (N_942,N_646,N_690);
or U943 (N_943,N_763,N_707);
xnor U944 (N_944,N_720,N_616);
or U945 (N_945,N_623,N_780);
xnor U946 (N_946,N_793,N_747);
nor U947 (N_947,N_610,N_723);
or U948 (N_948,N_739,N_610);
nor U949 (N_949,N_611,N_671);
nor U950 (N_950,N_681,N_729);
or U951 (N_951,N_651,N_617);
or U952 (N_952,N_600,N_694);
nand U953 (N_953,N_715,N_740);
nand U954 (N_954,N_602,N_656);
xnor U955 (N_955,N_680,N_795);
nand U956 (N_956,N_751,N_730);
nand U957 (N_957,N_752,N_730);
and U958 (N_958,N_684,N_666);
and U959 (N_959,N_761,N_645);
nor U960 (N_960,N_701,N_679);
and U961 (N_961,N_671,N_653);
and U962 (N_962,N_741,N_689);
nand U963 (N_963,N_639,N_634);
xor U964 (N_964,N_752,N_661);
nor U965 (N_965,N_666,N_725);
xor U966 (N_966,N_640,N_645);
xor U967 (N_967,N_607,N_673);
nor U968 (N_968,N_647,N_642);
nand U969 (N_969,N_613,N_780);
and U970 (N_970,N_685,N_680);
nor U971 (N_971,N_632,N_773);
nor U972 (N_972,N_792,N_723);
nand U973 (N_973,N_698,N_603);
nor U974 (N_974,N_625,N_648);
and U975 (N_975,N_620,N_628);
nand U976 (N_976,N_773,N_630);
or U977 (N_977,N_717,N_660);
nor U978 (N_978,N_790,N_643);
nand U979 (N_979,N_788,N_666);
nor U980 (N_980,N_751,N_757);
nor U981 (N_981,N_695,N_714);
nand U982 (N_982,N_773,N_703);
or U983 (N_983,N_674,N_694);
and U984 (N_984,N_624,N_701);
nor U985 (N_985,N_781,N_665);
and U986 (N_986,N_741,N_777);
nand U987 (N_987,N_758,N_795);
nand U988 (N_988,N_658,N_743);
nor U989 (N_989,N_790,N_659);
or U990 (N_990,N_614,N_617);
or U991 (N_991,N_764,N_637);
nor U992 (N_992,N_785,N_633);
xor U993 (N_993,N_716,N_701);
nor U994 (N_994,N_710,N_621);
and U995 (N_995,N_758,N_663);
nor U996 (N_996,N_659,N_699);
xor U997 (N_997,N_620,N_768);
and U998 (N_998,N_693,N_655);
xor U999 (N_999,N_652,N_674);
and U1000 (N_1000,N_822,N_999);
nor U1001 (N_1001,N_904,N_863);
or U1002 (N_1002,N_973,N_819);
and U1003 (N_1003,N_919,N_853);
and U1004 (N_1004,N_933,N_800);
nor U1005 (N_1005,N_900,N_955);
nand U1006 (N_1006,N_865,N_880);
and U1007 (N_1007,N_814,N_855);
nor U1008 (N_1008,N_846,N_917);
nor U1009 (N_1009,N_958,N_913);
and U1010 (N_1010,N_927,N_931);
xor U1011 (N_1011,N_861,N_829);
and U1012 (N_1012,N_983,N_964);
nor U1013 (N_1013,N_912,N_802);
and U1014 (N_1014,N_862,N_936);
nand U1015 (N_1015,N_868,N_804);
or U1016 (N_1016,N_997,N_873);
or U1017 (N_1017,N_911,N_872);
nand U1018 (N_1018,N_961,N_925);
nor U1019 (N_1019,N_817,N_810);
nor U1020 (N_1020,N_920,N_987);
or U1021 (N_1021,N_808,N_847);
and U1022 (N_1022,N_956,N_989);
or U1023 (N_1023,N_949,N_940);
xnor U1024 (N_1024,N_918,N_969);
or U1025 (N_1025,N_996,N_926);
nand U1026 (N_1026,N_893,N_851);
and U1027 (N_1027,N_994,N_903);
or U1028 (N_1028,N_857,N_944);
nand U1029 (N_1029,N_859,N_952);
or U1030 (N_1030,N_992,N_890);
nor U1031 (N_1031,N_897,N_832);
nor U1032 (N_1032,N_824,N_909);
or U1033 (N_1033,N_977,N_905);
nand U1034 (N_1034,N_823,N_833);
and U1035 (N_1035,N_948,N_801);
nor U1036 (N_1036,N_976,N_877);
nor U1037 (N_1037,N_916,N_886);
nand U1038 (N_1038,N_881,N_838);
nor U1039 (N_1039,N_860,N_806);
or U1040 (N_1040,N_813,N_840);
and U1041 (N_1041,N_842,N_929);
nor U1042 (N_1042,N_889,N_878);
and U1043 (N_1043,N_899,N_907);
or U1044 (N_1044,N_891,N_951);
and U1045 (N_1045,N_981,N_980);
nor U1046 (N_1046,N_979,N_852);
and U1047 (N_1047,N_908,N_963);
nand U1048 (N_1048,N_836,N_923);
or U1049 (N_1049,N_970,N_978);
nor U1050 (N_1050,N_953,N_870);
nor U1051 (N_1051,N_898,N_990);
nand U1052 (N_1052,N_820,N_812);
and U1053 (N_1053,N_966,N_837);
and U1054 (N_1054,N_867,N_968);
and U1055 (N_1055,N_883,N_835);
nand U1056 (N_1056,N_942,N_941);
nand U1057 (N_1057,N_938,N_975);
and U1058 (N_1058,N_845,N_807);
or U1059 (N_1059,N_910,N_848);
or U1060 (N_1060,N_945,N_932);
nand U1061 (N_1061,N_960,N_943);
or U1062 (N_1062,N_827,N_830);
or U1063 (N_1063,N_995,N_962);
or U1064 (N_1064,N_871,N_864);
nor U1065 (N_1065,N_826,N_869);
and U1066 (N_1066,N_998,N_831);
and U1067 (N_1067,N_858,N_825);
or U1068 (N_1068,N_967,N_985);
nand U1069 (N_1069,N_876,N_984);
and U1070 (N_1070,N_950,N_834);
or U1071 (N_1071,N_888,N_982);
and U1072 (N_1072,N_841,N_988);
and U1073 (N_1073,N_971,N_896);
nor U1074 (N_1074,N_914,N_928);
or U1075 (N_1075,N_875,N_843);
or U1076 (N_1076,N_991,N_887);
nor U1077 (N_1077,N_986,N_821);
nor U1078 (N_1078,N_818,N_906);
and U1079 (N_1079,N_902,N_828);
or U1080 (N_1080,N_965,N_922);
and U1081 (N_1081,N_885,N_805);
xor U1082 (N_1082,N_946,N_895);
nor U1083 (N_1083,N_957,N_882);
or U1084 (N_1084,N_839,N_879);
nor U1085 (N_1085,N_901,N_856);
nor U1086 (N_1086,N_935,N_947);
xnor U1087 (N_1087,N_803,N_866);
and U1088 (N_1088,N_816,N_972);
and U1089 (N_1089,N_939,N_934);
or U1090 (N_1090,N_930,N_915);
xor U1091 (N_1091,N_993,N_894);
nand U1092 (N_1092,N_809,N_850);
and U1093 (N_1093,N_921,N_811);
nand U1094 (N_1094,N_892,N_854);
nand U1095 (N_1095,N_844,N_849);
xor U1096 (N_1096,N_924,N_959);
nor U1097 (N_1097,N_974,N_937);
and U1098 (N_1098,N_874,N_954);
xnor U1099 (N_1099,N_884,N_815);
xnor U1100 (N_1100,N_989,N_965);
nand U1101 (N_1101,N_853,N_959);
xnor U1102 (N_1102,N_850,N_879);
and U1103 (N_1103,N_903,N_909);
nand U1104 (N_1104,N_978,N_982);
and U1105 (N_1105,N_846,N_952);
or U1106 (N_1106,N_839,N_830);
and U1107 (N_1107,N_850,N_992);
or U1108 (N_1108,N_919,N_993);
nand U1109 (N_1109,N_992,N_857);
nor U1110 (N_1110,N_909,N_813);
nand U1111 (N_1111,N_906,N_952);
nor U1112 (N_1112,N_837,N_877);
or U1113 (N_1113,N_983,N_961);
nand U1114 (N_1114,N_913,N_850);
and U1115 (N_1115,N_875,N_985);
nor U1116 (N_1116,N_804,N_927);
nand U1117 (N_1117,N_901,N_859);
or U1118 (N_1118,N_898,N_809);
nand U1119 (N_1119,N_865,N_967);
nor U1120 (N_1120,N_854,N_890);
nor U1121 (N_1121,N_827,N_962);
nor U1122 (N_1122,N_959,N_813);
and U1123 (N_1123,N_904,N_945);
nand U1124 (N_1124,N_825,N_873);
nand U1125 (N_1125,N_884,N_869);
xor U1126 (N_1126,N_981,N_899);
nor U1127 (N_1127,N_859,N_830);
xnor U1128 (N_1128,N_881,N_807);
or U1129 (N_1129,N_908,N_907);
nand U1130 (N_1130,N_931,N_989);
nand U1131 (N_1131,N_922,N_964);
and U1132 (N_1132,N_924,N_984);
and U1133 (N_1133,N_942,N_888);
and U1134 (N_1134,N_998,N_991);
and U1135 (N_1135,N_800,N_870);
nand U1136 (N_1136,N_930,N_816);
or U1137 (N_1137,N_964,N_903);
or U1138 (N_1138,N_825,N_965);
nand U1139 (N_1139,N_984,N_820);
nand U1140 (N_1140,N_997,N_838);
and U1141 (N_1141,N_852,N_970);
nand U1142 (N_1142,N_970,N_932);
or U1143 (N_1143,N_997,N_968);
and U1144 (N_1144,N_940,N_855);
nand U1145 (N_1145,N_997,N_912);
nand U1146 (N_1146,N_919,N_880);
or U1147 (N_1147,N_993,N_965);
nand U1148 (N_1148,N_972,N_906);
and U1149 (N_1149,N_965,N_808);
and U1150 (N_1150,N_806,N_851);
and U1151 (N_1151,N_929,N_910);
nand U1152 (N_1152,N_892,N_959);
nand U1153 (N_1153,N_813,N_873);
and U1154 (N_1154,N_955,N_928);
and U1155 (N_1155,N_850,N_934);
xnor U1156 (N_1156,N_907,N_946);
and U1157 (N_1157,N_899,N_974);
xor U1158 (N_1158,N_869,N_827);
and U1159 (N_1159,N_970,N_986);
nor U1160 (N_1160,N_905,N_926);
or U1161 (N_1161,N_847,N_889);
nand U1162 (N_1162,N_895,N_825);
nand U1163 (N_1163,N_965,N_830);
and U1164 (N_1164,N_809,N_968);
and U1165 (N_1165,N_991,N_800);
xor U1166 (N_1166,N_906,N_916);
nand U1167 (N_1167,N_834,N_994);
and U1168 (N_1168,N_934,N_883);
nand U1169 (N_1169,N_990,N_959);
nand U1170 (N_1170,N_872,N_965);
nand U1171 (N_1171,N_829,N_805);
and U1172 (N_1172,N_832,N_911);
nor U1173 (N_1173,N_903,N_938);
nor U1174 (N_1174,N_838,N_829);
or U1175 (N_1175,N_832,N_915);
and U1176 (N_1176,N_888,N_948);
or U1177 (N_1177,N_839,N_818);
xor U1178 (N_1178,N_881,N_889);
and U1179 (N_1179,N_988,N_888);
or U1180 (N_1180,N_966,N_825);
nand U1181 (N_1181,N_818,N_895);
or U1182 (N_1182,N_908,N_993);
or U1183 (N_1183,N_895,N_964);
and U1184 (N_1184,N_823,N_969);
nor U1185 (N_1185,N_941,N_906);
or U1186 (N_1186,N_843,N_894);
xor U1187 (N_1187,N_973,N_800);
nor U1188 (N_1188,N_905,N_911);
and U1189 (N_1189,N_920,N_901);
nand U1190 (N_1190,N_933,N_924);
or U1191 (N_1191,N_944,N_964);
and U1192 (N_1192,N_833,N_824);
and U1193 (N_1193,N_977,N_882);
or U1194 (N_1194,N_809,N_965);
xnor U1195 (N_1195,N_990,N_984);
nor U1196 (N_1196,N_961,N_844);
nand U1197 (N_1197,N_812,N_998);
nand U1198 (N_1198,N_971,N_911);
nand U1199 (N_1199,N_880,N_828);
or U1200 (N_1200,N_1103,N_1108);
or U1201 (N_1201,N_1088,N_1020);
nand U1202 (N_1202,N_1069,N_1021);
and U1203 (N_1203,N_1162,N_1083);
nor U1204 (N_1204,N_1125,N_1074);
nand U1205 (N_1205,N_1077,N_1024);
xnor U1206 (N_1206,N_1100,N_1138);
and U1207 (N_1207,N_1019,N_1065);
and U1208 (N_1208,N_1160,N_1058);
nand U1209 (N_1209,N_1163,N_1196);
or U1210 (N_1210,N_1165,N_1041);
nor U1211 (N_1211,N_1174,N_1142);
nor U1212 (N_1212,N_1008,N_1164);
or U1213 (N_1213,N_1183,N_1158);
nand U1214 (N_1214,N_1107,N_1050);
or U1215 (N_1215,N_1151,N_1131);
nor U1216 (N_1216,N_1113,N_1124);
and U1217 (N_1217,N_1015,N_1182);
nand U1218 (N_1218,N_1156,N_1010);
nor U1219 (N_1219,N_1187,N_1054);
nand U1220 (N_1220,N_1052,N_1130);
or U1221 (N_1221,N_1102,N_1153);
nand U1222 (N_1222,N_1172,N_1161);
or U1223 (N_1223,N_1176,N_1134);
xor U1224 (N_1224,N_1034,N_1147);
and U1225 (N_1225,N_1048,N_1145);
or U1226 (N_1226,N_1188,N_1004);
and U1227 (N_1227,N_1005,N_1013);
or U1228 (N_1228,N_1144,N_1146);
and U1229 (N_1229,N_1002,N_1136);
and U1230 (N_1230,N_1043,N_1132);
nand U1231 (N_1231,N_1084,N_1149);
nor U1232 (N_1232,N_1126,N_1189);
nand U1233 (N_1233,N_1135,N_1011);
and U1234 (N_1234,N_1025,N_1195);
nor U1235 (N_1235,N_1090,N_1167);
xor U1236 (N_1236,N_1118,N_1028);
nand U1237 (N_1237,N_1092,N_1110);
nand U1238 (N_1238,N_1022,N_1046);
nand U1239 (N_1239,N_1141,N_1061);
nor U1240 (N_1240,N_1119,N_1129);
and U1241 (N_1241,N_1199,N_1044);
nor U1242 (N_1242,N_1040,N_1081);
nor U1243 (N_1243,N_1097,N_1063);
and U1244 (N_1244,N_1076,N_1185);
nand U1245 (N_1245,N_1059,N_1042);
nand U1246 (N_1246,N_1095,N_1012);
nor U1247 (N_1247,N_1049,N_1093);
and U1248 (N_1248,N_1073,N_1056);
and U1249 (N_1249,N_1062,N_1036);
or U1250 (N_1250,N_1137,N_1009);
xnor U1251 (N_1251,N_1027,N_1068);
and U1252 (N_1252,N_1033,N_1096);
and U1253 (N_1253,N_1169,N_1079);
nand U1254 (N_1254,N_1099,N_1091);
or U1255 (N_1255,N_1072,N_1121);
nor U1256 (N_1256,N_1112,N_1152);
and U1257 (N_1257,N_1031,N_1191);
xnor U1258 (N_1258,N_1085,N_1150);
nor U1259 (N_1259,N_1111,N_1197);
nor U1260 (N_1260,N_1066,N_1157);
nand U1261 (N_1261,N_1087,N_1171);
xnor U1262 (N_1262,N_1082,N_1177);
or U1263 (N_1263,N_1045,N_1123);
nor U1264 (N_1264,N_1003,N_1078);
or U1265 (N_1265,N_1098,N_1181);
nor U1266 (N_1266,N_1075,N_1117);
nor U1267 (N_1267,N_1140,N_1198);
and U1268 (N_1268,N_1047,N_1070);
nand U1269 (N_1269,N_1071,N_1001);
or U1270 (N_1270,N_1175,N_1039);
or U1271 (N_1271,N_1037,N_1105);
and U1272 (N_1272,N_1128,N_1067);
and U1273 (N_1273,N_1026,N_1032);
and U1274 (N_1274,N_1064,N_1192);
or U1275 (N_1275,N_1116,N_1170);
nand U1276 (N_1276,N_1122,N_1055);
or U1277 (N_1277,N_1120,N_1057);
xnor U1278 (N_1278,N_1179,N_1060);
nor U1279 (N_1279,N_1133,N_1109);
xor U1280 (N_1280,N_1030,N_1173);
or U1281 (N_1281,N_1006,N_1094);
nor U1282 (N_1282,N_1086,N_1029);
nand U1283 (N_1283,N_1114,N_1080);
nor U1284 (N_1284,N_1155,N_1180);
nand U1285 (N_1285,N_1014,N_1053);
or U1286 (N_1286,N_1007,N_1193);
nand U1287 (N_1287,N_1184,N_1154);
or U1288 (N_1288,N_1186,N_1143);
nand U1289 (N_1289,N_1089,N_1035);
nor U1290 (N_1290,N_1106,N_1166);
or U1291 (N_1291,N_1104,N_1139);
and U1292 (N_1292,N_1159,N_1101);
or U1293 (N_1293,N_1023,N_1178);
nand U1294 (N_1294,N_1194,N_1168);
xnor U1295 (N_1295,N_1127,N_1016);
or U1296 (N_1296,N_1018,N_1000);
and U1297 (N_1297,N_1148,N_1190);
nor U1298 (N_1298,N_1051,N_1115);
nor U1299 (N_1299,N_1017,N_1038);
xnor U1300 (N_1300,N_1015,N_1086);
nand U1301 (N_1301,N_1028,N_1083);
or U1302 (N_1302,N_1167,N_1132);
nand U1303 (N_1303,N_1151,N_1099);
or U1304 (N_1304,N_1147,N_1021);
or U1305 (N_1305,N_1032,N_1056);
and U1306 (N_1306,N_1115,N_1074);
nand U1307 (N_1307,N_1014,N_1102);
and U1308 (N_1308,N_1006,N_1038);
and U1309 (N_1309,N_1125,N_1121);
and U1310 (N_1310,N_1042,N_1152);
and U1311 (N_1311,N_1112,N_1106);
nor U1312 (N_1312,N_1156,N_1102);
and U1313 (N_1313,N_1002,N_1020);
and U1314 (N_1314,N_1165,N_1034);
nand U1315 (N_1315,N_1107,N_1174);
nand U1316 (N_1316,N_1199,N_1047);
nand U1317 (N_1317,N_1140,N_1097);
nand U1318 (N_1318,N_1121,N_1099);
and U1319 (N_1319,N_1014,N_1147);
or U1320 (N_1320,N_1137,N_1139);
nor U1321 (N_1321,N_1076,N_1094);
or U1322 (N_1322,N_1184,N_1192);
or U1323 (N_1323,N_1103,N_1188);
nand U1324 (N_1324,N_1113,N_1033);
nand U1325 (N_1325,N_1037,N_1124);
nand U1326 (N_1326,N_1054,N_1163);
xor U1327 (N_1327,N_1173,N_1048);
nor U1328 (N_1328,N_1142,N_1027);
nand U1329 (N_1329,N_1048,N_1036);
or U1330 (N_1330,N_1065,N_1126);
and U1331 (N_1331,N_1198,N_1138);
nand U1332 (N_1332,N_1012,N_1060);
and U1333 (N_1333,N_1045,N_1138);
nand U1334 (N_1334,N_1037,N_1169);
nand U1335 (N_1335,N_1007,N_1183);
nand U1336 (N_1336,N_1057,N_1081);
or U1337 (N_1337,N_1087,N_1117);
and U1338 (N_1338,N_1020,N_1057);
nor U1339 (N_1339,N_1187,N_1155);
or U1340 (N_1340,N_1010,N_1124);
nand U1341 (N_1341,N_1168,N_1012);
or U1342 (N_1342,N_1057,N_1121);
and U1343 (N_1343,N_1123,N_1043);
and U1344 (N_1344,N_1145,N_1122);
nor U1345 (N_1345,N_1048,N_1007);
or U1346 (N_1346,N_1197,N_1091);
or U1347 (N_1347,N_1098,N_1065);
nor U1348 (N_1348,N_1146,N_1019);
or U1349 (N_1349,N_1174,N_1115);
and U1350 (N_1350,N_1151,N_1089);
nand U1351 (N_1351,N_1173,N_1077);
nor U1352 (N_1352,N_1015,N_1057);
nor U1353 (N_1353,N_1065,N_1079);
xnor U1354 (N_1354,N_1100,N_1026);
or U1355 (N_1355,N_1165,N_1028);
and U1356 (N_1356,N_1083,N_1115);
nor U1357 (N_1357,N_1087,N_1156);
nand U1358 (N_1358,N_1065,N_1035);
xor U1359 (N_1359,N_1031,N_1162);
nor U1360 (N_1360,N_1054,N_1150);
and U1361 (N_1361,N_1047,N_1105);
and U1362 (N_1362,N_1137,N_1072);
nor U1363 (N_1363,N_1154,N_1077);
nor U1364 (N_1364,N_1099,N_1079);
xor U1365 (N_1365,N_1176,N_1054);
nor U1366 (N_1366,N_1036,N_1186);
nand U1367 (N_1367,N_1142,N_1053);
nand U1368 (N_1368,N_1132,N_1045);
nand U1369 (N_1369,N_1063,N_1032);
nor U1370 (N_1370,N_1125,N_1153);
or U1371 (N_1371,N_1019,N_1002);
and U1372 (N_1372,N_1167,N_1114);
nand U1373 (N_1373,N_1064,N_1130);
xnor U1374 (N_1374,N_1070,N_1120);
or U1375 (N_1375,N_1030,N_1075);
and U1376 (N_1376,N_1139,N_1189);
nand U1377 (N_1377,N_1035,N_1036);
nor U1378 (N_1378,N_1196,N_1038);
nand U1379 (N_1379,N_1158,N_1190);
nor U1380 (N_1380,N_1037,N_1015);
nor U1381 (N_1381,N_1089,N_1023);
nand U1382 (N_1382,N_1184,N_1144);
or U1383 (N_1383,N_1187,N_1115);
xnor U1384 (N_1384,N_1000,N_1138);
or U1385 (N_1385,N_1133,N_1047);
or U1386 (N_1386,N_1053,N_1190);
nor U1387 (N_1387,N_1079,N_1183);
nand U1388 (N_1388,N_1005,N_1017);
and U1389 (N_1389,N_1070,N_1051);
nor U1390 (N_1390,N_1034,N_1020);
xor U1391 (N_1391,N_1177,N_1106);
and U1392 (N_1392,N_1193,N_1048);
and U1393 (N_1393,N_1013,N_1117);
or U1394 (N_1394,N_1178,N_1196);
xnor U1395 (N_1395,N_1153,N_1158);
and U1396 (N_1396,N_1106,N_1095);
nand U1397 (N_1397,N_1065,N_1089);
and U1398 (N_1398,N_1013,N_1093);
or U1399 (N_1399,N_1087,N_1013);
or U1400 (N_1400,N_1287,N_1328);
nand U1401 (N_1401,N_1395,N_1249);
or U1402 (N_1402,N_1312,N_1303);
or U1403 (N_1403,N_1238,N_1335);
or U1404 (N_1404,N_1280,N_1291);
or U1405 (N_1405,N_1355,N_1290);
xor U1406 (N_1406,N_1208,N_1219);
or U1407 (N_1407,N_1326,N_1314);
nor U1408 (N_1408,N_1285,N_1396);
and U1409 (N_1409,N_1352,N_1206);
and U1410 (N_1410,N_1286,N_1365);
nor U1411 (N_1411,N_1321,N_1283);
nand U1412 (N_1412,N_1348,N_1227);
xor U1413 (N_1413,N_1292,N_1302);
nor U1414 (N_1414,N_1251,N_1381);
nor U1415 (N_1415,N_1214,N_1334);
or U1416 (N_1416,N_1235,N_1250);
or U1417 (N_1417,N_1261,N_1360);
nor U1418 (N_1418,N_1324,N_1388);
and U1419 (N_1419,N_1346,N_1277);
nand U1420 (N_1420,N_1358,N_1268);
and U1421 (N_1421,N_1203,N_1323);
and U1422 (N_1422,N_1382,N_1344);
or U1423 (N_1423,N_1310,N_1308);
nand U1424 (N_1424,N_1253,N_1317);
nand U1425 (N_1425,N_1289,N_1376);
xor U1426 (N_1426,N_1378,N_1271);
or U1427 (N_1427,N_1331,N_1299);
and U1428 (N_1428,N_1359,N_1304);
nand U1429 (N_1429,N_1370,N_1345);
and U1430 (N_1430,N_1240,N_1263);
or U1431 (N_1431,N_1246,N_1297);
xnor U1432 (N_1432,N_1274,N_1296);
nor U1433 (N_1433,N_1354,N_1315);
and U1434 (N_1434,N_1230,N_1397);
nor U1435 (N_1435,N_1392,N_1247);
nand U1436 (N_1436,N_1260,N_1200);
xnor U1437 (N_1437,N_1361,N_1364);
nand U1438 (N_1438,N_1273,N_1363);
nand U1439 (N_1439,N_1337,N_1351);
nand U1440 (N_1440,N_1207,N_1209);
and U1441 (N_1441,N_1325,N_1272);
or U1442 (N_1442,N_1243,N_1329);
and U1443 (N_1443,N_1236,N_1225);
or U1444 (N_1444,N_1254,N_1343);
nand U1445 (N_1445,N_1228,N_1309);
nor U1446 (N_1446,N_1245,N_1284);
and U1447 (N_1447,N_1327,N_1362);
or U1448 (N_1448,N_1300,N_1233);
and U1449 (N_1449,N_1257,N_1269);
or U1450 (N_1450,N_1281,N_1379);
xnor U1451 (N_1451,N_1390,N_1305);
and U1452 (N_1452,N_1385,N_1342);
nor U1453 (N_1453,N_1393,N_1226);
and U1454 (N_1454,N_1377,N_1347);
or U1455 (N_1455,N_1231,N_1239);
and U1456 (N_1456,N_1366,N_1311);
or U1457 (N_1457,N_1237,N_1212);
nand U1458 (N_1458,N_1298,N_1338);
nand U1459 (N_1459,N_1202,N_1232);
and U1460 (N_1460,N_1371,N_1341);
or U1461 (N_1461,N_1234,N_1295);
nand U1462 (N_1462,N_1332,N_1220);
and U1463 (N_1463,N_1389,N_1213);
and U1464 (N_1464,N_1391,N_1221);
nand U1465 (N_1465,N_1340,N_1244);
and U1466 (N_1466,N_1383,N_1375);
nor U1467 (N_1467,N_1380,N_1216);
nor U1468 (N_1468,N_1356,N_1357);
nand U1469 (N_1469,N_1386,N_1204);
and U1470 (N_1470,N_1222,N_1294);
or U1471 (N_1471,N_1278,N_1248);
nor U1472 (N_1472,N_1374,N_1384);
or U1473 (N_1473,N_1394,N_1293);
or U1474 (N_1474,N_1282,N_1320);
or U1475 (N_1475,N_1242,N_1398);
xor U1476 (N_1476,N_1256,N_1372);
or U1477 (N_1477,N_1399,N_1223);
or U1478 (N_1478,N_1210,N_1313);
nand U1479 (N_1479,N_1264,N_1288);
xor U1480 (N_1480,N_1333,N_1275);
nor U1481 (N_1481,N_1316,N_1339);
nor U1482 (N_1482,N_1276,N_1217);
nor U1483 (N_1483,N_1307,N_1319);
nand U1484 (N_1484,N_1258,N_1215);
nand U1485 (N_1485,N_1205,N_1279);
nor U1486 (N_1486,N_1336,N_1229);
and U1487 (N_1487,N_1373,N_1224);
nand U1488 (N_1488,N_1218,N_1201);
or U1489 (N_1489,N_1318,N_1265);
nor U1490 (N_1490,N_1306,N_1259);
xor U1491 (N_1491,N_1255,N_1349);
and U1492 (N_1492,N_1322,N_1368);
nand U1493 (N_1493,N_1301,N_1350);
or U1494 (N_1494,N_1387,N_1266);
nor U1495 (N_1495,N_1367,N_1262);
and U1496 (N_1496,N_1241,N_1267);
xnor U1497 (N_1497,N_1270,N_1252);
and U1498 (N_1498,N_1330,N_1211);
and U1499 (N_1499,N_1369,N_1353);
nor U1500 (N_1500,N_1381,N_1282);
or U1501 (N_1501,N_1370,N_1303);
or U1502 (N_1502,N_1358,N_1262);
or U1503 (N_1503,N_1282,N_1342);
or U1504 (N_1504,N_1312,N_1324);
and U1505 (N_1505,N_1314,N_1298);
nand U1506 (N_1506,N_1385,N_1231);
nor U1507 (N_1507,N_1358,N_1290);
or U1508 (N_1508,N_1356,N_1297);
nand U1509 (N_1509,N_1274,N_1358);
and U1510 (N_1510,N_1346,N_1294);
nand U1511 (N_1511,N_1305,N_1287);
xnor U1512 (N_1512,N_1307,N_1247);
or U1513 (N_1513,N_1270,N_1248);
xor U1514 (N_1514,N_1373,N_1380);
and U1515 (N_1515,N_1262,N_1321);
nor U1516 (N_1516,N_1377,N_1386);
nand U1517 (N_1517,N_1228,N_1340);
nor U1518 (N_1518,N_1328,N_1215);
and U1519 (N_1519,N_1249,N_1285);
nor U1520 (N_1520,N_1356,N_1295);
or U1521 (N_1521,N_1339,N_1237);
nor U1522 (N_1522,N_1202,N_1288);
nor U1523 (N_1523,N_1329,N_1374);
nand U1524 (N_1524,N_1219,N_1356);
nand U1525 (N_1525,N_1209,N_1247);
and U1526 (N_1526,N_1244,N_1330);
or U1527 (N_1527,N_1371,N_1348);
and U1528 (N_1528,N_1282,N_1287);
and U1529 (N_1529,N_1384,N_1341);
and U1530 (N_1530,N_1373,N_1382);
nand U1531 (N_1531,N_1290,N_1250);
nor U1532 (N_1532,N_1363,N_1362);
nand U1533 (N_1533,N_1304,N_1321);
and U1534 (N_1534,N_1386,N_1270);
and U1535 (N_1535,N_1364,N_1210);
xnor U1536 (N_1536,N_1310,N_1269);
or U1537 (N_1537,N_1393,N_1298);
nand U1538 (N_1538,N_1310,N_1335);
nand U1539 (N_1539,N_1381,N_1360);
and U1540 (N_1540,N_1385,N_1305);
nand U1541 (N_1541,N_1231,N_1399);
nor U1542 (N_1542,N_1350,N_1333);
or U1543 (N_1543,N_1286,N_1392);
nand U1544 (N_1544,N_1332,N_1249);
and U1545 (N_1545,N_1344,N_1331);
and U1546 (N_1546,N_1255,N_1245);
xnor U1547 (N_1547,N_1343,N_1349);
and U1548 (N_1548,N_1217,N_1229);
or U1549 (N_1549,N_1351,N_1215);
or U1550 (N_1550,N_1325,N_1227);
nor U1551 (N_1551,N_1321,N_1367);
or U1552 (N_1552,N_1234,N_1229);
nand U1553 (N_1553,N_1392,N_1356);
nand U1554 (N_1554,N_1251,N_1241);
and U1555 (N_1555,N_1236,N_1247);
nand U1556 (N_1556,N_1358,N_1353);
or U1557 (N_1557,N_1387,N_1289);
nand U1558 (N_1558,N_1318,N_1297);
nor U1559 (N_1559,N_1228,N_1352);
or U1560 (N_1560,N_1306,N_1205);
and U1561 (N_1561,N_1218,N_1284);
nor U1562 (N_1562,N_1397,N_1313);
nor U1563 (N_1563,N_1381,N_1331);
nor U1564 (N_1564,N_1330,N_1338);
nand U1565 (N_1565,N_1285,N_1262);
xnor U1566 (N_1566,N_1343,N_1201);
or U1567 (N_1567,N_1300,N_1226);
xor U1568 (N_1568,N_1213,N_1350);
nand U1569 (N_1569,N_1267,N_1252);
nor U1570 (N_1570,N_1355,N_1321);
nor U1571 (N_1571,N_1323,N_1347);
nor U1572 (N_1572,N_1347,N_1319);
and U1573 (N_1573,N_1251,N_1362);
and U1574 (N_1574,N_1204,N_1356);
nand U1575 (N_1575,N_1308,N_1321);
and U1576 (N_1576,N_1323,N_1272);
nor U1577 (N_1577,N_1314,N_1377);
or U1578 (N_1578,N_1289,N_1373);
nor U1579 (N_1579,N_1316,N_1291);
or U1580 (N_1580,N_1272,N_1352);
and U1581 (N_1581,N_1253,N_1220);
nand U1582 (N_1582,N_1267,N_1275);
nand U1583 (N_1583,N_1217,N_1221);
nor U1584 (N_1584,N_1253,N_1290);
nor U1585 (N_1585,N_1224,N_1394);
and U1586 (N_1586,N_1214,N_1283);
nor U1587 (N_1587,N_1246,N_1279);
or U1588 (N_1588,N_1391,N_1352);
and U1589 (N_1589,N_1355,N_1295);
and U1590 (N_1590,N_1363,N_1398);
nor U1591 (N_1591,N_1270,N_1321);
or U1592 (N_1592,N_1302,N_1234);
and U1593 (N_1593,N_1304,N_1256);
nor U1594 (N_1594,N_1290,N_1329);
nor U1595 (N_1595,N_1265,N_1321);
nor U1596 (N_1596,N_1294,N_1281);
xor U1597 (N_1597,N_1324,N_1261);
and U1598 (N_1598,N_1222,N_1255);
nand U1599 (N_1599,N_1253,N_1314);
and U1600 (N_1600,N_1424,N_1412);
nor U1601 (N_1601,N_1594,N_1589);
nor U1602 (N_1602,N_1415,N_1497);
nor U1603 (N_1603,N_1441,N_1473);
and U1604 (N_1604,N_1530,N_1451);
nor U1605 (N_1605,N_1432,N_1492);
and U1606 (N_1606,N_1519,N_1513);
nor U1607 (N_1607,N_1572,N_1577);
or U1608 (N_1608,N_1459,N_1562);
nand U1609 (N_1609,N_1574,N_1510);
nor U1610 (N_1610,N_1579,N_1538);
xor U1611 (N_1611,N_1452,N_1410);
nor U1612 (N_1612,N_1467,N_1431);
and U1613 (N_1613,N_1484,N_1503);
nand U1614 (N_1614,N_1475,N_1563);
or U1615 (N_1615,N_1533,N_1541);
and U1616 (N_1616,N_1578,N_1546);
nor U1617 (N_1617,N_1550,N_1597);
and U1618 (N_1618,N_1458,N_1421);
and U1619 (N_1619,N_1444,N_1559);
xor U1620 (N_1620,N_1526,N_1486);
and U1621 (N_1621,N_1403,N_1543);
and U1622 (N_1622,N_1501,N_1442);
and U1623 (N_1623,N_1439,N_1437);
and U1624 (N_1624,N_1545,N_1419);
nor U1625 (N_1625,N_1581,N_1416);
and U1626 (N_1626,N_1407,N_1447);
or U1627 (N_1627,N_1434,N_1445);
and U1628 (N_1628,N_1402,N_1423);
nor U1629 (N_1629,N_1554,N_1518);
nor U1630 (N_1630,N_1469,N_1471);
or U1631 (N_1631,N_1435,N_1587);
nor U1632 (N_1632,N_1417,N_1567);
and U1633 (N_1633,N_1512,N_1551);
nor U1634 (N_1634,N_1590,N_1438);
and U1635 (N_1635,N_1524,N_1585);
nand U1636 (N_1636,N_1511,N_1548);
nor U1637 (N_1637,N_1496,N_1544);
or U1638 (N_1638,N_1599,N_1547);
and U1639 (N_1639,N_1427,N_1401);
and U1640 (N_1640,N_1422,N_1520);
or U1641 (N_1641,N_1558,N_1478);
or U1642 (N_1642,N_1506,N_1509);
xnor U1643 (N_1643,N_1549,N_1450);
nand U1644 (N_1644,N_1472,N_1517);
and U1645 (N_1645,N_1468,N_1528);
nand U1646 (N_1646,N_1476,N_1453);
and U1647 (N_1647,N_1536,N_1569);
nor U1648 (N_1648,N_1592,N_1428);
or U1649 (N_1649,N_1470,N_1464);
nand U1650 (N_1650,N_1540,N_1532);
nand U1651 (N_1651,N_1433,N_1502);
nand U1652 (N_1652,N_1571,N_1521);
nand U1653 (N_1653,N_1429,N_1454);
and U1654 (N_1654,N_1565,N_1515);
nor U1655 (N_1655,N_1523,N_1539);
and U1656 (N_1656,N_1570,N_1493);
and U1657 (N_1657,N_1534,N_1418);
and U1658 (N_1658,N_1556,N_1576);
xor U1659 (N_1659,N_1588,N_1583);
nand U1660 (N_1660,N_1568,N_1404);
or U1661 (N_1661,N_1440,N_1490);
and U1662 (N_1662,N_1552,N_1598);
nor U1663 (N_1663,N_1466,N_1408);
and U1664 (N_1664,N_1495,N_1593);
xor U1665 (N_1665,N_1531,N_1414);
nand U1666 (N_1666,N_1477,N_1595);
nor U1667 (N_1667,N_1500,N_1406);
nor U1668 (N_1668,N_1409,N_1487);
nand U1669 (N_1669,N_1505,N_1456);
and U1670 (N_1670,N_1553,N_1460);
nor U1671 (N_1671,N_1535,N_1436);
nand U1672 (N_1672,N_1516,N_1485);
nand U1673 (N_1673,N_1504,N_1465);
nor U1674 (N_1674,N_1480,N_1463);
nand U1675 (N_1675,N_1507,N_1482);
nor U1676 (N_1676,N_1474,N_1491);
nor U1677 (N_1677,N_1560,N_1455);
nor U1678 (N_1678,N_1529,N_1449);
and U1679 (N_1679,N_1596,N_1584);
nand U1680 (N_1680,N_1498,N_1555);
nand U1681 (N_1681,N_1413,N_1573);
and U1682 (N_1682,N_1446,N_1489);
nand U1683 (N_1683,N_1582,N_1425);
or U1684 (N_1684,N_1411,N_1448);
and U1685 (N_1685,N_1481,N_1400);
and U1686 (N_1686,N_1537,N_1580);
xnor U1687 (N_1687,N_1426,N_1483);
or U1688 (N_1688,N_1405,N_1586);
nor U1689 (N_1689,N_1542,N_1461);
nor U1690 (N_1690,N_1508,N_1457);
and U1691 (N_1691,N_1575,N_1479);
nand U1692 (N_1692,N_1420,N_1561);
xnor U1693 (N_1693,N_1430,N_1564);
and U1694 (N_1694,N_1499,N_1488);
and U1695 (N_1695,N_1462,N_1525);
nor U1696 (N_1696,N_1591,N_1443);
or U1697 (N_1697,N_1514,N_1522);
xnor U1698 (N_1698,N_1527,N_1494);
nor U1699 (N_1699,N_1566,N_1557);
nand U1700 (N_1700,N_1593,N_1463);
nor U1701 (N_1701,N_1574,N_1597);
nand U1702 (N_1702,N_1596,N_1512);
nand U1703 (N_1703,N_1500,N_1463);
or U1704 (N_1704,N_1414,N_1404);
nor U1705 (N_1705,N_1482,N_1590);
nor U1706 (N_1706,N_1517,N_1475);
nand U1707 (N_1707,N_1405,N_1457);
or U1708 (N_1708,N_1421,N_1515);
or U1709 (N_1709,N_1586,N_1503);
or U1710 (N_1710,N_1557,N_1407);
or U1711 (N_1711,N_1453,N_1427);
and U1712 (N_1712,N_1578,N_1423);
nand U1713 (N_1713,N_1452,N_1438);
or U1714 (N_1714,N_1475,N_1508);
or U1715 (N_1715,N_1463,N_1485);
or U1716 (N_1716,N_1476,N_1420);
nand U1717 (N_1717,N_1526,N_1462);
nand U1718 (N_1718,N_1591,N_1491);
nor U1719 (N_1719,N_1567,N_1436);
nor U1720 (N_1720,N_1537,N_1424);
and U1721 (N_1721,N_1546,N_1516);
and U1722 (N_1722,N_1499,N_1590);
nand U1723 (N_1723,N_1584,N_1490);
and U1724 (N_1724,N_1593,N_1461);
and U1725 (N_1725,N_1495,N_1472);
xor U1726 (N_1726,N_1586,N_1406);
and U1727 (N_1727,N_1499,N_1576);
or U1728 (N_1728,N_1594,N_1474);
and U1729 (N_1729,N_1553,N_1400);
nand U1730 (N_1730,N_1466,N_1523);
and U1731 (N_1731,N_1560,N_1482);
or U1732 (N_1732,N_1574,N_1414);
or U1733 (N_1733,N_1482,N_1461);
and U1734 (N_1734,N_1402,N_1590);
nand U1735 (N_1735,N_1538,N_1474);
and U1736 (N_1736,N_1527,N_1565);
xor U1737 (N_1737,N_1437,N_1415);
or U1738 (N_1738,N_1533,N_1520);
or U1739 (N_1739,N_1405,N_1577);
xor U1740 (N_1740,N_1573,N_1440);
nand U1741 (N_1741,N_1581,N_1585);
nand U1742 (N_1742,N_1552,N_1508);
nor U1743 (N_1743,N_1585,N_1423);
nand U1744 (N_1744,N_1437,N_1560);
and U1745 (N_1745,N_1512,N_1561);
or U1746 (N_1746,N_1445,N_1592);
or U1747 (N_1747,N_1448,N_1557);
xor U1748 (N_1748,N_1571,N_1543);
nor U1749 (N_1749,N_1587,N_1411);
or U1750 (N_1750,N_1459,N_1538);
nor U1751 (N_1751,N_1478,N_1521);
or U1752 (N_1752,N_1596,N_1590);
or U1753 (N_1753,N_1540,N_1446);
nand U1754 (N_1754,N_1536,N_1432);
or U1755 (N_1755,N_1432,N_1456);
and U1756 (N_1756,N_1569,N_1496);
and U1757 (N_1757,N_1573,N_1442);
or U1758 (N_1758,N_1460,N_1463);
nor U1759 (N_1759,N_1467,N_1409);
nor U1760 (N_1760,N_1530,N_1444);
and U1761 (N_1761,N_1568,N_1563);
xnor U1762 (N_1762,N_1530,N_1526);
xnor U1763 (N_1763,N_1482,N_1462);
nor U1764 (N_1764,N_1496,N_1468);
or U1765 (N_1765,N_1552,N_1577);
nor U1766 (N_1766,N_1524,N_1583);
nor U1767 (N_1767,N_1545,N_1598);
nand U1768 (N_1768,N_1420,N_1413);
nand U1769 (N_1769,N_1446,N_1408);
nand U1770 (N_1770,N_1461,N_1467);
or U1771 (N_1771,N_1409,N_1578);
nand U1772 (N_1772,N_1581,N_1505);
nand U1773 (N_1773,N_1472,N_1503);
or U1774 (N_1774,N_1561,N_1414);
or U1775 (N_1775,N_1440,N_1489);
nor U1776 (N_1776,N_1439,N_1580);
nand U1777 (N_1777,N_1462,N_1412);
and U1778 (N_1778,N_1414,N_1406);
or U1779 (N_1779,N_1572,N_1529);
nand U1780 (N_1780,N_1459,N_1466);
nor U1781 (N_1781,N_1580,N_1576);
and U1782 (N_1782,N_1538,N_1446);
nand U1783 (N_1783,N_1520,N_1441);
nand U1784 (N_1784,N_1445,N_1567);
nor U1785 (N_1785,N_1512,N_1496);
or U1786 (N_1786,N_1470,N_1475);
nor U1787 (N_1787,N_1518,N_1565);
nand U1788 (N_1788,N_1448,N_1582);
and U1789 (N_1789,N_1474,N_1592);
or U1790 (N_1790,N_1516,N_1495);
nor U1791 (N_1791,N_1550,N_1588);
nor U1792 (N_1792,N_1454,N_1463);
and U1793 (N_1793,N_1590,N_1562);
nand U1794 (N_1794,N_1561,N_1470);
xor U1795 (N_1795,N_1556,N_1434);
nor U1796 (N_1796,N_1575,N_1515);
xnor U1797 (N_1797,N_1488,N_1413);
and U1798 (N_1798,N_1418,N_1455);
nor U1799 (N_1799,N_1496,N_1442);
nor U1800 (N_1800,N_1624,N_1766);
nand U1801 (N_1801,N_1785,N_1795);
and U1802 (N_1802,N_1731,N_1799);
or U1803 (N_1803,N_1714,N_1675);
nor U1804 (N_1804,N_1782,N_1767);
nand U1805 (N_1805,N_1745,N_1733);
or U1806 (N_1806,N_1789,N_1706);
nand U1807 (N_1807,N_1752,N_1705);
and U1808 (N_1808,N_1640,N_1651);
xor U1809 (N_1809,N_1788,N_1792);
and U1810 (N_1810,N_1747,N_1654);
and U1811 (N_1811,N_1794,N_1650);
nand U1812 (N_1812,N_1718,N_1626);
nand U1813 (N_1813,N_1781,N_1719);
nand U1814 (N_1814,N_1703,N_1727);
and U1815 (N_1815,N_1647,N_1663);
and U1816 (N_1816,N_1771,N_1758);
or U1817 (N_1817,N_1638,N_1725);
nor U1818 (N_1818,N_1635,N_1760);
xor U1819 (N_1819,N_1688,N_1614);
nor U1820 (N_1820,N_1672,N_1797);
and U1821 (N_1821,N_1798,N_1658);
xor U1822 (N_1822,N_1625,N_1662);
nor U1823 (N_1823,N_1678,N_1777);
nor U1824 (N_1824,N_1632,N_1616);
and U1825 (N_1825,N_1699,N_1645);
and U1826 (N_1826,N_1677,N_1652);
or U1827 (N_1827,N_1716,N_1746);
or U1828 (N_1828,N_1622,N_1664);
nand U1829 (N_1829,N_1721,N_1791);
or U1830 (N_1830,N_1770,N_1611);
nor U1831 (N_1831,N_1708,N_1709);
or U1832 (N_1832,N_1659,N_1723);
nand U1833 (N_1833,N_1713,N_1786);
or U1834 (N_1834,N_1633,N_1690);
and U1835 (N_1835,N_1710,N_1685);
or U1836 (N_1836,N_1609,N_1780);
or U1837 (N_1837,N_1689,N_1748);
nand U1838 (N_1838,N_1682,N_1653);
nand U1839 (N_1839,N_1720,N_1742);
nor U1840 (N_1840,N_1793,N_1735);
nor U1841 (N_1841,N_1796,N_1759);
nand U1842 (N_1842,N_1617,N_1765);
nand U1843 (N_1843,N_1711,N_1667);
and U1844 (N_1844,N_1603,N_1665);
or U1845 (N_1845,N_1773,N_1755);
and U1846 (N_1846,N_1669,N_1750);
or U1847 (N_1847,N_1649,N_1743);
nand U1848 (N_1848,N_1737,N_1757);
and U1849 (N_1849,N_1631,N_1621);
and U1850 (N_1850,N_1637,N_1712);
or U1851 (N_1851,N_1787,N_1761);
and U1852 (N_1852,N_1643,N_1762);
and U1853 (N_1853,N_1671,N_1776);
or U1854 (N_1854,N_1676,N_1612);
and U1855 (N_1855,N_1661,N_1630);
and U1856 (N_1856,N_1692,N_1623);
nor U1857 (N_1857,N_1769,N_1768);
and U1858 (N_1858,N_1790,N_1604);
xor U1859 (N_1859,N_1724,N_1600);
and U1860 (N_1860,N_1702,N_1660);
or U1861 (N_1861,N_1754,N_1741);
and U1862 (N_1862,N_1687,N_1607);
and U1863 (N_1863,N_1608,N_1615);
and U1864 (N_1864,N_1666,N_1684);
xor U1865 (N_1865,N_1697,N_1779);
or U1866 (N_1866,N_1778,N_1681);
and U1867 (N_1867,N_1619,N_1772);
xnor U1868 (N_1868,N_1639,N_1634);
or U1869 (N_1869,N_1736,N_1618);
or U1870 (N_1870,N_1775,N_1646);
nand U1871 (N_1871,N_1739,N_1644);
or U1872 (N_1872,N_1693,N_1674);
nor U1873 (N_1873,N_1751,N_1715);
and U1874 (N_1874,N_1606,N_1694);
and U1875 (N_1875,N_1683,N_1628);
nand U1876 (N_1876,N_1749,N_1717);
or U1877 (N_1877,N_1601,N_1784);
and U1878 (N_1878,N_1701,N_1642);
or U1879 (N_1879,N_1679,N_1656);
nand U1880 (N_1880,N_1620,N_1691);
or U1881 (N_1881,N_1763,N_1695);
nor U1882 (N_1882,N_1655,N_1686);
or U1883 (N_1883,N_1738,N_1613);
nor U1884 (N_1884,N_1636,N_1698);
nor U1885 (N_1885,N_1764,N_1696);
or U1886 (N_1886,N_1627,N_1673);
or U1887 (N_1887,N_1657,N_1734);
nor U1888 (N_1888,N_1707,N_1774);
or U1889 (N_1889,N_1740,N_1729);
or U1890 (N_1890,N_1670,N_1732);
or U1891 (N_1891,N_1602,N_1753);
and U1892 (N_1892,N_1680,N_1605);
nand U1893 (N_1893,N_1648,N_1641);
nor U1894 (N_1894,N_1704,N_1700);
nand U1895 (N_1895,N_1629,N_1726);
nand U1896 (N_1896,N_1756,N_1722);
nor U1897 (N_1897,N_1610,N_1783);
nor U1898 (N_1898,N_1668,N_1728);
or U1899 (N_1899,N_1744,N_1730);
or U1900 (N_1900,N_1760,N_1770);
and U1901 (N_1901,N_1714,N_1652);
nor U1902 (N_1902,N_1637,N_1603);
or U1903 (N_1903,N_1686,N_1717);
nor U1904 (N_1904,N_1780,N_1761);
and U1905 (N_1905,N_1613,N_1611);
xor U1906 (N_1906,N_1760,N_1772);
or U1907 (N_1907,N_1700,N_1696);
or U1908 (N_1908,N_1701,N_1759);
and U1909 (N_1909,N_1646,N_1794);
xor U1910 (N_1910,N_1644,N_1678);
xor U1911 (N_1911,N_1738,N_1775);
xnor U1912 (N_1912,N_1662,N_1626);
or U1913 (N_1913,N_1790,N_1755);
nor U1914 (N_1914,N_1727,N_1761);
nor U1915 (N_1915,N_1727,N_1752);
nand U1916 (N_1916,N_1722,N_1606);
xor U1917 (N_1917,N_1635,N_1765);
or U1918 (N_1918,N_1659,N_1751);
and U1919 (N_1919,N_1610,N_1647);
or U1920 (N_1920,N_1751,N_1644);
or U1921 (N_1921,N_1718,N_1654);
or U1922 (N_1922,N_1668,N_1650);
or U1923 (N_1923,N_1799,N_1636);
nor U1924 (N_1924,N_1657,N_1797);
and U1925 (N_1925,N_1785,N_1656);
or U1926 (N_1926,N_1635,N_1781);
or U1927 (N_1927,N_1710,N_1666);
or U1928 (N_1928,N_1640,N_1675);
nor U1929 (N_1929,N_1644,N_1729);
and U1930 (N_1930,N_1743,N_1792);
and U1931 (N_1931,N_1687,N_1674);
and U1932 (N_1932,N_1756,N_1607);
nand U1933 (N_1933,N_1622,N_1607);
nand U1934 (N_1934,N_1617,N_1728);
xnor U1935 (N_1935,N_1662,N_1711);
or U1936 (N_1936,N_1649,N_1735);
or U1937 (N_1937,N_1678,N_1743);
nand U1938 (N_1938,N_1664,N_1705);
xnor U1939 (N_1939,N_1680,N_1691);
xnor U1940 (N_1940,N_1703,N_1707);
and U1941 (N_1941,N_1713,N_1775);
or U1942 (N_1942,N_1674,N_1716);
or U1943 (N_1943,N_1695,N_1682);
nor U1944 (N_1944,N_1627,N_1671);
nor U1945 (N_1945,N_1623,N_1752);
nor U1946 (N_1946,N_1613,N_1775);
or U1947 (N_1947,N_1600,N_1771);
and U1948 (N_1948,N_1687,N_1638);
nor U1949 (N_1949,N_1637,N_1725);
and U1950 (N_1950,N_1629,N_1723);
nand U1951 (N_1951,N_1626,N_1765);
or U1952 (N_1952,N_1757,N_1713);
nand U1953 (N_1953,N_1626,N_1614);
or U1954 (N_1954,N_1711,N_1697);
nand U1955 (N_1955,N_1660,N_1738);
nand U1956 (N_1956,N_1776,N_1708);
nor U1957 (N_1957,N_1636,N_1620);
nand U1958 (N_1958,N_1785,N_1743);
nand U1959 (N_1959,N_1709,N_1698);
nand U1960 (N_1960,N_1637,N_1672);
nand U1961 (N_1961,N_1624,N_1614);
nand U1962 (N_1962,N_1743,N_1725);
or U1963 (N_1963,N_1635,N_1639);
and U1964 (N_1964,N_1658,N_1651);
nor U1965 (N_1965,N_1722,N_1735);
nand U1966 (N_1966,N_1777,N_1765);
nor U1967 (N_1967,N_1635,N_1743);
or U1968 (N_1968,N_1779,N_1778);
nor U1969 (N_1969,N_1665,N_1776);
nor U1970 (N_1970,N_1705,N_1754);
and U1971 (N_1971,N_1711,N_1661);
nor U1972 (N_1972,N_1758,N_1682);
nand U1973 (N_1973,N_1795,N_1792);
nand U1974 (N_1974,N_1788,N_1743);
nand U1975 (N_1975,N_1787,N_1669);
xor U1976 (N_1976,N_1609,N_1634);
or U1977 (N_1977,N_1650,N_1692);
xor U1978 (N_1978,N_1770,N_1722);
xnor U1979 (N_1979,N_1673,N_1637);
and U1980 (N_1980,N_1677,N_1645);
or U1981 (N_1981,N_1715,N_1621);
or U1982 (N_1982,N_1603,N_1645);
nand U1983 (N_1983,N_1740,N_1705);
nand U1984 (N_1984,N_1769,N_1601);
or U1985 (N_1985,N_1627,N_1778);
nand U1986 (N_1986,N_1656,N_1645);
and U1987 (N_1987,N_1767,N_1797);
nor U1988 (N_1988,N_1760,N_1678);
or U1989 (N_1989,N_1764,N_1614);
nand U1990 (N_1990,N_1620,N_1642);
nor U1991 (N_1991,N_1747,N_1663);
and U1992 (N_1992,N_1739,N_1716);
nand U1993 (N_1993,N_1725,N_1797);
nand U1994 (N_1994,N_1799,N_1747);
or U1995 (N_1995,N_1694,N_1715);
or U1996 (N_1996,N_1672,N_1611);
xor U1997 (N_1997,N_1628,N_1613);
or U1998 (N_1998,N_1790,N_1798);
or U1999 (N_1999,N_1609,N_1628);
nor U2000 (N_2000,N_1935,N_1835);
nor U2001 (N_2001,N_1944,N_1998);
nand U2002 (N_2002,N_1918,N_1866);
nor U2003 (N_2003,N_1828,N_1829);
nand U2004 (N_2004,N_1851,N_1999);
or U2005 (N_2005,N_1968,N_1811);
or U2006 (N_2006,N_1960,N_1967);
nand U2007 (N_2007,N_1943,N_1834);
or U2008 (N_2008,N_1945,N_1982);
and U2009 (N_2009,N_1898,N_1959);
nor U2010 (N_2010,N_1821,N_1961);
nand U2011 (N_2011,N_1983,N_1876);
nand U2012 (N_2012,N_1849,N_1870);
and U2013 (N_2013,N_1936,N_1922);
or U2014 (N_2014,N_1810,N_1939);
and U2015 (N_2015,N_1885,N_1859);
nor U2016 (N_2016,N_1981,N_1956);
nand U2017 (N_2017,N_1823,N_1895);
nor U2018 (N_2018,N_1973,N_1817);
and U2019 (N_2019,N_1803,N_1932);
nor U2020 (N_2020,N_1862,N_1871);
nand U2021 (N_2021,N_1891,N_1873);
and U2022 (N_2022,N_1893,N_1839);
and U2023 (N_2023,N_1869,N_1984);
and U2024 (N_2024,N_1845,N_1822);
nand U2025 (N_2025,N_1814,N_1841);
nand U2026 (N_2026,N_1946,N_1934);
nand U2027 (N_2027,N_1825,N_1972);
and U2028 (N_2028,N_1970,N_1801);
and U2029 (N_2029,N_1903,N_1980);
xor U2030 (N_2030,N_1966,N_1996);
nor U2031 (N_2031,N_1975,N_1833);
nand U2032 (N_2032,N_1995,N_1800);
or U2033 (N_2033,N_1997,N_1824);
and U2034 (N_2034,N_1840,N_1872);
xor U2035 (N_2035,N_1954,N_1940);
and U2036 (N_2036,N_1897,N_1826);
nand U2037 (N_2037,N_1947,N_1853);
or U2038 (N_2038,N_1923,N_1938);
and U2039 (N_2039,N_1830,N_1908);
or U2040 (N_2040,N_1951,N_1950);
nand U2041 (N_2041,N_1921,N_1927);
nor U2042 (N_2042,N_1881,N_1877);
and U2043 (N_2043,N_1805,N_1924);
or U2044 (N_2044,N_1812,N_1847);
and U2045 (N_2045,N_1900,N_1925);
or U2046 (N_2046,N_1831,N_1875);
and U2047 (N_2047,N_1912,N_1916);
nor U2048 (N_2048,N_1978,N_1969);
or U2049 (N_2049,N_1902,N_1868);
or U2050 (N_2050,N_1974,N_1964);
or U2051 (N_2051,N_1994,N_1992);
nor U2052 (N_2052,N_1931,N_1990);
xor U2053 (N_2053,N_1977,N_1993);
nand U2054 (N_2054,N_1813,N_1878);
nor U2055 (N_2055,N_1929,N_1901);
nor U2056 (N_2056,N_1911,N_1941);
nand U2057 (N_2057,N_1819,N_1857);
nand U2058 (N_2058,N_1861,N_1986);
nand U2059 (N_2059,N_1842,N_1919);
and U2060 (N_2060,N_1848,N_1809);
or U2061 (N_2061,N_1899,N_1915);
nor U2062 (N_2062,N_1827,N_1856);
nor U2063 (N_2063,N_1926,N_1949);
or U2064 (N_2064,N_1913,N_1854);
nand U2065 (N_2065,N_1948,N_1883);
and U2066 (N_2066,N_1838,N_1955);
nand U2067 (N_2067,N_1879,N_1864);
nor U2068 (N_2068,N_1843,N_1888);
nand U2069 (N_2069,N_1815,N_1892);
nor U2070 (N_2070,N_1953,N_1928);
nand U2071 (N_2071,N_1820,N_1852);
nor U2072 (N_2072,N_1957,N_1965);
nor U2073 (N_2073,N_1958,N_1889);
nand U2074 (N_2074,N_1976,N_1952);
nand U2075 (N_2075,N_1904,N_1874);
nor U2076 (N_2076,N_1937,N_1985);
nand U2077 (N_2077,N_1989,N_1837);
nor U2078 (N_2078,N_1920,N_1880);
nor U2079 (N_2079,N_1867,N_1933);
nand U2080 (N_2080,N_1816,N_1832);
and U2081 (N_2081,N_1860,N_1846);
xor U2082 (N_2082,N_1887,N_1917);
nand U2083 (N_2083,N_1818,N_1930);
nor U2084 (N_2084,N_1806,N_1963);
nand U2085 (N_2085,N_1855,N_1910);
or U2086 (N_2086,N_1808,N_1909);
or U2087 (N_2087,N_1844,N_1905);
or U2088 (N_2088,N_1836,N_1804);
or U2089 (N_2089,N_1987,N_1971);
nand U2090 (N_2090,N_1962,N_1907);
xnor U2091 (N_2091,N_1914,N_1890);
nand U2092 (N_2092,N_1865,N_1896);
or U2093 (N_2093,N_1991,N_1882);
and U2094 (N_2094,N_1979,N_1802);
nand U2095 (N_2095,N_1886,N_1807);
nor U2096 (N_2096,N_1906,N_1988);
nor U2097 (N_2097,N_1863,N_1858);
and U2098 (N_2098,N_1894,N_1850);
and U2099 (N_2099,N_1942,N_1884);
nand U2100 (N_2100,N_1947,N_1883);
nor U2101 (N_2101,N_1972,N_1936);
or U2102 (N_2102,N_1959,N_1970);
nand U2103 (N_2103,N_1901,N_1981);
or U2104 (N_2104,N_1874,N_1856);
nand U2105 (N_2105,N_1968,N_1864);
nand U2106 (N_2106,N_1813,N_1981);
nand U2107 (N_2107,N_1928,N_1835);
nor U2108 (N_2108,N_1842,N_1859);
nand U2109 (N_2109,N_1847,N_1805);
and U2110 (N_2110,N_1867,N_1993);
and U2111 (N_2111,N_1895,N_1998);
and U2112 (N_2112,N_1971,N_1893);
nor U2113 (N_2113,N_1866,N_1815);
xnor U2114 (N_2114,N_1813,N_1974);
or U2115 (N_2115,N_1848,N_1966);
or U2116 (N_2116,N_1853,N_1832);
xnor U2117 (N_2117,N_1867,N_1927);
and U2118 (N_2118,N_1932,N_1802);
nand U2119 (N_2119,N_1982,N_1956);
nor U2120 (N_2120,N_1827,N_1937);
nand U2121 (N_2121,N_1935,N_1965);
or U2122 (N_2122,N_1985,N_1910);
nand U2123 (N_2123,N_1980,N_1853);
nor U2124 (N_2124,N_1929,N_1912);
nor U2125 (N_2125,N_1875,N_1837);
nor U2126 (N_2126,N_1986,N_1926);
nand U2127 (N_2127,N_1808,N_1903);
xnor U2128 (N_2128,N_1822,N_1842);
and U2129 (N_2129,N_1987,N_1886);
nor U2130 (N_2130,N_1931,N_1879);
xnor U2131 (N_2131,N_1966,N_1982);
nand U2132 (N_2132,N_1985,N_1890);
or U2133 (N_2133,N_1892,N_1811);
xor U2134 (N_2134,N_1834,N_1836);
or U2135 (N_2135,N_1943,N_1820);
xor U2136 (N_2136,N_1992,N_1927);
nand U2137 (N_2137,N_1842,N_1990);
or U2138 (N_2138,N_1909,N_1827);
nor U2139 (N_2139,N_1890,N_1835);
xnor U2140 (N_2140,N_1866,N_1926);
nor U2141 (N_2141,N_1818,N_1840);
nand U2142 (N_2142,N_1921,N_1995);
nor U2143 (N_2143,N_1969,N_1979);
nor U2144 (N_2144,N_1987,N_1965);
and U2145 (N_2145,N_1880,N_1957);
nor U2146 (N_2146,N_1863,N_1852);
or U2147 (N_2147,N_1856,N_1840);
nor U2148 (N_2148,N_1972,N_1978);
and U2149 (N_2149,N_1940,N_1809);
and U2150 (N_2150,N_1996,N_1939);
and U2151 (N_2151,N_1982,N_1815);
nand U2152 (N_2152,N_1916,N_1863);
or U2153 (N_2153,N_1974,N_1872);
and U2154 (N_2154,N_1933,N_1821);
or U2155 (N_2155,N_1821,N_1884);
nand U2156 (N_2156,N_1931,N_1938);
or U2157 (N_2157,N_1893,N_1991);
xnor U2158 (N_2158,N_1918,N_1987);
and U2159 (N_2159,N_1976,N_1993);
nand U2160 (N_2160,N_1831,N_1856);
and U2161 (N_2161,N_1951,N_1943);
or U2162 (N_2162,N_1805,N_1938);
or U2163 (N_2163,N_1818,N_1800);
nor U2164 (N_2164,N_1824,N_1853);
or U2165 (N_2165,N_1952,N_1893);
nand U2166 (N_2166,N_1840,N_1860);
or U2167 (N_2167,N_1969,N_1831);
or U2168 (N_2168,N_1815,N_1851);
xor U2169 (N_2169,N_1969,N_1871);
or U2170 (N_2170,N_1827,N_1826);
nor U2171 (N_2171,N_1945,N_1962);
nor U2172 (N_2172,N_1967,N_1936);
nor U2173 (N_2173,N_1984,N_1955);
or U2174 (N_2174,N_1992,N_1985);
and U2175 (N_2175,N_1889,N_1903);
nor U2176 (N_2176,N_1996,N_1891);
or U2177 (N_2177,N_1823,N_1923);
nor U2178 (N_2178,N_1861,N_1821);
nor U2179 (N_2179,N_1991,N_1937);
nand U2180 (N_2180,N_1862,N_1927);
nand U2181 (N_2181,N_1844,N_1830);
or U2182 (N_2182,N_1892,N_1898);
and U2183 (N_2183,N_1849,N_1837);
or U2184 (N_2184,N_1969,N_1829);
nor U2185 (N_2185,N_1928,N_1823);
xnor U2186 (N_2186,N_1819,N_1986);
and U2187 (N_2187,N_1839,N_1924);
nor U2188 (N_2188,N_1819,N_1998);
and U2189 (N_2189,N_1843,N_1816);
and U2190 (N_2190,N_1989,N_1963);
xor U2191 (N_2191,N_1991,N_1972);
or U2192 (N_2192,N_1801,N_1875);
nand U2193 (N_2193,N_1870,N_1845);
or U2194 (N_2194,N_1999,N_1913);
and U2195 (N_2195,N_1903,N_1938);
nor U2196 (N_2196,N_1844,N_1985);
xor U2197 (N_2197,N_1846,N_1842);
xnor U2198 (N_2198,N_1876,N_1821);
nand U2199 (N_2199,N_1857,N_1873);
and U2200 (N_2200,N_2115,N_2139);
xor U2201 (N_2201,N_2073,N_2154);
and U2202 (N_2202,N_2068,N_2042);
and U2203 (N_2203,N_2137,N_2004);
nor U2204 (N_2204,N_2003,N_2136);
nor U2205 (N_2205,N_2124,N_2030);
or U2206 (N_2206,N_2160,N_2100);
nor U2207 (N_2207,N_2118,N_2001);
nor U2208 (N_2208,N_2016,N_2049);
nor U2209 (N_2209,N_2191,N_2062);
nand U2210 (N_2210,N_2164,N_2149);
or U2211 (N_2211,N_2085,N_2086);
xor U2212 (N_2212,N_2040,N_2117);
nor U2213 (N_2213,N_2194,N_2091);
or U2214 (N_2214,N_2105,N_2186);
nor U2215 (N_2215,N_2190,N_2078);
nand U2216 (N_2216,N_2130,N_2132);
nand U2217 (N_2217,N_2083,N_2059);
nand U2218 (N_2218,N_2155,N_2039);
nand U2219 (N_2219,N_2008,N_2007);
nand U2220 (N_2220,N_2171,N_2022);
xor U2221 (N_2221,N_2097,N_2143);
nand U2222 (N_2222,N_2080,N_2052);
and U2223 (N_2223,N_2090,N_2046);
nor U2224 (N_2224,N_2138,N_2034);
xor U2225 (N_2225,N_2000,N_2168);
or U2226 (N_2226,N_2029,N_2157);
nor U2227 (N_2227,N_2065,N_2187);
nand U2228 (N_2228,N_2096,N_2076);
nand U2229 (N_2229,N_2174,N_2075);
or U2230 (N_2230,N_2082,N_2088);
xnor U2231 (N_2231,N_2113,N_2144);
nor U2232 (N_2232,N_2066,N_2167);
nor U2233 (N_2233,N_2189,N_2026);
nand U2234 (N_2234,N_2145,N_2162);
or U2235 (N_2235,N_2092,N_2010);
and U2236 (N_2236,N_2147,N_2192);
and U2237 (N_2237,N_2087,N_2125);
xnor U2238 (N_2238,N_2199,N_2079);
xor U2239 (N_2239,N_2027,N_2063);
xor U2240 (N_2240,N_2054,N_2110);
or U2241 (N_2241,N_2148,N_2181);
and U2242 (N_2242,N_2151,N_2089);
nor U2243 (N_2243,N_2146,N_2109);
or U2244 (N_2244,N_2107,N_2077);
or U2245 (N_2245,N_2177,N_2180);
xor U2246 (N_2246,N_2179,N_2178);
nand U2247 (N_2247,N_2018,N_2095);
nand U2248 (N_2248,N_2112,N_2102);
nand U2249 (N_2249,N_2128,N_2025);
xor U2250 (N_2250,N_2012,N_2058);
and U2251 (N_2251,N_2045,N_2158);
nor U2252 (N_2252,N_2099,N_2033);
nand U2253 (N_2253,N_2006,N_2044);
or U2254 (N_2254,N_2197,N_2056);
xor U2255 (N_2255,N_2094,N_2170);
and U2256 (N_2256,N_2084,N_2120);
nand U2257 (N_2257,N_2081,N_2067);
nor U2258 (N_2258,N_2198,N_2123);
and U2259 (N_2259,N_2126,N_2141);
and U2260 (N_2260,N_2013,N_2116);
nor U2261 (N_2261,N_2153,N_2176);
nand U2262 (N_2262,N_2037,N_2122);
or U2263 (N_2263,N_2093,N_2031);
nor U2264 (N_2264,N_2188,N_2161);
and U2265 (N_2265,N_2108,N_2048);
nor U2266 (N_2266,N_2043,N_2020);
and U2267 (N_2267,N_2057,N_2071);
or U2268 (N_2268,N_2142,N_2070);
or U2269 (N_2269,N_2182,N_2193);
or U2270 (N_2270,N_2053,N_2166);
and U2271 (N_2271,N_2002,N_2019);
nand U2272 (N_2272,N_2014,N_2009);
nand U2273 (N_2273,N_2172,N_2101);
xnor U2274 (N_2274,N_2061,N_2103);
xnor U2275 (N_2275,N_2055,N_2165);
nor U2276 (N_2276,N_2140,N_2129);
nor U2277 (N_2277,N_2185,N_2121);
nor U2278 (N_2278,N_2169,N_2047);
and U2279 (N_2279,N_2127,N_2038);
nor U2280 (N_2280,N_2111,N_2032);
xor U2281 (N_2281,N_2098,N_2131);
nor U2282 (N_2282,N_2011,N_2184);
nor U2283 (N_2283,N_2060,N_2050);
nand U2284 (N_2284,N_2106,N_2041);
and U2285 (N_2285,N_2021,N_2133);
nor U2286 (N_2286,N_2195,N_2159);
nor U2287 (N_2287,N_2175,N_2135);
nand U2288 (N_2288,N_2005,N_2064);
and U2289 (N_2289,N_2015,N_2035);
and U2290 (N_2290,N_2104,N_2163);
nand U2291 (N_2291,N_2074,N_2173);
or U2292 (N_2292,N_2183,N_2196);
or U2293 (N_2293,N_2134,N_2036);
nand U2294 (N_2294,N_2152,N_2150);
nand U2295 (N_2295,N_2017,N_2069);
and U2296 (N_2296,N_2156,N_2023);
or U2297 (N_2297,N_2072,N_2114);
nand U2298 (N_2298,N_2024,N_2028);
nand U2299 (N_2299,N_2119,N_2051);
and U2300 (N_2300,N_2089,N_2155);
nand U2301 (N_2301,N_2165,N_2174);
nor U2302 (N_2302,N_2082,N_2079);
nor U2303 (N_2303,N_2166,N_2054);
xor U2304 (N_2304,N_2018,N_2071);
nor U2305 (N_2305,N_2101,N_2073);
nor U2306 (N_2306,N_2106,N_2102);
xnor U2307 (N_2307,N_2008,N_2097);
nor U2308 (N_2308,N_2016,N_2191);
and U2309 (N_2309,N_2070,N_2158);
nand U2310 (N_2310,N_2179,N_2184);
nor U2311 (N_2311,N_2076,N_2145);
nand U2312 (N_2312,N_2184,N_2026);
and U2313 (N_2313,N_2054,N_2071);
or U2314 (N_2314,N_2057,N_2198);
and U2315 (N_2315,N_2192,N_2054);
nor U2316 (N_2316,N_2046,N_2012);
or U2317 (N_2317,N_2095,N_2187);
and U2318 (N_2318,N_2165,N_2192);
and U2319 (N_2319,N_2107,N_2069);
nand U2320 (N_2320,N_2092,N_2128);
nand U2321 (N_2321,N_2119,N_2009);
and U2322 (N_2322,N_2119,N_2115);
and U2323 (N_2323,N_2007,N_2027);
or U2324 (N_2324,N_2193,N_2116);
nand U2325 (N_2325,N_2144,N_2103);
nor U2326 (N_2326,N_2008,N_2157);
or U2327 (N_2327,N_2051,N_2041);
nor U2328 (N_2328,N_2188,N_2018);
and U2329 (N_2329,N_2009,N_2136);
nor U2330 (N_2330,N_2089,N_2149);
nand U2331 (N_2331,N_2058,N_2053);
nor U2332 (N_2332,N_2134,N_2195);
nor U2333 (N_2333,N_2187,N_2075);
nor U2334 (N_2334,N_2062,N_2090);
and U2335 (N_2335,N_2009,N_2112);
or U2336 (N_2336,N_2077,N_2112);
nand U2337 (N_2337,N_2020,N_2067);
or U2338 (N_2338,N_2059,N_2126);
or U2339 (N_2339,N_2100,N_2082);
nor U2340 (N_2340,N_2172,N_2064);
and U2341 (N_2341,N_2121,N_2079);
nor U2342 (N_2342,N_2010,N_2077);
and U2343 (N_2343,N_2012,N_2070);
nor U2344 (N_2344,N_2053,N_2105);
and U2345 (N_2345,N_2093,N_2199);
nor U2346 (N_2346,N_2003,N_2001);
and U2347 (N_2347,N_2131,N_2030);
or U2348 (N_2348,N_2167,N_2012);
or U2349 (N_2349,N_2158,N_2065);
nor U2350 (N_2350,N_2024,N_2124);
xnor U2351 (N_2351,N_2104,N_2160);
nor U2352 (N_2352,N_2138,N_2158);
nand U2353 (N_2353,N_2004,N_2029);
or U2354 (N_2354,N_2018,N_2077);
or U2355 (N_2355,N_2011,N_2063);
and U2356 (N_2356,N_2041,N_2175);
or U2357 (N_2357,N_2143,N_2141);
nand U2358 (N_2358,N_2050,N_2010);
and U2359 (N_2359,N_2050,N_2055);
nor U2360 (N_2360,N_2199,N_2139);
or U2361 (N_2361,N_2151,N_2133);
nor U2362 (N_2362,N_2067,N_2126);
nand U2363 (N_2363,N_2119,N_2043);
or U2364 (N_2364,N_2102,N_2002);
nand U2365 (N_2365,N_2145,N_2173);
nand U2366 (N_2366,N_2068,N_2074);
nand U2367 (N_2367,N_2099,N_2136);
xor U2368 (N_2368,N_2113,N_2107);
and U2369 (N_2369,N_2163,N_2099);
nor U2370 (N_2370,N_2185,N_2174);
and U2371 (N_2371,N_2044,N_2094);
and U2372 (N_2372,N_2130,N_2142);
nand U2373 (N_2373,N_2103,N_2075);
nor U2374 (N_2374,N_2123,N_2005);
nor U2375 (N_2375,N_2098,N_2130);
or U2376 (N_2376,N_2098,N_2052);
nand U2377 (N_2377,N_2116,N_2138);
nand U2378 (N_2378,N_2026,N_2013);
nand U2379 (N_2379,N_2017,N_2068);
nand U2380 (N_2380,N_2062,N_2064);
or U2381 (N_2381,N_2123,N_2040);
or U2382 (N_2382,N_2195,N_2122);
and U2383 (N_2383,N_2049,N_2129);
and U2384 (N_2384,N_2008,N_2196);
or U2385 (N_2385,N_2194,N_2018);
nand U2386 (N_2386,N_2134,N_2013);
or U2387 (N_2387,N_2026,N_2197);
or U2388 (N_2388,N_2076,N_2133);
nor U2389 (N_2389,N_2183,N_2030);
nand U2390 (N_2390,N_2152,N_2157);
nand U2391 (N_2391,N_2012,N_2006);
or U2392 (N_2392,N_2161,N_2059);
xor U2393 (N_2393,N_2104,N_2103);
nand U2394 (N_2394,N_2180,N_2136);
xnor U2395 (N_2395,N_2062,N_2155);
or U2396 (N_2396,N_2159,N_2103);
or U2397 (N_2397,N_2147,N_2056);
nand U2398 (N_2398,N_2131,N_2124);
nor U2399 (N_2399,N_2193,N_2162);
and U2400 (N_2400,N_2252,N_2390);
nand U2401 (N_2401,N_2357,N_2293);
and U2402 (N_2402,N_2386,N_2398);
nor U2403 (N_2403,N_2397,N_2335);
nand U2404 (N_2404,N_2200,N_2268);
nand U2405 (N_2405,N_2253,N_2388);
nor U2406 (N_2406,N_2230,N_2381);
and U2407 (N_2407,N_2221,N_2236);
nor U2408 (N_2408,N_2208,N_2322);
nand U2409 (N_2409,N_2326,N_2231);
and U2410 (N_2410,N_2389,N_2209);
and U2411 (N_2411,N_2399,N_2316);
or U2412 (N_2412,N_2233,N_2291);
or U2413 (N_2413,N_2393,N_2356);
or U2414 (N_2414,N_2224,N_2307);
nand U2415 (N_2415,N_2301,N_2262);
nor U2416 (N_2416,N_2330,N_2333);
xor U2417 (N_2417,N_2303,N_2368);
nand U2418 (N_2418,N_2258,N_2271);
and U2419 (N_2419,N_2275,N_2324);
nor U2420 (N_2420,N_2302,N_2225);
nand U2421 (N_2421,N_2338,N_2249);
and U2422 (N_2422,N_2371,N_2234);
or U2423 (N_2423,N_2396,N_2214);
nor U2424 (N_2424,N_2321,N_2286);
nor U2425 (N_2425,N_2319,N_2325);
or U2426 (N_2426,N_2384,N_2372);
nor U2427 (N_2427,N_2254,N_2220);
nand U2428 (N_2428,N_2212,N_2317);
nand U2429 (N_2429,N_2340,N_2226);
and U2430 (N_2430,N_2295,N_2240);
nand U2431 (N_2431,N_2279,N_2383);
nor U2432 (N_2432,N_2363,N_2243);
or U2433 (N_2433,N_2354,N_2277);
and U2434 (N_2434,N_2216,N_2255);
or U2435 (N_2435,N_2219,N_2395);
nor U2436 (N_2436,N_2203,N_2264);
nand U2437 (N_2437,N_2260,N_2201);
and U2438 (N_2438,N_2229,N_2353);
nand U2439 (N_2439,N_2362,N_2235);
nor U2440 (N_2440,N_2342,N_2288);
nor U2441 (N_2441,N_2223,N_2278);
or U2442 (N_2442,N_2211,N_2344);
nor U2443 (N_2443,N_2306,N_2210);
nor U2444 (N_2444,N_2334,N_2350);
and U2445 (N_2445,N_2366,N_2385);
nand U2446 (N_2446,N_2281,N_2289);
nor U2447 (N_2447,N_2348,N_2305);
nor U2448 (N_2448,N_2337,N_2375);
nor U2449 (N_2449,N_2245,N_2267);
nor U2450 (N_2450,N_2364,N_2308);
nor U2451 (N_2451,N_2373,N_2239);
xnor U2452 (N_2452,N_2232,N_2228);
xnor U2453 (N_2453,N_2358,N_2296);
or U2454 (N_2454,N_2273,N_2204);
or U2455 (N_2455,N_2251,N_2272);
xor U2456 (N_2456,N_2346,N_2367);
and U2457 (N_2457,N_2259,N_2377);
nand U2458 (N_2458,N_2343,N_2370);
nand U2459 (N_2459,N_2290,N_2311);
and U2460 (N_2460,N_2300,N_2365);
nand U2461 (N_2461,N_2270,N_2244);
and U2462 (N_2462,N_2359,N_2294);
xor U2463 (N_2463,N_2206,N_2394);
and U2464 (N_2464,N_2309,N_2352);
and U2465 (N_2465,N_2332,N_2292);
or U2466 (N_2466,N_2378,N_2285);
nor U2467 (N_2467,N_2360,N_2382);
nand U2468 (N_2468,N_2222,N_2287);
nor U2469 (N_2469,N_2246,N_2202);
nand U2470 (N_2470,N_2376,N_2282);
or U2471 (N_2471,N_2265,N_2274);
and U2472 (N_2472,N_2331,N_2261);
and U2473 (N_2473,N_2315,N_2256);
nor U2474 (N_2474,N_2218,N_2336);
and U2475 (N_2475,N_2345,N_2313);
nand U2476 (N_2476,N_2318,N_2276);
nand U2477 (N_2477,N_2238,N_2310);
and U2478 (N_2478,N_2263,N_2215);
or U2479 (N_2479,N_2349,N_2207);
nand U2480 (N_2480,N_2242,N_2379);
nor U2481 (N_2481,N_2347,N_2205);
nand U2482 (N_2482,N_2327,N_2392);
nor U2483 (N_2483,N_2237,N_2391);
nor U2484 (N_2484,N_2298,N_2351);
nand U2485 (N_2485,N_2312,N_2266);
nand U2486 (N_2486,N_2297,N_2257);
nor U2487 (N_2487,N_2374,N_2284);
and U2488 (N_2488,N_2241,N_2361);
nand U2489 (N_2489,N_2280,N_2250);
and U2490 (N_2490,N_2299,N_2320);
nand U2491 (N_2491,N_2248,N_2339);
or U2492 (N_2492,N_2328,N_2217);
nand U2493 (N_2493,N_2213,N_2329);
nor U2494 (N_2494,N_2304,N_2227);
and U2495 (N_2495,N_2380,N_2369);
xor U2496 (N_2496,N_2387,N_2323);
or U2497 (N_2497,N_2314,N_2283);
nor U2498 (N_2498,N_2269,N_2341);
or U2499 (N_2499,N_2355,N_2247);
nand U2500 (N_2500,N_2239,N_2353);
or U2501 (N_2501,N_2317,N_2349);
and U2502 (N_2502,N_2229,N_2342);
xor U2503 (N_2503,N_2223,N_2235);
nor U2504 (N_2504,N_2200,N_2318);
or U2505 (N_2505,N_2337,N_2315);
or U2506 (N_2506,N_2372,N_2354);
nor U2507 (N_2507,N_2250,N_2357);
or U2508 (N_2508,N_2263,N_2240);
xor U2509 (N_2509,N_2254,N_2299);
and U2510 (N_2510,N_2357,N_2235);
or U2511 (N_2511,N_2313,N_2355);
or U2512 (N_2512,N_2235,N_2387);
or U2513 (N_2513,N_2310,N_2257);
xnor U2514 (N_2514,N_2274,N_2389);
or U2515 (N_2515,N_2316,N_2326);
or U2516 (N_2516,N_2229,N_2386);
or U2517 (N_2517,N_2393,N_2366);
nand U2518 (N_2518,N_2374,N_2260);
nand U2519 (N_2519,N_2250,N_2325);
or U2520 (N_2520,N_2383,N_2312);
nor U2521 (N_2521,N_2387,N_2328);
xor U2522 (N_2522,N_2302,N_2266);
and U2523 (N_2523,N_2288,N_2256);
nor U2524 (N_2524,N_2217,N_2288);
or U2525 (N_2525,N_2300,N_2360);
and U2526 (N_2526,N_2215,N_2384);
and U2527 (N_2527,N_2346,N_2227);
and U2528 (N_2528,N_2284,N_2214);
or U2529 (N_2529,N_2262,N_2324);
and U2530 (N_2530,N_2341,N_2255);
nand U2531 (N_2531,N_2256,N_2298);
nor U2532 (N_2532,N_2205,N_2360);
and U2533 (N_2533,N_2277,N_2295);
or U2534 (N_2534,N_2362,N_2347);
nor U2535 (N_2535,N_2317,N_2264);
nand U2536 (N_2536,N_2248,N_2337);
xor U2537 (N_2537,N_2369,N_2277);
or U2538 (N_2538,N_2279,N_2231);
nand U2539 (N_2539,N_2375,N_2341);
or U2540 (N_2540,N_2390,N_2227);
or U2541 (N_2541,N_2256,N_2399);
nand U2542 (N_2542,N_2250,N_2267);
nand U2543 (N_2543,N_2389,N_2276);
nor U2544 (N_2544,N_2238,N_2335);
nor U2545 (N_2545,N_2300,N_2279);
and U2546 (N_2546,N_2298,N_2368);
or U2547 (N_2547,N_2233,N_2269);
nand U2548 (N_2548,N_2265,N_2390);
xor U2549 (N_2549,N_2387,N_2279);
or U2550 (N_2550,N_2239,N_2377);
or U2551 (N_2551,N_2330,N_2326);
nor U2552 (N_2552,N_2276,N_2329);
or U2553 (N_2553,N_2214,N_2376);
and U2554 (N_2554,N_2259,N_2241);
xnor U2555 (N_2555,N_2348,N_2270);
nor U2556 (N_2556,N_2313,N_2241);
xor U2557 (N_2557,N_2253,N_2232);
or U2558 (N_2558,N_2206,N_2289);
xnor U2559 (N_2559,N_2277,N_2223);
xor U2560 (N_2560,N_2330,N_2381);
nor U2561 (N_2561,N_2373,N_2370);
nor U2562 (N_2562,N_2223,N_2380);
nor U2563 (N_2563,N_2371,N_2352);
nor U2564 (N_2564,N_2397,N_2388);
nor U2565 (N_2565,N_2340,N_2260);
and U2566 (N_2566,N_2225,N_2358);
nor U2567 (N_2567,N_2392,N_2273);
and U2568 (N_2568,N_2353,N_2288);
and U2569 (N_2569,N_2296,N_2285);
and U2570 (N_2570,N_2228,N_2231);
or U2571 (N_2571,N_2224,N_2331);
xnor U2572 (N_2572,N_2228,N_2383);
nand U2573 (N_2573,N_2261,N_2248);
nand U2574 (N_2574,N_2382,N_2396);
nand U2575 (N_2575,N_2367,N_2327);
xor U2576 (N_2576,N_2331,N_2350);
nor U2577 (N_2577,N_2246,N_2337);
xor U2578 (N_2578,N_2361,N_2339);
and U2579 (N_2579,N_2285,N_2260);
nand U2580 (N_2580,N_2335,N_2235);
nor U2581 (N_2581,N_2258,N_2395);
and U2582 (N_2582,N_2291,N_2230);
nor U2583 (N_2583,N_2265,N_2283);
nor U2584 (N_2584,N_2252,N_2249);
nand U2585 (N_2585,N_2299,N_2274);
and U2586 (N_2586,N_2303,N_2212);
and U2587 (N_2587,N_2388,N_2235);
and U2588 (N_2588,N_2235,N_2266);
xnor U2589 (N_2589,N_2355,N_2203);
and U2590 (N_2590,N_2261,N_2357);
or U2591 (N_2591,N_2277,N_2211);
nor U2592 (N_2592,N_2270,N_2368);
nor U2593 (N_2593,N_2211,N_2236);
nor U2594 (N_2594,N_2235,N_2298);
or U2595 (N_2595,N_2288,N_2364);
or U2596 (N_2596,N_2325,N_2324);
nand U2597 (N_2597,N_2265,N_2329);
or U2598 (N_2598,N_2295,N_2223);
nor U2599 (N_2599,N_2365,N_2284);
and U2600 (N_2600,N_2417,N_2415);
or U2601 (N_2601,N_2496,N_2562);
nor U2602 (N_2602,N_2485,N_2502);
nor U2603 (N_2603,N_2536,N_2522);
xnor U2604 (N_2604,N_2526,N_2486);
or U2605 (N_2605,N_2494,N_2513);
nor U2606 (N_2606,N_2529,N_2487);
and U2607 (N_2607,N_2431,N_2473);
nor U2608 (N_2608,N_2515,N_2414);
nor U2609 (N_2609,N_2564,N_2576);
and U2610 (N_2610,N_2454,N_2461);
and U2611 (N_2611,N_2438,N_2514);
nor U2612 (N_2612,N_2488,N_2447);
or U2613 (N_2613,N_2533,N_2423);
or U2614 (N_2614,N_2409,N_2462);
and U2615 (N_2615,N_2538,N_2528);
nor U2616 (N_2616,N_2599,N_2455);
nor U2617 (N_2617,N_2521,N_2559);
nand U2618 (N_2618,N_2503,N_2586);
nor U2619 (N_2619,N_2540,N_2549);
or U2620 (N_2620,N_2491,N_2523);
or U2621 (N_2621,N_2553,N_2594);
or U2622 (N_2622,N_2580,N_2456);
nor U2623 (N_2623,N_2537,N_2499);
and U2624 (N_2624,N_2500,N_2505);
nand U2625 (N_2625,N_2495,N_2575);
nand U2626 (N_2626,N_2430,N_2589);
nor U2627 (N_2627,N_2452,N_2595);
xnor U2628 (N_2628,N_2565,N_2410);
nand U2629 (N_2629,N_2401,N_2466);
nand U2630 (N_2630,N_2403,N_2520);
xor U2631 (N_2631,N_2527,N_2463);
or U2632 (N_2632,N_2405,N_2437);
nor U2633 (N_2633,N_2518,N_2511);
nor U2634 (N_2634,N_2584,N_2420);
or U2635 (N_2635,N_2425,N_2546);
nand U2636 (N_2636,N_2411,N_2573);
and U2637 (N_2637,N_2539,N_2577);
or U2638 (N_2638,N_2552,N_2554);
and U2639 (N_2639,N_2571,N_2570);
or U2640 (N_2640,N_2459,N_2467);
nand U2641 (N_2641,N_2568,N_2510);
and U2642 (N_2642,N_2445,N_2555);
nor U2643 (N_2643,N_2561,N_2501);
or U2644 (N_2644,N_2479,N_2448);
and U2645 (N_2645,N_2464,N_2493);
and U2646 (N_2646,N_2442,N_2440);
nor U2647 (N_2647,N_2418,N_2524);
nor U2648 (N_2648,N_2444,N_2478);
nand U2649 (N_2649,N_2497,N_2531);
or U2650 (N_2650,N_2481,N_2413);
nor U2651 (N_2651,N_2406,N_2474);
nor U2652 (N_2652,N_2578,N_2412);
or U2653 (N_2653,N_2416,N_2422);
nand U2654 (N_2654,N_2460,N_2458);
nor U2655 (N_2655,N_2465,N_2548);
nor U2656 (N_2656,N_2534,N_2400);
nand U2657 (N_2657,N_2543,N_2434);
and U2658 (N_2658,N_2597,N_2408);
or U2659 (N_2659,N_2490,N_2402);
or U2660 (N_2660,N_2506,N_2446);
and U2661 (N_2661,N_2532,N_2483);
or U2662 (N_2662,N_2545,N_2590);
xor U2663 (N_2663,N_2482,N_2492);
nand U2664 (N_2664,N_2550,N_2419);
and U2665 (N_2665,N_2443,N_2551);
and U2666 (N_2666,N_2453,N_2591);
nand U2667 (N_2667,N_2489,N_2556);
nor U2668 (N_2668,N_2509,N_2484);
nand U2669 (N_2669,N_2579,N_2476);
nor U2670 (N_2670,N_2426,N_2572);
nand U2671 (N_2671,N_2581,N_2541);
or U2672 (N_2672,N_2433,N_2470);
and U2673 (N_2673,N_2566,N_2477);
and U2674 (N_2674,N_2471,N_2508);
and U2675 (N_2675,N_2435,N_2583);
and U2676 (N_2676,N_2424,N_2449);
or U2677 (N_2677,N_2432,N_2574);
xnor U2678 (N_2678,N_2441,N_2480);
and U2679 (N_2679,N_2450,N_2525);
xor U2680 (N_2680,N_2451,N_2530);
nor U2681 (N_2681,N_2468,N_2427);
nand U2682 (N_2682,N_2567,N_2588);
or U2683 (N_2683,N_2428,N_2421);
and U2684 (N_2684,N_2429,N_2596);
and U2685 (N_2685,N_2404,N_2582);
and U2686 (N_2686,N_2439,N_2569);
nor U2687 (N_2687,N_2563,N_2475);
xor U2688 (N_2688,N_2544,N_2592);
nor U2689 (N_2689,N_2472,N_2560);
or U2690 (N_2690,N_2547,N_2585);
nand U2691 (N_2691,N_2457,N_2407);
nor U2692 (N_2692,N_2558,N_2517);
nand U2693 (N_2693,N_2557,N_2469);
or U2694 (N_2694,N_2542,N_2498);
and U2695 (N_2695,N_2593,N_2512);
nand U2696 (N_2696,N_2535,N_2519);
or U2697 (N_2697,N_2587,N_2507);
nor U2698 (N_2698,N_2436,N_2598);
or U2699 (N_2699,N_2504,N_2516);
nand U2700 (N_2700,N_2537,N_2556);
nor U2701 (N_2701,N_2520,N_2531);
nand U2702 (N_2702,N_2434,N_2420);
nand U2703 (N_2703,N_2423,N_2544);
nor U2704 (N_2704,N_2580,N_2409);
nor U2705 (N_2705,N_2523,N_2517);
nand U2706 (N_2706,N_2591,N_2501);
or U2707 (N_2707,N_2432,N_2524);
and U2708 (N_2708,N_2471,N_2491);
nor U2709 (N_2709,N_2458,N_2415);
or U2710 (N_2710,N_2454,N_2410);
nand U2711 (N_2711,N_2512,N_2423);
or U2712 (N_2712,N_2539,N_2480);
and U2713 (N_2713,N_2493,N_2597);
nand U2714 (N_2714,N_2406,N_2475);
and U2715 (N_2715,N_2596,N_2540);
and U2716 (N_2716,N_2599,N_2558);
nor U2717 (N_2717,N_2509,N_2434);
and U2718 (N_2718,N_2406,N_2493);
nor U2719 (N_2719,N_2453,N_2441);
nor U2720 (N_2720,N_2487,N_2451);
nor U2721 (N_2721,N_2438,N_2580);
or U2722 (N_2722,N_2413,N_2505);
nor U2723 (N_2723,N_2494,N_2580);
and U2724 (N_2724,N_2596,N_2512);
or U2725 (N_2725,N_2584,N_2532);
and U2726 (N_2726,N_2579,N_2495);
or U2727 (N_2727,N_2501,N_2488);
nand U2728 (N_2728,N_2414,N_2403);
nor U2729 (N_2729,N_2417,N_2506);
nor U2730 (N_2730,N_2519,N_2572);
nand U2731 (N_2731,N_2470,N_2496);
nor U2732 (N_2732,N_2444,N_2531);
or U2733 (N_2733,N_2520,N_2538);
nand U2734 (N_2734,N_2470,N_2557);
nand U2735 (N_2735,N_2460,N_2448);
or U2736 (N_2736,N_2564,N_2571);
or U2737 (N_2737,N_2426,N_2436);
nor U2738 (N_2738,N_2478,N_2442);
and U2739 (N_2739,N_2581,N_2437);
nor U2740 (N_2740,N_2439,N_2525);
and U2741 (N_2741,N_2515,N_2436);
nor U2742 (N_2742,N_2416,N_2570);
nand U2743 (N_2743,N_2486,N_2411);
or U2744 (N_2744,N_2542,N_2433);
or U2745 (N_2745,N_2416,N_2455);
nor U2746 (N_2746,N_2541,N_2404);
nor U2747 (N_2747,N_2598,N_2437);
or U2748 (N_2748,N_2518,N_2527);
nand U2749 (N_2749,N_2464,N_2566);
nor U2750 (N_2750,N_2438,N_2494);
and U2751 (N_2751,N_2414,N_2469);
and U2752 (N_2752,N_2510,N_2584);
nor U2753 (N_2753,N_2437,N_2406);
or U2754 (N_2754,N_2515,N_2582);
or U2755 (N_2755,N_2527,N_2489);
or U2756 (N_2756,N_2589,N_2477);
or U2757 (N_2757,N_2436,N_2568);
nor U2758 (N_2758,N_2596,N_2513);
or U2759 (N_2759,N_2536,N_2514);
and U2760 (N_2760,N_2597,N_2480);
nand U2761 (N_2761,N_2411,N_2454);
and U2762 (N_2762,N_2441,N_2425);
nor U2763 (N_2763,N_2576,N_2570);
nand U2764 (N_2764,N_2515,N_2491);
xnor U2765 (N_2765,N_2485,N_2554);
nand U2766 (N_2766,N_2536,N_2412);
and U2767 (N_2767,N_2482,N_2564);
nor U2768 (N_2768,N_2440,N_2471);
nand U2769 (N_2769,N_2423,N_2539);
or U2770 (N_2770,N_2582,N_2446);
nor U2771 (N_2771,N_2414,N_2494);
nand U2772 (N_2772,N_2400,N_2499);
nand U2773 (N_2773,N_2516,N_2465);
nand U2774 (N_2774,N_2403,N_2569);
nand U2775 (N_2775,N_2550,N_2500);
nor U2776 (N_2776,N_2459,N_2537);
nand U2777 (N_2777,N_2456,N_2498);
nor U2778 (N_2778,N_2424,N_2534);
or U2779 (N_2779,N_2417,N_2561);
nand U2780 (N_2780,N_2523,N_2521);
xnor U2781 (N_2781,N_2538,N_2564);
nor U2782 (N_2782,N_2433,N_2405);
or U2783 (N_2783,N_2453,N_2540);
and U2784 (N_2784,N_2491,N_2460);
and U2785 (N_2785,N_2523,N_2447);
or U2786 (N_2786,N_2477,N_2438);
nor U2787 (N_2787,N_2449,N_2558);
and U2788 (N_2788,N_2593,N_2546);
and U2789 (N_2789,N_2430,N_2514);
and U2790 (N_2790,N_2595,N_2581);
xor U2791 (N_2791,N_2540,N_2572);
xor U2792 (N_2792,N_2515,N_2490);
or U2793 (N_2793,N_2418,N_2506);
and U2794 (N_2794,N_2462,N_2520);
nand U2795 (N_2795,N_2514,N_2554);
or U2796 (N_2796,N_2471,N_2497);
and U2797 (N_2797,N_2433,N_2503);
and U2798 (N_2798,N_2482,N_2472);
nand U2799 (N_2799,N_2495,N_2587);
or U2800 (N_2800,N_2603,N_2731);
xnor U2801 (N_2801,N_2625,N_2789);
nor U2802 (N_2802,N_2669,N_2650);
nand U2803 (N_2803,N_2707,N_2788);
nor U2804 (N_2804,N_2649,N_2615);
or U2805 (N_2805,N_2729,N_2609);
nand U2806 (N_2806,N_2613,N_2630);
nand U2807 (N_2807,N_2612,N_2602);
and U2808 (N_2808,N_2755,N_2720);
xor U2809 (N_2809,N_2699,N_2639);
nor U2810 (N_2810,N_2790,N_2620);
or U2811 (N_2811,N_2748,N_2618);
nand U2812 (N_2812,N_2757,N_2715);
and U2813 (N_2813,N_2647,N_2670);
nor U2814 (N_2814,N_2740,N_2698);
nor U2815 (N_2815,N_2733,N_2723);
nor U2816 (N_2816,N_2708,N_2721);
and U2817 (N_2817,N_2724,N_2605);
nand U2818 (N_2818,N_2738,N_2711);
nor U2819 (N_2819,N_2616,N_2750);
and U2820 (N_2820,N_2773,N_2712);
nand U2821 (N_2821,N_2744,N_2680);
nand U2822 (N_2822,N_2716,N_2726);
or U2823 (N_2823,N_2710,N_2795);
and U2824 (N_2824,N_2745,N_2791);
and U2825 (N_2825,N_2656,N_2766);
nor U2826 (N_2826,N_2659,N_2679);
and U2827 (N_2827,N_2737,N_2666);
and U2828 (N_2828,N_2621,N_2633);
nand U2829 (N_2829,N_2651,N_2783);
xnor U2830 (N_2830,N_2663,N_2617);
xnor U2831 (N_2831,N_2759,N_2683);
or U2832 (N_2832,N_2629,N_2754);
and U2833 (N_2833,N_2681,N_2718);
nand U2834 (N_2834,N_2743,N_2652);
or U2835 (N_2835,N_2717,N_2706);
xor U2836 (N_2836,N_2725,N_2760);
or U2837 (N_2837,N_2749,N_2753);
nor U2838 (N_2838,N_2636,N_2662);
nor U2839 (N_2839,N_2746,N_2628);
nand U2840 (N_2840,N_2665,N_2675);
nand U2841 (N_2841,N_2722,N_2688);
and U2842 (N_2842,N_2784,N_2682);
and U2843 (N_2843,N_2769,N_2763);
and U2844 (N_2844,N_2660,N_2781);
or U2845 (N_2845,N_2691,N_2770);
nand U2846 (N_2846,N_2654,N_2768);
nor U2847 (N_2847,N_2735,N_2673);
and U2848 (N_2848,N_2685,N_2661);
and U2849 (N_2849,N_2756,N_2727);
xor U2850 (N_2850,N_2799,N_2728);
or U2851 (N_2851,N_2701,N_2705);
nor U2852 (N_2852,N_2739,N_2765);
nand U2853 (N_2853,N_2657,N_2719);
or U2854 (N_2854,N_2697,N_2794);
nor U2855 (N_2855,N_2751,N_2690);
nand U2856 (N_2856,N_2645,N_2774);
nor U2857 (N_2857,N_2796,N_2792);
or U2858 (N_2858,N_2736,N_2704);
nand U2859 (N_2859,N_2668,N_2703);
and U2860 (N_2860,N_2742,N_2692);
and U2861 (N_2861,N_2655,N_2786);
nand U2862 (N_2862,N_2785,N_2611);
and U2863 (N_2863,N_2624,N_2653);
nand U2864 (N_2864,N_2713,N_2696);
and U2865 (N_2865,N_2644,N_2677);
or U2866 (N_2866,N_2782,N_2664);
and U2867 (N_2867,N_2637,N_2762);
nor U2868 (N_2868,N_2604,N_2600);
nand U2869 (N_2869,N_2787,N_2709);
or U2870 (N_2870,N_2632,N_2752);
and U2871 (N_2871,N_2608,N_2777);
nand U2872 (N_2872,N_2635,N_2747);
nand U2873 (N_2873,N_2658,N_2674);
and U2874 (N_2874,N_2642,N_2778);
and U2875 (N_2875,N_2693,N_2610);
or U2876 (N_2876,N_2672,N_2671);
or U2877 (N_2877,N_2614,N_2676);
xor U2878 (N_2878,N_2732,N_2695);
or U2879 (N_2879,N_2775,N_2684);
xor U2880 (N_2880,N_2689,N_2702);
or U2881 (N_2881,N_2601,N_2678);
or U2882 (N_2882,N_2730,N_2758);
and U2883 (N_2883,N_2779,N_2619);
and U2884 (N_2884,N_2714,N_2631);
nor U2885 (N_2885,N_2793,N_2626);
and U2886 (N_2886,N_2798,N_2771);
nand U2887 (N_2887,N_2634,N_2640);
and U2888 (N_2888,N_2622,N_2687);
and U2889 (N_2889,N_2646,N_2767);
and U2890 (N_2890,N_2606,N_2607);
nand U2891 (N_2891,N_2641,N_2667);
nor U2892 (N_2892,N_2700,N_2638);
and U2893 (N_2893,N_2686,N_2643);
nor U2894 (N_2894,N_2741,N_2627);
or U2895 (N_2895,N_2776,N_2764);
nand U2896 (N_2896,N_2734,N_2772);
xor U2897 (N_2897,N_2648,N_2694);
nor U2898 (N_2898,N_2780,N_2761);
and U2899 (N_2899,N_2797,N_2623);
nor U2900 (N_2900,N_2637,N_2635);
or U2901 (N_2901,N_2636,N_2718);
or U2902 (N_2902,N_2755,N_2733);
nand U2903 (N_2903,N_2656,N_2640);
nor U2904 (N_2904,N_2748,N_2789);
nor U2905 (N_2905,N_2647,N_2672);
nand U2906 (N_2906,N_2708,N_2737);
or U2907 (N_2907,N_2769,N_2627);
or U2908 (N_2908,N_2626,N_2797);
and U2909 (N_2909,N_2696,N_2790);
nor U2910 (N_2910,N_2664,N_2742);
nor U2911 (N_2911,N_2756,N_2726);
nand U2912 (N_2912,N_2769,N_2661);
nor U2913 (N_2913,N_2742,N_2796);
nor U2914 (N_2914,N_2788,N_2625);
or U2915 (N_2915,N_2734,N_2768);
and U2916 (N_2916,N_2646,N_2626);
xor U2917 (N_2917,N_2644,N_2742);
nand U2918 (N_2918,N_2797,N_2739);
nand U2919 (N_2919,N_2695,N_2758);
or U2920 (N_2920,N_2677,N_2788);
nor U2921 (N_2921,N_2774,N_2622);
or U2922 (N_2922,N_2693,N_2676);
or U2923 (N_2923,N_2644,N_2791);
and U2924 (N_2924,N_2794,N_2720);
or U2925 (N_2925,N_2609,N_2797);
nand U2926 (N_2926,N_2784,N_2640);
nand U2927 (N_2927,N_2625,N_2657);
or U2928 (N_2928,N_2787,N_2770);
or U2929 (N_2929,N_2689,N_2792);
nand U2930 (N_2930,N_2766,N_2720);
and U2931 (N_2931,N_2685,N_2606);
or U2932 (N_2932,N_2784,N_2630);
and U2933 (N_2933,N_2722,N_2674);
xnor U2934 (N_2934,N_2633,N_2660);
or U2935 (N_2935,N_2729,N_2682);
and U2936 (N_2936,N_2691,N_2632);
and U2937 (N_2937,N_2616,N_2608);
nand U2938 (N_2938,N_2706,N_2644);
nor U2939 (N_2939,N_2767,N_2790);
and U2940 (N_2940,N_2629,N_2710);
nand U2941 (N_2941,N_2788,N_2675);
nand U2942 (N_2942,N_2645,N_2784);
and U2943 (N_2943,N_2665,N_2645);
and U2944 (N_2944,N_2735,N_2688);
xor U2945 (N_2945,N_2609,N_2606);
nand U2946 (N_2946,N_2742,N_2695);
and U2947 (N_2947,N_2672,N_2630);
or U2948 (N_2948,N_2646,N_2608);
and U2949 (N_2949,N_2663,N_2630);
nor U2950 (N_2950,N_2681,N_2690);
and U2951 (N_2951,N_2681,N_2675);
or U2952 (N_2952,N_2723,N_2690);
and U2953 (N_2953,N_2791,N_2637);
xor U2954 (N_2954,N_2719,N_2778);
nand U2955 (N_2955,N_2786,N_2602);
and U2956 (N_2956,N_2736,N_2652);
xor U2957 (N_2957,N_2776,N_2624);
xor U2958 (N_2958,N_2785,N_2633);
nor U2959 (N_2959,N_2691,N_2766);
nor U2960 (N_2960,N_2710,N_2681);
xnor U2961 (N_2961,N_2693,N_2631);
or U2962 (N_2962,N_2760,N_2793);
or U2963 (N_2963,N_2745,N_2690);
xor U2964 (N_2964,N_2676,N_2792);
or U2965 (N_2965,N_2794,N_2760);
or U2966 (N_2966,N_2779,N_2756);
nor U2967 (N_2967,N_2719,N_2770);
nor U2968 (N_2968,N_2777,N_2767);
nand U2969 (N_2969,N_2736,N_2606);
and U2970 (N_2970,N_2698,N_2604);
nand U2971 (N_2971,N_2716,N_2776);
and U2972 (N_2972,N_2600,N_2669);
nand U2973 (N_2973,N_2779,N_2637);
and U2974 (N_2974,N_2775,N_2720);
nand U2975 (N_2975,N_2772,N_2782);
or U2976 (N_2976,N_2726,N_2739);
nor U2977 (N_2977,N_2798,N_2620);
or U2978 (N_2978,N_2701,N_2699);
nor U2979 (N_2979,N_2602,N_2756);
and U2980 (N_2980,N_2758,N_2778);
nand U2981 (N_2981,N_2734,N_2756);
nor U2982 (N_2982,N_2745,N_2613);
or U2983 (N_2983,N_2682,N_2636);
or U2984 (N_2984,N_2666,N_2709);
or U2985 (N_2985,N_2661,N_2607);
nor U2986 (N_2986,N_2734,N_2716);
nand U2987 (N_2987,N_2747,N_2783);
or U2988 (N_2988,N_2621,N_2687);
xor U2989 (N_2989,N_2684,N_2759);
xnor U2990 (N_2990,N_2676,N_2627);
or U2991 (N_2991,N_2748,N_2706);
and U2992 (N_2992,N_2707,N_2735);
nand U2993 (N_2993,N_2626,N_2684);
nor U2994 (N_2994,N_2711,N_2790);
xor U2995 (N_2995,N_2777,N_2631);
nand U2996 (N_2996,N_2703,N_2669);
and U2997 (N_2997,N_2713,N_2727);
nand U2998 (N_2998,N_2691,N_2762);
xor U2999 (N_2999,N_2609,N_2751);
and U3000 (N_3000,N_2867,N_2831);
nor U3001 (N_3001,N_2843,N_2824);
and U3002 (N_3002,N_2809,N_2922);
and U3003 (N_3003,N_2845,N_2817);
nor U3004 (N_3004,N_2820,N_2929);
nor U3005 (N_3005,N_2814,N_2996);
nand U3006 (N_3006,N_2813,N_2846);
nand U3007 (N_3007,N_2851,N_2837);
nor U3008 (N_3008,N_2967,N_2894);
nor U3009 (N_3009,N_2821,N_2947);
nand U3010 (N_3010,N_2892,N_2963);
nor U3011 (N_3011,N_2960,N_2966);
nor U3012 (N_3012,N_2871,N_2870);
or U3013 (N_3013,N_2921,N_2827);
nor U3014 (N_3014,N_2826,N_2957);
or U3015 (N_3015,N_2991,N_2898);
and U3016 (N_3016,N_2932,N_2866);
and U3017 (N_3017,N_2900,N_2984);
or U3018 (N_3018,N_2863,N_2876);
nor U3019 (N_3019,N_2971,N_2927);
xor U3020 (N_3020,N_2816,N_2990);
nor U3021 (N_3021,N_2834,N_2942);
xor U3022 (N_3022,N_2858,N_2958);
and U3023 (N_3023,N_2974,N_2877);
and U3024 (N_3024,N_2987,N_2986);
or U3025 (N_3025,N_2811,N_2976);
nor U3026 (N_3026,N_2950,N_2935);
or U3027 (N_3027,N_2838,N_2807);
nand U3028 (N_3028,N_2829,N_2856);
xor U3029 (N_3029,N_2994,N_2940);
nor U3030 (N_3030,N_2885,N_2879);
or U3031 (N_3031,N_2939,N_2938);
or U3032 (N_3032,N_2931,N_2890);
xor U3033 (N_3033,N_2906,N_2916);
xor U3034 (N_3034,N_2982,N_2886);
nand U3035 (N_3035,N_2860,N_2859);
and U3036 (N_3036,N_2954,N_2944);
xnor U3037 (N_3037,N_2806,N_2969);
nand U3038 (N_3038,N_2936,N_2904);
xor U3039 (N_3039,N_2854,N_2887);
nand U3040 (N_3040,N_2881,N_2853);
or U3041 (N_3041,N_2993,N_2998);
or U3042 (N_3042,N_2897,N_2839);
nand U3043 (N_3043,N_2874,N_2878);
nand U3044 (N_3044,N_2920,N_2889);
xnor U3045 (N_3045,N_2861,N_2835);
and U3046 (N_3046,N_2842,N_2872);
and U3047 (N_3047,N_2907,N_2905);
and U3048 (N_3048,N_2822,N_2955);
and U3049 (N_3049,N_2902,N_2959);
or U3050 (N_3050,N_2836,N_2924);
nor U3051 (N_3051,N_2961,N_2995);
xnor U3052 (N_3052,N_2808,N_2801);
nor U3053 (N_3053,N_2926,N_2825);
nand U3054 (N_3054,N_2802,N_2883);
and U3055 (N_3055,N_2953,N_2970);
or U3056 (N_3056,N_2864,N_2919);
and U3057 (N_3057,N_2997,N_2999);
or U3058 (N_3058,N_2981,N_2855);
or U3059 (N_3059,N_2928,N_2800);
nor U3060 (N_3060,N_2830,N_2896);
and U3061 (N_3061,N_2880,N_2891);
nor U3062 (N_3062,N_2983,N_2934);
nand U3063 (N_3063,N_2895,N_2930);
and U3064 (N_3064,N_2828,N_2818);
or U3065 (N_3065,N_2917,N_2979);
nand U3066 (N_3066,N_2968,N_2943);
nor U3067 (N_3067,N_2952,N_2908);
or U3068 (N_3068,N_2918,N_2914);
and U3069 (N_3069,N_2803,N_2847);
nand U3070 (N_3070,N_2949,N_2875);
nor U3071 (N_3071,N_2812,N_2850);
nand U3072 (N_3072,N_2980,N_2819);
nand U3073 (N_3073,N_2910,N_2862);
or U3074 (N_3074,N_2988,N_2840);
and U3075 (N_3075,N_2815,N_2868);
nand U3076 (N_3076,N_2989,N_2978);
nor U3077 (N_3077,N_2882,N_2956);
nor U3078 (N_3078,N_2972,N_2884);
and U3079 (N_3079,N_2823,N_2912);
and U3080 (N_3080,N_2911,N_2962);
nand U3081 (N_3081,N_2909,N_2888);
nor U3082 (N_3082,N_2893,N_2946);
or U3083 (N_3083,N_2841,N_2948);
nand U3084 (N_3084,N_2833,N_2869);
or U3085 (N_3085,N_2873,N_2832);
xnor U3086 (N_3086,N_2985,N_2915);
or U3087 (N_3087,N_2899,N_2977);
or U3088 (N_3088,N_2810,N_2913);
and U3089 (N_3089,N_2937,N_2975);
nor U3090 (N_3090,N_2805,N_2848);
nor U3091 (N_3091,N_2973,N_2945);
and U3092 (N_3092,N_2925,N_2965);
nor U3093 (N_3093,N_2941,N_2951);
nand U3094 (N_3094,N_2804,N_2865);
or U3095 (N_3095,N_2923,N_2852);
or U3096 (N_3096,N_2901,N_2857);
nor U3097 (N_3097,N_2964,N_2992);
nand U3098 (N_3098,N_2933,N_2903);
nand U3099 (N_3099,N_2849,N_2844);
xor U3100 (N_3100,N_2944,N_2833);
or U3101 (N_3101,N_2952,N_2827);
or U3102 (N_3102,N_2815,N_2916);
and U3103 (N_3103,N_2991,N_2899);
and U3104 (N_3104,N_2970,N_2841);
nand U3105 (N_3105,N_2948,N_2987);
nor U3106 (N_3106,N_2961,N_2990);
nor U3107 (N_3107,N_2957,N_2933);
or U3108 (N_3108,N_2809,N_2970);
or U3109 (N_3109,N_2822,N_2829);
and U3110 (N_3110,N_2916,N_2865);
nor U3111 (N_3111,N_2941,N_2888);
nor U3112 (N_3112,N_2929,N_2837);
and U3113 (N_3113,N_2809,N_2932);
or U3114 (N_3114,N_2904,N_2864);
or U3115 (N_3115,N_2937,N_2812);
nand U3116 (N_3116,N_2943,N_2921);
nor U3117 (N_3117,N_2949,N_2982);
or U3118 (N_3118,N_2923,N_2814);
and U3119 (N_3119,N_2851,N_2801);
or U3120 (N_3120,N_2905,N_2972);
and U3121 (N_3121,N_2831,N_2883);
or U3122 (N_3122,N_2826,N_2948);
or U3123 (N_3123,N_2854,N_2986);
or U3124 (N_3124,N_2924,N_2811);
nand U3125 (N_3125,N_2826,N_2802);
nand U3126 (N_3126,N_2899,N_2937);
or U3127 (N_3127,N_2975,N_2815);
and U3128 (N_3128,N_2845,N_2982);
xor U3129 (N_3129,N_2912,N_2881);
nor U3130 (N_3130,N_2800,N_2994);
xor U3131 (N_3131,N_2945,N_2977);
xor U3132 (N_3132,N_2832,N_2994);
nand U3133 (N_3133,N_2897,N_2991);
or U3134 (N_3134,N_2855,N_2871);
and U3135 (N_3135,N_2822,N_2885);
and U3136 (N_3136,N_2945,N_2867);
nand U3137 (N_3137,N_2888,N_2871);
or U3138 (N_3138,N_2976,N_2822);
nand U3139 (N_3139,N_2807,N_2841);
nand U3140 (N_3140,N_2913,N_2988);
xnor U3141 (N_3141,N_2808,N_2972);
nand U3142 (N_3142,N_2998,N_2937);
nand U3143 (N_3143,N_2808,N_2849);
and U3144 (N_3144,N_2870,N_2917);
and U3145 (N_3145,N_2884,N_2983);
nand U3146 (N_3146,N_2816,N_2857);
and U3147 (N_3147,N_2880,N_2823);
or U3148 (N_3148,N_2925,N_2967);
and U3149 (N_3149,N_2841,N_2855);
nand U3150 (N_3150,N_2929,N_2885);
nor U3151 (N_3151,N_2929,N_2821);
nor U3152 (N_3152,N_2823,N_2967);
nand U3153 (N_3153,N_2932,N_2834);
nand U3154 (N_3154,N_2934,N_2999);
nand U3155 (N_3155,N_2911,N_2902);
nor U3156 (N_3156,N_2885,N_2882);
nand U3157 (N_3157,N_2970,N_2964);
nand U3158 (N_3158,N_2802,N_2913);
or U3159 (N_3159,N_2964,N_2940);
nor U3160 (N_3160,N_2976,N_2828);
or U3161 (N_3161,N_2911,N_2888);
nor U3162 (N_3162,N_2819,N_2821);
or U3163 (N_3163,N_2879,N_2849);
and U3164 (N_3164,N_2960,N_2921);
nor U3165 (N_3165,N_2828,N_2853);
nand U3166 (N_3166,N_2953,N_2851);
or U3167 (N_3167,N_2939,N_2840);
and U3168 (N_3168,N_2838,N_2820);
or U3169 (N_3169,N_2840,N_2805);
or U3170 (N_3170,N_2803,N_2895);
and U3171 (N_3171,N_2992,N_2833);
and U3172 (N_3172,N_2899,N_2929);
nor U3173 (N_3173,N_2954,N_2931);
xor U3174 (N_3174,N_2860,N_2883);
nand U3175 (N_3175,N_2888,N_2814);
xnor U3176 (N_3176,N_2840,N_2994);
and U3177 (N_3177,N_2928,N_2936);
and U3178 (N_3178,N_2951,N_2894);
nor U3179 (N_3179,N_2985,N_2824);
nand U3180 (N_3180,N_2982,N_2995);
nand U3181 (N_3181,N_2829,N_2930);
xor U3182 (N_3182,N_2901,N_2902);
nor U3183 (N_3183,N_2993,N_2886);
nor U3184 (N_3184,N_2857,N_2973);
or U3185 (N_3185,N_2917,N_2850);
nand U3186 (N_3186,N_2835,N_2883);
and U3187 (N_3187,N_2923,N_2843);
nand U3188 (N_3188,N_2941,N_2926);
nor U3189 (N_3189,N_2916,N_2983);
or U3190 (N_3190,N_2906,N_2808);
nor U3191 (N_3191,N_2906,N_2873);
and U3192 (N_3192,N_2897,N_2818);
and U3193 (N_3193,N_2836,N_2815);
nor U3194 (N_3194,N_2844,N_2925);
and U3195 (N_3195,N_2802,N_2876);
and U3196 (N_3196,N_2819,N_2941);
xor U3197 (N_3197,N_2916,N_2827);
nor U3198 (N_3198,N_2858,N_2944);
nor U3199 (N_3199,N_2891,N_2817);
nor U3200 (N_3200,N_3028,N_3060);
and U3201 (N_3201,N_3024,N_3166);
nand U3202 (N_3202,N_3196,N_3186);
or U3203 (N_3203,N_3089,N_3106);
and U3204 (N_3204,N_3093,N_3088);
or U3205 (N_3205,N_3127,N_3039);
nand U3206 (N_3206,N_3094,N_3040);
or U3207 (N_3207,N_3097,N_3072);
nand U3208 (N_3208,N_3171,N_3055);
and U3209 (N_3209,N_3120,N_3095);
nor U3210 (N_3210,N_3063,N_3101);
or U3211 (N_3211,N_3012,N_3001);
nand U3212 (N_3212,N_3085,N_3168);
or U3213 (N_3213,N_3102,N_3086);
and U3214 (N_3214,N_3169,N_3020);
and U3215 (N_3215,N_3013,N_3172);
or U3216 (N_3216,N_3140,N_3021);
or U3217 (N_3217,N_3008,N_3135);
nand U3218 (N_3218,N_3134,N_3192);
and U3219 (N_3219,N_3098,N_3049);
nand U3220 (N_3220,N_3058,N_3099);
or U3221 (N_3221,N_3109,N_3051);
and U3222 (N_3222,N_3133,N_3184);
nor U3223 (N_3223,N_3119,N_3046);
nand U3224 (N_3224,N_3175,N_3074);
and U3225 (N_3225,N_3123,N_3079);
and U3226 (N_3226,N_3103,N_3062);
xnor U3227 (N_3227,N_3173,N_3083);
or U3228 (N_3228,N_3047,N_3026);
or U3229 (N_3229,N_3003,N_3155);
or U3230 (N_3230,N_3188,N_3193);
and U3231 (N_3231,N_3147,N_3068);
or U3232 (N_3232,N_3152,N_3071);
nor U3233 (N_3233,N_3032,N_3125);
and U3234 (N_3234,N_3131,N_3017);
xnor U3235 (N_3235,N_3112,N_3004);
nor U3236 (N_3236,N_3191,N_3044);
nor U3237 (N_3237,N_3042,N_3023);
nand U3238 (N_3238,N_3041,N_3078);
or U3239 (N_3239,N_3035,N_3170);
or U3240 (N_3240,N_3136,N_3164);
nor U3241 (N_3241,N_3077,N_3050);
or U3242 (N_3242,N_3163,N_3111);
and U3243 (N_3243,N_3145,N_3069);
nand U3244 (N_3244,N_3038,N_3137);
and U3245 (N_3245,N_3081,N_3199);
nor U3246 (N_3246,N_3174,N_3197);
nand U3247 (N_3247,N_3104,N_3151);
and U3248 (N_3248,N_3052,N_3000);
nor U3249 (N_3249,N_3198,N_3065);
or U3250 (N_3250,N_3146,N_3031);
nand U3251 (N_3251,N_3064,N_3033);
nand U3252 (N_3252,N_3084,N_3130);
nor U3253 (N_3253,N_3181,N_3156);
nand U3254 (N_3254,N_3053,N_3105);
and U3255 (N_3255,N_3179,N_3080);
nor U3256 (N_3256,N_3148,N_3182);
nand U3257 (N_3257,N_3185,N_3061);
nand U3258 (N_3258,N_3150,N_3177);
nor U3259 (N_3259,N_3019,N_3154);
nor U3260 (N_3260,N_3159,N_3195);
or U3261 (N_3261,N_3167,N_3036);
xnor U3262 (N_3262,N_3029,N_3121);
or U3263 (N_3263,N_3025,N_3030);
nor U3264 (N_3264,N_3022,N_3027);
or U3265 (N_3265,N_3189,N_3011);
or U3266 (N_3266,N_3082,N_3190);
nor U3267 (N_3267,N_3034,N_3009);
and U3268 (N_3268,N_3160,N_3005);
nand U3269 (N_3269,N_3092,N_3157);
and U3270 (N_3270,N_3116,N_3070);
nand U3271 (N_3271,N_3183,N_3124);
xnor U3272 (N_3272,N_3144,N_3141);
and U3273 (N_3273,N_3126,N_3162);
and U3274 (N_3274,N_3045,N_3073);
nand U3275 (N_3275,N_3096,N_3114);
or U3276 (N_3276,N_3100,N_3118);
nand U3277 (N_3277,N_3129,N_3067);
nand U3278 (N_3278,N_3007,N_3091);
nand U3279 (N_3279,N_3016,N_3138);
or U3280 (N_3280,N_3132,N_3054);
nor U3281 (N_3281,N_3194,N_3180);
or U3282 (N_3282,N_3165,N_3113);
nand U3283 (N_3283,N_3117,N_3110);
and U3284 (N_3284,N_3018,N_3014);
xnor U3285 (N_3285,N_3059,N_3108);
or U3286 (N_3286,N_3056,N_3187);
or U3287 (N_3287,N_3178,N_3010);
nand U3288 (N_3288,N_3087,N_3139);
nor U3289 (N_3289,N_3043,N_3143);
xnor U3290 (N_3290,N_3090,N_3122);
nor U3291 (N_3291,N_3115,N_3037);
nor U3292 (N_3292,N_3161,N_3142);
nor U3293 (N_3293,N_3153,N_3107);
nor U3294 (N_3294,N_3002,N_3066);
and U3295 (N_3295,N_3128,N_3075);
or U3296 (N_3296,N_3076,N_3149);
nor U3297 (N_3297,N_3057,N_3176);
or U3298 (N_3298,N_3158,N_3006);
or U3299 (N_3299,N_3048,N_3015);
nor U3300 (N_3300,N_3149,N_3053);
and U3301 (N_3301,N_3066,N_3059);
xnor U3302 (N_3302,N_3042,N_3016);
and U3303 (N_3303,N_3168,N_3134);
xor U3304 (N_3304,N_3028,N_3111);
or U3305 (N_3305,N_3143,N_3162);
nand U3306 (N_3306,N_3016,N_3150);
nand U3307 (N_3307,N_3160,N_3029);
nand U3308 (N_3308,N_3084,N_3046);
nand U3309 (N_3309,N_3079,N_3080);
nor U3310 (N_3310,N_3169,N_3093);
and U3311 (N_3311,N_3186,N_3175);
nor U3312 (N_3312,N_3163,N_3115);
nand U3313 (N_3313,N_3041,N_3046);
nand U3314 (N_3314,N_3021,N_3152);
or U3315 (N_3315,N_3149,N_3061);
nor U3316 (N_3316,N_3022,N_3104);
xor U3317 (N_3317,N_3107,N_3056);
and U3318 (N_3318,N_3031,N_3105);
or U3319 (N_3319,N_3123,N_3034);
and U3320 (N_3320,N_3084,N_3110);
or U3321 (N_3321,N_3199,N_3153);
or U3322 (N_3322,N_3063,N_3081);
or U3323 (N_3323,N_3068,N_3101);
or U3324 (N_3324,N_3029,N_3027);
nor U3325 (N_3325,N_3149,N_3089);
and U3326 (N_3326,N_3172,N_3139);
nor U3327 (N_3327,N_3139,N_3143);
xnor U3328 (N_3328,N_3091,N_3146);
xnor U3329 (N_3329,N_3124,N_3012);
nor U3330 (N_3330,N_3101,N_3170);
nor U3331 (N_3331,N_3017,N_3147);
or U3332 (N_3332,N_3147,N_3010);
nor U3333 (N_3333,N_3072,N_3112);
nor U3334 (N_3334,N_3034,N_3096);
nand U3335 (N_3335,N_3084,N_3138);
nor U3336 (N_3336,N_3196,N_3160);
and U3337 (N_3337,N_3168,N_3035);
or U3338 (N_3338,N_3068,N_3080);
or U3339 (N_3339,N_3069,N_3048);
or U3340 (N_3340,N_3123,N_3169);
or U3341 (N_3341,N_3019,N_3002);
and U3342 (N_3342,N_3044,N_3094);
nand U3343 (N_3343,N_3022,N_3167);
nand U3344 (N_3344,N_3160,N_3165);
xor U3345 (N_3345,N_3062,N_3149);
xnor U3346 (N_3346,N_3104,N_3189);
xor U3347 (N_3347,N_3135,N_3041);
xnor U3348 (N_3348,N_3149,N_3136);
and U3349 (N_3349,N_3034,N_3079);
nand U3350 (N_3350,N_3164,N_3184);
and U3351 (N_3351,N_3058,N_3028);
nand U3352 (N_3352,N_3148,N_3086);
nor U3353 (N_3353,N_3046,N_3168);
and U3354 (N_3354,N_3005,N_3105);
or U3355 (N_3355,N_3164,N_3143);
nor U3356 (N_3356,N_3129,N_3173);
nand U3357 (N_3357,N_3091,N_3070);
and U3358 (N_3358,N_3194,N_3022);
xor U3359 (N_3359,N_3058,N_3192);
nor U3360 (N_3360,N_3189,N_3109);
nor U3361 (N_3361,N_3120,N_3026);
nor U3362 (N_3362,N_3114,N_3104);
or U3363 (N_3363,N_3058,N_3055);
xnor U3364 (N_3364,N_3017,N_3173);
nand U3365 (N_3365,N_3008,N_3180);
nand U3366 (N_3366,N_3137,N_3032);
nor U3367 (N_3367,N_3197,N_3026);
or U3368 (N_3368,N_3184,N_3196);
and U3369 (N_3369,N_3147,N_3047);
nor U3370 (N_3370,N_3051,N_3156);
nor U3371 (N_3371,N_3000,N_3015);
nand U3372 (N_3372,N_3143,N_3090);
and U3373 (N_3373,N_3032,N_3105);
or U3374 (N_3374,N_3196,N_3038);
nor U3375 (N_3375,N_3146,N_3015);
nand U3376 (N_3376,N_3128,N_3028);
and U3377 (N_3377,N_3077,N_3122);
nor U3378 (N_3378,N_3019,N_3158);
and U3379 (N_3379,N_3139,N_3157);
nand U3380 (N_3380,N_3194,N_3065);
or U3381 (N_3381,N_3053,N_3125);
and U3382 (N_3382,N_3059,N_3187);
nor U3383 (N_3383,N_3070,N_3111);
nor U3384 (N_3384,N_3049,N_3160);
nor U3385 (N_3385,N_3185,N_3121);
nor U3386 (N_3386,N_3118,N_3193);
nor U3387 (N_3387,N_3000,N_3149);
nand U3388 (N_3388,N_3173,N_3151);
xnor U3389 (N_3389,N_3157,N_3019);
xnor U3390 (N_3390,N_3041,N_3065);
and U3391 (N_3391,N_3003,N_3005);
nand U3392 (N_3392,N_3030,N_3034);
xnor U3393 (N_3393,N_3152,N_3150);
nand U3394 (N_3394,N_3078,N_3056);
or U3395 (N_3395,N_3062,N_3058);
nand U3396 (N_3396,N_3061,N_3152);
nand U3397 (N_3397,N_3090,N_3015);
and U3398 (N_3398,N_3181,N_3025);
xor U3399 (N_3399,N_3152,N_3139);
or U3400 (N_3400,N_3324,N_3313);
nand U3401 (N_3401,N_3210,N_3302);
nand U3402 (N_3402,N_3222,N_3247);
or U3403 (N_3403,N_3328,N_3248);
nand U3404 (N_3404,N_3217,N_3297);
nor U3405 (N_3405,N_3218,N_3293);
nand U3406 (N_3406,N_3212,N_3318);
or U3407 (N_3407,N_3334,N_3374);
nand U3408 (N_3408,N_3332,N_3370);
and U3409 (N_3409,N_3269,N_3389);
and U3410 (N_3410,N_3258,N_3200);
and U3411 (N_3411,N_3230,N_3335);
nand U3412 (N_3412,N_3268,N_3331);
or U3413 (N_3413,N_3382,N_3301);
and U3414 (N_3414,N_3254,N_3341);
and U3415 (N_3415,N_3385,N_3311);
xor U3416 (N_3416,N_3315,N_3252);
nor U3417 (N_3417,N_3323,N_3359);
or U3418 (N_3418,N_3241,N_3291);
nor U3419 (N_3419,N_3215,N_3392);
nand U3420 (N_3420,N_3285,N_3366);
and U3421 (N_3421,N_3321,N_3387);
nor U3422 (N_3422,N_3242,N_3263);
and U3423 (N_3423,N_3279,N_3208);
and U3424 (N_3424,N_3253,N_3375);
and U3425 (N_3425,N_3283,N_3317);
and U3426 (N_3426,N_3362,N_3209);
nand U3427 (N_3427,N_3314,N_3277);
nor U3428 (N_3428,N_3342,N_3272);
and U3429 (N_3429,N_3207,N_3245);
nor U3430 (N_3430,N_3356,N_3264);
nand U3431 (N_3431,N_3244,N_3221);
or U3432 (N_3432,N_3363,N_3201);
and U3433 (N_3433,N_3224,N_3265);
nor U3434 (N_3434,N_3303,N_3288);
nor U3435 (N_3435,N_3239,N_3394);
nor U3436 (N_3436,N_3286,N_3231);
or U3437 (N_3437,N_3205,N_3300);
nor U3438 (N_3438,N_3262,N_3275);
nand U3439 (N_3439,N_3371,N_3384);
and U3440 (N_3440,N_3232,N_3347);
or U3441 (N_3441,N_3353,N_3310);
or U3442 (N_3442,N_3271,N_3284);
and U3443 (N_3443,N_3233,N_3227);
nor U3444 (N_3444,N_3278,N_3383);
or U3445 (N_3445,N_3266,N_3337);
and U3446 (N_3446,N_3348,N_3397);
and U3447 (N_3447,N_3364,N_3344);
nand U3448 (N_3448,N_3270,N_3246);
nand U3449 (N_3449,N_3309,N_3307);
xnor U3450 (N_3450,N_3280,N_3259);
nand U3451 (N_3451,N_3296,N_3249);
and U3452 (N_3452,N_3290,N_3398);
nand U3453 (N_3453,N_3237,N_3206);
or U3454 (N_3454,N_3260,N_3261);
and U3455 (N_3455,N_3308,N_3346);
and U3456 (N_3456,N_3257,N_3330);
xor U3457 (N_3457,N_3326,N_3343);
nor U3458 (N_3458,N_3267,N_3395);
xor U3459 (N_3459,N_3325,N_3372);
or U3460 (N_3460,N_3322,N_3281);
nor U3461 (N_3461,N_3204,N_3329);
and U3462 (N_3462,N_3352,N_3391);
and U3463 (N_3463,N_3214,N_3225);
nand U3464 (N_3464,N_3350,N_3319);
and U3465 (N_3465,N_3388,N_3333);
or U3466 (N_3466,N_3360,N_3379);
nor U3467 (N_3467,N_3213,N_3234);
xnor U3468 (N_3468,N_3377,N_3336);
and U3469 (N_3469,N_3236,N_3380);
and U3470 (N_3470,N_3273,N_3390);
and U3471 (N_3471,N_3312,N_3304);
or U3472 (N_3472,N_3282,N_3396);
nand U3473 (N_3473,N_3276,N_3351);
and U3474 (N_3474,N_3339,N_3289);
nand U3475 (N_3475,N_3367,N_3358);
or U3476 (N_3476,N_3294,N_3228);
nor U3477 (N_3477,N_3295,N_3373);
nor U3478 (N_3478,N_3251,N_3256);
nor U3479 (N_3479,N_3211,N_3355);
or U3480 (N_3480,N_3378,N_3365);
and U3481 (N_3481,N_3349,N_3229);
or U3482 (N_3482,N_3235,N_3274);
and U3483 (N_3483,N_3238,N_3345);
nand U3484 (N_3484,N_3393,N_3250);
and U3485 (N_3485,N_3386,N_3223);
or U3486 (N_3486,N_3203,N_3219);
nor U3487 (N_3487,N_3240,N_3255);
and U3488 (N_3488,N_3287,N_3292);
nand U3489 (N_3489,N_3340,N_3226);
nand U3490 (N_3490,N_3216,N_3354);
or U3491 (N_3491,N_3243,N_3202);
nand U3492 (N_3492,N_3320,N_3369);
or U3493 (N_3493,N_3368,N_3298);
and U3494 (N_3494,N_3327,N_3299);
or U3495 (N_3495,N_3338,N_3220);
and U3496 (N_3496,N_3376,N_3306);
and U3497 (N_3497,N_3399,N_3305);
or U3498 (N_3498,N_3316,N_3357);
xnor U3499 (N_3499,N_3361,N_3381);
or U3500 (N_3500,N_3322,N_3348);
nand U3501 (N_3501,N_3201,N_3337);
and U3502 (N_3502,N_3225,N_3317);
nand U3503 (N_3503,N_3337,N_3270);
nand U3504 (N_3504,N_3255,N_3371);
nor U3505 (N_3505,N_3387,N_3204);
nand U3506 (N_3506,N_3337,N_3239);
nand U3507 (N_3507,N_3383,N_3390);
and U3508 (N_3508,N_3398,N_3305);
or U3509 (N_3509,N_3284,N_3273);
and U3510 (N_3510,N_3243,N_3382);
xnor U3511 (N_3511,N_3290,N_3246);
nor U3512 (N_3512,N_3324,N_3306);
nor U3513 (N_3513,N_3343,N_3342);
or U3514 (N_3514,N_3220,N_3353);
and U3515 (N_3515,N_3260,N_3380);
nor U3516 (N_3516,N_3219,N_3305);
nor U3517 (N_3517,N_3220,N_3385);
or U3518 (N_3518,N_3204,N_3206);
and U3519 (N_3519,N_3352,N_3220);
nand U3520 (N_3520,N_3230,N_3208);
or U3521 (N_3521,N_3310,N_3363);
and U3522 (N_3522,N_3286,N_3363);
or U3523 (N_3523,N_3232,N_3328);
nand U3524 (N_3524,N_3337,N_3381);
and U3525 (N_3525,N_3354,N_3244);
and U3526 (N_3526,N_3373,N_3250);
xnor U3527 (N_3527,N_3296,N_3251);
nand U3528 (N_3528,N_3375,N_3373);
nand U3529 (N_3529,N_3285,N_3382);
or U3530 (N_3530,N_3292,N_3334);
xor U3531 (N_3531,N_3348,N_3283);
nor U3532 (N_3532,N_3341,N_3201);
and U3533 (N_3533,N_3214,N_3269);
xor U3534 (N_3534,N_3289,N_3371);
nor U3535 (N_3535,N_3292,N_3211);
and U3536 (N_3536,N_3288,N_3298);
and U3537 (N_3537,N_3356,N_3265);
nand U3538 (N_3538,N_3294,N_3346);
nor U3539 (N_3539,N_3309,N_3281);
nand U3540 (N_3540,N_3213,N_3352);
nor U3541 (N_3541,N_3340,N_3316);
and U3542 (N_3542,N_3320,N_3317);
and U3543 (N_3543,N_3342,N_3217);
and U3544 (N_3544,N_3272,N_3341);
nand U3545 (N_3545,N_3315,N_3249);
nor U3546 (N_3546,N_3377,N_3200);
nor U3547 (N_3547,N_3313,N_3261);
nor U3548 (N_3548,N_3233,N_3390);
nand U3549 (N_3549,N_3341,N_3397);
nand U3550 (N_3550,N_3280,N_3350);
or U3551 (N_3551,N_3394,N_3348);
nand U3552 (N_3552,N_3360,N_3396);
xnor U3553 (N_3553,N_3290,N_3232);
nor U3554 (N_3554,N_3274,N_3339);
and U3555 (N_3555,N_3284,N_3201);
or U3556 (N_3556,N_3352,N_3329);
and U3557 (N_3557,N_3205,N_3291);
or U3558 (N_3558,N_3224,N_3296);
and U3559 (N_3559,N_3374,N_3333);
nor U3560 (N_3560,N_3348,N_3213);
and U3561 (N_3561,N_3299,N_3298);
nor U3562 (N_3562,N_3285,N_3354);
and U3563 (N_3563,N_3242,N_3306);
nor U3564 (N_3564,N_3307,N_3242);
xor U3565 (N_3565,N_3292,N_3260);
and U3566 (N_3566,N_3246,N_3221);
or U3567 (N_3567,N_3216,N_3236);
nor U3568 (N_3568,N_3330,N_3270);
nor U3569 (N_3569,N_3335,N_3238);
nand U3570 (N_3570,N_3245,N_3375);
nand U3571 (N_3571,N_3314,N_3300);
and U3572 (N_3572,N_3236,N_3310);
or U3573 (N_3573,N_3226,N_3359);
nor U3574 (N_3574,N_3358,N_3260);
xnor U3575 (N_3575,N_3241,N_3333);
nor U3576 (N_3576,N_3364,N_3287);
nand U3577 (N_3577,N_3387,N_3325);
nand U3578 (N_3578,N_3378,N_3396);
nor U3579 (N_3579,N_3367,N_3247);
nor U3580 (N_3580,N_3364,N_3316);
and U3581 (N_3581,N_3308,N_3267);
or U3582 (N_3582,N_3349,N_3216);
nor U3583 (N_3583,N_3260,N_3304);
xor U3584 (N_3584,N_3324,N_3226);
nand U3585 (N_3585,N_3208,N_3391);
or U3586 (N_3586,N_3266,N_3214);
nand U3587 (N_3587,N_3350,N_3340);
nor U3588 (N_3588,N_3230,N_3397);
nand U3589 (N_3589,N_3354,N_3393);
nand U3590 (N_3590,N_3273,N_3298);
and U3591 (N_3591,N_3362,N_3325);
nor U3592 (N_3592,N_3207,N_3292);
nor U3593 (N_3593,N_3305,N_3279);
or U3594 (N_3594,N_3325,N_3243);
nor U3595 (N_3595,N_3211,N_3233);
xnor U3596 (N_3596,N_3226,N_3369);
and U3597 (N_3597,N_3386,N_3230);
nand U3598 (N_3598,N_3221,N_3363);
or U3599 (N_3599,N_3304,N_3310);
nor U3600 (N_3600,N_3554,N_3579);
nor U3601 (N_3601,N_3590,N_3480);
and U3602 (N_3602,N_3414,N_3584);
nand U3603 (N_3603,N_3420,N_3530);
xor U3604 (N_3604,N_3410,N_3587);
and U3605 (N_3605,N_3582,N_3560);
or U3606 (N_3606,N_3565,N_3424);
nor U3607 (N_3607,N_3514,N_3572);
nand U3608 (N_3608,N_3461,N_3562);
nand U3609 (N_3609,N_3526,N_3401);
or U3610 (N_3610,N_3434,N_3546);
and U3611 (N_3611,N_3559,N_3433);
nand U3612 (N_3612,N_3594,N_3495);
nor U3613 (N_3613,N_3501,N_3597);
and U3614 (N_3614,N_3586,N_3561);
nand U3615 (N_3615,N_3525,N_3459);
or U3616 (N_3616,N_3419,N_3599);
nand U3617 (N_3617,N_3441,N_3496);
nand U3618 (N_3618,N_3542,N_3485);
nor U3619 (N_3619,N_3598,N_3555);
nor U3620 (N_3620,N_3581,N_3446);
nor U3621 (N_3621,N_3457,N_3529);
or U3622 (N_3622,N_3479,N_3570);
and U3623 (N_3623,N_3557,N_3415);
nand U3624 (N_3624,N_3472,N_3558);
and U3625 (N_3625,N_3563,N_3406);
nand U3626 (N_3626,N_3504,N_3492);
xnor U3627 (N_3627,N_3426,N_3445);
nor U3628 (N_3628,N_3402,N_3456);
and U3629 (N_3629,N_3438,N_3413);
or U3630 (N_3630,N_3467,N_3512);
xnor U3631 (N_3631,N_3442,N_3425);
nor U3632 (N_3632,N_3444,N_3437);
nand U3633 (N_3633,N_3462,N_3528);
and U3634 (N_3634,N_3482,N_3469);
nand U3635 (N_3635,N_3538,N_3517);
or U3636 (N_3636,N_3483,N_3523);
nor U3637 (N_3637,N_3518,N_3547);
nor U3638 (N_3638,N_3533,N_3576);
nand U3639 (N_3639,N_3490,N_3405);
nand U3640 (N_3640,N_3503,N_3577);
and U3641 (N_3641,N_3478,N_3436);
or U3642 (N_3642,N_3564,N_3421);
nand U3643 (N_3643,N_3578,N_3535);
nor U3644 (N_3644,N_3511,N_3509);
or U3645 (N_3645,N_3493,N_3592);
nand U3646 (N_3646,N_3507,N_3431);
and U3647 (N_3647,N_3429,N_3536);
nand U3648 (N_3648,N_3596,N_3404);
nor U3649 (N_3649,N_3516,N_3502);
or U3650 (N_3650,N_3498,N_3423);
xor U3651 (N_3651,N_3400,N_3450);
and U3652 (N_3652,N_3476,N_3521);
and U3653 (N_3653,N_3453,N_3585);
and U3654 (N_3654,N_3447,N_3513);
and U3655 (N_3655,N_3574,N_3463);
nand U3656 (N_3656,N_3455,N_3544);
nand U3657 (N_3657,N_3540,N_3543);
nor U3658 (N_3658,N_3422,N_3417);
nand U3659 (N_3659,N_3487,N_3531);
xor U3660 (N_3660,N_3448,N_3566);
nand U3661 (N_3661,N_3534,N_3553);
or U3662 (N_3662,N_3588,N_3494);
nand U3663 (N_3663,N_3575,N_3499);
or U3664 (N_3664,N_3466,N_3428);
nor U3665 (N_3665,N_3593,N_3484);
or U3666 (N_3666,N_3500,N_3520);
or U3667 (N_3667,N_3549,N_3451);
and U3668 (N_3668,N_3403,N_3412);
or U3669 (N_3669,N_3460,N_3551);
nand U3670 (N_3670,N_3454,N_3411);
nand U3671 (N_3671,N_3573,N_3488);
or U3672 (N_3672,N_3548,N_3443);
nand U3673 (N_3673,N_3505,N_3477);
and U3674 (N_3674,N_3464,N_3432);
or U3675 (N_3675,N_3527,N_3583);
and U3676 (N_3676,N_3458,N_3473);
nand U3677 (N_3677,N_3427,N_3452);
nor U3678 (N_3678,N_3440,N_3435);
nand U3679 (N_3679,N_3515,N_3510);
and U3680 (N_3680,N_3475,N_3465);
nand U3681 (N_3681,N_3522,N_3418);
nor U3682 (N_3682,N_3489,N_3580);
nand U3683 (N_3683,N_3541,N_3471);
nor U3684 (N_3684,N_3591,N_3552);
and U3685 (N_3685,N_3539,N_3439);
nand U3686 (N_3686,N_3567,N_3491);
or U3687 (N_3687,N_3470,N_3556);
and U3688 (N_3688,N_3497,N_3486);
and U3689 (N_3689,N_3537,N_3508);
nand U3690 (N_3690,N_3409,N_3568);
xnor U3691 (N_3691,N_3506,N_3468);
nor U3692 (N_3692,N_3407,N_3416);
or U3693 (N_3693,N_3474,N_3449);
nor U3694 (N_3694,N_3571,N_3481);
or U3695 (N_3695,N_3532,N_3545);
and U3696 (N_3696,N_3595,N_3408);
or U3697 (N_3697,N_3430,N_3569);
nor U3698 (N_3698,N_3524,N_3589);
and U3699 (N_3699,N_3550,N_3519);
xor U3700 (N_3700,N_3525,N_3428);
or U3701 (N_3701,N_3453,N_3526);
nor U3702 (N_3702,N_3522,N_3463);
and U3703 (N_3703,N_3470,N_3487);
nor U3704 (N_3704,N_3509,N_3599);
nand U3705 (N_3705,N_3518,N_3450);
nand U3706 (N_3706,N_3590,N_3441);
nor U3707 (N_3707,N_3508,N_3593);
nor U3708 (N_3708,N_3414,N_3432);
nand U3709 (N_3709,N_3438,N_3511);
nand U3710 (N_3710,N_3549,N_3547);
and U3711 (N_3711,N_3554,N_3557);
nand U3712 (N_3712,N_3533,N_3479);
xor U3713 (N_3713,N_3562,N_3582);
and U3714 (N_3714,N_3490,N_3448);
xor U3715 (N_3715,N_3408,N_3445);
xnor U3716 (N_3716,N_3505,N_3569);
nand U3717 (N_3717,N_3515,N_3470);
nor U3718 (N_3718,N_3591,N_3561);
nor U3719 (N_3719,N_3417,N_3478);
nor U3720 (N_3720,N_3405,N_3456);
or U3721 (N_3721,N_3503,N_3595);
and U3722 (N_3722,N_3445,N_3571);
and U3723 (N_3723,N_3566,N_3437);
and U3724 (N_3724,N_3458,N_3402);
nor U3725 (N_3725,N_3598,N_3442);
nor U3726 (N_3726,N_3536,N_3523);
and U3727 (N_3727,N_3552,N_3599);
and U3728 (N_3728,N_3426,N_3550);
and U3729 (N_3729,N_3446,N_3580);
nor U3730 (N_3730,N_3463,N_3585);
and U3731 (N_3731,N_3512,N_3585);
nand U3732 (N_3732,N_3527,N_3480);
and U3733 (N_3733,N_3463,N_3569);
nor U3734 (N_3734,N_3433,N_3409);
nor U3735 (N_3735,N_3548,N_3466);
and U3736 (N_3736,N_3406,N_3465);
or U3737 (N_3737,N_3453,N_3452);
or U3738 (N_3738,N_3594,N_3548);
nand U3739 (N_3739,N_3430,N_3447);
nor U3740 (N_3740,N_3487,N_3536);
nand U3741 (N_3741,N_3507,N_3484);
nor U3742 (N_3742,N_3425,N_3437);
nand U3743 (N_3743,N_3447,N_3521);
nor U3744 (N_3744,N_3459,N_3435);
nand U3745 (N_3745,N_3496,N_3499);
nor U3746 (N_3746,N_3478,N_3408);
xor U3747 (N_3747,N_3486,N_3517);
and U3748 (N_3748,N_3411,N_3466);
and U3749 (N_3749,N_3548,N_3549);
nand U3750 (N_3750,N_3578,N_3576);
nor U3751 (N_3751,N_3597,N_3591);
and U3752 (N_3752,N_3442,N_3405);
nor U3753 (N_3753,N_3500,N_3554);
xor U3754 (N_3754,N_3426,N_3587);
or U3755 (N_3755,N_3503,N_3420);
nand U3756 (N_3756,N_3560,N_3555);
nand U3757 (N_3757,N_3498,N_3449);
xor U3758 (N_3758,N_3513,N_3477);
and U3759 (N_3759,N_3441,N_3410);
or U3760 (N_3760,N_3501,N_3591);
nand U3761 (N_3761,N_3485,N_3406);
nand U3762 (N_3762,N_3590,N_3586);
and U3763 (N_3763,N_3438,N_3478);
nor U3764 (N_3764,N_3545,N_3539);
nand U3765 (N_3765,N_3471,N_3464);
nor U3766 (N_3766,N_3553,N_3595);
nand U3767 (N_3767,N_3501,N_3504);
or U3768 (N_3768,N_3425,N_3514);
and U3769 (N_3769,N_3581,N_3503);
or U3770 (N_3770,N_3447,N_3474);
nor U3771 (N_3771,N_3507,N_3551);
nor U3772 (N_3772,N_3566,N_3578);
and U3773 (N_3773,N_3470,N_3533);
or U3774 (N_3774,N_3404,N_3571);
xnor U3775 (N_3775,N_3567,N_3428);
or U3776 (N_3776,N_3553,N_3499);
nand U3777 (N_3777,N_3444,N_3592);
nor U3778 (N_3778,N_3478,N_3531);
nor U3779 (N_3779,N_3511,N_3595);
nor U3780 (N_3780,N_3451,N_3534);
nor U3781 (N_3781,N_3428,N_3584);
xnor U3782 (N_3782,N_3539,N_3474);
nor U3783 (N_3783,N_3589,N_3431);
nand U3784 (N_3784,N_3592,N_3401);
xor U3785 (N_3785,N_3539,N_3522);
nand U3786 (N_3786,N_3449,N_3554);
nand U3787 (N_3787,N_3534,N_3560);
nor U3788 (N_3788,N_3532,N_3446);
nor U3789 (N_3789,N_3488,N_3537);
and U3790 (N_3790,N_3508,N_3474);
nand U3791 (N_3791,N_3522,N_3519);
nor U3792 (N_3792,N_3539,N_3402);
nor U3793 (N_3793,N_3518,N_3478);
and U3794 (N_3794,N_3447,N_3494);
nor U3795 (N_3795,N_3436,N_3520);
nor U3796 (N_3796,N_3576,N_3415);
nand U3797 (N_3797,N_3596,N_3576);
or U3798 (N_3798,N_3456,N_3527);
or U3799 (N_3799,N_3469,N_3546);
nor U3800 (N_3800,N_3745,N_3617);
nand U3801 (N_3801,N_3639,N_3691);
nor U3802 (N_3802,N_3604,N_3660);
nand U3803 (N_3803,N_3742,N_3695);
or U3804 (N_3804,N_3665,N_3730);
nand U3805 (N_3805,N_3788,N_3683);
nand U3806 (N_3806,N_3768,N_3608);
or U3807 (N_3807,N_3749,N_3711);
nand U3808 (N_3808,N_3731,N_3654);
nand U3809 (N_3809,N_3771,N_3629);
and U3810 (N_3810,N_3766,N_3670);
or U3811 (N_3811,N_3655,N_3661);
or U3812 (N_3812,N_3753,N_3770);
nor U3813 (N_3813,N_3638,N_3767);
xnor U3814 (N_3814,N_3758,N_3713);
and U3815 (N_3815,N_3652,N_3689);
nand U3816 (N_3816,N_3605,N_3757);
or U3817 (N_3817,N_3773,N_3725);
xor U3818 (N_3818,N_3791,N_3727);
or U3819 (N_3819,N_3677,N_3603);
nand U3820 (N_3820,N_3672,N_3615);
xor U3821 (N_3821,N_3649,N_3724);
nand U3822 (N_3822,N_3710,N_3795);
nor U3823 (N_3823,N_3612,N_3620);
nand U3824 (N_3824,N_3732,N_3675);
nand U3825 (N_3825,N_3776,N_3772);
and U3826 (N_3826,N_3721,N_3624);
and U3827 (N_3827,N_3626,N_3746);
xnor U3828 (N_3828,N_3799,N_3720);
nand U3829 (N_3829,N_3611,N_3671);
and U3830 (N_3830,N_3761,N_3700);
nor U3831 (N_3831,N_3636,N_3783);
nor U3832 (N_3832,N_3685,N_3687);
nor U3833 (N_3833,N_3778,N_3796);
or U3834 (N_3834,N_3667,N_3614);
nor U3835 (N_3835,N_3659,N_3719);
nand U3836 (N_3836,N_3769,N_3797);
nand U3837 (N_3837,N_3607,N_3748);
nand U3838 (N_3838,N_3676,N_3698);
nor U3839 (N_3839,N_3738,N_3723);
nor U3840 (N_3840,N_3760,N_3613);
nand U3841 (N_3841,N_3690,N_3646);
nor U3842 (N_3842,N_3790,N_3643);
or U3843 (N_3843,N_3680,N_3669);
xor U3844 (N_3844,N_3688,N_3755);
nand U3845 (N_3845,N_3627,N_3681);
nand U3846 (N_3846,N_3759,N_3609);
and U3847 (N_3847,N_3704,N_3702);
nand U3848 (N_3848,N_3621,N_3775);
nor U3849 (N_3849,N_3641,N_3674);
nand U3850 (N_3850,N_3717,N_3645);
or U3851 (N_3851,N_3792,N_3625);
and U3852 (N_3852,N_3618,N_3735);
and U3853 (N_3853,N_3662,N_3777);
nor U3854 (N_3854,N_3623,N_3763);
and U3855 (N_3855,N_3750,N_3779);
nand U3856 (N_3856,N_3786,N_3644);
and U3857 (N_3857,N_3606,N_3684);
and U3858 (N_3858,N_3679,N_3789);
or U3859 (N_3859,N_3648,N_3734);
nor U3860 (N_3860,N_3630,N_3635);
and U3861 (N_3861,N_3707,N_3600);
xor U3862 (N_3862,N_3632,N_3705);
and U3863 (N_3863,N_3754,N_3640);
or U3864 (N_3864,N_3764,N_3647);
xor U3865 (N_3865,N_3726,N_3631);
xnor U3866 (N_3866,N_3708,N_3642);
nand U3867 (N_3867,N_3653,N_3729);
and U3868 (N_3868,N_3781,N_3762);
and U3869 (N_3869,N_3628,N_3650);
and U3870 (N_3870,N_3601,N_3712);
nand U3871 (N_3871,N_3798,N_3780);
nor U3872 (N_3872,N_3739,N_3634);
nor U3873 (N_3873,N_3694,N_3787);
nand U3874 (N_3874,N_3663,N_3633);
nor U3875 (N_3875,N_3740,N_3701);
xnor U3876 (N_3876,N_3733,N_3741);
xnor U3877 (N_3877,N_3774,N_3651);
xor U3878 (N_3878,N_3658,N_3682);
and U3879 (N_3879,N_3744,N_3784);
or U3880 (N_3880,N_3637,N_3616);
nand U3881 (N_3881,N_3765,N_3782);
nand U3882 (N_3882,N_3697,N_3673);
or U3883 (N_3883,N_3686,N_3714);
nand U3884 (N_3884,N_3664,N_3756);
and U3885 (N_3885,N_3722,N_3657);
nand U3886 (N_3886,N_3678,N_3709);
and U3887 (N_3887,N_3668,N_3794);
nand U3888 (N_3888,N_3619,N_3602);
nand U3889 (N_3889,N_3706,N_3718);
or U3890 (N_3890,N_3743,N_3656);
nand U3891 (N_3891,N_3736,N_3699);
and U3892 (N_3892,N_3785,N_3728);
and U3893 (N_3893,N_3793,N_3696);
nand U3894 (N_3894,N_3622,N_3692);
nand U3895 (N_3895,N_3666,N_3693);
or U3896 (N_3896,N_3715,N_3610);
and U3897 (N_3897,N_3752,N_3751);
or U3898 (N_3898,N_3716,N_3737);
or U3899 (N_3899,N_3747,N_3703);
xor U3900 (N_3900,N_3705,N_3624);
nor U3901 (N_3901,N_3776,N_3736);
or U3902 (N_3902,N_3627,N_3746);
nand U3903 (N_3903,N_3700,N_3690);
or U3904 (N_3904,N_3755,N_3725);
and U3905 (N_3905,N_3704,N_3691);
nand U3906 (N_3906,N_3699,N_3658);
xor U3907 (N_3907,N_3734,N_3747);
and U3908 (N_3908,N_3707,N_3761);
or U3909 (N_3909,N_3619,N_3710);
nor U3910 (N_3910,N_3731,N_3715);
nand U3911 (N_3911,N_3612,N_3721);
nor U3912 (N_3912,N_3732,N_3651);
or U3913 (N_3913,N_3684,N_3615);
xnor U3914 (N_3914,N_3766,N_3691);
and U3915 (N_3915,N_3753,N_3798);
and U3916 (N_3916,N_3646,N_3718);
nand U3917 (N_3917,N_3688,N_3655);
nand U3918 (N_3918,N_3607,N_3605);
nand U3919 (N_3919,N_3783,N_3751);
nand U3920 (N_3920,N_3765,N_3635);
nor U3921 (N_3921,N_3763,N_3673);
nor U3922 (N_3922,N_3660,N_3737);
xnor U3923 (N_3923,N_3786,N_3655);
and U3924 (N_3924,N_3697,N_3675);
nor U3925 (N_3925,N_3785,N_3745);
nand U3926 (N_3926,N_3774,N_3617);
and U3927 (N_3927,N_3744,N_3650);
nand U3928 (N_3928,N_3749,N_3734);
xnor U3929 (N_3929,N_3668,N_3799);
xor U3930 (N_3930,N_3621,N_3681);
nor U3931 (N_3931,N_3613,N_3734);
xor U3932 (N_3932,N_3654,N_3701);
xor U3933 (N_3933,N_3734,N_3657);
nor U3934 (N_3934,N_3674,N_3784);
nand U3935 (N_3935,N_3659,N_3772);
nand U3936 (N_3936,N_3680,N_3790);
and U3937 (N_3937,N_3691,N_3742);
nor U3938 (N_3938,N_3768,N_3793);
nand U3939 (N_3939,N_3711,N_3790);
nor U3940 (N_3940,N_3657,N_3698);
and U3941 (N_3941,N_3621,N_3728);
nor U3942 (N_3942,N_3728,N_3643);
xor U3943 (N_3943,N_3680,N_3633);
nor U3944 (N_3944,N_3683,N_3717);
and U3945 (N_3945,N_3624,N_3688);
nand U3946 (N_3946,N_3634,N_3638);
nand U3947 (N_3947,N_3727,N_3783);
nand U3948 (N_3948,N_3732,N_3658);
xor U3949 (N_3949,N_3750,N_3739);
xor U3950 (N_3950,N_3679,N_3619);
or U3951 (N_3951,N_3619,N_3672);
nand U3952 (N_3952,N_3703,N_3625);
or U3953 (N_3953,N_3688,N_3728);
and U3954 (N_3954,N_3685,N_3700);
or U3955 (N_3955,N_3773,N_3778);
nand U3956 (N_3956,N_3691,N_3602);
xnor U3957 (N_3957,N_3723,N_3687);
xor U3958 (N_3958,N_3735,N_3722);
nor U3959 (N_3959,N_3689,N_3694);
or U3960 (N_3960,N_3744,N_3657);
nand U3961 (N_3961,N_3757,N_3619);
or U3962 (N_3962,N_3661,N_3703);
or U3963 (N_3963,N_3698,N_3684);
or U3964 (N_3964,N_3617,N_3621);
and U3965 (N_3965,N_3693,N_3650);
nor U3966 (N_3966,N_3627,N_3792);
nor U3967 (N_3967,N_3604,N_3691);
nand U3968 (N_3968,N_3656,N_3630);
nor U3969 (N_3969,N_3695,N_3606);
and U3970 (N_3970,N_3697,N_3743);
nand U3971 (N_3971,N_3657,N_3633);
nor U3972 (N_3972,N_3730,N_3633);
and U3973 (N_3973,N_3624,N_3744);
or U3974 (N_3974,N_3616,N_3778);
nand U3975 (N_3975,N_3779,N_3645);
xor U3976 (N_3976,N_3622,N_3726);
nor U3977 (N_3977,N_3748,N_3634);
nor U3978 (N_3978,N_3765,N_3612);
or U3979 (N_3979,N_3760,N_3631);
or U3980 (N_3980,N_3796,N_3661);
and U3981 (N_3981,N_3754,N_3694);
nand U3982 (N_3982,N_3695,N_3678);
xor U3983 (N_3983,N_3609,N_3792);
nand U3984 (N_3984,N_3781,N_3777);
nand U3985 (N_3985,N_3624,N_3727);
or U3986 (N_3986,N_3737,N_3691);
xor U3987 (N_3987,N_3668,N_3763);
xor U3988 (N_3988,N_3626,N_3655);
nand U3989 (N_3989,N_3689,N_3744);
or U3990 (N_3990,N_3613,N_3717);
nand U3991 (N_3991,N_3739,N_3655);
or U3992 (N_3992,N_3718,N_3645);
nand U3993 (N_3993,N_3672,N_3727);
nor U3994 (N_3994,N_3798,N_3680);
and U3995 (N_3995,N_3677,N_3762);
nor U3996 (N_3996,N_3668,N_3637);
and U3997 (N_3997,N_3746,N_3679);
nand U3998 (N_3998,N_3795,N_3693);
nor U3999 (N_3999,N_3612,N_3628);
nor U4000 (N_4000,N_3864,N_3866);
nor U4001 (N_4001,N_3846,N_3901);
and U4002 (N_4002,N_3944,N_3986);
or U4003 (N_4003,N_3899,N_3805);
nor U4004 (N_4004,N_3840,N_3961);
nand U4005 (N_4005,N_3824,N_3835);
and U4006 (N_4006,N_3843,N_3922);
nor U4007 (N_4007,N_3868,N_3971);
nor U4008 (N_4008,N_3998,N_3975);
xor U4009 (N_4009,N_3985,N_3948);
nand U4010 (N_4010,N_3919,N_3915);
and U4011 (N_4011,N_3976,N_3813);
or U4012 (N_4012,N_3987,N_3859);
xnor U4013 (N_4013,N_3946,N_3887);
xnor U4014 (N_4014,N_3810,N_3993);
nand U4015 (N_4015,N_3941,N_3822);
nor U4016 (N_4016,N_3829,N_3917);
nand U4017 (N_4017,N_3875,N_3804);
or U4018 (N_4018,N_3978,N_3955);
and U4019 (N_4019,N_3966,N_3897);
nor U4020 (N_4020,N_3881,N_3930);
nand U4021 (N_4021,N_3937,N_3850);
nor U4022 (N_4022,N_3823,N_3800);
and U4023 (N_4023,N_3984,N_3883);
nand U4024 (N_4024,N_3928,N_3817);
nor U4025 (N_4025,N_3953,N_3861);
or U4026 (N_4026,N_3841,N_3909);
xor U4027 (N_4027,N_3995,N_3990);
nand U4028 (N_4028,N_3906,N_3918);
nand U4029 (N_4029,N_3877,N_3807);
or U4030 (N_4030,N_3982,N_3972);
nand U4031 (N_4031,N_3924,N_3886);
and U4032 (N_4032,N_3852,N_3867);
and U4033 (N_4033,N_3942,N_3965);
nor U4034 (N_4034,N_3913,N_3838);
or U4035 (N_4035,N_3876,N_3851);
nor U4036 (N_4036,N_3960,N_3907);
and U4037 (N_4037,N_3834,N_3825);
and U4038 (N_4038,N_3855,N_3973);
and U4039 (N_4039,N_3951,N_3814);
and U4040 (N_4040,N_3974,N_3842);
nor U4041 (N_4041,N_3963,N_3812);
or U4042 (N_4042,N_3905,N_3977);
or U4043 (N_4043,N_3981,N_3957);
or U4044 (N_4044,N_3815,N_3903);
nand U4045 (N_4045,N_3819,N_3933);
xnor U4046 (N_4046,N_3929,N_3871);
and U4047 (N_4047,N_3895,N_3854);
nor U4048 (N_4048,N_3893,N_3904);
nand U4049 (N_4049,N_3908,N_3945);
nor U4050 (N_4050,N_3828,N_3935);
or U4051 (N_4051,N_3964,N_3940);
nand U4052 (N_4052,N_3931,N_3890);
nand U4053 (N_4053,N_3969,N_3880);
or U4054 (N_4054,N_3921,N_3956);
or U4055 (N_4055,N_3916,N_3832);
nor U4056 (N_4056,N_3896,N_3911);
and U4057 (N_4057,N_3970,N_3863);
or U4058 (N_4058,N_3839,N_3954);
or U4059 (N_4059,N_3902,N_3836);
and U4060 (N_4060,N_3934,N_3988);
or U4061 (N_4061,N_3959,N_3844);
and U4062 (N_4062,N_3991,N_3802);
or U4063 (N_4063,N_3927,N_3818);
nor U4064 (N_4064,N_3882,N_3808);
nor U4065 (N_4065,N_3892,N_3958);
nor U4066 (N_4066,N_3936,N_3857);
and U4067 (N_4067,N_3858,N_3809);
and U4068 (N_4068,N_3827,N_3938);
and U4069 (N_4069,N_3926,N_3900);
nor U4070 (N_4070,N_3849,N_3816);
or U4071 (N_4071,N_3820,N_3811);
and U4072 (N_4072,N_3845,N_3996);
and U4073 (N_4073,N_3950,N_3894);
and U4074 (N_4074,N_3856,N_3989);
nand U4075 (N_4075,N_3848,N_3878);
nor U4076 (N_4076,N_3806,N_3862);
or U4077 (N_4077,N_3884,N_3967);
nand U4078 (N_4078,N_3872,N_3943);
nand U4079 (N_4079,N_3865,N_3821);
and U4080 (N_4080,N_3939,N_3874);
and U4081 (N_4081,N_3831,N_3949);
nor U4082 (N_4082,N_3952,N_3962);
nand U4083 (N_4083,N_3920,N_3830);
nor U4084 (N_4084,N_3947,N_3891);
nor U4085 (N_4085,N_3914,N_3833);
nand U4086 (N_4086,N_3888,N_3826);
or U4087 (N_4087,N_3992,N_3912);
nand U4088 (N_4088,N_3847,N_3994);
nand U4089 (N_4089,N_3837,N_3932);
and U4090 (N_4090,N_3803,N_3889);
nor U4091 (N_4091,N_3910,N_3968);
nor U4092 (N_4092,N_3999,N_3879);
nand U4093 (N_4093,N_3898,N_3997);
and U4094 (N_4094,N_3923,N_3801);
nand U4095 (N_4095,N_3869,N_3870);
and U4096 (N_4096,N_3979,N_3980);
nor U4097 (N_4097,N_3885,N_3983);
nand U4098 (N_4098,N_3925,N_3853);
and U4099 (N_4099,N_3860,N_3873);
and U4100 (N_4100,N_3887,N_3925);
nor U4101 (N_4101,N_3971,N_3859);
or U4102 (N_4102,N_3816,N_3860);
nand U4103 (N_4103,N_3899,N_3848);
xor U4104 (N_4104,N_3994,N_3846);
nor U4105 (N_4105,N_3953,N_3828);
and U4106 (N_4106,N_3832,N_3860);
or U4107 (N_4107,N_3955,N_3981);
or U4108 (N_4108,N_3869,N_3807);
xnor U4109 (N_4109,N_3808,N_3851);
or U4110 (N_4110,N_3831,N_3809);
nand U4111 (N_4111,N_3979,N_3896);
nor U4112 (N_4112,N_3886,N_3842);
nand U4113 (N_4113,N_3865,N_3970);
or U4114 (N_4114,N_3984,N_3828);
nand U4115 (N_4115,N_3803,N_3972);
or U4116 (N_4116,N_3907,N_3920);
and U4117 (N_4117,N_3870,N_3939);
or U4118 (N_4118,N_3885,N_3886);
nand U4119 (N_4119,N_3865,N_3824);
and U4120 (N_4120,N_3856,N_3980);
or U4121 (N_4121,N_3913,N_3850);
xor U4122 (N_4122,N_3934,N_3993);
xnor U4123 (N_4123,N_3870,N_3843);
and U4124 (N_4124,N_3801,N_3860);
nand U4125 (N_4125,N_3943,N_3996);
or U4126 (N_4126,N_3829,N_3919);
nand U4127 (N_4127,N_3879,N_3810);
or U4128 (N_4128,N_3863,N_3873);
or U4129 (N_4129,N_3986,N_3836);
nand U4130 (N_4130,N_3956,N_3887);
nor U4131 (N_4131,N_3894,N_3819);
nor U4132 (N_4132,N_3992,N_3961);
nor U4133 (N_4133,N_3939,N_3882);
nor U4134 (N_4134,N_3954,N_3846);
and U4135 (N_4135,N_3876,N_3866);
or U4136 (N_4136,N_3934,N_3873);
nand U4137 (N_4137,N_3896,N_3851);
nand U4138 (N_4138,N_3959,N_3927);
nor U4139 (N_4139,N_3989,N_3871);
xnor U4140 (N_4140,N_3920,N_3983);
nor U4141 (N_4141,N_3809,N_3890);
nand U4142 (N_4142,N_3965,N_3881);
and U4143 (N_4143,N_3944,N_3861);
and U4144 (N_4144,N_3981,N_3978);
or U4145 (N_4145,N_3849,N_3892);
and U4146 (N_4146,N_3905,N_3995);
or U4147 (N_4147,N_3825,N_3947);
nand U4148 (N_4148,N_3856,N_3900);
xor U4149 (N_4149,N_3841,N_3939);
xnor U4150 (N_4150,N_3971,N_3883);
nand U4151 (N_4151,N_3974,N_3824);
and U4152 (N_4152,N_3916,N_3834);
nor U4153 (N_4153,N_3862,N_3990);
xnor U4154 (N_4154,N_3851,N_3929);
xnor U4155 (N_4155,N_3821,N_3838);
nand U4156 (N_4156,N_3853,N_3862);
nand U4157 (N_4157,N_3804,N_3824);
xor U4158 (N_4158,N_3824,N_3851);
or U4159 (N_4159,N_3899,N_3907);
or U4160 (N_4160,N_3817,N_3978);
nor U4161 (N_4161,N_3996,N_3941);
and U4162 (N_4162,N_3825,N_3954);
nand U4163 (N_4163,N_3891,N_3966);
or U4164 (N_4164,N_3967,N_3818);
or U4165 (N_4165,N_3905,N_3878);
or U4166 (N_4166,N_3951,N_3866);
or U4167 (N_4167,N_3918,N_3900);
nand U4168 (N_4168,N_3941,N_3995);
and U4169 (N_4169,N_3806,N_3822);
or U4170 (N_4170,N_3905,N_3836);
or U4171 (N_4171,N_3803,N_3990);
or U4172 (N_4172,N_3941,N_3899);
nor U4173 (N_4173,N_3865,N_3952);
or U4174 (N_4174,N_3817,N_3815);
or U4175 (N_4175,N_3861,N_3827);
nor U4176 (N_4176,N_3949,N_3905);
nand U4177 (N_4177,N_3986,N_3839);
nor U4178 (N_4178,N_3872,N_3800);
nor U4179 (N_4179,N_3974,N_3878);
nor U4180 (N_4180,N_3978,N_3961);
and U4181 (N_4181,N_3950,N_3931);
or U4182 (N_4182,N_3984,N_3946);
nor U4183 (N_4183,N_3849,N_3912);
or U4184 (N_4184,N_3891,N_3930);
and U4185 (N_4185,N_3975,N_3968);
nor U4186 (N_4186,N_3959,N_3810);
nor U4187 (N_4187,N_3847,N_3928);
or U4188 (N_4188,N_3805,N_3908);
and U4189 (N_4189,N_3938,N_3949);
xor U4190 (N_4190,N_3919,N_3846);
or U4191 (N_4191,N_3806,N_3813);
nor U4192 (N_4192,N_3935,N_3923);
and U4193 (N_4193,N_3864,N_3935);
and U4194 (N_4194,N_3819,N_3813);
nand U4195 (N_4195,N_3901,N_3837);
nand U4196 (N_4196,N_3949,N_3823);
or U4197 (N_4197,N_3874,N_3851);
and U4198 (N_4198,N_3836,N_3911);
xor U4199 (N_4199,N_3898,N_3833);
nor U4200 (N_4200,N_4181,N_4115);
nor U4201 (N_4201,N_4113,N_4071);
nand U4202 (N_4202,N_4096,N_4079);
or U4203 (N_4203,N_4029,N_4019);
nor U4204 (N_4204,N_4117,N_4042);
and U4205 (N_4205,N_4076,N_4165);
nand U4206 (N_4206,N_4020,N_4043);
nand U4207 (N_4207,N_4155,N_4039);
and U4208 (N_4208,N_4097,N_4158);
nor U4209 (N_4209,N_4195,N_4114);
nor U4210 (N_4210,N_4083,N_4037);
nor U4211 (N_4211,N_4028,N_4048);
nand U4212 (N_4212,N_4065,N_4151);
or U4213 (N_4213,N_4006,N_4170);
and U4214 (N_4214,N_4002,N_4157);
nand U4215 (N_4215,N_4093,N_4167);
or U4216 (N_4216,N_4090,N_4102);
nand U4217 (N_4217,N_4063,N_4031);
nand U4218 (N_4218,N_4112,N_4073);
nand U4219 (N_4219,N_4080,N_4138);
or U4220 (N_4220,N_4052,N_4058);
or U4221 (N_4221,N_4088,N_4130);
or U4222 (N_4222,N_4035,N_4030);
and U4223 (N_4223,N_4060,N_4056);
nand U4224 (N_4224,N_4160,N_4141);
xnor U4225 (N_4225,N_4055,N_4085);
nand U4226 (N_4226,N_4143,N_4180);
nand U4227 (N_4227,N_4182,N_4144);
nand U4228 (N_4228,N_4199,N_4150);
nand U4229 (N_4229,N_4021,N_4140);
nor U4230 (N_4230,N_4024,N_4045);
xor U4231 (N_4231,N_4166,N_4127);
nor U4232 (N_4232,N_4163,N_4059);
or U4233 (N_4233,N_4014,N_4010);
nand U4234 (N_4234,N_4069,N_4193);
or U4235 (N_4235,N_4168,N_4187);
or U4236 (N_4236,N_4162,N_4016);
nand U4237 (N_4237,N_4176,N_4095);
nand U4238 (N_4238,N_4082,N_4089);
or U4239 (N_4239,N_4017,N_4110);
nand U4240 (N_4240,N_4098,N_4190);
or U4241 (N_4241,N_4171,N_4178);
nand U4242 (N_4242,N_4186,N_4054);
xor U4243 (N_4243,N_4129,N_4120);
or U4244 (N_4244,N_4108,N_4156);
and U4245 (N_4245,N_4128,N_4111);
and U4246 (N_4246,N_4116,N_4012);
xnor U4247 (N_4247,N_4184,N_4027);
and U4248 (N_4248,N_4086,N_4041);
and U4249 (N_4249,N_4145,N_4146);
nand U4250 (N_4250,N_4173,N_4137);
or U4251 (N_4251,N_4040,N_4047);
nor U4252 (N_4252,N_4172,N_4044);
nand U4253 (N_4253,N_4196,N_4066);
nand U4254 (N_4254,N_4050,N_4148);
and U4255 (N_4255,N_4067,N_4009);
or U4256 (N_4256,N_4072,N_4007);
and U4257 (N_4257,N_4139,N_4084);
or U4258 (N_4258,N_4057,N_4136);
and U4259 (N_4259,N_4197,N_4174);
nand U4260 (N_4260,N_4034,N_4008);
xor U4261 (N_4261,N_4077,N_4126);
nor U4262 (N_4262,N_4049,N_4123);
nor U4263 (N_4263,N_4018,N_4154);
nand U4264 (N_4264,N_4061,N_4004);
nand U4265 (N_4265,N_4038,N_4122);
or U4266 (N_4266,N_4153,N_4124);
nor U4267 (N_4267,N_4001,N_4119);
or U4268 (N_4268,N_4164,N_4100);
and U4269 (N_4269,N_4051,N_4075);
or U4270 (N_4270,N_4081,N_4022);
and U4271 (N_4271,N_4125,N_4070);
xor U4272 (N_4272,N_4023,N_4152);
or U4273 (N_4273,N_4147,N_4099);
or U4274 (N_4274,N_4161,N_4087);
or U4275 (N_4275,N_4142,N_4194);
xor U4276 (N_4276,N_4198,N_4074);
nand U4277 (N_4277,N_4068,N_4000);
or U4278 (N_4278,N_4191,N_4091);
and U4279 (N_4279,N_4107,N_4106);
nand U4280 (N_4280,N_4131,N_4025);
xnor U4281 (N_4281,N_4132,N_4159);
and U4282 (N_4282,N_4177,N_4133);
nor U4283 (N_4283,N_4105,N_4005);
nor U4284 (N_4284,N_4053,N_4185);
xnor U4285 (N_4285,N_4013,N_4026);
or U4286 (N_4286,N_4192,N_4011);
nand U4287 (N_4287,N_4078,N_4092);
nand U4288 (N_4288,N_4046,N_4175);
xor U4289 (N_4289,N_4179,N_4094);
nor U4290 (N_4290,N_4134,N_4188);
and U4291 (N_4291,N_4003,N_4118);
nand U4292 (N_4292,N_4033,N_4103);
and U4293 (N_4293,N_4189,N_4101);
xnor U4294 (N_4294,N_4183,N_4169);
or U4295 (N_4295,N_4015,N_4064);
or U4296 (N_4296,N_4109,N_4121);
nand U4297 (N_4297,N_4032,N_4062);
xnor U4298 (N_4298,N_4104,N_4036);
and U4299 (N_4299,N_4149,N_4135);
or U4300 (N_4300,N_4094,N_4041);
nand U4301 (N_4301,N_4179,N_4126);
nand U4302 (N_4302,N_4160,N_4184);
nand U4303 (N_4303,N_4154,N_4093);
and U4304 (N_4304,N_4134,N_4186);
xor U4305 (N_4305,N_4010,N_4021);
or U4306 (N_4306,N_4130,N_4039);
xnor U4307 (N_4307,N_4095,N_4060);
nor U4308 (N_4308,N_4166,N_4053);
nand U4309 (N_4309,N_4092,N_4015);
and U4310 (N_4310,N_4127,N_4019);
nand U4311 (N_4311,N_4141,N_4083);
or U4312 (N_4312,N_4030,N_4070);
and U4313 (N_4313,N_4066,N_4043);
or U4314 (N_4314,N_4013,N_4151);
nor U4315 (N_4315,N_4119,N_4034);
nand U4316 (N_4316,N_4048,N_4040);
nor U4317 (N_4317,N_4144,N_4107);
nand U4318 (N_4318,N_4038,N_4011);
and U4319 (N_4319,N_4024,N_4199);
nor U4320 (N_4320,N_4076,N_4010);
nor U4321 (N_4321,N_4157,N_4052);
and U4322 (N_4322,N_4086,N_4169);
and U4323 (N_4323,N_4058,N_4075);
nor U4324 (N_4324,N_4161,N_4198);
nand U4325 (N_4325,N_4063,N_4056);
nor U4326 (N_4326,N_4104,N_4170);
nand U4327 (N_4327,N_4155,N_4061);
nor U4328 (N_4328,N_4086,N_4146);
nand U4329 (N_4329,N_4166,N_4027);
or U4330 (N_4330,N_4081,N_4177);
nand U4331 (N_4331,N_4122,N_4148);
and U4332 (N_4332,N_4034,N_4029);
nand U4333 (N_4333,N_4131,N_4129);
nand U4334 (N_4334,N_4047,N_4116);
nand U4335 (N_4335,N_4008,N_4167);
nor U4336 (N_4336,N_4169,N_4120);
nand U4337 (N_4337,N_4198,N_4036);
and U4338 (N_4338,N_4145,N_4124);
nor U4339 (N_4339,N_4132,N_4100);
and U4340 (N_4340,N_4100,N_4061);
nand U4341 (N_4341,N_4185,N_4138);
nand U4342 (N_4342,N_4029,N_4014);
nand U4343 (N_4343,N_4071,N_4029);
and U4344 (N_4344,N_4069,N_4165);
nor U4345 (N_4345,N_4187,N_4038);
nor U4346 (N_4346,N_4189,N_4043);
nor U4347 (N_4347,N_4189,N_4118);
and U4348 (N_4348,N_4146,N_4188);
nor U4349 (N_4349,N_4191,N_4086);
or U4350 (N_4350,N_4158,N_4091);
nand U4351 (N_4351,N_4186,N_4083);
and U4352 (N_4352,N_4052,N_4134);
or U4353 (N_4353,N_4133,N_4141);
nand U4354 (N_4354,N_4182,N_4132);
and U4355 (N_4355,N_4076,N_4086);
nand U4356 (N_4356,N_4086,N_4125);
nand U4357 (N_4357,N_4115,N_4148);
nand U4358 (N_4358,N_4179,N_4061);
and U4359 (N_4359,N_4099,N_4151);
nor U4360 (N_4360,N_4094,N_4108);
and U4361 (N_4361,N_4019,N_4005);
xnor U4362 (N_4362,N_4160,N_4047);
nor U4363 (N_4363,N_4147,N_4060);
or U4364 (N_4364,N_4135,N_4068);
or U4365 (N_4365,N_4052,N_4060);
nand U4366 (N_4366,N_4169,N_4121);
nor U4367 (N_4367,N_4144,N_4138);
nor U4368 (N_4368,N_4045,N_4064);
nor U4369 (N_4369,N_4073,N_4194);
nand U4370 (N_4370,N_4179,N_4035);
and U4371 (N_4371,N_4029,N_4058);
or U4372 (N_4372,N_4186,N_4123);
xor U4373 (N_4373,N_4175,N_4094);
nand U4374 (N_4374,N_4065,N_4093);
and U4375 (N_4375,N_4001,N_4163);
nor U4376 (N_4376,N_4091,N_4143);
nor U4377 (N_4377,N_4130,N_4192);
or U4378 (N_4378,N_4178,N_4176);
nand U4379 (N_4379,N_4119,N_4029);
nor U4380 (N_4380,N_4037,N_4092);
nor U4381 (N_4381,N_4061,N_4121);
and U4382 (N_4382,N_4133,N_4118);
or U4383 (N_4383,N_4153,N_4134);
and U4384 (N_4384,N_4135,N_4161);
and U4385 (N_4385,N_4055,N_4010);
or U4386 (N_4386,N_4013,N_4049);
and U4387 (N_4387,N_4093,N_4111);
nand U4388 (N_4388,N_4106,N_4025);
nor U4389 (N_4389,N_4196,N_4168);
nor U4390 (N_4390,N_4123,N_4162);
or U4391 (N_4391,N_4020,N_4013);
or U4392 (N_4392,N_4076,N_4108);
or U4393 (N_4393,N_4167,N_4140);
nor U4394 (N_4394,N_4115,N_4167);
nand U4395 (N_4395,N_4078,N_4050);
and U4396 (N_4396,N_4033,N_4006);
nor U4397 (N_4397,N_4126,N_4192);
and U4398 (N_4398,N_4121,N_4107);
nand U4399 (N_4399,N_4090,N_4113);
nor U4400 (N_4400,N_4330,N_4287);
or U4401 (N_4401,N_4202,N_4315);
and U4402 (N_4402,N_4301,N_4337);
or U4403 (N_4403,N_4246,N_4389);
xor U4404 (N_4404,N_4354,N_4295);
and U4405 (N_4405,N_4254,N_4227);
xor U4406 (N_4406,N_4364,N_4224);
and U4407 (N_4407,N_4359,N_4209);
and U4408 (N_4408,N_4268,N_4313);
and U4409 (N_4409,N_4264,N_4381);
and U4410 (N_4410,N_4323,N_4331);
nor U4411 (N_4411,N_4311,N_4373);
or U4412 (N_4412,N_4367,N_4297);
and U4413 (N_4413,N_4380,N_4365);
and U4414 (N_4414,N_4345,N_4258);
nand U4415 (N_4415,N_4274,N_4241);
and U4416 (N_4416,N_4387,N_4325);
nor U4417 (N_4417,N_4231,N_4397);
nand U4418 (N_4418,N_4296,N_4320);
and U4419 (N_4419,N_4277,N_4335);
nor U4420 (N_4420,N_4289,N_4235);
and U4421 (N_4421,N_4203,N_4360);
nor U4422 (N_4422,N_4234,N_4236);
nand U4423 (N_4423,N_4358,N_4378);
and U4424 (N_4424,N_4326,N_4303);
xnor U4425 (N_4425,N_4239,N_4271);
and U4426 (N_4426,N_4394,N_4267);
nor U4427 (N_4427,N_4272,N_4247);
or U4428 (N_4428,N_4379,N_4370);
nor U4429 (N_4429,N_4251,N_4217);
nor U4430 (N_4430,N_4392,N_4213);
or U4431 (N_4431,N_4314,N_4220);
or U4432 (N_4432,N_4218,N_4307);
and U4433 (N_4433,N_4372,N_4366);
or U4434 (N_4434,N_4346,N_4293);
and U4435 (N_4435,N_4350,N_4250);
or U4436 (N_4436,N_4255,N_4237);
and U4437 (N_4437,N_4362,N_4275);
nor U4438 (N_4438,N_4221,N_4273);
or U4439 (N_4439,N_4368,N_4200);
nand U4440 (N_4440,N_4279,N_4261);
or U4441 (N_4441,N_4386,N_4260);
nand U4442 (N_4442,N_4244,N_4294);
and U4443 (N_4443,N_4385,N_4399);
nor U4444 (N_4444,N_4396,N_4248);
nand U4445 (N_4445,N_4309,N_4369);
or U4446 (N_4446,N_4225,N_4351);
and U4447 (N_4447,N_4357,N_4349);
nor U4448 (N_4448,N_4222,N_4353);
and U4449 (N_4449,N_4310,N_4266);
or U4450 (N_4450,N_4333,N_4219);
nand U4451 (N_4451,N_4343,N_4252);
nand U4452 (N_4452,N_4259,N_4288);
or U4453 (N_4453,N_4253,N_4321);
and U4454 (N_4454,N_4329,N_4363);
and U4455 (N_4455,N_4201,N_4262);
or U4456 (N_4456,N_4327,N_4334);
nor U4457 (N_4457,N_4319,N_4398);
or U4458 (N_4458,N_4282,N_4214);
nor U4459 (N_4459,N_4230,N_4361);
and U4460 (N_4460,N_4382,N_4238);
or U4461 (N_4461,N_4376,N_4356);
nand U4462 (N_4462,N_4308,N_4245);
and U4463 (N_4463,N_4322,N_4375);
or U4464 (N_4464,N_4298,N_4280);
nand U4465 (N_4465,N_4284,N_4348);
or U4466 (N_4466,N_4223,N_4263);
nor U4467 (N_4467,N_4384,N_4383);
or U4468 (N_4468,N_4300,N_4332);
nor U4469 (N_4469,N_4229,N_4336);
nand U4470 (N_4470,N_4355,N_4216);
or U4471 (N_4471,N_4304,N_4233);
and U4472 (N_4472,N_4215,N_4205);
nor U4473 (N_4473,N_4318,N_4270);
nand U4474 (N_4474,N_4265,N_4306);
and U4475 (N_4475,N_4291,N_4212);
nand U4476 (N_4476,N_4257,N_4206);
nor U4477 (N_4477,N_4249,N_4240);
nand U4478 (N_4478,N_4276,N_4226);
or U4479 (N_4479,N_4338,N_4324);
nor U4480 (N_4480,N_4317,N_4395);
and U4481 (N_4481,N_4312,N_4228);
nand U4482 (N_4482,N_4347,N_4299);
nand U4483 (N_4483,N_4286,N_4344);
and U4484 (N_4484,N_4302,N_4208);
or U4485 (N_4485,N_4285,N_4281);
xnor U4486 (N_4486,N_4305,N_4341);
xor U4487 (N_4487,N_4374,N_4316);
nand U4488 (N_4488,N_4393,N_4242);
or U4489 (N_4489,N_4290,N_4352);
nand U4490 (N_4490,N_4328,N_4391);
xor U4491 (N_4491,N_4243,N_4339);
and U4492 (N_4492,N_4210,N_4211);
and U4493 (N_4493,N_4377,N_4292);
nand U4494 (N_4494,N_4371,N_4278);
nand U4495 (N_4495,N_4340,N_4342);
nor U4496 (N_4496,N_4388,N_4204);
or U4497 (N_4497,N_4283,N_4256);
nand U4498 (N_4498,N_4207,N_4232);
and U4499 (N_4499,N_4269,N_4390);
or U4500 (N_4500,N_4296,N_4267);
and U4501 (N_4501,N_4338,N_4326);
or U4502 (N_4502,N_4332,N_4365);
nand U4503 (N_4503,N_4385,N_4392);
or U4504 (N_4504,N_4338,N_4327);
nand U4505 (N_4505,N_4211,N_4257);
nor U4506 (N_4506,N_4250,N_4348);
nor U4507 (N_4507,N_4277,N_4240);
and U4508 (N_4508,N_4297,N_4360);
nor U4509 (N_4509,N_4304,N_4296);
nand U4510 (N_4510,N_4311,N_4218);
nand U4511 (N_4511,N_4230,N_4366);
nand U4512 (N_4512,N_4276,N_4382);
xor U4513 (N_4513,N_4337,N_4282);
nor U4514 (N_4514,N_4215,N_4352);
or U4515 (N_4515,N_4272,N_4353);
nor U4516 (N_4516,N_4218,N_4245);
nand U4517 (N_4517,N_4288,N_4203);
nor U4518 (N_4518,N_4387,N_4230);
and U4519 (N_4519,N_4328,N_4252);
xor U4520 (N_4520,N_4330,N_4364);
or U4521 (N_4521,N_4259,N_4252);
nor U4522 (N_4522,N_4313,N_4261);
nor U4523 (N_4523,N_4365,N_4335);
nand U4524 (N_4524,N_4275,N_4369);
nor U4525 (N_4525,N_4352,N_4229);
nor U4526 (N_4526,N_4284,N_4368);
xnor U4527 (N_4527,N_4227,N_4232);
nand U4528 (N_4528,N_4313,N_4286);
nor U4529 (N_4529,N_4395,N_4313);
nor U4530 (N_4530,N_4367,N_4229);
or U4531 (N_4531,N_4295,N_4276);
nor U4532 (N_4532,N_4334,N_4394);
or U4533 (N_4533,N_4203,N_4231);
or U4534 (N_4534,N_4259,N_4351);
or U4535 (N_4535,N_4379,N_4341);
and U4536 (N_4536,N_4289,N_4225);
nand U4537 (N_4537,N_4342,N_4200);
or U4538 (N_4538,N_4243,N_4226);
nor U4539 (N_4539,N_4236,N_4346);
nor U4540 (N_4540,N_4397,N_4364);
and U4541 (N_4541,N_4256,N_4398);
xor U4542 (N_4542,N_4383,N_4389);
or U4543 (N_4543,N_4223,N_4383);
or U4544 (N_4544,N_4263,N_4392);
nor U4545 (N_4545,N_4363,N_4276);
and U4546 (N_4546,N_4207,N_4399);
nor U4547 (N_4547,N_4360,N_4278);
nand U4548 (N_4548,N_4229,N_4368);
and U4549 (N_4549,N_4360,N_4213);
nand U4550 (N_4550,N_4306,N_4247);
nand U4551 (N_4551,N_4271,N_4231);
nor U4552 (N_4552,N_4284,N_4339);
nor U4553 (N_4553,N_4255,N_4214);
or U4554 (N_4554,N_4274,N_4329);
nand U4555 (N_4555,N_4243,N_4224);
xnor U4556 (N_4556,N_4361,N_4321);
and U4557 (N_4557,N_4394,N_4376);
nand U4558 (N_4558,N_4385,N_4212);
or U4559 (N_4559,N_4263,N_4284);
nor U4560 (N_4560,N_4328,N_4345);
or U4561 (N_4561,N_4218,N_4301);
xnor U4562 (N_4562,N_4249,N_4294);
nor U4563 (N_4563,N_4218,N_4347);
nand U4564 (N_4564,N_4361,N_4207);
nor U4565 (N_4565,N_4350,N_4223);
and U4566 (N_4566,N_4224,N_4381);
nor U4567 (N_4567,N_4201,N_4207);
or U4568 (N_4568,N_4279,N_4217);
nand U4569 (N_4569,N_4333,N_4361);
and U4570 (N_4570,N_4219,N_4352);
and U4571 (N_4571,N_4387,N_4296);
nor U4572 (N_4572,N_4396,N_4290);
or U4573 (N_4573,N_4270,N_4243);
xor U4574 (N_4574,N_4385,N_4243);
or U4575 (N_4575,N_4253,N_4280);
and U4576 (N_4576,N_4261,N_4332);
and U4577 (N_4577,N_4340,N_4306);
nor U4578 (N_4578,N_4223,N_4289);
and U4579 (N_4579,N_4233,N_4225);
and U4580 (N_4580,N_4289,N_4348);
nor U4581 (N_4581,N_4232,N_4313);
nand U4582 (N_4582,N_4392,N_4373);
nand U4583 (N_4583,N_4323,N_4259);
xor U4584 (N_4584,N_4273,N_4212);
nand U4585 (N_4585,N_4381,N_4331);
nor U4586 (N_4586,N_4222,N_4239);
and U4587 (N_4587,N_4345,N_4286);
and U4588 (N_4588,N_4210,N_4298);
nor U4589 (N_4589,N_4256,N_4233);
nand U4590 (N_4590,N_4393,N_4240);
or U4591 (N_4591,N_4316,N_4255);
or U4592 (N_4592,N_4394,N_4304);
nor U4593 (N_4593,N_4333,N_4307);
and U4594 (N_4594,N_4216,N_4214);
and U4595 (N_4595,N_4239,N_4337);
and U4596 (N_4596,N_4374,N_4266);
and U4597 (N_4597,N_4266,N_4361);
nand U4598 (N_4598,N_4376,N_4354);
or U4599 (N_4599,N_4230,N_4281);
nand U4600 (N_4600,N_4480,N_4420);
and U4601 (N_4601,N_4471,N_4440);
nand U4602 (N_4602,N_4421,N_4538);
nor U4603 (N_4603,N_4446,N_4563);
xor U4604 (N_4604,N_4579,N_4531);
nand U4605 (N_4605,N_4599,N_4404);
or U4606 (N_4606,N_4555,N_4546);
and U4607 (N_4607,N_4464,N_4477);
nor U4608 (N_4608,N_4499,N_4454);
or U4609 (N_4609,N_4574,N_4463);
nor U4610 (N_4610,N_4484,N_4447);
and U4611 (N_4611,N_4575,N_4510);
and U4612 (N_4612,N_4472,N_4549);
and U4613 (N_4613,N_4545,N_4565);
and U4614 (N_4614,N_4497,N_4543);
nor U4615 (N_4615,N_4473,N_4550);
or U4616 (N_4616,N_4490,N_4475);
nand U4617 (N_4617,N_4482,N_4413);
or U4618 (N_4618,N_4402,N_4569);
and U4619 (N_4619,N_4589,N_4529);
xor U4620 (N_4620,N_4594,N_4479);
nor U4621 (N_4621,N_4465,N_4562);
or U4622 (N_4622,N_4491,N_4564);
nand U4623 (N_4623,N_4485,N_4540);
nand U4624 (N_4624,N_4439,N_4415);
nand U4625 (N_4625,N_4584,N_4572);
nand U4626 (N_4626,N_4498,N_4432);
and U4627 (N_4627,N_4561,N_4532);
xor U4628 (N_4628,N_4578,N_4450);
nand U4629 (N_4629,N_4526,N_4528);
and U4630 (N_4630,N_4598,N_4583);
or U4631 (N_4631,N_4449,N_4592);
and U4632 (N_4632,N_4568,N_4448);
nor U4633 (N_4633,N_4542,N_4487);
or U4634 (N_4634,N_4533,N_4585);
or U4635 (N_4635,N_4500,N_4520);
and U4636 (N_4636,N_4516,N_4557);
nand U4637 (N_4637,N_4573,N_4438);
or U4638 (N_4638,N_4539,N_4582);
nor U4639 (N_4639,N_4504,N_4444);
and U4640 (N_4640,N_4428,N_4521);
nor U4641 (N_4641,N_4456,N_4547);
and U4642 (N_4642,N_4496,N_4481);
xnor U4643 (N_4643,N_4567,N_4527);
nor U4644 (N_4644,N_4408,N_4593);
nand U4645 (N_4645,N_4466,N_4452);
and U4646 (N_4646,N_4588,N_4576);
nand U4647 (N_4647,N_4541,N_4595);
nand U4648 (N_4648,N_4483,N_4581);
or U4649 (N_4649,N_4433,N_4519);
or U4650 (N_4650,N_4430,N_4434);
or U4651 (N_4651,N_4554,N_4458);
nand U4652 (N_4652,N_4431,N_4423);
nor U4653 (N_4653,N_4590,N_4492);
or U4654 (N_4654,N_4407,N_4426);
xor U4655 (N_4655,N_4486,N_4418);
and U4656 (N_4656,N_4414,N_4453);
nand U4657 (N_4657,N_4469,N_4451);
and U4658 (N_4658,N_4597,N_4468);
and U4659 (N_4659,N_4416,N_4551);
nor U4660 (N_4660,N_4559,N_4403);
nand U4661 (N_4661,N_4525,N_4400);
and U4662 (N_4662,N_4437,N_4474);
or U4663 (N_4663,N_4512,N_4457);
xor U4664 (N_4664,N_4422,N_4577);
and U4665 (N_4665,N_4523,N_4425);
nand U4666 (N_4666,N_4460,N_4560);
nand U4667 (N_4667,N_4455,N_4515);
nand U4668 (N_4668,N_4441,N_4461);
nand U4669 (N_4669,N_4427,N_4508);
nand U4670 (N_4670,N_4502,N_4534);
and U4671 (N_4671,N_4505,N_4405);
nand U4672 (N_4672,N_4459,N_4509);
nor U4673 (N_4673,N_4544,N_4406);
nor U4674 (N_4674,N_4411,N_4548);
and U4675 (N_4675,N_4443,N_4470);
xnor U4676 (N_4676,N_4511,N_4535);
or U4677 (N_4677,N_4596,N_4417);
or U4678 (N_4678,N_4591,N_4518);
and U4679 (N_4679,N_4552,N_4401);
nor U4680 (N_4680,N_4553,N_4410);
nand U4681 (N_4681,N_4493,N_4476);
and U4682 (N_4682,N_4556,N_4587);
or U4683 (N_4683,N_4489,N_4570);
nor U4684 (N_4684,N_4442,N_4409);
nor U4685 (N_4685,N_4501,N_4462);
or U4686 (N_4686,N_4580,N_4488);
or U4687 (N_4687,N_4524,N_4506);
and U4688 (N_4688,N_4566,N_4467);
and U4689 (N_4689,N_4445,N_4571);
nand U4690 (N_4690,N_4412,N_4558);
nor U4691 (N_4691,N_4435,N_4495);
and U4692 (N_4692,N_4436,N_4530);
xor U4693 (N_4693,N_4586,N_4537);
nand U4694 (N_4694,N_4494,N_4419);
or U4695 (N_4695,N_4522,N_4513);
or U4696 (N_4696,N_4429,N_4424);
or U4697 (N_4697,N_4507,N_4517);
nor U4698 (N_4698,N_4514,N_4503);
nor U4699 (N_4699,N_4536,N_4478);
nand U4700 (N_4700,N_4490,N_4566);
nor U4701 (N_4701,N_4558,N_4445);
and U4702 (N_4702,N_4458,N_4516);
or U4703 (N_4703,N_4472,N_4457);
nand U4704 (N_4704,N_4407,N_4503);
nand U4705 (N_4705,N_4493,N_4538);
and U4706 (N_4706,N_4587,N_4585);
nor U4707 (N_4707,N_4410,N_4527);
and U4708 (N_4708,N_4457,N_4578);
or U4709 (N_4709,N_4510,N_4443);
or U4710 (N_4710,N_4561,N_4470);
xnor U4711 (N_4711,N_4510,N_4481);
nor U4712 (N_4712,N_4513,N_4560);
nand U4713 (N_4713,N_4408,N_4403);
nand U4714 (N_4714,N_4438,N_4461);
nor U4715 (N_4715,N_4563,N_4576);
xnor U4716 (N_4716,N_4518,N_4477);
and U4717 (N_4717,N_4425,N_4544);
nor U4718 (N_4718,N_4545,N_4410);
and U4719 (N_4719,N_4517,N_4588);
nand U4720 (N_4720,N_4584,N_4432);
nor U4721 (N_4721,N_4427,N_4477);
nand U4722 (N_4722,N_4518,N_4539);
nor U4723 (N_4723,N_4445,N_4539);
nor U4724 (N_4724,N_4570,N_4487);
nor U4725 (N_4725,N_4578,N_4513);
or U4726 (N_4726,N_4481,N_4414);
nand U4727 (N_4727,N_4564,N_4511);
nor U4728 (N_4728,N_4498,N_4514);
or U4729 (N_4729,N_4541,N_4585);
and U4730 (N_4730,N_4589,N_4442);
or U4731 (N_4731,N_4464,N_4597);
nand U4732 (N_4732,N_4404,N_4479);
nand U4733 (N_4733,N_4583,N_4420);
xor U4734 (N_4734,N_4580,N_4418);
or U4735 (N_4735,N_4436,N_4596);
nor U4736 (N_4736,N_4496,N_4469);
nand U4737 (N_4737,N_4571,N_4538);
xor U4738 (N_4738,N_4566,N_4448);
nor U4739 (N_4739,N_4499,N_4462);
or U4740 (N_4740,N_4429,N_4446);
or U4741 (N_4741,N_4505,N_4498);
and U4742 (N_4742,N_4599,N_4508);
nand U4743 (N_4743,N_4421,N_4588);
nor U4744 (N_4744,N_4455,N_4568);
nand U4745 (N_4745,N_4462,N_4525);
and U4746 (N_4746,N_4411,N_4525);
and U4747 (N_4747,N_4555,N_4522);
nor U4748 (N_4748,N_4537,N_4595);
and U4749 (N_4749,N_4453,N_4450);
xnor U4750 (N_4750,N_4552,N_4447);
nor U4751 (N_4751,N_4554,N_4413);
or U4752 (N_4752,N_4429,N_4505);
or U4753 (N_4753,N_4588,N_4438);
or U4754 (N_4754,N_4465,N_4511);
nor U4755 (N_4755,N_4549,N_4540);
and U4756 (N_4756,N_4487,N_4552);
or U4757 (N_4757,N_4440,N_4461);
nor U4758 (N_4758,N_4489,N_4460);
and U4759 (N_4759,N_4471,N_4503);
and U4760 (N_4760,N_4569,N_4576);
and U4761 (N_4761,N_4480,N_4441);
and U4762 (N_4762,N_4593,N_4472);
nand U4763 (N_4763,N_4501,N_4504);
xor U4764 (N_4764,N_4498,N_4555);
nor U4765 (N_4765,N_4541,N_4418);
xnor U4766 (N_4766,N_4564,N_4527);
and U4767 (N_4767,N_4446,N_4407);
or U4768 (N_4768,N_4506,N_4458);
and U4769 (N_4769,N_4432,N_4442);
and U4770 (N_4770,N_4418,N_4563);
or U4771 (N_4771,N_4586,N_4426);
or U4772 (N_4772,N_4567,N_4495);
or U4773 (N_4773,N_4434,N_4422);
xnor U4774 (N_4774,N_4570,N_4507);
nand U4775 (N_4775,N_4539,N_4561);
nand U4776 (N_4776,N_4406,N_4480);
or U4777 (N_4777,N_4435,N_4468);
nor U4778 (N_4778,N_4524,N_4568);
or U4779 (N_4779,N_4430,N_4597);
nor U4780 (N_4780,N_4521,N_4540);
nor U4781 (N_4781,N_4404,N_4485);
and U4782 (N_4782,N_4457,N_4452);
nand U4783 (N_4783,N_4412,N_4548);
or U4784 (N_4784,N_4446,N_4508);
and U4785 (N_4785,N_4403,N_4547);
or U4786 (N_4786,N_4517,N_4584);
xnor U4787 (N_4787,N_4438,N_4437);
nor U4788 (N_4788,N_4413,N_4456);
and U4789 (N_4789,N_4587,N_4565);
or U4790 (N_4790,N_4459,N_4416);
nand U4791 (N_4791,N_4491,N_4551);
nand U4792 (N_4792,N_4560,N_4550);
or U4793 (N_4793,N_4531,N_4468);
and U4794 (N_4794,N_4491,N_4530);
nand U4795 (N_4795,N_4530,N_4588);
nor U4796 (N_4796,N_4447,N_4473);
or U4797 (N_4797,N_4503,N_4409);
or U4798 (N_4798,N_4409,N_4433);
and U4799 (N_4799,N_4447,N_4574);
nor U4800 (N_4800,N_4632,N_4777);
and U4801 (N_4801,N_4622,N_4648);
or U4802 (N_4802,N_4746,N_4658);
nor U4803 (N_4803,N_4751,N_4768);
and U4804 (N_4804,N_4742,N_4724);
or U4805 (N_4805,N_4625,N_4705);
and U4806 (N_4806,N_4698,N_4665);
nor U4807 (N_4807,N_4654,N_4602);
and U4808 (N_4808,N_4735,N_4781);
nor U4809 (N_4809,N_4772,N_4619);
nor U4810 (N_4810,N_4722,N_4604);
nand U4811 (N_4811,N_4655,N_4618);
nand U4812 (N_4812,N_4709,N_4701);
nand U4813 (N_4813,N_4643,N_4671);
and U4814 (N_4814,N_4757,N_4718);
and U4815 (N_4815,N_4710,N_4669);
xnor U4816 (N_4816,N_4630,N_4731);
nand U4817 (N_4817,N_4774,N_4651);
or U4818 (N_4818,N_4716,N_4797);
or U4819 (N_4819,N_4766,N_4747);
and U4820 (N_4820,N_4733,N_4695);
or U4821 (N_4821,N_4642,N_4694);
xor U4822 (N_4822,N_4761,N_4764);
nand U4823 (N_4823,N_4788,N_4667);
or U4824 (N_4824,N_4631,N_4762);
or U4825 (N_4825,N_4613,N_4726);
nand U4826 (N_4826,N_4795,N_4737);
nor U4827 (N_4827,N_4723,N_4711);
and U4828 (N_4828,N_4729,N_4616);
xnor U4829 (N_4829,N_4789,N_4699);
nor U4830 (N_4830,N_4779,N_4753);
or U4831 (N_4831,N_4706,N_4749);
and U4832 (N_4832,N_4689,N_4691);
nand U4833 (N_4833,N_4730,N_4783);
xor U4834 (N_4834,N_4672,N_4647);
or U4835 (N_4835,N_4629,N_4693);
or U4836 (N_4836,N_4639,N_4601);
or U4837 (N_4837,N_4785,N_4717);
nand U4838 (N_4838,N_4649,N_4745);
and U4839 (N_4839,N_4673,N_4721);
and U4840 (N_4840,N_4660,N_4646);
nand U4841 (N_4841,N_4623,N_4659);
or U4842 (N_4842,N_4703,N_4677);
and U4843 (N_4843,N_4775,N_4739);
or U4844 (N_4844,N_4617,N_4713);
and U4845 (N_4845,N_4637,N_4640);
nor U4846 (N_4846,N_4738,N_4678);
xnor U4847 (N_4847,N_4784,N_4606);
nand U4848 (N_4848,N_4635,N_4668);
and U4849 (N_4849,N_4771,N_4732);
nor U4850 (N_4850,N_4690,N_4798);
and U4851 (N_4851,N_4638,N_4687);
and U4852 (N_4852,N_4780,N_4799);
xor U4853 (N_4853,N_4776,N_4611);
and U4854 (N_4854,N_4657,N_4715);
nand U4855 (N_4855,N_4684,N_4670);
nor U4856 (N_4856,N_4750,N_4641);
nor U4857 (N_4857,N_4697,N_4708);
nor U4858 (N_4858,N_4661,N_4792);
or U4859 (N_4859,N_4719,N_4743);
nor U4860 (N_4860,N_4600,N_4692);
xnor U4861 (N_4861,N_4610,N_4712);
xor U4862 (N_4862,N_4787,N_4680);
xnor U4863 (N_4863,N_4790,N_4612);
nand U4864 (N_4864,N_4662,N_4767);
or U4865 (N_4865,N_4603,N_4759);
or U4866 (N_4866,N_4727,N_4796);
or U4867 (N_4867,N_4685,N_4688);
nand U4868 (N_4868,N_4728,N_4621);
or U4869 (N_4869,N_4614,N_4686);
or U4870 (N_4870,N_4791,N_4626);
nor U4871 (N_4871,N_4744,N_4734);
xor U4872 (N_4872,N_4714,N_4676);
xor U4873 (N_4873,N_4607,N_4652);
and U4874 (N_4874,N_4666,N_4696);
or U4875 (N_4875,N_4620,N_4605);
and U4876 (N_4876,N_4754,N_4704);
and U4877 (N_4877,N_4653,N_4702);
and U4878 (N_4878,N_4740,N_4679);
nor U4879 (N_4879,N_4609,N_4633);
and U4880 (N_4880,N_4674,N_4681);
or U4881 (N_4881,N_4650,N_4675);
xor U4882 (N_4882,N_4765,N_4778);
or U4883 (N_4883,N_4741,N_4663);
nand U4884 (N_4884,N_4720,N_4763);
nand U4885 (N_4885,N_4656,N_4773);
or U4886 (N_4886,N_4786,N_4707);
or U4887 (N_4887,N_4628,N_4758);
nor U4888 (N_4888,N_4634,N_4645);
nor U4889 (N_4889,N_4752,N_4700);
nor U4890 (N_4890,N_4793,N_4608);
nand U4891 (N_4891,N_4736,N_4682);
and U4892 (N_4892,N_4769,N_4756);
nor U4893 (N_4893,N_4794,N_4782);
nand U4894 (N_4894,N_4644,N_4636);
nor U4895 (N_4895,N_4683,N_4760);
or U4896 (N_4896,N_4755,N_4627);
nand U4897 (N_4897,N_4725,N_4748);
and U4898 (N_4898,N_4615,N_4664);
nor U4899 (N_4899,N_4624,N_4770);
nor U4900 (N_4900,N_4716,N_4786);
nor U4901 (N_4901,N_4674,N_4784);
nor U4902 (N_4902,N_4715,N_4639);
nor U4903 (N_4903,N_4759,N_4758);
or U4904 (N_4904,N_4642,N_4617);
xor U4905 (N_4905,N_4709,N_4678);
nand U4906 (N_4906,N_4615,N_4652);
or U4907 (N_4907,N_4704,N_4764);
nand U4908 (N_4908,N_4619,N_4604);
and U4909 (N_4909,N_4643,N_4677);
and U4910 (N_4910,N_4686,N_4781);
or U4911 (N_4911,N_4664,N_4723);
nor U4912 (N_4912,N_4795,N_4694);
and U4913 (N_4913,N_4747,N_4685);
nor U4914 (N_4914,N_4660,N_4650);
or U4915 (N_4915,N_4625,N_4710);
or U4916 (N_4916,N_4612,N_4651);
and U4917 (N_4917,N_4784,N_4700);
or U4918 (N_4918,N_4630,N_4750);
and U4919 (N_4919,N_4674,N_4654);
nand U4920 (N_4920,N_4670,N_4735);
or U4921 (N_4921,N_4696,N_4794);
nand U4922 (N_4922,N_4683,N_4667);
and U4923 (N_4923,N_4746,N_4767);
nor U4924 (N_4924,N_4672,N_4742);
nor U4925 (N_4925,N_4692,N_4626);
or U4926 (N_4926,N_4768,N_4641);
nand U4927 (N_4927,N_4707,N_4774);
nor U4928 (N_4928,N_4630,N_4789);
nand U4929 (N_4929,N_4695,N_4604);
or U4930 (N_4930,N_4628,N_4787);
nand U4931 (N_4931,N_4742,N_4653);
or U4932 (N_4932,N_4702,N_4652);
nand U4933 (N_4933,N_4618,N_4642);
nand U4934 (N_4934,N_4637,N_4616);
xnor U4935 (N_4935,N_4698,N_4736);
nand U4936 (N_4936,N_4616,N_4692);
nand U4937 (N_4937,N_4611,N_4795);
xor U4938 (N_4938,N_4767,N_4618);
nor U4939 (N_4939,N_4733,N_4615);
xnor U4940 (N_4940,N_4708,N_4640);
nor U4941 (N_4941,N_4650,N_4654);
and U4942 (N_4942,N_4787,N_4693);
and U4943 (N_4943,N_4626,N_4742);
nand U4944 (N_4944,N_4756,N_4713);
and U4945 (N_4945,N_4774,N_4760);
and U4946 (N_4946,N_4625,N_4701);
and U4947 (N_4947,N_4634,N_4669);
nand U4948 (N_4948,N_4608,N_4615);
or U4949 (N_4949,N_4689,N_4683);
nand U4950 (N_4950,N_4741,N_4738);
nor U4951 (N_4951,N_4778,N_4781);
and U4952 (N_4952,N_4770,N_4667);
nand U4953 (N_4953,N_4777,N_4620);
and U4954 (N_4954,N_4678,N_4752);
nand U4955 (N_4955,N_4618,N_4750);
and U4956 (N_4956,N_4783,N_4782);
and U4957 (N_4957,N_4737,N_4603);
or U4958 (N_4958,N_4663,N_4752);
or U4959 (N_4959,N_4662,N_4627);
nor U4960 (N_4960,N_4727,N_4610);
and U4961 (N_4961,N_4640,N_4745);
or U4962 (N_4962,N_4691,N_4678);
nor U4963 (N_4963,N_4620,N_4696);
or U4964 (N_4964,N_4767,N_4740);
or U4965 (N_4965,N_4716,N_4707);
xnor U4966 (N_4966,N_4685,N_4708);
nor U4967 (N_4967,N_4674,N_4636);
or U4968 (N_4968,N_4632,N_4750);
or U4969 (N_4969,N_4716,N_4603);
nor U4970 (N_4970,N_4680,N_4788);
or U4971 (N_4971,N_4712,N_4604);
nor U4972 (N_4972,N_4659,N_4616);
nor U4973 (N_4973,N_4611,N_4753);
nand U4974 (N_4974,N_4673,N_4792);
nand U4975 (N_4975,N_4639,N_4758);
or U4976 (N_4976,N_4746,N_4763);
nand U4977 (N_4977,N_4614,N_4722);
and U4978 (N_4978,N_4673,N_4647);
nor U4979 (N_4979,N_4647,N_4705);
xnor U4980 (N_4980,N_4600,N_4723);
or U4981 (N_4981,N_4635,N_4687);
nor U4982 (N_4982,N_4671,N_4677);
nor U4983 (N_4983,N_4765,N_4780);
or U4984 (N_4984,N_4610,N_4796);
or U4985 (N_4985,N_4706,N_4757);
nand U4986 (N_4986,N_4770,N_4773);
or U4987 (N_4987,N_4768,N_4718);
and U4988 (N_4988,N_4713,N_4685);
and U4989 (N_4989,N_4767,N_4789);
xor U4990 (N_4990,N_4705,N_4759);
nor U4991 (N_4991,N_4795,N_4725);
xnor U4992 (N_4992,N_4703,N_4742);
nand U4993 (N_4993,N_4669,N_4684);
nor U4994 (N_4994,N_4648,N_4785);
or U4995 (N_4995,N_4749,N_4726);
nand U4996 (N_4996,N_4704,N_4782);
and U4997 (N_4997,N_4655,N_4600);
or U4998 (N_4998,N_4698,N_4638);
and U4999 (N_4999,N_4790,N_4721);
nand UO_0 (O_0,N_4915,N_4821);
nor UO_1 (O_1,N_4959,N_4858);
nand UO_2 (O_2,N_4887,N_4846);
or UO_3 (O_3,N_4852,N_4820);
and UO_4 (O_4,N_4929,N_4981);
nand UO_5 (O_5,N_4965,N_4902);
nand UO_6 (O_6,N_4864,N_4810);
and UO_7 (O_7,N_4878,N_4939);
nand UO_8 (O_8,N_4917,N_4885);
xor UO_9 (O_9,N_4946,N_4963);
nand UO_10 (O_10,N_4900,N_4932);
or UO_11 (O_11,N_4837,N_4960);
nor UO_12 (O_12,N_4997,N_4854);
or UO_13 (O_13,N_4899,N_4978);
or UO_14 (O_14,N_4947,N_4862);
nand UO_15 (O_15,N_4880,N_4905);
or UO_16 (O_16,N_4800,N_4814);
and UO_17 (O_17,N_4881,N_4839);
and UO_18 (O_18,N_4938,N_4896);
nor UO_19 (O_19,N_4971,N_4955);
or UO_20 (O_20,N_4891,N_4926);
and UO_21 (O_21,N_4974,N_4865);
and UO_22 (O_22,N_4913,N_4819);
or UO_23 (O_23,N_4961,N_4859);
nor UO_24 (O_24,N_4931,N_4910);
or UO_25 (O_25,N_4869,N_4822);
and UO_26 (O_26,N_4901,N_4990);
nor UO_27 (O_27,N_4970,N_4906);
nand UO_28 (O_28,N_4824,N_4841);
and UO_29 (O_29,N_4886,N_4924);
xnor UO_30 (O_30,N_4835,N_4874);
or UO_31 (O_31,N_4879,N_4801);
and UO_32 (O_32,N_4934,N_4979);
nor UO_33 (O_33,N_4999,N_4956);
or UO_34 (O_34,N_4920,N_4912);
nand UO_35 (O_35,N_4830,N_4969);
and UO_36 (O_36,N_4804,N_4948);
xnor UO_37 (O_37,N_4903,N_4923);
xor UO_38 (O_38,N_4987,N_4895);
nor UO_39 (O_39,N_4855,N_4823);
or UO_40 (O_40,N_4863,N_4828);
or UO_41 (O_41,N_4953,N_4911);
nand UO_42 (O_42,N_4893,N_4817);
nand UO_43 (O_43,N_4843,N_4840);
nor UO_44 (O_44,N_4836,N_4838);
xor UO_45 (O_45,N_4827,N_4894);
and UO_46 (O_46,N_4813,N_4952);
nand UO_47 (O_47,N_4832,N_4847);
xnor UO_48 (O_48,N_4861,N_4933);
or UO_49 (O_49,N_4940,N_4802);
nor UO_50 (O_50,N_4921,N_4857);
nand UO_51 (O_51,N_4908,N_4851);
xor UO_52 (O_52,N_4898,N_4972);
and UO_53 (O_53,N_4909,N_4882);
nor UO_54 (O_54,N_4950,N_4811);
and UO_55 (O_55,N_4991,N_4975);
xnor UO_56 (O_56,N_4935,N_4967);
nand UO_57 (O_57,N_4809,N_4871);
nor UO_58 (O_58,N_4983,N_4829);
nand UO_59 (O_59,N_4844,N_4890);
nor UO_60 (O_60,N_4985,N_4848);
or UO_61 (O_61,N_4925,N_4936);
nor UO_62 (O_62,N_4989,N_4945);
or UO_63 (O_63,N_4966,N_4995);
nand UO_64 (O_64,N_4977,N_4842);
nand UO_65 (O_65,N_4876,N_4976);
and UO_66 (O_66,N_4954,N_4941);
and UO_67 (O_67,N_4870,N_4922);
xnor UO_68 (O_68,N_4884,N_4872);
and UO_69 (O_69,N_4888,N_4943);
nor UO_70 (O_70,N_4928,N_4850);
nand UO_71 (O_71,N_4867,N_4805);
and UO_72 (O_72,N_4986,N_4868);
xor UO_73 (O_73,N_4973,N_4951);
nor UO_74 (O_74,N_4988,N_4992);
nor UO_75 (O_75,N_4942,N_4815);
xor UO_76 (O_76,N_4834,N_4918);
or UO_77 (O_77,N_4944,N_4845);
nand UO_78 (O_78,N_4826,N_4873);
or UO_79 (O_79,N_4853,N_4883);
nor UO_80 (O_80,N_4833,N_4807);
and UO_81 (O_81,N_4993,N_4904);
xnor UO_82 (O_82,N_4927,N_4964);
nand UO_83 (O_83,N_4968,N_4892);
nand UO_84 (O_84,N_4919,N_4994);
and UO_85 (O_85,N_4860,N_4875);
nand UO_86 (O_86,N_4877,N_4949);
and UO_87 (O_87,N_4856,N_4825);
xnor UO_88 (O_88,N_4808,N_4958);
and UO_89 (O_89,N_4996,N_4907);
nand UO_90 (O_90,N_4982,N_4831);
xnor UO_91 (O_91,N_4930,N_4937);
and UO_92 (O_92,N_4998,N_4914);
and UO_93 (O_93,N_4889,N_4957);
or UO_94 (O_94,N_4984,N_4897);
and UO_95 (O_95,N_4866,N_4812);
nor UO_96 (O_96,N_4962,N_4916);
nand UO_97 (O_97,N_4980,N_4849);
or UO_98 (O_98,N_4803,N_4816);
nor UO_99 (O_99,N_4818,N_4806);
nor UO_100 (O_100,N_4961,N_4813);
nand UO_101 (O_101,N_4827,N_4829);
nand UO_102 (O_102,N_4996,N_4915);
or UO_103 (O_103,N_4806,N_4873);
nand UO_104 (O_104,N_4915,N_4872);
and UO_105 (O_105,N_4827,N_4916);
or UO_106 (O_106,N_4854,N_4912);
and UO_107 (O_107,N_4951,N_4926);
nand UO_108 (O_108,N_4800,N_4946);
or UO_109 (O_109,N_4819,N_4911);
and UO_110 (O_110,N_4978,N_4802);
xnor UO_111 (O_111,N_4890,N_4958);
or UO_112 (O_112,N_4813,N_4842);
and UO_113 (O_113,N_4833,N_4879);
or UO_114 (O_114,N_4860,N_4969);
nand UO_115 (O_115,N_4895,N_4950);
nor UO_116 (O_116,N_4895,N_4856);
nor UO_117 (O_117,N_4973,N_4835);
xor UO_118 (O_118,N_4989,N_4841);
xnor UO_119 (O_119,N_4897,N_4813);
nand UO_120 (O_120,N_4977,N_4997);
or UO_121 (O_121,N_4829,N_4914);
and UO_122 (O_122,N_4965,N_4933);
and UO_123 (O_123,N_4817,N_4939);
nor UO_124 (O_124,N_4856,N_4806);
and UO_125 (O_125,N_4804,N_4999);
and UO_126 (O_126,N_4931,N_4926);
and UO_127 (O_127,N_4867,N_4975);
and UO_128 (O_128,N_4801,N_4872);
or UO_129 (O_129,N_4917,N_4985);
and UO_130 (O_130,N_4937,N_4882);
nand UO_131 (O_131,N_4962,N_4825);
nor UO_132 (O_132,N_4903,N_4925);
or UO_133 (O_133,N_4873,N_4922);
or UO_134 (O_134,N_4919,N_4901);
xor UO_135 (O_135,N_4924,N_4884);
nor UO_136 (O_136,N_4890,N_4823);
nand UO_137 (O_137,N_4815,N_4985);
nand UO_138 (O_138,N_4812,N_4930);
or UO_139 (O_139,N_4889,N_4848);
nor UO_140 (O_140,N_4946,N_4834);
xor UO_141 (O_141,N_4999,N_4866);
nor UO_142 (O_142,N_4846,N_4836);
or UO_143 (O_143,N_4954,N_4988);
nor UO_144 (O_144,N_4835,N_4878);
nand UO_145 (O_145,N_4986,N_4822);
nor UO_146 (O_146,N_4843,N_4999);
and UO_147 (O_147,N_4841,N_4994);
or UO_148 (O_148,N_4925,N_4878);
nand UO_149 (O_149,N_4910,N_4800);
nand UO_150 (O_150,N_4971,N_4967);
nand UO_151 (O_151,N_4879,N_4815);
nand UO_152 (O_152,N_4944,N_4808);
and UO_153 (O_153,N_4980,N_4830);
or UO_154 (O_154,N_4913,N_4882);
nor UO_155 (O_155,N_4916,N_4988);
and UO_156 (O_156,N_4818,N_4984);
or UO_157 (O_157,N_4868,N_4944);
nor UO_158 (O_158,N_4913,N_4916);
nand UO_159 (O_159,N_4858,N_4948);
nand UO_160 (O_160,N_4899,N_4994);
nor UO_161 (O_161,N_4894,N_4884);
nand UO_162 (O_162,N_4922,N_4846);
nor UO_163 (O_163,N_4948,N_4852);
nor UO_164 (O_164,N_4807,N_4953);
nand UO_165 (O_165,N_4826,N_4870);
nand UO_166 (O_166,N_4927,N_4996);
xnor UO_167 (O_167,N_4829,N_4845);
nor UO_168 (O_168,N_4818,N_4869);
nor UO_169 (O_169,N_4845,N_4918);
nor UO_170 (O_170,N_4905,N_4911);
nor UO_171 (O_171,N_4916,N_4869);
and UO_172 (O_172,N_4988,N_4973);
xnor UO_173 (O_173,N_4877,N_4952);
and UO_174 (O_174,N_4974,N_4976);
nor UO_175 (O_175,N_4917,N_4979);
nor UO_176 (O_176,N_4935,N_4988);
or UO_177 (O_177,N_4865,N_4822);
or UO_178 (O_178,N_4900,N_4870);
and UO_179 (O_179,N_4977,N_4862);
nor UO_180 (O_180,N_4817,N_4987);
xnor UO_181 (O_181,N_4901,N_4876);
and UO_182 (O_182,N_4923,N_4965);
nor UO_183 (O_183,N_4974,N_4906);
or UO_184 (O_184,N_4941,N_4912);
or UO_185 (O_185,N_4800,N_4833);
nand UO_186 (O_186,N_4913,N_4892);
nand UO_187 (O_187,N_4804,N_4980);
xor UO_188 (O_188,N_4987,N_4901);
and UO_189 (O_189,N_4836,N_4998);
nor UO_190 (O_190,N_4841,N_4969);
nor UO_191 (O_191,N_4929,N_4820);
and UO_192 (O_192,N_4964,N_4872);
nand UO_193 (O_193,N_4995,N_4811);
xnor UO_194 (O_194,N_4820,N_4955);
nand UO_195 (O_195,N_4972,N_4948);
xnor UO_196 (O_196,N_4993,N_4954);
or UO_197 (O_197,N_4932,N_4925);
nor UO_198 (O_198,N_4982,N_4910);
nor UO_199 (O_199,N_4920,N_4904);
nand UO_200 (O_200,N_4960,N_4948);
or UO_201 (O_201,N_4893,N_4992);
and UO_202 (O_202,N_4999,N_4990);
nor UO_203 (O_203,N_4891,N_4855);
or UO_204 (O_204,N_4849,N_4976);
nand UO_205 (O_205,N_4951,N_4940);
and UO_206 (O_206,N_4900,N_4859);
nor UO_207 (O_207,N_4920,N_4894);
and UO_208 (O_208,N_4861,N_4803);
nor UO_209 (O_209,N_4857,N_4831);
and UO_210 (O_210,N_4926,N_4842);
and UO_211 (O_211,N_4814,N_4820);
nand UO_212 (O_212,N_4827,N_4921);
xnor UO_213 (O_213,N_4922,N_4857);
and UO_214 (O_214,N_4930,N_4913);
nor UO_215 (O_215,N_4885,N_4859);
and UO_216 (O_216,N_4806,N_4947);
and UO_217 (O_217,N_4854,N_4987);
nand UO_218 (O_218,N_4883,N_4861);
nand UO_219 (O_219,N_4979,N_4855);
and UO_220 (O_220,N_4892,N_4948);
and UO_221 (O_221,N_4909,N_4968);
or UO_222 (O_222,N_4884,N_4945);
nand UO_223 (O_223,N_4959,N_4839);
nand UO_224 (O_224,N_4959,N_4889);
and UO_225 (O_225,N_4925,N_4846);
nand UO_226 (O_226,N_4919,N_4899);
or UO_227 (O_227,N_4870,N_4925);
and UO_228 (O_228,N_4944,N_4937);
and UO_229 (O_229,N_4837,N_4853);
xnor UO_230 (O_230,N_4910,N_4952);
and UO_231 (O_231,N_4819,N_4914);
xnor UO_232 (O_232,N_4999,N_4860);
and UO_233 (O_233,N_4895,N_4913);
or UO_234 (O_234,N_4985,N_4850);
or UO_235 (O_235,N_4917,N_4932);
and UO_236 (O_236,N_4894,N_4971);
nor UO_237 (O_237,N_4860,N_4950);
or UO_238 (O_238,N_4961,N_4957);
xnor UO_239 (O_239,N_4897,N_4971);
or UO_240 (O_240,N_4937,N_4822);
nor UO_241 (O_241,N_4801,N_4916);
xor UO_242 (O_242,N_4992,N_4873);
nand UO_243 (O_243,N_4862,N_4972);
nand UO_244 (O_244,N_4860,N_4925);
and UO_245 (O_245,N_4821,N_4926);
or UO_246 (O_246,N_4890,N_4956);
nand UO_247 (O_247,N_4862,N_4845);
nor UO_248 (O_248,N_4979,N_4809);
and UO_249 (O_249,N_4930,N_4873);
and UO_250 (O_250,N_4817,N_4866);
nor UO_251 (O_251,N_4930,N_4942);
and UO_252 (O_252,N_4802,N_4839);
or UO_253 (O_253,N_4943,N_4835);
and UO_254 (O_254,N_4880,N_4942);
nor UO_255 (O_255,N_4845,N_4910);
and UO_256 (O_256,N_4815,N_4902);
and UO_257 (O_257,N_4956,N_4809);
nand UO_258 (O_258,N_4914,N_4894);
nand UO_259 (O_259,N_4800,N_4922);
or UO_260 (O_260,N_4813,N_4997);
nand UO_261 (O_261,N_4818,N_4808);
and UO_262 (O_262,N_4922,N_4973);
xor UO_263 (O_263,N_4993,N_4840);
nand UO_264 (O_264,N_4844,N_4917);
nand UO_265 (O_265,N_4987,N_4983);
nor UO_266 (O_266,N_4984,N_4935);
or UO_267 (O_267,N_4828,N_4997);
and UO_268 (O_268,N_4895,N_4830);
nor UO_269 (O_269,N_4986,N_4852);
and UO_270 (O_270,N_4826,N_4986);
and UO_271 (O_271,N_4841,N_4840);
or UO_272 (O_272,N_4855,N_4915);
and UO_273 (O_273,N_4974,N_4964);
and UO_274 (O_274,N_4950,N_4888);
or UO_275 (O_275,N_4951,N_4857);
nor UO_276 (O_276,N_4856,N_4823);
and UO_277 (O_277,N_4825,N_4905);
nand UO_278 (O_278,N_4956,N_4850);
nor UO_279 (O_279,N_4907,N_4858);
nor UO_280 (O_280,N_4978,N_4847);
or UO_281 (O_281,N_4907,N_4975);
nor UO_282 (O_282,N_4909,N_4826);
or UO_283 (O_283,N_4807,N_4906);
or UO_284 (O_284,N_4853,N_4836);
nand UO_285 (O_285,N_4956,N_4954);
nand UO_286 (O_286,N_4847,N_4819);
and UO_287 (O_287,N_4929,N_4992);
nand UO_288 (O_288,N_4930,N_4934);
nand UO_289 (O_289,N_4974,N_4857);
xnor UO_290 (O_290,N_4995,N_4946);
nand UO_291 (O_291,N_4884,N_4881);
nand UO_292 (O_292,N_4910,N_4993);
nand UO_293 (O_293,N_4833,N_4910);
nor UO_294 (O_294,N_4854,N_4969);
or UO_295 (O_295,N_4995,N_4898);
or UO_296 (O_296,N_4891,N_4854);
nand UO_297 (O_297,N_4831,N_4821);
or UO_298 (O_298,N_4824,N_4831);
nand UO_299 (O_299,N_4809,N_4907);
and UO_300 (O_300,N_4974,N_4951);
and UO_301 (O_301,N_4902,N_4891);
xor UO_302 (O_302,N_4946,N_4951);
nor UO_303 (O_303,N_4958,N_4818);
or UO_304 (O_304,N_4904,N_4934);
nand UO_305 (O_305,N_4815,N_4923);
and UO_306 (O_306,N_4870,N_4848);
or UO_307 (O_307,N_4983,N_4868);
nand UO_308 (O_308,N_4969,N_4817);
xor UO_309 (O_309,N_4876,N_4839);
nor UO_310 (O_310,N_4907,N_4890);
xor UO_311 (O_311,N_4987,N_4992);
nand UO_312 (O_312,N_4954,N_4892);
and UO_313 (O_313,N_4843,N_4938);
and UO_314 (O_314,N_4841,N_4819);
and UO_315 (O_315,N_4959,N_4866);
nor UO_316 (O_316,N_4917,N_4957);
or UO_317 (O_317,N_4960,N_4971);
xor UO_318 (O_318,N_4843,N_4967);
nor UO_319 (O_319,N_4922,N_4926);
and UO_320 (O_320,N_4884,N_4931);
nand UO_321 (O_321,N_4927,N_4916);
nor UO_322 (O_322,N_4995,N_4800);
and UO_323 (O_323,N_4988,N_4871);
nand UO_324 (O_324,N_4856,N_4926);
nor UO_325 (O_325,N_4826,N_4847);
or UO_326 (O_326,N_4858,N_4887);
nor UO_327 (O_327,N_4868,N_4962);
and UO_328 (O_328,N_4973,N_4826);
nor UO_329 (O_329,N_4835,N_4942);
and UO_330 (O_330,N_4944,N_4995);
nand UO_331 (O_331,N_4952,N_4931);
xnor UO_332 (O_332,N_4891,N_4851);
nand UO_333 (O_333,N_4923,N_4805);
and UO_334 (O_334,N_4909,N_4925);
and UO_335 (O_335,N_4827,N_4875);
nor UO_336 (O_336,N_4922,N_4899);
nand UO_337 (O_337,N_4904,N_4826);
or UO_338 (O_338,N_4950,N_4836);
nor UO_339 (O_339,N_4963,N_4887);
or UO_340 (O_340,N_4901,N_4815);
nand UO_341 (O_341,N_4810,N_4972);
or UO_342 (O_342,N_4909,N_4865);
or UO_343 (O_343,N_4998,N_4833);
nor UO_344 (O_344,N_4846,N_4820);
nand UO_345 (O_345,N_4831,N_4890);
nor UO_346 (O_346,N_4831,N_4986);
xnor UO_347 (O_347,N_4826,N_4969);
and UO_348 (O_348,N_4956,N_4831);
or UO_349 (O_349,N_4912,N_4992);
xnor UO_350 (O_350,N_4912,N_4931);
or UO_351 (O_351,N_4998,N_4802);
and UO_352 (O_352,N_4874,N_4946);
or UO_353 (O_353,N_4807,N_4936);
nand UO_354 (O_354,N_4916,N_4937);
or UO_355 (O_355,N_4974,N_4919);
and UO_356 (O_356,N_4925,N_4929);
nor UO_357 (O_357,N_4806,N_4925);
xor UO_358 (O_358,N_4816,N_4986);
nor UO_359 (O_359,N_4989,N_4871);
or UO_360 (O_360,N_4902,N_4936);
and UO_361 (O_361,N_4978,N_4897);
xnor UO_362 (O_362,N_4924,N_4882);
nand UO_363 (O_363,N_4995,N_4805);
and UO_364 (O_364,N_4929,N_4893);
nor UO_365 (O_365,N_4847,N_4924);
nand UO_366 (O_366,N_4809,N_4855);
nor UO_367 (O_367,N_4829,N_4952);
nor UO_368 (O_368,N_4944,N_4893);
nand UO_369 (O_369,N_4989,N_4817);
and UO_370 (O_370,N_4993,N_4858);
nand UO_371 (O_371,N_4937,N_4973);
and UO_372 (O_372,N_4949,N_4803);
xnor UO_373 (O_373,N_4807,N_4956);
nor UO_374 (O_374,N_4953,N_4861);
xnor UO_375 (O_375,N_4907,N_4909);
nor UO_376 (O_376,N_4858,N_4912);
nor UO_377 (O_377,N_4967,N_4864);
and UO_378 (O_378,N_4951,N_4855);
and UO_379 (O_379,N_4935,N_4920);
nand UO_380 (O_380,N_4871,N_4875);
or UO_381 (O_381,N_4846,N_4842);
and UO_382 (O_382,N_4877,N_4859);
xnor UO_383 (O_383,N_4817,N_4825);
nand UO_384 (O_384,N_4866,N_4820);
nand UO_385 (O_385,N_4927,N_4899);
nand UO_386 (O_386,N_4897,N_4960);
xor UO_387 (O_387,N_4955,N_4861);
nor UO_388 (O_388,N_4809,N_4808);
or UO_389 (O_389,N_4924,N_4853);
xor UO_390 (O_390,N_4993,N_4901);
and UO_391 (O_391,N_4879,N_4922);
nor UO_392 (O_392,N_4971,N_4925);
or UO_393 (O_393,N_4815,N_4917);
and UO_394 (O_394,N_4904,N_4880);
and UO_395 (O_395,N_4919,N_4906);
or UO_396 (O_396,N_4886,N_4822);
xor UO_397 (O_397,N_4801,N_4868);
and UO_398 (O_398,N_4968,N_4875);
nor UO_399 (O_399,N_4853,N_4882);
xor UO_400 (O_400,N_4819,N_4921);
or UO_401 (O_401,N_4903,N_4883);
xnor UO_402 (O_402,N_4861,N_4898);
and UO_403 (O_403,N_4837,N_4924);
nor UO_404 (O_404,N_4891,N_4886);
or UO_405 (O_405,N_4919,N_4811);
and UO_406 (O_406,N_4947,N_4923);
xor UO_407 (O_407,N_4842,N_4942);
and UO_408 (O_408,N_4865,N_4931);
and UO_409 (O_409,N_4879,N_4970);
nor UO_410 (O_410,N_4835,N_4979);
nand UO_411 (O_411,N_4880,N_4953);
xnor UO_412 (O_412,N_4904,N_4824);
or UO_413 (O_413,N_4805,N_4888);
nor UO_414 (O_414,N_4902,N_4904);
or UO_415 (O_415,N_4926,N_4997);
nand UO_416 (O_416,N_4928,N_4905);
xnor UO_417 (O_417,N_4818,N_4860);
or UO_418 (O_418,N_4832,N_4960);
nand UO_419 (O_419,N_4819,N_4970);
nor UO_420 (O_420,N_4952,N_4851);
nand UO_421 (O_421,N_4847,N_4804);
nand UO_422 (O_422,N_4875,N_4994);
nor UO_423 (O_423,N_4943,N_4912);
nand UO_424 (O_424,N_4842,N_4835);
nor UO_425 (O_425,N_4850,N_4821);
xnor UO_426 (O_426,N_4992,N_4976);
nand UO_427 (O_427,N_4873,N_4804);
nand UO_428 (O_428,N_4811,N_4882);
and UO_429 (O_429,N_4925,N_4919);
nand UO_430 (O_430,N_4963,N_4956);
or UO_431 (O_431,N_4872,N_4878);
and UO_432 (O_432,N_4943,N_4807);
nor UO_433 (O_433,N_4952,N_4891);
nand UO_434 (O_434,N_4848,N_4860);
nor UO_435 (O_435,N_4989,N_4983);
or UO_436 (O_436,N_4992,N_4839);
nand UO_437 (O_437,N_4918,N_4917);
nand UO_438 (O_438,N_4813,N_4994);
or UO_439 (O_439,N_4862,N_4980);
and UO_440 (O_440,N_4992,N_4814);
xor UO_441 (O_441,N_4847,N_4855);
xnor UO_442 (O_442,N_4844,N_4945);
nor UO_443 (O_443,N_4989,N_4881);
nand UO_444 (O_444,N_4825,N_4819);
nand UO_445 (O_445,N_4839,N_4979);
nand UO_446 (O_446,N_4803,N_4827);
and UO_447 (O_447,N_4946,N_4957);
and UO_448 (O_448,N_4996,N_4816);
nand UO_449 (O_449,N_4891,N_4969);
nand UO_450 (O_450,N_4919,N_4873);
xnor UO_451 (O_451,N_4999,N_4895);
nand UO_452 (O_452,N_4945,N_4858);
nand UO_453 (O_453,N_4821,N_4805);
or UO_454 (O_454,N_4815,N_4838);
xor UO_455 (O_455,N_4994,N_4983);
nor UO_456 (O_456,N_4804,N_4866);
or UO_457 (O_457,N_4818,N_4886);
xor UO_458 (O_458,N_4923,N_4877);
nand UO_459 (O_459,N_4905,N_4857);
nor UO_460 (O_460,N_4806,N_4984);
or UO_461 (O_461,N_4800,N_4926);
or UO_462 (O_462,N_4801,N_4800);
and UO_463 (O_463,N_4879,N_4895);
and UO_464 (O_464,N_4833,N_4957);
or UO_465 (O_465,N_4962,N_4992);
nor UO_466 (O_466,N_4870,N_4957);
nor UO_467 (O_467,N_4842,N_4811);
and UO_468 (O_468,N_4852,N_4865);
nor UO_469 (O_469,N_4856,N_4871);
or UO_470 (O_470,N_4829,N_4873);
nor UO_471 (O_471,N_4802,N_4872);
nor UO_472 (O_472,N_4954,N_4898);
and UO_473 (O_473,N_4810,N_4898);
nand UO_474 (O_474,N_4897,N_4908);
and UO_475 (O_475,N_4912,N_4813);
or UO_476 (O_476,N_4989,N_4961);
nand UO_477 (O_477,N_4954,N_4952);
or UO_478 (O_478,N_4986,N_4973);
or UO_479 (O_479,N_4824,N_4900);
or UO_480 (O_480,N_4852,N_4859);
nand UO_481 (O_481,N_4912,N_4897);
nand UO_482 (O_482,N_4848,N_4917);
xor UO_483 (O_483,N_4814,N_4931);
or UO_484 (O_484,N_4965,N_4858);
or UO_485 (O_485,N_4826,N_4958);
and UO_486 (O_486,N_4805,N_4807);
nor UO_487 (O_487,N_4803,N_4865);
nand UO_488 (O_488,N_4969,N_4896);
nor UO_489 (O_489,N_4882,N_4879);
or UO_490 (O_490,N_4886,N_4828);
and UO_491 (O_491,N_4980,N_4822);
and UO_492 (O_492,N_4919,N_4815);
and UO_493 (O_493,N_4843,N_4872);
nor UO_494 (O_494,N_4962,N_4986);
nor UO_495 (O_495,N_4842,N_4869);
and UO_496 (O_496,N_4942,N_4803);
or UO_497 (O_497,N_4837,N_4920);
and UO_498 (O_498,N_4979,N_4908);
nand UO_499 (O_499,N_4875,N_4867);
and UO_500 (O_500,N_4933,N_4959);
nor UO_501 (O_501,N_4969,N_4958);
and UO_502 (O_502,N_4943,N_4986);
nor UO_503 (O_503,N_4983,N_4905);
nand UO_504 (O_504,N_4926,N_4937);
nor UO_505 (O_505,N_4960,N_4899);
xor UO_506 (O_506,N_4987,N_4829);
nand UO_507 (O_507,N_4996,N_4904);
or UO_508 (O_508,N_4987,N_4980);
xor UO_509 (O_509,N_4950,N_4875);
and UO_510 (O_510,N_4952,N_4908);
or UO_511 (O_511,N_4815,N_4980);
xor UO_512 (O_512,N_4930,N_4811);
or UO_513 (O_513,N_4872,N_4831);
nor UO_514 (O_514,N_4829,N_4881);
nor UO_515 (O_515,N_4999,N_4877);
nor UO_516 (O_516,N_4983,N_4883);
nand UO_517 (O_517,N_4888,N_4912);
or UO_518 (O_518,N_4970,N_4890);
xor UO_519 (O_519,N_4986,N_4896);
and UO_520 (O_520,N_4967,N_4982);
and UO_521 (O_521,N_4854,N_4923);
nor UO_522 (O_522,N_4945,N_4846);
xnor UO_523 (O_523,N_4938,N_4998);
and UO_524 (O_524,N_4802,N_4917);
xor UO_525 (O_525,N_4829,N_4860);
nor UO_526 (O_526,N_4899,N_4824);
nand UO_527 (O_527,N_4903,N_4922);
and UO_528 (O_528,N_4901,N_4879);
nor UO_529 (O_529,N_4857,N_4836);
and UO_530 (O_530,N_4944,N_4814);
nand UO_531 (O_531,N_4919,N_4930);
and UO_532 (O_532,N_4867,N_4998);
nor UO_533 (O_533,N_4996,N_4899);
nand UO_534 (O_534,N_4835,N_4805);
and UO_535 (O_535,N_4980,N_4854);
and UO_536 (O_536,N_4919,N_4910);
or UO_537 (O_537,N_4834,N_4954);
and UO_538 (O_538,N_4808,N_4870);
nor UO_539 (O_539,N_4808,N_4976);
or UO_540 (O_540,N_4935,N_4978);
or UO_541 (O_541,N_4966,N_4977);
or UO_542 (O_542,N_4912,N_4910);
and UO_543 (O_543,N_4804,N_4933);
nor UO_544 (O_544,N_4848,N_4807);
and UO_545 (O_545,N_4831,N_4989);
nor UO_546 (O_546,N_4830,N_4909);
xnor UO_547 (O_547,N_4998,N_4818);
nor UO_548 (O_548,N_4920,N_4821);
nand UO_549 (O_549,N_4864,N_4922);
xor UO_550 (O_550,N_4953,N_4959);
nand UO_551 (O_551,N_4893,N_4964);
or UO_552 (O_552,N_4973,N_4901);
nor UO_553 (O_553,N_4963,N_4901);
xor UO_554 (O_554,N_4947,N_4913);
or UO_555 (O_555,N_4966,N_4885);
or UO_556 (O_556,N_4830,N_4801);
xor UO_557 (O_557,N_4994,N_4944);
xor UO_558 (O_558,N_4937,N_4962);
and UO_559 (O_559,N_4957,N_4842);
or UO_560 (O_560,N_4878,N_4988);
nor UO_561 (O_561,N_4912,N_4803);
nor UO_562 (O_562,N_4993,N_4964);
nand UO_563 (O_563,N_4868,N_4967);
and UO_564 (O_564,N_4943,N_4944);
or UO_565 (O_565,N_4987,N_4916);
and UO_566 (O_566,N_4912,N_4856);
nand UO_567 (O_567,N_4865,N_4895);
nand UO_568 (O_568,N_4825,N_4940);
and UO_569 (O_569,N_4931,N_4860);
xor UO_570 (O_570,N_4980,N_4843);
nor UO_571 (O_571,N_4971,N_4840);
nand UO_572 (O_572,N_4808,N_4929);
xor UO_573 (O_573,N_4870,N_4946);
and UO_574 (O_574,N_4886,N_4866);
or UO_575 (O_575,N_4965,N_4910);
and UO_576 (O_576,N_4921,N_4853);
nor UO_577 (O_577,N_4812,N_4819);
nand UO_578 (O_578,N_4947,N_4985);
nor UO_579 (O_579,N_4906,N_4966);
nor UO_580 (O_580,N_4865,N_4845);
and UO_581 (O_581,N_4858,N_4835);
and UO_582 (O_582,N_4875,N_4927);
nor UO_583 (O_583,N_4984,N_4837);
nand UO_584 (O_584,N_4815,N_4868);
xor UO_585 (O_585,N_4848,N_4955);
xnor UO_586 (O_586,N_4944,N_4910);
xor UO_587 (O_587,N_4840,N_4858);
or UO_588 (O_588,N_4918,N_4907);
and UO_589 (O_589,N_4909,N_4998);
and UO_590 (O_590,N_4970,N_4921);
or UO_591 (O_591,N_4802,N_4881);
and UO_592 (O_592,N_4823,N_4814);
or UO_593 (O_593,N_4833,N_4966);
xor UO_594 (O_594,N_4948,N_4815);
nand UO_595 (O_595,N_4938,N_4919);
or UO_596 (O_596,N_4991,N_4879);
or UO_597 (O_597,N_4814,N_4821);
nand UO_598 (O_598,N_4941,N_4976);
nor UO_599 (O_599,N_4811,N_4812);
nand UO_600 (O_600,N_4841,N_4868);
nand UO_601 (O_601,N_4877,N_4910);
nor UO_602 (O_602,N_4899,N_4835);
and UO_603 (O_603,N_4903,N_4878);
and UO_604 (O_604,N_4930,N_4965);
nand UO_605 (O_605,N_4899,N_4997);
and UO_606 (O_606,N_4986,N_4981);
nor UO_607 (O_607,N_4928,N_4813);
or UO_608 (O_608,N_4845,N_4806);
nor UO_609 (O_609,N_4858,N_4863);
nand UO_610 (O_610,N_4822,N_4845);
or UO_611 (O_611,N_4824,N_4819);
nor UO_612 (O_612,N_4999,N_4963);
and UO_613 (O_613,N_4892,N_4945);
xnor UO_614 (O_614,N_4952,N_4957);
or UO_615 (O_615,N_4830,N_4833);
and UO_616 (O_616,N_4857,N_4891);
or UO_617 (O_617,N_4898,N_4917);
and UO_618 (O_618,N_4888,N_4902);
nor UO_619 (O_619,N_4864,N_4901);
or UO_620 (O_620,N_4948,N_4918);
and UO_621 (O_621,N_4810,N_4919);
nand UO_622 (O_622,N_4806,N_4969);
xnor UO_623 (O_623,N_4933,N_4846);
or UO_624 (O_624,N_4941,N_4952);
nor UO_625 (O_625,N_4992,N_4910);
xnor UO_626 (O_626,N_4845,N_4950);
or UO_627 (O_627,N_4803,N_4878);
and UO_628 (O_628,N_4923,N_4881);
xor UO_629 (O_629,N_4852,N_4927);
nor UO_630 (O_630,N_4956,N_4976);
nand UO_631 (O_631,N_4933,N_4978);
and UO_632 (O_632,N_4841,N_4870);
nand UO_633 (O_633,N_4875,N_4975);
and UO_634 (O_634,N_4867,N_4874);
or UO_635 (O_635,N_4817,N_4922);
or UO_636 (O_636,N_4871,N_4953);
nor UO_637 (O_637,N_4997,N_4871);
nor UO_638 (O_638,N_4980,N_4970);
nor UO_639 (O_639,N_4957,N_4910);
nand UO_640 (O_640,N_4894,N_4885);
xnor UO_641 (O_641,N_4969,N_4919);
xor UO_642 (O_642,N_4974,N_4928);
or UO_643 (O_643,N_4992,N_4858);
nor UO_644 (O_644,N_4934,N_4801);
and UO_645 (O_645,N_4891,N_4945);
or UO_646 (O_646,N_4948,N_4959);
or UO_647 (O_647,N_4940,N_4932);
nand UO_648 (O_648,N_4828,N_4957);
nor UO_649 (O_649,N_4847,N_4983);
or UO_650 (O_650,N_4989,N_4900);
nand UO_651 (O_651,N_4885,N_4801);
nor UO_652 (O_652,N_4962,N_4927);
and UO_653 (O_653,N_4967,N_4863);
and UO_654 (O_654,N_4963,N_4957);
or UO_655 (O_655,N_4980,N_4891);
nor UO_656 (O_656,N_4934,N_4967);
and UO_657 (O_657,N_4982,N_4937);
or UO_658 (O_658,N_4958,N_4909);
or UO_659 (O_659,N_4882,N_4985);
nand UO_660 (O_660,N_4915,N_4930);
nor UO_661 (O_661,N_4916,N_4838);
nor UO_662 (O_662,N_4951,N_4815);
xnor UO_663 (O_663,N_4877,N_4885);
or UO_664 (O_664,N_4882,N_4992);
or UO_665 (O_665,N_4958,N_4876);
and UO_666 (O_666,N_4864,N_4949);
or UO_667 (O_667,N_4968,N_4881);
xor UO_668 (O_668,N_4953,N_4918);
and UO_669 (O_669,N_4853,N_4986);
nand UO_670 (O_670,N_4863,N_4988);
or UO_671 (O_671,N_4838,N_4858);
nand UO_672 (O_672,N_4844,N_4838);
nand UO_673 (O_673,N_4903,N_4909);
nand UO_674 (O_674,N_4995,N_4940);
and UO_675 (O_675,N_4864,N_4894);
xnor UO_676 (O_676,N_4903,N_4836);
xnor UO_677 (O_677,N_4987,N_4911);
and UO_678 (O_678,N_4935,N_4881);
nor UO_679 (O_679,N_4993,N_4973);
or UO_680 (O_680,N_4832,N_4983);
nor UO_681 (O_681,N_4903,N_4864);
nor UO_682 (O_682,N_4897,N_4821);
or UO_683 (O_683,N_4822,N_4946);
nand UO_684 (O_684,N_4875,N_4995);
nand UO_685 (O_685,N_4972,N_4956);
and UO_686 (O_686,N_4890,N_4863);
or UO_687 (O_687,N_4851,N_4850);
and UO_688 (O_688,N_4833,N_4931);
nor UO_689 (O_689,N_4960,N_4904);
xor UO_690 (O_690,N_4990,N_4923);
nor UO_691 (O_691,N_4914,N_4987);
nor UO_692 (O_692,N_4889,N_4910);
nand UO_693 (O_693,N_4846,N_4855);
nor UO_694 (O_694,N_4854,N_4973);
xor UO_695 (O_695,N_4802,N_4825);
and UO_696 (O_696,N_4973,N_4908);
and UO_697 (O_697,N_4883,N_4886);
xor UO_698 (O_698,N_4995,N_4984);
nor UO_699 (O_699,N_4819,N_4974);
nand UO_700 (O_700,N_4807,N_4939);
and UO_701 (O_701,N_4960,N_4876);
and UO_702 (O_702,N_4955,N_4926);
or UO_703 (O_703,N_4840,N_4915);
or UO_704 (O_704,N_4961,N_4804);
nand UO_705 (O_705,N_4919,N_4858);
nor UO_706 (O_706,N_4880,N_4997);
or UO_707 (O_707,N_4992,N_4980);
and UO_708 (O_708,N_4844,N_4867);
nor UO_709 (O_709,N_4806,N_4807);
xnor UO_710 (O_710,N_4937,N_4906);
xnor UO_711 (O_711,N_4985,N_4910);
nor UO_712 (O_712,N_4923,N_4813);
nor UO_713 (O_713,N_4935,N_4872);
nor UO_714 (O_714,N_4807,N_4901);
nor UO_715 (O_715,N_4938,N_4851);
and UO_716 (O_716,N_4808,N_4917);
and UO_717 (O_717,N_4978,N_4936);
and UO_718 (O_718,N_4957,N_4874);
nor UO_719 (O_719,N_4890,N_4880);
and UO_720 (O_720,N_4967,N_4849);
or UO_721 (O_721,N_4991,N_4846);
xnor UO_722 (O_722,N_4800,N_4935);
or UO_723 (O_723,N_4873,N_4978);
and UO_724 (O_724,N_4845,N_4869);
or UO_725 (O_725,N_4930,N_4958);
nand UO_726 (O_726,N_4997,N_4894);
nor UO_727 (O_727,N_4836,N_4973);
or UO_728 (O_728,N_4995,N_4937);
nor UO_729 (O_729,N_4951,N_4949);
and UO_730 (O_730,N_4828,N_4815);
xor UO_731 (O_731,N_4983,N_4852);
and UO_732 (O_732,N_4940,N_4901);
or UO_733 (O_733,N_4986,N_4904);
nor UO_734 (O_734,N_4916,N_4974);
nand UO_735 (O_735,N_4815,N_4955);
xor UO_736 (O_736,N_4960,N_4848);
nand UO_737 (O_737,N_4804,N_4890);
nor UO_738 (O_738,N_4839,N_4913);
and UO_739 (O_739,N_4955,N_4928);
nand UO_740 (O_740,N_4895,N_4994);
xnor UO_741 (O_741,N_4933,N_4888);
nor UO_742 (O_742,N_4915,N_4921);
nand UO_743 (O_743,N_4902,N_4952);
and UO_744 (O_744,N_4879,N_4946);
or UO_745 (O_745,N_4806,N_4819);
nand UO_746 (O_746,N_4993,N_4968);
nand UO_747 (O_747,N_4876,N_4944);
or UO_748 (O_748,N_4921,N_4896);
nand UO_749 (O_749,N_4831,N_4978);
nand UO_750 (O_750,N_4831,N_4870);
xnor UO_751 (O_751,N_4901,N_4937);
nand UO_752 (O_752,N_4951,N_4954);
nand UO_753 (O_753,N_4914,N_4879);
or UO_754 (O_754,N_4861,N_4892);
nor UO_755 (O_755,N_4939,N_4864);
or UO_756 (O_756,N_4972,N_4878);
nor UO_757 (O_757,N_4819,N_4977);
and UO_758 (O_758,N_4883,N_4881);
or UO_759 (O_759,N_4835,N_4920);
nand UO_760 (O_760,N_4852,N_4910);
nor UO_761 (O_761,N_4852,N_4947);
xor UO_762 (O_762,N_4845,N_4816);
or UO_763 (O_763,N_4921,N_4985);
nand UO_764 (O_764,N_4896,N_4850);
nor UO_765 (O_765,N_4824,N_4957);
nand UO_766 (O_766,N_4963,N_4897);
and UO_767 (O_767,N_4912,N_4864);
nor UO_768 (O_768,N_4868,N_4803);
and UO_769 (O_769,N_4848,N_4986);
or UO_770 (O_770,N_4947,N_4995);
nand UO_771 (O_771,N_4891,N_4899);
and UO_772 (O_772,N_4878,N_4952);
and UO_773 (O_773,N_4894,N_4980);
and UO_774 (O_774,N_4950,N_4859);
nand UO_775 (O_775,N_4821,N_4975);
xnor UO_776 (O_776,N_4991,N_4910);
nand UO_777 (O_777,N_4959,N_4925);
and UO_778 (O_778,N_4870,N_4892);
nor UO_779 (O_779,N_4830,N_4878);
or UO_780 (O_780,N_4920,N_4814);
and UO_781 (O_781,N_4993,N_4828);
nand UO_782 (O_782,N_4856,N_4933);
nand UO_783 (O_783,N_4894,N_4957);
nand UO_784 (O_784,N_4885,N_4854);
xnor UO_785 (O_785,N_4950,N_4831);
nand UO_786 (O_786,N_4816,N_4812);
or UO_787 (O_787,N_4822,N_4847);
xnor UO_788 (O_788,N_4866,N_4863);
xnor UO_789 (O_789,N_4980,N_4962);
nor UO_790 (O_790,N_4986,N_4984);
nand UO_791 (O_791,N_4855,N_4812);
nor UO_792 (O_792,N_4913,N_4831);
nor UO_793 (O_793,N_4947,N_4917);
and UO_794 (O_794,N_4945,N_4875);
nor UO_795 (O_795,N_4993,N_4935);
and UO_796 (O_796,N_4902,N_4939);
or UO_797 (O_797,N_4981,N_4809);
nor UO_798 (O_798,N_4843,N_4994);
or UO_799 (O_799,N_4894,N_4896);
and UO_800 (O_800,N_4838,N_4991);
nor UO_801 (O_801,N_4956,N_4819);
nand UO_802 (O_802,N_4808,N_4954);
nor UO_803 (O_803,N_4809,N_4803);
and UO_804 (O_804,N_4906,N_4829);
xnor UO_805 (O_805,N_4842,N_4850);
nand UO_806 (O_806,N_4997,N_4911);
nor UO_807 (O_807,N_4822,N_4913);
xnor UO_808 (O_808,N_4994,N_4890);
xnor UO_809 (O_809,N_4911,N_4922);
nand UO_810 (O_810,N_4849,N_4870);
or UO_811 (O_811,N_4967,N_4986);
nand UO_812 (O_812,N_4845,N_4833);
xor UO_813 (O_813,N_4925,N_4824);
and UO_814 (O_814,N_4952,N_4987);
nand UO_815 (O_815,N_4973,N_4891);
xnor UO_816 (O_816,N_4971,N_4987);
nand UO_817 (O_817,N_4858,N_4957);
nand UO_818 (O_818,N_4885,N_4829);
xor UO_819 (O_819,N_4804,N_4821);
nor UO_820 (O_820,N_4834,N_4817);
xnor UO_821 (O_821,N_4874,N_4973);
and UO_822 (O_822,N_4836,N_4848);
xnor UO_823 (O_823,N_4891,N_4961);
nand UO_824 (O_824,N_4940,N_4819);
nor UO_825 (O_825,N_4955,N_4913);
nor UO_826 (O_826,N_4832,N_4992);
or UO_827 (O_827,N_4954,N_4841);
nor UO_828 (O_828,N_4981,N_4988);
xor UO_829 (O_829,N_4933,N_4854);
nor UO_830 (O_830,N_4962,N_4984);
xnor UO_831 (O_831,N_4895,N_4926);
nor UO_832 (O_832,N_4845,N_4882);
nor UO_833 (O_833,N_4824,N_4947);
nor UO_834 (O_834,N_4806,N_4917);
nand UO_835 (O_835,N_4822,N_4902);
nand UO_836 (O_836,N_4841,N_4908);
nor UO_837 (O_837,N_4941,N_4979);
or UO_838 (O_838,N_4809,N_4864);
or UO_839 (O_839,N_4848,N_4899);
and UO_840 (O_840,N_4829,N_4922);
xor UO_841 (O_841,N_4949,N_4875);
and UO_842 (O_842,N_4915,N_4931);
xnor UO_843 (O_843,N_4930,N_4972);
nor UO_844 (O_844,N_4945,N_4809);
or UO_845 (O_845,N_4899,N_4826);
or UO_846 (O_846,N_4850,N_4815);
nor UO_847 (O_847,N_4820,N_4995);
or UO_848 (O_848,N_4931,N_4859);
nor UO_849 (O_849,N_4843,N_4963);
xnor UO_850 (O_850,N_4943,N_4977);
nand UO_851 (O_851,N_4841,N_4901);
xor UO_852 (O_852,N_4940,N_4910);
nor UO_853 (O_853,N_4816,N_4878);
nand UO_854 (O_854,N_4935,N_4835);
xor UO_855 (O_855,N_4845,N_4920);
nand UO_856 (O_856,N_4873,N_4842);
or UO_857 (O_857,N_4937,N_4931);
nand UO_858 (O_858,N_4974,N_4936);
or UO_859 (O_859,N_4847,N_4932);
nand UO_860 (O_860,N_4927,N_4991);
nand UO_861 (O_861,N_4830,N_4967);
or UO_862 (O_862,N_4927,N_4891);
and UO_863 (O_863,N_4835,N_4890);
xnor UO_864 (O_864,N_4922,N_4961);
and UO_865 (O_865,N_4858,N_4954);
nand UO_866 (O_866,N_4951,N_4909);
xor UO_867 (O_867,N_4808,N_4967);
xnor UO_868 (O_868,N_4883,N_4801);
and UO_869 (O_869,N_4937,N_4885);
and UO_870 (O_870,N_4934,N_4818);
nand UO_871 (O_871,N_4974,N_4937);
and UO_872 (O_872,N_4853,N_4917);
and UO_873 (O_873,N_4955,N_4986);
or UO_874 (O_874,N_4960,N_4922);
nand UO_875 (O_875,N_4866,N_4911);
or UO_876 (O_876,N_4924,N_4914);
and UO_877 (O_877,N_4856,N_4810);
or UO_878 (O_878,N_4967,N_4877);
and UO_879 (O_879,N_4885,N_4944);
nand UO_880 (O_880,N_4836,N_4983);
or UO_881 (O_881,N_4966,N_4943);
xor UO_882 (O_882,N_4954,N_4994);
nor UO_883 (O_883,N_4933,N_4869);
nand UO_884 (O_884,N_4849,N_4930);
and UO_885 (O_885,N_4930,N_4959);
and UO_886 (O_886,N_4979,N_4851);
nor UO_887 (O_887,N_4958,N_4875);
nand UO_888 (O_888,N_4838,N_4817);
nor UO_889 (O_889,N_4869,N_4912);
or UO_890 (O_890,N_4821,N_4971);
or UO_891 (O_891,N_4934,N_4835);
xnor UO_892 (O_892,N_4893,N_4855);
or UO_893 (O_893,N_4919,N_4897);
nand UO_894 (O_894,N_4974,N_4954);
nor UO_895 (O_895,N_4826,N_4984);
nor UO_896 (O_896,N_4837,N_4890);
nor UO_897 (O_897,N_4992,N_4906);
nand UO_898 (O_898,N_4918,N_4867);
or UO_899 (O_899,N_4816,N_4829);
or UO_900 (O_900,N_4935,N_4968);
and UO_901 (O_901,N_4950,N_4847);
nand UO_902 (O_902,N_4958,N_4898);
xnor UO_903 (O_903,N_4866,N_4842);
xor UO_904 (O_904,N_4856,N_4960);
or UO_905 (O_905,N_4919,N_4950);
or UO_906 (O_906,N_4818,N_4888);
nand UO_907 (O_907,N_4864,N_4823);
nand UO_908 (O_908,N_4935,N_4894);
nand UO_909 (O_909,N_4911,N_4810);
and UO_910 (O_910,N_4838,N_4911);
and UO_911 (O_911,N_4804,N_4991);
nand UO_912 (O_912,N_4881,N_4831);
or UO_913 (O_913,N_4838,N_4936);
and UO_914 (O_914,N_4921,N_4950);
nor UO_915 (O_915,N_4828,N_4972);
nor UO_916 (O_916,N_4894,N_4871);
nor UO_917 (O_917,N_4995,N_4933);
nand UO_918 (O_918,N_4965,N_4808);
and UO_919 (O_919,N_4916,N_4814);
nor UO_920 (O_920,N_4882,N_4990);
nor UO_921 (O_921,N_4830,N_4915);
nor UO_922 (O_922,N_4835,N_4898);
nand UO_923 (O_923,N_4994,N_4869);
nand UO_924 (O_924,N_4974,N_4807);
nor UO_925 (O_925,N_4947,N_4849);
nand UO_926 (O_926,N_4978,N_4975);
nor UO_927 (O_927,N_4987,N_4849);
or UO_928 (O_928,N_4832,N_4957);
and UO_929 (O_929,N_4939,N_4980);
and UO_930 (O_930,N_4835,N_4811);
nor UO_931 (O_931,N_4806,N_4823);
and UO_932 (O_932,N_4897,N_4842);
xnor UO_933 (O_933,N_4857,N_4982);
xor UO_934 (O_934,N_4866,N_4908);
and UO_935 (O_935,N_4962,N_4961);
or UO_936 (O_936,N_4852,N_4902);
or UO_937 (O_937,N_4862,N_4937);
and UO_938 (O_938,N_4828,N_4821);
nand UO_939 (O_939,N_4910,N_4857);
or UO_940 (O_940,N_4836,N_4959);
or UO_941 (O_941,N_4898,N_4838);
nand UO_942 (O_942,N_4854,N_4887);
and UO_943 (O_943,N_4825,N_4848);
nor UO_944 (O_944,N_4870,N_4887);
and UO_945 (O_945,N_4984,N_4941);
or UO_946 (O_946,N_4876,N_4941);
nand UO_947 (O_947,N_4848,N_4914);
xor UO_948 (O_948,N_4884,N_4822);
and UO_949 (O_949,N_4872,N_4813);
nand UO_950 (O_950,N_4836,N_4890);
and UO_951 (O_951,N_4965,N_4859);
and UO_952 (O_952,N_4995,N_4830);
nor UO_953 (O_953,N_4984,N_4963);
and UO_954 (O_954,N_4947,N_4952);
nor UO_955 (O_955,N_4975,N_4918);
nand UO_956 (O_956,N_4978,N_4843);
nor UO_957 (O_957,N_4887,N_4993);
nor UO_958 (O_958,N_4956,N_4996);
nor UO_959 (O_959,N_4861,N_4908);
nor UO_960 (O_960,N_4944,N_4989);
and UO_961 (O_961,N_4974,N_4903);
and UO_962 (O_962,N_4938,N_4869);
or UO_963 (O_963,N_4933,N_4918);
or UO_964 (O_964,N_4851,N_4852);
xnor UO_965 (O_965,N_4916,N_4857);
or UO_966 (O_966,N_4984,N_4974);
nand UO_967 (O_967,N_4916,N_4981);
nand UO_968 (O_968,N_4871,N_4813);
nand UO_969 (O_969,N_4889,N_4942);
nor UO_970 (O_970,N_4933,N_4805);
and UO_971 (O_971,N_4992,N_4903);
nand UO_972 (O_972,N_4970,N_4928);
and UO_973 (O_973,N_4959,N_4982);
and UO_974 (O_974,N_4920,N_4933);
and UO_975 (O_975,N_4963,N_4930);
and UO_976 (O_976,N_4885,N_4862);
or UO_977 (O_977,N_4915,N_4980);
or UO_978 (O_978,N_4875,N_4897);
xnor UO_979 (O_979,N_4801,N_4845);
nand UO_980 (O_980,N_4999,N_4929);
nor UO_981 (O_981,N_4828,N_4807);
nor UO_982 (O_982,N_4942,N_4897);
xnor UO_983 (O_983,N_4808,N_4856);
or UO_984 (O_984,N_4812,N_4938);
or UO_985 (O_985,N_4842,N_4852);
nor UO_986 (O_986,N_4882,N_4862);
nor UO_987 (O_987,N_4976,N_4830);
nand UO_988 (O_988,N_4927,N_4978);
or UO_989 (O_989,N_4920,N_4841);
xnor UO_990 (O_990,N_4856,N_4968);
or UO_991 (O_991,N_4831,N_4963);
and UO_992 (O_992,N_4924,N_4859);
or UO_993 (O_993,N_4991,N_4869);
xor UO_994 (O_994,N_4952,N_4824);
xor UO_995 (O_995,N_4869,N_4850);
or UO_996 (O_996,N_4950,N_4961);
and UO_997 (O_997,N_4998,N_4885);
nor UO_998 (O_998,N_4896,N_4826);
nand UO_999 (O_999,N_4905,N_4962);
endmodule