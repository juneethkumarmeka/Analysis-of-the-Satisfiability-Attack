module basic_750_5000_1000_2_levels_1xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2502,N_2503,N_2505,N_2506,N_2507,N_2509,N_2511,N_2512,N_2513,N_2516,N_2517,N_2518,N_2519,N_2520,N_2522,N_2523,N_2524,N_2525,N_2526,N_2529,N_2531,N_2535,N_2536,N_2537,N_2538,N_2540,N_2541,N_2543,N_2546,N_2547,N_2548,N_2550,N_2551,N_2552,N_2553,N_2556,N_2557,N_2558,N_2559,N_2560,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2589,N_2591,N_2594,N_2595,N_2596,N_2598,N_2599,N_2600,N_2601,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2615,N_2617,N_2618,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2630,N_2631,N_2633,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2642,N_2644,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2655,N_2656,N_2657,N_2660,N_2661,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2678,N_2679,N_2680,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2696,N_2698,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2707,N_2708,N_2709,N_2710,N_2714,N_2715,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2736,N_2737,N_2738,N_2740,N_2741,N_2743,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2815,N_2816,N_2818,N_2819,N_2821,N_2823,N_2824,N_2825,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2837,N_2839,N_2840,N_2841,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2858,N_2859,N_2860,N_2861,N_2863,N_2866,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2881,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2896,N_2897,N_2898,N_2900,N_2901,N_2902,N_2903,N_2905,N_2907,N_2908,N_2909,N_2910,N_2912,N_2913,N_2914,N_2916,N_2917,N_2918,N_2920,N_2921,N_2924,N_2925,N_2926,N_2928,N_2929,N_2933,N_2934,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2948,N_2949,N_2951,N_2952,N_2954,N_2955,N_2956,N_2957,N_2960,N_2961,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2988,N_2990,N_2991,N_2992,N_2996,N_2997,N_2998,N_3001,N_3002,N_3004,N_3005,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3021,N_3022,N_3023,N_3024,N_3025,N_3028,N_3029,N_3030,N_3031,N_3032,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3049,N_3051,N_3052,N_3053,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3064,N_3065,N_3066,N_3068,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3081,N_3083,N_3084,N_3085,N_3086,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3100,N_3101,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3136,N_3137,N_3138,N_3139,N_3141,N_3142,N_3144,N_3145,N_3146,N_3147,N_3148,N_3151,N_3152,N_3155,N_3157,N_3158,N_3159,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3169,N_3170,N_3171,N_3172,N_3173,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3183,N_3184,N_3185,N_3187,N_3188,N_3190,N_3191,N_3192,N_3193,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3235,N_3236,N_3238,N_3239,N_3240,N_3241,N_3243,N_3244,N_3245,N_3248,N_3249,N_3250,N_3252,N_3253,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3275,N_3276,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3306,N_3307,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3317,N_3318,N_3320,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3335,N_3336,N_3337,N_3338,N_3339,N_3341,N_3342,N_3343,N_3346,N_3347,N_3350,N_3352,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3370,N_3371,N_3372,N_3373,N_3375,N_3376,N_3377,N_3378,N_3379,N_3381,N_3382,N_3383,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3396,N_3397,N_3398,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3410,N_3411,N_3412,N_3413,N_3414,N_3416,N_3417,N_3419,N_3420,N_3422,N_3423,N_3424,N_3426,N_3427,N_3430,N_3432,N_3433,N_3434,N_3435,N_3437,N_3438,N_3439,N_3440,N_3441,N_3443,N_3445,N_3446,N_3448,N_3451,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3490,N_3492,N_3495,N_3496,N_3497,N_3498,N_3499,N_3502,N_3503,N_3504,N_3505,N_3506,N_3508,N_3509,N_3510,N_3511,N_3512,N_3514,N_3515,N_3518,N_3519,N_3520,N_3521,N_3522,N_3524,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3540,N_3541,N_3542,N_3544,N_3546,N_3547,N_3548,N_3549,N_3550,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3561,N_3562,N_3563,N_3566,N_3567,N_3568,N_3569,N_3571,N_3572,N_3573,N_3575,N_3576,N_3577,N_3578,N_3579,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3597,N_3598,N_3599,N_3600,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3615,N_3616,N_3619,N_3620,N_3621,N_3622,N_3623,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3632,N_3633,N_3634,N_3637,N_3638,N_3639,N_3640,N_3641,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3655,N_3656,N_3657,N_3659,N_3660,N_3661,N_3664,N_3665,N_3666,N_3668,N_3671,N_3672,N_3673,N_3676,N_3677,N_3678,N_3681,N_3682,N_3683,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3694,N_3695,N_3696,N_3697,N_3700,N_3701,N_3702,N_3703,N_3704,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3727,N_3728,N_3729,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3749,N_3751,N_3753,N_3756,N_3757,N_3758,N_3759,N_3760,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3775,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3786,N_3787,N_3788,N_3789,N_3791,N_3794,N_3795,N_3796,N_3798,N_3799,N_3800,N_3802,N_3803,N_3805,N_3806,N_3807,N_3809,N_3810,N_3811,N_3812,N_3813,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3857,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3871,N_3874,N_3875,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3898,N_3899,N_3900,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3926,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3935,N_3936,N_3937,N_3939,N_3940,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3967,N_3968,N_3969,N_3970,N_3972,N_3973,N_3974,N_3975,N_3977,N_3978,N_3980,N_3981,N_3982,N_3983,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3996,N_3997,N_3998,N_4000,N_4001,N_4002,N_4003,N_4005,N_4006,N_4008,N_4010,N_4011,N_4012,N_4013,N_4014,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4036,N_4037,N_4039,N_4041,N_4042,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4085,N_4086,N_4089,N_4092,N_4093,N_4095,N_4096,N_4097,N_4098,N_4100,N_4101,N_4102,N_4103,N_4104,N_4106,N_4107,N_4108,N_4109,N_4111,N_4112,N_4115,N_4116,N_4118,N_4119,N_4120,N_4121,N_4123,N_4124,N_4126,N_4127,N_4129,N_4131,N_4132,N_4133,N_4134,N_4135,N_4137,N_4138,N_4140,N_4141,N_4142,N_4143,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4152,N_4153,N_4154,N_4155,N_4156,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4187,N_4188,N_4191,N_4192,N_4193,N_4196,N_4197,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4252,N_4253,N_4254,N_4256,N_4258,N_4259,N_4261,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4285,N_4286,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4310,N_4311,N_4313,N_4314,N_4316,N_4317,N_4319,N_4320,N_4321,N_4322,N_4323,N_4328,N_4329,N_4331,N_4334,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4346,N_4347,N_4348,N_4349,N_4350,N_4352,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4385,N_4387,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4401,N_4402,N_4403,N_4404,N_4406,N_4407,N_4408,N_4409,N_4410,N_4412,N_4413,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4452,N_4454,N_4455,N_4456,N_4457,N_4458,N_4460,N_4461,N_4462,N_4463,N_4464,N_4466,N_4467,N_4468,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4481,N_4482,N_4483,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4494,N_4495,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4509,N_4510,N_4511,N_4513,N_4514,N_4515,N_4517,N_4518,N_4519,N_4520,N_4521,N_4523,N_4524,N_4525,N_4526,N_4527,N_4529,N_4530,N_4531,N_4533,N_4535,N_4537,N_4538,N_4540,N_4541,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4586,N_4587,N_4589,N_4590,N_4592,N_4593,N_4594,N_4595,N_4597,N_4598,N_4599,N_4600,N_4601,N_4603,N_4604,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4613,N_4614,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4634,N_4635,N_4636,N_4637,N_4638,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4653,N_4654,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4664,N_4665,N_4666,N_4667,N_4668,N_4670,N_4672,N_4673,N_4674,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4684,N_4685,N_4686,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4696,N_4697,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4721,N_4725,N_4726,N_4727,N_4728,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4763,N_4764,N_4766,N_4768,N_4769,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4815,N_4818,N_4819,N_4820,N_4822,N_4823,N_4825,N_4826,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4851,N_4852,N_4853,N_4854,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4870,N_4872,N_4873,N_4874,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4884,N_4885,N_4886,N_4887,N_4888,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4919,N_4923,N_4924,N_4926,N_4927,N_4928,N_4929,N_4931,N_4933,N_4934,N_4935,N_4937,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4954,N_4955,N_4956,N_4957,N_4958,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4979,N_4980,N_4981,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4998,N_4999;
nand U0 (N_0,In_724,In_485);
or U1 (N_1,In_443,In_481);
nand U2 (N_2,In_260,In_422);
nor U3 (N_3,In_43,In_339);
or U4 (N_4,In_577,In_384);
xnor U5 (N_5,In_52,In_711);
xnor U6 (N_6,In_446,In_746);
or U7 (N_7,In_202,In_328);
or U8 (N_8,In_487,In_373);
or U9 (N_9,In_381,In_92);
nand U10 (N_10,In_343,In_108);
nor U11 (N_11,In_147,In_473);
nand U12 (N_12,In_149,In_709);
nand U13 (N_13,In_488,In_122);
nand U14 (N_14,In_214,In_447);
or U15 (N_15,In_527,In_565);
and U16 (N_16,In_583,In_142);
nor U17 (N_17,In_164,In_67);
nand U18 (N_18,In_242,In_702);
nand U19 (N_19,In_528,In_564);
nand U20 (N_20,In_170,In_361);
nor U21 (N_21,In_17,In_167);
and U22 (N_22,In_448,In_492);
or U23 (N_23,In_595,In_687);
and U24 (N_24,In_203,In_249);
and U25 (N_25,In_582,In_347);
nand U26 (N_26,In_228,In_679);
or U27 (N_27,In_686,In_695);
xor U28 (N_28,In_340,In_174);
nand U29 (N_29,In_417,In_216);
nand U30 (N_30,In_737,In_662);
nor U31 (N_31,In_162,In_289);
nor U32 (N_32,In_639,In_199);
nor U33 (N_33,In_478,In_219);
or U34 (N_34,In_175,In_580);
and U35 (N_35,In_325,In_459);
nand U36 (N_36,In_96,In_543);
nand U37 (N_37,In_456,In_375);
nand U38 (N_38,In_4,In_101);
nor U39 (N_39,In_525,In_649);
nand U40 (N_40,In_41,In_93);
nand U41 (N_41,In_424,In_633);
and U42 (N_42,In_69,In_745);
or U43 (N_43,In_3,In_313);
and U44 (N_44,In_460,In_573);
nor U45 (N_45,In_246,In_55);
and U46 (N_46,In_638,In_689);
and U47 (N_47,In_708,In_282);
or U48 (N_48,In_269,In_120);
or U49 (N_49,In_342,In_676);
nor U50 (N_50,In_320,In_585);
nand U51 (N_51,In_698,In_561);
and U52 (N_52,In_178,In_66);
and U53 (N_53,In_379,In_226);
or U54 (N_54,In_465,In_501);
nand U55 (N_55,In_368,In_206);
nor U56 (N_56,In_427,In_376);
or U57 (N_57,In_499,In_441);
nand U58 (N_58,In_137,In_363);
and U59 (N_59,In_374,In_391);
or U60 (N_60,In_444,In_7);
nand U61 (N_61,In_400,In_539);
and U62 (N_62,In_90,In_97);
nand U63 (N_63,In_620,In_629);
and U64 (N_64,In_79,In_429);
and U65 (N_65,In_238,In_114);
or U66 (N_66,In_284,In_571);
or U67 (N_67,In_33,In_513);
nand U68 (N_68,In_84,In_109);
and U69 (N_69,In_378,In_404);
nor U70 (N_70,In_128,In_472);
or U71 (N_71,In_263,In_256);
and U72 (N_72,In_100,In_198);
nor U73 (N_73,In_644,In_551);
nor U74 (N_74,In_11,In_266);
and U75 (N_75,In_642,In_102);
nand U76 (N_76,In_454,In_602);
nor U77 (N_77,In_704,In_14);
or U78 (N_78,In_161,In_721);
nor U79 (N_79,In_218,In_222);
and U80 (N_80,In_537,In_184);
nor U81 (N_81,In_48,In_104);
or U82 (N_82,In_13,In_461);
or U83 (N_83,In_299,In_645);
nor U84 (N_84,In_450,In_383);
or U85 (N_85,In_237,In_418);
nor U86 (N_86,In_277,In_389);
or U87 (N_87,In_179,In_117);
nor U88 (N_88,In_557,In_394);
nor U89 (N_89,In_707,In_171);
and U90 (N_90,In_195,In_747);
or U91 (N_91,In_603,In_318);
and U92 (N_92,In_526,In_736);
and U93 (N_93,In_636,In_165);
nor U94 (N_94,In_24,In_223);
and U95 (N_95,In_37,In_32);
nor U96 (N_96,In_62,In_123);
nand U97 (N_97,In_519,In_230);
or U98 (N_98,In_684,In_29);
or U99 (N_99,In_156,In_319);
nor U100 (N_100,In_35,In_221);
nor U101 (N_101,In_601,In_477);
nor U102 (N_102,In_305,In_432);
nand U103 (N_103,In_30,In_64);
xnor U104 (N_104,In_598,In_484);
and U105 (N_105,In_209,In_316);
and U106 (N_106,In_452,In_262);
and U107 (N_107,In_393,In_713);
and U108 (N_108,In_245,In_421);
nor U109 (N_109,In_306,In_553);
and U110 (N_110,In_236,In_111);
nand U111 (N_111,In_185,In_89);
and U112 (N_112,In_99,In_307);
or U113 (N_113,In_480,In_207);
nor U114 (N_114,In_106,In_302);
nor U115 (N_115,In_398,In_303);
nor U116 (N_116,In_545,In_118);
or U117 (N_117,In_57,In_124);
nor U118 (N_118,In_58,In_344);
nand U119 (N_119,In_594,In_357);
and U120 (N_120,In_744,In_574);
or U121 (N_121,In_630,In_466);
nand U122 (N_122,In_436,In_570);
nand U123 (N_123,In_129,In_157);
nor U124 (N_124,In_433,In_483);
nor U125 (N_125,In_496,In_234);
or U126 (N_126,In_494,In_740);
and U127 (N_127,In_74,In_235);
nand U128 (N_128,In_489,In_412);
or U129 (N_129,In_188,In_233);
or U130 (N_130,In_270,In_294);
or U131 (N_131,In_608,In_469);
or U132 (N_132,In_81,In_591);
nor U133 (N_133,In_596,In_135);
or U134 (N_134,In_220,In_26);
or U135 (N_135,In_152,In_140);
xnor U136 (N_136,In_741,In_685);
or U137 (N_137,In_535,In_42);
and U138 (N_138,In_680,In_546);
or U139 (N_139,In_449,In_304);
and U140 (N_140,In_619,In_227);
nand U141 (N_141,In_738,In_430);
and U142 (N_142,In_244,In_669);
and U143 (N_143,In_309,In_654);
nand U144 (N_144,In_335,In_560);
nor U145 (N_145,In_20,In_604);
nor U146 (N_146,In_634,In_159);
nand U147 (N_147,In_498,In_27);
or U148 (N_148,In_336,In_440);
or U149 (N_149,In_650,In_590);
and U150 (N_150,In_193,In_211);
or U151 (N_151,In_366,In_315);
nor U152 (N_152,In_556,In_434);
or U153 (N_153,In_180,In_49);
nor U154 (N_154,In_416,In_212);
nand U155 (N_155,In_563,In_613);
and U156 (N_156,In_39,In_621);
or U157 (N_157,In_252,In_382);
nand U158 (N_158,In_46,In_665);
and U159 (N_159,In_80,In_190);
and U160 (N_160,In_646,In_321);
nor U161 (N_161,In_139,In_349);
nand U162 (N_162,In_224,In_54);
or U163 (N_163,In_355,In_438);
or U164 (N_164,In_281,In_749);
nand U165 (N_165,In_581,In_257);
nor U166 (N_166,In_200,In_362);
or U167 (N_167,In_622,In_247);
nor U168 (N_168,In_463,In_2);
or U169 (N_169,In_1,In_377);
and U170 (N_170,In_194,In_504);
and U171 (N_171,In_173,In_575);
nand U172 (N_172,In_356,In_176);
and U173 (N_173,In_158,In_548);
and U174 (N_174,In_442,In_593);
nor U175 (N_175,In_628,In_627);
or U176 (N_176,In_510,In_144);
or U177 (N_177,In_599,In_172);
nand U178 (N_178,In_61,In_82);
and U179 (N_179,In_134,In_291);
nor U180 (N_180,In_21,In_19);
xor U181 (N_181,In_166,In_664);
or U182 (N_182,In_559,In_395);
or U183 (N_183,In_215,In_431);
nor U184 (N_184,In_544,In_464);
and U185 (N_185,In_267,In_533);
nand U186 (N_186,In_723,In_632);
nor U187 (N_187,In_85,In_722);
or U188 (N_188,In_506,In_660);
xnor U189 (N_189,In_251,In_15);
and U190 (N_190,In_276,In_720);
nand U191 (N_191,In_338,In_516);
or U192 (N_192,In_503,In_133);
and U193 (N_193,In_201,In_453);
nor U194 (N_194,In_353,In_110);
or U195 (N_195,In_12,In_229);
or U196 (N_196,In_413,In_618);
or U197 (N_197,In_491,In_288);
or U198 (N_198,In_439,In_673);
nor U199 (N_199,In_587,In_568);
and U200 (N_200,In_131,In_177);
nor U201 (N_201,In_332,In_208);
nand U202 (N_202,In_196,In_584);
nand U203 (N_203,In_94,In_411);
nand U204 (N_204,In_502,In_712);
and U205 (N_205,In_701,In_44);
or U206 (N_206,In_264,In_72);
and U207 (N_207,In_652,In_314);
nor U208 (N_208,In_697,In_532);
nor U209 (N_209,In_141,In_95);
nor U210 (N_210,In_399,In_76);
nor U211 (N_211,In_530,In_125);
and U212 (N_212,In_243,In_495);
and U213 (N_213,In_426,In_225);
nand U214 (N_214,In_607,In_189);
nor U215 (N_215,In_107,In_589);
nor U216 (N_216,In_358,In_259);
and U217 (N_217,In_547,In_365);
and U218 (N_218,In_31,In_617);
nand U219 (N_219,In_369,In_88);
nand U220 (N_220,In_254,In_323);
nor U221 (N_221,In_540,In_408);
or U222 (N_222,In_730,In_523);
and U223 (N_223,In_324,In_348);
nand U224 (N_224,In_455,In_715);
xor U225 (N_225,In_51,In_345);
and U226 (N_226,In_396,In_612);
and U227 (N_227,In_169,In_40);
nor U228 (N_228,In_239,In_690);
or U229 (N_229,In_658,In_286);
and U230 (N_230,In_732,In_675);
and U231 (N_231,In_457,In_354);
nand U232 (N_232,In_522,In_609);
or U233 (N_233,In_677,In_409);
nand U234 (N_234,In_210,In_248);
and U235 (N_235,In_670,In_529);
nand U236 (N_236,In_330,In_705);
or U237 (N_237,In_719,In_626);
and U238 (N_238,In_470,In_588);
nor U239 (N_239,In_8,In_734);
nor U240 (N_240,In_91,In_663);
nor U241 (N_241,In_554,In_6);
or U242 (N_242,In_297,In_386);
nand U243 (N_243,In_428,In_60);
nor U244 (N_244,In_682,In_521);
and U245 (N_245,In_371,In_518);
nor U246 (N_246,In_367,In_146);
nand U247 (N_247,In_597,In_572);
xor U248 (N_248,In_205,In_414);
and U249 (N_249,In_163,In_531);
and U250 (N_250,In_435,In_611);
nor U251 (N_251,In_605,In_292);
or U252 (N_252,In_168,In_425);
and U253 (N_253,In_105,In_370);
nor U254 (N_254,In_160,In_748);
nor U255 (N_255,In_191,In_462);
and U256 (N_256,In_641,In_718);
or U257 (N_257,In_566,In_45);
nand U258 (N_258,In_616,In_648);
and U259 (N_259,In_327,In_23);
nor U260 (N_260,In_87,In_71);
and U261 (N_261,In_115,In_419);
or U262 (N_262,In_253,In_275);
nand U263 (N_263,In_651,In_28);
or U264 (N_264,In_655,In_541);
xnor U265 (N_265,In_490,In_717);
nand U266 (N_266,In_56,In_407);
nand U267 (N_267,In_5,In_538);
nand U268 (N_268,In_726,In_667);
or U269 (N_269,In_562,In_63);
nand U270 (N_270,In_467,In_241);
or U271 (N_271,In_273,In_143);
nor U272 (N_272,In_126,In_186);
nand U273 (N_273,In_520,In_271);
or U274 (N_274,In_372,In_265);
or U275 (N_275,In_390,In_555);
nor U276 (N_276,In_279,In_731);
and U277 (N_277,In_113,In_380);
or U278 (N_278,In_512,In_733);
nor U279 (N_279,In_507,In_192);
nor U280 (N_280,In_727,In_352);
nor U281 (N_281,In_696,In_514);
or U282 (N_282,In_714,In_668);
nand U283 (N_283,In_637,In_34);
or U284 (N_284,In_231,In_666);
or U285 (N_285,In_148,In_59);
nor U286 (N_286,In_197,In_661);
nand U287 (N_287,In_569,In_479);
nor U288 (N_288,In_742,In_25);
nor U289 (N_289,In_301,In_387);
nand U290 (N_290,In_683,In_402);
nor U291 (N_291,In_255,In_657);
nor U292 (N_292,In_656,In_83);
nand U293 (N_293,In_258,In_274);
nor U294 (N_294,In_0,In_360);
nand U295 (N_295,In_287,In_36);
and U296 (N_296,In_672,In_542);
nand U297 (N_297,In_153,In_415);
or U298 (N_298,In_725,In_341);
and U299 (N_299,In_739,In_614);
nor U300 (N_300,In_640,In_293);
or U301 (N_301,In_272,In_127);
nor U302 (N_302,In_280,In_471);
nor U303 (N_303,In_451,In_688);
nor U304 (N_304,In_331,In_624);
nand U305 (N_305,In_486,In_476);
or U306 (N_306,In_145,In_217);
nand U307 (N_307,In_116,In_567);
or U308 (N_308,In_295,In_623);
or U309 (N_309,In_317,In_392);
or U310 (N_310,In_610,In_524);
nand U311 (N_311,In_308,In_75);
or U312 (N_312,In_182,In_388);
nor U313 (N_313,In_334,In_710);
or U314 (N_314,In_549,In_16);
nand U315 (N_315,In_47,In_631);
or U316 (N_316,In_50,In_653);
nor U317 (N_317,In_300,In_517);
nor U318 (N_318,In_703,In_497);
nor U319 (N_319,In_385,In_311);
nor U320 (N_320,In_121,In_509);
or U321 (N_321,In_68,In_674);
nor U322 (N_322,In_671,In_728);
nand U323 (N_323,In_86,In_154);
nor U324 (N_324,In_10,In_458);
and U325 (N_325,In_296,In_445);
or U326 (N_326,In_183,In_22);
and U327 (N_327,In_474,In_681);
nor U328 (N_328,In_691,In_558);
nand U329 (N_329,In_678,In_729);
nor U330 (N_330,In_552,In_606);
and U331 (N_331,In_65,In_735);
or U332 (N_332,In_18,In_716);
nand U333 (N_333,In_550,In_643);
nor U334 (N_334,In_53,In_420);
or U335 (N_335,In_73,In_322);
or U336 (N_336,In_592,In_600);
and U337 (N_337,In_515,In_78);
nor U338 (N_338,In_181,In_406);
or U339 (N_339,In_694,In_351);
and U340 (N_340,In_150,In_500);
nand U341 (N_341,In_337,In_706);
and U342 (N_342,In_403,In_615);
and U343 (N_343,In_576,In_505);
and U344 (N_344,In_232,In_437);
nor U345 (N_345,In_77,In_397);
and U346 (N_346,In_285,In_468);
or U347 (N_347,In_423,In_700);
and U348 (N_348,In_482,In_635);
nand U349 (N_349,In_493,In_298);
or U350 (N_350,In_659,In_250);
or U351 (N_351,In_405,In_743);
and U352 (N_352,In_346,In_692);
nand U353 (N_353,In_70,In_103);
and U354 (N_354,In_699,In_359);
or U355 (N_355,In_579,In_625);
nor U356 (N_356,In_310,In_112);
and U357 (N_357,In_213,In_401);
nor U358 (N_358,In_155,In_261);
and U359 (N_359,In_278,In_586);
and U360 (N_360,In_98,In_536);
and U361 (N_361,In_511,In_534);
or U362 (N_362,In_132,In_333);
and U363 (N_363,In_290,In_268);
nor U364 (N_364,In_364,In_508);
nor U365 (N_365,In_647,In_283);
or U366 (N_366,In_350,In_136);
nand U367 (N_367,In_329,In_475);
or U368 (N_368,In_312,In_187);
or U369 (N_369,In_9,In_693);
or U370 (N_370,In_204,In_119);
nand U371 (N_371,In_130,In_410);
and U372 (N_372,In_326,In_151);
nor U373 (N_373,In_38,In_578);
and U374 (N_374,In_240,In_138);
nand U375 (N_375,In_433,In_153);
nand U376 (N_376,In_426,In_58);
or U377 (N_377,In_11,In_243);
nand U378 (N_378,In_713,In_29);
and U379 (N_379,In_354,In_486);
nand U380 (N_380,In_410,In_450);
nand U381 (N_381,In_414,In_430);
nor U382 (N_382,In_433,In_210);
nand U383 (N_383,In_620,In_383);
or U384 (N_384,In_34,In_629);
or U385 (N_385,In_142,In_446);
nor U386 (N_386,In_104,In_228);
nor U387 (N_387,In_272,In_361);
nor U388 (N_388,In_71,In_379);
nand U389 (N_389,In_603,In_193);
and U390 (N_390,In_583,In_743);
and U391 (N_391,In_507,In_365);
or U392 (N_392,In_62,In_627);
and U393 (N_393,In_560,In_2);
or U394 (N_394,In_316,In_613);
and U395 (N_395,In_569,In_354);
nand U396 (N_396,In_6,In_513);
and U397 (N_397,In_139,In_268);
or U398 (N_398,In_458,In_436);
or U399 (N_399,In_127,In_123);
or U400 (N_400,In_497,In_455);
or U401 (N_401,In_402,In_139);
or U402 (N_402,In_621,In_128);
nand U403 (N_403,In_412,In_384);
and U404 (N_404,In_53,In_689);
and U405 (N_405,In_407,In_68);
and U406 (N_406,In_508,In_352);
or U407 (N_407,In_542,In_10);
or U408 (N_408,In_577,In_606);
and U409 (N_409,In_356,In_475);
and U410 (N_410,In_165,In_211);
or U411 (N_411,In_379,In_271);
or U412 (N_412,In_680,In_686);
nand U413 (N_413,In_686,In_609);
nand U414 (N_414,In_403,In_43);
nand U415 (N_415,In_381,In_595);
nand U416 (N_416,In_121,In_212);
nand U417 (N_417,In_211,In_728);
nor U418 (N_418,In_144,In_336);
or U419 (N_419,In_383,In_362);
nor U420 (N_420,In_542,In_643);
nor U421 (N_421,In_690,In_158);
nand U422 (N_422,In_508,In_383);
nand U423 (N_423,In_562,In_688);
or U424 (N_424,In_442,In_681);
nor U425 (N_425,In_209,In_372);
nor U426 (N_426,In_331,In_223);
or U427 (N_427,In_168,In_539);
and U428 (N_428,In_140,In_476);
nand U429 (N_429,In_637,In_196);
nor U430 (N_430,In_585,In_229);
or U431 (N_431,In_488,In_251);
nand U432 (N_432,In_82,In_103);
nand U433 (N_433,In_573,In_627);
nand U434 (N_434,In_325,In_403);
and U435 (N_435,In_303,In_482);
or U436 (N_436,In_59,In_318);
nor U437 (N_437,In_714,In_707);
or U438 (N_438,In_481,In_523);
nor U439 (N_439,In_660,In_103);
nor U440 (N_440,In_363,In_737);
and U441 (N_441,In_228,In_388);
nor U442 (N_442,In_115,In_647);
or U443 (N_443,In_487,In_200);
nand U444 (N_444,In_508,In_280);
or U445 (N_445,In_441,In_354);
and U446 (N_446,In_590,In_417);
nor U447 (N_447,In_185,In_327);
nand U448 (N_448,In_595,In_418);
nand U449 (N_449,In_606,In_49);
nor U450 (N_450,In_364,In_116);
nand U451 (N_451,In_563,In_147);
nor U452 (N_452,In_190,In_744);
nand U453 (N_453,In_38,In_413);
nand U454 (N_454,In_413,In_659);
nor U455 (N_455,In_592,In_14);
and U456 (N_456,In_442,In_330);
nor U457 (N_457,In_478,In_378);
or U458 (N_458,In_557,In_188);
nor U459 (N_459,In_66,In_639);
nor U460 (N_460,In_728,In_503);
nor U461 (N_461,In_696,In_660);
and U462 (N_462,In_425,In_155);
nor U463 (N_463,In_216,In_79);
or U464 (N_464,In_565,In_558);
nand U465 (N_465,In_376,In_277);
or U466 (N_466,In_536,In_595);
and U467 (N_467,In_712,In_677);
nor U468 (N_468,In_125,In_340);
xnor U469 (N_469,In_586,In_19);
or U470 (N_470,In_114,In_715);
or U471 (N_471,In_393,In_360);
or U472 (N_472,In_260,In_609);
and U473 (N_473,In_613,In_596);
nor U474 (N_474,In_521,In_35);
and U475 (N_475,In_466,In_18);
and U476 (N_476,In_236,In_633);
nand U477 (N_477,In_723,In_213);
nor U478 (N_478,In_698,In_559);
nand U479 (N_479,In_329,In_609);
nand U480 (N_480,In_163,In_196);
and U481 (N_481,In_680,In_685);
nor U482 (N_482,In_83,In_406);
nor U483 (N_483,In_43,In_666);
nor U484 (N_484,In_711,In_523);
nand U485 (N_485,In_141,In_661);
or U486 (N_486,In_520,In_29);
nand U487 (N_487,In_317,In_417);
nand U488 (N_488,In_454,In_255);
and U489 (N_489,In_272,In_203);
or U490 (N_490,In_580,In_59);
nand U491 (N_491,In_17,In_104);
nand U492 (N_492,In_186,In_98);
nand U493 (N_493,In_537,In_465);
and U494 (N_494,In_669,In_300);
nand U495 (N_495,In_678,In_64);
or U496 (N_496,In_713,In_539);
or U497 (N_497,In_612,In_271);
nor U498 (N_498,In_580,In_275);
nor U499 (N_499,In_354,In_127);
and U500 (N_500,In_89,In_152);
xor U501 (N_501,In_476,In_0);
and U502 (N_502,In_375,In_618);
xnor U503 (N_503,In_75,In_561);
or U504 (N_504,In_289,In_33);
nor U505 (N_505,In_666,In_494);
nand U506 (N_506,In_301,In_614);
nand U507 (N_507,In_412,In_564);
nor U508 (N_508,In_247,In_49);
or U509 (N_509,In_230,In_547);
nand U510 (N_510,In_311,In_394);
nand U511 (N_511,In_646,In_19);
nor U512 (N_512,In_510,In_373);
nand U513 (N_513,In_728,In_160);
and U514 (N_514,In_141,In_36);
nand U515 (N_515,In_579,In_201);
nand U516 (N_516,In_705,In_479);
nand U517 (N_517,In_130,In_303);
nand U518 (N_518,In_34,In_291);
nor U519 (N_519,In_468,In_683);
nor U520 (N_520,In_646,In_204);
nand U521 (N_521,In_189,In_194);
or U522 (N_522,In_52,In_93);
and U523 (N_523,In_706,In_147);
or U524 (N_524,In_683,In_655);
or U525 (N_525,In_576,In_654);
and U526 (N_526,In_230,In_379);
nor U527 (N_527,In_207,In_313);
nand U528 (N_528,In_669,In_407);
or U529 (N_529,In_208,In_79);
and U530 (N_530,In_647,In_13);
or U531 (N_531,In_672,In_524);
nand U532 (N_532,In_716,In_197);
or U533 (N_533,In_417,In_329);
and U534 (N_534,In_71,In_441);
and U535 (N_535,In_464,In_400);
nor U536 (N_536,In_507,In_171);
or U537 (N_537,In_255,In_167);
and U538 (N_538,In_559,In_63);
nand U539 (N_539,In_469,In_435);
nor U540 (N_540,In_77,In_685);
nor U541 (N_541,In_132,In_562);
nand U542 (N_542,In_141,In_720);
nand U543 (N_543,In_141,In_38);
or U544 (N_544,In_440,In_30);
and U545 (N_545,In_82,In_381);
nand U546 (N_546,In_591,In_455);
or U547 (N_547,In_334,In_7);
or U548 (N_548,In_498,In_532);
nand U549 (N_549,In_487,In_558);
nand U550 (N_550,In_267,In_573);
nand U551 (N_551,In_709,In_396);
and U552 (N_552,In_8,In_724);
nand U553 (N_553,In_603,In_343);
nor U554 (N_554,In_194,In_76);
or U555 (N_555,In_228,In_155);
nor U556 (N_556,In_517,In_141);
and U557 (N_557,In_161,In_302);
and U558 (N_558,In_529,In_512);
or U559 (N_559,In_540,In_2);
nor U560 (N_560,In_477,In_429);
or U561 (N_561,In_331,In_158);
nand U562 (N_562,In_377,In_424);
or U563 (N_563,In_237,In_105);
and U564 (N_564,In_287,In_148);
nor U565 (N_565,In_414,In_561);
nor U566 (N_566,In_102,In_137);
nand U567 (N_567,In_155,In_34);
xnor U568 (N_568,In_664,In_562);
and U569 (N_569,In_157,In_559);
nand U570 (N_570,In_121,In_119);
nor U571 (N_571,In_700,In_248);
nand U572 (N_572,In_488,In_489);
nand U573 (N_573,In_367,In_439);
nor U574 (N_574,In_356,In_28);
nand U575 (N_575,In_734,In_147);
and U576 (N_576,In_355,In_542);
and U577 (N_577,In_700,In_380);
nor U578 (N_578,In_656,In_537);
nand U579 (N_579,In_557,In_593);
or U580 (N_580,In_47,In_349);
nor U581 (N_581,In_113,In_707);
and U582 (N_582,In_724,In_643);
nand U583 (N_583,In_323,In_609);
nor U584 (N_584,In_147,In_659);
nand U585 (N_585,In_426,In_502);
or U586 (N_586,In_557,In_116);
nand U587 (N_587,In_575,In_143);
nand U588 (N_588,In_572,In_249);
and U589 (N_589,In_467,In_48);
nand U590 (N_590,In_117,In_377);
or U591 (N_591,In_361,In_678);
nor U592 (N_592,In_594,In_449);
and U593 (N_593,In_111,In_197);
nand U594 (N_594,In_629,In_483);
and U595 (N_595,In_682,In_158);
nand U596 (N_596,In_295,In_633);
nand U597 (N_597,In_450,In_220);
or U598 (N_598,In_62,In_550);
and U599 (N_599,In_716,In_338);
or U600 (N_600,In_0,In_640);
nor U601 (N_601,In_218,In_242);
or U602 (N_602,In_33,In_267);
nor U603 (N_603,In_17,In_442);
and U604 (N_604,In_40,In_29);
and U605 (N_605,In_205,In_368);
or U606 (N_606,In_187,In_642);
and U607 (N_607,In_299,In_212);
and U608 (N_608,In_267,In_10);
or U609 (N_609,In_66,In_376);
nand U610 (N_610,In_354,In_76);
or U611 (N_611,In_684,In_184);
nor U612 (N_612,In_114,In_639);
and U613 (N_613,In_731,In_711);
nor U614 (N_614,In_579,In_312);
and U615 (N_615,In_652,In_560);
or U616 (N_616,In_416,In_183);
or U617 (N_617,In_410,In_713);
or U618 (N_618,In_624,In_550);
nand U619 (N_619,In_181,In_56);
nand U620 (N_620,In_649,In_268);
or U621 (N_621,In_79,In_397);
or U622 (N_622,In_504,In_184);
or U623 (N_623,In_437,In_515);
nor U624 (N_624,In_15,In_317);
nand U625 (N_625,In_711,In_576);
and U626 (N_626,In_581,In_173);
nand U627 (N_627,In_724,In_226);
or U628 (N_628,In_370,In_335);
or U629 (N_629,In_200,In_1);
and U630 (N_630,In_48,In_280);
nor U631 (N_631,In_144,In_190);
or U632 (N_632,In_289,In_599);
nand U633 (N_633,In_429,In_14);
nor U634 (N_634,In_576,In_23);
and U635 (N_635,In_401,In_438);
nand U636 (N_636,In_478,In_194);
nand U637 (N_637,In_9,In_236);
and U638 (N_638,In_640,In_241);
or U639 (N_639,In_686,In_606);
and U640 (N_640,In_653,In_674);
and U641 (N_641,In_27,In_655);
nand U642 (N_642,In_339,In_208);
or U643 (N_643,In_198,In_201);
and U644 (N_644,In_121,In_478);
nand U645 (N_645,In_308,In_91);
nor U646 (N_646,In_54,In_4);
or U647 (N_647,In_117,In_390);
or U648 (N_648,In_628,In_263);
nor U649 (N_649,In_218,In_301);
nand U650 (N_650,In_727,In_402);
and U651 (N_651,In_456,In_200);
and U652 (N_652,In_631,In_15);
or U653 (N_653,In_494,In_242);
and U654 (N_654,In_23,In_286);
nand U655 (N_655,In_5,In_7);
nand U656 (N_656,In_210,In_233);
and U657 (N_657,In_699,In_500);
and U658 (N_658,In_317,In_519);
and U659 (N_659,In_285,In_20);
nand U660 (N_660,In_451,In_278);
and U661 (N_661,In_90,In_174);
and U662 (N_662,In_739,In_25);
nor U663 (N_663,In_464,In_142);
nand U664 (N_664,In_580,In_572);
or U665 (N_665,In_35,In_404);
nor U666 (N_666,In_390,In_738);
and U667 (N_667,In_490,In_591);
or U668 (N_668,In_510,In_551);
nor U669 (N_669,In_577,In_103);
and U670 (N_670,In_158,In_5);
nand U671 (N_671,In_647,In_413);
and U672 (N_672,In_163,In_517);
or U673 (N_673,In_704,In_481);
nor U674 (N_674,In_565,In_11);
nor U675 (N_675,In_222,In_150);
nand U676 (N_676,In_380,In_92);
nand U677 (N_677,In_529,In_13);
or U678 (N_678,In_301,In_735);
or U679 (N_679,In_720,In_21);
nor U680 (N_680,In_389,In_547);
nand U681 (N_681,In_278,In_419);
or U682 (N_682,In_389,In_358);
or U683 (N_683,In_184,In_366);
and U684 (N_684,In_476,In_89);
and U685 (N_685,In_296,In_196);
nand U686 (N_686,In_17,In_672);
and U687 (N_687,In_628,In_248);
nor U688 (N_688,In_394,In_32);
nand U689 (N_689,In_221,In_446);
and U690 (N_690,In_365,In_552);
and U691 (N_691,In_354,In_717);
and U692 (N_692,In_306,In_244);
nand U693 (N_693,In_542,In_696);
nand U694 (N_694,In_740,In_133);
and U695 (N_695,In_505,In_178);
nand U696 (N_696,In_16,In_437);
nand U697 (N_697,In_263,In_211);
or U698 (N_698,In_467,In_420);
and U699 (N_699,In_212,In_418);
and U700 (N_700,In_578,In_316);
nor U701 (N_701,In_12,In_104);
or U702 (N_702,In_534,In_75);
nand U703 (N_703,In_26,In_101);
or U704 (N_704,In_381,In_550);
and U705 (N_705,In_674,In_235);
nor U706 (N_706,In_98,In_54);
and U707 (N_707,In_339,In_119);
and U708 (N_708,In_58,In_60);
and U709 (N_709,In_423,In_273);
and U710 (N_710,In_388,In_208);
nand U711 (N_711,In_163,In_253);
nor U712 (N_712,In_335,In_490);
nor U713 (N_713,In_395,In_558);
and U714 (N_714,In_211,In_398);
or U715 (N_715,In_496,In_145);
or U716 (N_716,In_258,In_701);
or U717 (N_717,In_484,In_500);
and U718 (N_718,In_333,In_592);
or U719 (N_719,In_416,In_743);
and U720 (N_720,In_556,In_707);
nor U721 (N_721,In_722,In_130);
and U722 (N_722,In_683,In_446);
nor U723 (N_723,In_305,In_371);
and U724 (N_724,In_663,In_40);
nor U725 (N_725,In_402,In_624);
and U726 (N_726,In_206,In_97);
nor U727 (N_727,In_4,In_234);
nand U728 (N_728,In_351,In_497);
or U729 (N_729,In_659,In_600);
and U730 (N_730,In_322,In_344);
nand U731 (N_731,In_719,In_270);
xor U732 (N_732,In_521,In_320);
nor U733 (N_733,In_402,In_562);
and U734 (N_734,In_471,In_327);
and U735 (N_735,In_350,In_75);
nand U736 (N_736,In_523,In_282);
nand U737 (N_737,In_207,In_695);
nor U738 (N_738,In_138,In_179);
nand U739 (N_739,In_36,In_50);
nand U740 (N_740,In_310,In_343);
and U741 (N_741,In_232,In_76);
nand U742 (N_742,In_389,In_118);
or U743 (N_743,In_117,In_161);
and U744 (N_744,In_201,In_258);
nand U745 (N_745,In_412,In_42);
nor U746 (N_746,In_562,In_198);
nor U747 (N_747,In_132,In_177);
nand U748 (N_748,In_309,In_300);
nand U749 (N_749,In_18,In_390);
nor U750 (N_750,In_74,In_731);
nand U751 (N_751,In_63,In_407);
or U752 (N_752,In_349,In_358);
nor U753 (N_753,In_50,In_263);
and U754 (N_754,In_585,In_683);
and U755 (N_755,In_519,In_122);
nand U756 (N_756,In_352,In_524);
or U757 (N_757,In_172,In_132);
nand U758 (N_758,In_35,In_29);
and U759 (N_759,In_305,In_444);
nand U760 (N_760,In_137,In_436);
nor U761 (N_761,In_481,In_110);
or U762 (N_762,In_294,In_8);
nor U763 (N_763,In_74,In_77);
and U764 (N_764,In_402,In_392);
nand U765 (N_765,In_147,In_22);
nor U766 (N_766,In_472,In_191);
and U767 (N_767,In_728,In_100);
nand U768 (N_768,In_291,In_270);
and U769 (N_769,In_461,In_475);
nor U770 (N_770,In_360,In_243);
and U771 (N_771,In_192,In_451);
nor U772 (N_772,In_399,In_336);
or U773 (N_773,In_551,In_689);
nor U774 (N_774,In_491,In_302);
and U775 (N_775,In_656,In_405);
nor U776 (N_776,In_271,In_548);
nand U777 (N_777,In_655,In_231);
nor U778 (N_778,In_304,In_694);
and U779 (N_779,In_25,In_201);
nor U780 (N_780,In_518,In_727);
nand U781 (N_781,In_214,In_441);
nor U782 (N_782,In_657,In_238);
nor U783 (N_783,In_217,In_501);
nand U784 (N_784,In_378,In_662);
or U785 (N_785,In_746,In_465);
or U786 (N_786,In_580,In_647);
nand U787 (N_787,In_389,In_246);
nand U788 (N_788,In_618,In_514);
nor U789 (N_789,In_676,In_608);
nand U790 (N_790,In_552,In_289);
or U791 (N_791,In_458,In_725);
nor U792 (N_792,In_192,In_544);
or U793 (N_793,In_393,In_689);
nor U794 (N_794,In_155,In_327);
nor U795 (N_795,In_440,In_175);
and U796 (N_796,In_652,In_420);
or U797 (N_797,In_480,In_136);
nand U798 (N_798,In_102,In_540);
nor U799 (N_799,In_311,In_71);
or U800 (N_800,In_165,In_331);
or U801 (N_801,In_602,In_461);
nor U802 (N_802,In_650,In_681);
nand U803 (N_803,In_213,In_224);
or U804 (N_804,In_241,In_266);
nand U805 (N_805,In_2,In_693);
nand U806 (N_806,In_104,In_418);
or U807 (N_807,In_145,In_493);
nand U808 (N_808,In_225,In_695);
and U809 (N_809,In_489,In_4);
or U810 (N_810,In_98,In_184);
nor U811 (N_811,In_414,In_252);
nor U812 (N_812,In_719,In_656);
nor U813 (N_813,In_28,In_5);
nor U814 (N_814,In_384,In_400);
nor U815 (N_815,In_325,In_250);
nor U816 (N_816,In_390,In_537);
or U817 (N_817,In_5,In_588);
nor U818 (N_818,In_103,In_135);
and U819 (N_819,In_16,In_66);
xor U820 (N_820,In_171,In_87);
nor U821 (N_821,In_280,In_732);
or U822 (N_822,In_343,In_222);
and U823 (N_823,In_358,In_676);
nand U824 (N_824,In_515,In_477);
and U825 (N_825,In_440,In_685);
nand U826 (N_826,In_728,In_659);
or U827 (N_827,In_632,In_278);
and U828 (N_828,In_349,In_228);
and U829 (N_829,In_256,In_87);
or U830 (N_830,In_307,In_288);
nor U831 (N_831,In_680,In_717);
and U832 (N_832,In_651,In_550);
or U833 (N_833,In_401,In_407);
and U834 (N_834,In_619,In_158);
and U835 (N_835,In_422,In_399);
nor U836 (N_836,In_546,In_300);
and U837 (N_837,In_363,In_127);
nor U838 (N_838,In_99,In_698);
nand U839 (N_839,In_212,In_134);
and U840 (N_840,In_412,In_212);
nand U841 (N_841,In_159,In_241);
nand U842 (N_842,In_243,In_356);
or U843 (N_843,In_396,In_479);
and U844 (N_844,In_100,In_288);
nand U845 (N_845,In_105,In_87);
or U846 (N_846,In_236,In_7);
and U847 (N_847,In_176,In_242);
and U848 (N_848,In_655,In_459);
and U849 (N_849,In_366,In_699);
or U850 (N_850,In_196,In_147);
nor U851 (N_851,In_722,In_426);
and U852 (N_852,In_406,In_111);
and U853 (N_853,In_12,In_76);
nand U854 (N_854,In_123,In_464);
or U855 (N_855,In_30,In_427);
and U856 (N_856,In_410,In_729);
nor U857 (N_857,In_46,In_559);
nand U858 (N_858,In_418,In_298);
and U859 (N_859,In_394,In_453);
and U860 (N_860,In_432,In_364);
and U861 (N_861,In_189,In_715);
or U862 (N_862,In_504,In_291);
nand U863 (N_863,In_319,In_5);
nand U864 (N_864,In_614,In_51);
and U865 (N_865,In_150,In_407);
or U866 (N_866,In_183,In_120);
and U867 (N_867,In_382,In_31);
and U868 (N_868,In_286,In_183);
nor U869 (N_869,In_403,In_458);
nor U870 (N_870,In_333,In_516);
nor U871 (N_871,In_562,In_259);
nand U872 (N_872,In_621,In_489);
nand U873 (N_873,In_473,In_303);
nor U874 (N_874,In_633,In_491);
nor U875 (N_875,In_391,In_406);
and U876 (N_876,In_419,In_532);
and U877 (N_877,In_40,In_167);
or U878 (N_878,In_143,In_317);
or U879 (N_879,In_728,In_412);
nand U880 (N_880,In_744,In_88);
nand U881 (N_881,In_608,In_552);
or U882 (N_882,In_545,In_363);
or U883 (N_883,In_722,In_349);
nand U884 (N_884,In_295,In_196);
nor U885 (N_885,In_10,In_406);
and U886 (N_886,In_623,In_725);
nor U887 (N_887,In_746,In_378);
or U888 (N_888,In_644,In_91);
nand U889 (N_889,In_500,In_301);
or U890 (N_890,In_472,In_418);
nor U891 (N_891,In_70,In_741);
nor U892 (N_892,In_417,In_382);
nor U893 (N_893,In_393,In_746);
nand U894 (N_894,In_529,In_280);
or U895 (N_895,In_555,In_282);
and U896 (N_896,In_373,In_476);
nor U897 (N_897,In_615,In_725);
nor U898 (N_898,In_66,In_465);
nand U899 (N_899,In_46,In_642);
and U900 (N_900,In_10,In_438);
nor U901 (N_901,In_280,In_581);
nand U902 (N_902,In_217,In_534);
and U903 (N_903,In_100,In_139);
and U904 (N_904,In_62,In_126);
and U905 (N_905,In_25,In_26);
nor U906 (N_906,In_445,In_647);
nor U907 (N_907,In_407,In_509);
nand U908 (N_908,In_267,In_583);
and U909 (N_909,In_646,In_424);
nand U910 (N_910,In_592,In_76);
or U911 (N_911,In_506,In_49);
or U912 (N_912,In_683,In_90);
and U913 (N_913,In_486,In_706);
nor U914 (N_914,In_213,In_120);
xnor U915 (N_915,In_155,In_252);
nor U916 (N_916,In_624,In_388);
or U917 (N_917,In_270,In_548);
nor U918 (N_918,In_301,In_375);
and U919 (N_919,In_463,In_462);
nand U920 (N_920,In_649,In_209);
or U921 (N_921,In_280,In_194);
or U922 (N_922,In_524,In_107);
or U923 (N_923,In_384,In_719);
or U924 (N_924,In_402,In_576);
nor U925 (N_925,In_303,In_676);
or U926 (N_926,In_493,In_469);
and U927 (N_927,In_180,In_607);
or U928 (N_928,In_123,In_615);
or U929 (N_929,In_605,In_204);
and U930 (N_930,In_323,In_601);
nand U931 (N_931,In_264,In_213);
nor U932 (N_932,In_324,In_533);
nor U933 (N_933,In_575,In_185);
and U934 (N_934,In_327,In_738);
or U935 (N_935,In_610,In_48);
and U936 (N_936,In_734,In_27);
or U937 (N_937,In_458,In_123);
nor U938 (N_938,In_364,In_102);
or U939 (N_939,In_241,In_717);
nand U940 (N_940,In_24,In_19);
and U941 (N_941,In_648,In_226);
nor U942 (N_942,In_611,In_226);
or U943 (N_943,In_137,In_357);
or U944 (N_944,In_188,In_118);
nor U945 (N_945,In_361,In_129);
nor U946 (N_946,In_685,In_438);
nor U947 (N_947,In_489,In_694);
or U948 (N_948,In_579,In_250);
nand U949 (N_949,In_536,In_140);
or U950 (N_950,In_30,In_682);
nand U951 (N_951,In_493,In_633);
nor U952 (N_952,In_454,In_88);
and U953 (N_953,In_69,In_399);
or U954 (N_954,In_715,In_630);
nor U955 (N_955,In_221,In_97);
or U956 (N_956,In_299,In_43);
nor U957 (N_957,In_76,In_622);
nor U958 (N_958,In_277,In_441);
nand U959 (N_959,In_139,In_307);
or U960 (N_960,In_262,In_439);
nand U961 (N_961,In_305,In_542);
nor U962 (N_962,In_210,In_468);
or U963 (N_963,In_697,In_59);
nand U964 (N_964,In_556,In_40);
or U965 (N_965,In_22,In_297);
nor U966 (N_966,In_86,In_738);
or U967 (N_967,In_729,In_8);
nor U968 (N_968,In_529,In_723);
and U969 (N_969,In_672,In_641);
nand U970 (N_970,In_489,In_172);
nand U971 (N_971,In_499,In_49);
nor U972 (N_972,In_402,In_550);
nor U973 (N_973,In_373,In_609);
and U974 (N_974,In_94,In_712);
or U975 (N_975,In_174,In_161);
and U976 (N_976,In_396,In_242);
xor U977 (N_977,In_319,In_141);
nor U978 (N_978,In_563,In_499);
and U979 (N_979,In_211,In_215);
xnor U980 (N_980,In_87,In_521);
and U981 (N_981,In_207,In_487);
xnor U982 (N_982,In_132,In_492);
and U983 (N_983,In_739,In_353);
or U984 (N_984,In_692,In_664);
nor U985 (N_985,In_569,In_452);
or U986 (N_986,In_548,In_65);
nand U987 (N_987,In_529,In_553);
nand U988 (N_988,In_353,In_720);
nor U989 (N_989,In_704,In_83);
nand U990 (N_990,In_471,In_293);
or U991 (N_991,In_375,In_476);
nand U992 (N_992,In_600,In_597);
or U993 (N_993,In_592,In_406);
nor U994 (N_994,In_44,In_257);
nand U995 (N_995,In_331,In_644);
nand U996 (N_996,In_313,In_288);
nor U997 (N_997,In_103,In_102);
or U998 (N_998,In_653,In_168);
and U999 (N_999,In_324,In_374);
and U1000 (N_1000,In_486,In_40);
nor U1001 (N_1001,In_655,In_1);
nand U1002 (N_1002,In_136,In_588);
nand U1003 (N_1003,In_14,In_185);
and U1004 (N_1004,In_93,In_400);
or U1005 (N_1005,In_214,In_517);
nand U1006 (N_1006,In_554,In_364);
nand U1007 (N_1007,In_679,In_422);
nand U1008 (N_1008,In_342,In_741);
nand U1009 (N_1009,In_468,In_85);
nand U1010 (N_1010,In_40,In_393);
nor U1011 (N_1011,In_65,In_478);
nand U1012 (N_1012,In_76,In_641);
nor U1013 (N_1013,In_4,In_679);
or U1014 (N_1014,In_128,In_735);
nor U1015 (N_1015,In_487,In_643);
or U1016 (N_1016,In_672,In_89);
or U1017 (N_1017,In_34,In_265);
and U1018 (N_1018,In_572,In_431);
nand U1019 (N_1019,In_709,In_336);
and U1020 (N_1020,In_146,In_52);
and U1021 (N_1021,In_579,In_110);
or U1022 (N_1022,In_288,In_672);
nor U1023 (N_1023,In_387,In_6);
nand U1024 (N_1024,In_408,In_26);
nor U1025 (N_1025,In_327,In_573);
and U1026 (N_1026,In_455,In_595);
and U1027 (N_1027,In_536,In_87);
and U1028 (N_1028,In_233,In_417);
nor U1029 (N_1029,In_89,In_169);
nand U1030 (N_1030,In_405,In_310);
nor U1031 (N_1031,In_675,In_194);
nor U1032 (N_1032,In_252,In_616);
and U1033 (N_1033,In_356,In_90);
or U1034 (N_1034,In_348,In_467);
nand U1035 (N_1035,In_346,In_81);
nor U1036 (N_1036,In_266,In_249);
or U1037 (N_1037,In_199,In_517);
nand U1038 (N_1038,In_399,In_322);
and U1039 (N_1039,In_629,In_130);
and U1040 (N_1040,In_377,In_509);
nor U1041 (N_1041,In_77,In_466);
and U1042 (N_1042,In_563,In_139);
nand U1043 (N_1043,In_566,In_291);
or U1044 (N_1044,In_285,In_86);
and U1045 (N_1045,In_136,In_710);
and U1046 (N_1046,In_341,In_96);
or U1047 (N_1047,In_85,In_447);
nor U1048 (N_1048,In_18,In_126);
nand U1049 (N_1049,In_447,In_585);
nor U1050 (N_1050,In_160,In_358);
or U1051 (N_1051,In_747,In_21);
nor U1052 (N_1052,In_452,In_290);
nor U1053 (N_1053,In_191,In_674);
and U1054 (N_1054,In_466,In_172);
and U1055 (N_1055,In_710,In_534);
and U1056 (N_1056,In_49,In_236);
and U1057 (N_1057,In_306,In_108);
or U1058 (N_1058,In_163,In_123);
nor U1059 (N_1059,In_585,In_157);
nand U1060 (N_1060,In_248,In_527);
xnor U1061 (N_1061,In_646,In_222);
nor U1062 (N_1062,In_398,In_732);
xor U1063 (N_1063,In_108,In_37);
nand U1064 (N_1064,In_613,In_264);
and U1065 (N_1065,In_574,In_368);
nand U1066 (N_1066,In_594,In_120);
nand U1067 (N_1067,In_513,In_241);
and U1068 (N_1068,In_45,In_594);
and U1069 (N_1069,In_704,In_589);
or U1070 (N_1070,In_566,In_449);
nand U1071 (N_1071,In_4,In_10);
nor U1072 (N_1072,In_345,In_114);
nor U1073 (N_1073,In_650,In_497);
or U1074 (N_1074,In_282,In_524);
nand U1075 (N_1075,In_36,In_602);
nor U1076 (N_1076,In_117,In_731);
or U1077 (N_1077,In_225,In_388);
nand U1078 (N_1078,In_449,In_570);
xnor U1079 (N_1079,In_748,In_352);
or U1080 (N_1080,In_65,In_49);
nand U1081 (N_1081,In_77,In_587);
and U1082 (N_1082,In_44,In_314);
nand U1083 (N_1083,In_14,In_129);
and U1084 (N_1084,In_17,In_302);
nor U1085 (N_1085,In_119,In_212);
and U1086 (N_1086,In_205,In_389);
and U1087 (N_1087,In_725,In_674);
nor U1088 (N_1088,In_74,In_128);
nand U1089 (N_1089,In_723,In_200);
or U1090 (N_1090,In_456,In_214);
nand U1091 (N_1091,In_462,In_291);
nand U1092 (N_1092,In_318,In_130);
nand U1093 (N_1093,In_482,In_23);
and U1094 (N_1094,In_431,In_422);
nand U1095 (N_1095,In_176,In_453);
nor U1096 (N_1096,In_84,In_575);
nand U1097 (N_1097,In_308,In_234);
and U1098 (N_1098,In_405,In_549);
nand U1099 (N_1099,In_610,In_679);
nand U1100 (N_1100,In_12,In_202);
xnor U1101 (N_1101,In_183,In_480);
nor U1102 (N_1102,In_67,In_620);
and U1103 (N_1103,In_586,In_203);
and U1104 (N_1104,In_112,In_462);
nand U1105 (N_1105,In_59,In_193);
or U1106 (N_1106,In_678,In_242);
nor U1107 (N_1107,In_197,In_415);
or U1108 (N_1108,In_454,In_450);
nand U1109 (N_1109,In_244,In_742);
or U1110 (N_1110,In_196,In_179);
or U1111 (N_1111,In_527,In_347);
nand U1112 (N_1112,In_93,In_42);
nand U1113 (N_1113,In_213,In_59);
or U1114 (N_1114,In_572,In_399);
and U1115 (N_1115,In_558,In_203);
nand U1116 (N_1116,In_468,In_69);
nor U1117 (N_1117,In_659,In_545);
and U1118 (N_1118,In_540,In_232);
nand U1119 (N_1119,In_100,In_736);
nand U1120 (N_1120,In_253,In_373);
or U1121 (N_1121,In_387,In_238);
or U1122 (N_1122,In_670,In_366);
xor U1123 (N_1123,In_422,In_226);
nand U1124 (N_1124,In_497,In_498);
and U1125 (N_1125,In_662,In_257);
nand U1126 (N_1126,In_366,In_455);
nand U1127 (N_1127,In_529,In_469);
nand U1128 (N_1128,In_26,In_4);
nor U1129 (N_1129,In_293,In_510);
nor U1130 (N_1130,In_76,In_306);
nor U1131 (N_1131,In_604,In_298);
nand U1132 (N_1132,In_446,In_745);
nor U1133 (N_1133,In_133,In_529);
or U1134 (N_1134,In_30,In_119);
nor U1135 (N_1135,In_413,In_341);
xnor U1136 (N_1136,In_518,In_308);
and U1137 (N_1137,In_264,In_118);
nand U1138 (N_1138,In_248,In_528);
nand U1139 (N_1139,In_158,In_224);
or U1140 (N_1140,In_129,In_687);
nand U1141 (N_1141,In_105,In_64);
and U1142 (N_1142,In_414,In_441);
or U1143 (N_1143,In_465,In_567);
and U1144 (N_1144,In_300,In_357);
nor U1145 (N_1145,In_150,In_295);
nor U1146 (N_1146,In_333,In_580);
and U1147 (N_1147,In_502,In_197);
nand U1148 (N_1148,In_135,In_35);
or U1149 (N_1149,In_368,In_30);
nand U1150 (N_1150,In_700,In_343);
or U1151 (N_1151,In_344,In_239);
and U1152 (N_1152,In_586,In_86);
nand U1153 (N_1153,In_715,In_674);
nand U1154 (N_1154,In_212,In_78);
or U1155 (N_1155,In_523,In_399);
or U1156 (N_1156,In_656,In_552);
nand U1157 (N_1157,In_503,In_223);
xor U1158 (N_1158,In_71,In_14);
nor U1159 (N_1159,In_613,In_637);
and U1160 (N_1160,In_412,In_173);
or U1161 (N_1161,In_516,In_690);
or U1162 (N_1162,In_207,In_241);
nor U1163 (N_1163,In_655,In_578);
nand U1164 (N_1164,In_644,In_405);
or U1165 (N_1165,In_528,In_621);
nor U1166 (N_1166,In_694,In_138);
or U1167 (N_1167,In_31,In_702);
nor U1168 (N_1168,In_162,In_411);
xor U1169 (N_1169,In_558,In_176);
nand U1170 (N_1170,In_471,In_648);
or U1171 (N_1171,In_351,In_140);
or U1172 (N_1172,In_158,In_388);
or U1173 (N_1173,In_732,In_738);
or U1174 (N_1174,In_580,In_173);
or U1175 (N_1175,In_80,In_564);
or U1176 (N_1176,In_139,In_633);
or U1177 (N_1177,In_653,In_457);
nand U1178 (N_1178,In_650,In_439);
or U1179 (N_1179,In_426,In_595);
nor U1180 (N_1180,In_12,In_262);
nor U1181 (N_1181,In_700,In_236);
nand U1182 (N_1182,In_343,In_512);
nand U1183 (N_1183,In_542,In_320);
xnor U1184 (N_1184,In_111,In_472);
nor U1185 (N_1185,In_391,In_230);
nor U1186 (N_1186,In_563,In_400);
nand U1187 (N_1187,In_563,In_743);
and U1188 (N_1188,In_570,In_730);
nand U1189 (N_1189,In_481,In_533);
and U1190 (N_1190,In_370,In_537);
or U1191 (N_1191,In_491,In_246);
nor U1192 (N_1192,In_674,In_743);
and U1193 (N_1193,In_188,In_315);
and U1194 (N_1194,In_719,In_159);
and U1195 (N_1195,In_656,In_371);
nor U1196 (N_1196,In_595,In_187);
nor U1197 (N_1197,In_235,In_654);
or U1198 (N_1198,In_340,In_280);
nand U1199 (N_1199,In_665,In_441);
and U1200 (N_1200,In_300,In_613);
and U1201 (N_1201,In_149,In_588);
or U1202 (N_1202,In_130,In_725);
nor U1203 (N_1203,In_352,In_415);
and U1204 (N_1204,In_114,In_109);
and U1205 (N_1205,In_731,In_640);
or U1206 (N_1206,In_709,In_542);
or U1207 (N_1207,In_191,In_123);
or U1208 (N_1208,In_195,In_108);
nor U1209 (N_1209,In_202,In_152);
or U1210 (N_1210,In_346,In_128);
nor U1211 (N_1211,In_544,In_337);
and U1212 (N_1212,In_320,In_706);
nor U1213 (N_1213,In_230,In_429);
or U1214 (N_1214,In_399,In_43);
and U1215 (N_1215,In_432,In_445);
or U1216 (N_1216,In_591,In_667);
nand U1217 (N_1217,In_418,In_60);
and U1218 (N_1218,In_383,In_196);
and U1219 (N_1219,In_690,In_463);
or U1220 (N_1220,In_598,In_147);
nand U1221 (N_1221,In_382,In_700);
nand U1222 (N_1222,In_431,In_628);
or U1223 (N_1223,In_356,In_428);
nand U1224 (N_1224,In_375,In_49);
nor U1225 (N_1225,In_704,In_541);
nand U1226 (N_1226,In_443,In_199);
or U1227 (N_1227,In_506,In_382);
nand U1228 (N_1228,In_688,In_214);
or U1229 (N_1229,In_728,In_328);
nor U1230 (N_1230,In_338,In_587);
nor U1231 (N_1231,In_121,In_47);
and U1232 (N_1232,In_559,In_311);
nor U1233 (N_1233,In_239,In_329);
or U1234 (N_1234,In_133,In_496);
nor U1235 (N_1235,In_212,In_188);
nand U1236 (N_1236,In_200,In_36);
or U1237 (N_1237,In_718,In_552);
and U1238 (N_1238,In_430,In_166);
nand U1239 (N_1239,In_617,In_318);
or U1240 (N_1240,In_162,In_267);
nand U1241 (N_1241,In_549,In_716);
xor U1242 (N_1242,In_113,In_606);
nand U1243 (N_1243,In_293,In_22);
and U1244 (N_1244,In_722,In_148);
nand U1245 (N_1245,In_347,In_704);
nand U1246 (N_1246,In_14,In_550);
nand U1247 (N_1247,In_749,In_493);
nor U1248 (N_1248,In_350,In_151);
nand U1249 (N_1249,In_83,In_65);
or U1250 (N_1250,In_600,In_656);
nand U1251 (N_1251,In_53,In_411);
nand U1252 (N_1252,In_200,In_138);
or U1253 (N_1253,In_74,In_72);
nor U1254 (N_1254,In_174,In_331);
or U1255 (N_1255,In_560,In_625);
nand U1256 (N_1256,In_266,In_707);
nor U1257 (N_1257,In_342,In_353);
or U1258 (N_1258,In_690,In_410);
nand U1259 (N_1259,In_319,In_722);
nor U1260 (N_1260,In_488,In_273);
and U1261 (N_1261,In_45,In_591);
nor U1262 (N_1262,In_536,In_283);
xnor U1263 (N_1263,In_217,In_630);
nor U1264 (N_1264,In_378,In_296);
nand U1265 (N_1265,In_654,In_130);
or U1266 (N_1266,In_360,In_264);
nand U1267 (N_1267,In_458,In_531);
and U1268 (N_1268,In_124,In_143);
and U1269 (N_1269,In_711,In_298);
nand U1270 (N_1270,In_255,In_508);
and U1271 (N_1271,In_309,In_334);
or U1272 (N_1272,In_268,In_232);
or U1273 (N_1273,In_577,In_699);
nand U1274 (N_1274,In_277,In_131);
and U1275 (N_1275,In_242,In_71);
nor U1276 (N_1276,In_402,In_537);
and U1277 (N_1277,In_521,In_700);
and U1278 (N_1278,In_160,In_462);
nand U1279 (N_1279,In_538,In_207);
and U1280 (N_1280,In_131,In_285);
and U1281 (N_1281,In_447,In_354);
nor U1282 (N_1282,In_532,In_632);
and U1283 (N_1283,In_394,In_604);
or U1284 (N_1284,In_503,In_308);
and U1285 (N_1285,In_37,In_749);
nor U1286 (N_1286,In_736,In_480);
nor U1287 (N_1287,In_463,In_28);
nand U1288 (N_1288,In_699,In_642);
or U1289 (N_1289,In_202,In_378);
and U1290 (N_1290,In_342,In_621);
or U1291 (N_1291,In_199,In_595);
and U1292 (N_1292,In_403,In_206);
nand U1293 (N_1293,In_271,In_150);
or U1294 (N_1294,In_519,In_600);
and U1295 (N_1295,In_539,In_428);
nand U1296 (N_1296,In_310,In_736);
or U1297 (N_1297,In_27,In_492);
nor U1298 (N_1298,In_20,In_586);
and U1299 (N_1299,In_626,In_717);
and U1300 (N_1300,In_490,In_135);
nand U1301 (N_1301,In_677,In_336);
and U1302 (N_1302,In_42,In_104);
nand U1303 (N_1303,In_139,In_10);
or U1304 (N_1304,In_678,In_236);
or U1305 (N_1305,In_623,In_308);
nand U1306 (N_1306,In_249,In_160);
or U1307 (N_1307,In_442,In_325);
or U1308 (N_1308,In_140,In_91);
nand U1309 (N_1309,In_599,In_223);
nor U1310 (N_1310,In_433,In_348);
and U1311 (N_1311,In_581,In_546);
nand U1312 (N_1312,In_235,In_584);
nor U1313 (N_1313,In_256,In_371);
or U1314 (N_1314,In_384,In_730);
nor U1315 (N_1315,In_286,In_648);
and U1316 (N_1316,In_610,In_226);
and U1317 (N_1317,In_94,In_28);
nand U1318 (N_1318,In_318,In_394);
nand U1319 (N_1319,In_119,In_580);
nand U1320 (N_1320,In_209,In_356);
and U1321 (N_1321,In_714,In_236);
nand U1322 (N_1322,In_74,In_674);
or U1323 (N_1323,In_682,In_454);
and U1324 (N_1324,In_566,In_406);
nand U1325 (N_1325,In_651,In_267);
or U1326 (N_1326,In_228,In_379);
nand U1327 (N_1327,In_426,In_511);
nor U1328 (N_1328,In_407,In_641);
xnor U1329 (N_1329,In_280,In_234);
nor U1330 (N_1330,In_100,In_290);
or U1331 (N_1331,In_407,In_704);
nand U1332 (N_1332,In_615,In_371);
nor U1333 (N_1333,In_382,In_487);
nor U1334 (N_1334,In_28,In_9);
and U1335 (N_1335,In_735,In_604);
nor U1336 (N_1336,In_682,In_82);
and U1337 (N_1337,In_284,In_228);
nand U1338 (N_1338,In_477,In_248);
or U1339 (N_1339,In_46,In_621);
or U1340 (N_1340,In_107,In_681);
and U1341 (N_1341,In_595,In_318);
and U1342 (N_1342,In_318,In_173);
or U1343 (N_1343,In_142,In_372);
and U1344 (N_1344,In_652,In_305);
or U1345 (N_1345,In_271,In_725);
nor U1346 (N_1346,In_410,In_176);
or U1347 (N_1347,In_292,In_466);
or U1348 (N_1348,In_168,In_572);
and U1349 (N_1349,In_519,In_88);
xnor U1350 (N_1350,In_667,In_603);
nand U1351 (N_1351,In_166,In_537);
nor U1352 (N_1352,In_446,In_727);
and U1353 (N_1353,In_528,In_70);
nor U1354 (N_1354,In_301,In_169);
or U1355 (N_1355,In_201,In_458);
and U1356 (N_1356,In_527,In_201);
and U1357 (N_1357,In_320,In_150);
or U1358 (N_1358,In_717,In_219);
nand U1359 (N_1359,In_341,In_192);
and U1360 (N_1360,In_633,In_470);
and U1361 (N_1361,In_460,In_717);
or U1362 (N_1362,In_553,In_503);
nand U1363 (N_1363,In_403,In_266);
and U1364 (N_1364,In_556,In_646);
nand U1365 (N_1365,In_51,In_451);
or U1366 (N_1366,In_524,In_135);
and U1367 (N_1367,In_366,In_679);
nor U1368 (N_1368,In_39,In_386);
nand U1369 (N_1369,In_451,In_191);
nand U1370 (N_1370,In_286,In_11);
nand U1371 (N_1371,In_114,In_95);
or U1372 (N_1372,In_246,In_549);
xor U1373 (N_1373,In_287,In_243);
and U1374 (N_1374,In_109,In_281);
nand U1375 (N_1375,In_294,In_37);
nor U1376 (N_1376,In_320,In_579);
xor U1377 (N_1377,In_655,In_432);
and U1378 (N_1378,In_417,In_212);
nor U1379 (N_1379,In_295,In_514);
xnor U1380 (N_1380,In_4,In_669);
or U1381 (N_1381,In_631,In_349);
nor U1382 (N_1382,In_33,In_609);
xor U1383 (N_1383,In_647,In_365);
and U1384 (N_1384,In_152,In_147);
or U1385 (N_1385,In_699,In_398);
nor U1386 (N_1386,In_287,In_521);
nand U1387 (N_1387,In_649,In_439);
or U1388 (N_1388,In_391,In_707);
or U1389 (N_1389,In_18,In_479);
nand U1390 (N_1390,In_491,In_547);
nor U1391 (N_1391,In_475,In_270);
or U1392 (N_1392,In_729,In_698);
nand U1393 (N_1393,In_543,In_266);
nand U1394 (N_1394,In_545,In_667);
and U1395 (N_1395,In_611,In_168);
nor U1396 (N_1396,In_443,In_178);
or U1397 (N_1397,In_456,In_385);
and U1398 (N_1398,In_660,In_529);
and U1399 (N_1399,In_343,In_322);
nor U1400 (N_1400,In_397,In_42);
and U1401 (N_1401,In_194,In_46);
or U1402 (N_1402,In_163,In_215);
xor U1403 (N_1403,In_379,In_375);
nand U1404 (N_1404,In_445,In_93);
nor U1405 (N_1405,In_738,In_481);
and U1406 (N_1406,In_2,In_510);
and U1407 (N_1407,In_378,In_526);
nand U1408 (N_1408,In_15,In_170);
or U1409 (N_1409,In_669,In_708);
nor U1410 (N_1410,In_524,In_260);
or U1411 (N_1411,In_232,In_45);
or U1412 (N_1412,In_675,In_310);
nor U1413 (N_1413,In_641,In_564);
nand U1414 (N_1414,In_308,In_321);
and U1415 (N_1415,In_29,In_310);
and U1416 (N_1416,In_1,In_486);
or U1417 (N_1417,In_473,In_583);
nand U1418 (N_1418,In_717,In_502);
nor U1419 (N_1419,In_97,In_19);
or U1420 (N_1420,In_651,In_713);
or U1421 (N_1421,In_252,In_182);
nor U1422 (N_1422,In_584,In_130);
nor U1423 (N_1423,In_449,In_708);
or U1424 (N_1424,In_17,In_529);
or U1425 (N_1425,In_546,In_713);
and U1426 (N_1426,In_722,In_409);
nand U1427 (N_1427,In_573,In_553);
and U1428 (N_1428,In_20,In_168);
nand U1429 (N_1429,In_460,In_316);
nor U1430 (N_1430,In_645,In_0);
nor U1431 (N_1431,In_176,In_105);
nand U1432 (N_1432,In_169,In_249);
nand U1433 (N_1433,In_664,In_491);
nor U1434 (N_1434,In_46,In_655);
and U1435 (N_1435,In_368,In_17);
or U1436 (N_1436,In_534,In_423);
or U1437 (N_1437,In_639,In_51);
nor U1438 (N_1438,In_656,In_318);
nor U1439 (N_1439,In_285,In_78);
or U1440 (N_1440,In_101,In_339);
nor U1441 (N_1441,In_126,In_663);
nor U1442 (N_1442,In_637,In_501);
or U1443 (N_1443,In_49,In_734);
or U1444 (N_1444,In_257,In_369);
and U1445 (N_1445,In_127,In_402);
nand U1446 (N_1446,In_27,In_352);
or U1447 (N_1447,In_477,In_442);
nor U1448 (N_1448,In_642,In_573);
xnor U1449 (N_1449,In_582,In_282);
and U1450 (N_1450,In_83,In_79);
or U1451 (N_1451,In_413,In_502);
nor U1452 (N_1452,In_263,In_574);
or U1453 (N_1453,In_647,In_199);
nor U1454 (N_1454,In_406,In_333);
or U1455 (N_1455,In_24,In_22);
and U1456 (N_1456,In_61,In_735);
or U1457 (N_1457,In_593,In_412);
nor U1458 (N_1458,In_576,In_405);
nand U1459 (N_1459,In_120,In_722);
nor U1460 (N_1460,In_401,In_688);
and U1461 (N_1461,In_18,In_747);
nor U1462 (N_1462,In_66,In_438);
or U1463 (N_1463,In_218,In_359);
nand U1464 (N_1464,In_710,In_676);
nor U1465 (N_1465,In_233,In_444);
nand U1466 (N_1466,In_130,In_481);
or U1467 (N_1467,In_144,In_532);
nand U1468 (N_1468,In_234,In_482);
nor U1469 (N_1469,In_447,In_702);
and U1470 (N_1470,In_225,In_655);
nor U1471 (N_1471,In_723,In_28);
or U1472 (N_1472,In_738,In_302);
nand U1473 (N_1473,In_262,In_122);
or U1474 (N_1474,In_307,In_556);
nand U1475 (N_1475,In_39,In_78);
or U1476 (N_1476,In_224,In_357);
nand U1477 (N_1477,In_694,In_698);
or U1478 (N_1478,In_461,In_94);
nand U1479 (N_1479,In_422,In_604);
and U1480 (N_1480,In_552,In_180);
or U1481 (N_1481,In_467,In_140);
nand U1482 (N_1482,In_704,In_519);
or U1483 (N_1483,In_711,In_338);
or U1484 (N_1484,In_669,In_730);
and U1485 (N_1485,In_26,In_445);
nor U1486 (N_1486,In_43,In_603);
nor U1487 (N_1487,In_49,In_661);
nand U1488 (N_1488,In_486,In_384);
nor U1489 (N_1489,In_596,In_516);
nor U1490 (N_1490,In_641,In_156);
nand U1491 (N_1491,In_377,In_454);
nor U1492 (N_1492,In_368,In_707);
or U1493 (N_1493,In_550,In_718);
and U1494 (N_1494,In_26,In_82);
nand U1495 (N_1495,In_663,In_509);
or U1496 (N_1496,In_581,In_377);
nor U1497 (N_1497,In_10,In_35);
and U1498 (N_1498,In_596,In_677);
and U1499 (N_1499,In_647,In_551);
or U1500 (N_1500,In_454,In_461);
nand U1501 (N_1501,In_440,In_492);
nand U1502 (N_1502,In_186,In_59);
nand U1503 (N_1503,In_64,In_376);
and U1504 (N_1504,In_307,In_508);
nor U1505 (N_1505,In_688,In_423);
or U1506 (N_1506,In_262,In_385);
or U1507 (N_1507,In_482,In_250);
nor U1508 (N_1508,In_83,In_51);
nor U1509 (N_1509,In_76,In_656);
or U1510 (N_1510,In_65,In_658);
nor U1511 (N_1511,In_435,In_599);
or U1512 (N_1512,In_585,In_166);
nor U1513 (N_1513,In_541,In_333);
or U1514 (N_1514,In_634,In_76);
or U1515 (N_1515,In_144,In_255);
or U1516 (N_1516,In_543,In_35);
nor U1517 (N_1517,In_221,In_222);
nor U1518 (N_1518,In_725,In_561);
and U1519 (N_1519,In_740,In_374);
and U1520 (N_1520,In_307,In_100);
or U1521 (N_1521,In_644,In_715);
and U1522 (N_1522,In_390,In_73);
and U1523 (N_1523,In_94,In_246);
and U1524 (N_1524,In_91,In_6);
nand U1525 (N_1525,In_722,In_608);
and U1526 (N_1526,In_476,In_565);
or U1527 (N_1527,In_587,In_215);
nor U1528 (N_1528,In_323,In_526);
nand U1529 (N_1529,In_748,In_489);
and U1530 (N_1530,In_565,In_320);
or U1531 (N_1531,In_165,In_438);
or U1532 (N_1532,In_162,In_472);
nor U1533 (N_1533,In_673,In_627);
nand U1534 (N_1534,In_697,In_146);
nor U1535 (N_1535,In_127,In_271);
and U1536 (N_1536,In_62,In_233);
or U1537 (N_1537,In_18,In_461);
nor U1538 (N_1538,In_362,In_562);
or U1539 (N_1539,In_635,In_316);
nor U1540 (N_1540,In_743,In_497);
nor U1541 (N_1541,In_568,In_676);
and U1542 (N_1542,In_16,In_347);
xor U1543 (N_1543,In_8,In_309);
nand U1544 (N_1544,In_660,In_86);
nand U1545 (N_1545,In_530,In_269);
nor U1546 (N_1546,In_170,In_43);
or U1547 (N_1547,In_327,In_557);
nor U1548 (N_1548,In_685,In_487);
nor U1549 (N_1549,In_540,In_392);
or U1550 (N_1550,In_86,In_621);
nor U1551 (N_1551,In_452,In_258);
and U1552 (N_1552,In_280,In_594);
nand U1553 (N_1553,In_177,In_426);
and U1554 (N_1554,In_268,In_424);
and U1555 (N_1555,In_126,In_746);
and U1556 (N_1556,In_496,In_345);
nand U1557 (N_1557,In_388,In_478);
and U1558 (N_1558,In_455,In_551);
nor U1559 (N_1559,In_573,In_504);
nor U1560 (N_1560,In_78,In_549);
or U1561 (N_1561,In_536,In_163);
xnor U1562 (N_1562,In_57,In_594);
and U1563 (N_1563,In_375,In_322);
nor U1564 (N_1564,In_288,In_423);
nand U1565 (N_1565,In_595,In_600);
or U1566 (N_1566,In_209,In_326);
or U1567 (N_1567,In_673,In_536);
nand U1568 (N_1568,In_264,In_14);
and U1569 (N_1569,In_691,In_330);
nand U1570 (N_1570,In_466,In_627);
nand U1571 (N_1571,In_12,In_689);
or U1572 (N_1572,In_619,In_636);
nor U1573 (N_1573,In_16,In_440);
or U1574 (N_1574,In_621,In_273);
and U1575 (N_1575,In_39,In_161);
or U1576 (N_1576,In_308,In_221);
or U1577 (N_1577,In_289,In_210);
nor U1578 (N_1578,In_325,In_103);
nor U1579 (N_1579,In_605,In_481);
nor U1580 (N_1580,In_274,In_717);
nor U1581 (N_1581,In_27,In_235);
nand U1582 (N_1582,In_345,In_598);
and U1583 (N_1583,In_532,In_138);
nor U1584 (N_1584,In_424,In_36);
or U1585 (N_1585,In_722,In_691);
nand U1586 (N_1586,In_444,In_53);
nor U1587 (N_1587,In_641,In_682);
nand U1588 (N_1588,In_642,In_281);
nand U1589 (N_1589,In_562,In_17);
or U1590 (N_1590,In_198,In_463);
nor U1591 (N_1591,In_580,In_731);
nand U1592 (N_1592,In_184,In_361);
nor U1593 (N_1593,In_388,In_670);
and U1594 (N_1594,In_742,In_659);
nand U1595 (N_1595,In_302,In_642);
nand U1596 (N_1596,In_635,In_217);
or U1597 (N_1597,In_99,In_413);
nor U1598 (N_1598,In_235,In_602);
or U1599 (N_1599,In_457,In_699);
nand U1600 (N_1600,In_291,In_339);
and U1601 (N_1601,In_75,In_336);
and U1602 (N_1602,In_44,In_210);
nor U1603 (N_1603,In_735,In_188);
nor U1604 (N_1604,In_415,In_111);
and U1605 (N_1605,In_594,In_484);
nand U1606 (N_1606,In_69,In_708);
and U1607 (N_1607,In_599,In_651);
xnor U1608 (N_1608,In_520,In_110);
or U1609 (N_1609,In_359,In_520);
or U1610 (N_1610,In_14,In_571);
or U1611 (N_1611,In_471,In_255);
nor U1612 (N_1612,In_293,In_267);
nor U1613 (N_1613,In_353,In_615);
and U1614 (N_1614,In_31,In_744);
nor U1615 (N_1615,In_65,In_206);
nand U1616 (N_1616,In_313,In_411);
nor U1617 (N_1617,In_501,In_116);
and U1618 (N_1618,In_525,In_13);
or U1619 (N_1619,In_517,In_458);
nor U1620 (N_1620,In_642,In_543);
or U1621 (N_1621,In_448,In_159);
nand U1622 (N_1622,In_429,In_535);
nor U1623 (N_1623,In_637,In_44);
nand U1624 (N_1624,In_217,In_416);
nand U1625 (N_1625,In_650,In_501);
nor U1626 (N_1626,In_133,In_604);
nor U1627 (N_1627,In_430,In_605);
nor U1628 (N_1628,In_643,In_611);
nand U1629 (N_1629,In_205,In_447);
and U1630 (N_1630,In_487,In_273);
and U1631 (N_1631,In_524,In_111);
nand U1632 (N_1632,In_293,In_682);
nand U1633 (N_1633,In_648,In_167);
or U1634 (N_1634,In_46,In_309);
and U1635 (N_1635,In_210,In_111);
or U1636 (N_1636,In_446,In_359);
nor U1637 (N_1637,In_21,In_302);
or U1638 (N_1638,In_53,In_453);
nand U1639 (N_1639,In_379,In_57);
or U1640 (N_1640,In_19,In_431);
nor U1641 (N_1641,In_400,In_42);
or U1642 (N_1642,In_221,In_160);
or U1643 (N_1643,In_510,In_9);
or U1644 (N_1644,In_336,In_521);
and U1645 (N_1645,In_317,In_666);
nor U1646 (N_1646,In_470,In_525);
nand U1647 (N_1647,In_410,In_32);
or U1648 (N_1648,In_433,In_676);
xor U1649 (N_1649,In_692,In_642);
nor U1650 (N_1650,In_724,In_237);
and U1651 (N_1651,In_544,In_288);
or U1652 (N_1652,In_49,In_59);
nand U1653 (N_1653,In_614,In_584);
and U1654 (N_1654,In_396,In_15);
nor U1655 (N_1655,In_666,In_143);
and U1656 (N_1656,In_38,In_192);
and U1657 (N_1657,In_366,In_704);
nand U1658 (N_1658,In_288,In_523);
nand U1659 (N_1659,In_382,In_308);
nand U1660 (N_1660,In_478,In_329);
nand U1661 (N_1661,In_162,In_663);
nand U1662 (N_1662,In_370,In_308);
and U1663 (N_1663,In_533,In_363);
or U1664 (N_1664,In_367,In_410);
nor U1665 (N_1665,In_538,In_379);
nand U1666 (N_1666,In_688,In_81);
nor U1667 (N_1667,In_199,In_33);
or U1668 (N_1668,In_632,In_342);
nor U1669 (N_1669,In_251,In_462);
nand U1670 (N_1670,In_609,In_392);
or U1671 (N_1671,In_52,In_241);
nor U1672 (N_1672,In_89,In_301);
and U1673 (N_1673,In_627,In_119);
or U1674 (N_1674,In_304,In_370);
nand U1675 (N_1675,In_583,In_682);
and U1676 (N_1676,In_630,In_634);
or U1677 (N_1677,In_507,In_631);
and U1678 (N_1678,In_129,In_127);
and U1679 (N_1679,In_729,In_96);
or U1680 (N_1680,In_453,In_155);
nor U1681 (N_1681,In_315,In_314);
and U1682 (N_1682,In_591,In_421);
nor U1683 (N_1683,In_305,In_203);
nand U1684 (N_1684,In_235,In_273);
or U1685 (N_1685,In_215,In_573);
nand U1686 (N_1686,In_4,In_428);
and U1687 (N_1687,In_736,In_731);
or U1688 (N_1688,In_222,In_100);
nor U1689 (N_1689,In_203,In_655);
nand U1690 (N_1690,In_516,In_275);
and U1691 (N_1691,In_60,In_578);
nand U1692 (N_1692,In_688,In_710);
or U1693 (N_1693,In_514,In_355);
or U1694 (N_1694,In_591,In_267);
and U1695 (N_1695,In_646,In_358);
nand U1696 (N_1696,In_682,In_346);
nor U1697 (N_1697,In_51,In_479);
nor U1698 (N_1698,In_488,In_632);
xor U1699 (N_1699,In_280,In_229);
nand U1700 (N_1700,In_628,In_428);
nand U1701 (N_1701,In_691,In_704);
or U1702 (N_1702,In_209,In_131);
nand U1703 (N_1703,In_370,In_21);
nand U1704 (N_1704,In_295,In_341);
or U1705 (N_1705,In_151,In_280);
nand U1706 (N_1706,In_382,In_643);
and U1707 (N_1707,In_121,In_155);
or U1708 (N_1708,In_304,In_343);
or U1709 (N_1709,In_360,In_565);
or U1710 (N_1710,In_336,In_285);
and U1711 (N_1711,In_91,In_479);
xor U1712 (N_1712,In_694,In_227);
and U1713 (N_1713,In_377,In_551);
and U1714 (N_1714,In_685,In_601);
and U1715 (N_1715,In_318,In_150);
nor U1716 (N_1716,In_434,In_668);
and U1717 (N_1717,In_597,In_664);
nand U1718 (N_1718,In_695,In_530);
nand U1719 (N_1719,In_201,In_505);
and U1720 (N_1720,In_745,In_470);
nand U1721 (N_1721,In_652,In_36);
nor U1722 (N_1722,In_338,In_119);
nor U1723 (N_1723,In_602,In_363);
nor U1724 (N_1724,In_415,In_74);
or U1725 (N_1725,In_574,In_223);
nand U1726 (N_1726,In_556,In_317);
nor U1727 (N_1727,In_256,In_439);
nor U1728 (N_1728,In_413,In_79);
and U1729 (N_1729,In_76,In_531);
nand U1730 (N_1730,In_723,In_6);
nor U1731 (N_1731,In_70,In_321);
and U1732 (N_1732,In_361,In_76);
or U1733 (N_1733,In_673,In_699);
or U1734 (N_1734,In_135,In_170);
or U1735 (N_1735,In_691,In_196);
nor U1736 (N_1736,In_334,In_238);
and U1737 (N_1737,In_184,In_535);
nor U1738 (N_1738,In_541,In_35);
nor U1739 (N_1739,In_317,In_734);
or U1740 (N_1740,In_24,In_76);
xnor U1741 (N_1741,In_124,In_636);
and U1742 (N_1742,In_278,In_363);
nor U1743 (N_1743,In_19,In_126);
or U1744 (N_1744,In_436,In_361);
nor U1745 (N_1745,In_626,In_593);
or U1746 (N_1746,In_435,In_61);
nand U1747 (N_1747,In_703,In_741);
and U1748 (N_1748,In_375,In_744);
and U1749 (N_1749,In_671,In_75);
or U1750 (N_1750,In_250,In_278);
nor U1751 (N_1751,In_349,In_611);
nand U1752 (N_1752,In_142,In_221);
and U1753 (N_1753,In_260,In_526);
or U1754 (N_1754,In_675,In_154);
and U1755 (N_1755,In_683,In_61);
or U1756 (N_1756,In_71,In_684);
nand U1757 (N_1757,In_679,In_533);
and U1758 (N_1758,In_126,In_69);
nor U1759 (N_1759,In_427,In_523);
nand U1760 (N_1760,In_283,In_598);
nand U1761 (N_1761,In_660,In_293);
or U1762 (N_1762,In_213,In_453);
nand U1763 (N_1763,In_633,In_181);
nand U1764 (N_1764,In_582,In_279);
or U1765 (N_1765,In_450,In_170);
nand U1766 (N_1766,In_161,In_403);
nor U1767 (N_1767,In_345,In_71);
or U1768 (N_1768,In_286,In_52);
and U1769 (N_1769,In_358,In_455);
or U1770 (N_1770,In_655,In_522);
nor U1771 (N_1771,In_56,In_596);
nor U1772 (N_1772,In_316,In_684);
nand U1773 (N_1773,In_217,In_32);
or U1774 (N_1774,In_311,In_473);
and U1775 (N_1775,In_504,In_496);
nand U1776 (N_1776,In_533,In_322);
and U1777 (N_1777,In_430,In_128);
nand U1778 (N_1778,In_621,In_257);
or U1779 (N_1779,In_426,In_72);
or U1780 (N_1780,In_647,In_612);
or U1781 (N_1781,In_475,In_483);
or U1782 (N_1782,In_444,In_558);
nor U1783 (N_1783,In_258,In_446);
nor U1784 (N_1784,In_248,In_278);
nand U1785 (N_1785,In_586,In_315);
nor U1786 (N_1786,In_547,In_181);
nor U1787 (N_1787,In_129,In_583);
nand U1788 (N_1788,In_99,In_185);
and U1789 (N_1789,In_399,In_224);
nor U1790 (N_1790,In_133,In_395);
or U1791 (N_1791,In_712,In_547);
or U1792 (N_1792,In_465,In_693);
and U1793 (N_1793,In_222,In_654);
nor U1794 (N_1794,In_663,In_421);
or U1795 (N_1795,In_726,In_199);
nor U1796 (N_1796,In_379,In_561);
or U1797 (N_1797,In_592,In_67);
or U1798 (N_1798,In_610,In_44);
nor U1799 (N_1799,In_689,In_362);
and U1800 (N_1800,In_65,In_139);
nor U1801 (N_1801,In_437,In_341);
nor U1802 (N_1802,In_261,In_482);
and U1803 (N_1803,In_411,In_661);
nor U1804 (N_1804,In_610,In_189);
or U1805 (N_1805,In_606,In_94);
and U1806 (N_1806,In_197,In_303);
and U1807 (N_1807,In_44,In_275);
nand U1808 (N_1808,In_708,In_218);
or U1809 (N_1809,In_13,In_44);
or U1810 (N_1810,In_209,In_599);
or U1811 (N_1811,In_457,In_79);
or U1812 (N_1812,In_513,In_272);
and U1813 (N_1813,In_354,In_559);
and U1814 (N_1814,In_134,In_355);
and U1815 (N_1815,In_224,In_344);
or U1816 (N_1816,In_95,In_677);
nor U1817 (N_1817,In_696,In_358);
or U1818 (N_1818,In_268,In_505);
nor U1819 (N_1819,In_16,In_23);
and U1820 (N_1820,In_266,In_151);
and U1821 (N_1821,In_365,In_706);
nor U1822 (N_1822,In_639,In_484);
nor U1823 (N_1823,In_484,In_356);
nor U1824 (N_1824,In_599,In_464);
nor U1825 (N_1825,In_189,In_29);
or U1826 (N_1826,In_515,In_446);
nor U1827 (N_1827,In_318,In_100);
nand U1828 (N_1828,In_101,In_269);
or U1829 (N_1829,In_246,In_49);
and U1830 (N_1830,In_113,In_335);
nor U1831 (N_1831,In_701,In_225);
nand U1832 (N_1832,In_435,In_140);
nor U1833 (N_1833,In_454,In_371);
and U1834 (N_1834,In_458,In_474);
nand U1835 (N_1835,In_439,In_306);
or U1836 (N_1836,In_235,In_416);
and U1837 (N_1837,In_247,In_337);
nor U1838 (N_1838,In_300,In_327);
and U1839 (N_1839,In_348,In_74);
nand U1840 (N_1840,In_448,In_63);
or U1841 (N_1841,In_141,In_267);
and U1842 (N_1842,In_207,In_450);
nor U1843 (N_1843,In_82,In_526);
or U1844 (N_1844,In_89,In_271);
nor U1845 (N_1845,In_279,In_347);
and U1846 (N_1846,In_602,In_533);
nor U1847 (N_1847,In_365,In_593);
or U1848 (N_1848,In_462,In_500);
nor U1849 (N_1849,In_690,In_506);
and U1850 (N_1850,In_78,In_522);
nor U1851 (N_1851,In_260,In_307);
or U1852 (N_1852,In_437,In_669);
nor U1853 (N_1853,In_579,In_584);
or U1854 (N_1854,In_643,In_698);
and U1855 (N_1855,In_543,In_34);
or U1856 (N_1856,In_407,In_577);
nor U1857 (N_1857,In_712,In_238);
and U1858 (N_1858,In_134,In_375);
or U1859 (N_1859,In_747,In_262);
nor U1860 (N_1860,In_41,In_561);
and U1861 (N_1861,In_535,In_225);
nand U1862 (N_1862,In_693,In_380);
nand U1863 (N_1863,In_196,In_140);
and U1864 (N_1864,In_677,In_479);
nand U1865 (N_1865,In_12,In_30);
nor U1866 (N_1866,In_389,In_643);
or U1867 (N_1867,In_579,In_175);
nand U1868 (N_1868,In_456,In_727);
nand U1869 (N_1869,In_622,In_303);
nor U1870 (N_1870,In_642,In_209);
nand U1871 (N_1871,In_552,In_112);
nor U1872 (N_1872,In_600,In_310);
or U1873 (N_1873,In_289,In_630);
nor U1874 (N_1874,In_155,In_329);
and U1875 (N_1875,In_40,In_591);
nand U1876 (N_1876,In_666,In_25);
or U1877 (N_1877,In_75,In_183);
nand U1878 (N_1878,In_749,In_349);
and U1879 (N_1879,In_509,In_301);
nor U1880 (N_1880,In_356,In_194);
nand U1881 (N_1881,In_639,In_201);
and U1882 (N_1882,In_212,In_104);
and U1883 (N_1883,In_106,In_597);
nand U1884 (N_1884,In_38,In_342);
or U1885 (N_1885,In_86,In_189);
nor U1886 (N_1886,In_304,In_396);
or U1887 (N_1887,In_404,In_732);
nor U1888 (N_1888,In_415,In_681);
nor U1889 (N_1889,In_356,In_737);
nand U1890 (N_1890,In_67,In_157);
and U1891 (N_1891,In_536,In_356);
nor U1892 (N_1892,In_31,In_128);
or U1893 (N_1893,In_113,In_285);
and U1894 (N_1894,In_161,In_362);
or U1895 (N_1895,In_548,In_576);
nand U1896 (N_1896,In_562,In_130);
or U1897 (N_1897,In_457,In_10);
nand U1898 (N_1898,In_389,In_642);
nand U1899 (N_1899,In_229,In_404);
nand U1900 (N_1900,In_568,In_48);
nand U1901 (N_1901,In_222,In_553);
and U1902 (N_1902,In_476,In_558);
nor U1903 (N_1903,In_169,In_255);
nor U1904 (N_1904,In_262,In_389);
and U1905 (N_1905,In_736,In_179);
nand U1906 (N_1906,In_732,In_622);
and U1907 (N_1907,In_55,In_334);
nor U1908 (N_1908,In_45,In_490);
or U1909 (N_1909,In_398,In_694);
or U1910 (N_1910,In_600,In_70);
and U1911 (N_1911,In_643,In_447);
and U1912 (N_1912,In_612,In_427);
nor U1913 (N_1913,In_713,In_293);
nand U1914 (N_1914,In_119,In_426);
nand U1915 (N_1915,In_295,In_329);
or U1916 (N_1916,In_660,In_96);
nor U1917 (N_1917,In_600,In_40);
nor U1918 (N_1918,In_162,In_194);
or U1919 (N_1919,In_275,In_569);
nand U1920 (N_1920,In_105,In_700);
nor U1921 (N_1921,In_168,In_7);
nor U1922 (N_1922,In_576,In_52);
or U1923 (N_1923,In_601,In_332);
nor U1924 (N_1924,In_64,In_34);
nor U1925 (N_1925,In_520,In_679);
nor U1926 (N_1926,In_238,In_290);
nand U1927 (N_1927,In_175,In_157);
or U1928 (N_1928,In_96,In_114);
or U1929 (N_1929,In_320,In_23);
or U1930 (N_1930,In_531,In_290);
nand U1931 (N_1931,In_521,In_648);
and U1932 (N_1932,In_205,In_217);
nand U1933 (N_1933,In_36,In_677);
and U1934 (N_1934,In_678,In_624);
nor U1935 (N_1935,In_128,In_456);
nand U1936 (N_1936,In_676,In_466);
xor U1937 (N_1937,In_369,In_712);
nand U1938 (N_1938,In_334,In_428);
nand U1939 (N_1939,In_669,In_610);
nand U1940 (N_1940,In_512,In_668);
xnor U1941 (N_1941,In_153,In_650);
nor U1942 (N_1942,In_368,In_251);
nand U1943 (N_1943,In_279,In_108);
nor U1944 (N_1944,In_417,In_564);
nor U1945 (N_1945,In_193,In_746);
nand U1946 (N_1946,In_498,In_210);
nand U1947 (N_1947,In_255,In_83);
nand U1948 (N_1948,In_454,In_274);
or U1949 (N_1949,In_706,In_406);
nor U1950 (N_1950,In_172,In_245);
nand U1951 (N_1951,In_133,In_429);
nand U1952 (N_1952,In_464,In_303);
nand U1953 (N_1953,In_658,In_201);
or U1954 (N_1954,In_91,In_61);
and U1955 (N_1955,In_679,In_88);
xor U1956 (N_1956,In_210,In_201);
nor U1957 (N_1957,In_554,In_57);
and U1958 (N_1958,In_174,In_181);
and U1959 (N_1959,In_739,In_173);
or U1960 (N_1960,In_185,In_239);
nor U1961 (N_1961,In_728,In_122);
and U1962 (N_1962,In_395,In_696);
or U1963 (N_1963,In_338,In_593);
or U1964 (N_1964,In_404,In_211);
and U1965 (N_1965,In_392,In_399);
and U1966 (N_1966,In_697,In_310);
or U1967 (N_1967,In_698,In_228);
nor U1968 (N_1968,In_204,In_183);
or U1969 (N_1969,In_513,In_737);
nand U1970 (N_1970,In_227,In_6);
nor U1971 (N_1971,In_470,In_689);
or U1972 (N_1972,In_647,In_107);
or U1973 (N_1973,In_117,In_115);
and U1974 (N_1974,In_320,In_498);
or U1975 (N_1975,In_521,In_133);
nor U1976 (N_1976,In_538,In_181);
or U1977 (N_1977,In_62,In_433);
and U1978 (N_1978,In_223,In_118);
nand U1979 (N_1979,In_178,In_303);
nor U1980 (N_1980,In_534,In_228);
or U1981 (N_1981,In_258,In_139);
nand U1982 (N_1982,In_155,In_611);
nand U1983 (N_1983,In_728,In_502);
or U1984 (N_1984,In_135,In_706);
and U1985 (N_1985,In_689,In_390);
and U1986 (N_1986,In_549,In_452);
or U1987 (N_1987,In_107,In_330);
nor U1988 (N_1988,In_422,In_415);
nand U1989 (N_1989,In_555,In_71);
nand U1990 (N_1990,In_235,In_282);
nor U1991 (N_1991,In_601,In_347);
nor U1992 (N_1992,In_208,In_343);
nor U1993 (N_1993,In_30,In_317);
nand U1994 (N_1994,In_451,In_109);
nor U1995 (N_1995,In_552,In_510);
or U1996 (N_1996,In_320,In_366);
nand U1997 (N_1997,In_734,In_399);
xnor U1998 (N_1998,In_234,In_390);
or U1999 (N_1999,In_47,In_616);
or U2000 (N_2000,In_235,In_531);
nand U2001 (N_2001,In_94,In_508);
or U2002 (N_2002,In_409,In_405);
nor U2003 (N_2003,In_184,In_214);
nand U2004 (N_2004,In_129,In_60);
or U2005 (N_2005,In_540,In_431);
nand U2006 (N_2006,In_657,In_257);
and U2007 (N_2007,In_106,In_3);
xor U2008 (N_2008,In_670,In_402);
and U2009 (N_2009,In_392,In_248);
or U2010 (N_2010,In_58,In_130);
nor U2011 (N_2011,In_664,In_42);
nor U2012 (N_2012,In_164,In_143);
and U2013 (N_2013,In_597,In_642);
nand U2014 (N_2014,In_671,In_449);
nor U2015 (N_2015,In_199,In_632);
or U2016 (N_2016,In_480,In_231);
nand U2017 (N_2017,In_319,In_339);
and U2018 (N_2018,In_455,In_357);
or U2019 (N_2019,In_385,In_265);
nor U2020 (N_2020,In_269,In_431);
nor U2021 (N_2021,In_136,In_105);
nand U2022 (N_2022,In_225,In_661);
or U2023 (N_2023,In_721,In_67);
or U2024 (N_2024,In_730,In_673);
nand U2025 (N_2025,In_702,In_136);
and U2026 (N_2026,In_45,In_379);
or U2027 (N_2027,In_519,In_58);
nand U2028 (N_2028,In_424,In_516);
nor U2029 (N_2029,In_147,In_49);
nand U2030 (N_2030,In_703,In_20);
and U2031 (N_2031,In_713,In_608);
nor U2032 (N_2032,In_415,In_227);
or U2033 (N_2033,In_638,In_209);
nor U2034 (N_2034,In_135,In_373);
nor U2035 (N_2035,In_576,In_749);
nand U2036 (N_2036,In_479,In_12);
and U2037 (N_2037,In_82,In_645);
nor U2038 (N_2038,In_493,In_668);
or U2039 (N_2039,In_742,In_55);
and U2040 (N_2040,In_561,In_273);
nand U2041 (N_2041,In_738,In_358);
nor U2042 (N_2042,In_708,In_467);
nor U2043 (N_2043,In_413,In_267);
or U2044 (N_2044,In_40,In_341);
nor U2045 (N_2045,In_693,In_674);
nor U2046 (N_2046,In_629,In_105);
nor U2047 (N_2047,In_290,In_125);
nor U2048 (N_2048,In_461,In_719);
or U2049 (N_2049,In_334,In_379);
and U2050 (N_2050,In_183,In_717);
nor U2051 (N_2051,In_236,In_443);
nor U2052 (N_2052,In_285,In_587);
nand U2053 (N_2053,In_430,In_684);
or U2054 (N_2054,In_571,In_150);
or U2055 (N_2055,In_222,In_442);
nand U2056 (N_2056,In_154,In_625);
or U2057 (N_2057,In_593,In_350);
and U2058 (N_2058,In_251,In_463);
nand U2059 (N_2059,In_484,In_54);
nor U2060 (N_2060,In_124,In_635);
and U2061 (N_2061,In_685,In_90);
or U2062 (N_2062,In_113,In_121);
nand U2063 (N_2063,In_283,In_204);
nor U2064 (N_2064,In_204,In_165);
and U2065 (N_2065,In_588,In_73);
nand U2066 (N_2066,In_548,In_538);
or U2067 (N_2067,In_128,In_221);
and U2068 (N_2068,In_579,In_427);
nor U2069 (N_2069,In_398,In_361);
nor U2070 (N_2070,In_527,In_420);
nand U2071 (N_2071,In_533,In_349);
xor U2072 (N_2072,In_739,In_548);
or U2073 (N_2073,In_641,In_368);
nor U2074 (N_2074,In_103,In_442);
nor U2075 (N_2075,In_535,In_713);
nor U2076 (N_2076,In_4,In_555);
nor U2077 (N_2077,In_601,In_619);
and U2078 (N_2078,In_667,In_581);
or U2079 (N_2079,In_739,In_484);
and U2080 (N_2080,In_184,In_224);
nor U2081 (N_2081,In_118,In_225);
nand U2082 (N_2082,In_576,In_140);
nand U2083 (N_2083,In_260,In_525);
and U2084 (N_2084,In_277,In_491);
nor U2085 (N_2085,In_467,In_383);
nand U2086 (N_2086,In_231,In_736);
or U2087 (N_2087,In_141,In_393);
nor U2088 (N_2088,In_97,In_646);
and U2089 (N_2089,In_464,In_630);
nor U2090 (N_2090,In_581,In_16);
and U2091 (N_2091,In_702,In_679);
nand U2092 (N_2092,In_629,In_214);
nor U2093 (N_2093,In_518,In_420);
and U2094 (N_2094,In_91,In_382);
or U2095 (N_2095,In_491,In_428);
or U2096 (N_2096,In_338,In_294);
and U2097 (N_2097,In_451,In_715);
nand U2098 (N_2098,In_503,In_718);
nor U2099 (N_2099,In_414,In_295);
or U2100 (N_2100,In_339,In_518);
nor U2101 (N_2101,In_253,In_380);
nand U2102 (N_2102,In_330,In_493);
and U2103 (N_2103,In_302,In_235);
nand U2104 (N_2104,In_19,In_516);
and U2105 (N_2105,In_76,In_235);
or U2106 (N_2106,In_66,In_584);
nand U2107 (N_2107,In_598,In_164);
or U2108 (N_2108,In_723,In_52);
nand U2109 (N_2109,In_351,In_1);
nor U2110 (N_2110,In_382,In_376);
and U2111 (N_2111,In_137,In_420);
or U2112 (N_2112,In_566,In_678);
or U2113 (N_2113,In_136,In_421);
or U2114 (N_2114,In_427,In_198);
nor U2115 (N_2115,In_509,In_471);
or U2116 (N_2116,In_319,In_175);
nor U2117 (N_2117,In_220,In_562);
or U2118 (N_2118,In_138,In_663);
nand U2119 (N_2119,In_174,In_89);
or U2120 (N_2120,In_588,In_682);
xor U2121 (N_2121,In_241,In_75);
nand U2122 (N_2122,In_335,In_243);
nand U2123 (N_2123,In_91,In_483);
and U2124 (N_2124,In_301,In_88);
or U2125 (N_2125,In_334,In_647);
or U2126 (N_2126,In_707,In_392);
nor U2127 (N_2127,In_139,In_133);
and U2128 (N_2128,In_201,In_397);
and U2129 (N_2129,In_109,In_521);
nor U2130 (N_2130,In_303,In_698);
nand U2131 (N_2131,In_455,In_749);
nor U2132 (N_2132,In_680,In_237);
or U2133 (N_2133,In_106,In_704);
nor U2134 (N_2134,In_737,In_115);
or U2135 (N_2135,In_76,In_300);
or U2136 (N_2136,In_314,In_334);
and U2137 (N_2137,In_29,In_459);
nor U2138 (N_2138,In_538,In_695);
nor U2139 (N_2139,In_70,In_360);
nand U2140 (N_2140,In_344,In_215);
nor U2141 (N_2141,In_214,In_52);
nor U2142 (N_2142,In_280,In_394);
nor U2143 (N_2143,In_443,In_619);
nor U2144 (N_2144,In_506,In_502);
nor U2145 (N_2145,In_121,In_715);
and U2146 (N_2146,In_586,In_701);
and U2147 (N_2147,In_456,In_690);
nor U2148 (N_2148,In_653,In_376);
nand U2149 (N_2149,In_154,In_304);
nor U2150 (N_2150,In_712,In_739);
nand U2151 (N_2151,In_657,In_603);
nand U2152 (N_2152,In_306,In_3);
and U2153 (N_2153,In_740,In_746);
xnor U2154 (N_2154,In_682,In_329);
nand U2155 (N_2155,In_615,In_330);
nand U2156 (N_2156,In_280,In_5);
and U2157 (N_2157,In_381,In_543);
nand U2158 (N_2158,In_446,In_582);
nand U2159 (N_2159,In_580,In_543);
and U2160 (N_2160,In_29,In_660);
nand U2161 (N_2161,In_387,In_556);
and U2162 (N_2162,In_403,In_452);
and U2163 (N_2163,In_594,In_166);
nand U2164 (N_2164,In_358,In_291);
nor U2165 (N_2165,In_27,In_322);
nand U2166 (N_2166,In_26,In_703);
nand U2167 (N_2167,In_88,In_397);
and U2168 (N_2168,In_424,In_616);
and U2169 (N_2169,In_376,In_377);
nand U2170 (N_2170,In_470,In_280);
nand U2171 (N_2171,In_590,In_534);
and U2172 (N_2172,In_236,In_741);
nand U2173 (N_2173,In_739,In_629);
or U2174 (N_2174,In_205,In_475);
nand U2175 (N_2175,In_310,In_524);
xor U2176 (N_2176,In_67,In_584);
nand U2177 (N_2177,In_19,In_468);
nand U2178 (N_2178,In_431,In_306);
or U2179 (N_2179,In_23,In_111);
xnor U2180 (N_2180,In_181,In_277);
and U2181 (N_2181,In_425,In_208);
nor U2182 (N_2182,In_546,In_363);
and U2183 (N_2183,In_92,In_146);
nor U2184 (N_2184,In_585,In_233);
and U2185 (N_2185,In_618,In_616);
nor U2186 (N_2186,In_505,In_382);
nor U2187 (N_2187,In_694,In_657);
and U2188 (N_2188,In_565,In_391);
and U2189 (N_2189,In_492,In_499);
or U2190 (N_2190,In_83,In_124);
or U2191 (N_2191,In_60,In_167);
nand U2192 (N_2192,In_660,In_378);
and U2193 (N_2193,In_572,In_686);
and U2194 (N_2194,In_16,In_14);
or U2195 (N_2195,In_562,In_312);
nor U2196 (N_2196,In_62,In_413);
xnor U2197 (N_2197,In_11,In_297);
nor U2198 (N_2198,In_274,In_656);
nand U2199 (N_2199,In_290,In_154);
and U2200 (N_2200,In_141,In_185);
or U2201 (N_2201,In_346,In_725);
or U2202 (N_2202,In_241,In_485);
or U2203 (N_2203,In_228,In_480);
or U2204 (N_2204,In_410,In_596);
or U2205 (N_2205,In_189,In_518);
nand U2206 (N_2206,In_504,In_395);
nand U2207 (N_2207,In_294,In_76);
nand U2208 (N_2208,In_363,In_181);
nor U2209 (N_2209,In_588,In_644);
nor U2210 (N_2210,In_399,In_185);
and U2211 (N_2211,In_245,In_31);
and U2212 (N_2212,In_335,In_550);
nand U2213 (N_2213,In_347,In_162);
nand U2214 (N_2214,In_112,In_230);
nand U2215 (N_2215,In_648,In_287);
and U2216 (N_2216,In_144,In_5);
or U2217 (N_2217,In_479,In_737);
xnor U2218 (N_2218,In_599,In_395);
nand U2219 (N_2219,In_31,In_360);
and U2220 (N_2220,In_269,In_536);
nor U2221 (N_2221,In_137,In_643);
nor U2222 (N_2222,In_662,In_438);
nor U2223 (N_2223,In_109,In_144);
or U2224 (N_2224,In_310,In_662);
nand U2225 (N_2225,In_234,In_322);
or U2226 (N_2226,In_736,In_548);
and U2227 (N_2227,In_733,In_24);
nand U2228 (N_2228,In_307,In_152);
and U2229 (N_2229,In_114,In_691);
nor U2230 (N_2230,In_504,In_365);
nor U2231 (N_2231,In_698,In_529);
nand U2232 (N_2232,In_132,In_445);
or U2233 (N_2233,In_485,In_330);
and U2234 (N_2234,In_659,In_683);
or U2235 (N_2235,In_108,In_120);
nor U2236 (N_2236,In_222,In_686);
nand U2237 (N_2237,In_255,In_217);
xor U2238 (N_2238,In_700,In_678);
or U2239 (N_2239,In_443,In_13);
or U2240 (N_2240,In_79,In_541);
nor U2241 (N_2241,In_248,In_745);
nand U2242 (N_2242,In_543,In_592);
nand U2243 (N_2243,In_263,In_294);
and U2244 (N_2244,In_715,In_178);
nand U2245 (N_2245,In_237,In_71);
and U2246 (N_2246,In_618,In_466);
and U2247 (N_2247,In_244,In_230);
nand U2248 (N_2248,In_663,In_392);
or U2249 (N_2249,In_372,In_245);
nor U2250 (N_2250,In_206,In_602);
nor U2251 (N_2251,In_631,In_409);
nand U2252 (N_2252,In_6,In_359);
nand U2253 (N_2253,In_683,In_89);
nor U2254 (N_2254,In_698,In_157);
nand U2255 (N_2255,In_579,In_716);
or U2256 (N_2256,In_394,In_440);
nor U2257 (N_2257,In_523,In_68);
or U2258 (N_2258,In_1,In_676);
and U2259 (N_2259,In_611,In_359);
or U2260 (N_2260,In_120,In_96);
and U2261 (N_2261,In_356,In_230);
nand U2262 (N_2262,In_358,In_310);
nand U2263 (N_2263,In_559,In_244);
nor U2264 (N_2264,In_489,In_589);
or U2265 (N_2265,In_730,In_554);
or U2266 (N_2266,In_306,In_623);
or U2267 (N_2267,In_727,In_137);
nand U2268 (N_2268,In_603,In_395);
nor U2269 (N_2269,In_282,In_600);
nand U2270 (N_2270,In_506,In_567);
nor U2271 (N_2271,In_84,In_711);
nor U2272 (N_2272,In_43,In_416);
nor U2273 (N_2273,In_549,In_46);
or U2274 (N_2274,In_63,In_542);
nand U2275 (N_2275,In_54,In_157);
nor U2276 (N_2276,In_733,In_592);
or U2277 (N_2277,In_51,In_723);
nor U2278 (N_2278,In_123,In_636);
nand U2279 (N_2279,In_87,In_19);
nor U2280 (N_2280,In_710,In_516);
and U2281 (N_2281,In_127,In_276);
and U2282 (N_2282,In_256,In_705);
nand U2283 (N_2283,In_102,In_125);
or U2284 (N_2284,In_421,In_26);
xnor U2285 (N_2285,In_581,In_471);
nand U2286 (N_2286,In_537,In_719);
nor U2287 (N_2287,In_587,In_179);
or U2288 (N_2288,In_122,In_67);
or U2289 (N_2289,In_86,In_155);
nand U2290 (N_2290,In_497,In_11);
or U2291 (N_2291,In_486,In_272);
nor U2292 (N_2292,In_243,In_266);
nand U2293 (N_2293,In_658,In_535);
or U2294 (N_2294,In_518,In_114);
or U2295 (N_2295,In_17,In_613);
or U2296 (N_2296,In_442,In_187);
nor U2297 (N_2297,In_128,In_646);
nor U2298 (N_2298,In_342,In_27);
and U2299 (N_2299,In_558,In_95);
and U2300 (N_2300,In_550,In_469);
nor U2301 (N_2301,In_242,In_550);
nor U2302 (N_2302,In_432,In_638);
nor U2303 (N_2303,In_326,In_282);
or U2304 (N_2304,In_473,In_327);
nor U2305 (N_2305,In_84,In_276);
nor U2306 (N_2306,In_399,In_536);
nand U2307 (N_2307,In_711,In_145);
or U2308 (N_2308,In_155,In_716);
nor U2309 (N_2309,In_131,In_527);
nor U2310 (N_2310,In_709,In_17);
and U2311 (N_2311,In_677,In_318);
nand U2312 (N_2312,In_711,In_510);
and U2313 (N_2313,In_563,In_619);
or U2314 (N_2314,In_187,In_89);
nand U2315 (N_2315,In_343,In_679);
nand U2316 (N_2316,In_344,In_595);
or U2317 (N_2317,In_222,In_264);
or U2318 (N_2318,In_506,In_193);
nor U2319 (N_2319,In_347,In_732);
nand U2320 (N_2320,In_302,In_684);
nand U2321 (N_2321,In_288,In_110);
or U2322 (N_2322,In_623,In_550);
nor U2323 (N_2323,In_397,In_521);
and U2324 (N_2324,In_94,In_146);
nor U2325 (N_2325,In_76,In_201);
or U2326 (N_2326,In_38,In_217);
and U2327 (N_2327,In_219,In_207);
nand U2328 (N_2328,In_674,In_87);
nor U2329 (N_2329,In_19,In_306);
nand U2330 (N_2330,In_395,In_746);
nand U2331 (N_2331,In_329,In_633);
nor U2332 (N_2332,In_528,In_710);
or U2333 (N_2333,In_428,In_399);
nand U2334 (N_2334,In_63,In_700);
and U2335 (N_2335,In_648,In_725);
nor U2336 (N_2336,In_28,In_248);
and U2337 (N_2337,In_236,In_140);
nor U2338 (N_2338,In_188,In_422);
or U2339 (N_2339,In_472,In_34);
nor U2340 (N_2340,In_370,In_32);
and U2341 (N_2341,In_137,In_744);
and U2342 (N_2342,In_739,In_310);
nor U2343 (N_2343,In_296,In_470);
or U2344 (N_2344,In_286,In_358);
nor U2345 (N_2345,In_235,In_303);
nand U2346 (N_2346,In_389,In_657);
nor U2347 (N_2347,In_701,In_213);
or U2348 (N_2348,In_278,In_526);
nor U2349 (N_2349,In_60,In_634);
or U2350 (N_2350,In_351,In_309);
nor U2351 (N_2351,In_246,In_384);
or U2352 (N_2352,In_456,In_626);
nand U2353 (N_2353,In_570,In_49);
nand U2354 (N_2354,In_626,In_35);
or U2355 (N_2355,In_514,In_30);
nand U2356 (N_2356,In_64,In_487);
or U2357 (N_2357,In_153,In_218);
nand U2358 (N_2358,In_605,In_388);
and U2359 (N_2359,In_284,In_47);
and U2360 (N_2360,In_39,In_593);
nor U2361 (N_2361,In_45,In_546);
nor U2362 (N_2362,In_259,In_263);
or U2363 (N_2363,In_737,In_163);
or U2364 (N_2364,In_386,In_602);
nand U2365 (N_2365,In_711,In_413);
and U2366 (N_2366,In_588,In_579);
nand U2367 (N_2367,In_261,In_42);
and U2368 (N_2368,In_403,In_93);
nand U2369 (N_2369,In_560,In_154);
or U2370 (N_2370,In_108,In_428);
nor U2371 (N_2371,In_371,In_124);
or U2372 (N_2372,In_272,In_573);
or U2373 (N_2373,In_718,In_656);
and U2374 (N_2374,In_566,In_609);
nand U2375 (N_2375,In_199,In_272);
nor U2376 (N_2376,In_56,In_130);
and U2377 (N_2377,In_100,In_88);
and U2378 (N_2378,In_554,In_545);
and U2379 (N_2379,In_636,In_585);
and U2380 (N_2380,In_414,In_357);
and U2381 (N_2381,In_521,In_652);
and U2382 (N_2382,In_504,In_418);
and U2383 (N_2383,In_704,In_585);
or U2384 (N_2384,In_25,In_575);
and U2385 (N_2385,In_665,In_678);
nor U2386 (N_2386,In_606,In_553);
or U2387 (N_2387,In_444,In_539);
and U2388 (N_2388,In_54,In_566);
and U2389 (N_2389,In_239,In_653);
or U2390 (N_2390,In_436,In_689);
or U2391 (N_2391,In_88,In_164);
nor U2392 (N_2392,In_417,In_718);
nand U2393 (N_2393,In_529,In_727);
nor U2394 (N_2394,In_524,In_729);
or U2395 (N_2395,In_681,In_530);
and U2396 (N_2396,In_643,In_710);
or U2397 (N_2397,In_166,In_329);
nor U2398 (N_2398,In_585,In_106);
and U2399 (N_2399,In_59,In_98);
and U2400 (N_2400,In_584,In_446);
nor U2401 (N_2401,In_639,In_32);
nand U2402 (N_2402,In_494,In_218);
nand U2403 (N_2403,In_616,In_418);
or U2404 (N_2404,In_434,In_457);
and U2405 (N_2405,In_585,In_153);
or U2406 (N_2406,In_219,In_152);
nand U2407 (N_2407,In_673,In_175);
nand U2408 (N_2408,In_736,In_403);
or U2409 (N_2409,In_460,In_79);
and U2410 (N_2410,In_367,In_65);
nand U2411 (N_2411,In_400,In_628);
and U2412 (N_2412,In_159,In_415);
nor U2413 (N_2413,In_745,In_557);
nor U2414 (N_2414,In_727,In_67);
nor U2415 (N_2415,In_68,In_52);
and U2416 (N_2416,In_696,In_295);
and U2417 (N_2417,In_458,In_739);
and U2418 (N_2418,In_625,In_359);
nand U2419 (N_2419,In_84,In_595);
or U2420 (N_2420,In_418,In_438);
and U2421 (N_2421,In_259,In_156);
and U2422 (N_2422,In_319,In_555);
nand U2423 (N_2423,In_84,In_334);
nand U2424 (N_2424,In_505,In_19);
nor U2425 (N_2425,In_333,In_49);
and U2426 (N_2426,In_282,In_336);
and U2427 (N_2427,In_499,In_391);
or U2428 (N_2428,In_291,In_467);
and U2429 (N_2429,In_168,In_666);
and U2430 (N_2430,In_275,In_59);
or U2431 (N_2431,In_727,In_147);
and U2432 (N_2432,In_81,In_342);
or U2433 (N_2433,In_740,In_111);
xnor U2434 (N_2434,In_274,In_502);
nor U2435 (N_2435,In_284,In_613);
nand U2436 (N_2436,In_478,In_498);
nand U2437 (N_2437,In_721,In_89);
nand U2438 (N_2438,In_229,In_537);
nor U2439 (N_2439,In_220,In_324);
nor U2440 (N_2440,In_199,In_568);
nand U2441 (N_2441,In_2,In_93);
nor U2442 (N_2442,In_482,In_259);
nand U2443 (N_2443,In_162,In_577);
and U2444 (N_2444,In_153,In_79);
or U2445 (N_2445,In_501,In_723);
nand U2446 (N_2446,In_417,In_572);
and U2447 (N_2447,In_361,In_195);
and U2448 (N_2448,In_394,In_50);
nand U2449 (N_2449,In_627,In_705);
nand U2450 (N_2450,In_705,In_338);
nand U2451 (N_2451,In_355,In_275);
nor U2452 (N_2452,In_177,In_165);
nand U2453 (N_2453,In_744,In_461);
or U2454 (N_2454,In_639,In_117);
or U2455 (N_2455,In_35,In_715);
nand U2456 (N_2456,In_374,In_541);
or U2457 (N_2457,In_35,In_509);
nand U2458 (N_2458,In_422,In_574);
or U2459 (N_2459,In_343,In_133);
nand U2460 (N_2460,In_151,In_671);
nand U2461 (N_2461,In_69,In_685);
or U2462 (N_2462,In_347,In_565);
nor U2463 (N_2463,In_470,In_417);
or U2464 (N_2464,In_620,In_644);
or U2465 (N_2465,In_205,In_306);
and U2466 (N_2466,In_275,In_96);
nor U2467 (N_2467,In_218,In_395);
nor U2468 (N_2468,In_447,In_368);
and U2469 (N_2469,In_111,In_605);
or U2470 (N_2470,In_277,In_228);
or U2471 (N_2471,In_608,In_332);
nor U2472 (N_2472,In_703,In_282);
and U2473 (N_2473,In_687,In_540);
or U2474 (N_2474,In_688,In_308);
nand U2475 (N_2475,In_364,In_4);
nand U2476 (N_2476,In_547,In_470);
and U2477 (N_2477,In_625,In_15);
or U2478 (N_2478,In_409,In_638);
nor U2479 (N_2479,In_306,In_156);
and U2480 (N_2480,In_611,In_399);
or U2481 (N_2481,In_401,In_612);
nand U2482 (N_2482,In_342,In_635);
or U2483 (N_2483,In_300,In_535);
or U2484 (N_2484,In_449,In_659);
nand U2485 (N_2485,In_527,In_366);
or U2486 (N_2486,In_227,In_188);
nor U2487 (N_2487,In_27,In_422);
nand U2488 (N_2488,In_481,In_506);
nand U2489 (N_2489,In_92,In_538);
or U2490 (N_2490,In_0,In_36);
and U2491 (N_2491,In_198,In_340);
or U2492 (N_2492,In_342,In_550);
nand U2493 (N_2493,In_454,In_324);
nor U2494 (N_2494,In_573,In_210);
and U2495 (N_2495,In_297,In_35);
nor U2496 (N_2496,In_352,In_442);
nand U2497 (N_2497,In_608,In_203);
nor U2498 (N_2498,In_238,In_360);
nor U2499 (N_2499,In_204,In_640);
or U2500 (N_2500,N_1223,N_1661);
and U2501 (N_2501,N_1444,N_1876);
or U2502 (N_2502,N_915,N_1492);
nand U2503 (N_2503,N_164,N_423);
and U2504 (N_2504,N_846,N_2198);
and U2505 (N_2505,N_1720,N_820);
nor U2506 (N_2506,N_1739,N_1451);
and U2507 (N_2507,N_2140,N_2155);
nor U2508 (N_2508,N_1425,N_2469);
or U2509 (N_2509,N_286,N_1855);
and U2510 (N_2510,N_1367,N_722);
nand U2511 (N_2511,N_141,N_359);
nor U2512 (N_2512,N_1788,N_1636);
nor U2513 (N_2513,N_1973,N_882);
or U2514 (N_2514,N_475,N_1795);
nand U2515 (N_2515,N_694,N_1481);
nand U2516 (N_2516,N_416,N_100);
nor U2517 (N_2517,N_2247,N_59);
nand U2518 (N_2518,N_218,N_2129);
nor U2519 (N_2519,N_1462,N_1774);
nor U2520 (N_2520,N_393,N_1963);
nand U2521 (N_2521,N_858,N_1067);
nor U2522 (N_2522,N_1009,N_2402);
and U2523 (N_2523,N_2318,N_58);
and U2524 (N_2524,N_1113,N_881);
nand U2525 (N_2525,N_1276,N_780);
nor U2526 (N_2526,N_352,N_388);
nand U2527 (N_2527,N_1230,N_1170);
or U2528 (N_2528,N_746,N_736);
and U2529 (N_2529,N_2072,N_829);
and U2530 (N_2530,N_1472,N_664);
and U2531 (N_2531,N_1868,N_436);
or U2532 (N_2532,N_1259,N_1524);
or U2533 (N_2533,N_248,N_1532);
or U2534 (N_2534,N_1769,N_252);
nor U2535 (N_2535,N_1742,N_815);
nor U2536 (N_2536,N_382,N_2310);
or U2537 (N_2537,N_1378,N_866);
nor U2538 (N_2538,N_1380,N_1646);
nor U2539 (N_2539,N_126,N_2455);
and U2540 (N_2540,N_823,N_1180);
or U2541 (N_2541,N_1995,N_2428);
and U2542 (N_2542,N_275,N_153);
nand U2543 (N_2543,N_1349,N_1423);
or U2544 (N_2544,N_266,N_1944);
nand U2545 (N_2545,N_1179,N_1333);
nand U2546 (N_2546,N_943,N_1169);
or U2547 (N_2547,N_2438,N_1517);
or U2548 (N_2548,N_1885,N_678);
and U2549 (N_2549,N_464,N_2342);
or U2550 (N_2550,N_1011,N_1718);
nand U2551 (N_2551,N_1657,N_1796);
nand U2552 (N_2552,N_1910,N_539);
xor U2553 (N_2553,N_2101,N_1779);
nor U2554 (N_2554,N_2341,N_327);
and U2555 (N_2555,N_1324,N_2167);
or U2556 (N_2556,N_1870,N_910);
nand U2557 (N_2557,N_263,N_917);
nor U2558 (N_2558,N_291,N_190);
nor U2559 (N_2559,N_732,N_4);
and U2560 (N_2560,N_101,N_1415);
or U2561 (N_2561,N_466,N_1049);
nor U2562 (N_2562,N_1695,N_1807);
nand U2563 (N_2563,N_1411,N_685);
or U2564 (N_2564,N_1780,N_482);
nor U2565 (N_2565,N_261,N_824);
and U2566 (N_2566,N_1212,N_353);
and U2567 (N_2567,N_2281,N_92);
or U2568 (N_2568,N_2163,N_609);
nor U2569 (N_2569,N_575,N_103);
nor U2570 (N_2570,N_634,N_524);
and U2571 (N_2571,N_2093,N_1773);
or U2572 (N_2572,N_2000,N_794);
nor U2573 (N_2573,N_508,N_1933);
and U2574 (N_2574,N_2189,N_1204);
and U2575 (N_2575,N_1967,N_874);
nor U2576 (N_2576,N_2203,N_90);
nand U2577 (N_2577,N_695,N_401);
nor U2578 (N_2578,N_1575,N_1390);
nand U2579 (N_2579,N_203,N_2109);
nand U2580 (N_2580,N_502,N_260);
nor U2581 (N_2581,N_1032,N_513);
and U2582 (N_2582,N_931,N_2490);
and U2583 (N_2583,N_1016,N_223);
nand U2584 (N_2584,N_2122,N_1790);
or U2585 (N_2585,N_648,N_813);
nor U2586 (N_2586,N_380,N_1108);
nor U2587 (N_2587,N_119,N_2498);
and U2588 (N_2588,N_1635,N_152);
or U2589 (N_2589,N_2021,N_1177);
nor U2590 (N_2590,N_1762,N_435);
and U2591 (N_2591,N_125,N_1019);
or U2592 (N_2592,N_1231,N_2376);
nor U2593 (N_2593,N_1610,N_178);
and U2594 (N_2594,N_1520,N_2314);
nor U2595 (N_2595,N_392,N_2266);
or U2596 (N_2596,N_1494,N_472);
and U2597 (N_2597,N_2124,N_939);
or U2598 (N_2598,N_1641,N_467);
and U2599 (N_2599,N_1474,N_1082);
nor U2600 (N_2600,N_967,N_1766);
nor U2601 (N_2601,N_1201,N_356);
and U2602 (N_2602,N_1012,N_364);
nor U2603 (N_2603,N_1961,N_2221);
or U2604 (N_2604,N_377,N_1529);
nand U2605 (N_2605,N_641,N_657);
and U2606 (N_2606,N_135,N_2042);
nand U2607 (N_2607,N_1284,N_1457);
nand U2608 (N_2608,N_188,N_2054);
nor U2609 (N_2609,N_1097,N_316);
and U2610 (N_2610,N_1731,N_398);
or U2611 (N_2611,N_287,N_2244);
nand U2612 (N_2612,N_1225,N_1136);
or U2613 (N_2613,N_1730,N_1332);
or U2614 (N_2614,N_509,N_895);
or U2615 (N_2615,N_268,N_2135);
or U2616 (N_2616,N_1834,N_2444);
nor U2617 (N_2617,N_1364,N_1063);
nand U2618 (N_2618,N_1543,N_439);
nand U2619 (N_2619,N_237,N_1841);
nor U2620 (N_2620,N_720,N_294);
and U2621 (N_2621,N_2009,N_2197);
or U2622 (N_2622,N_2174,N_592);
nor U2623 (N_2623,N_1768,N_702);
or U2624 (N_2624,N_578,N_432);
and U2625 (N_2625,N_2195,N_876);
or U2626 (N_2626,N_919,N_142);
or U2627 (N_2627,N_2278,N_1775);
nand U2628 (N_2628,N_1793,N_1533);
nor U2629 (N_2629,N_1835,N_474);
nand U2630 (N_2630,N_2029,N_308);
nor U2631 (N_2631,N_41,N_1343);
nand U2632 (N_2632,N_971,N_2141);
and U2633 (N_2633,N_45,N_434);
or U2634 (N_2634,N_2220,N_224);
nand U2635 (N_2635,N_2487,N_2245);
and U2636 (N_2636,N_1289,N_792);
or U2637 (N_2637,N_2262,N_1881);
and U2638 (N_2638,N_229,N_1250);
nor U2639 (N_2639,N_144,N_2338);
or U2640 (N_2640,N_1190,N_671);
nand U2641 (N_2641,N_1427,N_27);
and U2642 (N_2642,N_1662,N_1613);
and U2643 (N_2643,N_450,N_1549);
nand U2644 (N_2644,N_496,N_1561);
nand U2645 (N_2645,N_108,N_104);
and U2646 (N_2646,N_1936,N_2260);
nand U2647 (N_2647,N_2363,N_1865);
nand U2648 (N_2648,N_2156,N_580);
nor U2649 (N_2649,N_719,N_31);
xnor U2650 (N_2650,N_1687,N_2105);
and U2651 (N_2651,N_236,N_894);
nor U2652 (N_2652,N_1857,N_53);
and U2653 (N_2653,N_1597,N_673);
nor U2654 (N_2654,N_1329,N_511);
nand U2655 (N_2655,N_369,N_1569);
nand U2656 (N_2656,N_298,N_1678);
nand U2657 (N_2657,N_730,N_2465);
or U2658 (N_2658,N_447,N_24);
nor U2659 (N_2659,N_1106,N_1574);
and U2660 (N_2660,N_1948,N_683);
nand U2661 (N_2661,N_817,N_1041);
and U2662 (N_2662,N_449,N_756);
or U2663 (N_2663,N_389,N_568);
or U2664 (N_2664,N_2417,N_211);
or U2665 (N_2665,N_1907,N_777);
or U2666 (N_2666,N_184,N_35);
or U2667 (N_2667,N_1939,N_1402);
nand U2668 (N_2668,N_1658,N_2132);
nor U2669 (N_2669,N_1874,N_202);
and U2670 (N_2670,N_906,N_723);
nand U2671 (N_2671,N_1737,N_1847);
or U2672 (N_2672,N_699,N_1510);
and U2673 (N_2673,N_1837,N_787);
nor U2674 (N_2674,N_1003,N_834);
nor U2675 (N_2675,N_1157,N_1698);
and U2676 (N_2676,N_2261,N_504);
or U2677 (N_2677,N_2251,N_2048);
and U2678 (N_2678,N_738,N_1091);
nand U2679 (N_2679,N_1580,N_1585);
or U2680 (N_2680,N_216,N_519);
and U2681 (N_2681,N_577,N_1502);
and U2682 (N_2682,N_1304,N_1232);
nor U2683 (N_2683,N_681,N_2110);
or U2684 (N_2684,N_2304,N_1386);
nand U2685 (N_2685,N_2039,N_1290);
and U2686 (N_2686,N_923,N_1077);
nor U2687 (N_2687,N_1498,N_1830);
nand U2688 (N_2688,N_2431,N_282);
and U2689 (N_2689,N_1042,N_847);
or U2690 (N_2690,N_2329,N_1781);
nor U2691 (N_2691,N_1361,N_930);
and U2692 (N_2692,N_2117,N_2252);
or U2693 (N_2693,N_760,N_909);
nor U2694 (N_2694,N_1866,N_1392);
and U2695 (N_2695,N_620,N_1601);
and U2696 (N_2696,N_330,N_541);
and U2697 (N_2697,N_1383,N_182);
nand U2698 (N_2698,N_1149,N_650);
and U2699 (N_2699,N_1447,N_2120);
and U2700 (N_2700,N_1879,N_570);
and U2701 (N_2701,N_2420,N_507);
or U2702 (N_2702,N_2295,N_1104);
or U2703 (N_2703,N_373,N_400);
or U2704 (N_2704,N_1897,N_1856);
nor U2705 (N_2705,N_1776,N_959);
nor U2706 (N_2706,N_1515,N_1193);
nor U2707 (N_2707,N_1142,N_2183);
nor U2708 (N_2708,N_877,N_1504);
and U2709 (N_2709,N_2185,N_505);
and U2710 (N_2710,N_2446,N_2179);
and U2711 (N_2711,N_765,N_336);
nor U2712 (N_2712,N_148,N_1439);
nand U2713 (N_2713,N_1287,N_2415);
and U2714 (N_2714,N_234,N_1821);
nand U2715 (N_2715,N_49,N_527);
nand U2716 (N_2716,N_1320,N_2291);
or U2717 (N_2717,N_825,N_227);
nand U2718 (N_2718,N_1094,N_1213);
nand U2719 (N_2719,N_2225,N_1293);
or U2720 (N_2720,N_2300,N_515);
nor U2721 (N_2721,N_2254,N_1185);
nor U2722 (N_2722,N_833,N_415);
and U2723 (N_2723,N_2335,N_1203);
or U2724 (N_2724,N_2361,N_973);
nor U2725 (N_2725,N_1851,N_828);
and U2726 (N_2726,N_841,N_448);
and U2727 (N_2727,N_1676,N_879);
nor U2728 (N_2728,N_566,N_2137);
and U2729 (N_2729,N_2373,N_1126);
and U2730 (N_2730,N_168,N_347);
or U2731 (N_2731,N_2238,N_582);
or U2732 (N_2732,N_1491,N_471);
xnor U2733 (N_2733,N_1528,N_1556);
and U2734 (N_2734,N_399,N_1546);
nor U2735 (N_2735,N_456,N_1410);
nor U2736 (N_2736,N_129,N_95);
or U2737 (N_2737,N_921,N_2457);
nand U2738 (N_2738,N_1711,N_753);
nor U2739 (N_2739,N_2087,N_789);
nor U2740 (N_2740,N_2473,N_2035);
nor U2741 (N_2741,N_57,N_835);
and U2742 (N_2742,N_1810,N_19);
nor U2743 (N_2743,N_2068,N_731);
or U2744 (N_2744,N_1158,N_1634);
or U2745 (N_2745,N_2045,N_2234);
nand U2746 (N_2746,N_812,N_1323);
nor U2747 (N_2747,N_1633,N_257);
or U2748 (N_2748,N_2411,N_1120);
nand U2749 (N_2749,N_1396,N_1321);
xor U2750 (N_2750,N_413,N_1506);
or U2751 (N_2751,N_455,N_2052);
nor U2752 (N_2752,N_1909,N_2386);
nand U2753 (N_2753,N_2424,N_918);
nand U2754 (N_2754,N_1139,N_2483);
nor U2755 (N_2755,N_1838,N_600);
or U2756 (N_2756,N_1134,N_265);
and U2757 (N_2757,N_1466,N_395);
or U2758 (N_2758,N_2050,N_2392);
and U2759 (N_2759,N_2412,N_1461);
nor U2760 (N_2760,N_1391,N_936);
nand U2761 (N_2761,N_1668,N_995);
or U2762 (N_2762,N_637,N_561);
nor U2763 (N_2763,N_1589,N_2006);
or U2764 (N_2764,N_138,N_1014);
or U2765 (N_2765,N_1351,N_201);
nor U2766 (N_2766,N_2294,N_1235);
or U2767 (N_2767,N_659,N_17);
nor U2768 (N_2768,N_1872,N_2169);
or U2769 (N_2769,N_5,N_1432);
nor U2770 (N_2770,N_2100,N_1163);
nand U2771 (N_2771,N_2493,N_1783);
nand U2772 (N_2772,N_1708,N_1576);
or U2773 (N_2773,N_2089,N_1558);
nand U2774 (N_2774,N_441,N_2432);
and U2775 (N_2775,N_1602,N_420);
and U2776 (N_2776,N_2429,N_2389);
nor U2777 (N_2777,N_925,N_2257);
nor U2778 (N_2778,N_2485,N_486);
or U2779 (N_2779,N_1900,N_892);
nand U2780 (N_2780,N_891,N_2233);
or U2781 (N_2781,N_661,N_2463);
or U2782 (N_2782,N_2268,N_2401);
nor U2783 (N_2783,N_2046,N_529);
and U2784 (N_2784,N_1270,N_1412);
or U2785 (N_2785,N_2265,N_2382);
or U2786 (N_2786,N_215,N_2121);
nand U2787 (N_2787,N_1608,N_857);
and U2788 (N_2788,N_1105,N_603);
or U2789 (N_2789,N_868,N_2212);
nor U2790 (N_2790,N_2111,N_1281);
nand U2791 (N_2791,N_1189,N_636);
or U2792 (N_2792,N_1850,N_988);
and U2793 (N_2793,N_1819,N_7);
or U2794 (N_2794,N_797,N_1219);
and U2795 (N_2795,N_528,N_2482);
nand U2796 (N_2796,N_711,N_2336);
or U2797 (N_2797,N_2201,N_715);
or U2798 (N_2798,N_2014,N_1100);
nor U2799 (N_2799,N_1934,N_1224);
or U2800 (N_2800,N_2145,N_1171);
nor U2801 (N_2801,N_1080,N_1645);
and U2802 (N_2802,N_1034,N_983);
nor U2803 (N_2803,N_2370,N_1418);
and U2804 (N_2804,N_1369,N_2004);
or U2805 (N_2805,N_1467,N_1018);
nor U2806 (N_2806,N_1419,N_1651);
nor U2807 (N_2807,N_1000,N_2056);
xnor U2808 (N_2808,N_2194,N_2406);
or U2809 (N_2809,N_2041,N_288);
or U2810 (N_2810,N_1938,N_1717);
and U2811 (N_2811,N_2299,N_1022);
or U2812 (N_2812,N_734,N_2053);
nand U2813 (N_2813,N_1833,N_1437);
nand U2814 (N_2814,N_457,N_1184);
xnor U2815 (N_2815,N_1990,N_1187);
nand U2816 (N_2816,N_2285,N_1951);
nand U2817 (N_2817,N_771,N_91);
or U2818 (N_2818,N_642,N_2063);
or U2819 (N_2819,N_1751,N_1522);
nand U2820 (N_2820,N_150,N_665);
nor U2821 (N_2821,N_2393,N_446);
or U2822 (N_2822,N_1889,N_1846);
nor U2823 (N_2823,N_204,N_1802);
and U2824 (N_2824,N_1426,N_1195);
nor U2825 (N_2825,N_827,N_1537);
nor U2826 (N_2826,N_1536,N_157);
and U2827 (N_2827,N_1357,N_2377);
xor U2828 (N_2828,N_1697,N_2216);
nor U2829 (N_2829,N_1449,N_2139);
xor U2830 (N_2830,N_133,N_2489);
or U2831 (N_2831,N_2301,N_1355);
and U2832 (N_2832,N_1994,N_2467);
or U2833 (N_2833,N_821,N_2380);
and U2834 (N_2834,N_1860,N_1593);
nor U2835 (N_2835,N_721,N_186);
or U2836 (N_2836,N_1164,N_77);
nor U2837 (N_2837,N_344,N_493);
nor U2838 (N_2838,N_1372,N_226);
nand U2839 (N_2839,N_2351,N_1686);
or U2840 (N_2840,N_1424,N_1194);
nand U2841 (N_2841,N_1534,N_749);
nand U2842 (N_2842,N_2154,N_452);
nand U2843 (N_2843,N_1285,N_276);
nor U2844 (N_2844,N_300,N_1311);
and U2845 (N_2845,N_468,N_250);
nand U2846 (N_2846,N_385,N_2305);
and U2847 (N_2847,N_1538,N_1319);
and U2848 (N_2848,N_521,N_1214);
nor U2849 (N_2849,N_1121,N_2202);
nor U2850 (N_2850,N_1596,N_1976);
nor U2851 (N_2851,N_1409,N_1371);
nand U2852 (N_2852,N_1924,N_562);
and U2853 (N_2853,N_490,N_790);
nand U2854 (N_2854,N_1705,N_549);
or U2855 (N_2855,N_1625,N_501);
and U2856 (N_2856,N_590,N_1429);
nor U2857 (N_2857,N_759,N_796);
nand U2858 (N_2858,N_1572,N_1405);
and U2859 (N_2859,N_225,N_1197);
nand U2860 (N_2860,N_2086,N_1054);
and U2861 (N_2861,N_2456,N_2131);
nand U2862 (N_2862,N_1062,N_73);
or U2863 (N_2863,N_1283,N_412);
or U2864 (N_2864,N_1374,N_927);
or U2865 (N_2865,N_2325,N_2151);
and U2866 (N_2866,N_693,N_1297);
and U2867 (N_2867,N_1192,N_1033);
nor U2868 (N_2868,N_1594,N_955);
and U2869 (N_2869,N_1514,N_2475);
and U2870 (N_2870,N_2030,N_2027);
nor U2871 (N_2871,N_652,N_1068);
nand U2872 (N_2872,N_2462,N_938);
nor U2873 (N_2873,N_2001,N_1902);
or U2874 (N_2874,N_2492,N_1023);
nand U2875 (N_2875,N_323,N_2458);
nor U2876 (N_2876,N_2452,N_1854);
and U2877 (N_2877,N_705,N_680);
or U2878 (N_2878,N_2286,N_1366);
nand U2879 (N_2879,N_1053,N_1828);
and U2880 (N_2880,N_1825,N_376);
or U2881 (N_2881,N_2228,N_2011);
nand U2882 (N_2882,N_122,N_601);
nor U2883 (N_2883,N_1521,N_1044);
nor U2884 (N_2884,N_1935,N_1519);
and U2885 (N_2885,N_162,N_1562);
nand U2886 (N_2886,N_1791,N_1511);
nor U2887 (N_2887,N_72,N_2348);
and U2888 (N_2888,N_222,N_660);
and U2889 (N_2889,N_1770,N_1955);
nand U2890 (N_2890,N_2387,N_1986);
or U2891 (N_2891,N_633,N_84);
nor U2892 (N_2892,N_1478,N_1675);
nor U2893 (N_2893,N_1743,N_986);
nand U2894 (N_2894,N_1471,N_596);
nand U2895 (N_2895,N_1385,N_1918);
nand U2896 (N_2896,N_1677,N_818);
and U2897 (N_2897,N_361,N_2138);
nand U2898 (N_2898,N_2127,N_1926);
nor U2899 (N_2899,N_1591,N_1653);
and U2900 (N_2900,N_593,N_1020);
nor U2901 (N_2901,N_2084,N_8);
nand U2902 (N_2902,N_2430,N_905);
or U2903 (N_2903,N_1056,N_2359);
and U2904 (N_2904,N_343,N_1257);
nor U2905 (N_2905,N_1977,N_1128);
nor U2906 (N_2906,N_1923,N_552);
nand U2907 (N_2907,N_1709,N_889);
nor U2908 (N_2908,N_2479,N_1271);
nor U2909 (N_2909,N_1570,N_980);
nor U2910 (N_2910,N_2071,N_1337);
or U2911 (N_2911,N_1916,N_2184);
or U2912 (N_2912,N_484,N_1797);
and U2913 (N_2913,N_1229,N_349);
and U2914 (N_2914,N_755,N_1732);
nor U2915 (N_2915,N_213,N_2385);
and U2916 (N_2916,N_1119,N_1254);
and U2917 (N_2917,N_459,N_1959);
and U2918 (N_2918,N_709,N_1917);
and U2919 (N_2919,N_2017,N_1733);
nor U2920 (N_2920,N_581,N_2419);
or U2921 (N_2921,N_997,N_238);
or U2922 (N_2922,N_1239,N_458);
or U2923 (N_2923,N_1452,N_1244);
nor U2924 (N_2924,N_968,N_2047);
nor U2925 (N_2925,N_1740,N_1914);
nand U2926 (N_2926,N_1227,N_194);
nor U2927 (N_2927,N_16,N_279);
and U2928 (N_2928,N_2253,N_703);
nand U2929 (N_2929,N_1469,N_1503);
or U2930 (N_2930,N_741,N_219);
and U2931 (N_2931,N_791,N_1326);
and U2932 (N_2932,N_898,N_878);
nand U2933 (N_2933,N_2480,N_1037);
or U2934 (N_2934,N_560,N_757);
or U2935 (N_2935,N_411,N_1446);
or U2936 (N_2936,N_543,N_1359);
nor U2937 (N_2937,N_2319,N_1233);
or U2938 (N_2938,N_2049,N_599);
nor U2939 (N_2939,N_314,N_2024);
nor U2940 (N_2940,N_1688,N_217);
nor U2941 (N_2941,N_228,N_537);
or U2942 (N_2942,N_461,N_798);
nor U2943 (N_2943,N_1486,N_1665);
xnor U2944 (N_2944,N_1753,N_2303);
nor U2945 (N_2945,N_1960,N_1315);
nor U2946 (N_2946,N_2309,N_1871);
or U2947 (N_2947,N_161,N_1745);
and U2948 (N_2948,N_1508,N_500);
and U2949 (N_2949,N_1073,N_863);
and U2950 (N_2950,N_848,N_1084);
or U2951 (N_2951,N_1463,N_1911);
nand U2952 (N_2952,N_1714,N_56);
nor U2953 (N_2953,N_289,N_1399);
nand U2954 (N_2954,N_1761,N_2090);
and U2955 (N_2955,N_1109,N_2384);
nand U2956 (N_2956,N_900,N_1747);
nand U2957 (N_2957,N_1867,N_572);
and U2958 (N_2958,N_1612,N_2088);
and U2959 (N_2959,N_131,N_2075);
or U2960 (N_2960,N_1274,N_85);
nand U2961 (N_2961,N_2065,N_1729);
nand U2962 (N_2962,N_1925,N_1162);
and U2963 (N_2963,N_426,N_2269);
nand U2964 (N_2964,N_290,N_1669);
or U2965 (N_2965,N_497,N_644);
nor U2966 (N_2966,N_1767,N_859);
nand U2967 (N_2967,N_1309,N_530);
and U2968 (N_2968,N_1154,N_2400);
nand U2969 (N_2969,N_1495,N_1552);
or U2970 (N_2970,N_1667,N_1588);
or U2971 (N_2971,N_739,N_1518);
or U2972 (N_2972,N_1436,N_1308);
or U2973 (N_2973,N_1673,N_2275);
or U2974 (N_2974,N_2442,N_2057);
or U2975 (N_2975,N_536,N_10);
nor U2976 (N_2976,N_241,N_2150);
and U2977 (N_2977,N_1414,N_2488);
nor U2978 (N_2978,N_2322,N_811);
nor U2979 (N_2979,N_2157,N_123);
nand U2980 (N_2980,N_2153,N_1685);
nand U2981 (N_2981,N_1345,N_437);
nand U2982 (N_2982,N_2170,N_893);
nand U2983 (N_2983,N_107,N_1592);
and U2984 (N_2984,N_173,N_1978);
or U2985 (N_2985,N_1477,N_1307);
or U2986 (N_2986,N_1931,N_375);
or U2987 (N_2987,N_1252,N_2227);
or U2988 (N_2988,N_65,N_1347);
nor U2989 (N_2989,N_1291,N_1968);
nand U2990 (N_2990,N_591,N_2474);
or U2991 (N_2991,N_307,N_1942);
nand U2992 (N_2992,N_1674,N_1983);
and U2993 (N_2993,N_880,N_556);
and U2994 (N_2994,N_2059,N_1680);
and U2995 (N_2995,N_1937,N_1070);
and U2996 (N_2996,N_2378,N_18);
nor U2997 (N_2997,N_256,N_2128);
nand U2998 (N_2998,N_1175,N_2496);
nor U2999 (N_2999,N_158,N_476);
or U3000 (N_3000,N_1598,N_1778);
or U3001 (N_3001,N_1831,N_1215);
nand U3002 (N_3002,N_48,N_1406);
and U3003 (N_3003,N_302,N_1941);
and U3004 (N_3004,N_1306,N_1122);
nor U3005 (N_3005,N_311,N_1564);
and U3006 (N_3006,N_397,N_532);
nand U3007 (N_3007,N_1586,N_2007);
or U3008 (N_3008,N_2243,N_94);
and U3009 (N_3009,N_1131,N_935);
or U3010 (N_3010,N_1071,N_2395);
or U3011 (N_3011,N_506,N_1133);
and U3012 (N_3012,N_1784,N_235);
nor U3013 (N_3013,N_750,N_842);
and U3014 (N_3014,N_1387,N_576);
and U3015 (N_3015,N_2307,N_113);
or U3016 (N_3016,N_2199,N_831);
nand U3017 (N_3017,N_2437,N_1772);
nand U3018 (N_3018,N_1827,N_1027);
nor U3019 (N_3019,N_1389,N_1373);
nand U3020 (N_3020,N_838,N_1928);
or U3021 (N_3021,N_2413,N_405);
nor U3022 (N_3022,N_2160,N_1129);
and U3023 (N_3023,N_1736,N_629);
and U3024 (N_3024,N_74,N_1832);
or U3025 (N_3025,N_2346,N_2279);
and U3026 (N_3026,N_914,N_1824);
nand U3027 (N_3027,N_708,N_2312);
nor U3028 (N_3028,N_754,N_1932);
nor U3029 (N_3029,N_134,N_1039);
nand U3030 (N_3030,N_1339,N_2020);
nand U3031 (N_3031,N_1758,N_116);
nand U3032 (N_3032,N_2334,N_139);
and U3033 (N_3033,N_956,N_950);
or U3034 (N_3034,N_1905,N_643);
or U3035 (N_3035,N_1085,N_2186);
xnor U3036 (N_3036,N_573,N_806);
and U3037 (N_3037,N_1441,N_391);
or U3038 (N_3038,N_1222,N_503);
nand U3039 (N_3039,N_338,N_1701);
nand U3040 (N_3040,N_130,N_1573);
or U3041 (N_3041,N_1954,N_548);
or U3042 (N_3042,N_1176,N_998);
nand U3043 (N_3043,N_604,N_1985);
and U3044 (N_3044,N_1887,N_312);
nand U3045 (N_3045,N_735,N_1999);
or U3046 (N_3046,N_1899,N_2460);
and U3047 (N_3047,N_2345,N_804);
xnor U3048 (N_3048,N_803,N_247);
nand U3049 (N_3049,N_2073,N_1621);
and U3050 (N_3050,N_872,N_2226);
nand U3051 (N_3051,N_1453,N_1341);
or U3052 (N_3052,N_174,N_1246);
nand U3053 (N_3053,N_492,N_306);
or U3054 (N_3054,N_1280,N_903);
or U3055 (N_3055,N_2352,N_2107);
or U3056 (N_3056,N_1363,N_1305);
or U3057 (N_3057,N_1211,N_1420);
and U3058 (N_3058,N_1096,N_772);
nor U3059 (N_3059,N_773,N_554);
nand U3060 (N_3060,N_1117,N_2356);
xor U3061 (N_3061,N_800,N_2364);
or U3062 (N_3062,N_2394,N_1873);
nor U3063 (N_3063,N_1001,N_1663);
and U3064 (N_3064,N_105,N_309);
and U3065 (N_3065,N_481,N_2187);
or U3066 (N_3066,N_50,N_2478);
and U3067 (N_3067,N_1715,N_1947);
nor U3068 (N_3068,N_1482,N_1527);
xnor U3069 (N_3069,N_120,N_1431);
nor U3070 (N_3070,N_270,N_724);
and U3071 (N_3071,N_855,N_999);
or U3072 (N_3072,N_2369,N_2077);
and U3073 (N_3073,N_1880,N_1028);
or U3074 (N_3074,N_2449,N_292);
xor U3075 (N_3075,N_422,N_1883);
nor U3076 (N_3076,N_1058,N_167);
or U3077 (N_3077,N_691,N_1922);
nor U3078 (N_3078,N_1682,N_1125);
nor U3079 (N_3079,N_626,N_2350);
and U3080 (N_3080,N_1490,N_253);
or U3081 (N_3081,N_2083,N_1559);
nor U3082 (N_3082,N_2164,N_1236);
and U3083 (N_3083,N_2422,N_2302);
and U3084 (N_3084,N_1130,N_2263);
and U3085 (N_3085,N_1864,N_1272);
and U3086 (N_3086,N_55,N_1785);
or U3087 (N_3087,N_345,N_197);
or U3088 (N_3088,N_853,N_112);
or U3089 (N_3089,N_127,N_1792);
nor U3090 (N_3090,N_2255,N_654);
or U3091 (N_3091,N_1050,N_1587);
and U3092 (N_3092,N_1440,N_1505);
nand U3093 (N_3093,N_945,N_1583);
nor U3094 (N_3094,N_1801,N_1966);
nand U3095 (N_3095,N_2055,N_2218);
or U3096 (N_3096,N_408,N_1614);
or U3097 (N_3097,N_653,N_1135);
nand U3098 (N_3098,N_75,N_743);
and U3099 (N_3099,N_1724,N_1182);
nor U3100 (N_3100,N_1809,N_779);
nor U3101 (N_3101,N_179,N_890);
nand U3102 (N_3102,N_183,N_1310);
nand U3103 (N_3103,N_2242,N_2497);
nor U3104 (N_3104,N_1292,N_540);
and U3105 (N_3105,N_816,N_712);
nand U3106 (N_3106,N_1448,N_1550);
nand U3107 (N_3107,N_2108,N_922);
and U3108 (N_3108,N_1712,N_360);
nand U3109 (N_3109,N_2256,N_2371);
nor U3110 (N_3110,N_246,N_491);
and U3111 (N_3111,N_1408,N_278);
nand U3112 (N_3112,N_1859,N_299);
nor U3113 (N_3113,N_1974,N_2010);
or U3114 (N_3114,N_883,N_2470);
and U3115 (N_3115,N_2003,N_1813);
nand U3116 (N_3116,N_2330,N_1398);
or U3117 (N_3117,N_897,N_1799);
nor U3118 (N_3118,N_1262,N_960);
nand U3119 (N_3119,N_1862,N_1670);
nand U3120 (N_3120,N_2280,N_615);
nor U3121 (N_3121,N_1089,N_1590);
nor U3122 (N_3122,N_93,N_1719);
or U3123 (N_3123,N_1754,N_1464);
and U3124 (N_3124,N_2410,N_1208);
nand U3125 (N_3125,N_1107,N_1566);
or U3126 (N_3126,N_2028,N_1666);
or U3127 (N_3127,N_1487,N_295);
nor U3128 (N_3128,N_974,N_239);
or U3129 (N_3129,N_589,N_2188);
or U3130 (N_3130,N_2040,N_558);
and U3131 (N_3131,N_737,N_850);
nor U3132 (N_3132,N_498,N_1605);
or U3133 (N_3133,N_42,N_1760);
and U3134 (N_3134,N_1273,N_340);
nand U3135 (N_3135,N_2276,N_1264);
nor U3136 (N_3136,N_71,N_1765);
or U3137 (N_3137,N_1407,N_414);
nor U3138 (N_3138,N_362,N_1815);
nand U3139 (N_3139,N_386,N_2176);
and U3140 (N_3140,N_1734,N_928);
or U3141 (N_3141,N_2477,N_1888);
and U3142 (N_3142,N_2326,N_2142);
nand U3143 (N_3143,N_1322,N_1496);
nor U3144 (N_3144,N_208,N_1700);
nand U3145 (N_3145,N_975,N_370);
nor U3146 (N_3146,N_1604,N_649);
or U3147 (N_3147,N_1013,N_2388);
or U3148 (N_3148,N_1861,N_814);
nor U3149 (N_3149,N_1267,N_870);
and U3150 (N_3150,N_325,N_1806);
nand U3151 (N_3151,N_2207,N_443);
and U3152 (N_3152,N_1360,N_1087);
or U3153 (N_3153,N_1316,N_805);
nor U3154 (N_3154,N_1092,N_920);
nor U3155 (N_3155,N_1088,N_2096);
nor U3156 (N_3156,N_1168,N_713);
or U3157 (N_3157,N_2191,N_82);
nand U3158 (N_3158,N_1728,N_54);
nand U3159 (N_3159,N_1713,N_283);
or U3160 (N_3160,N_1615,N_667);
or U3161 (N_3161,N_209,N_1798);
nand U3162 (N_3162,N_111,N_836);
and U3163 (N_3163,N_1137,N_2208);
nor U3164 (N_3164,N_1563,N_579);
nor U3165 (N_3165,N_1863,N_1354);
nand U3166 (N_3166,N_2224,N_970);
nand U3167 (N_3167,N_1757,N_522);
or U3168 (N_3168,N_1997,N_145);
and U3169 (N_3169,N_143,N_2037);
nand U3170 (N_3170,N_869,N_1202);
or U3171 (N_3171,N_698,N_646);
and U3172 (N_3172,N_614,N_1913);
nand U3173 (N_3173,N_191,N_605);
or U3174 (N_3174,N_2230,N_2443);
and U3175 (N_3175,N_1927,N_1060);
and U3176 (N_3176,N_1206,N_1144);
nand U3177 (N_3177,N_1210,N_2130);
and U3178 (N_3178,N_2178,N_2425);
nand U3179 (N_3179,N_206,N_1186);
or U3180 (N_3180,N_1112,N_716);
and U3181 (N_3181,N_1702,N_329);
nor U3182 (N_3182,N_1268,N_1052);
or U3183 (N_3183,N_473,N_1632);
or U3184 (N_3184,N_2026,N_487);
nand U3185 (N_3185,N_433,N_2114);
and U3186 (N_3186,N_1970,N_602);
or U3187 (N_3187,N_1051,N_1413);
nand U3188 (N_3188,N_2283,N_1578);
and U3189 (N_3189,N_1660,N_2116);
and U3190 (N_3190,N_180,N_1965);
nand U3191 (N_3191,N_1624,N_583);
and U3192 (N_3192,N_1945,N_1637);
and U3193 (N_3193,N_799,N_2327);
nor U3194 (N_3194,N_2476,N_210);
and U3195 (N_3195,N_1340,N_953);
or U3196 (N_3196,N_1455,N_1400);
or U3197 (N_3197,N_1764,N_832);
nor U3198 (N_3198,N_1081,N_2019);
nand U3199 (N_3199,N_2403,N_1771);
nor U3200 (N_3200,N_1890,N_2204);
or U3201 (N_3201,N_63,N_2067);
or U3202 (N_3202,N_106,N_2229);
nand U3203 (N_3203,N_726,N_2158);
nand U3204 (N_3204,N_1099,N_1577);
or U3205 (N_3205,N_199,N_1330);
nor U3206 (N_3206,N_1288,N_2092);
or U3207 (N_3207,N_1852,N_1629);
and U3208 (N_3208,N_1836,N_2134);
nor U3209 (N_3209,N_1381,N_1755);
and U3210 (N_3210,N_704,N_1523);
nor U3211 (N_3211,N_1275,N_46);
and U3212 (N_3212,N_1979,N_1548);
nand U3213 (N_3213,N_1786,N_1816);
nor U3214 (N_3214,N_419,N_1489);
or U3215 (N_3215,N_2249,N_97);
nor U3216 (N_3216,N_1110,N_1393);
and U3217 (N_3217,N_1048,N_1443);
and U3218 (N_3218,N_214,N_1035);
nand U3219 (N_3219,N_2317,N_1992);
nor U3220 (N_3220,N_200,N_1286);
and U3221 (N_3221,N_1539,N_1350);
and U3222 (N_3222,N_2396,N_465);
nor U3223 (N_3223,N_977,N_2115);
and U3224 (N_3224,N_957,N_1299);
nand U3225 (N_3225,N_245,N_1445);
and U3226 (N_3226,N_864,N_1005);
and U3227 (N_3227,N_1582,N_304);
nand U3228 (N_3228,N_1545,N_1691);
nor U3229 (N_3229,N_371,N_1312);
nor U3230 (N_3230,N_2205,N_319);
nor U3231 (N_3231,N_355,N_994);
or U3232 (N_3232,N_402,N_1652);
nor U3233 (N_3233,N_2287,N_884);
or U3234 (N_3234,N_1706,N_1627);
or U3235 (N_3235,N_783,N_47);
or U3236 (N_3236,N_137,N_852);
nand U3237 (N_3237,N_2315,N_2357);
or U3238 (N_3238,N_1896,N_1093);
or U3239 (N_3239,N_326,N_383);
or U3240 (N_3240,N_1971,N_2106);
nor U3241 (N_3241,N_1998,N_1483);
or U3242 (N_3242,N_1683,N_745);
or U3243 (N_3243,N_952,N_840);
nor U3244 (N_3244,N_28,N_61);
nand U3245 (N_3245,N_390,N_366);
or U3246 (N_3246,N_916,N_2078);
nand U3247 (N_3247,N_469,N_1173);
and U3248 (N_3248,N_2213,N_744);
and U3249 (N_3249,N_1581,N_1912);
or U3250 (N_3250,N_2239,N_849);
and U3251 (N_3251,N_451,N_993);
nand U3252 (N_3252,N_1226,N_845);
or U3253 (N_3253,N_368,N_2450);
and U3254 (N_3254,N_2277,N_20);
nor U3255 (N_3255,N_1026,N_1102);
and U3256 (N_3256,N_1124,N_801);
and U3257 (N_3257,N_689,N_379);
or U3258 (N_3258,N_151,N_2259);
and U3259 (N_3259,N_494,N_1622);
nand U3260 (N_3260,N_60,N_616);
nor U3261 (N_3261,N_2397,N_1220);
nand U3262 (N_3262,N_163,N_632);
nor U3263 (N_3263,N_1241,N_969);
and U3264 (N_3264,N_1207,N_1148);
and U3265 (N_3265,N_546,N_69);
or U3266 (N_3266,N_154,N_2264);
nand U3267 (N_3267,N_822,N_885);
or U3268 (N_3268,N_1485,N_1165);
nor U3269 (N_3269,N_2102,N_2036);
or U3270 (N_3270,N_463,N_189);
or U3271 (N_3271,N_1095,N_2288);
nor U3272 (N_3272,N_1726,N_372);
and U3273 (N_3273,N_989,N_784);
or U3274 (N_3274,N_608,N_110);
nor U3275 (N_3275,N_424,N_1388);
or U3276 (N_3276,N_963,N_297);
nand U3277 (N_3277,N_417,N_1298);
and U3278 (N_3278,N_1010,N_1433);
xnor U3279 (N_3279,N_1972,N_2297);
or U3280 (N_3280,N_1218,N_320);
or U3281 (N_3281,N_1006,N_533);
nand U3282 (N_3282,N_2453,N_802);
nand U3283 (N_3283,N_778,N_1217);
nor U3284 (N_3284,N_1375,N_88);
and U3285 (N_3285,N_1161,N_2418);
and U3286 (N_3286,N_1693,N_315);
and U3287 (N_3287,N_947,N_688);
nor U3288 (N_3288,N_1156,N_1277);
nand U3289 (N_3289,N_553,N_1065);
and U3290 (N_3290,N_1829,N_1655);
nor U3291 (N_3291,N_1789,N_729);
nor U3292 (N_3292,N_1279,N_2355);
nand U3293 (N_3293,N_2070,N_2094);
and U3294 (N_3294,N_1008,N_1152);
and U3295 (N_3295,N_1525,N_567);
or U3296 (N_3296,N_2391,N_1710);
or U3297 (N_3297,N_2372,N_1692);
and U3298 (N_3298,N_2119,N_607);
and U3299 (N_3299,N_944,N_645);
and U3300 (N_3300,N_160,N_2211);
and U3301 (N_3301,N_2436,N_2113);
nand U3302 (N_3302,N_2033,N_2062);
or U3303 (N_3303,N_212,N_2353);
and U3304 (N_3304,N_2166,N_718);
and U3305 (N_3305,N_198,N_621);
nand U3306 (N_3306,N_334,N_254);
nand U3307 (N_3307,N_2399,N_2168);
nor U3308 (N_3308,N_1984,N_296);
nor U3309 (N_3309,N_485,N_1072);
and U3310 (N_3310,N_1328,N_32);
nand U3311 (N_3311,N_559,N_962);
or U3312 (N_3312,N_666,N_1317);
or U3313 (N_3313,N_2421,N_367);
nand U3314 (N_3314,N_109,N_2219);
xnor U3315 (N_3315,N_1151,N_1002);
nor U3316 (N_3316,N_2354,N_1442);
nand U3317 (N_3317,N_1991,N_488);
and U3318 (N_3318,N_2060,N_2149);
xnor U3319 (N_3319,N_2459,N_1982);
or U3320 (N_3320,N_132,N_1584);
or U3321 (N_3321,N_2308,N_1331);
nor U3322 (N_3322,N_1738,N_663);
nor U3323 (N_3323,N_929,N_912);
nand U3324 (N_3324,N_2367,N_677);
nor U3325 (N_3325,N_697,N_865);
and U3326 (N_3326,N_622,N_1261);
nand U3327 (N_3327,N_551,N_2484);
or U3328 (N_3328,N_114,N_1394);
or U3329 (N_3329,N_774,N_911);
nor U3330 (N_3330,N_39,N_1623);
nor U3331 (N_3331,N_193,N_810);
nor U3332 (N_3332,N_1147,N_686);
nor U3333 (N_3333,N_1314,N_2147);
and U3334 (N_3334,N_1266,N_87);
or U3335 (N_3335,N_310,N_1595);
nand U3336 (N_3336,N_1723,N_1541);
nor U3337 (N_3337,N_146,N_775);
or U3338 (N_3338,N_25,N_34);
and U3339 (N_3339,N_2112,N_1630);
nand U3340 (N_3340,N_656,N_1642);
nand U3341 (N_3341,N_717,N_23);
or U3342 (N_3342,N_1560,N_303);
nand U3343 (N_3343,N_9,N_538);
nor U3344 (N_3344,N_14,N_526);
nor U3345 (N_3345,N_1031,N_115);
nor U3346 (N_3346,N_1116,N_83);
or U3347 (N_3347,N_2217,N_40);
and U3348 (N_3348,N_2461,N_692);
and U3349 (N_3349,N_658,N_534);
and U3350 (N_3350,N_1384,N_942);
or U3351 (N_3351,N_670,N_33);
or U3352 (N_3352,N_1183,N_571);
or U3353 (N_3353,N_1240,N_147);
nor U3354 (N_3354,N_1814,N_1348);
and U3355 (N_3355,N_81,N_335);
nor U3356 (N_3356,N_1404,N_1435);
and U3357 (N_3357,N_322,N_1553);
nor U3358 (N_3358,N_585,N_862);
nand U3359 (N_3359,N_1221,N_2246);
nand U3360 (N_3360,N_29,N_1166);
and U3361 (N_3361,N_2241,N_2146);
and U3362 (N_3362,N_1150,N_429);
or U3363 (N_3363,N_421,N_1057);
nor U3364 (N_3364,N_597,N_195);
and U3365 (N_3365,N_1929,N_1869);
and U3366 (N_3366,N_2034,N_2210);
and U3367 (N_3367,N_2143,N_1282);
and U3368 (N_3368,N_518,N_155);
and U3369 (N_3369,N_1265,N_1043);
nor U3370 (N_3370,N_136,N_52);
and U3371 (N_3371,N_2144,N_333);
or U3372 (N_3372,N_976,N_1141);
nand U3373 (N_3373,N_696,N_187);
or U3374 (N_3374,N_2416,N_727);
nand U3375 (N_3375,N_1844,N_15);
or U3376 (N_3376,N_2439,N_768);
nor U3377 (N_3377,N_888,N_902);
nor U3378 (N_3378,N_1040,N_1296);
and U3379 (N_3379,N_690,N_1540);
and U3380 (N_3380,N_1644,N_1174);
and U3381 (N_3381,N_523,N_2451);
and U3382 (N_3382,N_2098,N_1205);
xor U3383 (N_3383,N_1460,N_1513);
or U3384 (N_3384,N_269,N_1066);
and U3385 (N_3385,N_255,N_1777);
nand U3386 (N_3386,N_1228,N_1294);
nand U3387 (N_3387,N_1886,N_1200);
nand U3388 (N_3388,N_170,N_1904);
nand U3389 (N_3389,N_937,N_318);
nand U3390 (N_3390,N_499,N_1609);
nor U3391 (N_3391,N_2267,N_1600);
nor U3392 (N_3392,N_873,N_196);
or U3393 (N_3393,N_1127,N_966);
or U3394 (N_3394,N_220,N_1346);
nor U3395 (N_3395,N_1376,N_785);
or U3396 (N_3396,N_1579,N_588);
nor U3397 (N_3397,N_1132,N_51);
nand U3398 (N_3398,N_2099,N_1964);
and U3399 (N_3399,N_844,N_933);
or U3400 (N_3400,N_758,N_1817);
nor U3401 (N_3401,N_675,N_2240);
or U3402 (N_3402,N_786,N_80);
nand U3403 (N_3403,N_886,N_495);
and U3404 (N_3404,N_351,N_1475);
xnor U3405 (N_3405,N_76,N_951);
nand U3406 (N_3406,N_2180,N_2464);
or U3407 (N_3407,N_748,N_1083);
nor U3408 (N_3408,N_1278,N_1327);
and U3409 (N_3409,N_990,N_1804);
nand U3410 (N_3410,N_946,N_332);
nand U3411 (N_3411,N_181,N_2405);
and U3412 (N_3412,N_1901,N_262);
xnor U3413 (N_3413,N_99,N_403);
nand U3414 (N_3414,N_669,N_1159);
and U3415 (N_3415,N_1358,N_594);
and U3416 (N_3416,N_1782,N_2408);
nand U3417 (N_3417,N_2435,N_1957);
and U3418 (N_3418,N_185,N_647);
nand U3419 (N_3419,N_1030,N_807);
nand U3420 (N_3420,N_477,N_489);
and U3421 (N_3421,N_1078,N_2080);
and U3422 (N_3422,N_725,N_258);
nor U3423 (N_3423,N_427,N_140);
nand U3424 (N_3424,N_982,N_2407);
or U3425 (N_3425,N_2022,N_1);
nand U3426 (N_3426,N_301,N_342);
nor U3427 (N_3427,N_2366,N_1024);
or U3428 (N_3428,N_1353,N_1516);
or U3429 (N_3429,N_36,N_462);
or U3430 (N_3430,N_1530,N_887);
or U3431 (N_3431,N_1535,N_1843);
nor U3432 (N_3432,N_1454,N_2079);
and U3433 (N_3433,N_175,N_2258);
or U3434 (N_3434,N_1365,N_707);
and U3435 (N_3435,N_1741,N_1716);
and U3436 (N_3436,N_1975,N_70);
nor U3437 (N_3437,N_259,N_1617);
or U3438 (N_3438,N_1654,N_2232);
and U3439 (N_3439,N_1055,N_1004);
nor U3440 (N_3440,N_1493,N_1153);
nor U3441 (N_3441,N_610,N_354);
and U3442 (N_3442,N_1989,N_2118);
nand U3443 (N_3443,N_2447,N_1946);
or U3444 (N_3444,N_1952,N_2181);
and U3445 (N_3445,N_761,N_98);
or U3446 (N_3446,N_2427,N_1438);
and U3447 (N_3447,N_1507,N_1146);
nor U3448 (N_3448,N_1958,N_1748);
nor U3449 (N_3449,N_2209,N_280);
nor U3450 (N_3450,N_706,N_1059);
and U3451 (N_3451,N_978,N_479);
nor U3452 (N_3452,N_1115,N_1237);
and U3453 (N_3453,N_2271,N_2379);
nor U3454 (N_3454,N_586,N_1090);
nand U3455 (N_3455,N_1480,N_328);
or U3456 (N_3456,N_2466,N_2190);
and U3457 (N_3457,N_769,N_740);
nand U3458 (N_3458,N_2344,N_2223);
nand U3459 (N_3459,N_2347,N_0);
nor U3460 (N_3460,N_662,N_2316);
and U3461 (N_3461,N_1921,N_2360);
and U3462 (N_3462,N_2192,N_752);
nand U3463 (N_3463,N_1401,N_1198);
nor U3464 (N_3464,N_66,N_701);
and U3465 (N_3465,N_896,N_584);
nor U3466 (N_3466,N_118,N_2058);
nand U3467 (N_3467,N_972,N_954);
nand U3468 (N_3468,N_1069,N_1512);
nor U3469 (N_3469,N_1845,N_1501);
nand U3470 (N_3470,N_2375,N_1877);
nor U3471 (N_3471,N_867,N_764);
nand U3472 (N_3472,N_826,N_1302);
nand U3473 (N_3473,N_1611,N_346);
and U3474 (N_3474,N_1639,N_2206);
and U3475 (N_3475,N_1342,N_782);
nand U3476 (N_3476,N_1416,N_714);
or U3477 (N_3477,N_2328,N_26);
or U3478 (N_3478,N_1079,N_674);
or U3479 (N_3479,N_2332,N_1664);
nor U3480 (N_3480,N_512,N_1258);
nor U3481 (N_3481,N_682,N_230);
and U3482 (N_3482,N_1746,N_89);
nand U3483 (N_3483,N_172,N_1571);
nand U3484 (N_3484,N_2270,N_2148);
and U3485 (N_3485,N_1145,N_531);
nor U3486 (N_3486,N_904,N_819);
nand U3487 (N_3487,N_964,N_1025);
and U3488 (N_3488,N_12,N_679);
and U3489 (N_3489,N_2340,N_1061);
nor U3490 (N_3490,N_1076,N_2284);
or U3491 (N_3491,N_1823,N_6);
and U3492 (N_3492,N_2311,N_2293);
nor U3493 (N_3493,N_2104,N_1750);
nand U3494 (N_3494,N_2324,N_1620);
or U3495 (N_3495,N_949,N_1465);
or U3496 (N_3496,N_991,N_1650);
xnor U3497 (N_3497,N_1749,N_617);
nor U3498 (N_3498,N_86,N_550);
nand U3499 (N_3499,N_240,N_428);
or U3500 (N_3500,N_2494,N_293);
nor U3501 (N_3501,N_843,N_1659);
nand U3502 (N_3502,N_460,N_1607);
nor U3503 (N_3503,N_672,N_1681);
and U3504 (N_3504,N_651,N_2337);
or U3505 (N_3505,N_264,N_1238);
nor U3506 (N_3506,N_766,N_2472);
nor U3507 (N_3507,N_1111,N_1599);
or U3508 (N_3508,N_1356,N_1118);
or U3509 (N_3509,N_1640,N_1722);
nand U3510 (N_3510,N_837,N_542);
or U3511 (N_3511,N_687,N_1017);
nand U3512 (N_3512,N_483,N_856);
and U3513 (N_3513,N_839,N_1808);
or U3514 (N_3514,N_1245,N_1468);
and U3515 (N_3515,N_128,N_243);
nand U3516 (N_3516,N_899,N_1763);
nor U3517 (N_3517,N_1428,N_444);
nor U3518 (N_3518,N_1842,N_324);
nand U3519 (N_3519,N_624,N_770);
nor U3520 (N_3520,N_1450,N_851);
nor U3521 (N_3521,N_640,N_2125);
and U3522 (N_3522,N_38,N_611);
nand U3523 (N_3523,N_2177,N_563);
or U3524 (N_3524,N_68,N_169);
and U3525 (N_3525,N_742,N_795);
nand U3526 (N_3526,N_1531,N_635);
or U3527 (N_3527,N_1618,N_1188);
and U3528 (N_3528,N_1143,N_728);
and U3529 (N_3529,N_1940,N_1029);
or U3530 (N_3530,N_285,N_78);
or U3531 (N_3531,N_1619,N_875);
or U3532 (N_3532,N_510,N_407);
or U3533 (N_3533,N_1555,N_404);
xnor U3534 (N_3534,N_2441,N_177);
or U3535 (N_3535,N_2448,N_932);
and U3536 (N_3536,N_2025,N_987);
and U3537 (N_3537,N_1334,N_2123);
or U3538 (N_3538,N_2236,N_62);
or U3539 (N_3539,N_1858,N_1626);
nand U3540 (N_3540,N_1047,N_924);
and U3541 (N_3541,N_2172,N_1853);
and U3542 (N_3542,N_2081,N_2235);
or U3543 (N_3543,N_2313,N_565);
nor U3544 (N_3544,N_961,N_1882);
nand U3545 (N_3545,N_2074,N_793);
or U3546 (N_3546,N_339,N_470);
and U3547 (N_3547,N_710,N_913);
or U3548 (N_3548,N_1943,N_861);
nand U3549 (N_3549,N_363,N_2390);
and U3550 (N_3550,N_480,N_1956);
nand U3551 (N_3551,N_2,N_623);
nand U3552 (N_3552,N_981,N_2362);
nor U3553 (N_3553,N_1894,N_1568);
nand U3554 (N_3554,N_1849,N_1694);
nand U3555 (N_3555,N_1547,N_1643);
xnor U3556 (N_3556,N_830,N_2214);
and U3557 (N_3557,N_535,N_1160);
nor U3558 (N_3558,N_1803,N_1382);
nor U3559 (N_3559,N_517,N_1962);
and U3560 (N_3560,N_628,N_934);
and U3561 (N_3561,N_348,N_1046);
or U3562 (N_3562,N_948,N_2159);
and U3563 (N_3563,N_1703,N_2193);
nand U3564 (N_3564,N_2044,N_2486);
nor U3565 (N_3565,N_587,N_1826);
or U3566 (N_3566,N_700,N_207);
nor U3567 (N_3567,N_668,N_776);
nand U3568 (N_3568,N_1509,N_2152);
nand U3569 (N_3569,N_1800,N_1671);
and U3570 (N_3570,N_2381,N_2468);
nand U3571 (N_3571,N_2349,N_2323);
or U3572 (N_3572,N_612,N_365);
nor U3573 (N_3573,N_231,N_2320);
and U3574 (N_3574,N_1403,N_2002);
and U3575 (N_3575,N_1735,N_2013);
nand U3576 (N_3576,N_2012,N_860);
and U3577 (N_3577,N_2085,N_1300);
nand U3578 (N_3578,N_1822,N_2200);
nor U3579 (N_3579,N_1488,N_2398);
nor U3580 (N_3580,N_13,N_244);
or U3581 (N_3581,N_445,N_1893);
nor U3582 (N_3582,N_1234,N_1903);
xnor U3583 (N_3583,N_1325,N_1253);
nor U3584 (N_3584,N_384,N_2434);
or U3585 (N_3585,N_808,N_2237);
nand U3586 (N_3586,N_1725,N_1648);
or U3587 (N_3587,N_2082,N_453);
nand U3588 (N_3588,N_102,N_2171);
nor U3589 (N_3589,N_871,N_516);
and U3590 (N_3590,N_547,N_1891);
nand U3591 (N_3591,N_2272,N_2032);
nor U3592 (N_3592,N_2222,N_1417);
or U3593 (N_3593,N_2076,N_2015);
and U3594 (N_3594,N_2165,N_2423);
and U3595 (N_3595,N_747,N_430);
or U3596 (N_3596,N_2274,N_1631);
nand U3597 (N_3597,N_926,N_1243);
and U3598 (N_3598,N_1542,N_2161);
and U3599 (N_3599,N_1209,N_1647);
nand U3600 (N_3600,N_2064,N_156);
or U3601 (N_3601,N_22,N_2250);
or U3602 (N_3602,N_1379,N_1335);
and U3603 (N_3603,N_564,N_11);
and U3604 (N_3604,N_2018,N_2126);
nand U3605 (N_3605,N_1015,N_1759);
and U3606 (N_3606,N_1260,N_1554);
nand U3607 (N_3607,N_79,N_387);
nand U3608 (N_3608,N_2365,N_1269);
nor U3609 (N_3609,N_2231,N_425);
nor U3610 (N_3610,N_454,N_2061);
and U3611 (N_3611,N_996,N_1987);
nand U3612 (N_3612,N_2173,N_1255);
and U3613 (N_3613,N_1470,N_317);
nor U3614 (N_3614,N_409,N_1138);
nand U3615 (N_3615,N_124,N_984);
nand U3616 (N_3616,N_2005,N_555);
nor U3617 (N_3617,N_1199,N_1397);
and U3618 (N_3618,N_627,N_221);
or U3619 (N_3619,N_557,N_733);
or U3620 (N_3620,N_2495,N_907);
nand U3621 (N_3621,N_233,N_619);
nand U3622 (N_3622,N_1434,N_1811);
nand U3623 (N_3623,N_1338,N_2368);
nor U3624 (N_3624,N_171,N_1638);
nand U3625 (N_3625,N_1036,N_1500);
nand U3626 (N_3626,N_2095,N_350);
or U3627 (N_3627,N_1805,N_277);
nor U3628 (N_3628,N_1473,N_958);
nand U3629 (N_3629,N_941,N_2404);
nor U3630 (N_3630,N_1649,N_2333);
and U3631 (N_3631,N_1892,N_1672);
or U3632 (N_3632,N_631,N_965);
and U3633 (N_3633,N_1256,N_1352);
nand U3634 (N_3634,N_2103,N_1021);
nor U3635 (N_3635,N_1075,N_1981);
and U3636 (N_3636,N_374,N_1603);
and U3637 (N_3637,N_30,N_2031);
nor U3638 (N_3638,N_1794,N_43);
nand U3639 (N_3639,N_1908,N_1884);
or U3640 (N_3640,N_1878,N_1459);
nand U3641 (N_3641,N_1606,N_545);
nor U3642 (N_3642,N_1950,N_2440);
nor U3643 (N_3643,N_1551,N_2445);
or U3644 (N_3644,N_1181,N_1458);
and U3645 (N_3645,N_410,N_2016);
nor U3646 (N_3646,N_1567,N_638);
or U3647 (N_3647,N_1616,N_1251);
or U3648 (N_3648,N_2289,N_1368);
nand U3649 (N_3649,N_525,N_781);
xor U3650 (N_3650,N_1969,N_1249);
nor U3651 (N_3651,N_313,N_1196);
nor U3652 (N_3652,N_1456,N_2043);
or U3653 (N_3653,N_242,N_166);
and U3654 (N_3654,N_1988,N_331);
and U3655 (N_3655,N_1839,N_1422);
or U3656 (N_3656,N_2273,N_2290);
nor U3657 (N_3657,N_478,N_1684);
and U3658 (N_3658,N_763,N_2097);
nand U3659 (N_3659,N_520,N_1953);
nor U3660 (N_3660,N_1178,N_1980);
and U3661 (N_3661,N_274,N_1699);
or U3662 (N_3662,N_514,N_305);
nand U3663 (N_3663,N_1915,N_1045);
nor U3664 (N_3664,N_341,N_1098);
nor U3665 (N_3665,N_1656,N_1696);
and U3666 (N_3666,N_809,N_1895);
or U3667 (N_3667,N_1263,N_655);
and U3668 (N_3668,N_251,N_281);
or U3669 (N_3669,N_2066,N_2038);
nand U3670 (N_3670,N_1344,N_2136);
or U3671 (N_3671,N_2196,N_2292);
and U3672 (N_3672,N_2133,N_272);
nor U3673 (N_3673,N_1544,N_569);
or U3674 (N_3674,N_2321,N_2414);
nor U3675 (N_3675,N_854,N_639);
and U3676 (N_3676,N_284,N_1526);
and U3677 (N_3677,N_1114,N_2051);
and U3678 (N_3678,N_1812,N_2162);
nand U3679 (N_3679,N_1101,N_2306);
or U3680 (N_3680,N_595,N_598);
or U3681 (N_3681,N_442,N_2426);
and U3682 (N_3682,N_2182,N_2248);
and U3683 (N_3683,N_1628,N_1744);
and U3684 (N_3684,N_1242,N_2454);
nand U3685 (N_3685,N_2008,N_2175);
and U3686 (N_3686,N_2343,N_985);
or U3687 (N_3687,N_2383,N_1704);
nand U3688 (N_3688,N_1707,N_1996);
nor U3689 (N_3689,N_1993,N_2358);
nand U3690 (N_3690,N_176,N_1295);
and U3691 (N_3691,N_1123,N_1499);
nand U3692 (N_3692,N_121,N_337);
nor U3693 (N_3693,N_979,N_751);
nor U3694 (N_3694,N_1074,N_788);
nor U3695 (N_3695,N_406,N_1930);
nor U3696 (N_3696,N_1313,N_1949);
nor U3697 (N_3697,N_1064,N_1370);
nor U3698 (N_3698,N_1301,N_1875);
and U3699 (N_3699,N_440,N_1818);
or U3700 (N_3700,N_1484,N_232);
nand U3701 (N_3701,N_2023,N_908);
or U3702 (N_3702,N_1247,N_321);
nor U3703 (N_3703,N_431,N_2296);
nor U3704 (N_3704,N_2298,N_1690);
and U3705 (N_3705,N_1155,N_1167);
and U3706 (N_3706,N_1103,N_2215);
nor U3707 (N_3707,N_1820,N_64);
nor U3708 (N_3708,N_1395,N_2433);
nand U3709 (N_3709,N_394,N_1318);
nand U3710 (N_3710,N_2339,N_149);
nor U3711 (N_3711,N_159,N_1787);
and U3712 (N_3712,N_2471,N_762);
xor U3713 (N_3713,N_613,N_1172);
and U3714 (N_3714,N_358,N_684);
nand U3715 (N_3715,N_1362,N_1377);
or U3716 (N_3716,N_1756,N_37);
or U3717 (N_3717,N_1086,N_767);
xnor U3718 (N_3718,N_1336,N_381);
and U3719 (N_3719,N_165,N_1840);
nand U3720 (N_3720,N_2374,N_1848);
or U3721 (N_3721,N_1007,N_2491);
nand U3722 (N_3722,N_574,N_676);
and U3723 (N_3723,N_117,N_1248);
and U3724 (N_3724,N_544,N_357);
nand U3725 (N_3725,N_618,N_1565);
nand U3726 (N_3726,N_44,N_267);
nor U3727 (N_3727,N_96,N_1898);
nand U3728 (N_3728,N_1721,N_1140);
nor U3729 (N_3729,N_67,N_21);
or U3730 (N_3730,N_418,N_1497);
and U3731 (N_3731,N_2091,N_1920);
nand U3732 (N_3732,N_1679,N_378);
and U3733 (N_3733,N_2499,N_1906);
and U3734 (N_3734,N_1038,N_2331);
nand U3735 (N_3735,N_396,N_625);
nand U3736 (N_3736,N_992,N_901);
and U3737 (N_3737,N_1689,N_606);
nand U3738 (N_3738,N_1191,N_1421);
nor U3739 (N_3739,N_2069,N_1919);
or U3740 (N_3740,N_1476,N_1216);
nor U3741 (N_3741,N_249,N_1479);
nor U3742 (N_3742,N_271,N_205);
and U3743 (N_3743,N_3,N_630);
nand U3744 (N_3744,N_1727,N_2409);
and U3745 (N_3745,N_2481,N_1557);
and U3746 (N_3746,N_1752,N_1430);
or U3747 (N_3747,N_273,N_2282);
nand U3748 (N_3748,N_438,N_1303);
and U3749 (N_3749,N_940,N_192);
nor U3750 (N_3750,N_2433,N_649);
and U3751 (N_3751,N_466,N_1500);
nand U3752 (N_3752,N_1509,N_1736);
or U3753 (N_3753,N_1087,N_886);
nand U3754 (N_3754,N_2468,N_1186);
nor U3755 (N_3755,N_1723,N_373);
nand U3756 (N_3756,N_776,N_623);
nor U3757 (N_3757,N_1359,N_2279);
nand U3758 (N_3758,N_1455,N_428);
nand U3759 (N_3759,N_1982,N_418);
nand U3760 (N_3760,N_711,N_1304);
nand U3761 (N_3761,N_1023,N_1891);
nand U3762 (N_3762,N_1193,N_1528);
nor U3763 (N_3763,N_1446,N_1793);
or U3764 (N_3764,N_2176,N_1482);
or U3765 (N_3765,N_2301,N_1623);
nor U3766 (N_3766,N_683,N_960);
xnor U3767 (N_3767,N_1881,N_518);
and U3768 (N_3768,N_1161,N_294);
nand U3769 (N_3769,N_508,N_1129);
or U3770 (N_3770,N_220,N_242);
or U3771 (N_3771,N_491,N_1918);
or U3772 (N_3772,N_1498,N_757);
nand U3773 (N_3773,N_998,N_192);
nor U3774 (N_3774,N_2380,N_682);
nand U3775 (N_3775,N_1679,N_915);
or U3776 (N_3776,N_299,N_2126);
or U3777 (N_3777,N_120,N_512);
or U3778 (N_3778,N_1946,N_1459);
nand U3779 (N_3779,N_127,N_1478);
nor U3780 (N_3780,N_1022,N_1968);
or U3781 (N_3781,N_909,N_945);
and U3782 (N_3782,N_1971,N_2059);
nor U3783 (N_3783,N_2165,N_2155);
nor U3784 (N_3784,N_119,N_2248);
nor U3785 (N_3785,N_341,N_1919);
and U3786 (N_3786,N_2128,N_341);
nor U3787 (N_3787,N_1983,N_1004);
and U3788 (N_3788,N_1617,N_546);
and U3789 (N_3789,N_1006,N_404);
or U3790 (N_3790,N_2486,N_1701);
nor U3791 (N_3791,N_1495,N_1029);
nand U3792 (N_3792,N_2123,N_2456);
nand U3793 (N_3793,N_583,N_1765);
nand U3794 (N_3794,N_32,N_789);
nor U3795 (N_3795,N_1462,N_190);
xnor U3796 (N_3796,N_1255,N_1791);
or U3797 (N_3797,N_250,N_931);
nor U3798 (N_3798,N_2094,N_2338);
or U3799 (N_3799,N_910,N_470);
and U3800 (N_3800,N_2105,N_1426);
nor U3801 (N_3801,N_2335,N_458);
or U3802 (N_3802,N_445,N_1703);
nor U3803 (N_3803,N_2184,N_122);
or U3804 (N_3804,N_552,N_1614);
or U3805 (N_3805,N_1716,N_1306);
and U3806 (N_3806,N_1247,N_2278);
and U3807 (N_3807,N_1942,N_1755);
nor U3808 (N_3808,N_2489,N_473);
xnor U3809 (N_3809,N_92,N_2238);
and U3810 (N_3810,N_1108,N_316);
or U3811 (N_3811,N_1878,N_751);
and U3812 (N_3812,N_947,N_1585);
nand U3813 (N_3813,N_698,N_966);
or U3814 (N_3814,N_268,N_1196);
or U3815 (N_3815,N_1046,N_276);
and U3816 (N_3816,N_713,N_522);
and U3817 (N_3817,N_664,N_63);
nor U3818 (N_3818,N_1687,N_250);
nand U3819 (N_3819,N_613,N_1994);
nor U3820 (N_3820,N_2390,N_78);
nor U3821 (N_3821,N_2439,N_1730);
nand U3822 (N_3822,N_420,N_323);
nand U3823 (N_3823,N_1210,N_1163);
or U3824 (N_3824,N_5,N_1646);
or U3825 (N_3825,N_505,N_1512);
or U3826 (N_3826,N_940,N_2);
nand U3827 (N_3827,N_1403,N_683);
or U3828 (N_3828,N_666,N_2248);
nand U3829 (N_3829,N_2389,N_1260);
or U3830 (N_3830,N_2243,N_1431);
nor U3831 (N_3831,N_423,N_1637);
nor U3832 (N_3832,N_224,N_362);
and U3833 (N_3833,N_2168,N_1800);
or U3834 (N_3834,N_755,N_902);
and U3835 (N_3835,N_2232,N_735);
nor U3836 (N_3836,N_1046,N_1882);
nand U3837 (N_3837,N_1405,N_151);
and U3838 (N_3838,N_425,N_2152);
or U3839 (N_3839,N_1824,N_1313);
and U3840 (N_3840,N_1961,N_1741);
or U3841 (N_3841,N_1010,N_1005);
or U3842 (N_3842,N_973,N_1915);
nor U3843 (N_3843,N_107,N_738);
nor U3844 (N_3844,N_89,N_789);
nor U3845 (N_3845,N_349,N_1150);
and U3846 (N_3846,N_1112,N_728);
nand U3847 (N_3847,N_2425,N_904);
and U3848 (N_3848,N_709,N_610);
and U3849 (N_3849,N_1000,N_2087);
or U3850 (N_3850,N_1807,N_2361);
and U3851 (N_3851,N_1878,N_2185);
nor U3852 (N_3852,N_706,N_1145);
nor U3853 (N_3853,N_311,N_1459);
and U3854 (N_3854,N_2361,N_1868);
nand U3855 (N_3855,N_1941,N_1940);
or U3856 (N_3856,N_2348,N_1392);
and U3857 (N_3857,N_444,N_47);
nor U3858 (N_3858,N_1645,N_1256);
nand U3859 (N_3859,N_713,N_1771);
and U3860 (N_3860,N_1465,N_2022);
and U3861 (N_3861,N_2107,N_691);
or U3862 (N_3862,N_1312,N_445);
or U3863 (N_3863,N_1350,N_2247);
and U3864 (N_3864,N_1070,N_2346);
nor U3865 (N_3865,N_1457,N_720);
nor U3866 (N_3866,N_984,N_1116);
nor U3867 (N_3867,N_282,N_1045);
or U3868 (N_3868,N_2495,N_1453);
nor U3869 (N_3869,N_2182,N_2214);
nor U3870 (N_3870,N_412,N_730);
and U3871 (N_3871,N_1943,N_2295);
and U3872 (N_3872,N_1072,N_738);
or U3873 (N_3873,N_1962,N_855);
and U3874 (N_3874,N_1615,N_1683);
nand U3875 (N_3875,N_433,N_1699);
nand U3876 (N_3876,N_2278,N_2070);
nand U3877 (N_3877,N_1060,N_856);
nor U3878 (N_3878,N_44,N_328);
or U3879 (N_3879,N_1989,N_1043);
nor U3880 (N_3880,N_1620,N_51);
or U3881 (N_3881,N_982,N_2098);
nor U3882 (N_3882,N_2058,N_588);
and U3883 (N_3883,N_2452,N_863);
or U3884 (N_3884,N_1783,N_195);
nand U3885 (N_3885,N_1544,N_2370);
nand U3886 (N_3886,N_664,N_861);
nor U3887 (N_3887,N_1652,N_1646);
and U3888 (N_3888,N_1656,N_1080);
nor U3889 (N_3889,N_2194,N_815);
nor U3890 (N_3890,N_2210,N_1526);
and U3891 (N_3891,N_2477,N_348);
xnor U3892 (N_3892,N_2142,N_1739);
and U3893 (N_3893,N_1931,N_247);
nor U3894 (N_3894,N_70,N_1893);
nor U3895 (N_3895,N_1264,N_1126);
and U3896 (N_3896,N_316,N_1323);
nor U3897 (N_3897,N_2441,N_2);
nand U3898 (N_3898,N_1330,N_1001);
nand U3899 (N_3899,N_1551,N_2018);
nand U3900 (N_3900,N_917,N_1081);
and U3901 (N_3901,N_2204,N_1008);
nand U3902 (N_3902,N_24,N_2424);
nand U3903 (N_3903,N_57,N_2112);
and U3904 (N_3904,N_534,N_2248);
nor U3905 (N_3905,N_1355,N_2455);
and U3906 (N_3906,N_1539,N_1596);
or U3907 (N_3907,N_1981,N_1744);
nand U3908 (N_3908,N_854,N_609);
and U3909 (N_3909,N_1024,N_1943);
or U3910 (N_3910,N_2042,N_2011);
or U3911 (N_3911,N_360,N_265);
or U3912 (N_3912,N_863,N_957);
nor U3913 (N_3913,N_902,N_2210);
and U3914 (N_3914,N_434,N_1949);
nor U3915 (N_3915,N_1996,N_815);
and U3916 (N_3916,N_2385,N_1014);
and U3917 (N_3917,N_1274,N_1993);
or U3918 (N_3918,N_2491,N_2163);
nor U3919 (N_3919,N_249,N_875);
or U3920 (N_3920,N_229,N_2198);
nand U3921 (N_3921,N_1340,N_1088);
and U3922 (N_3922,N_1309,N_1820);
and U3923 (N_3923,N_36,N_367);
and U3924 (N_3924,N_2355,N_1316);
nor U3925 (N_3925,N_16,N_1331);
or U3926 (N_3926,N_1099,N_1602);
or U3927 (N_3927,N_684,N_1045);
nand U3928 (N_3928,N_195,N_2040);
nor U3929 (N_3929,N_101,N_1156);
nor U3930 (N_3930,N_2204,N_2456);
and U3931 (N_3931,N_1103,N_212);
nand U3932 (N_3932,N_747,N_1116);
or U3933 (N_3933,N_1552,N_788);
or U3934 (N_3934,N_1481,N_265);
nor U3935 (N_3935,N_2030,N_203);
nor U3936 (N_3936,N_2451,N_794);
and U3937 (N_3937,N_10,N_2205);
or U3938 (N_3938,N_2051,N_168);
and U3939 (N_3939,N_1312,N_264);
nor U3940 (N_3940,N_2209,N_1371);
nor U3941 (N_3941,N_192,N_1394);
and U3942 (N_3942,N_141,N_1562);
and U3943 (N_3943,N_1859,N_340);
nand U3944 (N_3944,N_1218,N_924);
and U3945 (N_3945,N_2049,N_512);
or U3946 (N_3946,N_394,N_292);
and U3947 (N_3947,N_1204,N_1704);
and U3948 (N_3948,N_1676,N_2443);
and U3949 (N_3949,N_1760,N_1807);
nand U3950 (N_3950,N_2101,N_1807);
and U3951 (N_3951,N_472,N_1715);
or U3952 (N_3952,N_1412,N_1884);
and U3953 (N_3953,N_1570,N_2204);
nor U3954 (N_3954,N_986,N_1001);
or U3955 (N_3955,N_1542,N_1409);
and U3956 (N_3956,N_469,N_332);
or U3957 (N_3957,N_1586,N_784);
and U3958 (N_3958,N_2337,N_810);
nor U3959 (N_3959,N_1184,N_1949);
nor U3960 (N_3960,N_1206,N_2088);
nor U3961 (N_3961,N_2175,N_2027);
nand U3962 (N_3962,N_2241,N_2385);
and U3963 (N_3963,N_272,N_375);
and U3964 (N_3964,N_2278,N_197);
nand U3965 (N_3965,N_520,N_2253);
nor U3966 (N_3966,N_1260,N_1661);
and U3967 (N_3967,N_888,N_1857);
nand U3968 (N_3968,N_1220,N_1081);
nor U3969 (N_3969,N_32,N_2384);
nand U3970 (N_3970,N_630,N_647);
nor U3971 (N_3971,N_380,N_1709);
nor U3972 (N_3972,N_1727,N_408);
nor U3973 (N_3973,N_1668,N_1569);
and U3974 (N_3974,N_2485,N_363);
and U3975 (N_3975,N_1801,N_1881);
nor U3976 (N_3976,N_1042,N_1632);
nand U3977 (N_3977,N_591,N_2427);
nor U3978 (N_3978,N_183,N_1811);
and U3979 (N_3979,N_1393,N_1514);
or U3980 (N_3980,N_1925,N_1746);
nand U3981 (N_3981,N_2131,N_1080);
and U3982 (N_3982,N_2128,N_1845);
nand U3983 (N_3983,N_1181,N_103);
and U3984 (N_3984,N_2356,N_1787);
or U3985 (N_3985,N_1633,N_2254);
and U3986 (N_3986,N_1716,N_172);
or U3987 (N_3987,N_1281,N_1091);
nand U3988 (N_3988,N_1139,N_2210);
and U3989 (N_3989,N_636,N_1451);
or U3990 (N_3990,N_1709,N_332);
or U3991 (N_3991,N_947,N_814);
and U3992 (N_3992,N_1886,N_730);
and U3993 (N_3993,N_579,N_2193);
or U3994 (N_3994,N_1536,N_1317);
and U3995 (N_3995,N_2180,N_1427);
and U3996 (N_3996,N_592,N_809);
or U3997 (N_3997,N_1707,N_1703);
or U3998 (N_3998,N_651,N_2397);
nor U3999 (N_3999,N_398,N_710);
or U4000 (N_4000,N_1063,N_1554);
and U4001 (N_4001,N_1746,N_1021);
nor U4002 (N_4002,N_1201,N_646);
nor U4003 (N_4003,N_531,N_517);
nor U4004 (N_4004,N_658,N_1906);
or U4005 (N_4005,N_1649,N_1309);
or U4006 (N_4006,N_379,N_347);
and U4007 (N_4007,N_2170,N_217);
nor U4008 (N_4008,N_2318,N_39);
or U4009 (N_4009,N_618,N_1168);
or U4010 (N_4010,N_2359,N_1229);
or U4011 (N_4011,N_25,N_826);
and U4012 (N_4012,N_707,N_867);
nor U4013 (N_4013,N_1491,N_477);
or U4014 (N_4014,N_817,N_180);
nor U4015 (N_4015,N_931,N_2082);
or U4016 (N_4016,N_2015,N_501);
or U4017 (N_4017,N_1552,N_2002);
nand U4018 (N_4018,N_1065,N_2339);
and U4019 (N_4019,N_873,N_724);
or U4020 (N_4020,N_1888,N_2073);
nand U4021 (N_4021,N_850,N_134);
or U4022 (N_4022,N_643,N_2058);
nor U4023 (N_4023,N_2069,N_104);
and U4024 (N_4024,N_2378,N_914);
and U4025 (N_4025,N_1993,N_720);
nor U4026 (N_4026,N_933,N_792);
nand U4027 (N_4027,N_2183,N_23);
or U4028 (N_4028,N_2357,N_1674);
nand U4029 (N_4029,N_1233,N_1168);
nand U4030 (N_4030,N_1362,N_1425);
and U4031 (N_4031,N_1867,N_2142);
nor U4032 (N_4032,N_266,N_1996);
xor U4033 (N_4033,N_294,N_1811);
nand U4034 (N_4034,N_1210,N_2312);
or U4035 (N_4035,N_718,N_49);
nand U4036 (N_4036,N_480,N_1022);
nand U4037 (N_4037,N_612,N_752);
nor U4038 (N_4038,N_1861,N_2062);
and U4039 (N_4039,N_999,N_57);
nor U4040 (N_4040,N_802,N_1400);
or U4041 (N_4041,N_233,N_609);
and U4042 (N_4042,N_964,N_700);
and U4043 (N_4043,N_1701,N_225);
and U4044 (N_4044,N_929,N_104);
nand U4045 (N_4045,N_1245,N_2205);
nor U4046 (N_4046,N_1738,N_1799);
nor U4047 (N_4047,N_1519,N_1885);
nor U4048 (N_4048,N_748,N_708);
and U4049 (N_4049,N_685,N_1948);
nand U4050 (N_4050,N_67,N_1107);
and U4051 (N_4051,N_1377,N_1110);
and U4052 (N_4052,N_917,N_297);
or U4053 (N_4053,N_1981,N_1962);
or U4054 (N_4054,N_1493,N_522);
or U4055 (N_4055,N_1234,N_13);
and U4056 (N_4056,N_1206,N_60);
nand U4057 (N_4057,N_42,N_831);
or U4058 (N_4058,N_1477,N_826);
nand U4059 (N_4059,N_1663,N_2182);
or U4060 (N_4060,N_120,N_2379);
xnor U4061 (N_4061,N_596,N_1274);
or U4062 (N_4062,N_165,N_493);
nor U4063 (N_4063,N_972,N_2176);
nor U4064 (N_4064,N_1377,N_2175);
and U4065 (N_4065,N_1354,N_1325);
nor U4066 (N_4066,N_692,N_187);
or U4067 (N_4067,N_1497,N_1556);
or U4068 (N_4068,N_1951,N_2104);
nor U4069 (N_4069,N_1633,N_2040);
and U4070 (N_4070,N_1599,N_1473);
and U4071 (N_4071,N_538,N_153);
nor U4072 (N_4072,N_756,N_590);
nand U4073 (N_4073,N_1621,N_21);
or U4074 (N_4074,N_1051,N_124);
nand U4075 (N_4075,N_1655,N_1283);
and U4076 (N_4076,N_494,N_2340);
or U4077 (N_4077,N_1538,N_1732);
or U4078 (N_4078,N_1479,N_1631);
nor U4079 (N_4079,N_224,N_2022);
or U4080 (N_4080,N_1425,N_195);
nand U4081 (N_4081,N_2465,N_751);
nand U4082 (N_4082,N_1535,N_1508);
nor U4083 (N_4083,N_245,N_2073);
xor U4084 (N_4084,N_2139,N_960);
nor U4085 (N_4085,N_310,N_875);
nor U4086 (N_4086,N_1458,N_1971);
nand U4087 (N_4087,N_1569,N_1220);
or U4088 (N_4088,N_906,N_2010);
nand U4089 (N_4089,N_1096,N_1601);
nor U4090 (N_4090,N_13,N_1001);
or U4091 (N_4091,N_59,N_1280);
and U4092 (N_4092,N_1156,N_2464);
and U4093 (N_4093,N_2249,N_2092);
and U4094 (N_4094,N_1130,N_1391);
nor U4095 (N_4095,N_1973,N_1793);
or U4096 (N_4096,N_58,N_213);
nor U4097 (N_4097,N_674,N_1808);
and U4098 (N_4098,N_1241,N_897);
and U4099 (N_4099,N_1713,N_2134);
and U4100 (N_4100,N_96,N_493);
and U4101 (N_4101,N_1839,N_421);
nand U4102 (N_4102,N_2205,N_2305);
nor U4103 (N_4103,N_2257,N_2172);
or U4104 (N_4104,N_19,N_681);
nor U4105 (N_4105,N_2411,N_1567);
nor U4106 (N_4106,N_2383,N_1334);
nor U4107 (N_4107,N_1450,N_2264);
nand U4108 (N_4108,N_1527,N_1071);
or U4109 (N_4109,N_2159,N_1172);
nor U4110 (N_4110,N_234,N_2390);
nor U4111 (N_4111,N_955,N_1014);
or U4112 (N_4112,N_1031,N_1052);
or U4113 (N_4113,N_1707,N_1529);
nor U4114 (N_4114,N_1096,N_1810);
and U4115 (N_4115,N_1085,N_1113);
nand U4116 (N_4116,N_156,N_2432);
and U4117 (N_4117,N_846,N_1964);
or U4118 (N_4118,N_1454,N_1582);
nand U4119 (N_4119,N_32,N_2279);
nor U4120 (N_4120,N_153,N_1711);
nor U4121 (N_4121,N_108,N_206);
or U4122 (N_4122,N_1078,N_2112);
or U4123 (N_4123,N_332,N_860);
nor U4124 (N_4124,N_2262,N_226);
nand U4125 (N_4125,N_4,N_1520);
or U4126 (N_4126,N_2293,N_1487);
and U4127 (N_4127,N_1014,N_455);
or U4128 (N_4128,N_1030,N_2155);
and U4129 (N_4129,N_314,N_1431);
and U4130 (N_4130,N_1675,N_1491);
nand U4131 (N_4131,N_1408,N_800);
and U4132 (N_4132,N_1896,N_2108);
and U4133 (N_4133,N_335,N_1150);
or U4134 (N_4134,N_431,N_746);
nor U4135 (N_4135,N_464,N_194);
nand U4136 (N_4136,N_1020,N_1135);
nand U4137 (N_4137,N_397,N_2084);
nor U4138 (N_4138,N_114,N_1904);
nand U4139 (N_4139,N_2332,N_1732);
nor U4140 (N_4140,N_800,N_174);
nor U4141 (N_4141,N_512,N_826);
and U4142 (N_4142,N_522,N_1443);
or U4143 (N_4143,N_517,N_2447);
or U4144 (N_4144,N_1055,N_805);
and U4145 (N_4145,N_569,N_1356);
and U4146 (N_4146,N_2191,N_2436);
and U4147 (N_4147,N_1165,N_862);
and U4148 (N_4148,N_141,N_241);
and U4149 (N_4149,N_65,N_761);
nand U4150 (N_4150,N_1710,N_2465);
and U4151 (N_4151,N_922,N_199);
nor U4152 (N_4152,N_648,N_731);
nor U4153 (N_4153,N_1604,N_2006);
nor U4154 (N_4154,N_749,N_2479);
nand U4155 (N_4155,N_1668,N_160);
nand U4156 (N_4156,N_2059,N_1814);
nor U4157 (N_4157,N_1306,N_155);
and U4158 (N_4158,N_2060,N_1517);
nor U4159 (N_4159,N_1162,N_246);
nor U4160 (N_4160,N_793,N_1112);
or U4161 (N_4161,N_1762,N_612);
and U4162 (N_4162,N_994,N_1989);
nand U4163 (N_4163,N_709,N_708);
and U4164 (N_4164,N_971,N_2123);
nand U4165 (N_4165,N_1277,N_900);
or U4166 (N_4166,N_2138,N_801);
nor U4167 (N_4167,N_54,N_1906);
and U4168 (N_4168,N_474,N_1181);
or U4169 (N_4169,N_32,N_1032);
nand U4170 (N_4170,N_830,N_2016);
nand U4171 (N_4171,N_1051,N_2175);
or U4172 (N_4172,N_2099,N_948);
nor U4173 (N_4173,N_298,N_1495);
nor U4174 (N_4174,N_1696,N_928);
and U4175 (N_4175,N_694,N_625);
nand U4176 (N_4176,N_2388,N_27);
nor U4177 (N_4177,N_1847,N_61);
nor U4178 (N_4178,N_1505,N_1312);
nor U4179 (N_4179,N_1890,N_653);
and U4180 (N_4180,N_839,N_1730);
nor U4181 (N_4181,N_9,N_783);
nand U4182 (N_4182,N_980,N_932);
or U4183 (N_4183,N_2464,N_1297);
or U4184 (N_4184,N_2236,N_1278);
nand U4185 (N_4185,N_545,N_862);
xor U4186 (N_4186,N_482,N_1608);
nand U4187 (N_4187,N_1887,N_1551);
nor U4188 (N_4188,N_267,N_2205);
or U4189 (N_4189,N_2154,N_1277);
nand U4190 (N_4190,N_523,N_267);
or U4191 (N_4191,N_52,N_1775);
nor U4192 (N_4192,N_142,N_368);
nor U4193 (N_4193,N_471,N_1900);
and U4194 (N_4194,N_1866,N_1673);
and U4195 (N_4195,N_332,N_1920);
or U4196 (N_4196,N_2019,N_603);
or U4197 (N_4197,N_135,N_1575);
nand U4198 (N_4198,N_808,N_2102);
and U4199 (N_4199,N_1740,N_1165);
nand U4200 (N_4200,N_778,N_2115);
nand U4201 (N_4201,N_1512,N_2272);
nor U4202 (N_4202,N_912,N_1575);
nand U4203 (N_4203,N_1601,N_1295);
nor U4204 (N_4204,N_1270,N_2334);
nand U4205 (N_4205,N_1876,N_2225);
or U4206 (N_4206,N_567,N_1046);
nand U4207 (N_4207,N_1907,N_1839);
nand U4208 (N_4208,N_1568,N_950);
or U4209 (N_4209,N_389,N_2140);
nand U4210 (N_4210,N_1887,N_2351);
and U4211 (N_4211,N_315,N_2229);
nor U4212 (N_4212,N_90,N_2360);
and U4213 (N_4213,N_1497,N_1483);
or U4214 (N_4214,N_1493,N_1619);
nor U4215 (N_4215,N_985,N_166);
nor U4216 (N_4216,N_1264,N_2201);
or U4217 (N_4217,N_2098,N_1682);
and U4218 (N_4218,N_733,N_351);
or U4219 (N_4219,N_288,N_828);
or U4220 (N_4220,N_1457,N_927);
or U4221 (N_4221,N_1977,N_370);
or U4222 (N_4222,N_1451,N_1556);
xor U4223 (N_4223,N_366,N_1209);
nand U4224 (N_4224,N_1191,N_2377);
and U4225 (N_4225,N_106,N_419);
and U4226 (N_4226,N_1983,N_1514);
nor U4227 (N_4227,N_2445,N_356);
nand U4228 (N_4228,N_1506,N_1822);
and U4229 (N_4229,N_1188,N_1275);
nand U4230 (N_4230,N_1557,N_1409);
or U4231 (N_4231,N_443,N_277);
nand U4232 (N_4232,N_1704,N_121);
or U4233 (N_4233,N_2128,N_747);
nor U4234 (N_4234,N_2286,N_1690);
and U4235 (N_4235,N_1624,N_241);
nand U4236 (N_4236,N_1314,N_2363);
nor U4237 (N_4237,N_1516,N_2390);
and U4238 (N_4238,N_1812,N_2275);
nor U4239 (N_4239,N_2217,N_1063);
nor U4240 (N_4240,N_1430,N_983);
or U4241 (N_4241,N_483,N_2241);
or U4242 (N_4242,N_2391,N_209);
and U4243 (N_4243,N_1321,N_1783);
or U4244 (N_4244,N_1436,N_620);
nand U4245 (N_4245,N_662,N_1471);
and U4246 (N_4246,N_1568,N_349);
nor U4247 (N_4247,N_1236,N_524);
nor U4248 (N_4248,N_1158,N_1247);
and U4249 (N_4249,N_1666,N_233);
nand U4250 (N_4250,N_2443,N_277);
or U4251 (N_4251,N_79,N_2020);
nand U4252 (N_4252,N_2355,N_100);
nand U4253 (N_4253,N_22,N_2374);
and U4254 (N_4254,N_2069,N_1951);
nand U4255 (N_4255,N_1617,N_1715);
nand U4256 (N_4256,N_1567,N_1849);
nand U4257 (N_4257,N_1337,N_65);
nor U4258 (N_4258,N_783,N_1343);
nor U4259 (N_4259,N_409,N_1106);
nor U4260 (N_4260,N_520,N_2346);
and U4261 (N_4261,N_2406,N_2064);
xnor U4262 (N_4262,N_1668,N_1624);
or U4263 (N_4263,N_930,N_575);
and U4264 (N_4264,N_378,N_1471);
and U4265 (N_4265,N_481,N_827);
nor U4266 (N_4266,N_2083,N_254);
and U4267 (N_4267,N_447,N_1310);
and U4268 (N_4268,N_1202,N_1867);
and U4269 (N_4269,N_934,N_951);
nor U4270 (N_4270,N_2259,N_1864);
or U4271 (N_4271,N_1071,N_579);
xor U4272 (N_4272,N_2258,N_499);
and U4273 (N_4273,N_2353,N_577);
nor U4274 (N_4274,N_1693,N_1320);
nand U4275 (N_4275,N_1797,N_1840);
nor U4276 (N_4276,N_1483,N_475);
or U4277 (N_4277,N_169,N_418);
nor U4278 (N_4278,N_1469,N_1742);
or U4279 (N_4279,N_1970,N_256);
nor U4280 (N_4280,N_2228,N_1186);
nand U4281 (N_4281,N_830,N_634);
nor U4282 (N_4282,N_1298,N_1244);
nand U4283 (N_4283,N_1598,N_1546);
nand U4284 (N_4284,N_1855,N_1395);
nor U4285 (N_4285,N_1424,N_1591);
nor U4286 (N_4286,N_1799,N_1376);
and U4287 (N_4287,N_923,N_757);
nor U4288 (N_4288,N_2323,N_2054);
nor U4289 (N_4289,N_2075,N_1934);
nand U4290 (N_4290,N_29,N_2077);
nand U4291 (N_4291,N_2099,N_1547);
nor U4292 (N_4292,N_2315,N_290);
nand U4293 (N_4293,N_369,N_1734);
nand U4294 (N_4294,N_713,N_964);
nand U4295 (N_4295,N_44,N_1247);
or U4296 (N_4296,N_2398,N_1501);
and U4297 (N_4297,N_1499,N_144);
and U4298 (N_4298,N_1181,N_1285);
nor U4299 (N_4299,N_61,N_1218);
or U4300 (N_4300,N_2161,N_2003);
nand U4301 (N_4301,N_476,N_1157);
and U4302 (N_4302,N_1657,N_508);
nor U4303 (N_4303,N_2442,N_336);
nand U4304 (N_4304,N_575,N_2160);
nand U4305 (N_4305,N_752,N_400);
nor U4306 (N_4306,N_1680,N_1085);
nor U4307 (N_4307,N_1688,N_1644);
and U4308 (N_4308,N_2315,N_2466);
and U4309 (N_4309,N_1881,N_1204);
nor U4310 (N_4310,N_692,N_635);
nor U4311 (N_4311,N_2211,N_1849);
nor U4312 (N_4312,N_35,N_1502);
nand U4313 (N_4313,N_359,N_920);
nor U4314 (N_4314,N_759,N_1783);
nor U4315 (N_4315,N_1237,N_2180);
nor U4316 (N_4316,N_2303,N_2005);
nor U4317 (N_4317,N_921,N_1199);
and U4318 (N_4318,N_1477,N_430);
nand U4319 (N_4319,N_2479,N_1088);
nor U4320 (N_4320,N_960,N_48);
nand U4321 (N_4321,N_1784,N_2425);
nand U4322 (N_4322,N_2343,N_1227);
nor U4323 (N_4323,N_1290,N_2276);
nor U4324 (N_4324,N_1357,N_1396);
or U4325 (N_4325,N_1671,N_2415);
and U4326 (N_4326,N_420,N_1868);
nor U4327 (N_4327,N_1619,N_2471);
nand U4328 (N_4328,N_660,N_1781);
nor U4329 (N_4329,N_614,N_591);
or U4330 (N_4330,N_1641,N_1026);
and U4331 (N_4331,N_2471,N_2079);
and U4332 (N_4332,N_346,N_807);
nor U4333 (N_4333,N_202,N_2352);
nor U4334 (N_4334,N_2004,N_1152);
and U4335 (N_4335,N_629,N_1387);
or U4336 (N_4336,N_1560,N_513);
and U4337 (N_4337,N_1214,N_2296);
nor U4338 (N_4338,N_909,N_23);
or U4339 (N_4339,N_1970,N_482);
and U4340 (N_4340,N_2089,N_1945);
nor U4341 (N_4341,N_423,N_2053);
and U4342 (N_4342,N_2347,N_766);
nand U4343 (N_4343,N_1232,N_209);
nor U4344 (N_4344,N_2058,N_860);
nor U4345 (N_4345,N_1568,N_1791);
nand U4346 (N_4346,N_492,N_790);
nor U4347 (N_4347,N_856,N_824);
and U4348 (N_4348,N_142,N_797);
and U4349 (N_4349,N_1135,N_646);
or U4350 (N_4350,N_1398,N_1797);
and U4351 (N_4351,N_1934,N_2143);
or U4352 (N_4352,N_948,N_2028);
or U4353 (N_4353,N_2024,N_2213);
or U4354 (N_4354,N_167,N_1321);
or U4355 (N_4355,N_1215,N_2294);
and U4356 (N_4356,N_34,N_202);
or U4357 (N_4357,N_322,N_2207);
and U4358 (N_4358,N_1451,N_331);
and U4359 (N_4359,N_2010,N_1528);
or U4360 (N_4360,N_1029,N_1132);
or U4361 (N_4361,N_2434,N_2238);
nand U4362 (N_4362,N_366,N_1443);
and U4363 (N_4363,N_787,N_1955);
or U4364 (N_4364,N_59,N_2341);
nand U4365 (N_4365,N_2201,N_2394);
nor U4366 (N_4366,N_2045,N_2083);
nor U4367 (N_4367,N_559,N_1588);
nand U4368 (N_4368,N_1246,N_2056);
nand U4369 (N_4369,N_1721,N_2150);
and U4370 (N_4370,N_1945,N_2389);
nand U4371 (N_4371,N_142,N_66);
nand U4372 (N_4372,N_1736,N_2020);
and U4373 (N_4373,N_1083,N_1902);
and U4374 (N_4374,N_1584,N_1715);
or U4375 (N_4375,N_1531,N_159);
nor U4376 (N_4376,N_1758,N_2472);
nand U4377 (N_4377,N_1820,N_1450);
and U4378 (N_4378,N_472,N_884);
and U4379 (N_4379,N_305,N_1601);
nor U4380 (N_4380,N_1678,N_1689);
nand U4381 (N_4381,N_2011,N_1532);
nor U4382 (N_4382,N_235,N_1586);
nand U4383 (N_4383,N_2465,N_181);
nand U4384 (N_4384,N_608,N_1460);
nand U4385 (N_4385,N_2079,N_950);
nand U4386 (N_4386,N_1755,N_1398);
and U4387 (N_4387,N_40,N_2459);
nand U4388 (N_4388,N_573,N_2409);
and U4389 (N_4389,N_2127,N_186);
nand U4390 (N_4390,N_1249,N_510);
nand U4391 (N_4391,N_1399,N_1743);
and U4392 (N_4392,N_1204,N_1338);
or U4393 (N_4393,N_256,N_179);
and U4394 (N_4394,N_339,N_1299);
nor U4395 (N_4395,N_1280,N_2083);
and U4396 (N_4396,N_1123,N_1426);
xnor U4397 (N_4397,N_645,N_574);
and U4398 (N_4398,N_2194,N_860);
or U4399 (N_4399,N_2080,N_233);
or U4400 (N_4400,N_2198,N_2186);
nand U4401 (N_4401,N_1949,N_706);
or U4402 (N_4402,N_2254,N_2222);
and U4403 (N_4403,N_1088,N_389);
nor U4404 (N_4404,N_962,N_1168);
nor U4405 (N_4405,N_945,N_1202);
and U4406 (N_4406,N_2206,N_1568);
and U4407 (N_4407,N_2031,N_2312);
and U4408 (N_4408,N_2300,N_141);
nand U4409 (N_4409,N_894,N_1107);
and U4410 (N_4410,N_680,N_953);
and U4411 (N_4411,N_2434,N_83);
and U4412 (N_4412,N_2167,N_1614);
and U4413 (N_4413,N_1201,N_679);
or U4414 (N_4414,N_630,N_468);
and U4415 (N_4415,N_1582,N_2254);
nor U4416 (N_4416,N_2072,N_1134);
or U4417 (N_4417,N_821,N_212);
nand U4418 (N_4418,N_667,N_1802);
nand U4419 (N_4419,N_337,N_894);
nor U4420 (N_4420,N_398,N_1004);
nor U4421 (N_4421,N_2100,N_829);
and U4422 (N_4422,N_2107,N_2316);
or U4423 (N_4423,N_1147,N_1415);
nor U4424 (N_4424,N_1126,N_1105);
and U4425 (N_4425,N_258,N_249);
nor U4426 (N_4426,N_1223,N_1757);
or U4427 (N_4427,N_596,N_720);
nand U4428 (N_4428,N_1939,N_1433);
and U4429 (N_4429,N_589,N_795);
nand U4430 (N_4430,N_607,N_716);
nor U4431 (N_4431,N_2267,N_242);
nor U4432 (N_4432,N_2321,N_1492);
nor U4433 (N_4433,N_301,N_1604);
nor U4434 (N_4434,N_1405,N_1339);
and U4435 (N_4435,N_2484,N_1659);
or U4436 (N_4436,N_2184,N_1783);
nor U4437 (N_4437,N_1223,N_1165);
and U4438 (N_4438,N_1963,N_21);
nand U4439 (N_4439,N_521,N_423);
and U4440 (N_4440,N_689,N_2171);
nand U4441 (N_4441,N_1069,N_1640);
nor U4442 (N_4442,N_1071,N_1681);
and U4443 (N_4443,N_1198,N_791);
nand U4444 (N_4444,N_1377,N_1211);
nand U4445 (N_4445,N_1504,N_397);
or U4446 (N_4446,N_424,N_192);
nand U4447 (N_4447,N_1813,N_1165);
and U4448 (N_4448,N_606,N_2202);
nor U4449 (N_4449,N_1585,N_368);
nand U4450 (N_4450,N_2116,N_963);
nand U4451 (N_4451,N_252,N_87);
and U4452 (N_4452,N_859,N_1481);
or U4453 (N_4453,N_1191,N_217);
and U4454 (N_4454,N_2146,N_83);
and U4455 (N_4455,N_346,N_2154);
nand U4456 (N_4456,N_1916,N_1022);
or U4457 (N_4457,N_1590,N_1723);
or U4458 (N_4458,N_1632,N_571);
nand U4459 (N_4459,N_857,N_22);
and U4460 (N_4460,N_1034,N_173);
and U4461 (N_4461,N_1930,N_75);
nor U4462 (N_4462,N_626,N_2089);
and U4463 (N_4463,N_2178,N_1626);
and U4464 (N_4464,N_1876,N_1906);
nand U4465 (N_4465,N_831,N_342);
nand U4466 (N_4466,N_1088,N_44);
nor U4467 (N_4467,N_743,N_2197);
nand U4468 (N_4468,N_2245,N_1232);
or U4469 (N_4469,N_608,N_1904);
xor U4470 (N_4470,N_440,N_1388);
xnor U4471 (N_4471,N_838,N_1596);
nor U4472 (N_4472,N_309,N_1428);
nand U4473 (N_4473,N_1518,N_1475);
or U4474 (N_4474,N_237,N_479);
nand U4475 (N_4475,N_793,N_421);
or U4476 (N_4476,N_2190,N_1215);
and U4477 (N_4477,N_14,N_1878);
nor U4478 (N_4478,N_925,N_50);
and U4479 (N_4479,N_2478,N_1325);
nand U4480 (N_4480,N_1242,N_758);
or U4481 (N_4481,N_2105,N_1604);
and U4482 (N_4482,N_1343,N_731);
nor U4483 (N_4483,N_1801,N_1008);
or U4484 (N_4484,N_963,N_683);
nor U4485 (N_4485,N_2104,N_2049);
nor U4486 (N_4486,N_1903,N_956);
nor U4487 (N_4487,N_1510,N_1994);
nand U4488 (N_4488,N_2487,N_1701);
or U4489 (N_4489,N_1428,N_654);
or U4490 (N_4490,N_366,N_1680);
and U4491 (N_4491,N_528,N_1748);
nand U4492 (N_4492,N_2222,N_1082);
nand U4493 (N_4493,N_1722,N_1266);
and U4494 (N_4494,N_29,N_1016);
nand U4495 (N_4495,N_1912,N_2339);
nor U4496 (N_4496,N_2359,N_669);
and U4497 (N_4497,N_50,N_690);
nand U4498 (N_4498,N_2069,N_935);
nand U4499 (N_4499,N_246,N_1431);
or U4500 (N_4500,N_1523,N_1869);
nand U4501 (N_4501,N_1810,N_381);
or U4502 (N_4502,N_939,N_38);
nand U4503 (N_4503,N_1095,N_1869);
or U4504 (N_4504,N_2011,N_1903);
nor U4505 (N_4505,N_173,N_2242);
nand U4506 (N_4506,N_999,N_54);
or U4507 (N_4507,N_310,N_1011);
nor U4508 (N_4508,N_666,N_125);
nor U4509 (N_4509,N_328,N_482);
nor U4510 (N_4510,N_621,N_1683);
nand U4511 (N_4511,N_2370,N_842);
nor U4512 (N_4512,N_60,N_16);
or U4513 (N_4513,N_85,N_1600);
nand U4514 (N_4514,N_243,N_840);
nor U4515 (N_4515,N_318,N_2190);
and U4516 (N_4516,N_2442,N_1251);
nand U4517 (N_4517,N_1606,N_1607);
or U4518 (N_4518,N_762,N_746);
and U4519 (N_4519,N_591,N_135);
or U4520 (N_4520,N_1430,N_1148);
nor U4521 (N_4521,N_2316,N_1274);
nand U4522 (N_4522,N_675,N_47);
and U4523 (N_4523,N_80,N_1062);
nand U4524 (N_4524,N_1347,N_1779);
or U4525 (N_4525,N_485,N_330);
or U4526 (N_4526,N_1306,N_981);
or U4527 (N_4527,N_1758,N_895);
nand U4528 (N_4528,N_2366,N_2033);
nand U4529 (N_4529,N_313,N_1841);
nor U4530 (N_4530,N_2092,N_1307);
and U4531 (N_4531,N_1302,N_1429);
nor U4532 (N_4532,N_1460,N_335);
nand U4533 (N_4533,N_422,N_1902);
and U4534 (N_4534,N_1774,N_976);
nor U4535 (N_4535,N_67,N_369);
and U4536 (N_4536,N_668,N_2062);
nand U4537 (N_4537,N_1457,N_681);
nand U4538 (N_4538,N_1078,N_891);
and U4539 (N_4539,N_944,N_1144);
and U4540 (N_4540,N_1048,N_571);
or U4541 (N_4541,N_1405,N_1279);
nand U4542 (N_4542,N_890,N_251);
and U4543 (N_4543,N_1786,N_1108);
nor U4544 (N_4544,N_851,N_760);
or U4545 (N_4545,N_1085,N_791);
nand U4546 (N_4546,N_473,N_1172);
nand U4547 (N_4547,N_1392,N_1272);
nand U4548 (N_4548,N_965,N_936);
or U4549 (N_4549,N_1704,N_1175);
nor U4550 (N_4550,N_1806,N_2411);
nor U4551 (N_4551,N_456,N_2097);
xor U4552 (N_4552,N_231,N_1863);
nor U4553 (N_4553,N_265,N_1346);
and U4554 (N_4554,N_1359,N_481);
or U4555 (N_4555,N_978,N_2297);
and U4556 (N_4556,N_1467,N_1801);
nor U4557 (N_4557,N_824,N_1779);
or U4558 (N_4558,N_273,N_580);
or U4559 (N_4559,N_1316,N_1203);
nand U4560 (N_4560,N_1907,N_268);
nor U4561 (N_4561,N_1386,N_190);
nand U4562 (N_4562,N_2411,N_1371);
and U4563 (N_4563,N_290,N_1986);
or U4564 (N_4564,N_2498,N_62);
or U4565 (N_4565,N_591,N_1574);
and U4566 (N_4566,N_2312,N_2265);
nand U4567 (N_4567,N_2485,N_55);
and U4568 (N_4568,N_1709,N_1116);
nand U4569 (N_4569,N_1989,N_2219);
nor U4570 (N_4570,N_1708,N_2224);
or U4571 (N_4571,N_1147,N_875);
and U4572 (N_4572,N_353,N_1855);
or U4573 (N_4573,N_2354,N_2430);
nand U4574 (N_4574,N_2379,N_239);
nor U4575 (N_4575,N_353,N_909);
nand U4576 (N_4576,N_519,N_1850);
and U4577 (N_4577,N_692,N_1453);
nor U4578 (N_4578,N_1974,N_1762);
nor U4579 (N_4579,N_465,N_576);
nor U4580 (N_4580,N_1607,N_1770);
or U4581 (N_4581,N_1286,N_1959);
nor U4582 (N_4582,N_64,N_1526);
and U4583 (N_4583,N_1471,N_1436);
nand U4584 (N_4584,N_754,N_1714);
nor U4585 (N_4585,N_876,N_342);
or U4586 (N_4586,N_0,N_1899);
or U4587 (N_4587,N_140,N_62);
nor U4588 (N_4588,N_1759,N_938);
or U4589 (N_4589,N_626,N_2094);
nor U4590 (N_4590,N_1440,N_437);
and U4591 (N_4591,N_513,N_254);
nor U4592 (N_4592,N_1899,N_1191);
or U4593 (N_4593,N_2251,N_82);
and U4594 (N_4594,N_1354,N_1531);
and U4595 (N_4595,N_885,N_2034);
or U4596 (N_4596,N_2250,N_1945);
and U4597 (N_4597,N_1801,N_238);
or U4598 (N_4598,N_118,N_525);
or U4599 (N_4599,N_1123,N_607);
or U4600 (N_4600,N_180,N_767);
nor U4601 (N_4601,N_1754,N_664);
nand U4602 (N_4602,N_478,N_1902);
nor U4603 (N_4603,N_1834,N_990);
nand U4604 (N_4604,N_10,N_1699);
and U4605 (N_4605,N_1466,N_2232);
nor U4606 (N_4606,N_88,N_1465);
or U4607 (N_4607,N_1416,N_1659);
or U4608 (N_4608,N_2322,N_2345);
and U4609 (N_4609,N_1234,N_388);
and U4610 (N_4610,N_1451,N_1255);
nand U4611 (N_4611,N_801,N_654);
nor U4612 (N_4612,N_2376,N_139);
nand U4613 (N_4613,N_1300,N_808);
and U4614 (N_4614,N_143,N_1387);
nor U4615 (N_4615,N_253,N_901);
nor U4616 (N_4616,N_791,N_1357);
or U4617 (N_4617,N_1749,N_1052);
or U4618 (N_4618,N_1593,N_106);
nor U4619 (N_4619,N_2462,N_2344);
nand U4620 (N_4620,N_393,N_2100);
or U4621 (N_4621,N_1486,N_1792);
and U4622 (N_4622,N_862,N_1094);
nor U4623 (N_4623,N_173,N_864);
nor U4624 (N_4624,N_581,N_1739);
nand U4625 (N_4625,N_233,N_1731);
or U4626 (N_4626,N_2109,N_2363);
nand U4627 (N_4627,N_285,N_2435);
nand U4628 (N_4628,N_1969,N_123);
or U4629 (N_4629,N_1717,N_1080);
and U4630 (N_4630,N_793,N_1098);
or U4631 (N_4631,N_2427,N_2095);
and U4632 (N_4632,N_68,N_1051);
and U4633 (N_4633,N_1684,N_1047);
and U4634 (N_4634,N_1926,N_361);
nand U4635 (N_4635,N_1680,N_551);
and U4636 (N_4636,N_1001,N_1331);
or U4637 (N_4637,N_1494,N_1650);
or U4638 (N_4638,N_473,N_1580);
nand U4639 (N_4639,N_193,N_251);
or U4640 (N_4640,N_2399,N_1069);
and U4641 (N_4641,N_724,N_1675);
nor U4642 (N_4642,N_79,N_997);
nand U4643 (N_4643,N_1545,N_1686);
and U4644 (N_4644,N_1729,N_1426);
nand U4645 (N_4645,N_1307,N_504);
or U4646 (N_4646,N_2012,N_2382);
or U4647 (N_4647,N_2154,N_1927);
nand U4648 (N_4648,N_888,N_752);
and U4649 (N_4649,N_466,N_93);
nor U4650 (N_4650,N_20,N_1605);
and U4651 (N_4651,N_370,N_1095);
and U4652 (N_4652,N_1937,N_1784);
and U4653 (N_4653,N_684,N_1398);
or U4654 (N_4654,N_1810,N_1822);
nor U4655 (N_4655,N_862,N_2424);
nand U4656 (N_4656,N_734,N_2314);
or U4657 (N_4657,N_2200,N_737);
or U4658 (N_4658,N_494,N_1345);
or U4659 (N_4659,N_1277,N_258);
or U4660 (N_4660,N_1426,N_13);
or U4661 (N_4661,N_2376,N_2341);
nor U4662 (N_4662,N_1427,N_1947);
or U4663 (N_4663,N_1443,N_2300);
nor U4664 (N_4664,N_649,N_1407);
nand U4665 (N_4665,N_1850,N_1632);
nand U4666 (N_4666,N_371,N_1156);
and U4667 (N_4667,N_1605,N_2157);
nor U4668 (N_4668,N_317,N_2052);
nand U4669 (N_4669,N_265,N_1558);
nor U4670 (N_4670,N_2442,N_1760);
nor U4671 (N_4671,N_777,N_996);
nand U4672 (N_4672,N_194,N_1849);
or U4673 (N_4673,N_834,N_1309);
nor U4674 (N_4674,N_1549,N_2324);
nor U4675 (N_4675,N_1117,N_372);
nand U4676 (N_4676,N_1290,N_2281);
or U4677 (N_4677,N_1692,N_668);
nand U4678 (N_4678,N_193,N_1432);
or U4679 (N_4679,N_2411,N_2261);
nor U4680 (N_4680,N_965,N_66);
nor U4681 (N_4681,N_2209,N_1290);
and U4682 (N_4682,N_565,N_798);
xor U4683 (N_4683,N_448,N_877);
and U4684 (N_4684,N_666,N_1929);
and U4685 (N_4685,N_925,N_1428);
or U4686 (N_4686,N_1666,N_962);
and U4687 (N_4687,N_1822,N_198);
nor U4688 (N_4688,N_409,N_2);
and U4689 (N_4689,N_1307,N_1155);
nor U4690 (N_4690,N_2238,N_1113);
nand U4691 (N_4691,N_1073,N_2218);
and U4692 (N_4692,N_1444,N_1128);
nor U4693 (N_4693,N_1336,N_848);
nand U4694 (N_4694,N_1564,N_34);
or U4695 (N_4695,N_332,N_323);
or U4696 (N_4696,N_400,N_488);
nor U4697 (N_4697,N_1495,N_879);
and U4698 (N_4698,N_1046,N_751);
nand U4699 (N_4699,N_428,N_659);
and U4700 (N_4700,N_931,N_2371);
nand U4701 (N_4701,N_10,N_1228);
and U4702 (N_4702,N_231,N_2074);
and U4703 (N_4703,N_286,N_1965);
and U4704 (N_4704,N_1059,N_2034);
nand U4705 (N_4705,N_597,N_729);
nand U4706 (N_4706,N_1497,N_2022);
nor U4707 (N_4707,N_925,N_834);
nand U4708 (N_4708,N_1478,N_1957);
and U4709 (N_4709,N_81,N_182);
nor U4710 (N_4710,N_1813,N_1984);
xnor U4711 (N_4711,N_1475,N_676);
nor U4712 (N_4712,N_1576,N_1320);
and U4713 (N_4713,N_1712,N_1227);
and U4714 (N_4714,N_745,N_1054);
nand U4715 (N_4715,N_700,N_1732);
and U4716 (N_4716,N_700,N_1414);
or U4717 (N_4717,N_2259,N_2449);
nand U4718 (N_4718,N_1688,N_702);
or U4719 (N_4719,N_996,N_1254);
xor U4720 (N_4720,N_892,N_2067);
or U4721 (N_4721,N_63,N_2358);
or U4722 (N_4722,N_751,N_2179);
or U4723 (N_4723,N_2281,N_2024);
and U4724 (N_4724,N_239,N_1862);
nand U4725 (N_4725,N_617,N_127);
nand U4726 (N_4726,N_333,N_1396);
nor U4727 (N_4727,N_1724,N_2021);
and U4728 (N_4728,N_95,N_1210);
nor U4729 (N_4729,N_186,N_1708);
nand U4730 (N_4730,N_4,N_1532);
nand U4731 (N_4731,N_88,N_1599);
and U4732 (N_4732,N_2471,N_1378);
or U4733 (N_4733,N_1243,N_238);
or U4734 (N_4734,N_2352,N_317);
and U4735 (N_4735,N_584,N_1331);
and U4736 (N_4736,N_2310,N_229);
or U4737 (N_4737,N_1551,N_61);
or U4738 (N_4738,N_525,N_812);
and U4739 (N_4739,N_1436,N_1487);
or U4740 (N_4740,N_59,N_1514);
and U4741 (N_4741,N_171,N_785);
nand U4742 (N_4742,N_1029,N_1208);
or U4743 (N_4743,N_1681,N_783);
nand U4744 (N_4744,N_2324,N_1879);
nand U4745 (N_4745,N_2433,N_537);
and U4746 (N_4746,N_2212,N_1934);
and U4747 (N_4747,N_201,N_2452);
nor U4748 (N_4748,N_1505,N_2129);
and U4749 (N_4749,N_1400,N_1793);
and U4750 (N_4750,N_589,N_1395);
and U4751 (N_4751,N_1720,N_285);
or U4752 (N_4752,N_2450,N_660);
or U4753 (N_4753,N_1521,N_1069);
nor U4754 (N_4754,N_460,N_2079);
and U4755 (N_4755,N_439,N_1057);
or U4756 (N_4756,N_591,N_944);
nor U4757 (N_4757,N_789,N_1222);
nand U4758 (N_4758,N_1758,N_1596);
and U4759 (N_4759,N_400,N_2042);
nor U4760 (N_4760,N_2103,N_403);
or U4761 (N_4761,N_1716,N_820);
nand U4762 (N_4762,N_1717,N_1548);
or U4763 (N_4763,N_331,N_117);
nand U4764 (N_4764,N_312,N_1102);
or U4765 (N_4765,N_2015,N_1667);
or U4766 (N_4766,N_427,N_577);
or U4767 (N_4767,N_1042,N_2468);
nor U4768 (N_4768,N_2183,N_748);
and U4769 (N_4769,N_335,N_580);
nand U4770 (N_4770,N_898,N_1938);
and U4771 (N_4771,N_561,N_793);
and U4772 (N_4772,N_971,N_1400);
nor U4773 (N_4773,N_47,N_1657);
and U4774 (N_4774,N_1660,N_552);
and U4775 (N_4775,N_2233,N_221);
or U4776 (N_4776,N_1584,N_1222);
nand U4777 (N_4777,N_949,N_2088);
nand U4778 (N_4778,N_814,N_966);
and U4779 (N_4779,N_2485,N_1759);
and U4780 (N_4780,N_547,N_2178);
and U4781 (N_4781,N_1574,N_1651);
nand U4782 (N_4782,N_2252,N_1311);
and U4783 (N_4783,N_2225,N_630);
nand U4784 (N_4784,N_659,N_820);
nor U4785 (N_4785,N_489,N_1983);
and U4786 (N_4786,N_261,N_1733);
nand U4787 (N_4787,N_1692,N_2085);
or U4788 (N_4788,N_952,N_2461);
and U4789 (N_4789,N_2303,N_1157);
and U4790 (N_4790,N_1837,N_1748);
nor U4791 (N_4791,N_195,N_1602);
nor U4792 (N_4792,N_565,N_730);
or U4793 (N_4793,N_1205,N_1772);
nand U4794 (N_4794,N_352,N_2245);
nand U4795 (N_4795,N_986,N_1335);
and U4796 (N_4796,N_521,N_2163);
and U4797 (N_4797,N_2278,N_2119);
or U4798 (N_4798,N_511,N_2379);
nand U4799 (N_4799,N_1801,N_2426);
or U4800 (N_4800,N_415,N_2496);
and U4801 (N_4801,N_1723,N_2233);
and U4802 (N_4802,N_794,N_1399);
nor U4803 (N_4803,N_749,N_1179);
and U4804 (N_4804,N_1666,N_697);
or U4805 (N_4805,N_2167,N_1533);
nand U4806 (N_4806,N_1182,N_2230);
nor U4807 (N_4807,N_68,N_1988);
nor U4808 (N_4808,N_2017,N_2382);
or U4809 (N_4809,N_1920,N_169);
and U4810 (N_4810,N_1811,N_1678);
and U4811 (N_4811,N_987,N_2456);
or U4812 (N_4812,N_417,N_782);
or U4813 (N_4813,N_776,N_2144);
or U4814 (N_4814,N_2094,N_2311);
or U4815 (N_4815,N_2370,N_355);
nor U4816 (N_4816,N_859,N_1055);
nand U4817 (N_4817,N_2100,N_669);
or U4818 (N_4818,N_2449,N_942);
or U4819 (N_4819,N_865,N_896);
nand U4820 (N_4820,N_1080,N_2232);
xnor U4821 (N_4821,N_1439,N_1367);
and U4822 (N_4822,N_1643,N_2031);
or U4823 (N_4823,N_1160,N_2358);
nand U4824 (N_4824,N_2475,N_1023);
or U4825 (N_4825,N_2050,N_923);
nor U4826 (N_4826,N_2336,N_525);
nor U4827 (N_4827,N_994,N_205);
or U4828 (N_4828,N_1885,N_1694);
and U4829 (N_4829,N_2266,N_866);
or U4830 (N_4830,N_569,N_1607);
nor U4831 (N_4831,N_2042,N_998);
nand U4832 (N_4832,N_626,N_1476);
nand U4833 (N_4833,N_30,N_2124);
nor U4834 (N_4834,N_1183,N_2032);
nor U4835 (N_4835,N_1602,N_1000);
nor U4836 (N_4836,N_2265,N_140);
or U4837 (N_4837,N_411,N_2326);
nor U4838 (N_4838,N_2279,N_607);
or U4839 (N_4839,N_1646,N_85);
and U4840 (N_4840,N_246,N_245);
nor U4841 (N_4841,N_1906,N_8);
or U4842 (N_4842,N_1393,N_1867);
and U4843 (N_4843,N_321,N_1055);
nor U4844 (N_4844,N_2158,N_1716);
nand U4845 (N_4845,N_1906,N_1738);
and U4846 (N_4846,N_849,N_1505);
and U4847 (N_4847,N_1822,N_2366);
and U4848 (N_4848,N_1219,N_2322);
or U4849 (N_4849,N_505,N_2125);
nand U4850 (N_4850,N_2197,N_592);
nand U4851 (N_4851,N_723,N_2398);
nor U4852 (N_4852,N_1274,N_1302);
or U4853 (N_4853,N_2023,N_1417);
nor U4854 (N_4854,N_20,N_650);
and U4855 (N_4855,N_953,N_618);
nand U4856 (N_4856,N_364,N_174);
nor U4857 (N_4857,N_945,N_2363);
or U4858 (N_4858,N_1406,N_861);
nor U4859 (N_4859,N_964,N_1309);
and U4860 (N_4860,N_1309,N_2149);
nand U4861 (N_4861,N_2443,N_1694);
and U4862 (N_4862,N_840,N_1853);
or U4863 (N_4863,N_1310,N_1804);
and U4864 (N_4864,N_2084,N_2188);
nand U4865 (N_4865,N_2197,N_1957);
or U4866 (N_4866,N_836,N_968);
nor U4867 (N_4867,N_1761,N_1421);
nand U4868 (N_4868,N_1103,N_894);
and U4869 (N_4869,N_387,N_1424);
nor U4870 (N_4870,N_769,N_876);
or U4871 (N_4871,N_1447,N_1115);
nor U4872 (N_4872,N_551,N_2383);
and U4873 (N_4873,N_1797,N_1721);
or U4874 (N_4874,N_1582,N_293);
or U4875 (N_4875,N_2108,N_803);
nor U4876 (N_4876,N_2073,N_1031);
or U4877 (N_4877,N_125,N_1208);
and U4878 (N_4878,N_302,N_2455);
nand U4879 (N_4879,N_840,N_1227);
or U4880 (N_4880,N_1133,N_1903);
or U4881 (N_4881,N_523,N_1352);
and U4882 (N_4882,N_427,N_2095);
nor U4883 (N_4883,N_1141,N_1272);
and U4884 (N_4884,N_2043,N_334);
and U4885 (N_4885,N_853,N_2441);
or U4886 (N_4886,N_173,N_1193);
nor U4887 (N_4887,N_402,N_1245);
or U4888 (N_4888,N_2013,N_1756);
or U4889 (N_4889,N_2409,N_1383);
or U4890 (N_4890,N_354,N_43);
nor U4891 (N_4891,N_874,N_300);
and U4892 (N_4892,N_105,N_338);
and U4893 (N_4893,N_473,N_1171);
nor U4894 (N_4894,N_1439,N_585);
or U4895 (N_4895,N_556,N_700);
nor U4896 (N_4896,N_60,N_1939);
and U4897 (N_4897,N_95,N_2359);
nand U4898 (N_4898,N_2045,N_1906);
nor U4899 (N_4899,N_2145,N_845);
nor U4900 (N_4900,N_1595,N_877);
or U4901 (N_4901,N_1122,N_1261);
and U4902 (N_4902,N_393,N_248);
nand U4903 (N_4903,N_1040,N_1566);
nor U4904 (N_4904,N_1612,N_841);
nor U4905 (N_4905,N_2028,N_1551);
nand U4906 (N_4906,N_1507,N_1712);
and U4907 (N_4907,N_591,N_2412);
or U4908 (N_4908,N_687,N_630);
or U4909 (N_4909,N_265,N_531);
nand U4910 (N_4910,N_2151,N_1356);
nand U4911 (N_4911,N_62,N_476);
or U4912 (N_4912,N_1616,N_11);
nor U4913 (N_4913,N_2406,N_1289);
and U4914 (N_4914,N_1619,N_1898);
and U4915 (N_4915,N_389,N_427);
nor U4916 (N_4916,N_1100,N_1089);
nand U4917 (N_4917,N_1313,N_1012);
or U4918 (N_4918,N_1532,N_1528);
or U4919 (N_4919,N_1500,N_51);
xor U4920 (N_4920,N_2294,N_1893);
or U4921 (N_4921,N_2125,N_1675);
nor U4922 (N_4922,N_943,N_1857);
and U4923 (N_4923,N_23,N_527);
or U4924 (N_4924,N_1863,N_1421);
and U4925 (N_4925,N_1934,N_2449);
nor U4926 (N_4926,N_1477,N_1774);
nor U4927 (N_4927,N_2150,N_1443);
nor U4928 (N_4928,N_1044,N_1723);
nor U4929 (N_4929,N_2364,N_110);
nand U4930 (N_4930,N_841,N_1308);
nand U4931 (N_4931,N_610,N_1623);
nor U4932 (N_4932,N_1567,N_1727);
xnor U4933 (N_4933,N_184,N_2287);
nor U4934 (N_4934,N_768,N_1759);
nor U4935 (N_4935,N_23,N_1706);
nand U4936 (N_4936,N_1027,N_2347);
nor U4937 (N_4937,N_1863,N_612);
and U4938 (N_4938,N_892,N_694);
nor U4939 (N_4939,N_1485,N_1502);
nor U4940 (N_4940,N_2378,N_1882);
nand U4941 (N_4941,N_46,N_289);
nand U4942 (N_4942,N_2275,N_2033);
and U4943 (N_4943,N_927,N_892);
or U4944 (N_4944,N_287,N_836);
nor U4945 (N_4945,N_1379,N_871);
nand U4946 (N_4946,N_1720,N_2402);
nor U4947 (N_4947,N_383,N_1555);
and U4948 (N_4948,N_449,N_1092);
or U4949 (N_4949,N_398,N_1080);
and U4950 (N_4950,N_2115,N_357);
nor U4951 (N_4951,N_2076,N_1824);
or U4952 (N_4952,N_2225,N_2327);
nand U4953 (N_4953,N_2303,N_1344);
or U4954 (N_4954,N_1071,N_1052);
nand U4955 (N_4955,N_1239,N_1432);
and U4956 (N_4956,N_238,N_2226);
xor U4957 (N_4957,N_291,N_301);
nor U4958 (N_4958,N_1106,N_786);
and U4959 (N_4959,N_1103,N_1600);
or U4960 (N_4960,N_407,N_1437);
or U4961 (N_4961,N_2232,N_1715);
nand U4962 (N_4962,N_399,N_1606);
nand U4963 (N_4963,N_2116,N_137);
or U4964 (N_4964,N_1895,N_479);
nor U4965 (N_4965,N_2360,N_2236);
nand U4966 (N_4966,N_1481,N_1284);
nand U4967 (N_4967,N_931,N_948);
and U4968 (N_4968,N_2323,N_1688);
or U4969 (N_4969,N_95,N_1173);
nand U4970 (N_4970,N_655,N_286);
or U4971 (N_4971,N_1254,N_1352);
nor U4972 (N_4972,N_2193,N_2002);
nand U4973 (N_4973,N_3,N_14);
nor U4974 (N_4974,N_1139,N_2);
nand U4975 (N_4975,N_1134,N_809);
and U4976 (N_4976,N_2272,N_1035);
and U4977 (N_4977,N_504,N_2191);
or U4978 (N_4978,N_1461,N_1270);
or U4979 (N_4979,N_891,N_676);
and U4980 (N_4980,N_51,N_1357);
and U4981 (N_4981,N_832,N_407);
or U4982 (N_4982,N_1179,N_2136);
and U4983 (N_4983,N_1163,N_1249);
nor U4984 (N_4984,N_1176,N_792);
and U4985 (N_4985,N_1000,N_2472);
and U4986 (N_4986,N_580,N_1737);
or U4987 (N_4987,N_2320,N_765);
and U4988 (N_4988,N_971,N_1137);
nand U4989 (N_4989,N_458,N_2310);
or U4990 (N_4990,N_1363,N_604);
or U4991 (N_4991,N_2126,N_2386);
and U4992 (N_4992,N_678,N_2443);
nor U4993 (N_4993,N_2125,N_1057);
nand U4994 (N_4994,N_671,N_1645);
nand U4995 (N_4995,N_1216,N_75);
and U4996 (N_4996,N_231,N_1191);
nand U4997 (N_4997,N_85,N_1161);
and U4998 (N_4998,N_1804,N_1523);
or U4999 (N_4999,N_932,N_1686);
xnor UO_0 (O_0,N_3413,N_3366);
and UO_1 (O_1,N_4259,N_3460);
nand UO_2 (O_2,N_3383,N_3162);
nor UO_3 (O_3,N_3373,N_3304);
nand UO_4 (O_4,N_3495,N_4574);
or UO_5 (O_5,N_3338,N_3967);
nand UO_6 (O_6,N_4825,N_4823);
nor UO_7 (O_7,N_3830,N_2762);
nand UO_8 (O_8,N_3783,N_4713);
nor UO_9 (O_9,N_3928,N_4610);
nor UO_10 (O_10,N_3656,N_4937);
nor UO_11 (O_11,N_4048,N_3417);
or UO_12 (O_12,N_4111,N_2556);
nor UO_13 (O_13,N_3280,N_2771);
and UO_14 (O_14,N_4777,N_2934);
nor UO_15 (O_15,N_4763,N_3119);
nor UO_16 (O_16,N_2772,N_3248);
or UO_17 (O_17,N_2877,N_4576);
nand UO_18 (O_18,N_3621,N_3356);
or UO_19 (O_19,N_3147,N_3259);
nor UO_20 (O_20,N_4178,N_2566);
and UO_21 (O_21,N_4278,N_2780);
nor UO_22 (O_22,N_2828,N_2844);
nand UO_23 (O_23,N_3051,N_2548);
or UO_24 (O_24,N_2702,N_3066);
and UO_25 (O_25,N_4025,N_4566);
nand UO_26 (O_26,N_3952,N_4829);
nand UO_27 (O_27,N_3812,N_2547);
nand UO_28 (O_28,N_2581,N_4944);
nor UO_29 (O_29,N_4607,N_4448);
nor UO_30 (O_30,N_3567,N_3950);
or UO_31 (O_31,N_3296,N_4555);
xnor UO_32 (O_32,N_4244,N_4252);
and UO_33 (O_33,N_2748,N_4942);
and UO_34 (O_34,N_4630,N_4276);
nand UO_35 (O_35,N_4911,N_4220);
nor UO_36 (O_36,N_4563,N_4442);
or UO_37 (O_37,N_3687,N_3480);
or UO_38 (O_38,N_3266,N_3896);
or UO_39 (O_39,N_4005,N_4208);
and UO_40 (O_40,N_3419,N_2788);
or UO_41 (O_41,N_3968,N_2815);
nand UO_42 (O_42,N_3990,N_4867);
nand UO_43 (O_43,N_3841,N_3702);
nor UO_44 (O_44,N_4073,N_4894);
or UO_45 (O_45,N_3022,N_3879);
nor UO_46 (O_46,N_4933,N_2727);
or UO_47 (O_47,N_4134,N_3392);
nand UO_48 (O_48,N_4026,N_4965);
nor UO_49 (O_49,N_4372,N_3037);
and UO_50 (O_50,N_4461,N_4092);
nand UO_51 (O_51,N_3661,N_2678);
nor UO_52 (O_52,N_3007,N_2565);
nand UO_53 (O_53,N_3239,N_4104);
and UO_54 (O_54,N_3314,N_4217);
xnor UO_55 (O_55,N_3605,N_2823);
nor UO_56 (O_56,N_4664,N_3225);
nor UO_57 (O_57,N_3320,N_3258);
and UO_58 (O_58,N_3664,N_4975);
and UO_59 (O_59,N_2918,N_3944);
and UO_60 (O_60,N_4401,N_3512);
or UO_61 (O_61,N_3900,N_4527);
and UO_62 (O_62,N_4248,N_3298);
nand UO_63 (O_63,N_4914,N_4872);
or UO_64 (O_64,N_3433,N_4227);
nand UO_65 (O_65,N_3708,N_4019);
or UO_66 (O_66,N_2973,N_4055);
nor UO_67 (O_67,N_3671,N_2652);
and UO_68 (O_68,N_3167,N_2800);
or UO_69 (O_69,N_3573,N_3510);
nor UO_70 (O_70,N_4819,N_3332);
and UO_71 (O_71,N_3541,N_4558);
nand UO_72 (O_72,N_2770,N_3485);
or UO_73 (O_73,N_2980,N_3980);
and UO_74 (O_74,N_3172,N_4008);
nand UO_75 (O_75,N_4636,N_2990);
and UO_76 (O_76,N_2550,N_4185);
nand UO_77 (O_77,N_3279,N_3936);
nor UO_78 (O_78,N_2816,N_4988);
nand UO_79 (O_79,N_4844,N_3721);
nand UO_80 (O_80,N_4407,N_3659);
nand UO_81 (O_81,N_4733,N_3842);
nand UO_82 (O_82,N_2578,N_3355);
nand UO_83 (O_83,N_2878,N_4833);
and UO_84 (O_84,N_4483,N_2847);
nor UO_85 (O_85,N_4628,N_4960);
nand UO_86 (O_86,N_2537,N_3459);
and UO_87 (O_87,N_4583,N_4856);
and UO_88 (O_88,N_4868,N_3668);
nor UO_89 (O_89,N_3566,N_2975);
nand UO_90 (O_90,N_4826,N_3779);
nor UO_91 (O_91,N_2579,N_2608);
or UO_92 (O_92,N_4299,N_3041);
and UO_93 (O_93,N_3301,N_4486);
nand UO_94 (O_94,N_3973,N_4759);
and UO_95 (O_95,N_4804,N_4052);
nand UO_96 (O_96,N_3534,N_3499);
and UO_97 (O_97,N_3473,N_3477);
nor UO_98 (O_98,N_3773,N_4509);
nor UO_99 (O_99,N_3211,N_4041);
and UO_100 (O_100,N_4705,N_3268);
nor UO_101 (O_101,N_2759,N_4866);
nor UO_102 (O_102,N_2955,N_4155);
or UO_103 (O_103,N_3453,N_4112);
and UO_104 (O_104,N_3641,N_4556);
nand UO_105 (O_105,N_2688,N_4141);
nor UO_106 (O_106,N_4586,N_3244);
nor UO_107 (O_107,N_3583,N_4753);
nand UO_108 (O_108,N_2970,N_4143);
or UO_109 (O_109,N_3291,N_3337);
nor UO_110 (O_110,N_3029,N_2611);
or UO_111 (O_111,N_3847,N_3798);
nor UO_112 (O_112,N_4645,N_2840);
nand UO_113 (O_113,N_3427,N_4201);
and UO_114 (O_114,N_4694,N_3504);
nand UO_115 (O_115,N_3023,N_3262);
nand UO_116 (O_116,N_2852,N_4709);
or UO_117 (O_117,N_4156,N_2601);
or UO_118 (O_118,N_3745,N_4100);
nor UO_119 (O_119,N_4751,N_4375);
nand UO_120 (O_120,N_3974,N_4686);
nand UO_121 (O_121,N_3113,N_4462);
nor UO_122 (O_122,N_2791,N_4166);
or UO_123 (O_123,N_4885,N_4243);
nor UO_124 (O_124,N_4888,N_3331);
and UO_125 (O_125,N_3806,N_3249);
and UO_126 (O_126,N_2853,N_3053);
and UO_127 (O_127,N_4369,N_3892);
nand UO_128 (O_128,N_4828,N_3185);
xor UO_129 (O_129,N_2783,N_4848);
or UO_130 (O_130,N_4905,N_3620);
nand UO_131 (O_131,N_3908,N_4876);
or UO_132 (O_132,N_2781,N_3109);
and UO_133 (O_133,N_3749,N_3843);
and UO_134 (O_134,N_3025,N_4880);
nor UO_135 (O_135,N_4409,N_2982);
nor UO_136 (O_136,N_4608,N_4291);
or UO_137 (O_137,N_4096,N_3649);
and UO_138 (O_138,N_4993,N_4006);
and UO_139 (O_139,N_4510,N_3505);
or UO_140 (O_140,N_4487,N_2965);
nand UO_141 (O_141,N_2939,N_4801);
and UO_142 (O_142,N_2829,N_3329);
nor UO_143 (O_143,N_3177,N_2966);
nor UO_144 (O_144,N_4320,N_3002);
and UO_145 (O_145,N_3133,N_2551);
or UO_146 (O_146,N_3529,N_3275);
and UO_147 (O_147,N_4697,N_4758);
nand UO_148 (O_148,N_2956,N_4275);
or UO_149 (O_149,N_2804,N_2924);
nand UO_150 (O_150,N_4870,N_4183);
or UO_151 (O_151,N_4174,N_3179);
nand UO_152 (O_152,N_4233,N_4927);
nor UO_153 (O_153,N_4429,N_3619);
and UO_154 (O_154,N_3568,N_2807);
and UO_155 (O_155,N_4218,N_3956);
nand UO_156 (O_156,N_2763,N_4700);
and UO_157 (O_157,N_4050,N_3009);
or UO_158 (O_158,N_3100,N_3738);
nand UO_159 (O_159,N_3288,N_4367);
nor UO_160 (O_160,N_4648,N_3533);
and UO_161 (O_161,N_3891,N_4540);
or UO_162 (O_162,N_2715,N_4752);
or UO_163 (O_163,N_3508,N_4355);
or UO_164 (O_164,N_4443,N_2898);
and UO_165 (O_165,N_4343,N_3598);
nand UO_166 (O_166,N_2607,N_4000);
nand UO_167 (O_167,N_4650,N_3557);
nor UO_168 (O_168,N_2843,N_2701);
nor UO_169 (O_169,N_4270,N_4740);
or UO_170 (O_170,N_3412,N_3789);
and UO_171 (O_171,N_3562,N_3762);
nor UO_172 (O_172,N_4272,N_3608);
nor UO_173 (O_173,N_3056,N_4497);
nand UO_174 (O_174,N_4984,N_4891);
or UO_175 (O_175,N_4030,N_4097);
or UO_176 (O_176,N_4805,N_3389);
nand UO_177 (O_177,N_4860,N_3394);
nand UO_178 (O_178,N_2517,N_2996);
or UO_179 (O_179,N_3759,N_4377);
or UO_180 (O_180,N_4229,N_3817);
nand UO_181 (O_181,N_2576,N_3350);
nand UO_182 (O_182,N_4719,N_2949);
nor UO_183 (O_183,N_3229,N_3253);
nor UO_184 (O_184,N_3365,N_4624);
or UO_185 (O_185,N_2523,N_2796);
or UO_186 (O_186,N_2892,N_3126);
and UO_187 (O_187,N_4458,N_4051);
and UO_188 (O_188,N_4886,N_3914);
nand UO_189 (O_189,N_3420,N_4908);
or UO_190 (O_190,N_2631,N_4525);
nand UO_191 (O_191,N_4102,N_3955);
nor UO_192 (O_192,N_4444,N_3115);
nor UO_193 (O_193,N_3867,N_3929);
or UO_194 (O_194,N_4641,N_4895);
nor UO_195 (O_195,N_4661,N_3526);
nand UO_196 (O_196,N_4223,N_2974);
nor UO_197 (O_197,N_4614,N_4297);
nor UO_198 (O_198,N_2503,N_3352);
nand UO_199 (O_199,N_3197,N_4822);
or UO_200 (O_200,N_3678,N_4578);
nor UO_201 (O_201,N_4352,N_3245);
or UO_202 (O_202,N_2587,N_4154);
or UO_203 (O_203,N_3458,N_2893);
or UO_204 (O_204,N_4643,N_4169);
and UO_205 (O_205,N_4685,N_2967);
nor UO_206 (O_206,N_3853,N_2856);
nand UO_207 (O_207,N_3021,N_2988);
and UO_208 (O_208,N_2765,N_3723);
or UO_209 (O_209,N_3770,N_3486);
and UO_210 (O_210,N_3385,N_4994);
nand UO_211 (O_211,N_4507,N_3190);
nor UO_212 (O_212,N_2933,N_4795);
and UO_213 (O_213,N_4474,N_4376);
or UO_214 (O_214,N_3815,N_4140);
nor UO_215 (O_215,N_4403,N_3579);
and UO_216 (O_216,N_2552,N_3227);
and UO_217 (O_217,N_4359,N_4840);
or UO_218 (O_218,N_3488,N_3766);
nor UO_219 (O_219,N_4098,N_2937);
nor UO_220 (O_220,N_3238,N_3918);
and UO_221 (O_221,N_3295,N_3895);
and UO_222 (O_222,N_2546,N_4031);
nor UO_223 (O_223,N_3518,N_3665);
or UO_224 (O_224,N_4626,N_2595);
nor UO_225 (O_225,N_3386,N_3116);
nor UO_226 (O_226,N_3603,N_4726);
or UO_227 (O_227,N_2656,N_3809);
nor UO_228 (O_228,N_3595,N_4192);
or UO_229 (O_229,N_4964,N_2732);
or UO_230 (O_230,N_3623,N_4854);
nor UO_231 (O_231,N_2502,N_3014);
and UO_232 (O_232,N_3757,N_4533);
nand UO_233 (O_233,N_4635,N_3607);
or UO_234 (O_234,N_4929,N_4656);
and UO_235 (O_235,N_4604,N_2686);
nand UO_236 (O_236,N_4718,N_3722);
nor UO_237 (O_237,N_4773,N_3299);
nand UO_238 (O_238,N_2529,N_4592);
nand UO_239 (O_239,N_4363,N_3071);
nor UO_240 (O_240,N_3647,N_4342);
nor UO_241 (O_241,N_4587,N_2671);
nor UO_242 (O_242,N_3121,N_3556);
or UO_243 (O_243,N_3141,N_3276);
or UO_244 (O_244,N_4734,N_3923);
or UO_245 (O_245,N_4421,N_3200);
or UO_246 (O_246,N_4161,N_3131);
and UO_247 (O_247,N_4232,N_4133);
nor UO_248 (O_248,N_3088,N_2872);
nand UO_249 (O_249,N_4595,N_4057);
and UO_250 (O_250,N_2833,N_4809);
nand UO_251 (O_251,N_2693,N_3335);
and UO_252 (O_252,N_3840,N_3887);
nor UO_253 (O_253,N_4061,N_4518);
and UO_254 (O_254,N_3004,N_4360);
nor UO_255 (O_255,N_2505,N_3122);
and UO_256 (O_256,N_2986,N_2942);
nor UO_257 (O_257,N_4743,N_4464);
nand UO_258 (O_258,N_4657,N_3907);
nor UO_259 (O_259,N_4907,N_4909);
nand UO_260 (O_260,N_3457,N_3627);
nand UO_261 (O_261,N_3784,N_2705);
or UO_262 (O_262,N_2881,N_4678);
and UO_263 (O_263,N_4437,N_4884);
and UO_264 (O_264,N_4457,N_3904);
and UO_265 (O_265,N_4503,N_4247);
or UO_266 (O_266,N_3913,N_3470);
and UO_267 (O_267,N_4749,N_4799);
or UO_268 (O_268,N_2613,N_4422);
or UO_269 (O_269,N_4336,N_2700);
and UO_270 (O_270,N_2524,N_3905);
nor UO_271 (O_271,N_3969,N_2969);
or UO_272 (O_272,N_3865,N_2736);
nor UO_273 (O_273,N_4820,N_4766);
nand UO_274 (O_274,N_4940,N_3592);
or UO_275 (O_275,N_3343,N_4793);
or UO_276 (O_276,N_2926,N_4253);
or UO_277 (O_277,N_2809,N_4644);
or UO_278 (O_278,N_2622,N_2977);
and UO_279 (O_279,N_3866,N_4495);
and UO_280 (O_280,N_3093,N_3469);
and UO_281 (O_281,N_4370,N_4168);
nand UO_282 (O_282,N_4472,N_2596);
or UO_283 (O_283,N_3328,N_3173);
and UO_284 (O_284,N_3622,N_3035);
and UO_285 (O_285,N_3686,N_3581);
xnor UO_286 (O_286,N_2916,N_4812);
nor UO_287 (O_287,N_3701,N_4200);
nand UO_288 (O_288,N_4796,N_3039);
and UO_289 (O_289,N_3917,N_4261);
nor UO_290 (O_290,N_4502,N_4531);
nand UO_291 (O_291,N_2635,N_3448);
or UO_292 (O_292,N_3125,N_3078);
and UO_293 (O_293,N_3106,N_3192);
and UO_294 (O_294,N_3862,N_4433);
nand UO_295 (O_295,N_3281,N_4572);
and UO_296 (O_296,N_3371,N_4972);
and UO_297 (O_297,N_3068,N_3208);
nor UO_298 (O_298,N_4085,N_2626);
nand UO_299 (O_299,N_4955,N_3467);
or UO_300 (O_300,N_4666,N_2902);
and UO_301 (O_301,N_4392,N_3582);
nor UO_302 (O_302,N_2520,N_3933);
and UO_303 (O_303,N_3986,N_4836);
nor UO_304 (O_304,N_4281,N_2855);
or UO_305 (O_305,N_4832,N_2757);
and UO_306 (O_306,N_3293,N_3888);
nor UO_307 (O_307,N_3042,N_3552);
and UO_308 (O_308,N_3076,N_4980);
nor UO_309 (O_309,N_4676,N_3696);
and UO_310 (O_310,N_3228,N_3252);
and UO_311 (O_311,N_4845,N_4228);
and UO_312 (O_312,N_2961,N_3445);
or UO_313 (O_313,N_3184,N_3694);
and UO_314 (O_314,N_2870,N_2971);
and UO_315 (O_315,N_3171,N_4121);
or UO_316 (O_316,N_4441,N_2649);
and UO_317 (O_317,N_4941,N_3878);
nor UO_318 (O_318,N_3829,N_4950);
or UO_319 (O_319,N_2606,N_3800);
nand UO_320 (O_320,N_4835,N_4548);
and UO_321 (O_321,N_2875,N_4557);
and UO_322 (O_322,N_3796,N_4957);
or UO_323 (O_323,N_3610,N_4962);
nand UO_324 (O_324,N_3396,N_4300);
nor UO_325 (O_325,N_3920,N_2909);
nor UO_326 (O_326,N_4983,N_3820);
and UO_327 (O_327,N_3451,N_4689);
nor UO_328 (O_328,N_4732,N_3492);
nor UO_329 (O_329,N_2648,N_3993);
or UO_330 (O_330,N_3861,N_3786);
and UO_331 (O_331,N_4917,N_4488);
nand UO_332 (O_332,N_2564,N_3123);
nand UO_333 (O_333,N_2575,N_3768);
nand UO_334 (O_334,N_4191,N_4398);
or UO_335 (O_335,N_3751,N_3256);
or UO_336 (O_336,N_4598,N_2910);
nand UO_337 (O_337,N_4373,N_4438);
nor UO_338 (O_338,N_3871,N_3688);
nor UO_339 (O_339,N_4280,N_4919);
or UO_340 (O_340,N_4966,N_4273);
nand UO_341 (O_341,N_3958,N_3615);
or UO_342 (O_342,N_4118,N_3397);
or UO_343 (O_343,N_3965,N_2669);
and UO_344 (O_344,N_4665,N_3988);
and UO_345 (O_345,N_3416,N_4347);
and UO_346 (O_346,N_4044,N_3163);
nand UO_347 (O_347,N_4707,N_3821);
and UO_348 (O_348,N_4863,N_3544);
and UO_349 (O_349,N_3733,N_4452);
or UO_350 (O_350,N_3361,N_2751);
or UO_351 (O_351,N_3712,N_4361);
or UO_352 (O_352,N_4857,N_3833);
nor UO_353 (O_353,N_4774,N_3236);
nor UO_354 (O_354,N_2710,N_3286);
nand UO_355 (O_355,N_3132,N_3440);
or UO_356 (O_356,N_4670,N_4368);
nor UO_357 (O_357,N_3611,N_4163);
nor UO_358 (O_358,N_4390,N_4634);
or UO_359 (O_359,N_3695,N_4658);
and UO_360 (O_360,N_2719,N_3736);
nand UO_361 (O_361,N_4362,N_4688);
nand UO_362 (O_362,N_2605,N_3110);
nand UO_363 (O_363,N_2623,N_3760);
nor UO_364 (O_364,N_3519,N_4107);
nand UO_365 (O_365,N_3325,N_3481);
nand UO_366 (O_366,N_3038,N_4901);
nor UO_367 (O_367,N_3261,N_4292);
or UO_368 (O_368,N_3839,N_3138);
or UO_369 (O_369,N_2540,N_3880);
or UO_370 (O_370,N_3710,N_2983);
and UO_371 (O_371,N_4428,N_2683);
and UO_372 (O_372,N_3339,N_4446);
and UO_373 (O_373,N_3219,N_3576);
nor UO_374 (O_374,N_4268,N_2506);
nor UO_375 (O_375,N_3763,N_4056);
nor UO_376 (O_376,N_3217,N_3001);
nor UO_377 (O_377,N_3146,N_3503);
or UO_378 (O_378,N_2621,N_2873);
and UO_379 (O_379,N_2941,N_4313);
and UO_380 (O_380,N_4974,N_3922);
nand UO_381 (O_381,N_4449,N_2679);
nand UO_382 (O_382,N_4623,N_2509);
nand UO_383 (O_383,N_3218,N_4173);
or UO_384 (O_384,N_2812,N_3538);
or UO_385 (O_385,N_4410,N_4910);
nand UO_386 (O_386,N_3787,N_4176);
or UO_387 (O_387,N_3978,N_4788);
or UO_388 (O_388,N_4956,N_4171);
nand UO_389 (O_389,N_4838,N_3506);
nor UO_390 (O_390,N_4408,N_3443);
or UO_391 (O_391,N_3439,N_3711);
and UO_392 (O_392,N_4482,N_3059);
nand UO_393 (O_393,N_2536,N_3714);
xor UO_394 (O_394,N_4002,N_3832);
and UO_395 (O_395,N_4108,N_3463);
and UO_396 (O_396,N_3555,N_3364);
and UO_397 (O_397,N_4755,N_4447);
and UO_398 (O_398,N_4923,N_3307);
or UO_399 (O_399,N_4344,N_4704);
and UO_400 (O_400,N_4631,N_3764);
and UO_401 (O_401,N_3034,N_4089);
and UO_402 (O_402,N_3625,N_3882);
and UO_403 (O_403,N_3604,N_2795);
and UO_404 (O_404,N_4852,N_4830);
nor UO_405 (O_405,N_2912,N_3240);
or UO_406 (O_406,N_3169,N_2832);
nand UO_407 (O_407,N_4862,N_4581);
nor UO_408 (O_408,N_3893,N_3578);
xnor UO_409 (O_409,N_2985,N_3850);
or UO_410 (O_410,N_3260,N_4646);
nand UO_411 (O_411,N_4546,N_2714);
nor UO_412 (O_412,N_2704,N_3437);
or UO_413 (O_413,N_3962,N_4692);
nor UO_414 (O_414,N_2709,N_2753);
nand UO_415 (O_415,N_3036,N_2657);
nor UO_416 (O_416,N_3589,N_3716);
and UO_417 (O_417,N_4167,N_3692);
or UO_418 (O_418,N_4079,N_4394);
nor UO_419 (O_419,N_4584,N_2752);
or UO_420 (O_420,N_3537,N_2797);
or UO_421 (O_421,N_3257,N_2756);
or UO_422 (O_422,N_3393,N_4266);
and UO_423 (O_423,N_4137,N_4791);
or UO_424 (O_424,N_3294,N_3112);
or UO_425 (O_425,N_3731,N_4003);
nand UO_426 (O_426,N_3926,N_4834);
nand UO_427 (O_427,N_3137,N_4638);
nand UO_428 (O_428,N_2610,N_2689);
or UO_429 (O_429,N_4750,N_3464);
and UO_430 (O_430,N_4600,N_3209);
nor UO_431 (O_431,N_2598,N_2811);
or UO_432 (O_432,N_3390,N_2849);
nor UO_433 (O_433,N_3903,N_4306);
or UO_434 (O_434,N_2945,N_4491);
nor UO_435 (O_435,N_3780,N_4404);
nor UO_436 (O_436,N_3483,N_4783);
nand UO_437 (O_437,N_4395,N_3527);
nand UO_438 (O_438,N_3387,N_3709);
and UO_439 (O_439,N_2525,N_3089);
and UO_440 (O_440,N_4203,N_2584);
nor UO_441 (O_441,N_4505,N_3810);
or UO_442 (O_442,N_3231,N_4020);
nor UO_443 (O_443,N_4054,N_3697);
nand UO_444 (O_444,N_2696,N_2609);
nor UO_445 (O_445,N_3264,N_2951);
or UO_446 (O_446,N_2992,N_3430);
or UO_447 (O_447,N_3855,N_4622);
or UO_448 (O_448,N_2954,N_2786);
nand UO_449 (O_449,N_2936,N_4681);
nand UO_450 (O_450,N_3013,N_3199);
and UO_451 (O_451,N_4138,N_4568);
and UO_452 (O_452,N_4660,N_2894);
or UO_453 (O_453,N_3310,N_4209);
nor UO_454 (O_454,N_4045,N_2660);
nand UO_455 (O_455,N_4754,N_4011);
or UO_456 (O_456,N_4416,N_3105);
and UO_457 (O_457,N_4028,N_4890);
nand UO_458 (O_458,N_3554,N_2848);
nor UO_459 (O_459,N_3835,N_4684);
nand UO_460 (O_460,N_3859,N_3111);
and UO_461 (O_461,N_4014,N_3849);
or UO_462 (O_462,N_4577,N_3330);
or UO_463 (O_463,N_2903,N_4742);
and UO_464 (O_464,N_3575,N_3737);
or UO_465 (O_465,N_3183,N_4668);
or UO_466 (O_466,N_4477,N_3741);
nand UO_467 (O_467,N_2801,N_3426);
and UO_468 (O_468,N_4702,N_2766);
or UO_469 (O_469,N_3207,N_4594);
nor UO_470 (O_470,N_4846,N_3643);
or UO_471 (O_471,N_2998,N_3202);
nand UO_472 (O_472,N_3438,N_4786);
nand UO_473 (O_473,N_2760,N_4304);
and UO_474 (O_474,N_4708,N_3521);
or UO_475 (O_475,N_4498,N_2680);
or UO_476 (O_476,N_3875,N_3915);
nor UO_477 (O_477,N_4858,N_3290);
or UO_478 (O_478,N_4520,N_4339);
or UO_479 (O_479,N_3341,N_2925);
and UO_480 (O_480,N_4224,N_3378);
and UO_481 (O_481,N_2543,N_4934);
nor UO_482 (O_482,N_2774,N_3894);
nand UO_483 (O_483,N_4985,N_4439);
or UO_484 (O_484,N_4083,N_3289);
nor UO_485 (O_485,N_4931,N_2512);
and UO_486 (O_486,N_3572,N_3377);
nor UO_487 (O_487,N_3327,N_4188);
nand UO_488 (O_488,N_3454,N_3108);
or UO_489 (O_489,N_4948,N_2664);
nand UO_490 (O_490,N_3363,N_4987);
and UO_491 (O_491,N_3471,N_2707);
or UO_492 (O_492,N_2668,N_2617);
xor UO_493 (O_493,N_3632,N_4165);
or UO_494 (O_494,N_2835,N_4970);
nor UO_495 (O_495,N_4182,N_3657);
and UO_496 (O_496,N_3851,N_2733);
nor UO_497 (O_497,N_3948,N_3434);
nand UO_498 (O_498,N_4072,N_2745);
nand UO_499 (O_499,N_3478,N_3594);
nand UO_500 (O_500,N_3682,N_3874);
or UO_501 (O_501,N_3362,N_3062);
and UO_502 (O_502,N_2802,N_3101);
or UO_503 (O_503,N_4236,N_3531);
xnor UO_504 (O_504,N_4258,N_4715);
and UO_505 (O_505,N_3724,N_3886);
and UO_506 (O_506,N_3542,N_3588);
and UO_507 (O_507,N_2860,N_3498);
nand UO_508 (O_508,N_4882,N_2627);
nor UO_509 (O_509,N_2964,N_4541);
and UO_510 (O_510,N_3569,N_4747);
nor UO_511 (O_511,N_3302,N_4769);
or UO_512 (O_512,N_3791,N_4811);
or UO_513 (O_513,N_3852,N_4379);
and UO_514 (O_514,N_3411,N_4873);
nand UO_515 (O_515,N_4283,N_4331);
and UO_516 (O_516,N_3549,N_4036);
nor UO_517 (O_517,N_2782,N_3727);
or UO_518 (O_518,N_4659,N_3382);
or UO_519 (O_519,N_2615,N_4785);
nand UO_520 (O_520,N_3214,N_3370);
and UO_521 (O_521,N_4990,N_2559);
or UO_522 (O_522,N_2874,N_4293);
or UO_523 (O_523,N_4620,N_3474);
nand UO_524 (O_524,N_3472,N_2948);
and UO_525 (O_525,N_4149,N_2859);
and UO_526 (O_526,N_4562,N_4013);
or UO_527 (O_527,N_2871,N_2535);
nor UO_528 (O_528,N_4301,N_2518);
nand UO_529 (O_529,N_4517,N_4981);
xnor UO_530 (O_530,N_3819,N_3097);
or UO_531 (O_531,N_3609,N_4878);
nor UO_532 (O_532,N_3584,N_3511);
and UO_533 (O_533,N_2819,N_3313);
and UO_534 (O_534,N_4197,N_4371);
or UO_535 (O_535,N_3550,N_3103);
nor UO_536 (O_536,N_2861,N_4951);
and UO_537 (O_537,N_3144,N_3017);
nor UO_538 (O_538,N_4653,N_4431);
and UO_539 (O_539,N_2830,N_4492);
and UO_540 (O_540,N_2624,N_3828);
or UO_541 (O_541,N_3309,N_4989);
and UO_542 (O_542,N_3422,N_3306);
nor UO_543 (O_543,N_3388,N_4196);
nor UO_544 (O_544,N_3381,N_2572);
or UO_545 (O_545,N_4162,N_3127);
or UO_546 (O_546,N_4175,N_3728);
and UO_547 (O_547,N_2741,N_3939);
nor UO_548 (O_548,N_3530,N_4160);
or UO_549 (O_549,N_4357,N_3303);
nand UO_550 (O_550,N_3423,N_4784);
nand UO_551 (O_551,N_3753,N_3180);
or UO_552 (O_552,N_3899,N_4101);
nand UO_553 (O_553,N_4285,N_3646);
nor UO_554 (O_554,N_3825,N_4506);
and UO_555 (O_555,N_4109,N_3098);
or UO_556 (O_556,N_3193,N_2589);
or UO_557 (O_557,N_3010,N_4928);
nand UO_558 (O_558,N_3096,N_4338);
or UO_559 (O_559,N_2845,N_2775);
and UO_560 (O_560,N_3916,N_3585);
nor UO_561 (O_561,N_2580,N_4949);
and UO_562 (O_562,N_4348,N_2824);
or UO_563 (O_563,N_2722,N_2573);
nand UO_564 (O_564,N_4246,N_2717);
or UO_565 (O_565,N_2891,N_4730);
nor UO_566 (O_566,N_3672,N_4311);
nand UO_567 (O_567,N_3466,N_3482);
or UO_568 (O_568,N_4500,N_4146);
nor UO_569 (O_569,N_3981,N_3095);
nand UO_570 (O_570,N_3073,N_3271);
or UO_571 (O_571,N_4736,N_4690);
nor UO_572 (O_572,N_2738,N_3599);
or UO_573 (O_573,N_3799,N_3075);
nor UO_574 (O_574,N_2747,N_4419);
or UO_575 (O_575,N_4839,N_3957);
and UO_576 (O_576,N_2720,N_4735);
and UO_577 (O_577,N_4310,N_2897);
and UO_578 (O_578,N_4124,N_3060);
and UO_579 (O_579,N_3230,N_4609);
or UO_580 (O_580,N_4800,N_2500);
or UO_581 (O_581,N_3250,N_4103);
and UO_582 (O_582,N_3885,N_4837);
or UO_583 (O_583,N_2876,N_3951);
nor UO_584 (O_584,N_4712,N_4642);
nand UO_585 (O_585,N_3931,N_4393);
nand UO_586 (O_586,N_4815,N_4282);
or UO_587 (O_587,N_2798,N_4543);
and UO_588 (O_588,N_4537,N_4024);
nor UO_589 (O_589,N_4611,N_4998);
or UO_590 (O_590,N_2952,N_4307);
or UO_591 (O_591,N_4515,N_4120);
or UO_592 (O_592,N_2938,N_2585);
or UO_593 (O_593,N_3637,N_4637);
or UO_594 (O_594,N_4042,N_3586);
and UO_595 (O_595,N_3563,N_4211);
nor UO_596 (O_596,N_2698,N_3398);
xor UO_597 (O_597,N_4455,N_3520);
nor UO_598 (O_598,N_4467,N_4350);
nor UO_599 (O_599,N_4879,N_4991);
or UO_600 (O_600,N_4526,N_3414);
or UO_601 (O_601,N_4346,N_2981);
or UO_602 (O_602,N_3788,N_4322);
and UO_603 (O_603,N_3375,N_4947);
nor UO_604 (O_604,N_3124,N_3848);
and UO_605 (O_605,N_4967,N_3114);
or UO_606 (O_606,N_3232,N_3943);
and UO_607 (O_607,N_4068,N_4691);
nor UO_608 (O_608,N_4672,N_2703);
nand UO_609 (O_609,N_4771,N_4727);
or UO_610 (O_610,N_4436,N_4271);
nor UO_611 (O_611,N_4023,N_3717);
nor UO_612 (O_612,N_4230,N_2651);
or UO_613 (O_613,N_4216,N_3983);
or UO_614 (O_614,N_4744,N_3813);
and UO_615 (O_615,N_3558,N_3629);
or UO_616 (O_616,N_3318,N_3086);
nand UO_617 (O_617,N_4067,N_4625);
nand UO_618 (O_618,N_2633,N_2674);
and UO_619 (O_619,N_3987,N_3011);
or UO_620 (O_620,N_4575,N_2570);
or UO_621 (O_621,N_4818,N_2863);
nor UO_622 (O_622,N_4521,N_4831);
xor UO_623 (O_623,N_2917,N_2866);
or UO_624 (O_624,N_4295,N_3802);
nor UO_625 (O_625,N_2650,N_4971);
and UO_626 (O_626,N_2818,N_3765);
nor UO_627 (O_627,N_2900,N_4267);
nor UO_628 (O_628,N_4070,N_4460);
nor UO_629 (O_629,N_3940,N_3945);
nand UO_630 (O_630,N_3704,N_3175);
nor UO_631 (O_631,N_3906,N_4468);
and UO_632 (O_632,N_3778,N_2685);
nand UO_633 (O_633,N_3648,N_3213);
nor UO_634 (O_634,N_3408,N_4673);
or UO_635 (O_635,N_4086,N_3241);
and UO_636 (O_636,N_3359,N_4010);
or UO_637 (O_637,N_4412,N_2806);
nand UO_638 (O_638,N_4553,N_3405);
nand UO_639 (O_639,N_3315,N_3188);
or UO_640 (O_640,N_3120,N_4573);
nand UO_641 (O_641,N_4896,N_3742);
and UO_642 (O_642,N_4093,N_2675);
and UO_643 (O_643,N_3312,N_4570);
or UO_644 (O_644,N_3816,N_2630);
nor UO_645 (O_645,N_3729,N_3176);
or UO_646 (O_646,N_4613,N_4599);
nor UO_647 (O_647,N_3170,N_3461);
nor UO_648 (O_648,N_4127,N_4853);
and UO_649 (O_649,N_4142,N_3998);
or UO_650 (O_650,N_4877,N_3660);
nor UO_651 (O_651,N_4321,N_4046);
and UO_652 (O_652,N_3283,N_3775);
nand UO_653 (O_653,N_2655,N_4952);
and UO_654 (O_654,N_4423,N_4445);
nand UO_655 (O_655,N_4781,N_3805);
and UO_656 (O_656,N_3743,N_4706);
or UO_657 (O_657,N_4603,N_3811);
nand UO_658 (O_658,N_4680,N_4481);
and UO_659 (O_659,N_4679,N_3496);
nor UO_660 (O_660,N_3220,N_3502);
nor UO_661 (O_661,N_4899,N_4029);
nand UO_662 (O_662,N_4238,N_4693);
or UO_663 (O_663,N_2519,N_4892);
and UO_664 (O_664,N_3432,N_3024);
nor UO_665 (O_665,N_3165,N_3019);
nor UO_666 (O_666,N_4859,N_3532);
nand UO_667 (O_667,N_3152,N_3837);
and UO_668 (O_668,N_4340,N_4235);
nand UO_669 (O_669,N_2896,N_2746);
nor UO_670 (O_670,N_2851,N_3838);
or UO_671 (O_671,N_4221,N_4319);
and UO_672 (O_672,N_4999,N_2618);
nor UO_673 (O_673,N_4037,N_2513);
nand UO_674 (O_674,N_3781,N_4147);
and UO_675 (O_675,N_3406,N_2730);
and UO_676 (O_676,N_3989,N_2914);
or UO_677 (O_677,N_3326,N_4547);
or UO_678 (O_678,N_2787,N_2943);
nand UO_679 (O_679,N_4254,N_2511);
nor UO_680 (O_680,N_3357,N_4524);
nor UO_681 (O_681,N_3528,N_3201);
nor UO_682 (O_682,N_3522,N_4341);
nand UO_683 (O_683,N_2913,N_2644);
nor UO_684 (O_684,N_4152,N_2750);
nand UO_685 (O_685,N_4265,N_2854);
nand UO_686 (O_686,N_2694,N_3869);
nor UO_687 (O_687,N_4082,N_2568);
nor UO_688 (O_688,N_2968,N_3677);
nand UO_689 (O_689,N_3043,N_2604);
or UO_690 (O_690,N_3311,N_4897);
nor UO_691 (O_691,N_4946,N_4126);
and UO_692 (O_692,N_2743,N_3040);
and UO_693 (O_693,N_3638,N_4387);
nor UO_694 (O_694,N_3898,N_3597);
xor UO_695 (O_695,N_3854,N_3407);
nand UO_696 (O_696,N_3910,N_4903);
nor UO_697 (O_697,N_2640,N_4589);
nor UO_698 (O_698,N_4081,N_2665);
or UO_699 (O_699,N_3018,N_4001);
nand UO_700 (O_700,N_4119,N_3794);
and UO_701 (O_701,N_3651,N_3032);
and UO_702 (O_702,N_3718,N_4756);
or UO_703 (O_703,N_3591,N_3164);
or UO_704 (O_704,N_3058,N_4427);
or UO_705 (O_705,N_4504,N_4924);
nor UO_706 (O_706,N_3930,N_4080);
and UO_707 (O_707,N_4380,N_3720);
nand UO_708 (O_708,N_2603,N_4397);
nor UO_709 (O_709,N_3964,N_4456);
nand UO_710 (O_710,N_3807,N_3719);
and UO_711 (O_711,N_2562,N_3912);
or UO_712 (O_712,N_2583,N_4725);
and UO_713 (O_713,N_3735,N_2737);
nand UO_714 (O_714,N_4069,N_4768);
nor UO_715 (O_715,N_2991,N_2672);
or UO_716 (O_716,N_4470,N_2577);
xnor UO_717 (O_717,N_2789,N_2728);
and UO_718 (O_718,N_3616,N_2636);
or UO_719 (O_719,N_2773,N_4202);
nor UO_720 (O_720,N_2563,N_3064);
and UO_721 (O_721,N_2541,N_3970);
nor UO_722 (O_722,N_4549,N_3158);
and UO_723 (O_723,N_3602,N_3937);
nor UO_724 (O_724,N_2805,N_3536);
and UO_725 (O_725,N_3634,N_4544);
and UO_726 (O_726,N_4904,N_4780);
nor UO_727 (O_727,N_2673,N_3273);
or UO_728 (O_728,N_3997,N_4979);
nand UO_729 (O_729,N_2946,N_2740);
nand UO_730 (O_730,N_4454,N_2944);
or UO_731 (O_731,N_4682,N_3222);
and UO_732 (O_732,N_4797,N_4239);
nand UO_733 (O_733,N_3346,N_3278);
and UO_734 (O_734,N_4277,N_3836);
or UO_735 (O_735,N_2637,N_2724);
or UO_736 (O_736,N_3130,N_3546);
or UO_737 (O_737,N_3553,N_2997);
nand UO_738 (O_738,N_4861,N_3961);
and UO_739 (O_739,N_3379,N_4385);
or UO_740 (O_740,N_4286,N_4629);
or UO_741 (O_741,N_2639,N_4545);
or UO_742 (O_742,N_4728,N_4565);
or UO_743 (O_743,N_4205,N_4494);
nor UO_744 (O_744,N_4207,N_3782);
or UO_745 (O_745,N_4552,N_4760);
nand UO_746 (O_746,N_4364,N_4567);
nand UO_747 (O_747,N_4961,N_4187);
or UO_748 (O_748,N_4511,N_3673);
nand UO_749 (O_749,N_2839,N_3155);
or UO_750 (O_750,N_3734,N_3857);
nor UO_751 (O_751,N_2661,N_4034);
or UO_752 (O_752,N_4337,N_4329);
nor UO_753 (O_753,N_4204,N_4710);
nor UO_754 (O_754,N_4490,N_4737);
nand UO_755 (O_755,N_3889,N_4274);
or UO_756 (O_756,N_2825,N_4305);
nand UO_757 (O_757,N_3732,N_4378);
or UO_758 (O_758,N_2553,N_4264);
nor UO_759 (O_759,N_3410,N_4806);
and UO_760 (O_760,N_3877,N_2890);
nor UO_761 (O_761,N_4559,N_3831);
or UO_762 (O_762,N_4913,N_4032);
nand UO_763 (O_763,N_3424,N_4415);
or UO_764 (O_764,N_4426,N_4406);
and UO_765 (O_765,N_3404,N_4212);
and UO_766 (O_766,N_3991,N_4210);
nand UO_767 (O_767,N_2599,N_4153);
or UO_768 (O_768,N_2666,N_3666);
nor UO_769 (O_769,N_4906,N_3685);
and UO_770 (O_770,N_4748,N_4782);
or UO_771 (O_771,N_2784,N_3317);
and UO_772 (O_772,N_3403,N_4864);
and UO_773 (O_773,N_4674,N_3834);
nand UO_774 (O_774,N_2888,N_2869);
and UO_775 (O_775,N_3104,N_3747);
and UO_776 (O_776,N_4787,N_3090);
nor UO_777 (O_777,N_4926,N_3324);
nand UO_778 (O_778,N_3342,N_2886);
and UO_779 (O_779,N_2813,N_4485);
nand UO_780 (O_780,N_2921,N_3195);
or UO_781 (O_781,N_3600,N_4463);
nor UO_782 (O_782,N_3639,N_4213);
and UO_783 (O_783,N_2723,N_3644);
nand UO_784 (O_784,N_2984,N_3700);
nand UO_785 (O_785,N_3347,N_2516);
and UO_786 (O_786,N_3074,N_3476);
and UO_787 (O_787,N_3005,N_3157);
or UO_788 (O_788,N_3547,N_4640);
and UO_789 (O_789,N_3996,N_2901);
or UO_790 (O_790,N_4078,N_2885);
or UO_791 (O_791,N_4842,N_2749);
nand UO_792 (O_792,N_2850,N_3272);
or UO_793 (O_793,N_4738,N_3590);
nor UO_794 (O_794,N_4538,N_4746);
or UO_795 (O_795,N_2558,N_3142);
and UO_796 (O_796,N_4775,N_3963);
nand UO_797 (O_797,N_4039,N_3402);
and UO_798 (O_798,N_3181,N_4237);
nor UO_799 (O_799,N_2600,N_4417);
or UO_800 (O_800,N_3935,N_4954);
nor UO_801 (O_801,N_3676,N_4939);
and UO_802 (O_802,N_4181,N_4296);
or UO_803 (O_803,N_4302,N_3640);
nor UO_804 (O_804,N_4569,N_3300);
or UO_805 (O_805,N_4473,N_4619);
nand UO_806 (O_806,N_3884,N_3650);
and UO_807 (O_807,N_2531,N_2834);
and UO_808 (O_808,N_3826,N_4986);
nand UO_809 (O_809,N_4466,N_4915);
nor UO_810 (O_810,N_3030,N_4060);
and UO_811 (O_811,N_3772,N_2612);
or UO_812 (O_812,N_2790,N_3083);
or UO_813 (O_813,N_4810,N_4328);
or UO_814 (O_814,N_4701,N_4016);
and UO_815 (O_815,N_3216,N_3016);
nand UO_816 (O_816,N_4969,N_4807);
and UO_817 (O_817,N_3559,N_4849);
nand UO_818 (O_818,N_4530,N_4475);
nand UO_819 (O_819,N_3136,N_3827);
nand UO_820 (O_820,N_4294,N_2729);
and UO_821 (O_821,N_2692,N_4761);
and UO_822 (O_822,N_3094,N_3975);
nor UO_823 (O_823,N_4529,N_4131);
nand UO_824 (O_824,N_4402,N_4514);
nor UO_825 (O_825,N_4435,N_3129);
nand UO_826 (O_826,N_2928,N_3689);
and UO_827 (O_827,N_2591,N_2858);
or UO_828 (O_828,N_2690,N_3577);
nor UO_829 (O_829,N_4150,N_3691);
nand UO_830 (O_830,N_3221,N_4116);
nand UO_831 (O_831,N_3196,N_2647);
nand UO_832 (O_832,N_2582,N_2887);
nor UO_833 (O_833,N_4731,N_4135);
or UO_834 (O_834,N_3336,N_3883);
or UO_835 (O_835,N_3061,N_4269);
nor UO_836 (O_836,N_4551,N_2905);
or UO_837 (O_837,N_3084,N_2879);
nor UO_838 (O_838,N_3031,N_4714);
nand UO_839 (O_839,N_4047,N_4593);
nand UO_840 (O_840,N_4992,N_3468);
or UO_841 (O_841,N_2687,N_4049);
or UO_842 (O_842,N_3818,N_4349);
xor UO_843 (O_843,N_3739,N_4601);
and UO_844 (O_844,N_3487,N_4716);
and UO_845 (O_845,N_2708,N_2846);
nor UO_846 (O_846,N_4561,N_4148);
xor UO_847 (O_847,N_3191,N_3092);
and UO_848 (O_848,N_3333,N_3740);
or UO_849 (O_849,N_2628,N_2642);
or UO_850 (O_850,N_3166,N_3954);
nor UO_851 (O_851,N_4434,N_3215);
and UO_852 (O_852,N_3803,N_3593);
nor UO_853 (O_853,N_4647,N_2831);
nor UO_854 (O_854,N_2638,N_2808);
and UO_855 (O_855,N_3462,N_4772);
nand UO_856 (O_856,N_3391,N_2758);
nor UO_857 (O_857,N_4717,N_2526);
nand UO_858 (O_858,N_3270,N_4356);
nor UO_859 (O_859,N_4554,N_4018);
or UO_860 (O_860,N_3161,N_4095);
or UO_861 (O_861,N_4172,N_3012);
and UO_862 (O_862,N_3707,N_4290);
nand UO_863 (O_863,N_4115,N_2567);
or UO_864 (O_864,N_3358,N_4440);
nor UO_865 (O_865,N_3446,N_3864);
nand UO_866 (O_866,N_2667,N_3630);
nor UO_867 (O_867,N_3267,N_4222);
nor UO_868 (O_868,N_3769,N_4179);
nor UO_869 (O_869,N_4699,N_4973);
and UO_870 (O_870,N_3117,N_4424);
or UO_871 (O_871,N_3548,N_4240);
or UO_872 (O_872,N_4790,N_4627);
nand UO_873 (O_873,N_3484,N_3606);
or UO_874 (O_874,N_3921,N_4499);
or UO_875 (O_875,N_3159,N_4789);
nor UO_876 (O_876,N_2670,N_4303);
nor UO_877 (O_877,N_2684,N_4317);
nor UO_878 (O_878,N_4021,N_3645);
and UO_879 (O_879,N_4865,N_2764);
nor UO_880 (O_880,N_4316,N_4912);
or UO_881 (O_881,N_4798,N_3746);
or UO_882 (O_882,N_4184,N_4881);
nand UO_883 (O_883,N_4677,N_4289);
or UO_884 (O_884,N_4418,N_3479);
nor UO_885 (O_885,N_3151,N_3626);
nor UO_886 (O_886,N_4618,N_3128);
and UO_887 (O_887,N_3571,N_4245);
and UO_888 (O_888,N_4703,N_3860);
and UO_889 (O_889,N_3655,N_3015);
or UO_890 (O_890,N_3844,N_3206);
nor UO_891 (O_891,N_2960,N_3713);
nand UO_892 (O_892,N_4501,N_4225);
nand UO_893 (O_893,N_2837,N_4617);
nand UO_894 (O_894,N_3758,N_4413);
and UO_895 (O_895,N_3049,N_4170);
nor UO_896 (O_896,N_4033,N_4945);
and UO_897 (O_897,N_4058,N_4851);
and UO_898 (O_898,N_4199,N_4358);
nand UO_899 (O_899,N_2976,N_3715);
nand UO_900 (O_900,N_4792,N_2594);
or UO_901 (O_901,N_4471,N_3028);
nor UO_902 (O_902,N_2718,N_3953);
or UO_903 (O_903,N_4123,N_4314);
nand UO_904 (O_904,N_4902,N_4571);
xor UO_905 (O_905,N_3282,N_3284);
or UO_906 (O_906,N_2972,N_3509);
and UO_907 (O_907,N_3198,N_3233);
nand UO_908 (O_908,N_3148,N_2557);
or UO_909 (O_909,N_3942,N_4916);
and UO_910 (O_910,N_3455,N_3683);
or UO_911 (O_911,N_2963,N_3881);
nand UO_912 (O_912,N_2691,N_4808);
and UO_913 (O_913,N_3992,N_3845);
and UO_914 (O_914,N_4334,N_4059);
and UO_915 (O_915,N_3465,N_3919);
or UO_916 (O_916,N_2940,N_4523);
nor UO_917 (O_917,N_3947,N_4757);
nand UO_918 (O_918,N_2793,N_4071);
or UO_919 (O_919,N_3203,N_3756);
nand UO_920 (O_920,N_3360,N_2522);
nand UO_921 (O_921,N_4764,N_3497);
nor UO_922 (O_922,N_4180,N_4279);
nor UO_923 (O_923,N_3435,N_4739);
nor UO_924 (O_924,N_4391,N_4132);
nand UO_925 (O_925,N_3255,N_2507);
and UO_926 (O_926,N_3456,N_3187);
nand UO_927 (O_927,N_3085,N_4012);
nor UO_928 (O_928,N_4145,N_3863);
or UO_929 (O_929,N_3441,N_4935);
nand UO_930 (O_930,N_2794,N_4106);
nand UO_931 (O_931,N_4741,N_3911);
nor UO_932 (O_932,N_3091,N_4649);
nand UO_933 (O_933,N_4606,N_3287);
nand UO_934 (O_934,N_2868,N_3072);
nor UO_935 (O_935,N_2574,N_4621);
nor UO_936 (O_936,N_4893,N_2821);
nor UO_937 (O_937,N_4696,N_4721);
and UO_938 (O_938,N_2884,N_4129);
nor UO_939 (O_939,N_2761,N_3587);
nand UO_940 (O_940,N_3946,N_2889);
nand UO_941 (O_941,N_2625,N_2920);
nor UO_942 (O_942,N_3972,N_4017);
and UO_943 (O_943,N_2571,N_4396);
or UO_944 (O_944,N_3633,N_4976);
and UO_945 (O_945,N_3178,N_2731);
nand UO_946 (O_946,N_3514,N_3490);
nor UO_947 (O_947,N_4164,N_3924);
or UO_948 (O_948,N_3368,N_3367);
nand UO_949 (O_949,N_2676,N_4256);
nand UO_950 (O_950,N_2538,N_4579);
or UO_951 (O_951,N_3767,N_2978);
nor UO_952 (O_952,N_3134,N_2560);
and UO_953 (O_953,N_3628,N_4654);
nor UO_954 (O_954,N_3226,N_4535);
and UO_955 (O_955,N_3960,N_3824);
and UO_956 (O_956,N_3376,N_3540);
nor UO_957 (O_957,N_4847,N_4958);
nor UO_958 (O_958,N_3269,N_4803);
or UO_959 (O_959,N_2785,N_4263);
xor UO_960 (O_960,N_2929,N_4027);
and UO_961 (O_961,N_3777,N_2841);
nor UO_962 (O_962,N_3372,N_2776);
or UO_963 (O_963,N_4231,N_4802);
or UO_964 (O_964,N_4420,N_4580);
or UO_965 (O_965,N_4513,N_4943);
nor UO_966 (O_966,N_4077,N_4590);
and UO_967 (O_967,N_3145,N_2586);
nand UO_968 (O_968,N_3771,N_3932);
nand UO_969 (O_969,N_3535,N_3243);
nor UO_970 (O_970,N_3868,N_3890);
nor UO_971 (O_971,N_3139,N_4843);
nand UO_972 (O_972,N_4560,N_3077);
and UO_973 (O_973,N_3400,N_4776);
nor UO_974 (O_974,N_3235,N_3204);
nor UO_975 (O_975,N_3706,N_4323);
nand UO_976 (O_976,N_2682,N_4874);
nor UO_977 (O_977,N_2957,N_3323);
nor UO_978 (O_978,N_3065,N_3902);
or UO_979 (O_979,N_4219,N_3107);
or UO_980 (O_980,N_3223,N_3703);
and UO_981 (O_981,N_3652,N_3524);
nor UO_982 (O_982,N_4963,N_3285);
nand UO_983 (O_983,N_3401,N_3297);
or UO_984 (O_984,N_3265,N_4519);
nand UO_985 (O_985,N_4597,N_3052);
nand UO_986 (O_986,N_4366,N_3081);
and UO_987 (O_987,N_2810,N_3744);
or UO_988 (O_988,N_4430,N_4193);
nor UO_989 (O_989,N_3795,N_3982);
nand UO_990 (O_990,N_2908,N_3690);
nand UO_991 (O_991,N_4476,N_4887);
and UO_992 (O_992,N_2803,N_2907);
or UO_993 (O_993,N_3515,N_3008);
and UO_994 (O_994,N_4667,N_3681);
nand UO_995 (O_995,N_4900,N_2721);
or UO_996 (O_996,N_3977,N_3057);
or UO_997 (O_997,N_4582,N_4489);
nor UO_998 (O_998,N_3210,N_3725);
nand UO_999 (O_999,N_3561,N_4066);
endmodule