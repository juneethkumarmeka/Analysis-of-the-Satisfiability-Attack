module basic_500_3000_500_40_levels_1xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_439,In_151);
nand U1 (N_1,In_449,In_164);
nor U2 (N_2,In_401,In_233);
and U3 (N_3,In_306,In_297);
and U4 (N_4,In_180,In_432);
or U5 (N_5,In_413,In_222);
nor U6 (N_6,In_85,In_274);
nand U7 (N_7,In_157,In_205);
xor U8 (N_8,In_88,In_351);
nand U9 (N_9,In_345,In_440);
nand U10 (N_10,In_145,In_321);
or U11 (N_11,In_67,In_25);
and U12 (N_12,In_236,In_290);
nor U13 (N_13,In_135,In_53);
nor U14 (N_14,In_223,In_166);
or U15 (N_15,In_357,In_386);
or U16 (N_16,In_475,In_227);
nor U17 (N_17,In_150,In_387);
nand U18 (N_18,In_473,In_385);
nand U19 (N_19,In_260,In_395);
and U20 (N_20,In_352,In_450);
or U21 (N_21,In_396,In_244);
nand U22 (N_22,In_226,In_253);
nand U23 (N_23,In_86,In_111);
nand U24 (N_24,In_87,In_231);
nand U25 (N_25,In_437,In_415);
nor U26 (N_26,In_377,In_52);
or U27 (N_27,In_178,In_492);
or U28 (N_28,In_115,In_113);
nand U29 (N_29,In_142,In_106);
or U30 (N_30,In_208,In_441);
and U31 (N_31,In_248,In_144);
or U32 (N_32,In_105,In_262);
nand U33 (N_33,In_390,In_268);
and U34 (N_34,In_183,In_276);
nor U35 (N_35,In_232,In_489);
nand U36 (N_36,In_393,In_389);
and U37 (N_37,In_430,In_35);
and U38 (N_38,In_370,In_22);
or U39 (N_39,In_350,In_266);
or U40 (N_40,In_414,In_9);
and U41 (N_41,In_96,In_71);
and U42 (N_42,In_221,In_195);
nor U43 (N_43,In_355,In_36);
nor U44 (N_44,In_376,In_343);
or U45 (N_45,In_323,In_484);
nor U46 (N_46,In_291,In_495);
nand U47 (N_47,In_123,In_243);
nor U48 (N_48,In_407,In_270);
and U49 (N_49,In_126,In_131);
and U50 (N_50,In_313,In_33);
nor U51 (N_51,In_211,In_26);
and U52 (N_52,In_456,In_471);
and U53 (N_53,In_277,In_44);
or U54 (N_54,In_436,In_7);
nand U55 (N_55,In_30,In_104);
nor U56 (N_56,In_463,In_138);
and U57 (N_57,In_392,In_37);
and U58 (N_58,In_140,In_168);
or U59 (N_59,In_356,In_40);
nor U60 (N_60,In_491,In_483);
nor U61 (N_61,In_314,In_146);
nor U62 (N_62,In_46,In_127);
or U63 (N_63,In_259,In_280);
nor U64 (N_64,In_174,In_444);
and U65 (N_65,In_47,In_372);
and U66 (N_66,In_404,In_339);
and U67 (N_67,In_250,In_296);
and U68 (N_68,In_263,In_496);
nor U69 (N_69,In_51,In_284);
nand U70 (N_70,In_136,In_77);
or U71 (N_71,In_204,In_6);
or U72 (N_72,In_100,In_358);
and U73 (N_73,In_487,In_162);
or U74 (N_74,In_82,In_379);
nor U75 (N_75,N_56,N_40);
or U76 (N_76,In_287,In_464);
and U77 (N_77,In_416,In_428);
nand U78 (N_78,In_39,In_13);
and U79 (N_79,In_2,In_89);
and U80 (N_80,In_188,In_344);
and U81 (N_81,In_448,N_18);
or U82 (N_82,In_23,N_13);
or U83 (N_83,In_275,In_315);
nand U84 (N_84,In_490,In_454);
or U85 (N_85,In_118,N_68);
nor U86 (N_86,In_196,In_161);
and U87 (N_87,In_45,In_330);
nand U88 (N_88,N_14,In_417);
nand U89 (N_89,In_83,In_125);
nor U90 (N_90,In_272,In_353);
and U91 (N_91,In_337,In_310);
nand U92 (N_92,In_293,In_74);
or U93 (N_93,In_63,In_307);
nor U94 (N_94,In_299,In_203);
nand U95 (N_95,In_173,In_468);
xnor U96 (N_96,In_59,N_74);
and U97 (N_97,In_331,In_108);
or U98 (N_98,In_418,In_48);
nor U99 (N_99,In_497,In_478);
or U100 (N_100,In_175,N_21);
and U101 (N_101,In_476,N_39);
or U102 (N_102,In_420,In_317);
or U103 (N_103,In_300,N_72);
or U104 (N_104,N_28,In_4);
nand U105 (N_105,In_32,In_431);
or U106 (N_106,In_129,In_285);
and U107 (N_107,In_158,In_57);
nand U108 (N_108,In_119,In_15);
or U109 (N_109,In_316,In_419);
and U110 (N_110,In_271,In_455);
and U111 (N_111,In_206,In_187);
and U112 (N_112,In_470,In_303);
and U113 (N_113,In_499,N_41);
or U114 (N_114,In_324,In_384);
or U115 (N_115,In_27,In_247);
nor U116 (N_116,N_3,N_37);
or U117 (N_117,In_446,N_7);
nand U118 (N_118,In_170,In_381);
nor U119 (N_119,In_38,In_281);
or U120 (N_120,In_18,In_156);
and U121 (N_121,In_265,In_269);
nand U122 (N_122,In_477,N_50);
nand U123 (N_123,In_116,In_19);
or U124 (N_124,In_159,In_76);
nand U125 (N_125,In_101,In_371);
nor U126 (N_126,In_264,N_47);
nor U127 (N_127,N_38,N_36);
nand U128 (N_128,In_363,In_466);
nor U129 (N_129,In_383,In_242);
nor U130 (N_130,N_6,In_176);
nor U131 (N_131,In_434,In_273);
or U132 (N_132,In_172,In_254);
or U133 (N_133,In_238,In_219);
or U134 (N_134,In_132,In_325);
nor U135 (N_135,N_67,In_133);
and U136 (N_136,In_241,N_55);
nand U137 (N_137,In_124,In_334);
nand U138 (N_138,N_12,In_469);
nand U139 (N_139,In_305,In_453);
and U140 (N_140,In_34,In_72);
or U141 (N_141,In_309,In_286);
nand U142 (N_142,In_429,N_69);
or U143 (N_143,N_29,In_0);
nor U144 (N_144,In_267,In_197);
nor U145 (N_145,In_10,In_95);
or U146 (N_146,In_257,In_41);
and U147 (N_147,In_400,In_410);
and U148 (N_148,In_301,In_362);
nor U149 (N_149,In_399,In_341);
or U150 (N_150,In_163,In_128);
and U151 (N_151,In_348,N_60);
and U152 (N_152,N_4,N_61);
or U153 (N_153,N_90,In_75);
nand U154 (N_154,In_474,N_116);
or U155 (N_155,N_22,In_279);
nor U156 (N_156,In_402,In_452);
nand U157 (N_157,In_361,In_467);
nor U158 (N_158,In_423,In_93);
nand U159 (N_159,In_346,In_92);
nor U160 (N_160,N_93,In_143);
nor U161 (N_161,In_320,In_1);
and U162 (N_162,In_107,In_216);
and U163 (N_163,N_141,N_143);
or U164 (N_164,In_189,In_424);
nor U165 (N_165,N_46,In_283);
nor U166 (N_166,In_294,In_486);
nor U167 (N_167,N_5,In_3);
or U168 (N_168,In_65,In_167);
or U169 (N_169,In_398,In_69);
and U170 (N_170,In_459,In_29);
nand U171 (N_171,In_120,N_51);
and U172 (N_172,N_17,In_426);
nor U173 (N_173,In_5,In_185);
nor U174 (N_174,In_458,N_107);
and U175 (N_175,N_88,In_84);
nor U176 (N_176,In_148,In_465);
nor U177 (N_177,In_342,In_165);
nor U178 (N_178,In_494,N_97);
nand U179 (N_179,N_99,N_106);
nor U180 (N_180,N_87,In_112);
and U181 (N_181,In_54,In_179);
or U182 (N_182,In_328,In_472);
nor U183 (N_183,In_215,In_192);
nand U184 (N_184,N_65,N_117);
nand U185 (N_185,In_388,In_295);
nor U186 (N_186,In_493,In_457);
nand U187 (N_187,In_182,N_98);
and U188 (N_188,N_19,In_49);
and U189 (N_189,In_190,N_66);
or U190 (N_190,In_354,In_66);
nand U191 (N_191,In_249,In_368);
nand U192 (N_192,In_68,In_256);
or U193 (N_193,In_397,In_319);
nand U194 (N_194,In_336,In_31);
and U195 (N_195,N_118,In_246);
nor U196 (N_196,In_90,N_146);
and U197 (N_197,In_198,In_322);
nand U198 (N_198,In_169,N_43);
nor U199 (N_199,In_378,In_224);
xor U200 (N_200,N_59,N_103);
nor U201 (N_201,N_123,In_482);
nor U202 (N_202,In_16,In_405);
nand U203 (N_203,In_391,In_435);
and U204 (N_204,In_60,N_125);
nand U205 (N_205,N_0,In_79);
nand U206 (N_206,In_199,In_422);
nand U207 (N_207,In_421,N_79);
nand U208 (N_208,N_23,N_53);
nor U209 (N_209,In_230,In_160);
and U210 (N_210,In_193,In_427);
nor U211 (N_211,N_139,N_110);
nor U212 (N_212,N_140,In_8);
or U213 (N_213,In_382,In_134);
nor U214 (N_214,In_326,In_251);
nand U215 (N_215,In_261,In_17);
nand U216 (N_216,In_394,In_234);
nand U217 (N_217,In_409,N_86);
nand U218 (N_218,N_2,In_80);
or U219 (N_219,N_112,In_12);
or U220 (N_220,N_114,N_145);
nand U221 (N_221,In_365,In_403);
nor U222 (N_222,N_75,In_201);
nor U223 (N_223,N_52,In_335);
or U224 (N_224,In_97,In_239);
nor U225 (N_225,In_329,In_327);
or U226 (N_226,N_149,N_191);
and U227 (N_227,N_119,In_282);
nor U228 (N_228,N_176,N_54);
nand U229 (N_229,In_91,In_218);
or U230 (N_230,In_220,In_109);
nor U231 (N_231,In_406,In_21);
xnor U232 (N_232,In_438,In_153);
or U233 (N_233,In_99,N_91);
or U234 (N_234,In_318,N_152);
or U235 (N_235,N_174,N_63);
nand U236 (N_236,N_206,N_26);
nand U237 (N_237,In_240,N_58);
nand U238 (N_238,N_132,N_122);
or U239 (N_239,N_218,N_64);
or U240 (N_240,In_147,N_126);
and U241 (N_241,N_27,In_214);
nand U242 (N_242,N_81,N_92);
nand U243 (N_243,N_135,N_150);
nor U244 (N_244,N_163,N_222);
nor U245 (N_245,N_154,In_202);
nor U246 (N_246,In_117,In_207);
or U247 (N_247,N_73,In_408);
and U248 (N_248,In_364,N_210);
nand U249 (N_249,In_451,N_197);
and U250 (N_250,In_155,In_50);
and U251 (N_251,N_160,N_16);
or U252 (N_252,In_245,N_32);
nor U253 (N_253,In_338,N_205);
nor U254 (N_254,N_190,In_411);
nor U255 (N_255,N_105,In_62);
nor U256 (N_256,In_373,N_201);
and U257 (N_257,N_131,In_121);
nor U258 (N_258,N_184,N_215);
nor U259 (N_259,In_433,N_34);
nand U260 (N_260,In_171,N_82);
or U261 (N_261,N_129,In_258);
nand U262 (N_262,N_221,N_95);
or U263 (N_263,In_255,In_380);
nor U264 (N_264,N_155,N_151);
and U265 (N_265,N_166,N_102);
nand U266 (N_266,N_194,In_213);
or U267 (N_267,N_44,In_209);
and U268 (N_268,In_14,N_20);
and U269 (N_269,N_181,N_80);
or U270 (N_270,In_304,In_122);
nor U271 (N_271,In_184,N_77);
or U272 (N_272,In_20,N_156);
nand U273 (N_273,In_181,N_128);
nand U274 (N_274,N_165,N_169);
or U275 (N_275,In_442,N_168);
and U276 (N_276,N_157,N_164);
or U277 (N_277,In_24,N_1);
and U278 (N_278,N_183,In_11);
or U279 (N_279,In_137,In_102);
nand U280 (N_280,In_375,In_278);
and U281 (N_281,N_49,N_178);
or U282 (N_282,N_175,N_203);
or U283 (N_283,In_498,In_55);
xnor U284 (N_284,N_188,In_312);
or U285 (N_285,In_292,In_235);
nand U286 (N_286,N_124,In_366);
or U287 (N_287,N_192,N_24);
nor U288 (N_288,N_83,N_216);
and U289 (N_289,In_61,N_223);
and U290 (N_290,N_120,N_148);
nand U291 (N_291,N_180,In_228);
nor U292 (N_292,In_481,N_108);
nor U293 (N_293,In_200,In_488);
nor U294 (N_294,N_159,N_130);
or U295 (N_295,N_198,N_8);
and U296 (N_296,In_229,In_289);
nand U297 (N_297,N_153,N_76);
or U298 (N_298,N_10,In_177);
nand U299 (N_299,In_154,In_347);
nor U300 (N_300,N_162,N_255);
nand U301 (N_301,N_45,N_187);
nand U302 (N_302,N_287,N_109);
nand U303 (N_303,N_199,N_281);
and U304 (N_304,N_241,N_271);
nor U305 (N_305,N_84,N_239);
and U306 (N_306,N_250,In_237);
and U307 (N_307,In_114,N_247);
nand U308 (N_308,N_213,In_462);
and U309 (N_309,N_185,N_78);
or U310 (N_310,In_58,In_217);
and U311 (N_311,N_189,In_43);
or U312 (N_312,In_212,N_202);
nor U313 (N_313,In_332,N_147);
nand U314 (N_314,N_170,N_70);
or U315 (N_315,N_240,N_173);
nand U316 (N_316,In_443,N_224);
and U317 (N_317,N_207,N_217);
and U318 (N_318,N_278,In_302);
nor U319 (N_319,N_121,N_269);
nor U320 (N_320,N_133,N_249);
and U321 (N_321,N_204,N_288);
nor U322 (N_322,In_64,In_98);
nor U323 (N_323,N_134,N_274);
nand U324 (N_324,In_460,N_186);
nor U325 (N_325,In_340,N_48);
nand U326 (N_326,N_292,N_182);
nor U327 (N_327,N_11,N_233);
nand U328 (N_328,N_144,N_261);
nand U329 (N_329,N_283,In_152);
nor U330 (N_330,N_293,In_252);
or U331 (N_331,N_137,N_280);
or U332 (N_332,In_78,N_227);
nand U333 (N_333,In_81,N_256);
and U334 (N_334,N_289,In_461);
nor U335 (N_335,N_248,N_297);
or U336 (N_336,N_276,N_104);
nand U337 (N_337,N_295,In_42);
xor U338 (N_338,N_277,N_196);
nor U339 (N_339,N_42,N_267);
and U340 (N_340,N_253,N_177);
and U341 (N_341,In_485,N_279);
or U342 (N_342,N_229,N_262);
and U343 (N_343,N_214,In_480);
and U344 (N_344,N_291,In_186);
or U345 (N_345,N_193,In_139);
nor U346 (N_346,N_282,N_228);
nand U347 (N_347,In_308,N_113);
nor U348 (N_348,N_158,N_136);
or U349 (N_349,In_73,N_209);
and U350 (N_350,N_258,N_290);
nand U351 (N_351,N_96,N_161);
and U352 (N_352,N_296,In_369);
nor U353 (N_353,In_445,In_28);
and U354 (N_354,N_264,N_15);
or U355 (N_355,N_252,N_237);
or U356 (N_356,N_167,N_171);
nand U357 (N_357,N_89,N_259);
or U358 (N_358,N_211,N_115);
and U359 (N_359,N_298,N_235);
xnor U360 (N_360,N_263,In_149);
nor U361 (N_361,N_208,N_294);
nand U362 (N_362,In_130,In_110);
nor U363 (N_363,N_138,In_288);
and U364 (N_364,N_268,N_142);
or U365 (N_365,N_238,N_257);
or U366 (N_366,In_94,N_200);
and U367 (N_367,N_179,N_299);
nand U368 (N_368,N_244,N_260);
nor U369 (N_369,N_275,N_31);
or U370 (N_370,N_94,N_226);
and U371 (N_371,N_272,In_298);
or U372 (N_372,N_285,N_25);
nand U373 (N_373,N_243,N_127);
and U374 (N_374,N_212,N_270);
or U375 (N_375,N_62,N_349);
nand U376 (N_376,N_225,In_191);
nor U377 (N_377,N_326,N_339);
and U378 (N_378,N_306,N_308);
and U379 (N_379,N_246,N_360);
nor U380 (N_380,N_367,N_230);
or U381 (N_381,N_323,N_302);
nand U382 (N_382,N_301,N_366);
or U383 (N_383,In_210,N_370);
or U384 (N_384,N_361,N_356);
nor U385 (N_385,N_374,N_330);
nor U386 (N_386,N_220,N_245);
nand U387 (N_387,N_321,N_172);
and U388 (N_388,N_337,N_327);
and U389 (N_389,N_111,N_85);
and U390 (N_390,N_341,N_319);
nand U391 (N_391,N_336,N_325);
and U392 (N_392,N_320,N_317);
nor U393 (N_393,N_331,N_333);
nor U394 (N_394,N_101,N_373);
and U395 (N_395,N_346,N_266);
or U396 (N_396,In_447,N_219);
nand U397 (N_397,In_374,N_303);
nor U398 (N_398,N_9,N_33);
nor U399 (N_399,In_103,In_359);
nand U400 (N_400,N_236,N_355);
nand U401 (N_401,N_353,N_310);
nand U402 (N_402,N_340,N_304);
and U403 (N_403,N_311,N_329);
nor U404 (N_404,N_313,N_307);
nand U405 (N_405,In_425,In_367);
and U406 (N_406,N_57,N_322);
nand U407 (N_407,N_338,N_251);
nor U408 (N_408,N_365,N_305);
or U409 (N_409,In_412,N_350);
nand U410 (N_410,N_344,N_359);
nor U411 (N_411,N_232,N_30);
and U412 (N_412,N_35,N_100);
or U413 (N_413,N_286,N_347);
nand U414 (N_414,In_56,N_354);
or U415 (N_415,N_372,In_311);
and U416 (N_416,N_195,In_70);
nor U417 (N_417,N_351,N_368);
or U418 (N_418,N_265,N_318);
or U419 (N_419,N_358,In_194);
nand U420 (N_420,N_316,In_225);
nor U421 (N_421,N_312,N_369);
nand U422 (N_422,N_284,N_71);
or U423 (N_423,N_363,N_231);
nor U424 (N_424,N_234,N_357);
nor U425 (N_425,N_300,N_314);
or U426 (N_426,N_315,N_335);
or U427 (N_427,In_479,In_349);
and U428 (N_428,N_364,N_342);
nand U429 (N_429,N_254,N_328);
and U430 (N_430,N_309,In_141);
nand U431 (N_431,N_343,In_333);
and U432 (N_432,N_242,N_362);
and U433 (N_433,N_352,N_273);
and U434 (N_434,N_348,N_324);
nand U435 (N_435,N_334,N_332);
or U436 (N_436,N_345,In_360);
nor U437 (N_437,N_371,N_341);
or U438 (N_438,N_337,N_302);
nor U439 (N_439,N_362,N_266);
or U440 (N_440,N_317,N_332);
and U441 (N_441,N_306,N_346);
nand U442 (N_442,N_352,N_348);
nor U443 (N_443,N_284,N_326);
and U444 (N_444,N_302,In_349);
nor U445 (N_445,N_62,N_286);
and U446 (N_446,N_232,In_359);
or U447 (N_447,N_302,N_349);
or U448 (N_448,In_374,N_311);
nor U449 (N_449,N_195,In_103);
or U450 (N_450,N_441,N_407);
or U451 (N_451,N_401,N_411);
nand U452 (N_452,N_386,N_435);
nor U453 (N_453,N_396,N_379);
and U454 (N_454,N_445,N_437);
and U455 (N_455,N_378,N_399);
nor U456 (N_456,N_429,N_420);
or U457 (N_457,N_398,N_391);
and U458 (N_458,N_449,N_400);
or U459 (N_459,N_440,N_380);
nand U460 (N_460,N_418,N_434);
and U461 (N_461,N_447,N_405);
nor U462 (N_462,N_444,N_431);
and U463 (N_463,N_385,N_413);
and U464 (N_464,N_409,N_416);
nor U465 (N_465,N_443,N_448);
or U466 (N_466,N_439,N_415);
and U467 (N_467,N_424,N_423);
nor U468 (N_468,N_402,N_408);
or U469 (N_469,N_376,N_438);
nor U470 (N_470,N_442,N_406);
nor U471 (N_471,N_375,N_392);
or U472 (N_472,N_446,N_436);
nand U473 (N_473,N_395,N_382);
nor U474 (N_474,N_414,N_433);
and U475 (N_475,N_422,N_425);
and U476 (N_476,N_427,N_381);
nor U477 (N_477,N_388,N_389);
or U478 (N_478,N_419,N_387);
and U479 (N_479,N_432,N_383);
and U480 (N_480,N_430,N_394);
and U481 (N_481,N_384,N_397);
and U482 (N_482,N_410,N_390);
nor U483 (N_483,N_421,N_393);
or U484 (N_484,N_417,N_412);
or U485 (N_485,N_426,N_377);
or U486 (N_486,N_404,N_403);
nor U487 (N_487,N_428,N_389);
or U488 (N_488,N_387,N_408);
and U489 (N_489,N_419,N_392);
or U490 (N_490,N_416,N_431);
nor U491 (N_491,N_428,N_397);
nor U492 (N_492,N_447,N_418);
nor U493 (N_493,N_431,N_415);
nor U494 (N_494,N_376,N_429);
nand U495 (N_495,N_414,N_392);
and U496 (N_496,N_415,N_384);
and U497 (N_497,N_422,N_408);
nand U498 (N_498,N_404,N_424);
or U499 (N_499,N_439,N_411);
or U500 (N_500,N_433,N_378);
nor U501 (N_501,N_390,N_378);
and U502 (N_502,N_431,N_418);
nor U503 (N_503,N_431,N_421);
nor U504 (N_504,N_395,N_397);
nand U505 (N_505,N_449,N_397);
or U506 (N_506,N_385,N_399);
nor U507 (N_507,N_420,N_389);
or U508 (N_508,N_394,N_393);
or U509 (N_509,N_376,N_414);
and U510 (N_510,N_440,N_384);
or U511 (N_511,N_423,N_383);
nor U512 (N_512,N_407,N_429);
nand U513 (N_513,N_386,N_388);
and U514 (N_514,N_426,N_390);
or U515 (N_515,N_425,N_442);
and U516 (N_516,N_399,N_411);
and U517 (N_517,N_431,N_427);
nand U518 (N_518,N_411,N_398);
nand U519 (N_519,N_408,N_390);
nor U520 (N_520,N_418,N_395);
nor U521 (N_521,N_382,N_437);
and U522 (N_522,N_382,N_402);
and U523 (N_523,N_386,N_403);
and U524 (N_524,N_410,N_422);
and U525 (N_525,N_511,N_502);
nand U526 (N_526,N_454,N_519);
and U527 (N_527,N_453,N_452);
or U528 (N_528,N_503,N_516);
or U529 (N_529,N_471,N_523);
nand U530 (N_530,N_476,N_500);
and U531 (N_531,N_496,N_462);
and U532 (N_532,N_463,N_477);
or U533 (N_533,N_497,N_470);
nor U534 (N_534,N_484,N_509);
nand U535 (N_535,N_507,N_451);
or U536 (N_536,N_512,N_473);
nand U537 (N_537,N_455,N_521);
or U538 (N_538,N_475,N_514);
or U539 (N_539,N_506,N_460);
nor U540 (N_540,N_450,N_491);
and U541 (N_541,N_459,N_482);
and U542 (N_542,N_478,N_488);
and U543 (N_543,N_481,N_495);
nor U544 (N_544,N_504,N_472);
nor U545 (N_545,N_524,N_490);
or U546 (N_546,N_483,N_498);
nor U547 (N_547,N_466,N_510);
or U548 (N_548,N_505,N_517);
nor U549 (N_549,N_465,N_487);
nand U550 (N_550,N_515,N_468);
nor U551 (N_551,N_492,N_486);
nand U552 (N_552,N_461,N_501);
or U553 (N_553,N_493,N_467);
or U554 (N_554,N_474,N_480);
or U555 (N_555,N_513,N_518);
or U556 (N_556,N_520,N_457);
or U557 (N_557,N_479,N_456);
and U558 (N_558,N_489,N_494);
nand U559 (N_559,N_458,N_485);
nor U560 (N_560,N_464,N_499);
nor U561 (N_561,N_522,N_469);
nand U562 (N_562,N_508,N_515);
nor U563 (N_563,N_483,N_512);
nand U564 (N_564,N_491,N_462);
nand U565 (N_565,N_514,N_488);
and U566 (N_566,N_484,N_476);
nor U567 (N_567,N_511,N_460);
nand U568 (N_568,N_518,N_485);
and U569 (N_569,N_492,N_465);
nor U570 (N_570,N_493,N_453);
or U571 (N_571,N_493,N_509);
or U572 (N_572,N_466,N_518);
nand U573 (N_573,N_508,N_513);
or U574 (N_574,N_515,N_489);
nor U575 (N_575,N_509,N_474);
or U576 (N_576,N_512,N_474);
or U577 (N_577,N_460,N_478);
nand U578 (N_578,N_469,N_484);
or U579 (N_579,N_518,N_493);
nand U580 (N_580,N_499,N_480);
or U581 (N_581,N_450,N_484);
or U582 (N_582,N_465,N_476);
or U583 (N_583,N_466,N_509);
and U584 (N_584,N_484,N_473);
nor U585 (N_585,N_516,N_486);
or U586 (N_586,N_464,N_459);
nand U587 (N_587,N_517,N_477);
and U588 (N_588,N_463,N_516);
or U589 (N_589,N_500,N_488);
nor U590 (N_590,N_496,N_495);
and U591 (N_591,N_502,N_457);
nor U592 (N_592,N_524,N_471);
nand U593 (N_593,N_477,N_498);
nand U594 (N_594,N_520,N_459);
nor U595 (N_595,N_492,N_456);
nor U596 (N_596,N_507,N_496);
and U597 (N_597,N_480,N_450);
nand U598 (N_598,N_515,N_482);
nand U599 (N_599,N_499,N_478);
nor U600 (N_600,N_582,N_560);
and U601 (N_601,N_598,N_527);
nor U602 (N_602,N_587,N_531);
nor U603 (N_603,N_558,N_562);
nor U604 (N_604,N_557,N_528);
or U605 (N_605,N_547,N_545);
and U606 (N_606,N_551,N_579);
and U607 (N_607,N_581,N_544);
nor U608 (N_608,N_566,N_572);
and U609 (N_609,N_596,N_585);
nand U610 (N_610,N_556,N_537);
nor U611 (N_611,N_567,N_561);
nor U612 (N_612,N_574,N_569);
nor U613 (N_613,N_535,N_563);
and U614 (N_614,N_588,N_534);
or U615 (N_615,N_526,N_536);
nand U616 (N_616,N_577,N_549);
or U617 (N_617,N_533,N_599);
nor U618 (N_618,N_594,N_559);
nand U619 (N_619,N_525,N_552);
or U620 (N_620,N_539,N_593);
or U621 (N_621,N_554,N_586);
nor U622 (N_622,N_592,N_550);
nand U623 (N_623,N_548,N_575);
nand U624 (N_624,N_584,N_589);
and U625 (N_625,N_529,N_564);
or U626 (N_626,N_597,N_530);
nor U627 (N_627,N_590,N_595);
nand U628 (N_628,N_532,N_583);
nand U629 (N_629,N_565,N_546);
or U630 (N_630,N_538,N_576);
nand U631 (N_631,N_543,N_571);
and U632 (N_632,N_580,N_541);
and U633 (N_633,N_568,N_553);
and U634 (N_634,N_542,N_573);
nand U635 (N_635,N_540,N_578);
nor U636 (N_636,N_570,N_555);
and U637 (N_637,N_591,N_567);
or U638 (N_638,N_580,N_530);
or U639 (N_639,N_547,N_542);
or U640 (N_640,N_566,N_583);
and U641 (N_641,N_596,N_592);
xor U642 (N_642,N_530,N_581);
and U643 (N_643,N_572,N_579);
nor U644 (N_644,N_559,N_579);
and U645 (N_645,N_595,N_556);
and U646 (N_646,N_536,N_543);
nor U647 (N_647,N_579,N_528);
xnor U648 (N_648,N_599,N_547);
or U649 (N_649,N_559,N_533);
nor U650 (N_650,N_543,N_574);
nor U651 (N_651,N_583,N_550);
and U652 (N_652,N_595,N_575);
nand U653 (N_653,N_562,N_560);
nand U654 (N_654,N_576,N_562);
nand U655 (N_655,N_571,N_595);
and U656 (N_656,N_581,N_582);
and U657 (N_657,N_567,N_599);
nand U658 (N_658,N_531,N_579);
and U659 (N_659,N_597,N_548);
or U660 (N_660,N_557,N_590);
and U661 (N_661,N_543,N_562);
nor U662 (N_662,N_528,N_597);
nand U663 (N_663,N_582,N_588);
nand U664 (N_664,N_561,N_542);
or U665 (N_665,N_575,N_584);
and U666 (N_666,N_570,N_550);
or U667 (N_667,N_583,N_591);
or U668 (N_668,N_547,N_595);
and U669 (N_669,N_592,N_553);
nor U670 (N_670,N_586,N_599);
and U671 (N_671,N_526,N_551);
and U672 (N_672,N_557,N_560);
nor U673 (N_673,N_555,N_533);
and U674 (N_674,N_545,N_552);
nand U675 (N_675,N_628,N_617);
or U676 (N_676,N_669,N_660);
nor U677 (N_677,N_621,N_664);
nand U678 (N_678,N_646,N_615);
and U679 (N_679,N_637,N_606);
nand U680 (N_680,N_661,N_663);
nand U681 (N_681,N_657,N_608);
or U682 (N_682,N_612,N_642);
nand U683 (N_683,N_619,N_659);
nand U684 (N_684,N_647,N_620);
nand U685 (N_685,N_600,N_668);
and U686 (N_686,N_633,N_611);
or U687 (N_687,N_671,N_601);
nand U688 (N_688,N_662,N_635);
and U689 (N_689,N_665,N_672);
nand U690 (N_690,N_618,N_610);
nor U691 (N_691,N_638,N_624);
nand U692 (N_692,N_616,N_605);
and U693 (N_693,N_652,N_629);
and U694 (N_694,N_653,N_667);
and U695 (N_695,N_632,N_666);
and U696 (N_696,N_648,N_656);
nand U697 (N_697,N_636,N_673);
and U698 (N_698,N_640,N_604);
or U699 (N_699,N_623,N_603);
and U700 (N_700,N_602,N_607);
nand U701 (N_701,N_609,N_631);
nand U702 (N_702,N_655,N_626);
and U703 (N_703,N_649,N_639);
or U704 (N_704,N_650,N_674);
nand U705 (N_705,N_641,N_614);
nand U706 (N_706,N_622,N_630);
nor U707 (N_707,N_644,N_658);
or U708 (N_708,N_627,N_613);
or U709 (N_709,N_634,N_651);
and U710 (N_710,N_654,N_625);
nand U711 (N_711,N_645,N_670);
nor U712 (N_712,N_643,N_656);
nor U713 (N_713,N_624,N_613);
nor U714 (N_714,N_621,N_641);
or U715 (N_715,N_602,N_654);
or U716 (N_716,N_607,N_614);
and U717 (N_717,N_616,N_670);
and U718 (N_718,N_647,N_670);
and U719 (N_719,N_653,N_664);
or U720 (N_720,N_631,N_654);
and U721 (N_721,N_600,N_648);
nor U722 (N_722,N_639,N_613);
and U723 (N_723,N_656,N_642);
and U724 (N_724,N_604,N_607);
or U725 (N_725,N_637,N_639);
nand U726 (N_726,N_631,N_630);
nor U727 (N_727,N_642,N_624);
nor U728 (N_728,N_609,N_603);
or U729 (N_729,N_601,N_670);
and U730 (N_730,N_600,N_607);
or U731 (N_731,N_652,N_640);
nor U732 (N_732,N_657,N_632);
nor U733 (N_733,N_666,N_641);
or U734 (N_734,N_612,N_616);
or U735 (N_735,N_645,N_610);
or U736 (N_736,N_638,N_621);
or U737 (N_737,N_619,N_607);
nand U738 (N_738,N_635,N_659);
nor U739 (N_739,N_620,N_651);
and U740 (N_740,N_645,N_649);
nand U741 (N_741,N_636,N_638);
and U742 (N_742,N_631,N_665);
nor U743 (N_743,N_617,N_648);
nor U744 (N_744,N_666,N_621);
nor U745 (N_745,N_635,N_664);
nor U746 (N_746,N_637,N_664);
nor U747 (N_747,N_630,N_666);
and U748 (N_748,N_612,N_602);
nand U749 (N_749,N_616,N_615);
or U750 (N_750,N_730,N_728);
nor U751 (N_751,N_729,N_737);
and U752 (N_752,N_712,N_704);
nand U753 (N_753,N_710,N_681);
nand U754 (N_754,N_718,N_719);
nand U755 (N_755,N_694,N_708);
nor U756 (N_756,N_740,N_697);
nand U757 (N_757,N_701,N_709);
or U758 (N_758,N_675,N_692);
nor U759 (N_759,N_723,N_748);
nand U760 (N_760,N_745,N_679);
nand U761 (N_761,N_683,N_749);
and U762 (N_762,N_680,N_682);
nand U763 (N_763,N_686,N_731);
or U764 (N_764,N_688,N_726);
or U765 (N_765,N_707,N_700);
nor U766 (N_766,N_744,N_720);
nor U767 (N_767,N_742,N_698);
or U768 (N_768,N_732,N_734);
nand U769 (N_769,N_727,N_690);
nor U770 (N_770,N_715,N_691);
or U771 (N_771,N_721,N_677);
nor U772 (N_772,N_703,N_747);
or U773 (N_773,N_724,N_706);
and U774 (N_774,N_687,N_739);
nand U775 (N_775,N_725,N_699);
and U776 (N_776,N_696,N_746);
nor U777 (N_777,N_693,N_738);
nor U778 (N_778,N_685,N_678);
nor U779 (N_779,N_684,N_695);
and U780 (N_780,N_713,N_743);
and U781 (N_781,N_711,N_722);
nor U782 (N_782,N_705,N_676);
and U783 (N_783,N_714,N_741);
or U784 (N_784,N_689,N_702);
or U785 (N_785,N_733,N_735);
nand U786 (N_786,N_736,N_717);
nand U787 (N_787,N_716,N_729);
and U788 (N_788,N_744,N_699);
or U789 (N_789,N_679,N_741);
nand U790 (N_790,N_699,N_687);
nor U791 (N_791,N_736,N_704);
or U792 (N_792,N_745,N_743);
nor U793 (N_793,N_697,N_695);
nand U794 (N_794,N_744,N_716);
nor U795 (N_795,N_716,N_689);
or U796 (N_796,N_706,N_729);
and U797 (N_797,N_692,N_680);
nor U798 (N_798,N_743,N_740);
or U799 (N_799,N_701,N_740);
and U800 (N_800,N_730,N_718);
nor U801 (N_801,N_709,N_714);
nand U802 (N_802,N_691,N_725);
or U803 (N_803,N_683,N_708);
or U804 (N_804,N_728,N_691);
or U805 (N_805,N_717,N_696);
nor U806 (N_806,N_698,N_708);
or U807 (N_807,N_725,N_731);
nand U808 (N_808,N_684,N_720);
and U809 (N_809,N_687,N_746);
nand U810 (N_810,N_709,N_723);
nor U811 (N_811,N_682,N_676);
nand U812 (N_812,N_725,N_677);
and U813 (N_813,N_683,N_709);
and U814 (N_814,N_737,N_716);
nor U815 (N_815,N_675,N_684);
and U816 (N_816,N_682,N_702);
and U817 (N_817,N_701,N_710);
nand U818 (N_818,N_735,N_732);
nand U819 (N_819,N_704,N_698);
nor U820 (N_820,N_702,N_735);
or U821 (N_821,N_707,N_693);
or U822 (N_822,N_708,N_725);
and U823 (N_823,N_727,N_707);
nand U824 (N_824,N_741,N_700);
nor U825 (N_825,N_811,N_795);
or U826 (N_826,N_796,N_792);
or U827 (N_827,N_814,N_770);
and U828 (N_828,N_807,N_800);
or U829 (N_829,N_752,N_753);
or U830 (N_830,N_763,N_824);
and U831 (N_831,N_809,N_816);
nand U832 (N_832,N_790,N_756);
and U833 (N_833,N_799,N_755);
nand U834 (N_834,N_784,N_821);
nor U835 (N_835,N_810,N_759);
and U836 (N_836,N_766,N_757);
nor U837 (N_837,N_822,N_771);
nand U838 (N_838,N_789,N_804);
nand U839 (N_839,N_778,N_802);
or U840 (N_840,N_791,N_794);
and U841 (N_841,N_761,N_793);
nor U842 (N_842,N_768,N_803);
and U843 (N_843,N_758,N_798);
nand U844 (N_844,N_783,N_750);
or U845 (N_845,N_808,N_805);
nor U846 (N_846,N_817,N_820);
nand U847 (N_847,N_787,N_754);
nor U848 (N_848,N_786,N_764);
nand U849 (N_849,N_801,N_773);
or U850 (N_850,N_772,N_806);
or U851 (N_851,N_813,N_797);
nand U852 (N_852,N_819,N_760);
xor U853 (N_853,N_812,N_815);
and U854 (N_854,N_785,N_769);
and U855 (N_855,N_762,N_774);
nand U856 (N_856,N_780,N_775);
nor U857 (N_857,N_777,N_767);
nor U858 (N_858,N_781,N_818);
nand U859 (N_859,N_751,N_776);
nor U860 (N_860,N_782,N_765);
or U861 (N_861,N_823,N_779);
nand U862 (N_862,N_788,N_798);
nand U863 (N_863,N_765,N_798);
nand U864 (N_864,N_792,N_809);
or U865 (N_865,N_750,N_823);
and U866 (N_866,N_816,N_807);
and U867 (N_867,N_817,N_753);
and U868 (N_868,N_814,N_764);
and U869 (N_869,N_783,N_795);
nor U870 (N_870,N_820,N_766);
and U871 (N_871,N_778,N_777);
nor U872 (N_872,N_801,N_804);
nand U873 (N_873,N_791,N_787);
or U874 (N_874,N_789,N_758);
or U875 (N_875,N_788,N_792);
nor U876 (N_876,N_805,N_815);
and U877 (N_877,N_770,N_780);
or U878 (N_878,N_770,N_758);
and U879 (N_879,N_757,N_810);
or U880 (N_880,N_772,N_811);
nor U881 (N_881,N_820,N_753);
nor U882 (N_882,N_783,N_819);
and U883 (N_883,N_790,N_800);
nand U884 (N_884,N_759,N_778);
or U885 (N_885,N_796,N_795);
nor U886 (N_886,N_782,N_820);
and U887 (N_887,N_792,N_763);
or U888 (N_888,N_784,N_812);
nor U889 (N_889,N_768,N_774);
and U890 (N_890,N_756,N_797);
nor U891 (N_891,N_789,N_763);
nor U892 (N_892,N_817,N_821);
and U893 (N_893,N_781,N_785);
or U894 (N_894,N_792,N_802);
nand U895 (N_895,N_767,N_816);
and U896 (N_896,N_752,N_792);
or U897 (N_897,N_808,N_754);
nand U898 (N_898,N_760,N_821);
or U899 (N_899,N_755,N_798);
xor U900 (N_900,N_843,N_850);
nand U901 (N_901,N_836,N_859);
and U902 (N_902,N_887,N_839);
nand U903 (N_903,N_861,N_832);
or U904 (N_904,N_898,N_825);
nand U905 (N_905,N_838,N_860);
or U906 (N_906,N_841,N_896);
or U907 (N_907,N_846,N_870);
or U908 (N_908,N_842,N_873);
or U909 (N_909,N_894,N_869);
nand U910 (N_910,N_875,N_837);
or U911 (N_911,N_888,N_835);
and U912 (N_912,N_874,N_857);
nand U913 (N_913,N_880,N_895);
nand U914 (N_914,N_897,N_872);
and U915 (N_915,N_866,N_852);
nor U916 (N_916,N_854,N_844);
nor U917 (N_917,N_881,N_868);
nor U918 (N_918,N_876,N_884);
and U919 (N_919,N_851,N_871);
nor U920 (N_920,N_856,N_885);
nor U921 (N_921,N_865,N_879);
nor U922 (N_922,N_891,N_886);
or U923 (N_923,N_826,N_877);
nand U924 (N_924,N_853,N_829);
nand U925 (N_925,N_867,N_834);
and U926 (N_926,N_833,N_830);
xnor U927 (N_927,N_899,N_858);
and U928 (N_928,N_892,N_864);
or U929 (N_929,N_849,N_840);
nand U930 (N_930,N_855,N_862);
nand U931 (N_931,N_890,N_883);
and U932 (N_932,N_831,N_848);
nand U933 (N_933,N_878,N_889);
nand U934 (N_934,N_893,N_827);
and U935 (N_935,N_863,N_828);
nor U936 (N_936,N_845,N_847);
nand U937 (N_937,N_882,N_896);
and U938 (N_938,N_827,N_881);
or U939 (N_939,N_861,N_849);
nand U940 (N_940,N_864,N_888);
and U941 (N_941,N_826,N_870);
and U942 (N_942,N_831,N_828);
and U943 (N_943,N_845,N_888);
nand U944 (N_944,N_841,N_837);
nor U945 (N_945,N_882,N_834);
nand U946 (N_946,N_876,N_841);
or U947 (N_947,N_854,N_868);
nand U948 (N_948,N_883,N_882);
or U949 (N_949,N_894,N_880);
nand U950 (N_950,N_830,N_895);
or U951 (N_951,N_846,N_859);
nor U952 (N_952,N_832,N_897);
nand U953 (N_953,N_894,N_877);
nand U954 (N_954,N_865,N_897);
xor U955 (N_955,N_831,N_849);
nand U956 (N_956,N_832,N_847);
and U957 (N_957,N_869,N_865);
nand U958 (N_958,N_890,N_896);
nor U959 (N_959,N_842,N_852);
nor U960 (N_960,N_846,N_839);
or U961 (N_961,N_839,N_876);
and U962 (N_962,N_871,N_827);
and U963 (N_963,N_847,N_895);
nand U964 (N_964,N_866,N_869);
or U965 (N_965,N_866,N_846);
or U966 (N_966,N_866,N_893);
nor U967 (N_967,N_896,N_831);
or U968 (N_968,N_843,N_839);
nor U969 (N_969,N_866,N_844);
and U970 (N_970,N_858,N_861);
nor U971 (N_971,N_854,N_873);
nand U972 (N_972,N_883,N_880);
or U973 (N_973,N_859,N_858);
nor U974 (N_974,N_829,N_836);
xnor U975 (N_975,N_943,N_971);
or U976 (N_976,N_944,N_915);
nor U977 (N_977,N_932,N_960);
and U978 (N_978,N_946,N_927);
nand U979 (N_979,N_925,N_939);
nand U980 (N_980,N_967,N_964);
or U981 (N_981,N_924,N_937);
or U982 (N_982,N_917,N_948);
nand U983 (N_983,N_938,N_968);
nor U984 (N_984,N_909,N_903);
or U985 (N_985,N_953,N_906);
nand U986 (N_986,N_931,N_929);
nor U987 (N_987,N_956,N_974);
or U988 (N_988,N_904,N_969);
and U989 (N_989,N_911,N_950);
nand U990 (N_990,N_942,N_907);
nor U991 (N_991,N_926,N_936);
nand U992 (N_992,N_908,N_973);
nor U993 (N_993,N_940,N_947);
and U994 (N_994,N_919,N_912);
nand U995 (N_995,N_902,N_928);
and U996 (N_996,N_935,N_955);
and U997 (N_997,N_901,N_961);
nand U998 (N_998,N_965,N_930);
or U999 (N_999,N_957,N_951);
nor U1000 (N_1000,N_923,N_966);
or U1001 (N_1001,N_922,N_949);
nand U1002 (N_1002,N_914,N_963);
nor U1003 (N_1003,N_972,N_920);
nand U1004 (N_1004,N_945,N_918);
or U1005 (N_1005,N_934,N_933);
or U1006 (N_1006,N_916,N_913);
and U1007 (N_1007,N_954,N_905);
and U1008 (N_1008,N_952,N_962);
nand U1009 (N_1009,N_921,N_910);
and U1010 (N_1010,N_941,N_970);
and U1011 (N_1011,N_958,N_900);
or U1012 (N_1012,N_959,N_926);
nand U1013 (N_1013,N_944,N_934);
and U1014 (N_1014,N_913,N_938);
and U1015 (N_1015,N_919,N_938);
or U1016 (N_1016,N_911,N_927);
or U1017 (N_1017,N_939,N_920);
and U1018 (N_1018,N_927,N_960);
and U1019 (N_1019,N_974,N_973);
nor U1020 (N_1020,N_945,N_913);
nand U1021 (N_1021,N_918,N_960);
nand U1022 (N_1022,N_973,N_925);
nor U1023 (N_1023,N_941,N_918);
nand U1024 (N_1024,N_920,N_922);
nand U1025 (N_1025,N_961,N_939);
or U1026 (N_1026,N_949,N_934);
and U1027 (N_1027,N_945,N_947);
nand U1028 (N_1028,N_935,N_902);
nand U1029 (N_1029,N_952,N_967);
or U1030 (N_1030,N_964,N_902);
nand U1031 (N_1031,N_973,N_940);
nand U1032 (N_1032,N_920,N_923);
and U1033 (N_1033,N_911,N_907);
nor U1034 (N_1034,N_912,N_938);
and U1035 (N_1035,N_904,N_970);
nor U1036 (N_1036,N_943,N_966);
or U1037 (N_1037,N_945,N_943);
or U1038 (N_1038,N_971,N_923);
nand U1039 (N_1039,N_943,N_969);
nand U1040 (N_1040,N_931,N_933);
nand U1041 (N_1041,N_948,N_936);
nor U1042 (N_1042,N_905,N_974);
nand U1043 (N_1043,N_948,N_932);
nor U1044 (N_1044,N_917,N_905);
and U1045 (N_1045,N_927,N_941);
nor U1046 (N_1046,N_962,N_949);
nand U1047 (N_1047,N_973,N_913);
nand U1048 (N_1048,N_967,N_902);
nor U1049 (N_1049,N_917,N_916);
nand U1050 (N_1050,N_1014,N_1024);
nand U1051 (N_1051,N_1040,N_1002);
and U1052 (N_1052,N_1003,N_999);
nand U1053 (N_1053,N_994,N_996);
nor U1054 (N_1054,N_1011,N_1017);
and U1055 (N_1055,N_1042,N_993);
nand U1056 (N_1056,N_983,N_986);
nor U1057 (N_1057,N_988,N_1048);
nand U1058 (N_1058,N_1044,N_979);
or U1059 (N_1059,N_1047,N_975);
or U1060 (N_1060,N_976,N_978);
nand U1061 (N_1061,N_1037,N_1009);
nor U1062 (N_1062,N_1018,N_1021);
nor U1063 (N_1063,N_1036,N_989);
nor U1064 (N_1064,N_1007,N_1046);
and U1065 (N_1065,N_1005,N_1041);
nor U1066 (N_1066,N_1029,N_1008);
nand U1067 (N_1067,N_1026,N_995);
nand U1068 (N_1068,N_981,N_985);
nor U1069 (N_1069,N_1028,N_1022);
nand U1070 (N_1070,N_984,N_1001);
or U1071 (N_1071,N_1016,N_1013);
nand U1072 (N_1072,N_1032,N_992);
and U1073 (N_1073,N_980,N_991);
or U1074 (N_1074,N_1049,N_1034);
nand U1075 (N_1075,N_1045,N_997);
or U1076 (N_1076,N_1010,N_1000);
nor U1077 (N_1077,N_1027,N_1023);
or U1078 (N_1078,N_987,N_1004);
nor U1079 (N_1079,N_1030,N_982);
nor U1080 (N_1080,N_1015,N_1012);
and U1081 (N_1081,N_990,N_1031);
and U1082 (N_1082,N_1035,N_1025);
nor U1083 (N_1083,N_1019,N_977);
nor U1084 (N_1084,N_1038,N_1039);
nand U1085 (N_1085,N_1006,N_1033);
or U1086 (N_1086,N_1020,N_1043);
and U1087 (N_1087,N_998,N_1028);
and U1088 (N_1088,N_1003,N_976);
or U1089 (N_1089,N_1027,N_1031);
xnor U1090 (N_1090,N_1043,N_982);
and U1091 (N_1091,N_985,N_1044);
and U1092 (N_1092,N_1025,N_1044);
nand U1093 (N_1093,N_1002,N_976);
nand U1094 (N_1094,N_1024,N_1018);
nor U1095 (N_1095,N_1039,N_975);
nand U1096 (N_1096,N_1031,N_1037);
or U1097 (N_1097,N_1031,N_1046);
and U1098 (N_1098,N_1019,N_1036);
nand U1099 (N_1099,N_1034,N_1042);
nor U1100 (N_1100,N_1016,N_1028);
nand U1101 (N_1101,N_1038,N_1025);
nor U1102 (N_1102,N_1028,N_985);
nor U1103 (N_1103,N_1035,N_1028);
nand U1104 (N_1104,N_1041,N_1043);
nor U1105 (N_1105,N_1019,N_1001);
nor U1106 (N_1106,N_1038,N_1021);
nor U1107 (N_1107,N_981,N_1048);
or U1108 (N_1108,N_1022,N_1046);
nor U1109 (N_1109,N_984,N_1020);
nor U1110 (N_1110,N_1030,N_989);
and U1111 (N_1111,N_987,N_1046);
or U1112 (N_1112,N_1022,N_1027);
or U1113 (N_1113,N_1035,N_1034);
or U1114 (N_1114,N_1012,N_982);
nor U1115 (N_1115,N_992,N_991);
or U1116 (N_1116,N_1025,N_977);
nand U1117 (N_1117,N_1033,N_1017);
or U1118 (N_1118,N_982,N_999);
nor U1119 (N_1119,N_1021,N_1045);
or U1120 (N_1120,N_976,N_1012);
nor U1121 (N_1121,N_1008,N_1022);
nand U1122 (N_1122,N_1001,N_983);
nor U1123 (N_1123,N_1038,N_993);
nand U1124 (N_1124,N_1048,N_1031);
nand U1125 (N_1125,N_1104,N_1051);
nor U1126 (N_1126,N_1110,N_1061);
and U1127 (N_1127,N_1066,N_1052);
or U1128 (N_1128,N_1090,N_1081);
and U1129 (N_1129,N_1123,N_1067);
or U1130 (N_1130,N_1055,N_1078);
and U1131 (N_1131,N_1088,N_1060);
nand U1132 (N_1132,N_1114,N_1120);
nand U1133 (N_1133,N_1062,N_1112);
and U1134 (N_1134,N_1094,N_1086);
or U1135 (N_1135,N_1108,N_1065);
or U1136 (N_1136,N_1124,N_1053);
nor U1137 (N_1137,N_1101,N_1099);
nor U1138 (N_1138,N_1115,N_1095);
and U1139 (N_1139,N_1113,N_1117);
nor U1140 (N_1140,N_1092,N_1068);
nand U1141 (N_1141,N_1084,N_1091);
and U1142 (N_1142,N_1076,N_1070);
and U1143 (N_1143,N_1057,N_1079);
xnor U1144 (N_1144,N_1058,N_1111);
nand U1145 (N_1145,N_1085,N_1100);
nor U1146 (N_1146,N_1121,N_1116);
or U1147 (N_1147,N_1119,N_1071);
and U1148 (N_1148,N_1082,N_1074);
or U1149 (N_1149,N_1109,N_1054);
nor U1150 (N_1150,N_1107,N_1122);
or U1151 (N_1151,N_1050,N_1080);
nand U1152 (N_1152,N_1063,N_1087);
nor U1153 (N_1153,N_1105,N_1097);
or U1154 (N_1154,N_1083,N_1089);
or U1155 (N_1155,N_1102,N_1106);
nand U1156 (N_1156,N_1118,N_1103);
and U1157 (N_1157,N_1093,N_1098);
nor U1158 (N_1158,N_1073,N_1077);
or U1159 (N_1159,N_1069,N_1075);
nor U1160 (N_1160,N_1056,N_1059);
and U1161 (N_1161,N_1064,N_1072);
nand U1162 (N_1162,N_1096,N_1063);
nand U1163 (N_1163,N_1124,N_1083);
or U1164 (N_1164,N_1057,N_1112);
nand U1165 (N_1165,N_1081,N_1054);
and U1166 (N_1166,N_1096,N_1059);
nor U1167 (N_1167,N_1088,N_1111);
nand U1168 (N_1168,N_1087,N_1062);
or U1169 (N_1169,N_1121,N_1067);
and U1170 (N_1170,N_1077,N_1053);
and U1171 (N_1171,N_1050,N_1109);
nor U1172 (N_1172,N_1106,N_1062);
or U1173 (N_1173,N_1050,N_1122);
or U1174 (N_1174,N_1059,N_1065);
nand U1175 (N_1175,N_1119,N_1073);
and U1176 (N_1176,N_1091,N_1081);
nor U1177 (N_1177,N_1099,N_1110);
and U1178 (N_1178,N_1089,N_1057);
and U1179 (N_1179,N_1106,N_1117);
and U1180 (N_1180,N_1075,N_1124);
or U1181 (N_1181,N_1057,N_1118);
nor U1182 (N_1182,N_1068,N_1081);
and U1183 (N_1183,N_1124,N_1086);
or U1184 (N_1184,N_1114,N_1075);
nand U1185 (N_1185,N_1091,N_1065);
or U1186 (N_1186,N_1050,N_1065);
or U1187 (N_1187,N_1110,N_1078);
or U1188 (N_1188,N_1084,N_1109);
nand U1189 (N_1189,N_1059,N_1114);
or U1190 (N_1190,N_1102,N_1087);
or U1191 (N_1191,N_1092,N_1105);
and U1192 (N_1192,N_1102,N_1055);
or U1193 (N_1193,N_1059,N_1116);
nor U1194 (N_1194,N_1052,N_1099);
and U1195 (N_1195,N_1064,N_1059);
nor U1196 (N_1196,N_1121,N_1081);
and U1197 (N_1197,N_1102,N_1064);
nor U1198 (N_1198,N_1101,N_1122);
or U1199 (N_1199,N_1060,N_1100);
or U1200 (N_1200,N_1193,N_1137);
nand U1201 (N_1201,N_1198,N_1176);
or U1202 (N_1202,N_1136,N_1186);
nand U1203 (N_1203,N_1132,N_1185);
nand U1204 (N_1204,N_1190,N_1152);
nand U1205 (N_1205,N_1135,N_1199);
nor U1206 (N_1206,N_1169,N_1160);
nand U1207 (N_1207,N_1195,N_1177);
nor U1208 (N_1208,N_1197,N_1138);
nor U1209 (N_1209,N_1155,N_1191);
xor U1210 (N_1210,N_1142,N_1173);
nand U1211 (N_1211,N_1146,N_1178);
or U1212 (N_1212,N_1148,N_1157);
or U1213 (N_1213,N_1140,N_1175);
nor U1214 (N_1214,N_1130,N_1150);
nor U1215 (N_1215,N_1188,N_1134);
or U1216 (N_1216,N_1127,N_1168);
nor U1217 (N_1217,N_1192,N_1171);
nor U1218 (N_1218,N_1158,N_1180);
nor U1219 (N_1219,N_1174,N_1179);
or U1220 (N_1220,N_1167,N_1147);
nor U1221 (N_1221,N_1166,N_1165);
nand U1222 (N_1222,N_1170,N_1145);
and U1223 (N_1223,N_1156,N_1129);
and U1224 (N_1224,N_1172,N_1125);
or U1225 (N_1225,N_1189,N_1161);
or U1226 (N_1226,N_1143,N_1159);
and U1227 (N_1227,N_1154,N_1163);
nor U1228 (N_1228,N_1128,N_1149);
nor U1229 (N_1229,N_1126,N_1162);
or U1230 (N_1230,N_1182,N_1184);
nor U1231 (N_1231,N_1194,N_1141);
nor U1232 (N_1232,N_1153,N_1187);
or U1233 (N_1233,N_1144,N_1151);
and U1234 (N_1234,N_1181,N_1183);
or U1235 (N_1235,N_1133,N_1139);
nor U1236 (N_1236,N_1196,N_1131);
nand U1237 (N_1237,N_1164,N_1132);
or U1238 (N_1238,N_1183,N_1151);
nand U1239 (N_1239,N_1176,N_1159);
nor U1240 (N_1240,N_1179,N_1194);
nand U1241 (N_1241,N_1168,N_1146);
nand U1242 (N_1242,N_1172,N_1199);
nor U1243 (N_1243,N_1185,N_1151);
and U1244 (N_1244,N_1141,N_1134);
or U1245 (N_1245,N_1186,N_1163);
nor U1246 (N_1246,N_1149,N_1177);
or U1247 (N_1247,N_1190,N_1127);
and U1248 (N_1248,N_1173,N_1149);
and U1249 (N_1249,N_1189,N_1193);
nor U1250 (N_1250,N_1198,N_1174);
and U1251 (N_1251,N_1179,N_1129);
and U1252 (N_1252,N_1195,N_1145);
xnor U1253 (N_1253,N_1145,N_1155);
nor U1254 (N_1254,N_1156,N_1132);
nand U1255 (N_1255,N_1196,N_1189);
nand U1256 (N_1256,N_1169,N_1165);
and U1257 (N_1257,N_1185,N_1138);
nand U1258 (N_1258,N_1177,N_1180);
and U1259 (N_1259,N_1130,N_1138);
nand U1260 (N_1260,N_1193,N_1169);
and U1261 (N_1261,N_1142,N_1190);
nand U1262 (N_1262,N_1193,N_1197);
and U1263 (N_1263,N_1169,N_1174);
nor U1264 (N_1264,N_1199,N_1126);
nor U1265 (N_1265,N_1194,N_1168);
or U1266 (N_1266,N_1174,N_1191);
and U1267 (N_1267,N_1187,N_1199);
or U1268 (N_1268,N_1199,N_1192);
nand U1269 (N_1269,N_1160,N_1157);
nor U1270 (N_1270,N_1194,N_1157);
nor U1271 (N_1271,N_1143,N_1136);
nor U1272 (N_1272,N_1179,N_1151);
or U1273 (N_1273,N_1164,N_1198);
nand U1274 (N_1274,N_1169,N_1168);
and U1275 (N_1275,N_1214,N_1220);
or U1276 (N_1276,N_1253,N_1256);
nand U1277 (N_1277,N_1259,N_1252);
nor U1278 (N_1278,N_1247,N_1250);
or U1279 (N_1279,N_1237,N_1274);
or U1280 (N_1280,N_1246,N_1216);
nor U1281 (N_1281,N_1263,N_1249);
nand U1282 (N_1282,N_1265,N_1210);
nand U1283 (N_1283,N_1255,N_1224);
or U1284 (N_1284,N_1257,N_1226);
nand U1285 (N_1285,N_1206,N_1262);
or U1286 (N_1286,N_1228,N_1215);
or U1287 (N_1287,N_1231,N_1230);
nor U1288 (N_1288,N_1201,N_1269);
or U1289 (N_1289,N_1258,N_1222);
nor U1290 (N_1290,N_1273,N_1208);
nor U1291 (N_1291,N_1232,N_1207);
nand U1292 (N_1292,N_1219,N_1209);
or U1293 (N_1293,N_1203,N_1213);
nor U1294 (N_1294,N_1248,N_1240);
and U1295 (N_1295,N_1233,N_1221);
nor U1296 (N_1296,N_1243,N_1217);
nand U1297 (N_1297,N_1200,N_1254);
nand U1298 (N_1298,N_1267,N_1238);
nor U1299 (N_1299,N_1239,N_1211);
xor U1300 (N_1300,N_1271,N_1225);
nor U1301 (N_1301,N_1235,N_1266);
and U1302 (N_1302,N_1218,N_1261);
nor U1303 (N_1303,N_1223,N_1236);
nand U1304 (N_1304,N_1244,N_1270);
nor U1305 (N_1305,N_1264,N_1212);
nor U1306 (N_1306,N_1227,N_1204);
or U1307 (N_1307,N_1268,N_1241);
and U1308 (N_1308,N_1272,N_1242);
nor U1309 (N_1309,N_1205,N_1202);
nand U1310 (N_1310,N_1234,N_1245);
or U1311 (N_1311,N_1260,N_1251);
nand U1312 (N_1312,N_1229,N_1265);
or U1313 (N_1313,N_1248,N_1249);
nor U1314 (N_1314,N_1217,N_1214);
and U1315 (N_1315,N_1262,N_1201);
and U1316 (N_1316,N_1209,N_1227);
or U1317 (N_1317,N_1259,N_1200);
or U1318 (N_1318,N_1260,N_1236);
and U1319 (N_1319,N_1236,N_1212);
or U1320 (N_1320,N_1228,N_1229);
and U1321 (N_1321,N_1264,N_1274);
nor U1322 (N_1322,N_1267,N_1268);
nand U1323 (N_1323,N_1228,N_1209);
nand U1324 (N_1324,N_1225,N_1205);
nor U1325 (N_1325,N_1264,N_1217);
nand U1326 (N_1326,N_1208,N_1254);
or U1327 (N_1327,N_1224,N_1218);
and U1328 (N_1328,N_1216,N_1267);
nor U1329 (N_1329,N_1232,N_1271);
and U1330 (N_1330,N_1224,N_1262);
or U1331 (N_1331,N_1226,N_1272);
nand U1332 (N_1332,N_1255,N_1256);
and U1333 (N_1333,N_1241,N_1258);
and U1334 (N_1334,N_1238,N_1260);
and U1335 (N_1335,N_1218,N_1214);
nor U1336 (N_1336,N_1247,N_1245);
and U1337 (N_1337,N_1210,N_1268);
or U1338 (N_1338,N_1269,N_1233);
and U1339 (N_1339,N_1272,N_1269);
or U1340 (N_1340,N_1235,N_1233);
nand U1341 (N_1341,N_1260,N_1219);
and U1342 (N_1342,N_1226,N_1210);
nor U1343 (N_1343,N_1256,N_1268);
or U1344 (N_1344,N_1221,N_1222);
or U1345 (N_1345,N_1216,N_1210);
nor U1346 (N_1346,N_1239,N_1271);
nor U1347 (N_1347,N_1202,N_1245);
nor U1348 (N_1348,N_1259,N_1270);
nand U1349 (N_1349,N_1247,N_1233);
and U1350 (N_1350,N_1347,N_1287);
nand U1351 (N_1351,N_1275,N_1313);
nand U1352 (N_1352,N_1283,N_1284);
and U1353 (N_1353,N_1339,N_1288);
or U1354 (N_1354,N_1315,N_1299);
nor U1355 (N_1355,N_1335,N_1334);
nor U1356 (N_1356,N_1331,N_1308);
nor U1357 (N_1357,N_1338,N_1297);
and U1358 (N_1358,N_1319,N_1342);
nor U1359 (N_1359,N_1281,N_1344);
nor U1360 (N_1360,N_1329,N_1300);
or U1361 (N_1361,N_1324,N_1290);
nand U1362 (N_1362,N_1305,N_1349);
nand U1363 (N_1363,N_1320,N_1298);
nor U1364 (N_1364,N_1337,N_1276);
and U1365 (N_1365,N_1279,N_1317);
nor U1366 (N_1366,N_1278,N_1291);
and U1367 (N_1367,N_1327,N_1332);
or U1368 (N_1368,N_1336,N_1285);
xnor U1369 (N_1369,N_1302,N_1312);
and U1370 (N_1370,N_1293,N_1340);
nor U1371 (N_1371,N_1306,N_1295);
nor U1372 (N_1372,N_1341,N_1343);
nand U1373 (N_1373,N_1328,N_1345);
or U1374 (N_1374,N_1321,N_1346);
and U1375 (N_1375,N_1307,N_1322);
and U1376 (N_1376,N_1277,N_1348);
nor U1377 (N_1377,N_1280,N_1323);
and U1378 (N_1378,N_1286,N_1309);
nand U1379 (N_1379,N_1294,N_1330);
and U1380 (N_1380,N_1318,N_1304);
nor U1381 (N_1381,N_1303,N_1282);
nand U1382 (N_1382,N_1296,N_1292);
or U1383 (N_1383,N_1310,N_1333);
and U1384 (N_1384,N_1289,N_1326);
or U1385 (N_1385,N_1316,N_1314);
or U1386 (N_1386,N_1311,N_1325);
nor U1387 (N_1387,N_1301,N_1275);
nor U1388 (N_1388,N_1336,N_1295);
nor U1389 (N_1389,N_1343,N_1333);
and U1390 (N_1390,N_1325,N_1321);
or U1391 (N_1391,N_1336,N_1305);
nand U1392 (N_1392,N_1330,N_1331);
nand U1393 (N_1393,N_1313,N_1328);
or U1394 (N_1394,N_1323,N_1301);
or U1395 (N_1395,N_1308,N_1346);
nand U1396 (N_1396,N_1315,N_1326);
nand U1397 (N_1397,N_1308,N_1333);
xor U1398 (N_1398,N_1313,N_1291);
nand U1399 (N_1399,N_1286,N_1281);
nand U1400 (N_1400,N_1279,N_1340);
and U1401 (N_1401,N_1330,N_1344);
or U1402 (N_1402,N_1288,N_1326);
and U1403 (N_1403,N_1324,N_1320);
nand U1404 (N_1404,N_1322,N_1280);
nor U1405 (N_1405,N_1299,N_1348);
nand U1406 (N_1406,N_1313,N_1278);
and U1407 (N_1407,N_1294,N_1319);
or U1408 (N_1408,N_1298,N_1319);
nand U1409 (N_1409,N_1284,N_1324);
nand U1410 (N_1410,N_1327,N_1337);
nand U1411 (N_1411,N_1330,N_1293);
nor U1412 (N_1412,N_1312,N_1339);
or U1413 (N_1413,N_1301,N_1288);
or U1414 (N_1414,N_1285,N_1282);
or U1415 (N_1415,N_1334,N_1284);
nand U1416 (N_1416,N_1282,N_1322);
nor U1417 (N_1417,N_1282,N_1294);
or U1418 (N_1418,N_1348,N_1312);
nor U1419 (N_1419,N_1345,N_1324);
nor U1420 (N_1420,N_1345,N_1300);
nand U1421 (N_1421,N_1280,N_1275);
and U1422 (N_1422,N_1276,N_1342);
and U1423 (N_1423,N_1284,N_1319);
and U1424 (N_1424,N_1306,N_1344);
and U1425 (N_1425,N_1423,N_1392);
or U1426 (N_1426,N_1370,N_1373);
nor U1427 (N_1427,N_1360,N_1400);
nor U1428 (N_1428,N_1354,N_1412);
or U1429 (N_1429,N_1351,N_1355);
or U1430 (N_1430,N_1368,N_1389);
nand U1431 (N_1431,N_1372,N_1383);
nor U1432 (N_1432,N_1363,N_1406);
and U1433 (N_1433,N_1409,N_1366);
xnor U1434 (N_1434,N_1410,N_1393);
or U1435 (N_1435,N_1407,N_1353);
and U1436 (N_1436,N_1413,N_1384);
or U1437 (N_1437,N_1405,N_1358);
or U1438 (N_1438,N_1402,N_1361);
nand U1439 (N_1439,N_1350,N_1378);
and U1440 (N_1440,N_1388,N_1369);
nand U1441 (N_1441,N_1422,N_1411);
and U1442 (N_1442,N_1352,N_1382);
and U1443 (N_1443,N_1379,N_1394);
or U1444 (N_1444,N_1401,N_1395);
and U1445 (N_1445,N_1424,N_1385);
and U1446 (N_1446,N_1415,N_1356);
nand U1447 (N_1447,N_1419,N_1416);
or U1448 (N_1448,N_1420,N_1398);
or U1449 (N_1449,N_1421,N_1377);
nand U1450 (N_1450,N_1417,N_1367);
nand U1451 (N_1451,N_1397,N_1396);
nor U1452 (N_1452,N_1359,N_1418);
nor U1453 (N_1453,N_1381,N_1376);
and U1454 (N_1454,N_1408,N_1365);
nand U1455 (N_1455,N_1364,N_1374);
nand U1456 (N_1456,N_1362,N_1391);
nand U1457 (N_1457,N_1414,N_1403);
nand U1458 (N_1458,N_1386,N_1399);
or U1459 (N_1459,N_1390,N_1380);
or U1460 (N_1460,N_1371,N_1357);
or U1461 (N_1461,N_1387,N_1404);
nor U1462 (N_1462,N_1375,N_1385);
and U1463 (N_1463,N_1374,N_1350);
nor U1464 (N_1464,N_1376,N_1421);
nor U1465 (N_1465,N_1402,N_1356);
nand U1466 (N_1466,N_1380,N_1384);
nand U1467 (N_1467,N_1371,N_1424);
or U1468 (N_1468,N_1409,N_1421);
nand U1469 (N_1469,N_1389,N_1374);
nand U1470 (N_1470,N_1390,N_1352);
and U1471 (N_1471,N_1352,N_1422);
or U1472 (N_1472,N_1407,N_1409);
and U1473 (N_1473,N_1359,N_1411);
and U1474 (N_1474,N_1372,N_1414);
and U1475 (N_1475,N_1366,N_1356);
and U1476 (N_1476,N_1384,N_1421);
nand U1477 (N_1477,N_1389,N_1350);
nor U1478 (N_1478,N_1414,N_1375);
nor U1479 (N_1479,N_1354,N_1405);
and U1480 (N_1480,N_1386,N_1392);
nor U1481 (N_1481,N_1414,N_1394);
and U1482 (N_1482,N_1386,N_1372);
nand U1483 (N_1483,N_1406,N_1403);
xor U1484 (N_1484,N_1415,N_1412);
and U1485 (N_1485,N_1374,N_1367);
nand U1486 (N_1486,N_1409,N_1385);
nand U1487 (N_1487,N_1351,N_1386);
and U1488 (N_1488,N_1357,N_1382);
nand U1489 (N_1489,N_1392,N_1367);
nand U1490 (N_1490,N_1422,N_1364);
nand U1491 (N_1491,N_1381,N_1392);
nand U1492 (N_1492,N_1412,N_1408);
nand U1493 (N_1493,N_1404,N_1359);
nand U1494 (N_1494,N_1378,N_1391);
nand U1495 (N_1495,N_1357,N_1373);
nor U1496 (N_1496,N_1390,N_1356);
nor U1497 (N_1497,N_1358,N_1381);
and U1498 (N_1498,N_1417,N_1354);
and U1499 (N_1499,N_1389,N_1371);
or U1500 (N_1500,N_1472,N_1476);
and U1501 (N_1501,N_1489,N_1473);
and U1502 (N_1502,N_1433,N_1493);
nor U1503 (N_1503,N_1474,N_1475);
nand U1504 (N_1504,N_1445,N_1442);
nor U1505 (N_1505,N_1468,N_1457);
nor U1506 (N_1506,N_1430,N_1479);
nand U1507 (N_1507,N_1483,N_1432);
and U1508 (N_1508,N_1448,N_1497);
nor U1509 (N_1509,N_1467,N_1494);
nand U1510 (N_1510,N_1495,N_1485);
or U1511 (N_1511,N_1449,N_1487);
nand U1512 (N_1512,N_1471,N_1438);
nand U1513 (N_1513,N_1431,N_1486);
nor U1514 (N_1514,N_1456,N_1429);
and U1515 (N_1515,N_1450,N_1490);
nor U1516 (N_1516,N_1481,N_1464);
nor U1517 (N_1517,N_1439,N_1466);
and U1518 (N_1518,N_1446,N_1480);
or U1519 (N_1519,N_1454,N_1434);
nand U1520 (N_1520,N_1435,N_1465);
and U1521 (N_1521,N_1478,N_1496);
nand U1522 (N_1522,N_1428,N_1499);
and U1523 (N_1523,N_1427,N_1425);
or U1524 (N_1524,N_1426,N_1462);
and U1525 (N_1525,N_1453,N_1443);
and U1526 (N_1526,N_1477,N_1459);
nor U1527 (N_1527,N_1460,N_1482);
and U1528 (N_1528,N_1444,N_1458);
nand U1529 (N_1529,N_1436,N_1440);
nand U1530 (N_1530,N_1437,N_1452);
nor U1531 (N_1531,N_1484,N_1447);
or U1532 (N_1532,N_1441,N_1470);
nor U1533 (N_1533,N_1461,N_1469);
or U1534 (N_1534,N_1488,N_1491);
nor U1535 (N_1535,N_1463,N_1498);
nor U1536 (N_1536,N_1455,N_1451);
nand U1537 (N_1537,N_1492,N_1442);
or U1538 (N_1538,N_1478,N_1497);
nand U1539 (N_1539,N_1437,N_1426);
nor U1540 (N_1540,N_1482,N_1452);
or U1541 (N_1541,N_1425,N_1491);
nand U1542 (N_1542,N_1461,N_1436);
nor U1543 (N_1543,N_1426,N_1428);
nor U1544 (N_1544,N_1435,N_1463);
and U1545 (N_1545,N_1473,N_1469);
and U1546 (N_1546,N_1475,N_1430);
and U1547 (N_1547,N_1473,N_1437);
and U1548 (N_1548,N_1450,N_1465);
nor U1549 (N_1549,N_1439,N_1425);
or U1550 (N_1550,N_1440,N_1472);
nand U1551 (N_1551,N_1431,N_1425);
nand U1552 (N_1552,N_1491,N_1492);
nor U1553 (N_1553,N_1427,N_1477);
nor U1554 (N_1554,N_1474,N_1493);
or U1555 (N_1555,N_1475,N_1478);
and U1556 (N_1556,N_1459,N_1473);
or U1557 (N_1557,N_1483,N_1481);
nand U1558 (N_1558,N_1494,N_1492);
and U1559 (N_1559,N_1473,N_1445);
or U1560 (N_1560,N_1482,N_1465);
nor U1561 (N_1561,N_1491,N_1440);
nand U1562 (N_1562,N_1484,N_1457);
nor U1563 (N_1563,N_1428,N_1454);
nand U1564 (N_1564,N_1464,N_1467);
nand U1565 (N_1565,N_1441,N_1427);
nor U1566 (N_1566,N_1426,N_1472);
nor U1567 (N_1567,N_1432,N_1492);
nor U1568 (N_1568,N_1444,N_1489);
nand U1569 (N_1569,N_1464,N_1474);
nand U1570 (N_1570,N_1431,N_1482);
or U1571 (N_1571,N_1446,N_1458);
and U1572 (N_1572,N_1492,N_1495);
nor U1573 (N_1573,N_1443,N_1432);
nor U1574 (N_1574,N_1486,N_1480);
nand U1575 (N_1575,N_1528,N_1549);
nand U1576 (N_1576,N_1547,N_1513);
nand U1577 (N_1577,N_1571,N_1570);
nor U1578 (N_1578,N_1502,N_1524);
nand U1579 (N_1579,N_1512,N_1506);
or U1580 (N_1580,N_1566,N_1569);
nand U1581 (N_1581,N_1522,N_1501);
and U1582 (N_1582,N_1533,N_1546);
and U1583 (N_1583,N_1523,N_1573);
nand U1584 (N_1584,N_1505,N_1520);
and U1585 (N_1585,N_1525,N_1510);
and U1586 (N_1586,N_1517,N_1529);
or U1587 (N_1587,N_1557,N_1553);
nor U1588 (N_1588,N_1564,N_1500);
or U1589 (N_1589,N_1530,N_1540);
nand U1590 (N_1590,N_1572,N_1516);
or U1591 (N_1591,N_1556,N_1511);
and U1592 (N_1592,N_1503,N_1514);
nand U1593 (N_1593,N_1507,N_1565);
nand U1594 (N_1594,N_1550,N_1574);
and U1595 (N_1595,N_1545,N_1521);
or U1596 (N_1596,N_1518,N_1541);
or U1597 (N_1597,N_1563,N_1539);
nand U1598 (N_1598,N_1515,N_1537);
nor U1599 (N_1599,N_1508,N_1551);
or U1600 (N_1600,N_1568,N_1561);
or U1601 (N_1601,N_1555,N_1509);
nor U1602 (N_1602,N_1504,N_1552);
nand U1603 (N_1603,N_1526,N_1535);
nor U1604 (N_1604,N_1536,N_1543);
or U1605 (N_1605,N_1527,N_1558);
nor U1606 (N_1606,N_1548,N_1534);
and U1607 (N_1607,N_1562,N_1560);
nor U1608 (N_1608,N_1519,N_1531);
and U1609 (N_1609,N_1542,N_1554);
or U1610 (N_1610,N_1544,N_1532);
nand U1611 (N_1611,N_1567,N_1559);
nor U1612 (N_1612,N_1538,N_1511);
and U1613 (N_1613,N_1517,N_1501);
nor U1614 (N_1614,N_1555,N_1535);
nor U1615 (N_1615,N_1572,N_1502);
or U1616 (N_1616,N_1527,N_1531);
and U1617 (N_1617,N_1561,N_1526);
and U1618 (N_1618,N_1509,N_1510);
nor U1619 (N_1619,N_1536,N_1554);
and U1620 (N_1620,N_1544,N_1553);
nor U1621 (N_1621,N_1547,N_1507);
nor U1622 (N_1622,N_1536,N_1556);
or U1623 (N_1623,N_1513,N_1525);
nor U1624 (N_1624,N_1549,N_1574);
and U1625 (N_1625,N_1564,N_1567);
nor U1626 (N_1626,N_1520,N_1569);
or U1627 (N_1627,N_1503,N_1548);
nand U1628 (N_1628,N_1572,N_1555);
nor U1629 (N_1629,N_1509,N_1529);
or U1630 (N_1630,N_1503,N_1552);
and U1631 (N_1631,N_1506,N_1550);
nand U1632 (N_1632,N_1510,N_1544);
nand U1633 (N_1633,N_1572,N_1536);
and U1634 (N_1634,N_1555,N_1537);
or U1635 (N_1635,N_1566,N_1531);
and U1636 (N_1636,N_1571,N_1541);
and U1637 (N_1637,N_1548,N_1539);
or U1638 (N_1638,N_1545,N_1520);
or U1639 (N_1639,N_1511,N_1559);
nand U1640 (N_1640,N_1506,N_1514);
nand U1641 (N_1641,N_1539,N_1516);
nand U1642 (N_1642,N_1553,N_1562);
and U1643 (N_1643,N_1530,N_1541);
and U1644 (N_1644,N_1566,N_1547);
or U1645 (N_1645,N_1509,N_1512);
nor U1646 (N_1646,N_1526,N_1544);
nor U1647 (N_1647,N_1548,N_1519);
and U1648 (N_1648,N_1506,N_1560);
nor U1649 (N_1649,N_1550,N_1544);
nor U1650 (N_1650,N_1618,N_1627);
and U1651 (N_1651,N_1608,N_1637);
nand U1652 (N_1652,N_1602,N_1646);
or U1653 (N_1653,N_1645,N_1624);
nand U1654 (N_1654,N_1613,N_1576);
nor U1655 (N_1655,N_1599,N_1600);
or U1656 (N_1656,N_1582,N_1580);
and U1657 (N_1657,N_1587,N_1579);
or U1658 (N_1658,N_1581,N_1594);
or U1659 (N_1659,N_1612,N_1577);
or U1660 (N_1660,N_1639,N_1605);
nor U1661 (N_1661,N_1621,N_1638);
and U1662 (N_1662,N_1597,N_1586);
nand U1663 (N_1663,N_1589,N_1575);
nor U1664 (N_1664,N_1635,N_1631);
nand U1665 (N_1665,N_1648,N_1607);
or U1666 (N_1666,N_1634,N_1584);
and U1667 (N_1667,N_1616,N_1578);
nand U1668 (N_1668,N_1595,N_1644);
and U1669 (N_1669,N_1628,N_1610);
and U1670 (N_1670,N_1626,N_1593);
or U1671 (N_1671,N_1643,N_1617);
or U1672 (N_1672,N_1640,N_1598);
nand U1673 (N_1673,N_1622,N_1588);
nor U1674 (N_1674,N_1629,N_1633);
or U1675 (N_1675,N_1641,N_1604);
and U1676 (N_1676,N_1636,N_1615);
nand U1677 (N_1677,N_1603,N_1630);
and U1678 (N_1678,N_1609,N_1583);
nand U1679 (N_1679,N_1647,N_1590);
nor U1680 (N_1680,N_1620,N_1601);
nor U1681 (N_1681,N_1642,N_1625);
and U1682 (N_1682,N_1614,N_1596);
or U1683 (N_1683,N_1592,N_1649);
and U1684 (N_1684,N_1632,N_1611);
nor U1685 (N_1685,N_1606,N_1623);
nor U1686 (N_1686,N_1591,N_1619);
and U1687 (N_1687,N_1585,N_1596);
and U1688 (N_1688,N_1637,N_1647);
or U1689 (N_1689,N_1587,N_1580);
or U1690 (N_1690,N_1612,N_1645);
and U1691 (N_1691,N_1582,N_1646);
and U1692 (N_1692,N_1591,N_1609);
and U1693 (N_1693,N_1640,N_1594);
nor U1694 (N_1694,N_1626,N_1635);
or U1695 (N_1695,N_1598,N_1607);
and U1696 (N_1696,N_1599,N_1598);
or U1697 (N_1697,N_1576,N_1598);
and U1698 (N_1698,N_1637,N_1636);
and U1699 (N_1699,N_1605,N_1647);
nor U1700 (N_1700,N_1577,N_1623);
and U1701 (N_1701,N_1648,N_1596);
or U1702 (N_1702,N_1637,N_1596);
nor U1703 (N_1703,N_1641,N_1588);
or U1704 (N_1704,N_1622,N_1575);
nand U1705 (N_1705,N_1637,N_1638);
and U1706 (N_1706,N_1584,N_1603);
or U1707 (N_1707,N_1589,N_1577);
nor U1708 (N_1708,N_1581,N_1605);
nor U1709 (N_1709,N_1601,N_1635);
nor U1710 (N_1710,N_1605,N_1606);
or U1711 (N_1711,N_1603,N_1582);
nand U1712 (N_1712,N_1602,N_1626);
and U1713 (N_1713,N_1649,N_1622);
or U1714 (N_1714,N_1600,N_1603);
and U1715 (N_1715,N_1644,N_1645);
nand U1716 (N_1716,N_1611,N_1606);
nand U1717 (N_1717,N_1578,N_1598);
nand U1718 (N_1718,N_1597,N_1643);
nor U1719 (N_1719,N_1613,N_1630);
nor U1720 (N_1720,N_1616,N_1634);
nor U1721 (N_1721,N_1608,N_1615);
nand U1722 (N_1722,N_1593,N_1577);
and U1723 (N_1723,N_1623,N_1632);
and U1724 (N_1724,N_1634,N_1633);
or U1725 (N_1725,N_1719,N_1695);
nor U1726 (N_1726,N_1717,N_1650);
nor U1727 (N_1727,N_1721,N_1697);
and U1728 (N_1728,N_1704,N_1699);
and U1729 (N_1729,N_1657,N_1690);
or U1730 (N_1730,N_1675,N_1662);
nand U1731 (N_1731,N_1714,N_1689);
or U1732 (N_1732,N_1718,N_1679);
nand U1733 (N_1733,N_1659,N_1668);
and U1734 (N_1734,N_1674,N_1684);
nand U1735 (N_1735,N_1709,N_1687);
nor U1736 (N_1736,N_1683,N_1722);
nand U1737 (N_1737,N_1670,N_1661);
and U1738 (N_1738,N_1715,N_1658);
nor U1739 (N_1739,N_1681,N_1691);
nand U1740 (N_1740,N_1677,N_1685);
and U1741 (N_1741,N_1724,N_1678);
and U1742 (N_1742,N_1676,N_1688);
nand U1743 (N_1743,N_1655,N_1696);
and U1744 (N_1744,N_1652,N_1713);
nor U1745 (N_1745,N_1651,N_1694);
or U1746 (N_1746,N_1692,N_1700);
nor U1747 (N_1747,N_1663,N_1667);
nand U1748 (N_1748,N_1708,N_1660);
nor U1749 (N_1749,N_1707,N_1716);
nand U1750 (N_1750,N_1712,N_1710);
nor U1751 (N_1751,N_1720,N_1706);
or U1752 (N_1752,N_1664,N_1671);
and U1753 (N_1753,N_1693,N_1654);
nor U1754 (N_1754,N_1673,N_1723);
nand U1755 (N_1755,N_1682,N_1702);
nand U1756 (N_1756,N_1680,N_1703);
nor U1757 (N_1757,N_1665,N_1672);
nand U1758 (N_1758,N_1653,N_1705);
or U1759 (N_1759,N_1698,N_1669);
nand U1760 (N_1760,N_1701,N_1686);
and U1761 (N_1761,N_1666,N_1656);
and U1762 (N_1762,N_1711,N_1674);
nand U1763 (N_1763,N_1689,N_1713);
nand U1764 (N_1764,N_1720,N_1683);
nand U1765 (N_1765,N_1650,N_1697);
xnor U1766 (N_1766,N_1673,N_1670);
nor U1767 (N_1767,N_1676,N_1661);
nand U1768 (N_1768,N_1666,N_1679);
nor U1769 (N_1769,N_1690,N_1720);
nor U1770 (N_1770,N_1652,N_1659);
and U1771 (N_1771,N_1667,N_1718);
or U1772 (N_1772,N_1717,N_1687);
or U1773 (N_1773,N_1717,N_1692);
nor U1774 (N_1774,N_1678,N_1710);
or U1775 (N_1775,N_1669,N_1703);
or U1776 (N_1776,N_1718,N_1720);
or U1777 (N_1777,N_1651,N_1698);
nor U1778 (N_1778,N_1707,N_1706);
nand U1779 (N_1779,N_1697,N_1668);
nand U1780 (N_1780,N_1708,N_1687);
or U1781 (N_1781,N_1656,N_1650);
or U1782 (N_1782,N_1682,N_1677);
and U1783 (N_1783,N_1668,N_1715);
nor U1784 (N_1784,N_1718,N_1659);
and U1785 (N_1785,N_1675,N_1694);
and U1786 (N_1786,N_1672,N_1654);
nand U1787 (N_1787,N_1668,N_1685);
and U1788 (N_1788,N_1695,N_1666);
nand U1789 (N_1789,N_1682,N_1716);
and U1790 (N_1790,N_1683,N_1712);
nor U1791 (N_1791,N_1677,N_1683);
nand U1792 (N_1792,N_1704,N_1701);
nand U1793 (N_1793,N_1684,N_1675);
or U1794 (N_1794,N_1723,N_1665);
or U1795 (N_1795,N_1658,N_1687);
and U1796 (N_1796,N_1679,N_1669);
and U1797 (N_1797,N_1656,N_1667);
nor U1798 (N_1798,N_1653,N_1665);
or U1799 (N_1799,N_1710,N_1677);
or U1800 (N_1800,N_1774,N_1757);
nand U1801 (N_1801,N_1733,N_1781);
nor U1802 (N_1802,N_1770,N_1787);
nand U1803 (N_1803,N_1795,N_1755);
nor U1804 (N_1804,N_1732,N_1785);
and U1805 (N_1805,N_1739,N_1740);
nor U1806 (N_1806,N_1764,N_1746);
nor U1807 (N_1807,N_1744,N_1793);
nor U1808 (N_1808,N_1737,N_1762);
and U1809 (N_1809,N_1741,N_1751);
and U1810 (N_1810,N_1756,N_1745);
nand U1811 (N_1811,N_1731,N_1782);
nor U1812 (N_1812,N_1771,N_1761);
and U1813 (N_1813,N_1767,N_1777);
and U1814 (N_1814,N_1799,N_1738);
and U1815 (N_1815,N_1736,N_1754);
and U1816 (N_1816,N_1766,N_1749);
nand U1817 (N_1817,N_1769,N_1778);
or U1818 (N_1818,N_1752,N_1760);
and U1819 (N_1819,N_1789,N_1788);
nand U1820 (N_1820,N_1790,N_1758);
nor U1821 (N_1821,N_1725,N_1776);
or U1822 (N_1822,N_1742,N_1779);
or U1823 (N_1823,N_1797,N_1775);
nand U1824 (N_1824,N_1796,N_1759);
and U1825 (N_1825,N_1780,N_1791);
and U1826 (N_1826,N_1753,N_1747);
nand U1827 (N_1827,N_1792,N_1794);
nor U1828 (N_1828,N_1783,N_1729);
nor U1829 (N_1829,N_1750,N_1763);
nand U1830 (N_1830,N_1730,N_1735);
nor U1831 (N_1831,N_1734,N_1786);
and U1832 (N_1832,N_1727,N_1765);
and U1833 (N_1833,N_1798,N_1768);
nand U1834 (N_1834,N_1773,N_1728);
nor U1835 (N_1835,N_1748,N_1784);
or U1836 (N_1836,N_1726,N_1772);
or U1837 (N_1837,N_1743,N_1757);
and U1838 (N_1838,N_1773,N_1757);
nand U1839 (N_1839,N_1764,N_1791);
or U1840 (N_1840,N_1792,N_1734);
nor U1841 (N_1841,N_1766,N_1789);
nor U1842 (N_1842,N_1740,N_1799);
nand U1843 (N_1843,N_1740,N_1734);
or U1844 (N_1844,N_1798,N_1780);
or U1845 (N_1845,N_1731,N_1780);
or U1846 (N_1846,N_1796,N_1767);
and U1847 (N_1847,N_1730,N_1770);
nor U1848 (N_1848,N_1771,N_1747);
and U1849 (N_1849,N_1782,N_1789);
and U1850 (N_1850,N_1797,N_1785);
nor U1851 (N_1851,N_1760,N_1740);
and U1852 (N_1852,N_1760,N_1751);
or U1853 (N_1853,N_1798,N_1748);
and U1854 (N_1854,N_1779,N_1727);
nand U1855 (N_1855,N_1776,N_1769);
and U1856 (N_1856,N_1750,N_1766);
and U1857 (N_1857,N_1729,N_1747);
and U1858 (N_1858,N_1765,N_1730);
nand U1859 (N_1859,N_1776,N_1755);
or U1860 (N_1860,N_1740,N_1765);
nor U1861 (N_1861,N_1731,N_1761);
xnor U1862 (N_1862,N_1751,N_1781);
or U1863 (N_1863,N_1743,N_1786);
or U1864 (N_1864,N_1759,N_1729);
xor U1865 (N_1865,N_1745,N_1741);
nand U1866 (N_1866,N_1785,N_1747);
nor U1867 (N_1867,N_1749,N_1771);
nand U1868 (N_1868,N_1784,N_1766);
or U1869 (N_1869,N_1734,N_1737);
or U1870 (N_1870,N_1741,N_1795);
nand U1871 (N_1871,N_1772,N_1797);
or U1872 (N_1872,N_1737,N_1795);
or U1873 (N_1873,N_1743,N_1785);
and U1874 (N_1874,N_1798,N_1791);
nor U1875 (N_1875,N_1824,N_1811);
nand U1876 (N_1876,N_1800,N_1815);
or U1877 (N_1877,N_1820,N_1842);
and U1878 (N_1878,N_1864,N_1869);
or U1879 (N_1879,N_1867,N_1808);
or U1880 (N_1880,N_1821,N_1816);
nand U1881 (N_1881,N_1831,N_1865);
nand U1882 (N_1882,N_1841,N_1839);
nand U1883 (N_1883,N_1849,N_1830);
nand U1884 (N_1884,N_1857,N_1818);
and U1885 (N_1885,N_1833,N_1827);
and U1886 (N_1886,N_1840,N_1826);
nor U1887 (N_1887,N_1859,N_1870);
nand U1888 (N_1888,N_1806,N_1866);
or U1889 (N_1889,N_1862,N_1814);
or U1890 (N_1890,N_1810,N_1868);
or U1891 (N_1891,N_1874,N_1858);
or U1892 (N_1892,N_1838,N_1871);
nor U1893 (N_1893,N_1837,N_1863);
or U1894 (N_1894,N_1846,N_1835);
nor U1895 (N_1895,N_1812,N_1804);
nor U1896 (N_1896,N_1834,N_1817);
nor U1897 (N_1897,N_1850,N_1802);
nand U1898 (N_1898,N_1809,N_1805);
or U1899 (N_1899,N_1825,N_1853);
and U1900 (N_1900,N_1836,N_1848);
nand U1901 (N_1901,N_1844,N_1801);
nor U1902 (N_1902,N_1873,N_1819);
nand U1903 (N_1903,N_1860,N_1822);
and U1904 (N_1904,N_1813,N_1845);
and U1905 (N_1905,N_1855,N_1861);
and U1906 (N_1906,N_1851,N_1854);
and U1907 (N_1907,N_1872,N_1856);
nand U1908 (N_1908,N_1843,N_1823);
or U1909 (N_1909,N_1828,N_1807);
nand U1910 (N_1910,N_1803,N_1829);
nand U1911 (N_1911,N_1832,N_1852);
and U1912 (N_1912,N_1847,N_1800);
or U1913 (N_1913,N_1840,N_1800);
and U1914 (N_1914,N_1812,N_1861);
or U1915 (N_1915,N_1804,N_1851);
or U1916 (N_1916,N_1819,N_1870);
nand U1917 (N_1917,N_1808,N_1801);
nor U1918 (N_1918,N_1800,N_1818);
nand U1919 (N_1919,N_1838,N_1825);
nand U1920 (N_1920,N_1839,N_1806);
or U1921 (N_1921,N_1867,N_1830);
nand U1922 (N_1922,N_1812,N_1859);
nand U1923 (N_1923,N_1852,N_1807);
nor U1924 (N_1924,N_1819,N_1827);
and U1925 (N_1925,N_1864,N_1802);
nand U1926 (N_1926,N_1846,N_1842);
or U1927 (N_1927,N_1834,N_1841);
nor U1928 (N_1928,N_1820,N_1867);
nor U1929 (N_1929,N_1866,N_1861);
xnor U1930 (N_1930,N_1834,N_1803);
nand U1931 (N_1931,N_1863,N_1830);
and U1932 (N_1932,N_1823,N_1840);
or U1933 (N_1933,N_1803,N_1816);
nor U1934 (N_1934,N_1810,N_1829);
nor U1935 (N_1935,N_1815,N_1857);
or U1936 (N_1936,N_1848,N_1829);
or U1937 (N_1937,N_1849,N_1857);
or U1938 (N_1938,N_1814,N_1801);
and U1939 (N_1939,N_1863,N_1850);
or U1940 (N_1940,N_1852,N_1848);
or U1941 (N_1941,N_1825,N_1844);
and U1942 (N_1942,N_1868,N_1803);
and U1943 (N_1943,N_1818,N_1827);
nor U1944 (N_1944,N_1840,N_1844);
or U1945 (N_1945,N_1823,N_1834);
and U1946 (N_1946,N_1830,N_1828);
or U1947 (N_1947,N_1833,N_1811);
nor U1948 (N_1948,N_1856,N_1861);
nand U1949 (N_1949,N_1858,N_1848);
or U1950 (N_1950,N_1921,N_1917);
nor U1951 (N_1951,N_1876,N_1889);
nand U1952 (N_1952,N_1924,N_1900);
nand U1953 (N_1953,N_1909,N_1937);
and U1954 (N_1954,N_1911,N_1920);
nor U1955 (N_1955,N_1894,N_1925);
nor U1956 (N_1956,N_1904,N_1930);
and U1957 (N_1957,N_1929,N_1932);
nor U1958 (N_1958,N_1877,N_1885);
nor U1959 (N_1959,N_1880,N_1934);
nor U1960 (N_1960,N_1914,N_1933);
or U1961 (N_1961,N_1918,N_1893);
nor U1962 (N_1962,N_1940,N_1888);
nand U1963 (N_1963,N_1936,N_1903);
and U1964 (N_1964,N_1946,N_1891);
and U1965 (N_1965,N_1898,N_1901);
or U1966 (N_1966,N_1916,N_1890);
nor U1967 (N_1967,N_1927,N_1944);
nand U1968 (N_1968,N_1886,N_1947);
nand U1969 (N_1969,N_1912,N_1941);
nor U1970 (N_1970,N_1949,N_1881);
or U1971 (N_1971,N_1910,N_1943);
or U1972 (N_1972,N_1895,N_1919);
nor U1973 (N_1973,N_1931,N_1906);
or U1974 (N_1974,N_1899,N_1948);
nand U1975 (N_1975,N_1882,N_1935);
nand U1976 (N_1976,N_1878,N_1913);
nand U1977 (N_1977,N_1945,N_1887);
and U1978 (N_1978,N_1908,N_1905);
nor U1979 (N_1979,N_1923,N_1875);
nand U1980 (N_1980,N_1938,N_1879);
or U1981 (N_1981,N_1942,N_1922);
or U1982 (N_1982,N_1928,N_1897);
nand U1983 (N_1983,N_1883,N_1884);
and U1984 (N_1984,N_1892,N_1907);
and U1985 (N_1985,N_1902,N_1896);
nor U1986 (N_1986,N_1939,N_1915);
nor U1987 (N_1987,N_1926,N_1911);
nand U1988 (N_1988,N_1883,N_1894);
nand U1989 (N_1989,N_1918,N_1897);
nor U1990 (N_1990,N_1923,N_1876);
nor U1991 (N_1991,N_1886,N_1877);
or U1992 (N_1992,N_1921,N_1908);
or U1993 (N_1993,N_1922,N_1896);
and U1994 (N_1994,N_1878,N_1898);
or U1995 (N_1995,N_1913,N_1911);
or U1996 (N_1996,N_1936,N_1923);
nand U1997 (N_1997,N_1883,N_1887);
nand U1998 (N_1998,N_1928,N_1922);
xnor U1999 (N_1999,N_1881,N_1888);
and U2000 (N_2000,N_1899,N_1901);
nand U2001 (N_2001,N_1910,N_1914);
and U2002 (N_2002,N_1882,N_1924);
and U2003 (N_2003,N_1921,N_1923);
and U2004 (N_2004,N_1890,N_1937);
or U2005 (N_2005,N_1896,N_1947);
or U2006 (N_2006,N_1926,N_1933);
and U2007 (N_2007,N_1894,N_1880);
or U2008 (N_2008,N_1892,N_1929);
nor U2009 (N_2009,N_1914,N_1918);
nor U2010 (N_2010,N_1892,N_1927);
nand U2011 (N_2011,N_1889,N_1907);
or U2012 (N_2012,N_1904,N_1941);
nand U2013 (N_2013,N_1939,N_1937);
nand U2014 (N_2014,N_1923,N_1885);
and U2015 (N_2015,N_1892,N_1895);
nand U2016 (N_2016,N_1937,N_1920);
or U2017 (N_2017,N_1919,N_1909);
and U2018 (N_2018,N_1881,N_1941);
nand U2019 (N_2019,N_1889,N_1936);
nor U2020 (N_2020,N_1927,N_1935);
nand U2021 (N_2021,N_1885,N_1930);
or U2022 (N_2022,N_1891,N_1913);
or U2023 (N_2023,N_1946,N_1898);
nand U2024 (N_2024,N_1938,N_1932);
and U2025 (N_2025,N_2015,N_1950);
nand U2026 (N_2026,N_1951,N_1955);
and U2027 (N_2027,N_2022,N_1987);
nor U2028 (N_2028,N_1982,N_1977);
or U2029 (N_2029,N_1989,N_1962);
or U2030 (N_2030,N_1973,N_1970);
or U2031 (N_2031,N_1958,N_1980);
nand U2032 (N_2032,N_1998,N_2021);
and U2033 (N_2033,N_1996,N_1992);
and U2034 (N_2034,N_2013,N_2004);
nand U2035 (N_2035,N_1984,N_2024);
or U2036 (N_2036,N_2023,N_1956);
nor U2037 (N_2037,N_2007,N_1993);
or U2038 (N_2038,N_1957,N_2002);
nand U2039 (N_2039,N_1974,N_1981);
nor U2040 (N_2040,N_2000,N_1988);
nand U2041 (N_2041,N_1986,N_2020);
and U2042 (N_2042,N_1966,N_1979);
or U2043 (N_2043,N_2005,N_2018);
xnor U2044 (N_2044,N_1972,N_1968);
nor U2045 (N_2045,N_1960,N_1995);
or U2046 (N_2046,N_1969,N_1976);
nand U2047 (N_2047,N_2009,N_1952);
nor U2048 (N_2048,N_1997,N_1985);
and U2049 (N_2049,N_2011,N_1975);
or U2050 (N_2050,N_2006,N_1990);
nand U2051 (N_2051,N_2014,N_1959);
and U2052 (N_2052,N_1999,N_1991);
or U2053 (N_2053,N_2010,N_1961);
and U2054 (N_2054,N_1967,N_1994);
nand U2055 (N_2055,N_1964,N_1983);
nand U2056 (N_2056,N_1954,N_1965);
nor U2057 (N_2057,N_2019,N_2017);
nor U2058 (N_2058,N_2016,N_1978);
or U2059 (N_2059,N_2003,N_2008);
or U2060 (N_2060,N_2001,N_1963);
xnor U2061 (N_2061,N_1971,N_1953);
xor U2062 (N_2062,N_2012,N_1950);
nand U2063 (N_2063,N_1955,N_2003);
nor U2064 (N_2064,N_1954,N_2000);
nor U2065 (N_2065,N_2000,N_1953);
nor U2066 (N_2066,N_2002,N_2021);
xor U2067 (N_2067,N_2019,N_1981);
nor U2068 (N_2068,N_1982,N_2008);
nor U2069 (N_2069,N_2020,N_1972);
nand U2070 (N_2070,N_2006,N_1983);
and U2071 (N_2071,N_1977,N_1951);
nand U2072 (N_2072,N_1999,N_1951);
nor U2073 (N_2073,N_2023,N_1953);
nor U2074 (N_2074,N_2012,N_2018);
or U2075 (N_2075,N_2001,N_1982);
nand U2076 (N_2076,N_1954,N_1953);
and U2077 (N_2077,N_2016,N_2005);
nor U2078 (N_2078,N_2007,N_1963);
and U2079 (N_2079,N_1983,N_2017);
nand U2080 (N_2080,N_1990,N_1996);
and U2081 (N_2081,N_1959,N_1964);
nand U2082 (N_2082,N_1968,N_1980);
nand U2083 (N_2083,N_1984,N_1979);
or U2084 (N_2084,N_1972,N_1960);
nand U2085 (N_2085,N_2024,N_1966);
and U2086 (N_2086,N_1964,N_1962);
and U2087 (N_2087,N_1985,N_2011);
nand U2088 (N_2088,N_2005,N_2010);
or U2089 (N_2089,N_1955,N_2010);
and U2090 (N_2090,N_1961,N_1970);
nand U2091 (N_2091,N_2013,N_1970);
nor U2092 (N_2092,N_1983,N_1969);
nand U2093 (N_2093,N_1980,N_1974);
nor U2094 (N_2094,N_1980,N_2016);
xor U2095 (N_2095,N_1959,N_1983);
and U2096 (N_2096,N_2000,N_1972);
nand U2097 (N_2097,N_1975,N_1954);
or U2098 (N_2098,N_1995,N_1992);
or U2099 (N_2099,N_1982,N_2006);
nor U2100 (N_2100,N_2085,N_2078);
and U2101 (N_2101,N_2079,N_2056);
or U2102 (N_2102,N_2096,N_2083);
and U2103 (N_2103,N_2034,N_2051);
and U2104 (N_2104,N_2072,N_2077);
nor U2105 (N_2105,N_2059,N_2087);
nand U2106 (N_2106,N_2026,N_2065);
or U2107 (N_2107,N_2029,N_2094);
nand U2108 (N_2108,N_2047,N_2097);
nand U2109 (N_2109,N_2074,N_2063);
or U2110 (N_2110,N_2060,N_2042);
nand U2111 (N_2111,N_2032,N_2061);
or U2112 (N_2112,N_2095,N_2088);
nor U2113 (N_2113,N_2076,N_2046);
or U2114 (N_2114,N_2052,N_2071);
nor U2115 (N_2115,N_2067,N_2038);
or U2116 (N_2116,N_2058,N_2027);
nor U2117 (N_2117,N_2073,N_2036);
and U2118 (N_2118,N_2090,N_2098);
and U2119 (N_2119,N_2080,N_2082);
or U2120 (N_2120,N_2070,N_2064);
and U2121 (N_2121,N_2093,N_2057);
or U2122 (N_2122,N_2062,N_2035);
or U2123 (N_2123,N_2048,N_2025);
nor U2124 (N_2124,N_2066,N_2037);
nand U2125 (N_2125,N_2068,N_2055);
and U2126 (N_2126,N_2040,N_2069);
or U2127 (N_2127,N_2091,N_2053);
and U2128 (N_2128,N_2039,N_2075);
or U2129 (N_2129,N_2033,N_2031);
and U2130 (N_2130,N_2049,N_2081);
nand U2131 (N_2131,N_2030,N_2092);
or U2132 (N_2132,N_2084,N_2044);
nor U2133 (N_2133,N_2054,N_2028);
or U2134 (N_2134,N_2050,N_2045);
nor U2135 (N_2135,N_2043,N_2089);
nor U2136 (N_2136,N_2041,N_2086);
nand U2137 (N_2137,N_2099,N_2088);
nor U2138 (N_2138,N_2036,N_2092);
nor U2139 (N_2139,N_2035,N_2076);
nand U2140 (N_2140,N_2051,N_2046);
and U2141 (N_2141,N_2095,N_2052);
and U2142 (N_2142,N_2083,N_2058);
nor U2143 (N_2143,N_2071,N_2078);
nand U2144 (N_2144,N_2058,N_2055);
nor U2145 (N_2145,N_2026,N_2078);
nor U2146 (N_2146,N_2040,N_2052);
and U2147 (N_2147,N_2051,N_2064);
nor U2148 (N_2148,N_2099,N_2060);
nand U2149 (N_2149,N_2071,N_2031);
or U2150 (N_2150,N_2096,N_2067);
and U2151 (N_2151,N_2053,N_2068);
nand U2152 (N_2152,N_2096,N_2074);
and U2153 (N_2153,N_2043,N_2061);
nor U2154 (N_2154,N_2061,N_2046);
nand U2155 (N_2155,N_2085,N_2092);
or U2156 (N_2156,N_2031,N_2082);
nand U2157 (N_2157,N_2050,N_2067);
or U2158 (N_2158,N_2092,N_2080);
and U2159 (N_2159,N_2098,N_2025);
nor U2160 (N_2160,N_2036,N_2063);
or U2161 (N_2161,N_2089,N_2047);
and U2162 (N_2162,N_2065,N_2083);
or U2163 (N_2163,N_2088,N_2038);
and U2164 (N_2164,N_2030,N_2061);
nand U2165 (N_2165,N_2097,N_2079);
or U2166 (N_2166,N_2065,N_2038);
nor U2167 (N_2167,N_2088,N_2056);
nor U2168 (N_2168,N_2085,N_2091);
nor U2169 (N_2169,N_2026,N_2097);
nor U2170 (N_2170,N_2037,N_2060);
nand U2171 (N_2171,N_2063,N_2043);
nor U2172 (N_2172,N_2090,N_2060);
or U2173 (N_2173,N_2071,N_2039);
and U2174 (N_2174,N_2032,N_2064);
nor U2175 (N_2175,N_2133,N_2138);
nor U2176 (N_2176,N_2103,N_2158);
nand U2177 (N_2177,N_2117,N_2129);
nand U2178 (N_2178,N_2113,N_2152);
nor U2179 (N_2179,N_2110,N_2105);
or U2180 (N_2180,N_2121,N_2155);
nand U2181 (N_2181,N_2116,N_2130);
or U2182 (N_2182,N_2128,N_2170);
and U2183 (N_2183,N_2101,N_2114);
nand U2184 (N_2184,N_2115,N_2125);
or U2185 (N_2185,N_2111,N_2123);
nor U2186 (N_2186,N_2166,N_2150);
or U2187 (N_2187,N_2104,N_2160);
nor U2188 (N_2188,N_2161,N_2109);
nand U2189 (N_2189,N_2157,N_2174);
and U2190 (N_2190,N_2102,N_2132);
nor U2191 (N_2191,N_2100,N_2119);
or U2192 (N_2192,N_2134,N_2145);
or U2193 (N_2193,N_2147,N_2149);
nand U2194 (N_2194,N_2124,N_2146);
nor U2195 (N_2195,N_2107,N_2137);
or U2196 (N_2196,N_2141,N_2159);
nand U2197 (N_2197,N_2168,N_2106);
nor U2198 (N_2198,N_2165,N_2140);
nand U2199 (N_2199,N_2126,N_2167);
nand U2200 (N_2200,N_2122,N_2148);
or U2201 (N_2201,N_2156,N_2144);
or U2202 (N_2202,N_2118,N_2153);
nor U2203 (N_2203,N_2154,N_2131);
and U2204 (N_2204,N_2112,N_2169);
and U2205 (N_2205,N_2163,N_2172);
or U2206 (N_2206,N_2136,N_2151);
nand U2207 (N_2207,N_2108,N_2135);
nand U2208 (N_2208,N_2173,N_2127);
nor U2209 (N_2209,N_2171,N_2139);
or U2210 (N_2210,N_2164,N_2142);
nand U2211 (N_2211,N_2162,N_2143);
and U2212 (N_2212,N_2120,N_2160);
and U2213 (N_2213,N_2104,N_2161);
or U2214 (N_2214,N_2144,N_2145);
or U2215 (N_2215,N_2158,N_2119);
or U2216 (N_2216,N_2168,N_2117);
and U2217 (N_2217,N_2149,N_2166);
nor U2218 (N_2218,N_2133,N_2123);
nand U2219 (N_2219,N_2156,N_2159);
and U2220 (N_2220,N_2158,N_2170);
nor U2221 (N_2221,N_2107,N_2157);
nor U2222 (N_2222,N_2109,N_2155);
nand U2223 (N_2223,N_2132,N_2170);
nand U2224 (N_2224,N_2130,N_2168);
or U2225 (N_2225,N_2134,N_2156);
nand U2226 (N_2226,N_2128,N_2143);
nor U2227 (N_2227,N_2169,N_2114);
or U2228 (N_2228,N_2153,N_2129);
nor U2229 (N_2229,N_2129,N_2173);
nand U2230 (N_2230,N_2130,N_2158);
nor U2231 (N_2231,N_2169,N_2146);
nand U2232 (N_2232,N_2126,N_2134);
and U2233 (N_2233,N_2148,N_2135);
and U2234 (N_2234,N_2160,N_2168);
and U2235 (N_2235,N_2131,N_2158);
nand U2236 (N_2236,N_2157,N_2172);
nand U2237 (N_2237,N_2167,N_2159);
or U2238 (N_2238,N_2172,N_2127);
and U2239 (N_2239,N_2172,N_2123);
nor U2240 (N_2240,N_2103,N_2135);
nand U2241 (N_2241,N_2106,N_2112);
and U2242 (N_2242,N_2158,N_2102);
or U2243 (N_2243,N_2145,N_2128);
and U2244 (N_2244,N_2154,N_2104);
nor U2245 (N_2245,N_2121,N_2158);
nand U2246 (N_2246,N_2141,N_2144);
nand U2247 (N_2247,N_2155,N_2135);
nor U2248 (N_2248,N_2162,N_2132);
or U2249 (N_2249,N_2151,N_2138);
nor U2250 (N_2250,N_2217,N_2220);
and U2251 (N_2251,N_2231,N_2216);
and U2252 (N_2252,N_2242,N_2221);
nor U2253 (N_2253,N_2239,N_2190);
nand U2254 (N_2254,N_2248,N_2212);
xor U2255 (N_2255,N_2246,N_2204);
nand U2256 (N_2256,N_2227,N_2215);
nor U2257 (N_2257,N_2200,N_2247);
nand U2258 (N_2258,N_2222,N_2178);
and U2259 (N_2259,N_2186,N_2223);
nor U2260 (N_2260,N_2233,N_2238);
and U2261 (N_2261,N_2224,N_2201);
nor U2262 (N_2262,N_2209,N_2214);
nor U2263 (N_2263,N_2218,N_2240);
nand U2264 (N_2264,N_2185,N_2203);
nor U2265 (N_2265,N_2191,N_2189);
nand U2266 (N_2266,N_2243,N_2177);
and U2267 (N_2267,N_2241,N_2194);
and U2268 (N_2268,N_2188,N_2187);
and U2269 (N_2269,N_2175,N_2226);
nand U2270 (N_2270,N_2234,N_2228);
and U2271 (N_2271,N_2202,N_2198);
and U2272 (N_2272,N_2181,N_2225);
nand U2273 (N_2273,N_2207,N_2229);
and U2274 (N_2274,N_2195,N_2249);
nor U2275 (N_2275,N_2208,N_2219);
and U2276 (N_2276,N_2236,N_2193);
nand U2277 (N_2277,N_2232,N_2210);
and U2278 (N_2278,N_2205,N_2179);
nor U2279 (N_2279,N_2180,N_2182);
or U2280 (N_2280,N_2237,N_2230);
or U2281 (N_2281,N_2176,N_2211);
nor U2282 (N_2282,N_2235,N_2245);
and U2283 (N_2283,N_2197,N_2184);
and U2284 (N_2284,N_2192,N_2199);
nand U2285 (N_2285,N_2196,N_2206);
nor U2286 (N_2286,N_2213,N_2244);
nor U2287 (N_2287,N_2183,N_2215);
nor U2288 (N_2288,N_2209,N_2183);
and U2289 (N_2289,N_2249,N_2192);
or U2290 (N_2290,N_2193,N_2243);
or U2291 (N_2291,N_2209,N_2202);
and U2292 (N_2292,N_2215,N_2237);
nor U2293 (N_2293,N_2212,N_2205);
or U2294 (N_2294,N_2190,N_2199);
or U2295 (N_2295,N_2197,N_2248);
nor U2296 (N_2296,N_2221,N_2183);
and U2297 (N_2297,N_2243,N_2223);
nor U2298 (N_2298,N_2213,N_2239);
nand U2299 (N_2299,N_2243,N_2179);
or U2300 (N_2300,N_2190,N_2178);
and U2301 (N_2301,N_2216,N_2218);
nand U2302 (N_2302,N_2184,N_2186);
and U2303 (N_2303,N_2230,N_2231);
nand U2304 (N_2304,N_2204,N_2235);
nor U2305 (N_2305,N_2232,N_2240);
nor U2306 (N_2306,N_2209,N_2178);
nor U2307 (N_2307,N_2183,N_2205);
nand U2308 (N_2308,N_2207,N_2241);
nor U2309 (N_2309,N_2212,N_2193);
nor U2310 (N_2310,N_2183,N_2227);
nor U2311 (N_2311,N_2193,N_2214);
nand U2312 (N_2312,N_2198,N_2183);
or U2313 (N_2313,N_2179,N_2211);
and U2314 (N_2314,N_2245,N_2217);
and U2315 (N_2315,N_2199,N_2231);
and U2316 (N_2316,N_2178,N_2189);
nand U2317 (N_2317,N_2196,N_2230);
nand U2318 (N_2318,N_2217,N_2229);
nor U2319 (N_2319,N_2198,N_2219);
or U2320 (N_2320,N_2206,N_2238);
and U2321 (N_2321,N_2241,N_2247);
xnor U2322 (N_2322,N_2245,N_2226);
and U2323 (N_2323,N_2232,N_2248);
nor U2324 (N_2324,N_2193,N_2181);
and U2325 (N_2325,N_2271,N_2251);
or U2326 (N_2326,N_2286,N_2272);
and U2327 (N_2327,N_2263,N_2259);
nand U2328 (N_2328,N_2267,N_2309);
or U2329 (N_2329,N_2289,N_2288);
nor U2330 (N_2330,N_2266,N_2306);
nand U2331 (N_2331,N_2300,N_2297);
or U2332 (N_2332,N_2301,N_2275);
nand U2333 (N_2333,N_2285,N_2257);
nand U2334 (N_2334,N_2305,N_2299);
and U2335 (N_2335,N_2296,N_2256);
or U2336 (N_2336,N_2254,N_2302);
or U2337 (N_2337,N_2294,N_2321);
or U2338 (N_2338,N_2320,N_2313);
and U2339 (N_2339,N_2274,N_2304);
and U2340 (N_2340,N_2269,N_2255);
or U2341 (N_2341,N_2282,N_2322);
nor U2342 (N_2342,N_2250,N_2287);
and U2343 (N_2343,N_2261,N_2292);
or U2344 (N_2344,N_2298,N_2277);
and U2345 (N_2345,N_2315,N_2310);
nor U2346 (N_2346,N_2253,N_2281);
nand U2347 (N_2347,N_2324,N_2308);
nand U2348 (N_2348,N_2270,N_2279);
and U2349 (N_2349,N_2268,N_2284);
and U2350 (N_2350,N_2323,N_2252);
or U2351 (N_2351,N_2283,N_2318);
or U2352 (N_2352,N_2290,N_2280);
and U2353 (N_2353,N_2293,N_2307);
or U2354 (N_2354,N_2278,N_2276);
or U2355 (N_2355,N_2314,N_2317);
nor U2356 (N_2356,N_2295,N_2258);
nand U2357 (N_2357,N_2264,N_2291);
and U2358 (N_2358,N_2262,N_2303);
nor U2359 (N_2359,N_2260,N_2312);
nand U2360 (N_2360,N_2319,N_2273);
and U2361 (N_2361,N_2316,N_2265);
nor U2362 (N_2362,N_2311,N_2314);
nand U2363 (N_2363,N_2266,N_2278);
or U2364 (N_2364,N_2297,N_2275);
nand U2365 (N_2365,N_2270,N_2269);
nor U2366 (N_2366,N_2289,N_2299);
and U2367 (N_2367,N_2314,N_2301);
or U2368 (N_2368,N_2265,N_2272);
nand U2369 (N_2369,N_2315,N_2283);
and U2370 (N_2370,N_2285,N_2291);
nor U2371 (N_2371,N_2269,N_2264);
nor U2372 (N_2372,N_2293,N_2319);
and U2373 (N_2373,N_2316,N_2308);
nor U2374 (N_2374,N_2259,N_2308);
and U2375 (N_2375,N_2303,N_2311);
nor U2376 (N_2376,N_2273,N_2321);
nor U2377 (N_2377,N_2300,N_2308);
or U2378 (N_2378,N_2321,N_2323);
or U2379 (N_2379,N_2287,N_2254);
nor U2380 (N_2380,N_2289,N_2290);
or U2381 (N_2381,N_2253,N_2289);
and U2382 (N_2382,N_2251,N_2301);
nor U2383 (N_2383,N_2272,N_2263);
or U2384 (N_2384,N_2316,N_2305);
nor U2385 (N_2385,N_2289,N_2267);
and U2386 (N_2386,N_2283,N_2268);
nor U2387 (N_2387,N_2262,N_2250);
or U2388 (N_2388,N_2269,N_2311);
nand U2389 (N_2389,N_2320,N_2294);
and U2390 (N_2390,N_2266,N_2267);
and U2391 (N_2391,N_2274,N_2261);
and U2392 (N_2392,N_2261,N_2267);
or U2393 (N_2393,N_2299,N_2266);
nor U2394 (N_2394,N_2315,N_2293);
nand U2395 (N_2395,N_2263,N_2268);
or U2396 (N_2396,N_2273,N_2316);
xor U2397 (N_2397,N_2321,N_2310);
nand U2398 (N_2398,N_2281,N_2301);
and U2399 (N_2399,N_2298,N_2288);
nand U2400 (N_2400,N_2349,N_2366);
nand U2401 (N_2401,N_2399,N_2359);
nor U2402 (N_2402,N_2350,N_2344);
and U2403 (N_2403,N_2326,N_2390);
or U2404 (N_2404,N_2378,N_2361);
nor U2405 (N_2405,N_2340,N_2391);
or U2406 (N_2406,N_2379,N_2398);
or U2407 (N_2407,N_2395,N_2362);
nor U2408 (N_2408,N_2346,N_2354);
nor U2409 (N_2409,N_2355,N_2338);
nor U2410 (N_2410,N_2364,N_2363);
nand U2411 (N_2411,N_2392,N_2375);
or U2412 (N_2412,N_2384,N_2393);
nand U2413 (N_2413,N_2358,N_2357);
nand U2414 (N_2414,N_2333,N_2342);
and U2415 (N_2415,N_2337,N_2351);
or U2416 (N_2416,N_2341,N_2329);
or U2417 (N_2417,N_2352,N_2397);
and U2418 (N_2418,N_2331,N_2386);
nand U2419 (N_2419,N_2381,N_2365);
and U2420 (N_2420,N_2353,N_2382);
or U2421 (N_2421,N_2383,N_2387);
or U2422 (N_2422,N_2377,N_2336);
and U2423 (N_2423,N_2325,N_2335);
nor U2424 (N_2424,N_2396,N_2327);
nor U2425 (N_2425,N_2394,N_2369);
nand U2426 (N_2426,N_2388,N_2380);
nor U2427 (N_2427,N_2374,N_2389);
nand U2428 (N_2428,N_2339,N_2367);
and U2429 (N_2429,N_2372,N_2343);
nand U2430 (N_2430,N_2345,N_2370);
and U2431 (N_2431,N_2373,N_2330);
or U2432 (N_2432,N_2368,N_2332);
and U2433 (N_2433,N_2334,N_2360);
or U2434 (N_2434,N_2348,N_2385);
nor U2435 (N_2435,N_2328,N_2371);
and U2436 (N_2436,N_2376,N_2347);
and U2437 (N_2437,N_2356,N_2333);
nor U2438 (N_2438,N_2331,N_2392);
nor U2439 (N_2439,N_2392,N_2384);
or U2440 (N_2440,N_2381,N_2368);
nand U2441 (N_2441,N_2366,N_2397);
and U2442 (N_2442,N_2384,N_2382);
nand U2443 (N_2443,N_2376,N_2334);
nor U2444 (N_2444,N_2348,N_2342);
or U2445 (N_2445,N_2371,N_2352);
and U2446 (N_2446,N_2372,N_2396);
and U2447 (N_2447,N_2370,N_2332);
nand U2448 (N_2448,N_2382,N_2375);
and U2449 (N_2449,N_2341,N_2345);
and U2450 (N_2450,N_2386,N_2338);
and U2451 (N_2451,N_2363,N_2378);
and U2452 (N_2452,N_2386,N_2394);
and U2453 (N_2453,N_2357,N_2331);
or U2454 (N_2454,N_2359,N_2349);
and U2455 (N_2455,N_2336,N_2395);
or U2456 (N_2456,N_2362,N_2356);
nor U2457 (N_2457,N_2361,N_2391);
nand U2458 (N_2458,N_2373,N_2363);
and U2459 (N_2459,N_2386,N_2367);
or U2460 (N_2460,N_2368,N_2367);
nor U2461 (N_2461,N_2329,N_2338);
xnor U2462 (N_2462,N_2351,N_2328);
xnor U2463 (N_2463,N_2353,N_2351);
nand U2464 (N_2464,N_2356,N_2345);
and U2465 (N_2465,N_2355,N_2379);
and U2466 (N_2466,N_2353,N_2348);
nand U2467 (N_2467,N_2388,N_2377);
and U2468 (N_2468,N_2370,N_2394);
nor U2469 (N_2469,N_2390,N_2327);
and U2470 (N_2470,N_2397,N_2383);
and U2471 (N_2471,N_2342,N_2349);
nor U2472 (N_2472,N_2391,N_2331);
nand U2473 (N_2473,N_2393,N_2327);
or U2474 (N_2474,N_2347,N_2354);
nand U2475 (N_2475,N_2430,N_2401);
and U2476 (N_2476,N_2452,N_2444);
and U2477 (N_2477,N_2420,N_2458);
and U2478 (N_2478,N_2465,N_2436);
and U2479 (N_2479,N_2445,N_2432);
or U2480 (N_2480,N_2414,N_2433);
or U2481 (N_2481,N_2450,N_2426);
or U2482 (N_2482,N_2466,N_2428);
nor U2483 (N_2483,N_2459,N_2408);
and U2484 (N_2484,N_2447,N_2413);
nor U2485 (N_2485,N_2441,N_2409);
nand U2486 (N_2486,N_2440,N_2470);
and U2487 (N_2487,N_2422,N_2404);
nand U2488 (N_2488,N_2443,N_2423);
and U2489 (N_2489,N_2427,N_2457);
and U2490 (N_2490,N_2403,N_2410);
or U2491 (N_2491,N_2461,N_2415);
nand U2492 (N_2492,N_2446,N_2406);
nand U2493 (N_2493,N_2454,N_2417);
nand U2494 (N_2494,N_2431,N_2456);
and U2495 (N_2495,N_2471,N_2451);
nand U2496 (N_2496,N_2405,N_2469);
xnor U2497 (N_2497,N_2439,N_2418);
and U2498 (N_2498,N_2460,N_2402);
and U2499 (N_2499,N_2425,N_2424);
xor U2500 (N_2500,N_2435,N_2411);
nor U2501 (N_2501,N_2438,N_2472);
nand U2502 (N_2502,N_2419,N_2437);
or U2503 (N_2503,N_2468,N_2467);
nor U2504 (N_2504,N_2448,N_2453);
nor U2505 (N_2505,N_2421,N_2462);
or U2506 (N_2506,N_2474,N_2429);
nor U2507 (N_2507,N_2473,N_2407);
and U2508 (N_2508,N_2442,N_2434);
or U2509 (N_2509,N_2464,N_2463);
nor U2510 (N_2510,N_2449,N_2416);
or U2511 (N_2511,N_2400,N_2455);
nor U2512 (N_2512,N_2412,N_2434);
nor U2513 (N_2513,N_2429,N_2462);
and U2514 (N_2514,N_2449,N_2450);
or U2515 (N_2515,N_2459,N_2462);
and U2516 (N_2516,N_2424,N_2419);
and U2517 (N_2517,N_2469,N_2430);
or U2518 (N_2518,N_2411,N_2417);
nor U2519 (N_2519,N_2423,N_2410);
or U2520 (N_2520,N_2409,N_2422);
or U2521 (N_2521,N_2455,N_2471);
nand U2522 (N_2522,N_2472,N_2423);
nand U2523 (N_2523,N_2458,N_2474);
or U2524 (N_2524,N_2422,N_2474);
nor U2525 (N_2525,N_2440,N_2436);
nand U2526 (N_2526,N_2466,N_2460);
nor U2527 (N_2527,N_2429,N_2436);
nand U2528 (N_2528,N_2432,N_2470);
nand U2529 (N_2529,N_2427,N_2455);
and U2530 (N_2530,N_2447,N_2474);
and U2531 (N_2531,N_2457,N_2424);
or U2532 (N_2532,N_2446,N_2425);
xnor U2533 (N_2533,N_2405,N_2403);
nand U2534 (N_2534,N_2418,N_2470);
nand U2535 (N_2535,N_2443,N_2468);
and U2536 (N_2536,N_2459,N_2404);
and U2537 (N_2537,N_2464,N_2428);
or U2538 (N_2538,N_2432,N_2407);
nand U2539 (N_2539,N_2444,N_2405);
nor U2540 (N_2540,N_2474,N_2463);
nand U2541 (N_2541,N_2440,N_2451);
and U2542 (N_2542,N_2444,N_2468);
or U2543 (N_2543,N_2461,N_2405);
nand U2544 (N_2544,N_2461,N_2451);
or U2545 (N_2545,N_2452,N_2459);
and U2546 (N_2546,N_2441,N_2434);
or U2547 (N_2547,N_2442,N_2454);
or U2548 (N_2548,N_2431,N_2455);
and U2549 (N_2549,N_2406,N_2402);
or U2550 (N_2550,N_2529,N_2525);
nand U2551 (N_2551,N_2512,N_2516);
nand U2552 (N_2552,N_2517,N_2532);
or U2553 (N_2553,N_2487,N_2544);
nor U2554 (N_2554,N_2542,N_2493);
or U2555 (N_2555,N_2479,N_2481);
or U2556 (N_2556,N_2477,N_2527);
or U2557 (N_2557,N_2496,N_2475);
nand U2558 (N_2558,N_2518,N_2480);
nand U2559 (N_2559,N_2491,N_2483);
and U2560 (N_2560,N_2526,N_2519);
nor U2561 (N_2561,N_2485,N_2503);
or U2562 (N_2562,N_2488,N_2507);
or U2563 (N_2563,N_2520,N_2509);
and U2564 (N_2564,N_2500,N_2549);
or U2565 (N_2565,N_2514,N_2522);
or U2566 (N_2566,N_2504,N_2494);
or U2567 (N_2567,N_2510,N_2533);
and U2568 (N_2568,N_2538,N_2535);
nor U2569 (N_2569,N_2476,N_2501);
nor U2570 (N_2570,N_2548,N_2534);
nor U2571 (N_2571,N_2508,N_2545);
nor U2572 (N_2572,N_2521,N_2543);
nor U2573 (N_2573,N_2511,N_2482);
nand U2574 (N_2574,N_2523,N_2528);
and U2575 (N_2575,N_2540,N_2486);
nand U2576 (N_2576,N_2489,N_2515);
nor U2577 (N_2577,N_2490,N_2513);
nor U2578 (N_2578,N_2484,N_2547);
or U2579 (N_2579,N_2531,N_2530);
or U2580 (N_2580,N_2546,N_2497);
nand U2581 (N_2581,N_2524,N_2499);
or U2582 (N_2582,N_2506,N_2537);
nor U2583 (N_2583,N_2502,N_2492);
nor U2584 (N_2584,N_2539,N_2505);
and U2585 (N_2585,N_2541,N_2495);
nand U2586 (N_2586,N_2536,N_2478);
nor U2587 (N_2587,N_2498,N_2543);
or U2588 (N_2588,N_2505,N_2493);
and U2589 (N_2589,N_2482,N_2541);
nor U2590 (N_2590,N_2519,N_2493);
or U2591 (N_2591,N_2549,N_2493);
nor U2592 (N_2592,N_2526,N_2523);
nor U2593 (N_2593,N_2524,N_2546);
and U2594 (N_2594,N_2483,N_2475);
nor U2595 (N_2595,N_2523,N_2515);
nand U2596 (N_2596,N_2504,N_2545);
xnor U2597 (N_2597,N_2507,N_2501);
or U2598 (N_2598,N_2517,N_2475);
nor U2599 (N_2599,N_2543,N_2528);
and U2600 (N_2600,N_2478,N_2527);
nor U2601 (N_2601,N_2524,N_2490);
nor U2602 (N_2602,N_2548,N_2494);
or U2603 (N_2603,N_2494,N_2476);
and U2604 (N_2604,N_2542,N_2528);
and U2605 (N_2605,N_2545,N_2512);
nand U2606 (N_2606,N_2524,N_2512);
nand U2607 (N_2607,N_2523,N_2518);
and U2608 (N_2608,N_2542,N_2506);
nor U2609 (N_2609,N_2480,N_2516);
or U2610 (N_2610,N_2492,N_2480);
nor U2611 (N_2611,N_2547,N_2480);
nand U2612 (N_2612,N_2487,N_2522);
or U2613 (N_2613,N_2509,N_2548);
nor U2614 (N_2614,N_2496,N_2480);
nor U2615 (N_2615,N_2496,N_2503);
and U2616 (N_2616,N_2480,N_2504);
or U2617 (N_2617,N_2505,N_2542);
or U2618 (N_2618,N_2489,N_2514);
or U2619 (N_2619,N_2546,N_2548);
or U2620 (N_2620,N_2500,N_2505);
or U2621 (N_2621,N_2529,N_2516);
or U2622 (N_2622,N_2547,N_2527);
nor U2623 (N_2623,N_2481,N_2475);
nand U2624 (N_2624,N_2503,N_2519);
and U2625 (N_2625,N_2592,N_2561);
nand U2626 (N_2626,N_2602,N_2562);
and U2627 (N_2627,N_2573,N_2570);
nand U2628 (N_2628,N_2621,N_2610);
nand U2629 (N_2629,N_2567,N_2571);
or U2630 (N_2630,N_2558,N_2555);
nor U2631 (N_2631,N_2553,N_2593);
or U2632 (N_2632,N_2560,N_2590);
nand U2633 (N_2633,N_2589,N_2582);
nor U2634 (N_2634,N_2597,N_2576);
or U2635 (N_2635,N_2591,N_2584);
and U2636 (N_2636,N_2557,N_2565);
and U2637 (N_2637,N_2566,N_2550);
and U2638 (N_2638,N_2568,N_2616);
nand U2639 (N_2639,N_2603,N_2594);
and U2640 (N_2640,N_2605,N_2579);
and U2641 (N_2641,N_2585,N_2618);
nand U2642 (N_2642,N_2607,N_2596);
nand U2643 (N_2643,N_2624,N_2600);
nand U2644 (N_2644,N_2564,N_2572);
or U2645 (N_2645,N_2613,N_2604);
and U2646 (N_2646,N_2583,N_2612);
nand U2647 (N_2647,N_2575,N_2588);
nand U2648 (N_2648,N_2559,N_2554);
or U2649 (N_2649,N_2577,N_2620);
nor U2650 (N_2650,N_2623,N_2587);
nor U2651 (N_2651,N_2586,N_2574);
nand U2652 (N_2652,N_2601,N_2599);
nand U2653 (N_2653,N_2569,N_2611);
nor U2654 (N_2654,N_2606,N_2580);
nand U2655 (N_2655,N_2578,N_2617);
nor U2656 (N_2656,N_2552,N_2615);
nor U2657 (N_2657,N_2614,N_2563);
and U2658 (N_2658,N_2609,N_2608);
nor U2659 (N_2659,N_2551,N_2556);
nor U2660 (N_2660,N_2595,N_2581);
and U2661 (N_2661,N_2619,N_2598);
nor U2662 (N_2662,N_2622,N_2550);
or U2663 (N_2663,N_2619,N_2623);
nand U2664 (N_2664,N_2577,N_2610);
and U2665 (N_2665,N_2550,N_2611);
or U2666 (N_2666,N_2564,N_2594);
or U2667 (N_2667,N_2580,N_2598);
or U2668 (N_2668,N_2597,N_2618);
and U2669 (N_2669,N_2556,N_2616);
or U2670 (N_2670,N_2590,N_2562);
or U2671 (N_2671,N_2589,N_2565);
nor U2672 (N_2672,N_2610,N_2571);
nor U2673 (N_2673,N_2580,N_2573);
nor U2674 (N_2674,N_2602,N_2586);
nand U2675 (N_2675,N_2595,N_2588);
nor U2676 (N_2676,N_2568,N_2555);
and U2677 (N_2677,N_2583,N_2574);
or U2678 (N_2678,N_2576,N_2622);
nor U2679 (N_2679,N_2587,N_2619);
nand U2680 (N_2680,N_2600,N_2603);
nor U2681 (N_2681,N_2607,N_2614);
or U2682 (N_2682,N_2558,N_2601);
or U2683 (N_2683,N_2579,N_2588);
nor U2684 (N_2684,N_2623,N_2563);
and U2685 (N_2685,N_2564,N_2608);
and U2686 (N_2686,N_2589,N_2621);
or U2687 (N_2687,N_2624,N_2606);
nor U2688 (N_2688,N_2624,N_2554);
nand U2689 (N_2689,N_2575,N_2583);
or U2690 (N_2690,N_2561,N_2566);
nor U2691 (N_2691,N_2624,N_2558);
or U2692 (N_2692,N_2572,N_2616);
or U2693 (N_2693,N_2577,N_2575);
or U2694 (N_2694,N_2603,N_2613);
or U2695 (N_2695,N_2596,N_2584);
nand U2696 (N_2696,N_2565,N_2598);
nand U2697 (N_2697,N_2565,N_2615);
nand U2698 (N_2698,N_2613,N_2576);
nor U2699 (N_2699,N_2594,N_2566);
nor U2700 (N_2700,N_2654,N_2634);
nor U2701 (N_2701,N_2667,N_2633);
nor U2702 (N_2702,N_2668,N_2647);
nand U2703 (N_2703,N_2689,N_2658);
nor U2704 (N_2704,N_2691,N_2665);
xor U2705 (N_2705,N_2662,N_2646);
nor U2706 (N_2706,N_2661,N_2684);
nand U2707 (N_2707,N_2630,N_2653);
and U2708 (N_2708,N_2695,N_2686);
nand U2709 (N_2709,N_2674,N_2688);
nand U2710 (N_2710,N_2659,N_2671);
and U2711 (N_2711,N_2676,N_2670);
and U2712 (N_2712,N_2679,N_2655);
nand U2713 (N_2713,N_2645,N_2643);
and U2714 (N_2714,N_2685,N_2664);
nor U2715 (N_2715,N_2699,N_2680);
and U2716 (N_2716,N_2637,N_2669);
or U2717 (N_2717,N_2675,N_2650);
nand U2718 (N_2718,N_2638,N_2666);
and U2719 (N_2719,N_2656,N_2636);
or U2720 (N_2720,N_2629,N_2694);
nor U2721 (N_2721,N_2628,N_2677);
and U2722 (N_2722,N_2651,N_2660);
and U2723 (N_2723,N_2683,N_2657);
nor U2724 (N_2724,N_2641,N_2698);
and U2725 (N_2725,N_2692,N_2642);
nor U2726 (N_2726,N_2673,N_2693);
or U2727 (N_2727,N_2697,N_2672);
and U2728 (N_2728,N_2648,N_2639);
nand U2729 (N_2729,N_2632,N_2652);
or U2730 (N_2730,N_2635,N_2631);
nand U2731 (N_2731,N_2626,N_2681);
and U2732 (N_2732,N_2649,N_2678);
and U2733 (N_2733,N_2627,N_2625);
and U2734 (N_2734,N_2640,N_2687);
nand U2735 (N_2735,N_2682,N_2644);
or U2736 (N_2736,N_2696,N_2690);
nor U2737 (N_2737,N_2663,N_2662);
nand U2738 (N_2738,N_2666,N_2635);
nand U2739 (N_2739,N_2666,N_2678);
nand U2740 (N_2740,N_2664,N_2667);
nand U2741 (N_2741,N_2680,N_2696);
nor U2742 (N_2742,N_2666,N_2647);
and U2743 (N_2743,N_2682,N_2645);
or U2744 (N_2744,N_2627,N_2678);
and U2745 (N_2745,N_2652,N_2639);
nand U2746 (N_2746,N_2648,N_2655);
and U2747 (N_2747,N_2658,N_2629);
or U2748 (N_2748,N_2625,N_2687);
or U2749 (N_2749,N_2636,N_2683);
and U2750 (N_2750,N_2676,N_2652);
or U2751 (N_2751,N_2688,N_2656);
nand U2752 (N_2752,N_2649,N_2691);
and U2753 (N_2753,N_2653,N_2631);
and U2754 (N_2754,N_2690,N_2640);
and U2755 (N_2755,N_2671,N_2682);
nor U2756 (N_2756,N_2676,N_2655);
and U2757 (N_2757,N_2640,N_2678);
nor U2758 (N_2758,N_2690,N_2642);
nand U2759 (N_2759,N_2683,N_2658);
nor U2760 (N_2760,N_2651,N_2696);
nand U2761 (N_2761,N_2662,N_2658);
nand U2762 (N_2762,N_2660,N_2668);
nand U2763 (N_2763,N_2687,N_2674);
nor U2764 (N_2764,N_2664,N_2686);
nand U2765 (N_2765,N_2648,N_2669);
and U2766 (N_2766,N_2657,N_2643);
and U2767 (N_2767,N_2629,N_2642);
and U2768 (N_2768,N_2684,N_2671);
or U2769 (N_2769,N_2690,N_2695);
nor U2770 (N_2770,N_2687,N_2659);
nor U2771 (N_2771,N_2638,N_2646);
xnor U2772 (N_2772,N_2662,N_2683);
and U2773 (N_2773,N_2698,N_2686);
nor U2774 (N_2774,N_2629,N_2641);
and U2775 (N_2775,N_2747,N_2712);
or U2776 (N_2776,N_2730,N_2754);
and U2777 (N_2777,N_2752,N_2715);
or U2778 (N_2778,N_2753,N_2716);
or U2779 (N_2779,N_2718,N_2773);
and U2780 (N_2780,N_2760,N_2749);
and U2781 (N_2781,N_2736,N_2726);
nor U2782 (N_2782,N_2758,N_2744);
or U2783 (N_2783,N_2717,N_2738);
nor U2784 (N_2784,N_2741,N_2766);
nand U2785 (N_2785,N_2774,N_2770);
nor U2786 (N_2786,N_2725,N_2746);
and U2787 (N_2787,N_2732,N_2723);
and U2788 (N_2788,N_2722,N_2714);
xor U2789 (N_2789,N_2710,N_2751);
nor U2790 (N_2790,N_2750,N_2740);
nor U2791 (N_2791,N_2762,N_2761);
nand U2792 (N_2792,N_2757,N_2743);
and U2793 (N_2793,N_2704,N_2734);
nand U2794 (N_2794,N_2745,N_2768);
or U2795 (N_2795,N_2756,N_2700);
nor U2796 (N_2796,N_2703,N_2764);
nand U2797 (N_2797,N_2735,N_2769);
or U2798 (N_2798,N_2706,N_2713);
nor U2799 (N_2799,N_2731,N_2772);
nor U2800 (N_2800,N_2707,N_2763);
nor U2801 (N_2801,N_2765,N_2724);
nand U2802 (N_2802,N_2767,N_2709);
nor U2803 (N_2803,N_2755,N_2727);
xor U2804 (N_2804,N_2719,N_2733);
nor U2805 (N_2805,N_2728,N_2711);
or U2806 (N_2806,N_2742,N_2729);
and U2807 (N_2807,N_2737,N_2701);
and U2808 (N_2808,N_2739,N_2705);
nor U2809 (N_2809,N_2702,N_2708);
nor U2810 (N_2810,N_2721,N_2759);
or U2811 (N_2811,N_2771,N_2748);
and U2812 (N_2812,N_2720,N_2773);
nor U2813 (N_2813,N_2754,N_2737);
nor U2814 (N_2814,N_2774,N_2748);
or U2815 (N_2815,N_2761,N_2729);
and U2816 (N_2816,N_2747,N_2763);
xor U2817 (N_2817,N_2703,N_2741);
or U2818 (N_2818,N_2722,N_2761);
or U2819 (N_2819,N_2731,N_2773);
and U2820 (N_2820,N_2772,N_2702);
and U2821 (N_2821,N_2708,N_2722);
nor U2822 (N_2822,N_2769,N_2720);
nand U2823 (N_2823,N_2761,N_2768);
or U2824 (N_2824,N_2723,N_2704);
or U2825 (N_2825,N_2705,N_2768);
nor U2826 (N_2826,N_2747,N_2760);
nand U2827 (N_2827,N_2742,N_2726);
or U2828 (N_2828,N_2732,N_2749);
nor U2829 (N_2829,N_2733,N_2706);
or U2830 (N_2830,N_2742,N_2735);
nand U2831 (N_2831,N_2736,N_2769);
and U2832 (N_2832,N_2769,N_2754);
nor U2833 (N_2833,N_2745,N_2742);
nor U2834 (N_2834,N_2773,N_2723);
nand U2835 (N_2835,N_2725,N_2754);
xor U2836 (N_2836,N_2711,N_2768);
nor U2837 (N_2837,N_2740,N_2709);
nand U2838 (N_2838,N_2751,N_2735);
or U2839 (N_2839,N_2743,N_2756);
or U2840 (N_2840,N_2748,N_2713);
nand U2841 (N_2841,N_2726,N_2711);
or U2842 (N_2842,N_2717,N_2712);
nor U2843 (N_2843,N_2721,N_2708);
nand U2844 (N_2844,N_2739,N_2759);
and U2845 (N_2845,N_2763,N_2771);
and U2846 (N_2846,N_2759,N_2770);
nor U2847 (N_2847,N_2747,N_2754);
and U2848 (N_2848,N_2724,N_2700);
or U2849 (N_2849,N_2762,N_2751);
nand U2850 (N_2850,N_2837,N_2780);
nand U2851 (N_2851,N_2797,N_2804);
nor U2852 (N_2852,N_2802,N_2819);
or U2853 (N_2853,N_2808,N_2839);
nor U2854 (N_2854,N_2836,N_2788);
or U2855 (N_2855,N_2838,N_2799);
nand U2856 (N_2856,N_2801,N_2830);
nor U2857 (N_2857,N_2825,N_2820);
nand U2858 (N_2858,N_2835,N_2823);
or U2859 (N_2859,N_2807,N_2785);
nor U2860 (N_2860,N_2822,N_2798);
nor U2861 (N_2861,N_2789,N_2817);
and U2862 (N_2862,N_2843,N_2834);
or U2863 (N_2863,N_2810,N_2813);
nand U2864 (N_2864,N_2794,N_2841);
nand U2865 (N_2865,N_2806,N_2779);
and U2866 (N_2866,N_2787,N_2827);
nand U2867 (N_2867,N_2840,N_2784);
and U2868 (N_2868,N_2792,N_2814);
nor U2869 (N_2869,N_2815,N_2781);
or U2870 (N_2870,N_2821,N_2809);
or U2871 (N_2871,N_2777,N_2782);
or U2872 (N_2872,N_2800,N_2786);
or U2873 (N_2873,N_2791,N_2849);
and U2874 (N_2874,N_2796,N_2818);
or U2875 (N_2875,N_2783,N_2842);
nand U2876 (N_2876,N_2805,N_2812);
nor U2877 (N_2877,N_2828,N_2803);
or U2878 (N_2878,N_2816,N_2847);
nand U2879 (N_2879,N_2826,N_2831);
xnor U2880 (N_2880,N_2844,N_2811);
nor U2881 (N_2881,N_2778,N_2845);
nand U2882 (N_2882,N_2824,N_2793);
nand U2883 (N_2883,N_2776,N_2795);
nand U2884 (N_2884,N_2848,N_2790);
or U2885 (N_2885,N_2833,N_2829);
nor U2886 (N_2886,N_2775,N_2846);
xor U2887 (N_2887,N_2832,N_2798);
or U2888 (N_2888,N_2791,N_2827);
and U2889 (N_2889,N_2820,N_2777);
and U2890 (N_2890,N_2817,N_2842);
and U2891 (N_2891,N_2783,N_2833);
nor U2892 (N_2892,N_2825,N_2806);
nor U2893 (N_2893,N_2805,N_2794);
nand U2894 (N_2894,N_2810,N_2816);
nand U2895 (N_2895,N_2821,N_2828);
and U2896 (N_2896,N_2800,N_2835);
or U2897 (N_2897,N_2791,N_2837);
nand U2898 (N_2898,N_2816,N_2803);
and U2899 (N_2899,N_2806,N_2831);
nand U2900 (N_2900,N_2804,N_2805);
nor U2901 (N_2901,N_2828,N_2816);
nor U2902 (N_2902,N_2845,N_2791);
or U2903 (N_2903,N_2845,N_2792);
and U2904 (N_2904,N_2807,N_2788);
nand U2905 (N_2905,N_2847,N_2821);
and U2906 (N_2906,N_2821,N_2806);
nand U2907 (N_2907,N_2808,N_2840);
nor U2908 (N_2908,N_2828,N_2830);
nand U2909 (N_2909,N_2802,N_2810);
nand U2910 (N_2910,N_2788,N_2795);
nand U2911 (N_2911,N_2828,N_2781);
or U2912 (N_2912,N_2783,N_2809);
or U2913 (N_2913,N_2835,N_2809);
and U2914 (N_2914,N_2822,N_2818);
or U2915 (N_2915,N_2810,N_2775);
or U2916 (N_2916,N_2775,N_2828);
or U2917 (N_2917,N_2812,N_2794);
nand U2918 (N_2918,N_2797,N_2840);
and U2919 (N_2919,N_2786,N_2835);
nor U2920 (N_2920,N_2807,N_2831);
nor U2921 (N_2921,N_2848,N_2803);
nor U2922 (N_2922,N_2781,N_2831);
or U2923 (N_2923,N_2834,N_2806);
nand U2924 (N_2924,N_2798,N_2825);
nand U2925 (N_2925,N_2880,N_2886);
nor U2926 (N_2926,N_2876,N_2870);
nor U2927 (N_2927,N_2919,N_2852);
and U2928 (N_2928,N_2853,N_2922);
or U2929 (N_2929,N_2865,N_2858);
nand U2930 (N_2930,N_2854,N_2860);
nor U2931 (N_2931,N_2859,N_2917);
nand U2932 (N_2932,N_2873,N_2893);
nand U2933 (N_2933,N_2881,N_2850);
nor U2934 (N_2934,N_2861,N_2921);
nand U2935 (N_2935,N_2874,N_2877);
nand U2936 (N_2936,N_2899,N_2871);
or U2937 (N_2937,N_2875,N_2896);
nor U2938 (N_2938,N_2855,N_2885);
nor U2939 (N_2939,N_2869,N_2863);
and U2940 (N_2940,N_2879,N_2912);
or U2941 (N_2941,N_2868,N_2898);
nor U2942 (N_2942,N_2914,N_2857);
nor U2943 (N_2943,N_2867,N_2909);
or U2944 (N_2944,N_2910,N_2907);
nand U2945 (N_2945,N_2906,N_2872);
nor U2946 (N_2946,N_2883,N_2892);
and U2947 (N_2947,N_2864,N_2918);
nor U2948 (N_2948,N_2866,N_2894);
nand U2949 (N_2949,N_2900,N_2913);
and U2950 (N_2950,N_2887,N_2890);
nand U2951 (N_2951,N_2862,N_2923);
nor U2952 (N_2952,N_2901,N_2905);
or U2953 (N_2953,N_2908,N_2902);
nand U2954 (N_2954,N_2911,N_2856);
nor U2955 (N_2955,N_2882,N_2851);
nand U2956 (N_2956,N_2895,N_2891);
or U2957 (N_2957,N_2878,N_2920);
nand U2958 (N_2958,N_2915,N_2904);
nor U2959 (N_2959,N_2884,N_2897);
nor U2960 (N_2960,N_2924,N_2889);
or U2961 (N_2961,N_2903,N_2888);
xnor U2962 (N_2962,N_2916,N_2882);
or U2963 (N_2963,N_2911,N_2868);
nand U2964 (N_2964,N_2872,N_2850);
nand U2965 (N_2965,N_2864,N_2858);
nand U2966 (N_2966,N_2920,N_2870);
nor U2967 (N_2967,N_2894,N_2923);
nor U2968 (N_2968,N_2916,N_2876);
nor U2969 (N_2969,N_2871,N_2874);
or U2970 (N_2970,N_2854,N_2893);
nand U2971 (N_2971,N_2905,N_2861);
or U2972 (N_2972,N_2909,N_2905);
nor U2973 (N_2973,N_2918,N_2868);
nor U2974 (N_2974,N_2850,N_2893);
nand U2975 (N_2975,N_2897,N_2852);
and U2976 (N_2976,N_2912,N_2922);
nor U2977 (N_2977,N_2883,N_2915);
or U2978 (N_2978,N_2885,N_2865);
or U2979 (N_2979,N_2869,N_2899);
or U2980 (N_2980,N_2874,N_2858);
nor U2981 (N_2981,N_2870,N_2921);
nand U2982 (N_2982,N_2906,N_2889);
nor U2983 (N_2983,N_2867,N_2863);
and U2984 (N_2984,N_2895,N_2919);
or U2985 (N_2985,N_2870,N_2913);
or U2986 (N_2986,N_2870,N_2856);
nand U2987 (N_2987,N_2882,N_2893);
or U2988 (N_2988,N_2851,N_2853);
xnor U2989 (N_2989,N_2898,N_2853);
or U2990 (N_2990,N_2882,N_2892);
nor U2991 (N_2991,N_2883,N_2918);
nor U2992 (N_2992,N_2875,N_2867);
nor U2993 (N_2993,N_2870,N_2889);
and U2994 (N_2994,N_2901,N_2880);
or U2995 (N_2995,N_2870,N_2861);
nand U2996 (N_2996,N_2892,N_2885);
or U2997 (N_2997,N_2916,N_2919);
nor U2998 (N_2998,N_2890,N_2867);
and U2999 (N_2999,N_2876,N_2924);
and UO_0 (O_0,N_2995,N_2954);
or UO_1 (O_1,N_2937,N_2976);
or UO_2 (O_2,N_2998,N_2941);
or UO_3 (O_3,N_2936,N_2970);
nor UO_4 (O_4,N_2945,N_2953);
nand UO_5 (O_5,N_2928,N_2982);
nand UO_6 (O_6,N_2971,N_2932);
nor UO_7 (O_7,N_2957,N_2997);
and UO_8 (O_8,N_2975,N_2965);
or UO_9 (O_9,N_2931,N_2947);
or UO_10 (O_10,N_2952,N_2940);
or UO_11 (O_11,N_2996,N_2993);
nand UO_12 (O_12,N_2978,N_2973);
and UO_13 (O_13,N_2938,N_2999);
and UO_14 (O_14,N_2979,N_2949);
and UO_15 (O_15,N_2935,N_2991);
or UO_16 (O_16,N_2948,N_2925);
nor UO_17 (O_17,N_2981,N_2966);
nand UO_18 (O_18,N_2967,N_2988);
or UO_19 (O_19,N_2962,N_2933);
and UO_20 (O_20,N_2939,N_2959);
and UO_21 (O_21,N_2950,N_2955);
and UO_22 (O_22,N_2934,N_2930);
and UO_23 (O_23,N_2960,N_2942);
nor UO_24 (O_24,N_2992,N_2972);
and UO_25 (O_25,N_2984,N_2944);
or UO_26 (O_26,N_2946,N_2958);
nand UO_27 (O_27,N_2987,N_2968);
and UO_28 (O_28,N_2986,N_2926);
and UO_29 (O_29,N_2974,N_2951);
nor UO_30 (O_30,N_2927,N_2977);
nor UO_31 (O_31,N_2963,N_2961);
and UO_32 (O_32,N_2980,N_2983);
and UO_33 (O_33,N_2964,N_2969);
or UO_34 (O_34,N_2929,N_2943);
or UO_35 (O_35,N_2985,N_2990);
or UO_36 (O_36,N_2956,N_2989);
nand UO_37 (O_37,N_2994,N_2952);
nor UO_38 (O_38,N_2968,N_2995);
nand UO_39 (O_39,N_2942,N_2967);
or UO_40 (O_40,N_2945,N_2955);
and UO_41 (O_41,N_2988,N_2925);
or UO_42 (O_42,N_2938,N_2976);
and UO_43 (O_43,N_2969,N_2935);
and UO_44 (O_44,N_2981,N_2965);
or UO_45 (O_45,N_2990,N_2926);
or UO_46 (O_46,N_2995,N_2994);
and UO_47 (O_47,N_2940,N_2979);
and UO_48 (O_48,N_2984,N_2951);
or UO_49 (O_49,N_2930,N_2996);
and UO_50 (O_50,N_2930,N_2942);
and UO_51 (O_51,N_2936,N_2980);
and UO_52 (O_52,N_2961,N_2925);
and UO_53 (O_53,N_2938,N_2972);
nor UO_54 (O_54,N_2971,N_2942);
and UO_55 (O_55,N_2944,N_2958);
or UO_56 (O_56,N_2977,N_2951);
nor UO_57 (O_57,N_2943,N_2948);
nor UO_58 (O_58,N_2938,N_2958);
nor UO_59 (O_59,N_2994,N_2957);
and UO_60 (O_60,N_2940,N_2965);
or UO_61 (O_61,N_2927,N_2983);
nand UO_62 (O_62,N_2994,N_2930);
xor UO_63 (O_63,N_2938,N_2980);
and UO_64 (O_64,N_2957,N_2971);
and UO_65 (O_65,N_2995,N_2958);
or UO_66 (O_66,N_2937,N_2932);
nand UO_67 (O_67,N_2971,N_2997);
nand UO_68 (O_68,N_2995,N_2961);
and UO_69 (O_69,N_2969,N_2997);
or UO_70 (O_70,N_2971,N_2984);
and UO_71 (O_71,N_2983,N_2979);
or UO_72 (O_72,N_2959,N_2927);
nand UO_73 (O_73,N_2952,N_2939);
and UO_74 (O_74,N_2936,N_2958);
nand UO_75 (O_75,N_2955,N_2982);
and UO_76 (O_76,N_2992,N_2963);
nor UO_77 (O_77,N_2937,N_2952);
and UO_78 (O_78,N_2950,N_2972);
or UO_79 (O_79,N_2930,N_2941);
nand UO_80 (O_80,N_2981,N_2991);
nor UO_81 (O_81,N_2937,N_2943);
nand UO_82 (O_82,N_2962,N_2927);
nor UO_83 (O_83,N_2987,N_2997);
and UO_84 (O_84,N_2976,N_2948);
or UO_85 (O_85,N_2951,N_2962);
nand UO_86 (O_86,N_2930,N_2985);
nor UO_87 (O_87,N_2998,N_2950);
nor UO_88 (O_88,N_2998,N_2969);
nand UO_89 (O_89,N_2957,N_2989);
nor UO_90 (O_90,N_2952,N_2990);
nor UO_91 (O_91,N_2967,N_2948);
nor UO_92 (O_92,N_2929,N_2985);
nand UO_93 (O_93,N_2972,N_2951);
or UO_94 (O_94,N_2934,N_2978);
or UO_95 (O_95,N_2987,N_2972);
nor UO_96 (O_96,N_2966,N_2931);
or UO_97 (O_97,N_2939,N_2969);
nand UO_98 (O_98,N_2972,N_2997);
nor UO_99 (O_99,N_2963,N_2942);
or UO_100 (O_100,N_2960,N_2964);
xor UO_101 (O_101,N_2989,N_2954);
or UO_102 (O_102,N_2953,N_2981);
and UO_103 (O_103,N_2972,N_2953);
or UO_104 (O_104,N_2983,N_2976);
or UO_105 (O_105,N_2977,N_2968);
nand UO_106 (O_106,N_2994,N_2998);
nor UO_107 (O_107,N_2959,N_2973);
nand UO_108 (O_108,N_2936,N_2969);
nor UO_109 (O_109,N_2927,N_2925);
nor UO_110 (O_110,N_2950,N_2953);
or UO_111 (O_111,N_2990,N_2975);
or UO_112 (O_112,N_2934,N_2981);
nor UO_113 (O_113,N_2976,N_2994);
nor UO_114 (O_114,N_2942,N_2972);
nor UO_115 (O_115,N_2991,N_2986);
or UO_116 (O_116,N_2980,N_2995);
nand UO_117 (O_117,N_2973,N_2948);
or UO_118 (O_118,N_2974,N_2966);
nand UO_119 (O_119,N_2982,N_2927);
nor UO_120 (O_120,N_2926,N_2934);
nor UO_121 (O_121,N_2963,N_2983);
nand UO_122 (O_122,N_2938,N_2929);
and UO_123 (O_123,N_2948,N_2966);
and UO_124 (O_124,N_2949,N_2946);
nor UO_125 (O_125,N_2941,N_2994);
nor UO_126 (O_126,N_2973,N_2934);
and UO_127 (O_127,N_2930,N_2938);
and UO_128 (O_128,N_2952,N_2976);
and UO_129 (O_129,N_2946,N_2964);
nand UO_130 (O_130,N_2943,N_2977);
nor UO_131 (O_131,N_2955,N_2951);
nor UO_132 (O_132,N_2950,N_2981);
nor UO_133 (O_133,N_2993,N_2987);
nor UO_134 (O_134,N_2983,N_2955);
or UO_135 (O_135,N_2933,N_2949);
or UO_136 (O_136,N_2957,N_2975);
nand UO_137 (O_137,N_2995,N_2943);
and UO_138 (O_138,N_2928,N_2926);
nor UO_139 (O_139,N_2999,N_2956);
nand UO_140 (O_140,N_2984,N_2959);
xnor UO_141 (O_141,N_2929,N_2991);
nand UO_142 (O_142,N_2985,N_2995);
nor UO_143 (O_143,N_2998,N_2943);
or UO_144 (O_144,N_2993,N_2944);
nand UO_145 (O_145,N_2989,N_2987);
or UO_146 (O_146,N_2942,N_2973);
nand UO_147 (O_147,N_2943,N_2925);
and UO_148 (O_148,N_2975,N_2930);
or UO_149 (O_149,N_2929,N_2960);
or UO_150 (O_150,N_2953,N_2991);
and UO_151 (O_151,N_2996,N_2976);
nor UO_152 (O_152,N_2960,N_2928);
or UO_153 (O_153,N_2948,N_2961);
nand UO_154 (O_154,N_2943,N_2945);
xor UO_155 (O_155,N_2934,N_2995);
nand UO_156 (O_156,N_2956,N_2929);
nand UO_157 (O_157,N_2969,N_2976);
or UO_158 (O_158,N_2983,N_2940);
nor UO_159 (O_159,N_2932,N_2955);
nor UO_160 (O_160,N_2965,N_2943);
nor UO_161 (O_161,N_2955,N_2988);
nor UO_162 (O_162,N_2991,N_2985);
and UO_163 (O_163,N_2982,N_2980);
and UO_164 (O_164,N_2932,N_2992);
nand UO_165 (O_165,N_2967,N_2993);
and UO_166 (O_166,N_2974,N_2989);
and UO_167 (O_167,N_2986,N_2925);
nand UO_168 (O_168,N_2940,N_2980);
or UO_169 (O_169,N_2985,N_2931);
and UO_170 (O_170,N_2937,N_2980);
nand UO_171 (O_171,N_2943,N_2953);
nand UO_172 (O_172,N_2957,N_2970);
and UO_173 (O_173,N_2990,N_2945);
xor UO_174 (O_174,N_2945,N_2977);
and UO_175 (O_175,N_2991,N_2965);
nand UO_176 (O_176,N_2943,N_2940);
nand UO_177 (O_177,N_2973,N_2954);
nor UO_178 (O_178,N_2999,N_2990);
or UO_179 (O_179,N_2966,N_2968);
nand UO_180 (O_180,N_2954,N_2983);
nor UO_181 (O_181,N_2973,N_2960);
or UO_182 (O_182,N_2926,N_2963);
nor UO_183 (O_183,N_2934,N_2940);
and UO_184 (O_184,N_2932,N_2961);
or UO_185 (O_185,N_2928,N_2983);
and UO_186 (O_186,N_2987,N_2959);
nor UO_187 (O_187,N_2932,N_2988);
and UO_188 (O_188,N_2982,N_2950);
or UO_189 (O_189,N_2980,N_2957);
nor UO_190 (O_190,N_2956,N_2936);
and UO_191 (O_191,N_2945,N_2927);
nor UO_192 (O_192,N_2928,N_2953);
and UO_193 (O_193,N_2930,N_2970);
and UO_194 (O_194,N_2936,N_2964);
nor UO_195 (O_195,N_2935,N_2964);
or UO_196 (O_196,N_2979,N_2938);
nand UO_197 (O_197,N_2934,N_2957);
and UO_198 (O_198,N_2946,N_2931);
and UO_199 (O_199,N_2975,N_2998);
nand UO_200 (O_200,N_2949,N_2999);
and UO_201 (O_201,N_2989,N_2962);
and UO_202 (O_202,N_2939,N_2964);
or UO_203 (O_203,N_2960,N_2949);
nor UO_204 (O_204,N_2944,N_2998);
and UO_205 (O_205,N_2967,N_2998);
or UO_206 (O_206,N_2944,N_2983);
nor UO_207 (O_207,N_2940,N_2988);
nand UO_208 (O_208,N_2934,N_2992);
nor UO_209 (O_209,N_2977,N_2925);
or UO_210 (O_210,N_2963,N_2995);
nand UO_211 (O_211,N_2933,N_2967);
and UO_212 (O_212,N_2993,N_2995);
and UO_213 (O_213,N_2959,N_2982);
nor UO_214 (O_214,N_2931,N_2936);
nand UO_215 (O_215,N_2933,N_2979);
nor UO_216 (O_216,N_2987,N_2927);
or UO_217 (O_217,N_2969,N_2931);
nor UO_218 (O_218,N_2957,N_2943);
nand UO_219 (O_219,N_2962,N_2957);
and UO_220 (O_220,N_2937,N_2939);
nand UO_221 (O_221,N_2942,N_2957);
and UO_222 (O_222,N_2962,N_2963);
nor UO_223 (O_223,N_2927,N_2967);
nand UO_224 (O_224,N_2990,N_2944);
nand UO_225 (O_225,N_2993,N_2992);
nand UO_226 (O_226,N_2983,N_2987);
nor UO_227 (O_227,N_2931,N_2945);
or UO_228 (O_228,N_2990,N_2961);
or UO_229 (O_229,N_2954,N_2999);
nand UO_230 (O_230,N_2933,N_2963);
nand UO_231 (O_231,N_2950,N_2939);
nor UO_232 (O_232,N_2980,N_2976);
xnor UO_233 (O_233,N_2995,N_2974);
nor UO_234 (O_234,N_2951,N_2986);
or UO_235 (O_235,N_2925,N_2969);
nor UO_236 (O_236,N_2990,N_2995);
and UO_237 (O_237,N_2933,N_2930);
nand UO_238 (O_238,N_2980,N_2934);
nand UO_239 (O_239,N_2973,N_2984);
nor UO_240 (O_240,N_2970,N_2934);
and UO_241 (O_241,N_2999,N_2939);
and UO_242 (O_242,N_2944,N_2934);
nor UO_243 (O_243,N_2952,N_2931);
and UO_244 (O_244,N_2956,N_2935);
nand UO_245 (O_245,N_2931,N_2972);
nor UO_246 (O_246,N_2976,N_2929);
nand UO_247 (O_247,N_2977,N_2979);
and UO_248 (O_248,N_2950,N_2967);
nor UO_249 (O_249,N_2961,N_2944);
and UO_250 (O_250,N_2954,N_2979);
nand UO_251 (O_251,N_2936,N_2987);
and UO_252 (O_252,N_2929,N_2994);
nor UO_253 (O_253,N_2938,N_2948);
nand UO_254 (O_254,N_2986,N_2930);
or UO_255 (O_255,N_2930,N_2993);
nor UO_256 (O_256,N_2958,N_2951);
or UO_257 (O_257,N_2999,N_2967);
nor UO_258 (O_258,N_2927,N_2949);
and UO_259 (O_259,N_2963,N_2959);
or UO_260 (O_260,N_2970,N_2964);
nor UO_261 (O_261,N_2952,N_2971);
and UO_262 (O_262,N_2981,N_2968);
nand UO_263 (O_263,N_2935,N_2933);
nand UO_264 (O_264,N_2928,N_2929);
nor UO_265 (O_265,N_2938,N_2988);
nand UO_266 (O_266,N_2933,N_2982);
or UO_267 (O_267,N_2932,N_2987);
and UO_268 (O_268,N_2927,N_2971);
and UO_269 (O_269,N_2971,N_2993);
nand UO_270 (O_270,N_2942,N_2978);
or UO_271 (O_271,N_2979,N_2956);
nor UO_272 (O_272,N_2931,N_2981);
or UO_273 (O_273,N_2937,N_2948);
or UO_274 (O_274,N_2971,N_2974);
nand UO_275 (O_275,N_2943,N_2951);
and UO_276 (O_276,N_2987,N_2970);
nor UO_277 (O_277,N_2927,N_2942);
nor UO_278 (O_278,N_2955,N_2963);
nor UO_279 (O_279,N_2994,N_2931);
and UO_280 (O_280,N_2945,N_2951);
nand UO_281 (O_281,N_2994,N_2965);
or UO_282 (O_282,N_2998,N_2981);
and UO_283 (O_283,N_2963,N_2953);
and UO_284 (O_284,N_2974,N_2948);
or UO_285 (O_285,N_2969,N_2999);
nor UO_286 (O_286,N_2933,N_2999);
nor UO_287 (O_287,N_2949,N_2970);
nand UO_288 (O_288,N_2944,N_2926);
nor UO_289 (O_289,N_2951,N_2969);
nand UO_290 (O_290,N_2996,N_2950);
nand UO_291 (O_291,N_2983,N_2931);
and UO_292 (O_292,N_2948,N_2952);
and UO_293 (O_293,N_2935,N_2948);
and UO_294 (O_294,N_2938,N_2942);
and UO_295 (O_295,N_2943,N_2990);
or UO_296 (O_296,N_2994,N_2991);
nand UO_297 (O_297,N_2931,N_2973);
and UO_298 (O_298,N_2974,N_2978);
and UO_299 (O_299,N_2937,N_2933);
and UO_300 (O_300,N_2927,N_2968);
nand UO_301 (O_301,N_2949,N_2926);
nor UO_302 (O_302,N_2929,N_2926);
nor UO_303 (O_303,N_2938,N_2952);
and UO_304 (O_304,N_2947,N_2940);
nand UO_305 (O_305,N_2951,N_2950);
and UO_306 (O_306,N_2958,N_2989);
nand UO_307 (O_307,N_2985,N_2934);
and UO_308 (O_308,N_2993,N_2951);
nand UO_309 (O_309,N_2951,N_2997);
and UO_310 (O_310,N_2986,N_2977);
nor UO_311 (O_311,N_2949,N_2945);
nand UO_312 (O_312,N_2999,N_2931);
or UO_313 (O_313,N_2975,N_2926);
and UO_314 (O_314,N_2968,N_2963);
nor UO_315 (O_315,N_2980,N_2951);
or UO_316 (O_316,N_2965,N_2973);
and UO_317 (O_317,N_2991,N_2988);
or UO_318 (O_318,N_2998,N_2937);
nand UO_319 (O_319,N_2946,N_2997);
nor UO_320 (O_320,N_2975,N_2925);
or UO_321 (O_321,N_2999,N_2958);
or UO_322 (O_322,N_2994,N_2962);
nor UO_323 (O_323,N_2955,N_2996);
nand UO_324 (O_324,N_2932,N_2960);
nand UO_325 (O_325,N_2980,N_2961);
nor UO_326 (O_326,N_2954,N_2946);
nor UO_327 (O_327,N_2941,N_2972);
nand UO_328 (O_328,N_2942,N_2988);
nor UO_329 (O_329,N_2974,N_2972);
nor UO_330 (O_330,N_2939,N_2991);
nand UO_331 (O_331,N_2948,N_2999);
nor UO_332 (O_332,N_2949,N_2929);
nand UO_333 (O_333,N_2936,N_2983);
nand UO_334 (O_334,N_2953,N_2929);
and UO_335 (O_335,N_2951,N_2976);
nand UO_336 (O_336,N_2945,N_2933);
nand UO_337 (O_337,N_2979,N_2957);
nand UO_338 (O_338,N_2998,N_2948);
nor UO_339 (O_339,N_2987,N_2953);
nand UO_340 (O_340,N_2963,N_2999);
and UO_341 (O_341,N_2980,N_2994);
nand UO_342 (O_342,N_2926,N_2952);
or UO_343 (O_343,N_2993,N_2975);
or UO_344 (O_344,N_2928,N_2998);
or UO_345 (O_345,N_2981,N_2945);
and UO_346 (O_346,N_2995,N_2956);
nor UO_347 (O_347,N_2967,N_2972);
nand UO_348 (O_348,N_2965,N_2948);
or UO_349 (O_349,N_2984,N_2934);
and UO_350 (O_350,N_2968,N_2979);
or UO_351 (O_351,N_2930,N_2969);
or UO_352 (O_352,N_2929,N_2952);
or UO_353 (O_353,N_2925,N_2928);
nand UO_354 (O_354,N_2936,N_2999);
or UO_355 (O_355,N_2983,N_2972);
nand UO_356 (O_356,N_2994,N_2993);
and UO_357 (O_357,N_2927,N_2939);
nor UO_358 (O_358,N_2984,N_2989);
and UO_359 (O_359,N_2928,N_2986);
and UO_360 (O_360,N_2973,N_2937);
and UO_361 (O_361,N_2998,N_2936);
and UO_362 (O_362,N_2999,N_2968);
or UO_363 (O_363,N_2983,N_2958);
and UO_364 (O_364,N_2966,N_2998);
nand UO_365 (O_365,N_2979,N_2974);
nor UO_366 (O_366,N_2941,N_2950);
and UO_367 (O_367,N_2963,N_2971);
or UO_368 (O_368,N_2981,N_2995);
or UO_369 (O_369,N_2930,N_2984);
or UO_370 (O_370,N_2957,N_2982);
nand UO_371 (O_371,N_2973,N_2933);
nand UO_372 (O_372,N_2938,N_2994);
nor UO_373 (O_373,N_2962,N_2926);
and UO_374 (O_374,N_2960,N_2978);
and UO_375 (O_375,N_2993,N_2988);
or UO_376 (O_376,N_2952,N_2944);
nand UO_377 (O_377,N_2938,N_2946);
and UO_378 (O_378,N_2985,N_2951);
nand UO_379 (O_379,N_2989,N_2946);
nor UO_380 (O_380,N_2938,N_2966);
nand UO_381 (O_381,N_2995,N_2972);
or UO_382 (O_382,N_2970,N_2933);
nor UO_383 (O_383,N_2941,N_2934);
nand UO_384 (O_384,N_2948,N_2997);
or UO_385 (O_385,N_2935,N_2988);
nor UO_386 (O_386,N_2964,N_2967);
or UO_387 (O_387,N_2938,N_2956);
xnor UO_388 (O_388,N_2949,N_2939);
or UO_389 (O_389,N_2978,N_2980);
nand UO_390 (O_390,N_2966,N_2997);
and UO_391 (O_391,N_2982,N_2965);
nand UO_392 (O_392,N_2995,N_2973);
nand UO_393 (O_393,N_2973,N_2993);
nand UO_394 (O_394,N_2978,N_2996);
or UO_395 (O_395,N_2948,N_2987);
or UO_396 (O_396,N_2945,N_2995);
nand UO_397 (O_397,N_2980,N_2925);
nor UO_398 (O_398,N_2954,N_2926);
or UO_399 (O_399,N_2931,N_2955);
nand UO_400 (O_400,N_2999,N_2950);
nor UO_401 (O_401,N_2982,N_2952);
nand UO_402 (O_402,N_2993,N_2941);
nor UO_403 (O_403,N_2930,N_2943);
nor UO_404 (O_404,N_2994,N_2932);
or UO_405 (O_405,N_2929,N_2951);
or UO_406 (O_406,N_2968,N_2973);
nand UO_407 (O_407,N_2951,N_2991);
nor UO_408 (O_408,N_2933,N_2940);
or UO_409 (O_409,N_2980,N_2952);
nand UO_410 (O_410,N_2979,N_2964);
nand UO_411 (O_411,N_2982,N_2940);
nand UO_412 (O_412,N_2945,N_2971);
or UO_413 (O_413,N_2986,N_2934);
nor UO_414 (O_414,N_2941,N_2980);
nor UO_415 (O_415,N_2977,N_2991);
and UO_416 (O_416,N_2955,N_2971);
nor UO_417 (O_417,N_2980,N_2958);
or UO_418 (O_418,N_2943,N_2971);
nor UO_419 (O_419,N_2971,N_2934);
or UO_420 (O_420,N_2973,N_2977);
nor UO_421 (O_421,N_2967,N_2965);
nand UO_422 (O_422,N_2943,N_2947);
and UO_423 (O_423,N_2948,N_2957);
and UO_424 (O_424,N_2974,N_2953);
and UO_425 (O_425,N_2967,N_2941);
or UO_426 (O_426,N_2928,N_2994);
nor UO_427 (O_427,N_2941,N_2966);
and UO_428 (O_428,N_2927,N_2935);
or UO_429 (O_429,N_2929,N_2932);
nor UO_430 (O_430,N_2990,N_2972);
nor UO_431 (O_431,N_2953,N_2937);
nand UO_432 (O_432,N_2935,N_2934);
nand UO_433 (O_433,N_2929,N_2986);
nor UO_434 (O_434,N_2975,N_2941);
nor UO_435 (O_435,N_2972,N_2981);
or UO_436 (O_436,N_2966,N_2976);
nor UO_437 (O_437,N_2941,N_2935);
or UO_438 (O_438,N_2943,N_2935);
nor UO_439 (O_439,N_2986,N_2942);
nand UO_440 (O_440,N_2939,N_2963);
and UO_441 (O_441,N_2940,N_2972);
and UO_442 (O_442,N_2984,N_2939);
nor UO_443 (O_443,N_2969,N_2971);
or UO_444 (O_444,N_2995,N_2971);
nand UO_445 (O_445,N_2952,N_2964);
nor UO_446 (O_446,N_2990,N_2994);
or UO_447 (O_447,N_2986,N_2952);
nor UO_448 (O_448,N_2976,N_2928);
and UO_449 (O_449,N_2993,N_2949);
and UO_450 (O_450,N_2961,N_2974);
nor UO_451 (O_451,N_2969,N_2948);
nor UO_452 (O_452,N_2969,N_2992);
nand UO_453 (O_453,N_2929,N_2995);
nand UO_454 (O_454,N_2972,N_2959);
nor UO_455 (O_455,N_2936,N_2955);
and UO_456 (O_456,N_2996,N_2980);
or UO_457 (O_457,N_2973,N_2963);
nand UO_458 (O_458,N_2936,N_2974);
or UO_459 (O_459,N_2946,N_2975);
or UO_460 (O_460,N_2991,N_2979);
and UO_461 (O_461,N_2942,N_2956);
nand UO_462 (O_462,N_2952,N_2954);
or UO_463 (O_463,N_2987,N_2957);
and UO_464 (O_464,N_2959,N_2940);
or UO_465 (O_465,N_2975,N_2968);
or UO_466 (O_466,N_2940,N_2974);
or UO_467 (O_467,N_2988,N_2977);
nand UO_468 (O_468,N_2976,N_2972);
nor UO_469 (O_469,N_2957,N_2932);
nand UO_470 (O_470,N_2940,N_2945);
and UO_471 (O_471,N_2966,N_2946);
nand UO_472 (O_472,N_2966,N_2964);
and UO_473 (O_473,N_2947,N_2986);
or UO_474 (O_474,N_2948,N_2928);
or UO_475 (O_475,N_2971,N_2937);
and UO_476 (O_476,N_2931,N_2932);
or UO_477 (O_477,N_2970,N_2960);
or UO_478 (O_478,N_2995,N_2947);
and UO_479 (O_479,N_2966,N_2943);
and UO_480 (O_480,N_2925,N_2991);
xnor UO_481 (O_481,N_2976,N_2958);
nor UO_482 (O_482,N_2962,N_2966);
and UO_483 (O_483,N_2979,N_2955);
nor UO_484 (O_484,N_2995,N_2949);
nor UO_485 (O_485,N_2991,N_2952);
nor UO_486 (O_486,N_2978,N_2947);
nand UO_487 (O_487,N_2930,N_2947);
or UO_488 (O_488,N_2971,N_2994);
nand UO_489 (O_489,N_2958,N_2955);
nor UO_490 (O_490,N_2934,N_2949);
nor UO_491 (O_491,N_2984,N_2942);
and UO_492 (O_492,N_2988,N_2943);
nand UO_493 (O_493,N_2987,N_2946);
nor UO_494 (O_494,N_2950,N_2959);
or UO_495 (O_495,N_2970,N_2972);
and UO_496 (O_496,N_2927,N_2929);
or UO_497 (O_497,N_2935,N_2953);
and UO_498 (O_498,N_2953,N_2982);
nand UO_499 (O_499,N_2968,N_2955);
endmodule