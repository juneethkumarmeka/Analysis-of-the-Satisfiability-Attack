module basic_1500_15000_2000_15_levels_5xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
or U0 (N_0,In_929,In_654);
nand U1 (N_1,In_111,In_1008);
and U2 (N_2,In_134,In_1085);
nor U3 (N_3,In_1057,In_81);
or U4 (N_4,In_1275,In_609);
and U5 (N_5,In_980,In_736);
or U6 (N_6,In_1016,In_535);
nor U7 (N_7,In_375,In_246);
or U8 (N_8,In_35,In_363);
or U9 (N_9,In_770,In_700);
or U10 (N_10,In_1491,In_1392);
nor U11 (N_11,In_651,In_718);
nand U12 (N_12,In_1409,In_785);
nand U13 (N_13,In_1256,In_48);
or U14 (N_14,In_1340,In_790);
and U15 (N_15,In_1031,In_553);
and U16 (N_16,In_323,In_653);
and U17 (N_17,In_892,In_1399);
and U18 (N_18,In_1395,In_478);
nor U19 (N_19,In_1377,In_703);
and U20 (N_20,In_429,In_978);
and U21 (N_21,In_300,In_1437);
nor U22 (N_22,In_831,In_1);
or U23 (N_23,In_328,In_24);
or U24 (N_24,In_905,In_251);
nand U25 (N_25,In_925,In_1483);
and U26 (N_26,In_1133,In_249);
nand U27 (N_27,In_171,In_150);
or U28 (N_28,In_602,In_1312);
xor U29 (N_29,In_567,In_356);
and U30 (N_30,In_1481,In_738);
nand U31 (N_31,In_159,In_1067);
and U32 (N_32,In_722,In_219);
nor U33 (N_33,In_1035,In_874);
xor U34 (N_34,In_118,In_489);
and U35 (N_35,In_934,In_1131);
nor U36 (N_36,In_1447,In_232);
or U37 (N_37,In_1114,In_165);
and U38 (N_38,In_841,In_1320);
nand U39 (N_39,In_1358,In_979);
xor U40 (N_40,In_256,In_1476);
nand U41 (N_41,In_792,In_997);
xor U42 (N_42,In_1170,In_1211);
and U43 (N_43,In_221,In_336);
xnor U44 (N_44,In_822,In_410);
or U45 (N_45,In_1064,In_926);
nand U46 (N_46,In_1363,In_915);
xnor U47 (N_47,In_864,In_1339);
nor U48 (N_48,In_107,In_484);
xnor U49 (N_49,In_1189,In_5);
nand U50 (N_50,In_682,In_26);
and U51 (N_51,In_1072,In_487);
nand U52 (N_52,In_1279,In_327);
nor U53 (N_53,In_786,In_475);
and U54 (N_54,In_1194,In_1243);
xor U55 (N_55,In_470,In_1391);
xor U56 (N_56,In_1285,In_56);
xor U57 (N_57,In_1019,In_228);
nand U58 (N_58,In_183,In_64);
nor U59 (N_59,In_523,In_359);
xor U60 (N_60,In_223,In_143);
nor U61 (N_61,In_1207,In_261);
and U62 (N_62,In_170,In_503);
and U63 (N_63,In_899,In_1315);
nor U64 (N_64,In_746,In_1466);
nand U65 (N_65,In_571,In_1038);
nand U66 (N_66,In_1247,In_519);
nand U67 (N_67,In_304,In_999);
or U68 (N_68,In_1368,In_1144);
and U69 (N_69,In_724,In_906);
and U70 (N_70,In_975,In_775);
nor U71 (N_71,In_1010,In_276);
nor U72 (N_72,In_1098,In_283);
xor U73 (N_73,In_393,In_1028);
xnor U74 (N_74,In_617,In_54);
xor U75 (N_75,In_868,In_1383);
or U76 (N_76,In_633,In_959);
nor U77 (N_77,In_1222,In_1390);
nand U78 (N_78,In_575,In_1278);
or U79 (N_79,In_139,In_1029);
and U80 (N_80,In_793,In_41);
or U81 (N_81,In_869,In_1193);
nand U82 (N_82,In_582,In_153);
or U83 (N_83,In_259,In_1054);
and U84 (N_84,In_883,In_275);
and U85 (N_85,In_384,In_1096);
xnor U86 (N_86,In_1322,In_546);
or U87 (N_87,In_1431,In_401);
nor U88 (N_88,In_1484,In_1337);
nand U89 (N_89,In_605,In_162);
and U90 (N_90,In_1369,In_124);
and U91 (N_91,In_1271,In_108);
nand U92 (N_92,In_993,In_187);
or U93 (N_93,In_396,In_345);
and U94 (N_94,In_1365,In_342);
nand U95 (N_95,In_1226,In_1348);
or U96 (N_96,In_268,In_757);
or U97 (N_97,In_326,In_65);
and U98 (N_98,In_302,In_483);
nand U99 (N_99,In_235,In_1152);
and U100 (N_100,In_1236,In_32);
nor U101 (N_101,In_989,In_1324);
or U102 (N_102,In_636,In_303);
nor U103 (N_103,In_1300,In_1490);
or U104 (N_104,In_1117,In_603);
or U105 (N_105,In_974,In_699);
or U106 (N_106,In_619,In_1341);
and U107 (N_107,In_74,In_202);
or U108 (N_108,In_1313,In_110);
nand U109 (N_109,In_15,In_257);
and U110 (N_110,In_1355,In_40);
or U111 (N_111,In_1349,In_1406);
and U112 (N_112,In_167,In_307);
nor U113 (N_113,In_1308,In_986);
or U114 (N_114,In_1219,In_1148);
nor U115 (N_115,In_876,In_579);
or U116 (N_116,In_474,In_463);
nand U117 (N_117,In_679,In_587);
nand U118 (N_118,In_237,In_325);
nor U119 (N_119,In_390,In_966);
nand U120 (N_120,In_253,In_1077);
nand U121 (N_121,In_1023,In_96);
or U122 (N_122,In_743,In_1232);
nand U123 (N_123,In_683,In_1066);
or U124 (N_124,In_727,In_1204);
nor U125 (N_125,In_835,In_1069);
nor U126 (N_126,In_1145,In_773);
xor U127 (N_127,In_885,In_1276);
nor U128 (N_128,In_229,In_1311);
nand U129 (N_129,In_1418,In_1494);
and U130 (N_130,In_1007,In_1060);
or U131 (N_131,In_901,In_838);
and U132 (N_132,In_897,In_719);
and U133 (N_133,In_182,In_1089);
nand U134 (N_134,In_1497,In_676);
or U135 (N_135,In_1456,In_1137);
nand U136 (N_136,In_729,In_1327);
or U137 (N_137,In_627,In_665);
and U138 (N_138,In_155,In_115);
nand U139 (N_139,In_294,In_84);
nand U140 (N_140,In_1142,In_753);
nand U141 (N_141,In_560,In_371);
and U142 (N_142,In_1469,In_873);
nor U143 (N_143,In_642,In_392);
or U144 (N_144,In_1055,In_531);
and U145 (N_145,In_502,In_563);
or U146 (N_146,In_127,In_696);
xnor U147 (N_147,In_333,In_961);
and U148 (N_148,In_825,In_1161);
or U149 (N_149,In_1331,In_70);
and U150 (N_150,In_339,In_1020);
nor U151 (N_151,In_1353,In_511);
or U152 (N_152,In_1043,In_1479);
and U153 (N_153,In_570,In_595);
and U154 (N_154,In_528,In_426);
nor U155 (N_155,In_1199,In_953);
or U156 (N_156,In_1128,In_947);
nor U157 (N_157,In_626,In_123);
nor U158 (N_158,In_1171,In_1006);
or U159 (N_159,In_151,In_52);
and U160 (N_160,In_550,In_128);
and U161 (N_161,In_852,In_49);
and U162 (N_162,In_774,In_436);
and U163 (N_163,In_1159,In_1467);
nor U164 (N_164,In_674,In_880);
nor U165 (N_165,In_1013,In_1021);
and U166 (N_166,In_1173,In_260);
nor U167 (N_167,In_591,In_341);
nand U168 (N_168,In_44,In_1046);
nor U169 (N_169,In_1407,In_197);
xnor U170 (N_170,In_208,In_840);
and U171 (N_171,In_416,In_849);
and U172 (N_172,In_577,In_981);
nor U173 (N_173,In_344,In_378);
or U174 (N_174,In_542,In_1345);
nand U175 (N_175,In_1295,In_1472);
and U176 (N_176,In_1178,In_1328);
nand U177 (N_177,In_4,In_1231);
nand U178 (N_178,In_1239,In_494);
nand U179 (N_179,In_547,In_1041);
nand U180 (N_180,In_62,In_17);
and U181 (N_181,In_661,In_1044);
xnor U182 (N_182,In_920,In_188);
nor U183 (N_183,In_317,In_413);
and U184 (N_184,In_488,In_1492);
or U185 (N_185,In_1319,In_781);
and U186 (N_186,In_1306,In_269);
or U187 (N_187,In_1323,In_606);
xor U188 (N_188,In_1124,In_362);
nand U189 (N_189,In_1011,In_763);
xnor U190 (N_190,In_551,In_610);
and U191 (N_191,In_860,In_723);
or U192 (N_192,In_505,In_1286);
nor U193 (N_193,In_666,In_1493);
nor U194 (N_194,In_506,In_1386);
and U195 (N_195,In_239,In_879);
nor U196 (N_196,In_71,In_100);
or U197 (N_197,In_1335,In_675);
nor U198 (N_198,In_367,In_102);
and U199 (N_199,In_122,In_1183);
and U200 (N_200,In_278,In_114);
and U201 (N_201,In_106,In_184);
nor U202 (N_202,In_600,In_126);
or U203 (N_203,In_1334,In_286);
nand U204 (N_204,In_258,In_225);
nand U205 (N_205,In_690,In_1411);
and U206 (N_206,In_417,In_1326);
nand U207 (N_207,In_2,In_98);
and U208 (N_208,In_6,In_1423);
nor U209 (N_209,In_263,In_408);
xnor U210 (N_210,In_660,In_1445);
nand U211 (N_211,In_645,In_942);
nand U212 (N_212,In_705,In_43);
or U213 (N_213,In_465,In_923);
xor U214 (N_214,In_1428,In_394);
and U215 (N_215,In_1366,In_209);
nand U216 (N_216,In_1362,In_376);
or U217 (N_217,In_1037,In_1420);
nor U218 (N_218,In_662,In_1158);
nand U219 (N_219,In_433,In_308);
and U220 (N_220,In_148,In_827);
or U221 (N_221,In_1113,In_632);
nand U222 (N_222,In_60,In_569);
or U223 (N_223,In_224,In_819);
xnor U224 (N_224,In_295,In_1346);
nor U225 (N_225,In_101,In_1487);
or U226 (N_226,In_388,In_136);
and U227 (N_227,In_596,In_316);
and U228 (N_228,In_614,In_764);
xnor U229 (N_229,In_78,In_1053);
nor U230 (N_230,In_669,In_844);
or U231 (N_231,In_836,In_28);
and U232 (N_232,In_1138,In_889);
and U233 (N_233,In_808,In_1242);
nand U234 (N_234,In_843,In_190);
nor U235 (N_235,In_214,In_8);
xnor U236 (N_236,In_497,In_1174);
and U237 (N_237,In_572,In_900);
or U238 (N_238,In_990,In_717);
and U239 (N_239,In_266,In_320);
xnor U240 (N_240,In_444,In_14);
nor U241 (N_241,In_409,In_552);
and U242 (N_242,In_33,In_291);
nor U243 (N_243,In_1121,In_305);
xor U244 (N_244,In_391,In_647);
nand U245 (N_245,In_1419,In_315);
nand U246 (N_246,In_721,In_783);
xor U247 (N_247,In_370,In_1241);
xor U248 (N_248,In_807,In_1426);
nor U249 (N_249,In_1301,In_298);
xnor U250 (N_250,In_161,In_967);
nor U251 (N_251,In_1238,In_805);
nor U252 (N_252,In_462,In_772);
nor U253 (N_253,In_29,In_1156);
or U254 (N_254,In_881,In_1022);
or U255 (N_255,In_1024,In_374);
xnor U256 (N_256,In_66,In_105);
nor U257 (N_257,In_46,In_1000);
and U258 (N_258,In_347,In_1208);
nor U259 (N_259,In_586,In_1187);
nand U260 (N_260,In_539,In_911);
or U261 (N_261,In_765,In_580);
nor U262 (N_262,In_103,In_1403);
xnor U263 (N_263,In_313,In_1485);
nand U264 (N_264,In_79,In_812);
xor U265 (N_265,In_1080,In_1436);
or U266 (N_266,In_476,In_787);
nor U267 (N_267,In_958,In_1297);
or U268 (N_268,In_544,In_839);
nand U269 (N_269,In_527,In_594);
or U270 (N_270,In_467,In_557);
nand U271 (N_271,In_893,In_789);
or U272 (N_272,In_69,In_638);
or U273 (N_273,In_310,In_18);
or U274 (N_274,In_890,In_1318);
xor U275 (N_275,In_309,In_1017);
nor U276 (N_276,In_1482,In_1457);
nor U277 (N_277,In_499,In_1270);
or U278 (N_278,In_941,In_658);
or U279 (N_279,In_1062,In_67);
and U280 (N_280,In_760,In_1294);
or U281 (N_281,In_189,In_762);
or U282 (N_282,In_725,In_833);
or U283 (N_283,In_361,In_566);
xnor U284 (N_284,In_279,In_121);
xor U285 (N_285,In_1203,In_450);
and U286 (N_286,In_1387,In_973);
and U287 (N_287,In_1224,In_985);
or U288 (N_288,In_3,In_493);
or U289 (N_289,In_425,In_1450);
xor U290 (N_290,In_210,In_1052);
xor U291 (N_291,In_262,In_241);
nor U292 (N_292,In_704,In_1047);
nor U293 (N_293,In_916,In_92);
and U294 (N_294,In_332,In_460);
and U295 (N_295,In_293,In_1273);
and U296 (N_296,In_1460,In_55);
and U297 (N_297,In_1277,In_1255);
and U298 (N_298,In_533,In_962);
or U299 (N_299,In_1237,In_185);
nand U300 (N_300,In_576,In_368);
nand U301 (N_301,In_346,In_1040);
nand U302 (N_302,In_829,In_203);
nor U303 (N_303,In_635,In_630);
or U304 (N_304,In_383,In_1120);
nor U305 (N_305,In_853,In_1119);
and U306 (N_306,In_1112,In_971);
nor U307 (N_307,In_377,In_797);
or U308 (N_308,In_856,In_991);
or U309 (N_309,In_521,In_61);
nor U310 (N_310,In_1215,In_265);
or U311 (N_311,In_846,In_1015);
xnor U312 (N_312,In_1050,In_956);
and U313 (N_313,In_697,In_1453);
xor U314 (N_314,In_299,In_943);
and U315 (N_315,In_855,In_629);
or U316 (N_316,In_198,In_117);
nor U317 (N_317,In_671,In_1109);
xor U318 (N_318,In_357,In_23);
and U319 (N_319,In_1150,In_922);
xnor U320 (N_320,In_640,In_284);
nand U321 (N_321,In_73,In_964);
and U322 (N_322,In_1027,In_581);
and U323 (N_323,In_1176,In_1091);
and U324 (N_324,In_621,In_1107);
nor U325 (N_325,In_1087,In_1293);
or U326 (N_326,In_1065,In_945);
or U327 (N_327,In_933,In_1032);
or U328 (N_328,In_340,In_1108);
and U329 (N_329,In_398,In_1162);
nand U330 (N_330,In_1234,In_862);
xor U331 (N_331,In_684,In_434);
nand U332 (N_332,In_495,In_976);
and U333 (N_333,In_354,In_886);
nor U334 (N_334,In_432,In_716);
nand U335 (N_335,In_407,In_1051);
or U336 (N_336,In_420,In_1364);
or U337 (N_337,In_1225,In_749);
or U338 (N_338,In_1260,In_1220);
nor U339 (N_339,In_94,In_334);
nor U340 (N_340,In_509,In_932);
or U341 (N_341,In_1036,In_1459);
or U342 (N_342,In_623,In_1134);
nor U343 (N_343,In_1001,In_1136);
or U344 (N_344,In_548,In_1444);
and U345 (N_345,In_747,In_404);
nand U346 (N_346,In_1004,In_292);
and U347 (N_347,In_1042,In_1287);
and U348 (N_348,In_1415,In_1100);
nand U349 (N_349,In_77,In_711);
or U350 (N_350,In_794,In_702);
or U351 (N_351,In_944,In_954);
and U352 (N_352,In_1421,In_1382);
or U353 (N_353,In_125,In_248);
or U354 (N_354,In_1425,In_447);
xnor U355 (N_355,In_1321,In_937);
nand U356 (N_356,In_1026,In_498);
nor U357 (N_357,In_778,In_211);
nand U358 (N_358,In_1201,In_828);
nand U359 (N_359,In_1367,In_227);
nand U360 (N_360,In_146,In_842);
and U361 (N_361,In_803,In_352);
nor U362 (N_362,In_353,In_694);
nor U363 (N_363,In_11,In_965);
or U364 (N_364,In_86,In_813);
and U365 (N_365,In_443,In_281);
nor U366 (N_366,In_192,In_598);
and U367 (N_367,In_31,In_656);
or U368 (N_368,In_592,In_996);
and U369 (N_369,In_501,In_1179);
and U370 (N_370,In_250,In_1443);
and U371 (N_371,In_1265,In_688);
or U372 (N_372,In_744,In_1446);
or U373 (N_373,In_510,In_1081);
or U374 (N_374,In_205,In_983);
nand U375 (N_375,In_806,In_903);
nand U376 (N_376,In_421,In_1427);
nand U377 (N_377,In_321,In_400);
nor U378 (N_378,In_649,In_1342);
nor U379 (N_379,In_754,In_273);
and U380 (N_380,In_1251,In_1116);
or U381 (N_381,In_565,In_1442);
and U382 (N_382,In_244,In_464);
nor U383 (N_383,In_863,In_597);
nand U384 (N_384,In_1169,In_750);
and U385 (N_385,In_365,In_473);
nor U386 (N_386,In_708,In_274);
or U387 (N_387,In_648,In_1477);
and U388 (N_388,In_245,In_379);
nand U389 (N_389,In_424,In_720);
or U390 (N_390,In_924,In_1303);
or U391 (N_391,In_496,In_1099);
nand U392 (N_392,In_1048,In_364);
nand U393 (N_393,In_512,In_952);
xor U394 (N_394,In_848,In_1402);
xor U395 (N_395,In_1106,In_1408);
nand U396 (N_396,In_604,In_1218);
or U397 (N_397,In_518,In_908);
xor U398 (N_398,In_1325,In_691);
and U399 (N_399,In_532,In_1304);
nand U400 (N_400,In_455,In_492);
and U401 (N_401,In_1448,In_1249);
and U402 (N_402,In_1405,In_1317);
nand U403 (N_403,In_1292,In_1097);
or U404 (N_404,In_714,In_319);
or U405 (N_405,In_1400,In_935);
nand U406 (N_406,In_360,In_685);
nand U407 (N_407,In_1094,In_769);
nor U408 (N_408,In_1186,In_1282);
xor U409 (N_409,In_1473,In_130);
nand U410 (N_410,In_1433,In_524);
and U411 (N_411,In_1059,In_677);
or U412 (N_412,In_173,In_540);
nor U413 (N_413,In_1248,In_854);
or U414 (N_414,In_977,In_948);
nor U415 (N_415,In_385,In_1200);
nand U416 (N_416,In_1118,In_620);
nand U417 (N_417,In_220,In_734);
or U418 (N_418,In_441,In_608);
and U419 (N_419,In_1244,In_695);
or U420 (N_420,In_157,In_1149);
or U421 (N_421,In_145,In_1141);
xnor U422 (N_422,In_1309,In_453);
or U423 (N_423,In_1375,In_1123);
xor U424 (N_424,In_931,In_427);
nor U425 (N_425,In_402,In_199);
xnor U426 (N_426,In_82,In_625);
nor U427 (N_427,In_38,In_859);
xor U428 (N_428,In_928,In_1263);
nor U429 (N_429,In_514,In_1458);
or U430 (N_430,In_850,In_1185);
nor U431 (N_431,In_80,In_439);
xor U432 (N_432,In_449,In_927);
and U433 (N_433,In_779,In_280);
nor U434 (N_434,In_1468,In_1196);
or U435 (N_435,In_381,In_89);
or U436 (N_436,In_814,In_1155);
or U437 (N_437,In_1360,In_1361);
and U438 (N_438,In_709,In_607);
nand U439 (N_439,In_713,In_201);
and U440 (N_440,In_919,In_784);
nand U441 (N_441,In_272,In_585);
or U442 (N_442,In_1350,In_1165);
xnor U443 (N_443,In_1122,In_120);
nand U444 (N_444,In_1267,In_1259);
nand U445 (N_445,In_438,In_1478);
xnor U446 (N_446,In_176,In_50);
nor U447 (N_447,In_1359,In_1430);
xor U448 (N_448,In_1465,In_593);
nor U449 (N_449,In_804,In_504);
nand U450 (N_450,In_826,In_914);
and U451 (N_451,In_1463,In_147);
nor U452 (N_452,In_1274,In_373);
or U453 (N_453,In_57,In_884);
nand U454 (N_454,In_1240,In_196);
and U455 (N_455,In_329,In_918);
and U456 (N_456,In_1254,In_599);
or U457 (N_457,In_45,In_1132);
xnor U458 (N_458,In_1332,In_243);
nand U459 (N_459,In_1167,In_556);
nand U460 (N_460,In_1412,In_659);
or U461 (N_461,In_53,In_950);
and U462 (N_462,In_692,In_330);
or U463 (N_463,In_878,In_418);
nand U464 (N_464,In_680,In_289);
nand U465 (N_465,In_739,In_1164);
nand U466 (N_466,In_758,In_264);
nand U467 (N_467,In_1221,In_358);
and U468 (N_468,In_1129,In_380);
nand U469 (N_469,In_578,In_898);
and U470 (N_470,In_657,In_12);
and U471 (N_471,In_1143,In_963);
nand U472 (N_472,In_76,In_1389);
and U473 (N_473,In_1115,In_1197);
and U474 (N_474,In_1033,In_1449);
nand U475 (N_475,In_16,In_681);
and U476 (N_476,In_795,In_780);
and U477 (N_477,In_1495,In_821);
and U478 (N_478,In_1045,In_534);
nand U479 (N_479,In_761,In_1058);
xnor U480 (N_480,In_175,In_1356);
and U481 (N_481,In_397,In_768);
nor U482 (N_482,In_451,In_1281);
or U483 (N_483,In_1451,In_777);
and U484 (N_484,In_917,In_133);
and U485 (N_485,In_177,In_1250);
xnor U486 (N_486,In_1212,In_255);
and U487 (N_487,In_655,In_1296);
or U488 (N_488,In_1370,In_1330);
xnor U489 (N_489,In_1432,In_431);
or U490 (N_490,In_445,In_242);
nand U491 (N_491,In_851,In_297);
nor U492 (N_492,In_1252,In_174);
xnor U493 (N_493,In_456,In_998);
or U494 (N_494,In_141,In_1351);
xnor U495 (N_495,In_559,In_58);
nor U496 (N_496,In_1381,In_1498);
and U497 (N_497,In_446,In_222);
nor U498 (N_498,In_930,In_1268);
nand U499 (N_499,In_154,In_109);
nor U500 (N_500,In_386,In_351);
or U501 (N_501,In_584,In_231);
nor U502 (N_502,In_1126,In_1086);
xnor U503 (N_503,In_472,In_179);
and U504 (N_504,In_1266,In_399);
nor U505 (N_505,In_664,In_796);
or U506 (N_506,In_686,In_522);
xnor U507 (N_507,In_382,In_1075);
and U508 (N_508,In_887,In_296);
nand U509 (N_509,In_865,In_1214);
and U510 (N_510,In_1307,In_454);
and U511 (N_511,In_1217,In_1262);
nor U512 (N_512,In_672,In_631);
or U513 (N_513,In_628,In_1352);
nor U514 (N_514,In_545,In_217);
xnor U515 (N_515,In_1455,In_491);
and U516 (N_516,In_1003,In_1229);
or U517 (N_517,In_290,In_663);
nor U518 (N_518,In_168,In_767);
nand U519 (N_519,In_1233,In_195);
nand U520 (N_520,In_1235,In_37);
and U521 (N_521,In_1347,In_830);
or U522 (N_522,In_322,In_834);
or U523 (N_523,In_1338,In_311);
nand U524 (N_524,In_907,In_1213);
nand U525 (N_525,In_1230,In_156);
nand U526 (N_526,In_13,In_233);
nor U527 (N_527,In_1147,In_47);
and U528 (N_528,In_508,In_1486);
xnor U529 (N_529,In_987,In_215);
xnor U530 (N_530,In_562,In_68);
or U531 (N_531,In_637,In_163);
nor U532 (N_532,In_823,In_728);
nand U533 (N_533,In_1191,In_537);
and U534 (N_534,In_1014,In_1088);
nor U535 (N_535,In_1401,In_1374);
or U536 (N_536,In_1413,In_588);
nand U537 (N_537,In_240,In_1439);
or U538 (N_538,In_613,In_536);
nor U539 (N_539,In_1452,In_87);
or U540 (N_540,In_1475,In_1385);
xnor U541 (N_541,In_1499,In_1394);
nor U542 (N_542,In_1216,In_318);
nor U543 (N_543,In_1210,In_1462);
nor U544 (N_544,In_164,In_1461);
nor U545 (N_545,In_1049,In_216);
nor U546 (N_546,In_751,In_403);
nand U547 (N_547,In_938,In_1269);
or U548 (N_548,In_574,In_1298);
nor U549 (N_549,In_896,In_618);
and U550 (N_550,In_1206,In_554);
nor U551 (N_551,In_1329,In_138);
nor U552 (N_552,In_583,In_555);
xnor U553 (N_553,In_940,In_90);
nand U554 (N_554,In_815,In_1095);
and U555 (N_555,In_969,In_701);
xor U556 (N_556,In_448,In_589);
nand U557 (N_557,In_1034,In_1414);
nor U558 (N_558,In_1025,In_1344);
and U559 (N_559,In_1410,In_191);
nand U560 (N_560,In_91,In_324);
and U561 (N_561,In_1333,In_1074);
xnor U562 (N_562,In_477,In_1076);
nand U563 (N_563,In_1154,In_1079);
or U564 (N_564,In_1223,In_689);
nor U565 (N_565,In_788,In_238);
or U566 (N_566,In_207,In_206);
or U567 (N_567,In_471,In_355);
or U568 (N_568,In_1068,In_817);
and U569 (N_569,In_9,In_212);
or U570 (N_570,In_1272,In_271);
or U571 (N_571,In_564,In_678);
or U572 (N_572,In_314,In_461);
nor U573 (N_573,In_481,In_135);
and U574 (N_574,In_1157,In_25);
and U575 (N_575,In_349,In_939);
and U576 (N_576,In_234,In_372);
or U577 (N_577,In_1188,In_1093);
nor U578 (N_578,In_236,In_1082);
or U579 (N_579,In_1258,In_1435);
nand U580 (N_580,In_913,In_1184);
nand U581 (N_581,In_673,In_837);
xor U582 (N_582,In_706,In_1177);
nor U583 (N_583,In_1102,In_1464);
nor U584 (N_584,In_1388,In_1125);
and U585 (N_585,In_1496,In_142);
or U586 (N_586,In_343,In_1371);
nand U587 (N_587,In_858,In_1380);
or U588 (N_588,In_646,In_1316);
or U589 (N_589,In_158,In_160);
and U590 (N_590,In_538,In_348);
nor U591 (N_591,In_34,In_411);
xnor U592 (N_592,In_301,In_615);
xor U593 (N_593,In_909,In_1130);
or U594 (N_594,In_1398,In_759);
or U595 (N_595,In_1302,In_641);
nor U596 (N_596,In_816,In_818);
nor U597 (N_597,In_992,In_1198);
or U598 (N_598,In_847,In_288);
nand U599 (N_599,In_1018,In_549);
nor U600 (N_600,In_824,In_1283);
or U601 (N_601,In_652,In_104);
nand U602 (N_602,In_1146,In_366);
xnor U603 (N_603,In_1379,In_995);
or U604 (N_604,In_1291,In_1314);
nand U605 (N_605,In_1376,In_137);
nor U606 (N_606,In_482,In_1253);
xnor U607 (N_607,In_337,In_912);
nand U608 (N_608,In_590,In_601);
nor U609 (N_609,In_218,In_277);
nand U610 (N_610,In_960,In_1105);
and U611 (N_611,In_1002,In_335);
or U612 (N_612,In_832,In_1488);
and U613 (N_613,In_479,In_1429);
nor U614 (N_614,In_984,In_895);
xor U615 (N_615,In_857,In_1299);
xor U616 (N_616,In_710,In_1227);
nor U617 (N_617,In_415,In_186);
nor U618 (N_618,In_1378,In_369);
nand U619 (N_619,In_132,In_644);
nand U620 (N_620,In_1151,In_1310);
nand U621 (N_621,In_766,In_1202);
nand U622 (N_622,In_752,In_193);
nor U623 (N_623,In_800,In_811);
nand U624 (N_624,In_1396,In_1092);
nand U625 (N_625,In_1063,In_515);
xor U626 (N_626,In_740,In_994);
nand U627 (N_627,In_63,In_643);
or U628 (N_628,In_1290,In_1441);
and U629 (N_629,In_507,In_1160);
and U630 (N_630,In_1440,In_802);
and U631 (N_631,In_181,In_526);
and U632 (N_632,In_480,In_810);
nand U633 (N_633,In_1139,In_875);
nor U634 (N_634,In_338,In_946);
or U635 (N_635,In_513,In_1101);
nor U636 (N_636,In_1195,In_458);
nor U637 (N_637,In_1163,In_882);
or U638 (N_638,In_1245,In_745);
or U639 (N_639,In_1454,In_712);
nor U640 (N_640,In_698,In_748);
or U641 (N_641,In_140,In_1357);
and U642 (N_642,In_1373,In_22);
nor U643 (N_643,In_891,In_85);
nand U644 (N_644,In_442,In_1417);
nand U645 (N_645,In_1209,In_204);
or U646 (N_646,In_1180,In_19);
and U647 (N_647,In_972,In_670);
or U648 (N_648,In_350,In_194);
and U649 (N_649,In_968,In_693);
and U650 (N_650,In_1422,In_129);
nor U651 (N_651,In_634,In_1261);
or U652 (N_652,In_1336,In_1061);
nor U653 (N_653,In_957,In_490);
nand U654 (N_654,In_872,In_247);
nor U655 (N_655,In_866,In_1289);
and U656 (N_656,In_541,In_112);
nand U657 (N_657,In_611,In_430);
and U658 (N_658,In_7,In_622);
nor U659 (N_659,In_955,In_782);
nand U660 (N_660,In_1005,In_93);
or U661 (N_661,In_72,In_1111);
or U662 (N_662,In_707,In_200);
nand U663 (N_663,In_525,In_715);
and U664 (N_664,In_668,In_1175);
and U665 (N_665,In_39,In_667);
nand U666 (N_666,In_520,In_867);
and U667 (N_667,In_452,In_406);
or U668 (N_668,In_732,In_1480);
or U669 (N_669,In_285,In_131);
nand U670 (N_670,In_500,In_1424);
and U671 (N_671,In_116,In_733);
or U672 (N_672,In_419,In_97);
nor U673 (N_673,In_1190,In_771);
xor U674 (N_674,In_1153,In_113);
nor U675 (N_675,In_1257,In_801);
nand U676 (N_676,In_755,In_558);
nor U677 (N_677,In_904,In_42);
xnor U678 (N_678,In_0,In_144);
or U679 (N_679,In_312,In_820);
and U680 (N_680,In_423,In_1438);
and U681 (N_681,In_970,In_1397);
and U682 (N_682,In_51,In_1246);
or U683 (N_683,In_756,In_422);
and U684 (N_684,In_435,In_639);
nor U685 (N_685,In_27,In_516);
and U686 (N_686,In_226,In_888);
and U687 (N_687,In_1354,In_988);
nand U688 (N_688,In_1078,In_1181);
nand U689 (N_689,In_1084,In_21);
nand U690 (N_690,In_1470,In_798);
and U691 (N_691,In_440,In_252);
and U692 (N_692,In_119,In_405);
or U693 (N_693,In_1030,In_1393);
nor U694 (N_694,In_1056,In_99);
nand U695 (N_695,In_861,In_270);
and U696 (N_696,In_650,In_169);
nor U697 (N_697,In_517,In_1182);
or U698 (N_698,In_742,In_149);
or U699 (N_699,In_75,In_1104);
or U700 (N_700,In_871,In_414);
nor U701 (N_701,In_735,In_230);
nand U702 (N_702,In_877,In_331);
and U703 (N_703,In_1343,In_1012);
or U704 (N_704,In_1009,In_459);
nand U705 (N_705,In_287,In_1039);
or U706 (N_706,In_1384,In_59);
nor U707 (N_707,In_1434,In_1280);
nor U708 (N_708,In_1090,In_1071);
nand U709 (N_709,In_1471,In_529);
nand U710 (N_710,In_902,In_951);
or U711 (N_711,In_1110,In_166);
nor U712 (N_712,In_1168,In_178);
nor U713 (N_713,In_1192,In_457);
or U714 (N_714,In_83,In_1103);
xor U715 (N_715,In_36,In_1135);
and U716 (N_716,In_845,In_1205);
nand U717 (N_717,In_870,In_1404);
and U718 (N_718,In_731,In_387);
or U719 (N_719,In_624,In_776);
or U720 (N_720,In_389,In_1127);
or U721 (N_721,In_791,In_737);
xnor U722 (N_722,In_10,In_530);
and U723 (N_723,In_428,In_468);
or U724 (N_724,In_1140,In_687);
nor U725 (N_725,In_936,In_485);
nand U726 (N_726,In_486,In_1284);
nor U727 (N_727,In_306,In_561);
nand U728 (N_728,In_95,In_1083);
and U729 (N_729,In_395,In_730);
nand U730 (N_730,In_152,In_1288);
or U731 (N_731,In_1073,In_30);
or U732 (N_732,In_543,In_180);
or U733 (N_733,In_1172,In_1474);
nand U734 (N_734,In_1070,In_254);
or U735 (N_735,In_921,In_894);
nor U736 (N_736,In_809,In_573);
and U737 (N_737,In_469,In_172);
xnor U738 (N_738,In_799,In_1372);
xor U739 (N_739,In_612,In_1166);
or U740 (N_740,In_20,In_437);
nand U741 (N_741,In_267,In_88);
or U742 (N_742,In_726,In_949);
nand U743 (N_743,In_568,In_1264);
nor U744 (N_744,In_282,In_1489);
or U745 (N_745,In_982,In_1305);
nor U746 (N_746,In_1228,In_616);
and U747 (N_747,In_466,In_213);
nand U748 (N_748,In_1416,In_741);
nor U749 (N_749,In_412,In_910);
and U750 (N_750,In_1162,In_80);
xnor U751 (N_751,In_1271,In_35);
nand U752 (N_752,In_304,In_429);
and U753 (N_753,In_601,In_1250);
or U754 (N_754,In_42,In_509);
or U755 (N_755,In_69,In_1423);
or U756 (N_756,In_1431,In_312);
and U757 (N_757,In_719,In_1103);
and U758 (N_758,In_1124,In_96);
nor U759 (N_759,In_258,In_1483);
or U760 (N_760,In_358,In_563);
or U761 (N_761,In_452,In_1009);
nor U762 (N_762,In_1309,In_1323);
xor U763 (N_763,In_66,In_1413);
xor U764 (N_764,In_924,In_450);
nand U765 (N_765,In_440,In_235);
and U766 (N_766,In_1149,In_443);
or U767 (N_767,In_805,In_1201);
nor U768 (N_768,In_550,In_476);
or U769 (N_769,In_1108,In_640);
nand U770 (N_770,In_1213,In_165);
nand U771 (N_771,In_434,In_516);
or U772 (N_772,In_1424,In_1259);
or U773 (N_773,In_151,In_1262);
and U774 (N_774,In_525,In_610);
or U775 (N_775,In_611,In_76);
nand U776 (N_776,In_1386,In_929);
or U777 (N_777,In_376,In_1370);
nor U778 (N_778,In_1064,In_1287);
xnor U779 (N_779,In_586,In_897);
or U780 (N_780,In_424,In_451);
nand U781 (N_781,In_946,In_1002);
nor U782 (N_782,In_286,In_1185);
or U783 (N_783,In_1260,In_923);
or U784 (N_784,In_97,In_23);
nor U785 (N_785,In_943,In_930);
nor U786 (N_786,In_269,In_125);
nand U787 (N_787,In_75,In_1174);
xnor U788 (N_788,In_650,In_658);
nor U789 (N_789,In_722,In_553);
nand U790 (N_790,In_975,In_721);
or U791 (N_791,In_923,In_1288);
nor U792 (N_792,In_1193,In_1126);
nand U793 (N_793,In_1200,In_170);
or U794 (N_794,In_1132,In_88);
nor U795 (N_795,In_387,In_97);
xor U796 (N_796,In_92,In_1336);
nor U797 (N_797,In_964,In_767);
or U798 (N_798,In_107,In_1438);
nor U799 (N_799,In_984,In_947);
and U800 (N_800,In_192,In_930);
xnor U801 (N_801,In_163,In_79);
nor U802 (N_802,In_19,In_127);
or U803 (N_803,In_557,In_510);
or U804 (N_804,In_1220,In_1349);
or U805 (N_805,In_433,In_469);
nand U806 (N_806,In_193,In_399);
or U807 (N_807,In_1125,In_768);
or U808 (N_808,In_504,In_1047);
nand U809 (N_809,In_559,In_1060);
or U810 (N_810,In_1063,In_880);
and U811 (N_811,In_920,In_675);
and U812 (N_812,In_125,In_468);
nor U813 (N_813,In_819,In_133);
or U814 (N_814,In_1216,In_193);
nand U815 (N_815,In_329,In_117);
or U816 (N_816,In_450,In_1328);
nand U817 (N_817,In_263,In_20);
or U818 (N_818,In_1344,In_1246);
nor U819 (N_819,In_1404,In_711);
or U820 (N_820,In_697,In_241);
or U821 (N_821,In_22,In_758);
or U822 (N_822,In_1200,In_1015);
nand U823 (N_823,In_1338,In_514);
nand U824 (N_824,In_1445,In_1356);
nor U825 (N_825,In_1147,In_974);
or U826 (N_826,In_1445,In_126);
nand U827 (N_827,In_110,In_1440);
and U828 (N_828,In_664,In_1002);
nor U829 (N_829,In_288,In_376);
nor U830 (N_830,In_1438,In_822);
nor U831 (N_831,In_263,In_25);
xnor U832 (N_832,In_332,In_1121);
and U833 (N_833,In_283,In_1258);
nand U834 (N_834,In_166,In_852);
or U835 (N_835,In_560,In_981);
and U836 (N_836,In_614,In_1018);
nand U837 (N_837,In_635,In_874);
or U838 (N_838,In_826,In_1398);
nor U839 (N_839,In_1125,In_1187);
nor U840 (N_840,In_477,In_936);
or U841 (N_841,In_1116,In_1121);
and U842 (N_842,In_625,In_1204);
or U843 (N_843,In_1018,In_794);
nor U844 (N_844,In_1174,In_615);
nand U845 (N_845,In_1386,In_738);
xnor U846 (N_846,In_458,In_1351);
and U847 (N_847,In_1274,In_361);
and U848 (N_848,In_644,In_841);
and U849 (N_849,In_1254,In_335);
xnor U850 (N_850,In_124,In_1238);
nand U851 (N_851,In_1316,In_698);
xor U852 (N_852,In_33,In_512);
and U853 (N_853,In_593,In_1452);
xor U854 (N_854,In_1386,In_288);
nor U855 (N_855,In_718,In_470);
or U856 (N_856,In_1441,In_964);
nor U857 (N_857,In_834,In_960);
or U858 (N_858,In_505,In_1228);
nand U859 (N_859,In_830,In_941);
and U860 (N_860,In_651,In_931);
nand U861 (N_861,In_430,In_851);
or U862 (N_862,In_450,In_1205);
nor U863 (N_863,In_946,In_1151);
and U864 (N_864,In_353,In_808);
nand U865 (N_865,In_498,In_1341);
nor U866 (N_866,In_1426,In_657);
nand U867 (N_867,In_1081,In_1229);
nor U868 (N_868,In_218,In_968);
or U869 (N_869,In_864,In_265);
and U870 (N_870,In_1128,In_1390);
nand U871 (N_871,In_138,In_1337);
and U872 (N_872,In_1329,In_1244);
and U873 (N_873,In_729,In_384);
nor U874 (N_874,In_1354,In_937);
and U875 (N_875,In_1300,In_964);
and U876 (N_876,In_1023,In_83);
xor U877 (N_877,In_1470,In_477);
nand U878 (N_878,In_1252,In_556);
nor U879 (N_879,In_355,In_840);
nand U880 (N_880,In_403,In_420);
nand U881 (N_881,In_726,In_912);
and U882 (N_882,In_996,In_1070);
nor U883 (N_883,In_212,In_556);
nor U884 (N_884,In_845,In_1368);
nor U885 (N_885,In_462,In_658);
and U886 (N_886,In_1482,In_694);
nor U887 (N_887,In_253,In_858);
or U888 (N_888,In_0,In_641);
or U889 (N_889,In_941,In_1092);
or U890 (N_890,In_632,In_703);
nor U891 (N_891,In_1393,In_241);
xor U892 (N_892,In_1488,In_750);
or U893 (N_893,In_761,In_925);
or U894 (N_894,In_319,In_229);
and U895 (N_895,In_677,In_360);
nor U896 (N_896,In_1023,In_1229);
nor U897 (N_897,In_1116,In_1174);
or U898 (N_898,In_1129,In_41);
nor U899 (N_899,In_1055,In_1010);
or U900 (N_900,In_384,In_800);
nor U901 (N_901,In_1150,In_210);
xor U902 (N_902,In_1342,In_778);
nor U903 (N_903,In_1275,In_838);
or U904 (N_904,In_648,In_324);
nand U905 (N_905,In_1133,In_666);
nand U906 (N_906,In_14,In_1384);
nand U907 (N_907,In_638,In_959);
or U908 (N_908,In_962,In_52);
or U909 (N_909,In_880,In_107);
nand U910 (N_910,In_230,In_915);
nor U911 (N_911,In_789,In_945);
nand U912 (N_912,In_1454,In_388);
nand U913 (N_913,In_1125,In_616);
xnor U914 (N_914,In_1341,In_790);
or U915 (N_915,In_1452,In_581);
xnor U916 (N_916,In_246,In_619);
and U917 (N_917,In_744,In_604);
nor U918 (N_918,In_1087,In_761);
nor U919 (N_919,In_1210,In_147);
or U920 (N_920,In_268,In_682);
xor U921 (N_921,In_1165,In_163);
and U922 (N_922,In_170,In_237);
nor U923 (N_923,In_193,In_1466);
nand U924 (N_924,In_171,In_1231);
or U925 (N_925,In_1291,In_932);
and U926 (N_926,In_1136,In_659);
nor U927 (N_927,In_123,In_1358);
and U928 (N_928,In_1050,In_1367);
and U929 (N_929,In_992,In_269);
and U930 (N_930,In_705,In_840);
or U931 (N_931,In_1376,In_505);
nand U932 (N_932,In_357,In_590);
and U933 (N_933,In_441,In_296);
or U934 (N_934,In_698,In_1072);
or U935 (N_935,In_1264,In_315);
nand U936 (N_936,In_441,In_716);
and U937 (N_937,In_1025,In_1305);
or U938 (N_938,In_72,In_1498);
nor U939 (N_939,In_996,In_398);
nor U940 (N_940,In_52,In_1053);
nand U941 (N_941,In_256,In_668);
nand U942 (N_942,In_338,In_187);
xor U943 (N_943,In_115,In_1445);
and U944 (N_944,In_332,In_826);
or U945 (N_945,In_155,In_1417);
nor U946 (N_946,In_1243,In_552);
and U947 (N_947,In_1358,In_120);
nor U948 (N_948,In_366,In_1443);
and U949 (N_949,In_749,In_970);
xor U950 (N_950,In_640,In_1144);
and U951 (N_951,In_1473,In_309);
nand U952 (N_952,In_931,In_1138);
xor U953 (N_953,In_1163,In_1045);
nand U954 (N_954,In_738,In_1048);
nand U955 (N_955,In_952,In_637);
nor U956 (N_956,In_1116,In_703);
and U957 (N_957,In_942,In_41);
and U958 (N_958,In_1455,In_1234);
or U959 (N_959,In_226,In_150);
nor U960 (N_960,In_517,In_273);
nand U961 (N_961,In_612,In_467);
xor U962 (N_962,In_918,In_1033);
nor U963 (N_963,In_1049,In_721);
or U964 (N_964,In_828,In_1475);
or U965 (N_965,In_1176,In_199);
xor U966 (N_966,In_1233,In_1004);
nor U967 (N_967,In_518,In_1223);
and U968 (N_968,In_1286,In_401);
xor U969 (N_969,In_157,In_214);
nand U970 (N_970,In_118,In_312);
and U971 (N_971,In_390,In_1327);
and U972 (N_972,In_676,In_1172);
or U973 (N_973,In_1469,In_1075);
nor U974 (N_974,In_729,In_114);
nor U975 (N_975,In_1110,In_422);
xnor U976 (N_976,In_146,In_1132);
nor U977 (N_977,In_960,In_1267);
nor U978 (N_978,In_1044,In_526);
nor U979 (N_979,In_552,In_283);
xnor U980 (N_980,In_1207,In_1306);
nor U981 (N_981,In_348,In_1077);
nor U982 (N_982,In_976,In_394);
or U983 (N_983,In_584,In_893);
nand U984 (N_984,In_653,In_657);
xnor U985 (N_985,In_517,In_332);
and U986 (N_986,In_472,In_1425);
nor U987 (N_987,In_948,In_955);
and U988 (N_988,In_703,In_1357);
or U989 (N_989,In_80,In_1035);
and U990 (N_990,In_925,In_1295);
and U991 (N_991,In_573,In_1100);
or U992 (N_992,In_1253,In_1453);
nand U993 (N_993,In_461,In_726);
xor U994 (N_994,In_723,In_184);
xor U995 (N_995,In_335,In_509);
nand U996 (N_996,In_867,In_671);
xor U997 (N_997,In_617,In_235);
and U998 (N_998,In_439,In_557);
and U999 (N_999,In_106,In_689);
or U1000 (N_1000,N_807,N_904);
or U1001 (N_1001,N_269,N_975);
or U1002 (N_1002,N_552,N_474);
and U1003 (N_1003,N_72,N_683);
or U1004 (N_1004,N_422,N_828);
or U1005 (N_1005,N_594,N_829);
nor U1006 (N_1006,N_387,N_735);
nand U1007 (N_1007,N_968,N_528);
or U1008 (N_1008,N_251,N_709);
nor U1009 (N_1009,N_942,N_383);
and U1010 (N_1010,N_515,N_997);
or U1011 (N_1011,N_164,N_281);
or U1012 (N_1012,N_498,N_682);
xnor U1013 (N_1013,N_410,N_283);
and U1014 (N_1014,N_108,N_938);
xor U1015 (N_1015,N_761,N_712);
nor U1016 (N_1016,N_230,N_687);
nand U1017 (N_1017,N_122,N_192);
nor U1018 (N_1018,N_670,N_597);
and U1019 (N_1019,N_977,N_535);
nor U1020 (N_1020,N_981,N_789);
nor U1021 (N_1021,N_943,N_423);
or U1022 (N_1022,N_16,N_660);
and U1023 (N_1023,N_179,N_431);
and U1024 (N_1024,N_638,N_45);
or U1025 (N_1025,N_113,N_727);
nand U1026 (N_1026,N_900,N_915);
nand U1027 (N_1027,N_188,N_126);
or U1028 (N_1028,N_489,N_249);
nand U1029 (N_1029,N_110,N_842);
nand U1030 (N_1030,N_825,N_152);
nand U1031 (N_1031,N_551,N_123);
nor U1032 (N_1032,N_166,N_394);
nor U1033 (N_1033,N_362,N_624);
and U1034 (N_1034,N_823,N_395);
nand U1035 (N_1035,N_637,N_458);
nand U1036 (N_1036,N_701,N_169);
nor U1037 (N_1037,N_949,N_689);
and U1038 (N_1038,N_416,N_768);
nand U1039 (N_1039,N_506,N_534);
nor U1040 (N_1040,N_974,N_71);
or U1041 (N_1041,N_128,N_565);
and U1042 (N_1042,N_725,N_457);
nand U1043 (N_1043,N_103,N_722);
nand U1044 (N_1044,N_559,N_767);
and U1045 (N_1045,N_634,N_56);
xor U1046 (N_1046,N_325,N_928);
nand U1047 (N_1047,N_958,N_412);
or U1048 (N_1048,N_878,N_293);
or U1049 (N_1049,N_414,N_479);
nand U1050 (N_1050,N_966,N_496);
nor U1051 (N_1051,N_11,N_539);
and U1052 (N_1052,N_445,N_577);
nand U1053 (N_1053,N_906,N_77);
xnor U1054 (N_1054,N_935,N_702);
or U1055 (N_1055,N_610,N_830);
nand U1056 (N_1056,N_619,N_833);
nor U1057 (N_1057,N_875,N_891);
nand U1058 (N_1058,N_208,N_766);
nand U1059 (N_1059,N_247,N_973);
and U1060 (N_1060,N_4,N_163);
nand U1061 (N_1061,N_76,N_724);
nand U1062 (N_1062,N_596,N_23);
nand U1063 (N_1063,N_932,N_644);
and U1064 (N_1064,N_363,N_581);
or U1065 (N_1065,N_65,N_522);
nand U1066 (N_1066,N_814,N_694);
and U1067 (N_1067,N_959,N_476);
nand U1068 (N_1068,N_526,N_0);
and U1069 (N_1069,N_843,N_693);
and U1070 (N_1070,N_918,N_354);
or U1071 (N_1071,N_599,N_125);
and U1072 (N_1072,N_576,N_824);
or U1073 (N_1073,N_1,N_503);
nand U1074 (N_1074,N_834,N_554);
and U1075 (N_1075,N_628,N_510);
or U1076 (N_1076,N_73,N_36);
nor U1077 (N_1077,N_386,N_282);
nand U1078 (N_1078,N_519,N_51);
nor U1079 (N_1079,N_266,N_730);
nor U1080 (N_1080,N_334,N_140);
nor U1081 (N_1081,N_157,N_224);
nor U1082 (N_1082,N_186,N_81);
nor U1083 (N_1083,N_517,N_780);
or U1084 (N_1084,N_7,N_490);
or U1085 (N_1085,N_323,N_390);
nor U1086 (N_1086,N_415,N_425);
or U1087 (N_1087,N_35,N_172);
and U1088 (N_1088,N_237,N_575);
or U1089 (N_1089,N_792,N_37);
and U1090 (N_1090,N_254,N_305);
and U1091 (N_1091,N_376,N_561);
nor U1092 (N_1092,N_233,N_289);
nor U1093 (N_1093,N_819,N_226);
nor U1094 (N_1094,N_105,N_89);
xnor U1095 (N_1095,N_483,N_221);
nor U1096 (N_1096,N_146,N_527);
nand U1097 (N_1097,N_868,N_936);
or U1098 (N_1098,N_132,N_661);
nand U1099 (N_1099,N_967,N_826);
nand U1100 (N_1100,N_751,N_54);
nand U1101 (N_1101,N_46,N_207);
nand U1102 (N_1102,N_288,N_436);
nor U1103 (N_1103,N_742,N_889);
nor U1104 (N_1104,N_240,N_782);
nand U1105 (N_1105,N_337,N_351);
and U1106 (N_1106,N_846,N_516);
nor U1107 (N_1107,N_839,N_700);
nand U1108 (N_1108,N_443,N_264);
nand U1109 (N_1109,N_741,N_899);
nand U1110 (N_1110,N_631,N_642);
nand U1111 (N_1111,N_950,N_450);
nand U1112 (N_1112,N_406,N_646);
nor U1113 (N_1113,N_931,N_570);
and U1114 (N_1114,N_276,N_707);
or U1115 (N_1115,N_12,N_990);
and U1116 (N_1116,N_107,N_513);
or U1117 (N_1117,N_389,N_74);
or U1118 (N_1118,N_769,N_69);
or U1119 (N_1119,N_862,N_428);
or U1120 (N_1120,N_524,N_442);
nand U1121 (N_1121,N_426,N_630);
nand U1122 (N_1122,N_691,N_111);
nand U1123 (N_1123,N_781,N_505);
xor U1124 (N_1124,N_259,N_796);
nand U1125 (N_1125,N_137,N_220);
nor U1126 (N_1126,N_130,N_155);
nand U1127 (N_1127,N_40,N_794);
and U1128 (N_1128,N_468,N_292);
nand U1129 (N_1129,N_316,N_518);
nand U1130 (N_1130,N_972,N_867);
and U1131 (N_1131,N_655,N_598);
nor U1132 (N_1132,N_866,N_507);
and U1133 (N_1133,N_898,N_752);
nor U1134 (N_1134,N_589,N_718);
nor U1135 (N_1135,N_896,N_665);
or U1136 (N_1136,N_326,N_333);
and U1137 (N_1137,N_229,N_222);
and U1138 (N_1138,N_921,N_234);
and U1139 (N_1139,N_705,N_461);
and U1140 (N_1140,N_708,N_307);
and U1141 (N_1141,N_897,N_438);
nand U1142 (N_1142,N_135,N_338);
nor U1143 (N_1143,N_421,N_800);
nand U1144 (N_1144,N_852,N_262);
and U1145 (N_1145,N_348,N_61);
nand U1146 (N_1146,N_783,N_948);
or U1147 (N_1147,N_719,N_165);
nand U1148 (N_1148,N_378,N_855);
nand U1149 (N_1149,N_710,N_717);
or U1150 (N_1150,N_15,N_44);
or U1151 (N_1151,N_19,N_198);
nand U1152 (N_1152,N_941,N_9);
and U1153 (N_1153,N_388,N_758);
nor U1154 (N_1154,N_699,N_564);
nor U1155 (N_1155,N_881,N_555);
and U1156 (N_1156,N_568,N_494);
or U1157 (N_1157,N_245,N_303);
or U1158 (N_1158,N_466,N_80);
or U1159 (N_1159,N_678,N_347);
or U1160 (N_1160,N_360,N_189);
nor U1161 (N_1161,N_121,N_753);
nand U1162 (N_1162,N_716,N_558);
and U1163 (N_1163,N_120,N_971);
and U1164 (N_1164,N_956,N_593);
xor U1165 (N_1165,N_178,N_314);
or U1166 (N_1166,N_432,N_676);
and U1167 (N_1167,N_41,N_225);
xor U1168 (N_1168,N_848,N_744);
nand U1169 (N_1169,N_817,N_999);
nand U1170 (N_1170,N_812,N_860);
nor U1171 (N_1171,N_877,N_25);
nor U1172 (N_1172,N_374,N_215);
or U1173 (N_1173,N_210,N_560);
nand U1174 (N_1174,N_185,N_777);
nor U1175 (N_1175,N_181,N_879);
and U1176 (N_1176,N_850,N_984);
or U1177 (N_1177,N_925,N_601);
nand U1178 (N_1178,N_695,N_979);
nor U1179 (N_1179,N_297,N_42);
nand U1180 (N_1180,N_930,N_441);
and U1181 (N_1181,N_754,N_641);
nor U1182 (N_1182,N_223,N_652);
and U1183 (N_1183,N_549,N_116);
nor U1184 (N_1184,N_190,N_690);
and U1185 (N_1185,N_119,N_521);
nor U1186 (N_1186,N_344,N_501);
nor U1187 (N_1187,N_547,N_703);
nor U1188 (N_1188,N_33,N_329);
or U1189 (N_1189,N_308,N_34);
or U1190 (N_1190,N_924,N_893);
xor U1191 (N_1191,N_985,N_550);
nand U1192 (N_1192,N_562,N_541);
and U1193 (N_1193,N_32,N_439);
nor U1194 (N_1194,N_579,N_615);
nor U1195 (N_1195,N_733,N_58);
nor U1196 (N_1196,N_202,N_158);
nand U1197 (N_1197,N_890,N_171);
and U1198 (N_1198,N_109,N_926);
nor U1199 (N_1199,N_377,N_454);
or U1200 (N_1200,N_726,N_317);
nor U1201 (N_1201,N_847,N_255);
nand U1202 (N_1202,N_148,N_804);
or U1203 (N_1203,N_684,N_173);
and U1204 (N_1204,N_774,N_745);
nor U1205 (N_1205,N_131,N_573);
xnor U1206 (N_1206,N_728,N_865);
nand U1207 (N_1207,N_732,N_480);
and U1208 (N_1208,N_658,N_982);
or U1209 (N_1209,N_844,N_304);
or U1210 (N_1210,N_393,N_238);
nor U1211 (N_1211,N_47,N_664);
nor U1212 (N_1212,N_470,N_153);
and U1213 (N_1213,N_291,N_557);
or U1214 (N_1214,N_248,N_219);
nand U1215 (N_1215,N_986,N_82);
or U1216 (N_1216,N_149,N_663);
xor U1217 (N_1217,N_681,N_231);
nor U1218 (N_1218,N_402,N_244);
or U1219 (N_1219,N_270,N_413);
or U1220 (N_1220,N_488,N_75);
or U1221 (N_1221,N_349,N_493);
nand U1222 (N_1222,N_908,N_500);
nand U1223 (N_1223,N_688,N_662);
and U1224 (N_1224,N_391,N_204);
nand U1225 (N_1225,N_22,N_335);
or U1226 (N_1226,N_159,N_711);
xnor U1227 (N_1227,N_647,N_757);
nand U1228 (N_1228,N_242,N_706);
and U1229 (N_1229,N_680,N_100);
nand U1230 (N_1230,N_160,N_584);
and U1231 (N_1231,N_913,N_617);
nor U1232 (N_1232,N_21,N_95);
nand U1233 (N_1233,N_407,N_648);
xnor U1234 (N_1234,N_820,N_63);
nand U1235 (N_1235,N_427,N_668);
and U1236 (N_1236,N_548,N_485);
or U1237 (N_1237,N_639,N_57);
nor U1238 (N_1238,N_187,N_998);
xnor U1239 (N_1239,N_626,N_531);
and U1240 (N_1240,N_912,N_39);
and U1241 (N_1241,N_671,N_749);
nand U1242 (N_1242,N_858,N_937);
and U1243 (N_1243,N_704,N_371);
nand U1244 (N_1244,N_154,N_467);
and U1245 (N_1245,N_404,N_837);
and U1246 (N_1246,N_478,N_98);
and U1247 (N_1247,N_271,N_606);
nand U1248 (N_1248,N_49,N_306);
and U1249 (N_1249,N_286,N_954);
and U1250 (N_1250,N_434,N_471);
and U1251 (N_1251,N_696,N_243);
and U1252 (N_1252,N_94,N_26);
nand U1253 (N_1253,N_88,N_365);
or U1254 (N_1254,N_300,N_995);
nor U1255 (N_1255,N_731,N_327);
nor U1256 (N_1256,N_805,N_978);
and U1257 (N_1257,N_760,N_13);
and U1258 (N_1258,N_600,N_87);
or U1259 (N_1259,N_755,N_603);
and U1260 (N_1260,N_545,N_616);
nand U1261 (N_1261,N_235,N_359);
xor U1262 (N_1262,N_330,N_78);
or U1263 (N_1263,N_880,N_299);
and U1264 (N_1264,N_836,N_813);
nand U1265 (N_1265,N_963,N_232);
or U1266 (N_1266,N_28,N_318);
nand U1267 (N_1267,N_411,N_136);
and U1268 (N_1268,N_272,N_70);
nor U1269 (N_1269,N_882,N_373);
and U1270 (N_1270,N_141,N_544);
nand U1271 (N_1271,N_290,N_964);
or U1272 (N_1272,N_955,N_418);
or U1273 (N_1273,N_66,N_993);
nor U1274 (N_1274,N_633,N_713);
nand U1275 (N_1275,N_151,N_295);
or U1276 (N_1276,N_885,N_275);
or U1277 (N_1277,N_563,N_83);
nor U1278 (N_1278,N_933,N_692);
and U1279 (N_1279,N_460,N_771);
nand U1280 (N_1280,N_408,N_571);
xor U1281 (N_1281,N_736,N_864);
or U1282 (N_1282,N_375,N_6);
nand U1283 (N_1283,N_784,N_167);
nor U1284 (N_1284,N_324,N_538);
xnor U1285 (N_1285,N_93,N_162);
nand U1286 (N_1286,N_84,N_504);
and U1287 (N_1287,N_260,N_980);
nand U1288 (N_1288,N_572,N_267);
and U1289 (N_1289,N_20,N_320);
nor U1290 (N_1290,N_632,N_352);
nor U1291 (N_1291,N_650,N_779);
and U1292 (N_1292,N_346,N_640);
and U1293 (N_1293,N_734,N_910);
nor U1294 (N_1294,N_473,N_795);
nand U1295 (N_1295,N_118,N_969);
nor U1296 (N_1296,N_588,N_205);
xnor U1297 (N_1297,N_43,N_86);
or U1298 (N_1298,N_482,N_622);
or U1299 (N_1299,N_144,N_685);
or U1300 (N_1300,N_48,N_509);
nor U1301 (N_1301,N_659,N_604);
nand U1302 (N_1302,N_623,N_367);
and U1303 (N_1303,N_673,N_499);
and U1304 (N_1304,N_380,N_145);
nand U1305 (N_1305,N_602,N_298);
nor U1306 (N_1306,N_675,N_284);
nand U1307 (N_1307,N_355,N_112);
nand U1308 (N_1308,N_366,N_495);
nor U1309 (N_1309,N_793,N_952);
nor U1310 (N_1310,N_369,N_991);
and U1311 (N_1311,N_729,N_31);
and U1312 (N_1312,N_553,N_677);
nor U1313 (N_1313,N_651,N_193);
nor U1314 (N_1314,N_236,N_854);
nand U1315 (N_1315,N_339,N_902);
nand U1316 (N_1316,N_486,N_472);
or U1317 (N_1317,N_127,N_184);
nand U1318 (N_1318,N_511,N_951);
nor U1319 (N_1319,N_29,N_775);
nor U1320 (N_1320,N_133,N_294);
or U1321 (N_1321,N_627,N_456);
and U1322 (N_1322,N_961,N_279);
or U1323 (N_1323,N_940,N_916);
nor U1324 (N_1324,N_200,N_419);
xor U1325 (N_1325,N_96,N_216);
and U1326 (N_1326,N_191,N_392);
or U1327 (N_1327,N_310,N_117);
nand U1328 (N_1328,N_401,N_872);
and U1329 (N_1329,N_252,N_525);
and U1330 (N_1330,N_183,N_372);
or U1331 (N_1331,N_399,N_529);
or U1332 (N_1332,N_947,N_649);
xor U1333 (N_1333,N_840,N_253);
and U1334 (N_1334,N_497,N_321);
xnor U1335 (N_1335,N_962,N_440);
xnor U1336 (N_1336,N_201,N_876);
nor U1337 (N_1337,N_91,N_429);
or U1338 (N_1338,N_625,N_430);
or U1339 (N_1339,N_405,N_124);
and U1340 (N_1340,N_927,N_802);
nand U1341 (N_1341,N_832,N_853);
nand U1342 (N_1342,N_206,N_492);
nand U1343 (N_1343,N_543,N_988);
nor U1344 (N_1344,N_566,N_608);
nor U1345 (N_1345,N_356,N_987);
nor U1346 (N_1346,N_798,N_739);
or U1347 (N_1347,N_241,N_134);
and U1348 (N_1348,N_512,N_869);
or U1349 (N_1349,N_945,N_811);
or U1350 (N_1350,N_772,N_328);
and U1351 (N_1351,N_398,N_556);
and U1352 (N_1352,N_720,N_520);
and U1353 (N_1353,N_53,N_309);
nor U1354 (N_1354,N_475,N_542);
nor U1355 (N_1355,N_740,N_332);
nand U1356 (N_1356,N_546,N_274);
nand U1357 (N_1357,N_340,N_801);
and U1358 (N_1358,N_342,N_643);
nor U1359 (N_1359,N_285,N_523);
nand U1360 (N_1360,N_992,N_368);
nor U1361 (N_1361,N_838,N_976);
or U1362 (N_1362,N_903,N_487);
nand U1363 (N_1363,N_433,N_629);
nand U1364 (N_1364,N_815,N_382);
xnor U1365 (N_1365,N_67,N_656);
xor U1366 (N_1366,N_278,N_821);
and U1367 (N_1367,N_64,N_883);
or U1368 (N_1368,N_370,N_591);
nand U1369 (N_1369,N_960,N_62);
nor U1370 (N_1370,N_384,N_756);
or U1371 (N_1371,N_217,N_806);
nor U1372 (N_1372,N_763,N_5);
xnor U1373 (N_1373,N_669,N_447);
nor U1374 (N_1374,N_586,N_861);
nor U1375 (N_1375,N_462,N_147);
and U1376 (N_1376,N_199,N_743);
xor U1377 (N_1377,N_453,N_533);
and U1378 (N_1378,N_55,N_409);
xnor U1379 (N_1379,N_239,N_312);
and U1380 (N_1380,N_379,N_831);
nor U1381 (N_1381,N_827,N_27);
nor U1382 (N_1382,N_79,N_311);
nor U1383 (N_1383,N_686,N_613);
and U1384 (N_1384,N_180,N_750);
or U1385 (N_1385,N_585,N_764);
and U1386 (N_1386,N_574,N_358);
or U1387 (N_1387,N_901,N_50);
xor U1388 (N_1388,N_14,N_150);
nand U1389 (N_1389,N_922,N_18);
nor U1390 (N_1390,N_203,N_451);
and U1391 (N_1391,N_540,N_770);
or U1392 (N_1392,N_477,N_788);
and U1393 (N_1393,N_965,N_569);
nor U1394 (N_1394,N_52,N_30);
nor U1395 (N_1395,N_983,N_621);
or U1396 (N_1396,N_331,N_674);
nand U1397 (N_1397,N_592,N_580);
nor U1398 (N_1398,N_177,N_914);
and U1399 (N_1399,N_213,N_273);
and U1400 (N_1400,N_653,N_851);
nor U1401 (N_1401,N_946,N_381);
nor U1402 (N_1402,N_636,N_277);
and U1403 (N_1403,N_578,N_759);
and U1404 (N_1404,N_666,N_114);
and U1405 (N_1405,N_449,N_892);
and U1406 (N_1406,N_609,N_280);
or U1407 (N_1407,N_38,N_502);
nand U1408 (N_1408,N_212,N_747);
or U1409 (N_1409,N_508,N_92);
or U1410 (N_1410,N_104,N_8);
nor U1411 (N_1411,N_994,N_481);
xor U1412 (N_1412,N_870,N_156);
nand U1413 (N_1413,N_818,N_532);
or U1414 (N_1414,N_197,N_444);
and U1415 (N_1415,N_59,N_841);
xor U1416 (N_1416,N_341,N_888);
nor U1417 (N_1417,N_265,N_361);
or U1418 (N_1418,N_799,N_929);
nor U1419 (N_1419,N_920,N_459);
xnor U1420 (N_1420,N_797,N_364);
or U1421 (N_1421,N_301,N_143);
nand U1422 (N_1422,N_99,N_618);
nor U1423 (N_1423,N_776,N_970);
or U1424 (N_1424,N_424,N_808);
and U1425 (N_1425,N_196,N_263);
or U1426 (N_1426,N_863,N_791);
nor U1427 (N_1427,N_170,N_385);
xnor U1428 (N_1428,N_620,N_345);
nor U1429 (N_1429,N_778,N_287);
and U1430 (N_1430,N_464,N_455);
xnor U1431 (N_1431,N_895,N_679);
nor U1432 (N_1432,N_773,N_319);
nand U1433 (N_1433,N_996,N_17);
nor U1434 (N_1434,N_583,N_667);
or U1435 (N_1435,N_463,N_874);
and U1436 (N_1436,N_336,N_715);
nor U1437 (N_1437,N_437,N_810);
or U1438 (N_1438,N_400,N_917);
nand U1439 (N_1439,N_420,N_721);
nand U1440 (N_1440,N_296,N_115);
xor U1441 (N_1441,N_484,N_194);
and U1442 (N_1442,N_491,N_85);
xor U1443 (N_1443,N_258,N_138);
and U1444 (N_1444,N_469,N_397);
or U1445 (N_1445,N_919,N_612);
or U1446 (N_1446,N_857,N_887);
or U1447 (N_1447,N_214,N_582);
nand U1448 (N_1448,N_905,N_60);
or U1449 (N_1449,N_909,N_849);
nand U1450 (N_1450,N_246,N_698);
or U1451 (N_1451,N_765,N_989);
nor U1452 (N_1452,N_446,N_322);
nor U1453 (N_1453,N_261,N_873);
nor U1454 (N_1454,N_785,N_822);
xor U1455 (N_1455,N_257,N_738);
nor U1456 (N_1456,N_809,N_106);
nand U1457 (N_1457,N_657,N_786);
or U1458 (N_1458,N_803,N_886);
and U1459 (N_1459,N_465,N_714);
or U1460 (N_1460,N_907,N_587);
and U1461 (N_1461,N_923,N_605);
or U1462 (N_1462,N_313,N_939);
nor U1463 (N_1463,N_934,N_343);
and U1464 (N_1464,N_218,N_530);
xor U1465 (N_1465,N_845,N_3);
or U1466 (N_1466,N_452,N_102);
and U1467 (N_1467,N_353,N_567);
or U1468 (N_1468,N_168,N_590);
or U1469 (N_1469,N_403,N_315);
or U1470 (N_1470,N_856,N_10);
and U1471 (N_1471,N_607,N_209);
xnor U1472 (N_1472,N_97,N_835);
nor U1473 (N_1473,N_174,N_211);
nand U1474 (N_1474,N_536,N_250);
xnor U1475 (N_1475,N_357,N_175);
nor U1476 (N_1476,N_195,N_762);
xor U1477 (N_1477,N_816,N_161);
or U1478 (N_1478,N_654,N_256);
nor U1479 (N_1479,N_884,N_957);
and U1480 (N_1480,N_101,N_90);
and U1481 (N_1481,N_448,N_614);
or U1482 (N_1482,N_514,N_672);
nor U1483 (N_1483,N_68,N_176);
nor U1484 (N_1484,N_228,N_350);
and U1485 (N_1485,N_227,N_645);
and U1486 (N_1486,N_182,N_911);
and U1487 (N_1487,N_944,N_746);
nand U1488 (N_1488,N_129,N_723);
or U1489 (N_1489,N_894,N_302);
or U1490 (N_1490,N_748,N_417);
or U1491 (N_1491,N_790,N_871);
nor U1492 (N_1492,N_635,N_787);
nor U1493 (N_1493,N_142,N_268);
nand U1494 (N_1494,N_859,N_396);
or U1495 (N_1495,N_953,N_537);
nand U1496 (N_1496,N_611,N_737);
or U1497 (N_1497,N_435,N_2);
xnor U1498 (N_1498,N_697,N_139);
or U1499 (N_1499,N_24,N_595);
nor U1500 (N_1500,N_354,N_369);
nor U1501 (N_1501,N_265,N_952);
nand U1502 (N_1502,N_271,N_22);
or U1503 (N_1503,N_461,N_328);
nor U1504 (N_1504,N_772,N_543);
and U1505 (N_1505,N_332,N_922);
nor U1506 (N_1506,N_812,N_691);
or U1507 (N_1507,N_855,N_594);
or U1508 (N_1508,N_100,N_669);
or U1509 (N_1509,N_675,N_968);
nor U1510 (N_1510,N_675,N_517);
or U1511 (N_1511,N_309,N_692);
nand U1512 (N_1512,N_562,N_54);
nand U1513 (N_1513,N_467,N_996);
and U1514 (N_1514,N_956,N_467);
or U1515 (N_1515,N_829,N_578);
or U1516 (N_1516,N_709,N_410);
and U1517 (N_1517,N_383,N_680);
or U1518 (N_1518,N_444,N_482);
xnor U1519 (N_1519,N_374,N_137);
and U1520 (N_1520,N_938,N_778);
nor U1521 (N_1521,N_307,N_817);
nand U1522 (N_1522,N_813,N_632);
nand U1523 (N_1523,N_831,N_426);
or U1524 (N_1524,N_691,N_660);
nand U1525 (N_1525,N_659,N_704);
nand U1526 (N_1526,N_191,N_513);
and U1527 (N_1527,N_223,N_571);
nand U1528 (N_1528,N_920,N_999);
nor U1529 (N_1529,N_144,N_568);
and U1530 (N_1530,N_371,N_368);
and U1531 (N_1531,N_249,N_366);
nand U1532 (N_1532,N_289,N_177);
xnor U1533 (N_1533,N_300,N_615);
nor U1534 (N_1534,N_978,N_247);
nand U1535 (N_1535,N_921,N_431);
nor U1536 (N_1536,N_555,N_516);
nor U1537 (N_1537,N_142,N_881);
and U1538 (N_1538,N_234,N_996);
or U1539 (N_1539,N_0,N_984);
and U1540 (N_1540,N_648,N_726);
and U1541 (N_1541,N_791,N_847);
or U1542 (N_1542,N_507,N_308);
and U1543 (N_1543,N_720,N_847);
and U1544 (N_1544,N_79,N_675);
nor U1545 (N_1545,N_801,N_931);
xor U1546 (N_1546,N_966,N_1);
and U1547 (N_1547,N_93,N_167);
nor U1548 (N_1548,N_245,N_401);
or U1549 (N_1549,N_319,N_475);
nand U1550 (N_1550,N_804,N_266);
or U1551 (N_1551,N_491,N_60);
nand U1552 (N_1552,N_347,N_314);
nor U1553 (N_1553,N_529,N_561);
or U1554 (N_1554,N_109,N_437);
nor U1555 (N_1555,N_341,N_958);
and U1556 (N_1556,N_448,N_262);
or U1557 (N_1557,N_711,N_514);
nand U1558 (N_1558,N_769,N_540);
nor U1559 (N_1559,N_534,N_69);
or U1560 (N_1560,N_406,N_352);
nor U1561 (N_1561,N_784,N_360);
xor U1562 (N_1562,N_424,N_842);
and U1563 (N_1563,N_995,N_356);
or U1564 (N_1564,N_678,N_866);
and U1565 (N_1565,N_319,N_774);
nor U1566 (N_1566,N_167,N_845);
nand U1567 (N_1567,N_797,N_804);
nand U1568 (N_1568,N_24,N_701);
nand U1569 (N_1569,N_575,N_73);
nand U1570 (N_1570,N_129,N_615);
xor U1571 (N_1571,N_86,N_78);
nor U1572 (N_1572,N_111,N_3);
and U1573 (N_1573,N_129,N_234);
or U1574 (N_1574,N_725,N_245);
or U1575 (N_1575,N_848,N_885);
or U1576 (N_1576,N_877,N_241);
nand U1577 (N_1577,N_377,N_429);
or U1578 (N_1578,N_529,N_249);
and U1579 (N_1579,N_373,N_35);
and U1580 (N_1580,N_570,N_937);
or U1581 (N_1581,N_471,N_324);
nand U1582 (N_1582,N_361,N_504);
and U1583 (N_1583,N_460,N_133);
nand U1584 (N_1584,N_491,N_402);
nor U1585 (N_1585,N_495,N_546);
or U1586 (N_1586,N_381,N_960);
nand U1587 (N_1587,N_676,N_606);
and U1588 (N_1588,N_636,N_864);
and U1589 (N_1589,N_362,N_347);
and U1590 (N_1590,N_967,N_558);
or U1591 (N_1591,N_964,N_902);
or U1592 (N_1592,N_780,N_337);
or U1593 (N_1593,N_736,N_502);
nand U1594 (N_1594,N_444,N_263);
nor U1595 (N_1595,N_339,N_240);
nor U1596 (N_1596,N_948,N_531);
or U1597 (N_1597,N_309,N_583);
or U1598 (N_1598,N_820,N_126);
or U1599 (N_1599,N_84,N_774);
nand U1600 (N_1600,N_292,N_293);
xor U1601 (N_1601,N_620,N_73);
nand U1602 (N_1602,N_155,N_966);
nand U1603 (N_1603,N_470,N_751);
nand U1604 (N_1604,N_416,N_39);
or U1605 (N_1605,N_122,N_518);
nor U1606 (N_1606,N_575,N_464);
and U1607 (N_1607,N_932,N_68);
and U1608 (N_1608,N_982,N_151);
and U1609 (N_1609,N_464,N_644);
nor U1610 (N_1610,N_645,N_496);
or U1611 (N_1611,N_745,N_142);
and U1612 (N_1612,N_528,N_856);
nand U1613 (N_1613,N_204,N_16);
or U1614 (N_1614,N_989,N_803);
xor U1615 (N_1615,N_227,N_883);
and U1616 (N_1616,N_951,N_402);
or U1617 (N_1617,N_704,N_646);
nand U1618 (N_1618,N_521,N_311);
or U1619 (N_1619,N_769,N_886);
nand U1620 (N_1620,N_600,N_427);
nor U1621 (N_1621,N_545,N_708);
and U1622 (N_1622,N_542,N_599);
and U1623 (N_1623,N_295,N_489);
nor U1624 (N_1624,N_436,N_10);
nand U1625 (N_1625,N_946,N_471);
or U1626 (N_1626,N_676,N_863);
or U1627 (N_1627,N_321,N_298);
nand U1628 (N_1628,N_752,N_10);
nand U1629 (N_1629,N_263,N_149);
or U1630 (N_1630,N_544,N_955);
nand U1631 (N_1631,N_167,N_166);
and U1632 (N_1632,N_30,N_299);
nand U1633 (N_1633,N_979,N_770);
nand U1634 (N_1634,N_479,N_22);
and U1635 (N_1635,N_879,N_530);
nand U1636 (N_1636,N_244,N_165);
nand U1637 (N_1637,N_601,N_459);
nand U1638 (N_1638,N_509,N_251);
or U1639 (N_1639,N_787,N_270);
and U1640 (N_1640,N_309,N_114);
nand U1641 (N_1641,N_652,N_14);
nand U1642 (N_1642,N_346,N_189);
nand U1643 (N_1643,N_531,N_526);
and U1644 (N_1644,N_947,N_603);
and U1645 (N_1645,N_703,N_761);
and U1646 (N_1646,N_692,N_897);
or U1647 (N_1647,N_877,N_373);
or U1648 (N_1648,N_423,N_180);
or U1649 (N_1649,N_807,N_999);
nand U1650 (N_1650,N_753,N_497);
or U1651 (N_1651,N_628,N_910);
xor U1652 (N_1652,N_600,N_740);
or U1653 (N_1653,N_130,N_694);
nand U1654 (N_1654,N_191,N_303);
or U1655 (N_1655,N_795,N_643);
nand U1656 (N_1656,N_868,N_194);
or U1657 (N_1657,N_700,N_10);
nand U1658 (N_1658,N_758,N_493);
and U1659 (N_1659,N_138,N_900);
and U1660 (N_1660,N_763,N_4);
xnor U1661 (N_1661,N_413,N_859);
nor U1662 (N_1662,N_325,N_35);
nand U1663 (N_1663,N_792,N_869);
or U1664 (N_1664,N_678,N_751);
xor U1665 (N_1665,N_765,N_177);
nor U1666 (N_1666,N_823,N_217);
and U1667 (N_1667,N_196,N_923);
or U1668 (N_1668,N_459,N_623);
nor U1669 (N_1669,N_552,N_836);
or U1670 (N_1670,N_517,N_406);
nor U1671 (N_1671,N_742,N_132);
nor U1672 (N_1672,N_87,N_873);
or U1673 (N_1673,N_935,N_240);
or U1674 (N_1674,N_376,N_720);
nand U1675 (N_1675,N_844,N_554);
or U1676 (N_1676,N_61,N_634);
nor U1677 (N_1677,N_446,N_865);
and U1678 (N_1678,N_538,N_899);
nand U1679 (N_1679,N_33,N_35);
nand U1680 (N_1680,N_246,N_882);
or U1681 (N_1681,N_7,N_822);
or U1682 (N_1682,N_241,N_392);
nor U1683 (N_1683,N_83,N_534);
and U1684 (N_1684,N_732,N_832);
xnor U1685 (N_1685,N_783,N_833);
and U1686 (N_1686,N_798,N_802);
nand U1687 (N_1687,N_820,N_611);
nand U1688 (N_1688,N_727,N_574);
or U1689 (N_1689,N_355,N_521);
nor U1690 (N_1690,N_849,N_374);
or U1691 (N_1691,N_307,N_352);
xor U1692 (N_1692,N_226,N_678);
and U1693 (N_1693,N_471,N_932);
or U1694 (N_1694,N_651,N_441);
or U1695 (N_1695,N_454,N_371);
nor U1696 (N_1696,N_30,N_872);
nand U1697 (N_1697,N_774,N_30);
nor U1698 (N_1698,N_509,N_581);
and U1699 (N_1699,N_689,N_409);
and U1700 (N_1700,N_963,N_261);
nor U1701 (N_1701,N_492,N_860);
nor U1702 (N_1702,N_992,N_601);
nand U1703 (N_1703,N_142,N_451);
or U1704 (N_1704,N_402,N_882);
or U1705 (N_1705,N_562,N_725);
nand U1706 (N_1706,N_329,N_635);
nand U1707 (N_1707,N_722,N_796);
and U1708 (N_1708,N_748,N_813);
nand U1709 (N_1709,N_599,N_881);
or U1710 (N_1710,N_763,N_899);
nor U1711 (N_1711,N_852,N_257);
nand U1712 (N_1712,N_943,N_552);
and U1713 (N_1713,N_507,N_133);
nor U1714 (N_1714,N_988,N_831);
and U1715 (N_1715,N_992,N_861);
or U1716 (N_1716,N_666,N_87);
and U1717 (N_1717,N_668,N_590);
nor U1718 (N_1718,N_51,N_259);
nand U1719 (N_1719,N_41,N_793);
nor U1720 (N_1720,N_305,N_215);
and U1721 (N_1721,N_70,N_599);
xor U1722 (N_1722,N_316,N_430);
xor U1723 (N_1723,N_118,N_782);
nand U1724 (N_1724,N_788,N_603);
and U1725 (N_1725,N_141,N_515);
nand U1726 (N_1726,N_67,N_465);
nand U1727 (N_1727,N_369,N_371);
or U1728 (N_1728,N_990,N_151);
and U1729 (N_1729,N_528,N_212);
nor U1730 (N_1730,N_622,N_918);
nor U1731 (N_1731,N_138,N_879);
and U1732 (N_1732,N_365,N_524);
xor U1733 (N_1733,N_996,N_748);
xnor U1734 (N_1734,N_928,N_873);
nor U1735 (N_1735,N_416,N_262);
nor U1736 (N_1736,N_172,N_470);
xnor U1737 (N_1737,N_522,N_238);
nand U1738 (N_1738,N_584,N_220);
nand U1739 (N_1739,N_713,N_850);
nand U1740 (N_1740,N_8,N_265);
and U1741 (N_1741,N_121,N_739);
nand U1742 (N_1742,N_871,N_290);
nand U1743 (N_1743,N_436,N_639);
and U1744 (N_1744,N_933,N_857);
nor U1745 (N_1745,N_136,N_133);
nand U1746 (N_1746,N_899,N_792);
or U1747 (N_1747,N_405,N_116);
or U1748 (N_1748,N_34,N_42);
nor U1749 (N_1749,N_142,N_406);
nand U1750 (N_1750,N_339,N_109);
and U1751 (N_1751,N_683,N_274);
or U1752 (N_1752,N_548,N_411);
nor U1753 (N_1753,N_331,N_718);
or U1754 (N_1754,N_927,N_76);
xnor U1755 (N_1755,N_546,N_620);
and U1756 (N_1756,N_514,N_465);
nor U1757 (N_1757,N_558,N_356);
and U1758 (N_1758,N_765,N_62);
xor U1759 (N_1759,N_940,N_167);
or U1760 (N_1760,N_922,N_171);
nand U1761 (N_1761,N_44,N_194);
or U1762 (N_1762,N_426,N_664);
nand U1763 (N_1763,N_491,N_597);
nor U1764 (N_1764,N_918,N_937);
or U1765 (N_1765,N_426,N_897);
xor U1766 (N_1766,N_577,N_473);
xnor U1767 (N_1767,N_438,N_989);
xnor U1768 (N_1768,N_538,N_43);
and U1769 (N_1769,N_973,N_41);
nor U1770 (N_1770,N_215,N_902);
and U1771 (N_1771,N_670,N_91);
nand U1772 (N_1772,N_481,N_253);
and U1773 (N_1773,N_392,N_767);
or U1774 (N_1774,N_218,N_730);
nand U1775 (N_1775,N_270,N_84);
xor U1776 (N_1776,N_289,N_758);
or U1777 (N_1777,N_275,N_924);
or U1778 (N_1778,N_594,N_994);
nor U1779 (N_1779,N_888,N_265);
and U1780 (N_1780,N_175,N_687);
and U1781 (N_1781,N_293,N_982);
or U1782 (N_1782,N_170,N_606);
nand U1783 (N_1783,N_522,N_225);
or U1784 (N_1784,N_712,N_924);
nand U1785 (N_1785,N_554,N_126);
or U1786 (N_1786,N_964,N_621);
and U1787 (N_1787,N_157,N_468);
or U1788 (N_1788,N_89,N_597);
nor U1789 (N_1789,N_13,N_119);
and U1790 (N_1790,N_479,N_994);
and U1791 (N_1791,N_874,N_237);
nand U1792 (N_1792,N_801,N_856);
or U1793 (N_1793,N_410,N_619);
nand U1794 (N_1794,N_201,N_125);
xnor U1795 (N_1795,N_807,N_603);
or U1796 (N_1796,N_392,N_799);
nor U1797 (N_1797,N_575,N_80);
nor U1798 (N_1798,N_48,N_768);
nor U1799 (N_1799,N_832,N_549);
nor U1800 (N_1800,N_248,N_628);
and U1801 (N_1801,N_915,N_8);
or U1802 (N_1802,N_149,N_772);
or U1803 (N_1803,N_474,N_988);
or U1804 (N_1804,N_530,N_606);
and U1805 (N_1805,N_784,N_368);
and U1806 (N_1806,N_37,N_885);
or U1807 (N_1807,N_383,N_71);
nand U1808 (N_1808,N_446,N_833);
nand U1809 (N_1809,N_611,N_817);
and U1810 (N_1810,N_2,N_573);
nor U1811 (N_1811,N_150,N_122);
nand U1812 (N_1812,N_163,N_248);
and U1813 (N_1813,N_26,N_327);
nor U1814 (N_1814,N_560,N_714);
nand U1815 (N_1815,N_472,N_935);
nor U1816 (N_1816,N_302,N_714);
or U1817 (N_1817,N_552,N_38);
nor U1818 (N_1818,N_882,N_828);
and U1819 (N_1819,N_791,N_819);
nand U1820 (N_1820,N_370,N_227);
or U1821 (N_1821,N_876,N_813);
or U1822 (N_1822,N_551,N_386);
or U1823 (N_1823,N_950,N_455);
xnor U1824 (N_1824,N_914,N_539);
nor U1825 (N_1825,N_809,N_634);
nor U1826 (N_1826,N_831,N_219);
and U1827 (N_1827,N_166,N_843);
and U1828 (N_1828,N_440,N_466);
or U1829 (N_1829,N_328,N_659);
nor U1830 (N_1830,N_933,N_450);
nand U1831 (N_1831,N_441,N_577);
and U1832 (N_1832,N_845,N_998);
xor U1833 (N_1833,N_826,N_163);
xnor U1834 (N_1834,N_903,N_49);
nor U1835 (N_1835,N_459,N_72);
nand U1836 (N_1836,N_232,N_690);
or U1837 (N_1837,N_523,N_281);
nand U1838 (N_1838,N_181,N_771);
xnor U1839 (N_1839,N_625,N_861);
and U1840 (N_1840,N_22,N_167);
or U1841 (N_1841,N_678,N_36);
or U1842 (N_1842,N_961,N_46);
or U1843 (N_1843,N_436,N_511);
xor U1844 (N_1844,N_905,N_1);
or U1845 (N_1845,N_460,N_494);
xor U1846 (N_1846,N_205,N_305);
nor U1847 (N_1847,N_588,N_363);
nor U1848 (N_1848,N_731,N_927);
and U1849 (N_1849,N_758,N_844);
and U1850 (N_1850,N_44,N_924);
and U1851 (N_1851,N_673,N_622);
xnor U1852 (N_1852,N_354,N_228);
xor U1853 (N_1853,N_772,N_324);
or U1854 (N_1854,N_941,N_3);
or U1855 (N_1855,N_936,N_527);
nand U1856 (N_1856,N_36,N_64);
and U1857 (N_1857,N_170,N_897);
or U1858 (N_1858,N_728,N_105);
and U1859 (N_1859,N_552,N_141);
xor U1860 (N_1860,N_491,N_607);
or U1861 (N_1861,N_876,N_444);
or U1862 (N_1862,N_701,N_690);
nand U1863 (N_1863,N_726,N_777);
nand U1864 (N_1864,N_304,N_511);
and U1865 (N_1865,N_453,N_109);
and U1866 (N_1866,N_991,N_490);
nor U1867 (N_1867,N_951,N_504);
or U1868 (N_1868,N_822,N_614);
xor U1869 (N_1869,N_567,N_774);
and U1870 (N_1870,N_829,N_568);
and U1871 (N_1871,N_863,N_236);
or U1872 (N_1872,N_581,N_169);
nand U1873 (N_1873,N_399,N_232);
or U1874 (N_1874,N_942,N_129);
nor U1875 (N_1875,N_787,N_479);
and U1876 (N_1876,N_74,N_92);
xor U1877 (N_1877,N_713,N_613);
nor U1878 (N_1878,N_360,N_100);
nor U1879 (N_1879,N_890,N_353);
xor U1880 (N_1880,N_269,N_391);
and U1881 (N_1881,N_43,N_597);
nor U1882 (N_1882,N_607,N_613);
nor U1883 (N_1883,N_979,N_822);
xor U1884 (N_1884,N_785,N_660);
and U1885 (N_1885,N_321,N_138);
or U1886 (N_1886,N_661,N_305);
nor U1887 (N_1887,N_177,N_586);
nand U1888 (N_1888,N_544,N_459);
nand U1889 (N_1889,N_667,N_433);
or U1890 (N_1890,N_697,N_147);
or U1891 (N_1891,N_896,N_62);
or U1892 (N_1892,N_874,N_980);
nor U1893 (N_1893,N_883,N_927);
and U1894 (N_1894,N_497,N_987);
nor U1895 (N_1895,N_741,N_620);
and U1896 (N_1896,N_222,N_89);
nor U1897 (N_1897,N_99,N_726);
nor U1898 (N_1898,N_115,N_219);
nor U1899 (N_1899,N_460,N_160);
and U1900 (N_1900,N_2,N_125);
and U1901 (N_1901,N_743,N_993);
xnor U1902 (N_1902,N_530,N_971);
nor U1903 (N_1903,N_577,N_566);
xor U1904 (N_1904,N_73,N_123);
or U1905 (N_1905,N_918,N_219);
and U1906 (N_1906,N_539,N_755);
or U1907 (N_1907,N_759,N_580);
nor U1908 (N_1908,N_273,N_989);
nand U1909 (N_1909,N_917,N_727);
or U1910 (N_1910,N_681,N_666);
nor U1911 (N_1911,N_907,N_136);
nand U1912 (N_1912,N_679,N_696);
xor U1913 (N_1913,N_392,N_425);
or U1914 (N_1914,N_363,N_670);
nand U1915 (N_1915,N_984,N_461);
and U1916 (N_1916,N_222,N_41);
nor U1917 (N_1917,N_671,N_714);
nor U1918 (N_1918,N_471,N_91);
or U1919 (N_1919,N_183,N_831);
and U1920 (N_1920,N_801,N_451);
nor U1921 (N_1921,N_613,N_506);
xor U1922 (N_1922,N_17,N_708);
nor U1923 (N_1923,N_18,N_638);
or U1924 (N_1924,N_496,N_243);
and U1925 (N_1925,N_445,N_220);
or U1926 (N_1926,N_537,N_795);
or U1927 (N_1927,N_849,N_349);
nand U1928 (N_1928,N_233,N_986);
and U1929 (N_1929,N_334,N_880);
nor U1930 (N_1930,N_702,N_746);
nand U1931 (N_1931,N_94,N_819);
nand U1932 (N_1932,N_183,N_976);
nand U1933 (N_1933,N_998,N_192);
xor U1934 (N_1934,N_496,N_957);
nor U1935 (N_1935,N_152,N_142);
or U1936 (N_1936,N_886,N_363);
nand U1937 (N_1937,N_802,N_425);
nand U1938 (N_1938,N_353,N_92);
nand U1939 (N_1939,N_64,N_615);
nand U1940 (N_1940,N_758,N_21);
and U1941 (N_1941,N_766,N_757);
nand U1942 (N_1942,N_233,N_97);
and U1943 (N_1943,N_281,N_269);
nor U1944 (N_1944,N_345,N_187);
nor U1945 (N_1945,N_894,N_203);
or U1946 (N_1946,N_116,N_817);
nand U1947 (N_1947,N_49,N_67);
xnor U1948 (N_1948,N_217,N_481);
nor U1949 (N_1949,N_997,N_368);
and U1950 (N_1950,N_918,N_172);
nor U1951 (N_1951,N_582,N_704);
or U1952 (N_1952,N_49,N_509);
or U1953 (N_1953,N_339,N_367);
or U1954 (N_1954,N_12,N_717);
nor U1955 (N_1955,N_482,N_656);
or U1956 (N_1956,N_764,N_584);
nor U1957 (N_1957,N_981,N_953);
and U1958 (N_1958,N_208,N_266);
nor U1959 (N_1959,N_689,N_798);
xor U1960 (N_1960,N_299,N_853);
nor U1961 (N_1961,N_760,N_194);
or U1962 (N_1962,N_454,N_279);
or U1963 (N_1963,N_518,N_561);
or U1964 (N_1964,N_340,N_794);
or U1965 (N_1965,N_422,N_306);
and U1966 (N_1966,N_408,N_549);
and U1967 (N_1967,N_39,N_787);
or U1968 (N_1968,N_465,N_553);
nor U1969 (N_1969,N_316,N_174);
nor U1970 (N_1970,N_84,N_840);
or U1971 (N_1971,N_717,N_933);
xor U1972 (N_1972,N_59,N_389);
and U1973 (N_1973,N_485,N_432);
or U1974 (N_1974,N_881,N_709);
xnor U1975 (N_1975,N_884,N_229);
and U1976 (N_1976,N_544,N_454);
nand U1977 (N_1977,N_923,N_941);
or U1978 (N_1978,N_854,N_681);
nand U1979 (N_1979,N_639,N_87);
or U1980 (N_1980,N_112,N_526);
and U1981 (N_1981,N_148,N_127);
xor U1982 (N_1982,N_687,N_355);
or U1983 (N_1983,N_820,N_579);
and U1984 (N_1984,N_273,N_404);
nor U1985 (N_1985,N_642,N_867);
nand U1986 (N_1986,N_144,N_557);
nor U1987 (N_1987,N_810,N_702);
and U1988 (N_1988,N_510,N_758);
nor U1989 (N_1989,N_337,N_358);
nand U1990 (N_1990,N_760,N_88);
nor U1991 (N_1991,N_784,N_970);
or U1992 (N_1992,N_727,N_71);
and U1993 (N_1993,N_663,N_364);
nor U1994 (N_1994,N_33,N_832);
nand U1995 (N_1995,N_947,N_533);
nand U1996 (N_1996,N_283,N_248);
nand U1997 (N_1997,N_759,N_24);
nand U1998 (N_1998,N_558,N_420);
and U1999 (N_1999,N_951,N_370);
nand U2000 (N_2000,N_1167,N_1270);
nand U2001 (N_2001,N_1768,N_1140);
or U2002 (N_2002,N_1112,N_1147);
nand U2003 (N_2003,N_1141,N_1089);
and U2004 (N_2004,N_1446,N_1781);
or U2005 (N_2005,N_1379,N_1169);
and U2006 (N_2006,N_1833,N_1544);
or U2007 (N_2007,N_1670,N_1235);
and U2008 (N_2008,N_1259,N_1420);
nand U2009 (N_2009,N_1333,N_1569);
nor U2010 (N_2010,N_1965,N_1646);
xor U2011 (N_2011,N_1184,N_1972);
or U2012 (N_2012,N_1488,N_1536);
nand U2013 (N_2013,N_1051,N_1860);
xor U2014 (N_2014,N_1880,N_1439);
nor U2015 (N_2015,N_1025,N_1717);
nor U2016 (N_2016,N_1776,N_1729);
and U2017 (N_2017,N_1579,N_1399);
or U2018 (N_2018,N_1194,N_1118);
nor U2019 (N_2019,N_1904,N_1384);
or U2020 (N_2020,N_1176,N_1044);
and U2021 (N_2021,N_1899,N_1999);
nand U2022 (N_2022,N_1724,N_1907);
nor U2023 (N_2023,N_1419,N_1257);
or U2024 (N_2024,N_1738,N_1816);
nand U2025 (N_2025,N_1897,N_1137);
nor U2026 (N_2026,N_1269,N_1351);
nor U2027 (N_2027,N_1819,N_1489);
and U2028 (N_2028,N_1688,N_1566);
and U2029 (N_2029,N_1913,N_1283);
nor U2030 (N_2030,N_1593,N_1626);
or U2031 (N_2031,N_1725,N_1540);
nor U2032 (N_2032,N_1769,N_1404);
nand U2033 (N_2033,N_1634,N_1844);
nor U2034 (N_2034,N_1715,N_1039);
nor U2035 (N_2035,N_1504,N_1817);
or U2036 (N_2036,N_1726,N_1499);
and U2037 (N_2037,N_1629,N_1614);
and U2038 (N_2038,N_1452,N_1706);
and U2039 (N_2039,N_1124,N_1615);
nor U2040 (N_2040,N_1402,N_1014);
and U2041 (N_2041,N_1699,N_1881);
and U2042 (N_2042,N_1335,N_1791);
nand U2043 (N_2043,N_1122,N_1209);
nand U2044 (N_2044,N_1447,N_1422);
and U2045 (N_2045,N_1797,N_1808);
or U2046 (N_2046,N_1391,N_1567);
nor U2047 (N_2047,N_1970,N_1749);
and U2048 (N_2048,N_1697,N_1502);
xnor U2049 (N_2049,N_1211,N_1893);
nand U2050 (N_2050,N_1059,N_1728);
nand U2051 (N_2051,N_1467,N_1950);
or U2052 (N_2052,N_1490,N_1623);
nor U2053 (N_2053,N_1500,N_1457);
and U2054 (N_2054,N_1459,N_1521);
and U2055 (N_2055,N_1081,N_1123);
nand U2056 (N_2056,N_1493,N_1694);
nor U2057 (N_2057,N_1120,N_1707);
and U2058 (N_2058,N_1066,N_1621);
or U2059 (N_2059,N_1216,N_1324);
nor U2060 (N_2060,N_1591,N_1840);
nand U2061 (N_2061,N_1987,N_1747);
or U2062 (N_2062,N_1932,N_1849);
nand U2063 (N_2063,N_1556,N_1896);
nor U2064 (N_2064,N_1698,N_1622);
xor U2065 (N_2065,N_1170,N_1474);
nor U2066 (N_2066,N_1874,N_1071);
and U2067 (N_2067,N_1289,N_1055);
and U2068 (N_2068,N_1426,N_1338);
and U2069 (N_2069,N_1941,N_1921);
and U2070 (N_2070,N_1546,N_1889);
nand U2071 (N_2071,N_1590,N_1718);
nor U2072 (N_2072,N_1804,N_1319);
nand U2073 (N_2073,N_1928,N_1454);
or U2074 (N_2074,N_1523,N_1280);
nor U2075 (N_2075,N_1750,N_1487);
nand U2076 (N_2076,N_1246,N_1101);
xor U2077 (N_2077,N_1349,N_1665);
and U2078 (N_2078,N_1719,N_1413);
xor U2079 (N_2079,N_1796,N_1472);
nor U2080 (N_2080,N_1631,N_1919);
xor U2081 (N_2081,N_1260,N_1119);
or U2082 (N_2082,N_1735,N_1346);
nor U2083 (N_2083,N_1641,N_1938);
nor U2084 (N_2084,N_1412,N_1832);
nor U2085 (N_2085,N_1818,N_1037);
nand U2086 (N_2086,N_1966,N_1276);
nand U2087 (N_2087,N_1662,N_1254);
and U2088 (N_2088,N_1625,N_1933);
or U2089 (N_2089,N_1217,N_1787);
nand U2090 (N_2090,N_1857,N_1495);
nand U2091 (N_2091,N_1403,N_1027);
or U2092 (N_2092,N_1755,N_1191);
nand U2093 (N_2093,N_1294,N_1166);
or U2094 (N_2094,N_1786,N_1416);
nand U2095 (N_2095,N_1279,N_1421);
and U2096 (N_2096,N_1160,N_1092);
nand U2097 (N_2097,N_1978,N_1182);
nor U2098 (N_2098,N_1958,N_1618);
nor U2099 (N_2099,N_1858,N_1383);
xor U2100 (N_2100,N_1063,N_1129);
nand U2101 (N_2101,N_1664,N_1306);
nor U2102 (N_2102,N_1390,N_1883);
nand U2103 (N_2103,N_1485,N_1125);
xnor U2104 (N_2104,N_1173,N_1539);
nor U2105 (N_2105,N_1853,N_1721);
nor U2106 (N_2106,N_1589,N_1028);
or U2107 (N_2107,N_1049,N_1660);
and U2108 (N_2108,N_1627,N_1636);
and U2109 (N_2109,N_1464,N_1759);
nor U2110 (N_2110,N_1237,N_1056);
or U2111 (N_2111,N_1630,N_1240);
and U2112 (N_2112,N_1741,N_1638);
and U2113 (N_2113,N_1821,N_1088);
xnor U2114 (N_2114,N_1076,N_1054);
and U2115 (N_2115,N_1115,N_1005);
nand U2116 (N_2116,N_1770,N_1991);
nand U2117 (N_2117,N_1701,N_1795);
nor U2118 (N_2118,N_1829,N_1514);
or U2119 (N_2119,N_1994,N_1029);
and U2120 (N_2120,N_1744,N_1470);
nor U2121 (N_2121,N_1764,N_1099);
nor U2122 (N_2122,N_1117,N_1372);
and U2123 (N_2123,N_1854,N_1106);
and U2124 (N_2124,N_1183,N_1923);
nor U2125 (N_2125,N_1633,N_1207);
or U2126 (N_2126,N_1433,N_1350);
or U2127 (N_2127,N_1090,N_1036);
xor U2128 (N_2128,N_1313,N_1130);
nor U2129 (N_2129,N_1398,N_1830);
and U2130 (N_2130,N_1766,N_1165);
nor U2131 (N_2131,N_1355,N_1518);
or U2132 (N_2132,N_1971,N_1551);
nor U2133 (N_2133,N_1435,N_1834);
and U2134 (N_2134,N_1332,N_1916);
or U2135 (N_2135,N_1850,N_1836);
nand U2136 (N_2136,N_1864,N_1451);
nor U2137 (N_2137,N_1347,N_1599);
nand U2138 (N_2138,N_1922,N_1802);
nor U2139 (N_2139,N_1152,N_1613);
and U2140 (N_2140,N_1360,N_1050);
and U2141 (N_2141,N_1803,N_1100);
and U2142 (N_2142,N_1924,N_1132);
or U2143 (N_2143,N_1077,N_1678);
nor U2144 (N_2144,N_1676,N_1554);
or U2145 (N_2145,N_1230,N_1918);
or U2146 (N_2146,N_1975,N_1073);
nor U2147 (N_2147,N_1635,N_1146);
nand U2148 (N_2148,N_1023,N_1507);
or U2149 (N_2149,N_1900,N_1233);
xnor U2150 (N_2150,N_1440,N_1263);
nand U2151 (N_2151,N_1714,N_1377);
and U2152 (N_2152,N_1743,N_1837);
or U2153 (N_2153,N_1356,N_1410);
and U2154 (N_2154,N_1592,N_1131);
nand U2155 (N_2155,N_1415,N_1365);
nor U2156 (N_2156,N_1920,N_1189);
and U2157 (N_2157,N_1878,N_1305);
nand U2158 (N_2158,N_1689,N_1091);
nor U2159 (N_2159,N_1597,N_1656);
nand U2160 (N_2160,N_1297,N_1926);
xnor U2161 (N_2161,N_1103,N_1142);
and U2162 (N_2162,N_1150,N_1954);
or U2163 (N_2163,N_1652,N_1847);
nand U2164 (N_2164,N_1018,N_1486);
nand U2165 (N_2165,N_1555,N_1097);
nand U2166 (N_2166,N_1534,N_1208);
xor U2167 (N_2167,N_1952,N_1824);
and U2168 (N_2168,N_1887,N_1713);
nand U2169 (N_2169,N_1530,N_1159);
or U2170 (N_2170,N_1946,N_1158);
and U2171 (N_2171,N_1058,N_1370);
and U2172 (N_2172,N_1577,N_1892);
or U2173 (N_2173,N_1595,N_1730);
and U2174 (N_2174,N_1337,N_1387);
xnor U2175 (N_2175,N_1047,N_1033);
nor U2176 (N_2176,N_1835,N_1229);
or U2177 (N_2177,N_1760,N_1069);
nand U2178 (N_2178,N_1407,N_1957);
and U2179 (N_2179,N_1161,N_1777);
nor U2180 (N_2180,N_1441,N_1692);
xnor U2181 (N_2181,N_1234,N_1790);
nor U2182 (N_2182,N_1448,N_1848);
or U2183 (N_2183,N_1449,N_1468);
or U2184 (N_2184,N_1675,N_1262);
nand U2185 (N_2185,N_1481,N_1806);
or U2186 (N_2186,N_1906,N_1855);
and U2187 (N_2187,N_1344,N_1329);
and U2188 (N_2188,N_1397,N_1653);
nand U2189 (N_2189,N_1084,N_1411);
nand U2190 (N_2190,N_1560,N_1043);
nand U2191 (N_2191,N_1248,N_1369);
xor U2192 (N_2192,N_1594,N_1484);
or U2193 (N_2193,N_1133,N_1608);
or U2194 (N_2194,N_1019,N_1282);
xor U2195 (N_2195,N_1643,N_1221);
and U2196 (N_2196,N_1982,N_1583);
and U2197 (N_2197,N_1529,N_1378);
or U2198 (N_2198,N_1375,N_1362);
or U2199 (N_2199,N_1288,N_1973);
xnor U2200 (N_2200,N_1072,N_1496);
or U2201 (N_2201,N_1574,N_1578);
nand U2202 (N_2202,N_1174,N_1308);
and U2203 (N_2203,N_1995,N_1564);
nand U2204 (N_2204,N_1515,N_1438);
nand U2205 (N_2205,N_1466,N_1767);
or U2206 (N_2206,N_1558,N_1265);
xor U2207 (N_2207,N_1526,N_1761);
or U2208 (N_2208,N_1985,N_1542);
and U2209 (N_2209,N_1060,N_1671);
or U2210 (N_2210,N_1527,N_1805);
and U2211 (N_2211,N_1709,N_1181);
or U2212 (N_2212,N_1107,N_1609);
and U2213 (N_2213,N_1061,N_1242);
nor U2214 (N_2214,N_1733,N_1748);
or U2215 (N_2215,N_1256,N_1396);
nor U2216 (N_2216,N_1205,N_1967);
nor U2217 (N_2217,N_1710,N_1992);
xnor U2218 (N_2218,N_1222,N_1223);
and U2219 (N_2219,N_1245,N_1116);
and U2220 (N_2220,N_1284,N_1648);
nor U2221 (N_2221,N_1295,N_1655);
and U2222 (N_2222,N_1762,N_1443);
nand U2223 (N_2223,N_1114,N_1164);
xnor U2224 (N_2224,N_1460,N_1911);
or U2225 (N_2225,N_1550,N_1580);
nand U2226 (N_2226,N_1996,N_1644);
nand U2227 (N_2227,N_1204,N_1405);
and U2228 (N_2228,N_1079,N_1619);
nand U2229 (N_2229,N_1884,N_1666);
or U2230 (N_2230,N_1353,N_1559);
and U2231 (N_2231,N_1156,N_1153);
or U2232 (N_2232,N_1364,N_1075);
nor U2233 (N_2233,N_1693,N_1068);
nand U2234 (N_2234,N_1905,N_1668);
xnor U2235 (N_2235,N_1311,N_1048);
nand U2236 (N_2236,N_1974,N_1557);
nand U2237 (N_2237,N_1684,N_1322);
nor U2238 (N_2238,N_1010,N_1026);
nor U2239 (N_2239,N_1732,N_1494);
nand U2240 (N_2240,N_1030,N_1479);
or U2241 (N_2241,N_1267,N_1929);
nand U2242 (N_2242,N_1022,N_1310);
and U2243 (N_2243,N_1571,N_1238);
nor U2244 (N_2244,N_1782,N_1431);
nor U2245 (N_2245,N_1154,N_1838);
xor U2246 (N_2246,N_1015,N_1581);
nand U2247 (N_2247,N_1620,N_1231);
nor U2248 (N_2248,N_1483,N_1669);
nor U2249 (N_2249,N_1930,N_1007);
and U2250 (N_2250,N_1549,N_1570);
nand U2251 (N_2251,N_1392,N_1197);
and U2252 (N_2252,N_1788,N_1745);
or U2253 (N_2253,N_1345,N_1323);
and U2254 (N_2254,N_1936,N_1406);
nor U2255 (N_2255,N_1136,N_1381);
and U2256 (N_2256,N_1192,N_1908);
nand U2257 (N_2257,N_1193,N_1417);
or U2258 (N_2258,N_1702,N_1927);
nand U2259 (N_2259,N_1888,N_1111);
and U2260 (N_2260,N_1606,N_1179);
and U2261 (N_2261,N_1374,N_1510);
or U2262 (N_2262,N_1772,N_1011);
and U2263 (N_2263,N_1842,N_1980);
or U2264 (N_2264,N_1976,N_1385);
nor U2265 (N_2265,N_1427,N_1942);
and U2266 (N_2266,N_1541,N_1278);
or U2267 (N_2267,N_1603,N_1408);
nand U2268 (N_2268,N_1708,N_1820);
and U2269 (N_2269,N_1104,N_1587);
nand U2270 (N_2270,N_1865,N_1752);
nand U2271 (N_2271,N_1241,N_1009);
nor U2272 (N_2272,N_1645,N_1582);
and U2273 (N_2273,N_1272,N_1863);
and U2274 (N_2274,N_1145,N_1418);
and U2275 (N_2275,N_1517,N_1841);
or U2276 (N_2276,N_1151,N_1754);
nand U2277 (N_2277,N_1040,N_1016);
nand U2278 (N_2278,N_1758,N_1774);
nor U2279 (N_2279,N_1846,N_1309);
xnor U2280 (N_2280,N_1711,N_1651);
and U2281 (N_2281,N_1963,N_1687);
nor U2282 (N_2282,N_1703,N_1196);
nand U2283 (N_2283,N_1912,N_1809);
and U2284 (N_2284,N_1988,N_1219);
nor U2285 (N_2285,N_1757,N_1607);
nand U2286 (N_2286,N_1180,N_1052);
nand U2287 (N_2287,N_1914,N_1303);
xor U2288 (N_2288,N_1003,N_1792);
nor U2289 (N_2289,N_1143,N_1243);
and U2290 (N_2290,N_1109,N_1255);
or U2291 (N_2291,N_1328,N_1409);
nor U2292 (N_2292,N_1469,N_1340);
nor U2293 (N_2293,N_1098,N_1281);
xor U2294 (N_2294,N_1610,N_1366);
nand U2295 (N_2295,N_1727,N_1984);
and U2296 (N_2296,N_1501,N_1685);
nand U2297 (N_2297,N_1139,N_1895);
or U2298 (N_2298,N_1277,N_1827);
nand U2299 (N_2299,N_1186,N_1178);
nor U2300 (N_2300,N_1690,N_1312);
nor U2301 (N_2301,N_1831,N_1087);
or U2302 (N_2302,N_1258,N_1909);
or U2303 (N_2303,N_1823,N_1828);
or U2304 (N_2304,N_1035,N_1275);
or U2305 (N_2305,N_1006,N_1261);
nand U2306 (N_2306,N_1352,N_1320);
or U2307 (N_2307,N_1915,N_1250);
nand U2308 (N_2308,N_1673,N_1814);
and U2309 (N_2309,N_1508,N_1882);
nor U2310 (N_2310,N_1497,N_1065);
or U2311 (N_2311,N_1017,N_1220);
or U2312 (N_2312,N_1696,N_1704);
nand U2313 (N_2313,N_1478,N_1813);
nand U2314 (N_2314,N_1773,N_1659);
or U2315 (N_2315,N_1012,N_1304);
nand U2316 (N_2316,N_1172,N_1428);
and U2317 (N_2317,N_1680,N_1198);
and U2318 (N_2318,N_1512,N_1845);
xnor U2319 (N_2319,N_1314,N_1547);
or U2320 (N_2320,N_1959,N_1476);
and U2321 (N_2321,N_1868,N_1239);
and U2322 (N_2322,N_1461,N_1095);
nand U2323 (N_2323,N_1552,N_1244);
nand U2324 (N_2324,N_1784,N_1712);
and U2325 (N_2325,N_1455,N_1851);
nor U2326 (N_2326,N_1657,N_1401);
nor U2327 (N_2327,N_1382,N_1981);
or U2328 (N_2328,N_1126,N_1424);
or U2329 (N_2329,N_1601,N_1299);
and U2330 (N_2330,N_1642,N_1810);
xor U2331 (N_2331,N_1249,N_1436);
nand U2332 (N_2332,N_1948,N_1867);
nand U2333 (N_2333,N_1292,N_1894);
xnor U2334 (N_2334,N_1336,N_1856);
nor U2335 (N_2335,N_1127,N_1661);
nand U2336 (N_2336,N_1667,N_1538);
or U2337 (N_2337,N_1826,N_1201);
or U2338 (N_2338,N_1031,N_1935);
and U2339 (N_2339,N_1640,N_1902);
nor U2340 (N_2340,N_1575,N_1765);
nand U2341 (N_2341,N_1751,N_1674);
or U2342 (N_2342,N_1519,N_1187);
nand U2343 (N_2343,N_1086,N_1825);
nor U2344 (N_2344,N_1094,N_1785);
or U2345 (N_2345,N_1380,N_1977);
or U2346 (N_2346,N_1168,N_1898);
or U2347 (N_2347,N_1993,N_1775);
or U2348 (N_2348,N_1753,N_1202);
or U2349 (N_2349,N_1979,N_1503);
xor U2350 (N_2350,N_1232,N_1064);
nand U2351 (N_2351,N_1944,N_1171);
nor U2352 (N_2352,N_1175,N_1683);
nand U2353 (N_2353,N_1799,N_1331);
nand U2354 (N_2354,N_1742,N_1839);
and U2355 (N_2355,N_1213,N_1144);
and U2356 (N_2356,N_1686,N_1548);
or U2357 (N_2357,N_1989,N_1533);
nor U2358 (N_2358,N_1389,N_1444);
and U2359 (N_2359,N_1528,N_1327);
or U2360 (N_2360,N_1866,N_1339);
nand U2361 (N_2361,N_1869,N_1600);
nand U2362 (N_2362,N_1628,N_1214);
or U2363 (N_2363,N_1298,N_1394);
or U2364 (N_2364,N_1070,N_1482);
nor U2365 (N_2365,N_1511,N_1388);
xnor U2366 (N_2366,N_1588,N_1287);
xnor U2367 (N_2367,N_1227,N_1423);
nand U2368 (N_2368,N_1074,N_1330);
nor U2369 (N_2369,N_1373,N_1870);
or U2370 (N_2370,N_1225,N_1998);
xor U2371 (N_2371,N_1334,N_1203);
or U2372 (N_2372,N_1325,N_1465);
and U2373 (N_2373,N_1218,N_1273);
and U2374 (N_2374,N_1852,N_1506);
and U2375 (N_2375,N_1135,N_1990);
and U2376 (N_2376,N_1442,N_1290);
xor U2377 (N_2377,N_1509,N_1793);
or U2378 (N_2378,N_1801,N_1157);
or U2379 (N_2379,N_1113,N_1736);
and U2380 (N_2380,N_1639,N_1199);
and U2381 (N_2381,N_1871,N_1236);
and U2382 (N_2382,N_1498,N_1962);
or U2383 (N_2383,N_1917,N_1955);
nor U2384 (N_2384,N_1960,N_1522);
or U2385 (N_2385,N_1096,N_1341);
and U2386 (N_2386,N_1318,N_1617);
or U2387 (N_2387,N_1940,N_1602);
nor U2388 (N_2388,N_1021,N_1002);
or U2389 (N_2389,N_1361,N_1317);
or U2390 (N_2390,N_1315,N_1800);
xnor U2391 (N_2391,N_1085,N_1471);
nand U2392 (N_2392,N_1672,N_1080);
or U2393 (N_2393,N_1247,N_1705);
and U2394 (N_2394,N_1939,N_1654);
or U2395 (N_2395,N_1682,N_1274);
xnor U2396 (N_2396,N_1034,N_1425);
and U2397 (N_2397,N_1524,N_1149);
nand U2398 (N_2398,N_1969,N_1658);
or U2399 (N_2399,N_1268,N_1434);
nor U2400 (N_2400,N_1343,N_1045);
nor U2401 (N_2401,N_1565,N_1576);
and U2402 (N_2402,N_1105,N_1024);
or U2403 (N_2403,N_1695,N_1462);
nand U2404 (N_2404,N_1553,N_1062);
or U2405 (N_2405,N_1445,N_1177);
and U2406 (N_2406,N_1492,N_1224);
nand U2407 (N_2407,N_1649,N_1458);
nor U2408 (N_2408,N_1739,N_1505);
and U2409 (N_2409,N_1001,N_1368);
nor U2410 (N_2410,N_1188,N_1363);
nor U2411 (N_2411,N_1376,N_1949);
and U2412 (N_2412,N_1811,N_1301);
nand U2413 (N_2413,N_1901,N_1525);
nand U2414 (N_2414,N_1945,N_1128);
nor U2415 (N_2415,N_1480,N_1367);
xnor U2416 (N_2416,N_1110,N_1561);
nor U2417 (N_2417,N_1212,N_1535);
nand U2418 (N_2418,N_1545,N_1041);
and U2419 (N_2419,N_1302,N_1450);
nor U2420 (N_2420,N_1596,N_1108);
and U2421 (N_2421,N_1134,N_1612);
or U2422 (N_2422,N_1798,N_1326);
or U2423 (N_2423,N_1354,N_1563);
nor U2424 (N_2424,N_1266,N_1605);
nor U2425 (N_2425,N_1291,N_1700);
nor U2426 (N_2426,N_1253,N_1947);
nor U2427 (N_2427,N_1677,N_1093);
nor U2428 (N_2428,N_1121,N_1843);
or U2429 (N_2429,N_1138,N_1964);
and U2430 (N_2430,N_1020,N_1162);
nand U2431 (N_2431,N_1604,N_1862);
and U2432 (N_2432,N_1453,N_1516);
or U2433 (N_2433,N_1082,N_1585);
and U2434 (N_2434,N_1475,N_1456);
xor U2435 (N_2435,N_1780,N_1859);
and U2436 (N_2436,N_1190,N_1046);
nand U2437 (N_2437,N_1910,N_1778);
nor U2438 (N_2438,N_1543,N_1042);
and U2439 (N_2439,N_1986,N_1934);
or U2440 (N_2440,N_1432,N_1632);
and U2441 (N_2441,N_1067,N_1572);
nand U2442 (N_2442,N_1357,N_1163);
xor U2443 (N_2443,N_1053,N_1206);
and U2444 (N_2444,N_1763,N_1358);
nand U2445 (N_2445,N_1891,N_1386);
nand U2446 (N_2446,N_1956,N_1722);
and U2447 (N_2447,N_1861,N_1885);
nand U2448 (N_2448,N_1740,N_1943);
nand U2449 (N_2449,N_1348,N_1890);
nand U2450 (N_2450,N_1395,N_1251);
nor U2451 (N_2451,N_1584,N_1477);
and U2452 (N_2452,N_1437,N_1771);
and U2453 (N_2453,N_1807,N_1271);
nand U2454 (N_2454,N_1731,N_1215);
nand U2455 (N_2455,N_1537,N_1210);
or U2456 (N_2456,N_1873,N_1285);
nand U2457 (N_2457,N_1815,N_1393);
and U2458 (N_2458,N_1877,N_1568);
nand U2459 (N_2459,N_1647,N_1200);
and U2460 (N_2460,N_1195,N_1812);
or U2461 (N_2461,N_1562,N_1371);
nand U2462 (N_2462,N_1886,N_1307);
or U2463 (N_2463,N_1650,N_1228);
or U2464 (N_2464,N_1875,N_1185);
and U2465 (N_2465,N_1783,N_1513);
xnor U2466 (N_2466,N_1746,N_1252);
or U2467 (N_2467,N_1316,N_1637);
nand U2468 (N_2468,N_1720,N_1903);
nor U2469 (N_2469,N_1794,N_1879);
and U2470 (N_2470,N_1155,N_1983);
or U2471 (N_2471,N_1681,N_1414);
and U2472 (N_2472,N_1078,N_1000);
nor U2473 (N_2473,N_1961,N_1057);
or U2474 (N_2474,N_1359,N_1463);
or U2475 (N_2475,N_1429,N_1679);
nand U2476 (N_2476,N_1756,N_1931);
and U2477 (N_2477,N_1008,N_1038);
nor U2478 (N_2478,N_1737,N_1822);
nand U2479 (N_2479,N_1473,N_1573);
nor U2480 (N_2480,N_1953,N_1296);
nand U2481 (N_2481,N_1321,N_1937);
and U2482 (N_2482,N_1586,N_1598);
nor U2483 (N_2483,N_1691,N_1723);
or U2484 (N_2484,N_1148,N_1789);
or U2485 (N_2485,N_1716,N_1734);
or U2486 (N_2486,N_1872,N_1624);
nand U2487 (N_2487,N_1616,N_1876);
and U2488 (N_2488,N_1226,N_1531);
or U2489 (N_2489,N_1013,N_1951);
or U2490 (N_2490,N_1430,N_1400);
nand U2491 (N_2491,N_1925,N_1032);
nor U2492 (N_2492,N_1300,N_1491);
nand U2493 (N_2493,N_1997,N_1264);
and U2494 (N_2494,N_1342,N_1102);
and U2495 (N_2495,N_1004,N_1663);
nand U2496 (N_2496,N_1083,N_1779);
xnor U2497 (N_2497,N_1286,N_1520);
nand U2498 (N_2498,N_1532,N_1293);
nor U2499 (N_2499,N_1968,N_1611);
nor U2500 (N_2500,N_1958,N_1140);
xor U2501 (N_2501,N_1204,N_1422);
or U2502 (N_2502,N_1447,N_1010);
xnor U2503 (N_2503,N_1397,N_1880);
nor U2504 (N_2504,N_1838,N_1830);
or U2505 (N_2505,N_1301,N_1818);
xor U2506 (N_2506,N_1785,N_1142);
nand U2507 (N_2507,N_1982,N_1478);
and U2508 (N_2508,N_1615,N_1940);
or U2509 (N_2509,N_1781,N_1475);
or U2510 (N_2510,N_1993,N_1284);
or U2511 (N_2511,N_1486,N_1996);
xnor U2512 (N_2512,N_1377,N_1393);
nand U2513 (N_2513,N_1225,N_1121);
nand U2514 (N_2514,N_1833,N_1781);
or U2515 (N_2515,N_1656,N_1273);
or U2516 (N_2516,N_1287,N_1470);
or U2517 (N_2517,N_1926,N_1548);
or U2518 (N_2518,N_1626,N_1632);
xor U2519 (N_2519,N_1516,N_1972);
and U2520 (N_2520,N_1452,N_1769);
and U2521 (N_2521,N_1255,N_1456);
or U2522 (N_2522,N_1167,N_1407);
nand U2523 (N_2523,N_1445,N_1908);
nor U2524 (N_2524,N_1909,N_1238);
and U2525 (N_2525,N_1810,N_1888);
or U2526 (N_2526,N_1489,N_1252);
and U2527 (N_2527,N_1406,N_1262);
and U2528 (N_2528,N_1592,N_1167);
or U2529 (N_2529,N_1457,N_1728);
or U2530 (N_2530,N_1012,N_1204);
xnor U2531 (N_2531,N_1548,N_1753);
nor U2532 (N_2532,N_1497,N_1038);
nand U2533 (N_2533,N_1138,N_1579);
or U2534 (N_2534,N_1576,N_1215);
or U2535 (N_2535,N_1111,N_1545);
nor U2536 (N_2536,N_1415,N_1091);
nand U2537 (N_2537,N_1621,N_1792);
nor U2538 (N_2538,N_1403,N_1103);
nor U2539 (N_2539,N_1136,N_1081);
and U2540 (N_2540,N_1797,N_1223);
xor U2541 (N_2541,N_1331,N_1625);
nand U2542 (N_2542,N_1086,N_1920);
xnor U2543 (N_2543,N_1858,N_1692);
nor U2544 (N_2544,N_1531,N_1970);
xnor U2545 (N_2545,N_1351,N_1352);
and U2546 (N_2546,N_1327,N_1813);
or U2547 (N_2547,N_1978,N_1222);
nand U2548 (N_2548,N_1367,N_1810);
and U2549 (N_2549,N_1580,N_1696);
xnor U2550 (N_2550,N_1775,N_1252);
nor U2551 (N_2551,N_1860,N_1786);
nand U2552 (N_2552,N_1009,N_1954);
or U2553 (N_2553,N_1155,N_1585);
or U2554 (N_2554,N_1415,N_1114);
or U2555 (N_2555,N_1831,N_1671);
and U2556 (N_2556,N_1243,N_1866);
nor U2557 (N_2557,N_1357,N_1343);
or U2558 (N_2558,N_1647,N_1813);
nand U2559 (N_2559,N_1819,N_1269);
nor U2560 (N_2560,N_1517,N_1089);
and U2561 (N_2561,N_1425,N_1271);
nand U2562 (N_2562,N_1989,N_1529);
nand U2563 (N_2563,N_1679,N_1180);
or U2564 (N_2564,N_1488,N_1681);
and U2565 (N_2565,N_1046,N_1700);
and U2566 (N_2566,N_1996,N_1788);
nand U2567 (N_2567,N_1285,N_1018);
nor U2568 (N_2568,N_1839,N_1607);
and U2569 (N_2569,N_1561,N_1623);
nand U2570 (N_2570,N_1394,N_1328);
or U2571 (N_2571,N_1135,N_1375);
nand U2572 (N_2572,N_1574,N_1794);
or U2573 (N_2573,N_1792,N_1779);
or U2574 (N_2574,N_1915,N_1553);
nor U2575 (N_2575,N_1366,N_1291);
nor U2576 (N_2576,N_1590,N_1918);
and U2577 (N_2577,N_1089,N_1228);
nand U2578 (N_2578,N_1483,N_1708);
and U2579 (N_2579,N_1515,N_1541);
or U2580 (N_2580,N_1581,N_1519);
nand U2581 (N_2581,N_1878,N_1023);
or U2582 (N_2582,N_1148,N_1254);
nand U2583 (N_2583,N_1104,N_1111);
and U2584 (N_2584,N_1550,N_1545);
or U2585 (N_2585,N_1927,N_1503);
or U2586 (N_2586,N_1654,N_1759);
and U2587 (N_2587,N_1411,N_1990);
and U2588 (N_2588,N_1364,N_1746);
nand U2589 (N_2589,N_1132,N_1004);
nor U2590 (N_2590,N_1348,N_1015);
nand U2591 (N_2591,N_1999,N_1511);
xor U2592 (N_2592,N_1744,N_1066);
and U2593 (N_2593,N_1105,N_1874);
nor U2594 (N_2594,N_1049,N_1839);
nand U2595 (N_2595,N_1442,N_1668);
nand U2596 (N_2596,N_1655,N_1075);
and U2597 (N_2597,N_1913,N_1555);
and U2598 (N_2598,N_1434,N_1265);
and U2599 (N_2599,N_1457,N_1931);
xnor U2600 (N_2600,N_1015,N_1495);
or U2601 (N_2601,N_1094,N_1146);
or U2602 (N_2602,N_1135,N_1476);
and U2603 (N_2603,N_1346,N_1166);
nand U2604 (N_2604,N_1920,N_1891);
xnor U2605 (N_2605,N_1888,N_1727);
or U2606 (N_2606,N_1009,N_1515);
or U2607 (N_2607,N_1730,N_1055);
nor U2608 (N_2608,N_1633,N_1668);
xnor U2609 (N_2609,N_1588,N_1220);
or U2610 (N_2610,N_1616,N_1336);
or U2611 (N_2611,N_1652,N_1571);
and U2612 (N_2612,N_1260,N_1853);
nand U2613 (N_2613,N_1263,N_1289);
or U2614 (N_2614,N_1661,N_1044);
nor U2615 (N_2615,N_1316,N_1337);
and U2616 (N_2616,N_1342,N_1256);
nor U2617 (N_2617,N_1504,N_1625);
nor U2618 (N_2618,N_1186,N_1613);
or U2619 (N_2619,N_1585,N_1134);
nand U2620 (N_2620,N_1537,N_1296);
and U2621 (N_2621,N_1589,N_1604);
and U2622 (N_2622,N_1738,N_1193);
nand U2623 (N_2623,N_1012,N_1351);
nor U2624 (N_2624,N_1474,N_1450);
or U2625 (N_2625,N_1531,N_1246);
or U2626 (N_2626,N_1949,N_1615);
xnor U2627 (N_2627,N_1842,N_1298);
nor U2628 (N_2628,N_1208,N_1040);
nor U2629 (N_2629,N_1913,N_1520);
nor U2630 (N_2630,N_1534,N_1958);
nand U2631 (N_2631,N_1541,N_1801);
and U2632 (N_2632,N_1935,N_1926);
or U2633 (N_2633,N_1923,N_1137);
and U2634 (N_2634,N_1642,N_1663);
or U2635 (N_2635,N_1171,N_1795);
or U2636 (N_2636,N_1329,N_1734);
or U2637 (N_2637,N_1103,N_1622);
nor U2638 (N_2638,N_1956,N_1856);
or U2639 (N_2639,N_1247,N_1899);
and U2640 (N_2640,N_1642,N_1293);
or U2641 (N_2641,N_1581,N_1564);
nor U2642 (N_2642,N_1261,N_1052);
or U2643 (N_2643,N_1553,N_1026);
nand U2644 (N_2644,N_1839,N_1236);
nor U2645 (N_2645,N_1569,N_1211);
xor U2646 (N_2646,N_1340,N_1711);
or U2647 (N_2647,N_1704,N_1532);
and U2648 (N_2648,N_1461,N_1737);
or U2649 (N_2649,N_1091,N_1677);
and U2650 (N_2650,N_1216,N_1595);
or U2651 (N_2651,N_1260,N_1076);
and U2652 (N_2652,N_1883,N_1776);
or U2653 (N_2653,N_1712,N_1016);
nand U2654 (N_2654,N_1663,N_1579);
xnor U2655 (N_2655,N_1890,N_1936);
nor U2656 (N_2656,N_1668,N_1068);
or U2657 (N_2657,N_1992,N_1615);
and U2658 (N_2658,N_1663,N_1080);
and U2659 (N_2659,N_1349,N_1994);
nand U2660 (N_2660,N_1065,N_1972);
nand U2661 (N_2661,N_1587,N_1207);
xor U2662 (N_2662,N_1139,N_1062);
or U2663 (N_2663,N_1145,N_1834);
or U2664 (N_2664,N_1784,N_1806);
and U2665 (N_2665,N_1240,N_1989);
or U2666 (N_2666,N_1397,N_1727);
nand U2667 (N_2667,N_1403,N_1718);
nand U2668 (N_2668,N_1039,N_1743);
nor U2669 (N_2669,N_1235,N_1829);
nor U2670 (N_2670,N_1718,N_1166);
xnor U2671 (N_2671,N_1051,N_1700);
nand U2672 (N_2672,N_1129,N_1407);
or U2673 (N_2673,N_1833,N_1879);
nand U2674 (N_2674,N_1952,N_1664);
and U2675 (N_2675,N_1951,N_1526);
and U2676 (N_2676,N_1079,N_1499);
or U2677 (N_2677,N_1189,N_1996);
nand U2678 (N_2678,N_1820,N_1352);
nor U2679 (N_2679,N_1582,N_1587);
nor U2680 (N_2680,N_1807,N_1824);
and U2681 (N_2681,N_1386,N_1942);
and U2682 (N_2682,N_1286,N_1460);
xor U2683 (N_2683,N_1398,N_1967);
nand U2684 (N_2684,N_1904,N_1488);
or U2685 (N_2685,N_1084,N_1690);
and U2686 (N_2686,N_1570,N_1578);
or U2687 (N_2687,N_1762,N_1244);
xor U2688 (N_2688,N_1692,N_1687);
nor U2689 (N_2689,N_1816,N_1269);
nand U2690 (N_2690,N_1058,N_1324);
nand U2691 (N_2691,N_1952,N_1010);
nor U2692 (N_2692,N_1093,N_1847);
or U2693 (N_2693,N_1957,N_1868);
or U2694 (N_2694,N_1962,N_1642);
nor U2695 (N_2695,N_1359,N_1308);
xor U2696 (N_2696,N_1725,N_1770);
or U2697 (N_2697,N_1066,N_1888);
nor U2698 (N_2698,N_1993,N_1133);
nor U2699 (N_2699,N_1047,N_1890);
nor U2700 (N_2700,N_1433,N_1987);
and U2701 (N_2701,N_1328,N_1540);
xnor U2702 (N_2702,N_1606,N_1330);
and U2703 (N_2703,N_1505,N_1010);
or U2704 (N_2704,N_1549,N_1596);
and U2705 (N_2705,N_1904,N_1598);
and U2706 (N_2706,N_1960,N_1644);
nand U2707 (N_2707,N_1891,N_1643);
or U2708 (N_2708,N_1198,N_1385);
nand U2709 (N_2709,N_1603,N_1613);
or U2710 (N_2710,N_1990,N_1483);
nand U2711 (N_2711,N_1904,N_1298);
and U2712 (N_2712,N_1059,N_1276);
and U2713 (N_2713,N_1762,N_1055);
or U2714 (N_2714,N_1326,N_1219);
or U2715 (N_2715,N_1440,N_1955);
xor U2716 (N_2716,N_1837,N_1066);
nand U2717 (N_2717,N_1849,N_1997);
and U2718 (N_2718,N_1241,N_1916);
xnor U2719 (N_2719,N_1330,N_1281);
or U2720 (N_2720,N_1474,N_1161);
and U2721 (N_2721,N_1121,N_1955);
nand U2722 (N_2722,N_1149,N_1920);
nor U2723 (N_2723,N_1377,N_1651);
nand U2724 (N_2724,N_1260,N_1035);
nor U2725 (N_2725,N_1891,N_1361);
nand U2726 (N_2726,N_1641,N_1727);
or U2727 (N_2727,N_1356,N_1474);
and U2728 (N_2728,N_1389,N_1237);
or U2729 (N_2729,N_1695,N_1135);
or U2730 (N_2730,N_1748,N_1540);
nand U2731 (N_2731,N_1444,N_1534);
or U2732 (N_2732,N_1949,N_1309);
nor U2733 (N_2733,N_1761,N_1763);
and U2734 (N_2734,N_1942,N_1018);
and U2735 (N_2735,N_1682,N_1930);
nor U2736 (N_2736,N_1686,N_1905);
nand U2737 (N_2737,N_1975,N_1308);
or U2738 (N_2738,N_1867,N_1271);
nand U2739 (N_2739,N_1768,N_1827);
nor U2740 (N_2740,N_1850,N_1084);
or U2741 (N_2741,N_1975,N_1589);
or U2742 (N_2742,N_1148,N_1931);
and U2743 (N_2743,N_1420,N_1062);
nand U2744 (N_2744,N_1416,N_1190);
nand U2745 (N_2745,N_1199,N_1936);
nand U2746 (N_2746,N_1041,N_1134);
and U2747 (N_2747,N_1727,N_1899);
nor U2748 (N_2748,N_1372,N_1936);
or U2749 (N_2749,N_1367,N_1394);
or U2750 (N_2750,N_1297,N_1686);
or U2751 (N_2751,N_1048,N_1162);
nor U2752 (N_2752,N_1453,N_1816);
nor U2753 (N_2753,N_1236,N_1862);
nor U2754 (N_2754,N_1776,N_1301);
nor U2755 (N_2755,N_1776,N_1553);
nand U2756 (N_2756,N_1473,N_1836);
xor U2757 (N_2757,N_1310,N_1837);
and U2758 (N_2758,N_1644,N_1219);
and U2759 (N_2759,N_1230,N_1871);
or U2760 (N_2760,N_1359,N_1380);
or U2761 (N_2761,N_1696,N_1279);
nand U2762 (N_2762,N_1699,N_1848);
and U2763 (N_2763,N_1971,N_1879);
nor U2764 (N_2764,N_1465,N_1441);
and U2765 (N_2765,N_1809,N_1333);
nand U2766 (N_2766,N_1009,N_1357);
nand U2767 (N_2767,N_1083,N_1454);
and U2768 (N_2768,N_1956,N_1158);
xor U2769 (N_2769,N_1306,N_1808);
or U2770 (N_2770,N_1175,N_1216);
nor U2771 (N_2771,N_1351,N_1577);
or U2772 (N_2772,N_1231,N_1731);
or U2773 (N_2773,N_1917,N_1180);
nor U2774 (N_2774,N_1068,N_1378);
nand U2775 (N_2775,N_1365,N_1760);
and U2776 (N_2776,N_1487,N_1356);
nand U2777 (N_2777,N_1883,N_1190);
and U2778 (N_2778,N_1566,N_1326);
nand U2779 (N_2779,N_1452,N_1444);
or U2780 (N_2780,N_1867,N_1487);
xor U2781 (N_2781,N_1001,N_1235);
nand U2782 (N_2782,N_1299,N_1194);
nor U2783 (N_2783,N_1028,N_1230);
and U2784 (N_2784,N_1217,N_1653);
nor U2785 (N_2785,N_1573,N_1815);
or U2786 (N_2786,N_1189,N_1651);
nor U2787 (N_2787,N_1783,N_1083);
nor U2788 (N_2788,N_1775,N_1600);
nor U2789 (N_2789,N_1457,N_1864);
xor U2790 (N_2790,N_1231,N_1725);
xor U2791 (N_2791,N_1733,N_1085);
xor U2792 (N_2792,N_1499,N_1943);
and U2793 (N_2793,N_1512,N_1457);
nand U2794 (N_2794,N_1523,N_1811);
xor U2795 (N_2795,N_1542,N_1476);
or U2796 (N_2796,N_1022,N_1777);
and U2797 (N_2797,N_1167,N_1450);
and U2798 (N_2798,N_1394,N_1353);
nor U2799 (N_2799,N_1518,N_1090);
and U2800 (N_2800,N_1380,N_1573);
nand U2801 (N_2801,N_1774,N_1631);
and U2802 (N_2802,N_1980,N_1046);
and U2803 (N_2803,N_1679,N_1963);
and U2804 (N_2804,N_1972,N_1952);
or U2805 (N_2805,N_1878,N_1875);
nand U2806 (N_2806,N_1322,N_1053);
and U2807 (N_2807,N_1729,N_1828);
or U2808 (N_2808,N_1432,N_1761);
and U2809 (N_2809,N_1442,N_1814);
nor U2810 (N_2810,N_1969,N_1913);
nand U2811 (N_2811,N_1329,N_1362);
or U2812 (N_2812,N_1477,N_1262);
and U2813 (N_2813,N_1600,N_1373);
or U2814 (N_2814,N_1077,N_1355);
and U2815 (N_2815,N_1398,N_1404);
or U2816 (N_2816,N_1507,N_1027);
xor U2817 (N_2817,N_1060,N_1338);
and U2818 (N_2818,N_1049,N_1051);
nor U2819 (N_2819,N_1994,N_1152);
and U2820 (N_2820,N_1576,N_1736);
or U2821 (N_2821,N_1806,N_1128);
nand U2822 (N_2822,N_1551,N_1432);
and U2823 (N_2823,N_1445,N_1568);
or U2824 (N_2824,N_1878,N_1439);
or U2825 (N_2825,N_1470,N_1516);
xnor U2826 (N_2826,N_1597,N_1698);
and U2827 (N_2827,N_1875,N_1902);
nand U2828 (N_2828,N_1307,N_1906);
and U2829 (N_2829,N_1204,N_1578);
nand U2830 (N_2830,N_1114,N_1684);
xor U2831 (N_2831,N_1408,N_1179);
nand U2832 (N_2832,N_1456,N_1350);
and U2833 (N_2833,N_1647,N_1277);
xnor U2834 (N_2834,N_1042,N_1714);
and U2835 (N_2835,N_1488,N_1693);
or U2836 (N_2836,N_1969,N_1475);
or U2837 (N_2837,N_1457,N_1580);
or U2838 (N_2838,N_1096,N_1585);
and U2839 (N_2839,N_1834,N_1116);
xnor U2840 (N_2840,N_1981,N_1759);
and U2841 (N_2841,N_1105,N_1888);
and U2842 (N_2842,N_1127,N_1893);
or U2843 (N_2843,N_1221,N_1146);
or U2844 (N_2844,N_1558,N_1945);
and U2845 (N_2845,N_1861,N_1851);
nand U2846 (N_2846,N_1818,N_1010);
or U2847 (N_2847,N_1277,N_1026);
and U2848 (N_2848,N_1546,N_1503);
nand U2849 (N_2849,N_1002,N_1086);
nor U2850 (N_2850,N_1072,N_1279);
or U2851 (N_2851,N_1670,N_1961);
or U2852 (N_2852,N_1771,N_1951);
nor U2853 (N_2853,N_1490,N_1071);
nand U2854 (N_2854,N_1051,N_1599);
nand U2855 (N_2855,N_1880,N_1996);
nor U2856 (N_2856,N_1635,N_1473);
nand U2857 (N_2857,N_1322,N_1161);
nor U2858 (N_2858,N_1180,N_1103);
or U2859 (N_2859,N_1826,N_1186);
or U2860 (N_2860,N_1996,N_1589);
nor U2861 (N_2861,N_1938,N_1703);
and U2862 (N_2862,N_1654,N_1821);
or U2863 (N_2863,N_1525,N_1029);
or U2864 (N_2864,N_1996,N_1403);
nor U2865 (N_2865,N_1203,N_1099);
and U2866 (N_2866,N_1782,N_1755);
nor U2867 (N_2867,N_1931,N_1503);
nand U2868 (N_2868,N_1994,N_1446);
and U2869 (N_2869,N_1198,N_1582);
xor U2870 (N_2870,N_1395,N_1065);
nand U2871 (N_2871,N_1586,N_1280);
xor U2872 (N_2872,N_1679,N_1833);
and U2873 (N_2873,N_1246,N_1536);
nor U2874 (N_2874,N_1936,N_1457);
and U2875 (N_2875,N_1441,N_1220);
and U2876 (N_2876,N_1973,N_1904);
nor U2877 (N_2877,N_1883,N_1862);
and U2878 (N_2878,N_1297,N_1214);
nor U2879 (N_2879,N_1848,N_1042);
xor U2880 (N_2880,N_1802,N_1743);
nor U2881 (N_2881,N_1554,N_1742);
and U2882 (N_2882,N_1111,N_1779);
nand U2883 (N_2883,N_1282,N_1659);
and U2884 (N_2884,N_1337,N_1604);
and U2885 (N_2885,N_1374,N_1082);
nand U2886 (N_2886,N_1361,N_1204);
and U2887 (N_2887,N_1585,N_1067);
and U2888 (N_2888,N_1181,N_1584);
nor U2889 (N_2889,N_1631,N_1065);
nand U2890 (N_2890,N_1443,N_1759);
nor U2891 (N_2891,N_1658,N_1425);
xnor U2892 (N_2892,N_1121,N_1957);
nand U2893 (N_2893,N_1785,N_1616);
or U2894 (N_2894,N_1363,N_1936);
nor U2895 (N_2895,N_1425,N_1717);
or U2896 (N_2896,N_1010,N_1117);
and U2897 (N_2897,N_1530,N_1481);
and U2898 (N_2898,N_1564,N_1369);
or U2899 (N_2899,N_1432,N_1544);
nand U2900 (N_2900,N_1847,N_1443);
nor U2901 (N_2901,N_1562,N_1190);
nor U2902 (N_2902,N_1667,N_1457);
nand U2903 (N_2903,N_1383,N_1534);
nand U2904 (N_2904,N_1790,N_1746);
nor U2905 (N_2905,N_1767,N_1627);
nor U2906 (N_2906,N_1716,N_1040);
nor U2907 (N_2907,N_1455,N_1765);
or U2908 (N_2908,N_1145,N_1047);
and U2909 (N_2909,N_1973,N_1515);
or U2910 (N_2910,N_1230,N_1248);
nor U2911 (N_2911,N_1881,N_1297);
and U2912 (N_2912,N_1871,N_1164);
and U2913 (N_2913,N_1818,N_1065);
nor U2914 (N_2914,N_1428,N_1847);
or U2915 (N_2915,N_1499,N_1092);
nor U2916 (N_2916,N_1268,N_1637);
nand U2917 (N_2917,N_1134,N_1779);
or U2918 (N_2918,N_1630,N_1351);
nor U2919 (N_2919,N_1538,N_1442);
nor U2920 (N_2920,N_1280,N_1950);
nor U2921 (N_2921,N_1444,N_1753);
nand U2922 (N_2922,N_1712,N_1257);
nand U2923 (N_2923,N_1039,N_1215);
nor U2924 (N_2924,N_1883,N_1197);
nand U2925 (N_2925,N_1704,N_1461);
or U2926 (N_2926,N_1274,N_1208);
or U2927 (N_2927,N_1389,N_1149);
nor U2928 (N_2928,N_1313,N_1542);
nor U2929 (N_2929,N_1748,N_1766);
and U2930 (N_2930,N_1226,N_1323);
or U2931 (N_2931,N_1269,N_1931);
or U2932 (N_2932,N_1620,N_1862);
nand U2933 (N_2933,N_1569,N_1705);
xor U2934 (N_2934,N_1287,N_1139);
and U2935 (N_2935,N_1277,N_1080);
nand U2936 (N_2936,N_1242,N_1283);
nand U2937 (N_2937,N_1021,N_1763);
nand U2938 (N_2938,N_1095,N_1711);
xor U2939 (N_2939,N_1804,N_1338);
nand U2940 (N_2940,N_1332,N_1706);
nand U2941 (N_2941,N_1023,N_1700);
nand U2942 (N_2942,N_1308,N_1606);
nor U2943 (N_2943,N_1711,N_1493);
nand U2944 (N_2944,N_1759,N_1670);
nor U2945 (N_2945,N_1898,N_1215);
and U2946 (N_2946,N_1534,N_1010);
or U2947 (N_2947,N_1891,N_1587);
nand U2948 (N_2948,N_1452,N_1504);
nor U2949 (N_2949,N_1366,N_1715);
or U2950 (N_2950,N_1293,N_1343);
or U2951 (N_2951,N_1088,N_1438);
nand U2952 (N_2952,N_1760,N_1279);
or U2953 (N_2953,N_1048,N_1547);
nand U2954 (N_2954,N_1889,N_1893);
xnor U2955 (N_2955,N_1952,N_1861);
or U2956 (N_2956,N_1550,N_1651);
and U2957 (N_2957,N_1551,N_1787);
xnor U2958 (N_2958,N_1860,N_1968);
nand U2959 (N_2959,N_1797,N_1781);
nor U2960 (N_2960,N_1591,N_1582);
nor U2961 (N_2961,N_1282,N_1437);
nand U2962 (N_2962,N_1514,N_1950);
or U2963 (N_2963,N_1602,N_1690);
nand U2964 (N_2964,N_1513,N_1435);
or U2965 (N_2965,N_1825,N_1557);
and U2966 (N_2966,N_1075,N_1156);
and U2967 (N_2967,N_1834,N_1287);
and U2968 (N_2968,N_1395,N_1067);
nand U2969 (N_2969,N_1569,N_1064);
nand U2970 (N_2970,N_1282,N_1693);
nor U2971 (N_2971,N_1473,N_1221);
and U2972 (N_2972,N_1929,N_1928);
nor U2973 (N_2973,N_1974,N_1611);
or U2974 (N_2974,N_1402,N_1070);
and U2975 (N_2975,N_1654,N_1570);
or U2976 (N_2976,N_1574,N_1802);
xor U2977 (N_2977,N_1808,N_1349);
or U2978 (N_2978,N_1538,N_1722);
or U2979 (N_2979,N_1177,N_1338);
and U2980 (N_2980,N_1716,N_1826);
nor U2981 (N_2981,N_1056,N_1533);
and U2982 (N_2982,N_1349,N_1696);
and U2983 (N_2983,N_1806,N_1940);
or U2984 (N_2984,N_1260,N_1572);
nor U2985 (N_2985,N_1848,N_1345);
nor U2986 (N_2986,N_1625,N_1836);
and U2987 (N_2987,N_1141,N_1157);
or U2988 (N_2988,N_1605,N_1227);
nor U2989 (N_2989,N_1104,N_1442);
nand U2990 (N_2990,N_1468,N_1025);
nor U2991 (N_2991,N_1838,N_1530);
and U2992 (N_2992,N_1680,N_1886);
nor U2993 (N_2993,N_1402,N_1927);
or U2994 (N_2994,N_1742,N_1841);
nand U2995 (N_2995,N_1071,N_1869);
nor U2996 (N_2996,N_1780,N_1679);
nand U2997 (N_2997,N_1050,N_1618);
nor U2998 (N_2998,N_1906,N_1164);
nor U2999 (N_2999,N_1938,N_1484);
nand U3000 (N_3000,N_2584,N_2776);
or U3001 (N_3001,N_2550,N_2624);
and U3002 (N_3002,N_2299,N_2231);
and U3003 (N_3003,N_2449,N_2842);
nor U3004 (N_3004,N_2951,N_2756);
nand U3005 (N_3005,N_2938,N_2676);
nand U3006 (N_3006,N_2293,N_2044);
nor U3007 (N_3007,N_2450,N_2249);
nand U3008 (N_3008,N_2551,N_2937);
or U3009 (N_3009,N_2899,N_2996);
nand U3010 (N_3010,N_2944,N_2482);
nor U3011 (N_3011,N_2206,N_2385);
or U3012 (N_3012,N_2542,N_2272);
nand U3013 (N_3013,N_2397,N_2039);
nor U3014 (N_3014,N_2957,N_2443);
xnor U3015 (N_3015,N_2400,N_2049);
and U3016 (N_3016,N_2330,N_2140);
and U3017 (N_3017,N_2526,N_2532);
xor U3018 (N_3018,N_2749,N_2402);
or U3019 (N_3019,N_2611,N_2530);
and U3020 (N_3020,N_2343,N_2429);
and U3021 (N_3021,N_2979,N_2621);
nor U3022 (N_3022,N_2900,N_2619);
nand U3023 (N_3023,N_2052,N_2080);
or U3024 (N_3024,N_2399,N_2314);
nand U3025 (N_3025,N_2684,N_2216);
nand U3026 (N_3026,N_2856,N_2181);
and U3027 (N_3027,N_2794,N_2269);
xnor U3028 (N_3028,N_2728,N_2253);
or U3029 (N_3029,N_2960,N_2552);
xnor U3030 (N_3030,N_2256,N_2566);
xor U3031 (N_3031,N_2377,N_2348);
and U3032 (N_3032,N_2378,N_2345);
xnor U3033 (N_3033,N_2664,N_2178);
and U3034 (N_3034,N_2753,N_2485);
nor U3035 (N_3035,N_2817,N_2438);
or U3036 (N_3036,N_2693,N_2478);
and U3037 (N_3037,N_2075,N_2800);
xor U3038 (N_3038,N_2025,N_2763);
or U3039 (N_3039,N_2157,N_2329);
or U3040 (N_3040,N_2846,N_2685);
nor U3041 (N_3041,N_2074,N_2189);
nand U3042 (N_3042,N_2701,N_2302);
or U3043 (N_3043,N_2872,N_2695);
and U3044 (N_3044,N_2120,N_2204);
or U3045 (N_3045,N_2839,N_2850);
and U3046 (N_3046,N_2183,N_2285);
and U3047 (N_3047,N_2862,N_2026);
and U3048 (N_3048,N_2230,N_2413);
nor U3049 (N_3049,N_2655,N_2056);
and U3050 (N_3050,N_2561,N_2512);
nor U3051 (N_3051,N_2962,N_2681);
xor U3052 (N_3052,N_2738,N_2803);
nand U3053 (N_3053,N_2018,N_2337);
nor U3054 (N_3054,N_2246,N_2130);
nor U3055 (N_3055,N_2636,N_2940);
xnor U3056 (N_3056,N_2974,N_2132);
and U3057 (N_3057,N_2755,N_2033);
nor U3058 (N_3058,N_2404,N_2241);
nand U3059 (N_3059,N_2370,N_2227);
xor U3060 (N_3060,N_2304,N_2367);
and U3061 (N_3061,N_2386,N_2929);
and U3062 (N_3062,N_2000,N_2963);
and U3063 (N_3063,N_2381,N_2912);
and U3064 (N_3064,N_2435,N_2011);
nand U3065 (N_3065,N_2459,N_2760);
nor U3066 (N_3066,N_2836,N_2423);
nor U3067 (N_3067,N_2765,N_2106);
nor U3068 (N_3068,N_2827,N_2516);
and U3069 (N_3069,N_2600,N_2163);
nand U3070 (N_3070,N_2895,N_2745);
nor U3071 (N_3071,N_2508,N_2406);
nand U3072 (N_3072,N_2631,N_2818);
and U3073 (N_3073,N_2838,N_2312);
nor U3074 (N_3074,N_2514,N_2292);
nor U3075 (N_3075,N_2109,N_2094);
and U3076 (N_3076,N_2647,N_2830);
nand U3077 (N_3077,N_2534,N_2855);
nor U3078 (N_3078,N_2139,N_2637);
nor U3079 (N_3079,N_2283,N_2721);
nand U3080 (N_3080,N_2129,N_2126);
or U3081 (N_3081,N_2644,N_2692);
and U3082 (N_3082,N_2320,N_2570);
nand U3083 (N_3083,N_2474,N_2672);
and U3084 (N_3084,N_2175,N_2034);
and U3085 (N_3085,N_2807,N_2757);
or U3086 (N_3086,N_2977,N_2980);
and U3087 (N_3087,N_2475,N_2607);
and U3088 (N_3088,N_2654,N_2324);
and U3089 (N_3089,N_2792,N_2209);
xnor U3090 (N_3090,N_2686,N_2610);
and U3091 (N_3091,N_2270,N_2440);
nand U3092 (N_3092,N_2079,N_2562);
nand U3093 (N_3093,N_2070,N_2017);
nor U3094 (N_3094,N_2541,N_2748);
or U3095 (N_3095,N_2196,N_2061);
xor U3096 (N_3096,N_2028,N_2487);
nor U3097 (N_3097,N_2113,N_2328);
nand U3098 (N_3098,N_2003,N_2789);
nand U3099 (N_3099,N_2703,N_2766);
and U3100 (N_3100,N_2221,N_2517);
and U3101 (N_3101,N_2360,N_2316);
or U3102 (N_3102,N_2356,N_2252);
and U3103 (N_3103,N_2323,N_2633);
nor U3104 (N_3104,N_2319,N_2265);
and U3105 (N_3105,N_2281,N_2573);
nor U3106 (N_3106,N_2146,N_2590);
nor U3107 (N_3107,N_2945,N_2583);
or U3108 (N_3108,N_2863,N_2086);
nand U3109 (N_3109,N_2531,N_2840);
nand U3110 (N_3110,N_2630,N_2769);
or U3111 (N_3111,N_2066,N_2407);
nand U3112 (N_3112,N_2786,N_2122);
nor U3113 (N_3113,N_2545,N_2207);
or U3114 (N_3114,N_2232,N_2772);
nand U3115 (N_3115,N_2188,N_2095);
xor U3116 (N_3116,N_2923,N_2300);
nand U3117 (N_3117,N_2499,N_2511);
nand U3118 (N_3118,N_2696,N_2100);
nor U3119 (N_3119,N_2920,N_2298);
nor U3120 (N_3120,N_2428,N_2331);
nor U3121 (N_3121,N_2442,N_2102);
nor U3122 (N_3122,N_2403,N_2362);
xnor U3123 (N_3123,N_2159,N_2361);
nor U3124 (N_3124,N_2059,N_2612);
or U3125 (N_3125,N_2816,N_2578);
nand U3126 (N_3126,N_2373,N_2812);
and U3127 (N_3127,N_2747,N_2024);
nor U3128 (N_3128,N_2355,N_2040);
nand U3129 (N_3129,N_2935,N_2447);
nand U3130 (N_3130,N_2031,N_2501);
and U3131 (N_3131,N_2649,N_2058);
nor U3132 (N_3132,N_2988,N_2617);
and U3133 (N_3133,N_2332,N_2198);
or U3134 (N_3134,N_2093,N_2942);
and U3135 (N_3135,N_2809,N_2726);
or U3136 (N_3136,N_2211,N_2594);
or U3137 (N_3137,N_2480,N_2083);
or U3138 (N_3138,N_2483,N_2598);
or U3139 (N_3139,N_2821,N_2567);
and U3140 (N_3140,N_2651,N_2173);
nor U3141 (N_3141,N_2675,N_2326);
and U3142 (N_3142,N_2767,N_2525);
or U3143 (N_3143,N_2953,N_2796);
or U3144 (N_3144,N_2894,N_2710);
or U3145 (N_3145,N_2883,N_2868);
or U3146 (N_3146,N_2089,N_2325);
xnor U3147 (N_3147,N_2553,N_2012);
or U3148 (N_3148,N_2053,N_2363);
and U3149 (N_3149,N_2461,N_2013);
nor U3150 (N_3150,N_2489,N_2847);
and U3151 (N_3151,N_2687,N_2714);
or U3152 (N_3152,N_2973,N_2983);
nor U3153 (N_3153,N_2698,N_2110);
and U3154 (N_3154,N_2214,N_2162);
nand U3155 (N_3155,N_2743,N_2364);
and U3156 (N_3156,N_2793,N_2949);
or U3157 (N_3157,N_2683,N_2864);
nand U3158 (N_3158,N_2699,N_2466);
xnor U3159 (N_3159,N_2941,N_2679);
nand U3160 (N_3160,N_2242,N_2019);
nor U3161 (N_3161,N_2690,N_2503);
and U3162 (N_3162,N_2712,N_2874);
xor U3163 (N_3163,N_2295,N_2245);
xor U3164 (N_3164,N_2563,N_2497);
and U3165 (N_3165,N_2491,N_2050);
nor U3166 (N_3166,N_2932,N_2277);
nor U3167 (N_3167,N_2990,N_2632);
nor U3168 (N_3168,N_2829,N_2455);
and U3169 (N_3169,N_2338,N_2853);
or U3170 (N_3170,N_2903,N_2898);
and U3171 (N_3171,N_2841,N_2490);
and U3172 (N_3172,N_2097,N_2010);
nor U3173 (N_3173,N_2981,N_2673);
xor U3174 (N_3174,N_2549,N_2153);
nand U3175 (N_3175,N_2218,N_2301);
xnor U3176 (N_3176,N_2509,N_2802);
or U3177 (N_3177,N_2740,N_2462);
nor U3178 (N_3178,N_2603,N_2865);
nor U3179 (N_3179,N_2365,N_2742);
xnor U3180 (N_3180,N_2523,N_2035);
and U3181 (N_3181,N_2946,N_2824);
nor U3182 (N_3182,N_2544,N_2961);
or U3183 (N_3183,N_2296,N_2234);
nand U3184 (N_3184,N_2801,N_2844);
nor U3185 (N_3185,N_2777,N_2237);
and U3186 (N_3186,N_2614,N_2652);
xor U3187 (N_3187,N_2752,N_2764);
nand U3188 (N_3188,N_2170,N_2869);
nand U3189 (N_3189,N_2638,N_2925);
nor U3190 (N_3190,N_2472,N_2306);
nand U3191 (N_3191,N_2422,N_2174);
xnor U3192 (N_3192,N_2891,N_2959);
nor U3193 (N_3193,N_2092,N_2339);
or U3194 (N_3194,N_2254,N_2613);
or U3195 (N_3195,N_2599,N_2248);
and U3196 (N_3196,N_2557,N_2885);
or U3197 (N_3197,N_2914,N_2433);
xnor U3198 (N_3198,N_2375,N_2084);
and U3199 (N_3199,N_2507,N_2782);
nor U3200 (N_3200,N_2833,N_2032);
or U3201 (N_3201,N_2352,N_2791);
nand U3202 (N_3202,N_2448,N_2555);
and U3203 (N_3203,N_2444,N_2145);
xnor U3204 (N_3204,N_2493,N_2190);
nor U3205 (N_3205,N_2470,N_2351);
or U3206 (N_3206,N_2741,N_2484);
nor U3207 (N_3207,N_2797,N_2057);
nand U3208 (N_3208,N_2203,N_2441);
or U3209 (N_3209,N_2294,N_2458);
and U3210 (N_3210,N_2823,N_2985);
or U3211 (N_3211,N_2975,N_2371);
nor U3212 (N_3212,N_2870,N_2185);
nor U3213 (N_3213,N_2917,N_2678);
and U3214 (N_3214,N_2054,N_2144);
and U3215 (N_3215,N_2349,N_2719);
or U3216 (N_3216,N_2473,N_2989);
nand U3217 (N_3217,N_2704,N_2222);
nand U3218 (N_3218,N_2783,N_2620);
or U3219 (N_3219,N_2430,N_2579);
or U3220 (N_3220,N_2987,N_2892);
nand U3221 (N_3221,N_2219,N_2434);
and U3222 (N_3222,N_2063,N_2727);
xor U3223 (N_3223,N_2498,N_2233);
nand U3224 (N_3224,N_2588,N_2119);
and U3225 (N_3225,N_2592,N_2795);
nand U3226 (N_3226,N_2528,N_2533);
and U3227 (N_3227,N_2717,N_2837);
nor U3228 (N_3228,N_2608,N_2148);
nand U3229 (N_3229,N_2004,N_2504);
nor U3230 (N_3230,N_2926,N_2554);
xnor U3231 (N_3231,N_2055,N_2315);
nand U3232 (N_3232,N_2142,N_2014);
nor U3233 (N_3233,N_2276,N_2904);
nand U3234 (N_3234,N_2723,N_2496);
and U3235 (N_3235,N_2901,N_2906);
nor U3236 (N_3236,N_2187,N_2825);
or U3237 (N_3237,N_2984,N_2918);
nand U3238 (N_3238,N_2096,N_2041);
xnor U3239 (N_3239,N_2194,N_2814);
or U3240 (N_3240,N_2569,N_2605);
nand U3241 (N_3241,N_2813,N_2069);
xor U3242 (N_3242,N_2804,N_2682);
and U3243 (N_3243,N_2280,N_2668);
or U3244 (N_3244,N_2410,N_2008);
and U3245 (N_3245,N_2709,N_2191);
nand U3246 (N_3246,N_2724,N_2849);
or U3247 (N_3247,N_2860,N_2601);
or U3248 (N_3248,N_2966,N_2597);
or U3249 (N_3249,N_2262,N_2424);
and U3250 (N_3250,N_2297,N_2820);
nor U3251 (N_3251,N_2151,N_2143);
nand U3252 (N_3252,N_2875,N_2715);
nand U3253 (N_3253,N_2284,N_2288);
or U3254 (N_3254,N_2409,N_2215);
or U3255 (N_3255,N_2273,N_2716);
or U3256 (N_3256,N_2379,N_2662);
nand U3257 (N_3257,N_2006,N_2425);
and U3258 (N_3258,N_2537,N_2972);
nor U3259 (N_3259,N_2858,N_2346);
and U3260 (N_3260,N_2971,N_2733);
nand U3261 (N_3261,N_2398,N_2778);
and U3262 (N_3262,N_2759,N_2832);
and U3263 (N_3263,N_2595,N_2744);
and U3264 (N_3264,N_2604,N_2477);
nand U3265 (N_3265,N_2088,N_2780);
or U3266 (N_3266,N_2394,N_2307);
nor U3267 (N_3267,N_2111,N_2546);
or U3268 (N_3268,N_2002,N_2958);
or U3269 (N_3269,N_2943,N_2226);
or U3270 (N_3270,N_2609,N_2691);
nor U3271 (N_3271,N_2420,N_2736);
nand U3272 (N_3272,N_2665,N_2656);
and U3273 (N_3273,N_2457,N_2411);
and U3274 (N_3274,N_2939,N_2529);
nor U3275 (N_3275,N_2171,N_2910);
nor U3276 (N_3276,N_2141,N_2043);
xnor U3277 (N_3277,N_2009,N_2626);
or U3278 (N_3278,N_2176,N_2581);
nor U3279 (N_3279,N_2852,N_2392);
and U3280 (N_3280,N_2826,N_2197);
and U3281 (N_3281,N_2382,N_2225);
and U3282 (N_3282,N_2166,N_2785);
or U3283 (N_3283,N_2368,N_2967);
and U3284 (N_3284,N_2065,N_2118);
or U3285 (N_3285,N_2660,N_2488);
xor U3286 (N_3286,N_2916,N_2154);
and U3287 (N_3287,N_2469,N_2634);
or U3288 (N_3288,N_2815,N_2229);
and U3289 (N_3289,N_2344,N_2384);
nor U3290 (N_3290,N_2155,N_2418);
nand U3291 (N_3291,N_2463,N_2124);
nand U3292 (N_3292,N_2282,N_2150);
nor U3293 (N_3293,N_2376,N_2762);
or U3294 (N_3294,N_2205,N_2027);
or U3295 (N_3295,N_2831,N_2341);
nand U3296 (N_3296,N_2495,N_2152);
nand U3297 (N_3297,N_2184,N_2164);
and U3298 (N_3298,N_2243,N_2548);
or U3299 (N_3299,N_2720,N_2628);
nor U3300 (N_3300,N_2125,N_2543);
xor U3301 (N_3301,N_2771,N_2890);
or U3302 (N_3302,N_2915,N_2730);
xnor U3303 (N_3303,N_2121,N_2342);
and U3304 (N_3304,N_2414,N_2072);
and U3305 (N_3305,N_2774,N_2224);
xor U3306 (N_3306,N_2133,N_2580);
nor U3307 (N_3307,N_2560,N_2201);
nor U3308 (N_3308,N_2278,N_2023);
nand U3309 (N_3309,N_2635,N_2082);
or U3310 (N_3310,N_2020,N_2305);
nand U3311 (N_3311,N_2978,N_2258);
xor U3312 (N_3312,N_2922,N_2212);
and U3313 (N_3313,N_2689,N_2021);
and U3314 (N_3314,N_2822,N_2286);
and U3315 (N_3315,N_2976,N_2811);
nor U3316 (N_3316,N_2471,N_2706);
nor U3317 (N_3317,N_2108,N_2220);
xnor U3318 (N_3318,N_2333,N_2536);
and U3319 (N_3319,N_2653,N_2334);
or U3320 (N_3320,N_2722,N_2453);
nand U3321 (N_3321,N_2643,N_2354);
nor U3322 (N_3322,N_2454,N_2877);
nand U3323 (N_3323,N_2876,N_2582);
and U3324 (N_3324,N_2415,N_2629);
or U3325 (N_3325,N_2456,N_2993);
nor U3326 (N_3326,N_2167,N_2257);
or U3327 (N_3327,N_2623,N_2880);
or U3328 (N_3328,N_2650,N_2436);
and U3329 (N_3329,N_2700,N_2213);
and U3330 (N_3330,N_2437,N_2930);
nand U3331 (N_3331,N_2587,N_2103);
nor U3332 (N_3332,N_2357,N_2029);
nand U3333 (N_3333,N_2866,N_2223);
or U3334 (N_3334,N_2734,N_2663);
and U3335 (N_3335,N_2161,N_2513);
or U3336 (N_3336,N_2835,N_2287);
and U3337 (N_3337,N_2107,N_2138);
or U3338 (N_3338,N_2834,N_2098);
nor U3339 (N_3339,N_2640,N_2073);
nand U3340 (N_3340,N_2547,N_2087);
and U3341 (N_3341,N_2688,N_2347);
nand U3342 (N_3342,N_2431,N_2998);
or U3343 (N_3343,N_2228,N_2666);
nor U3344 (N_3344,N_2558,N_2136);
nor U3345 (N_3345,N_2182,N_2001);
nand U3346 (N_3346,N_2535,N_2180);
or U3347 (N_3347,N_2947,N_2193);
nor U3348 (N_3348,N_2905,N_2538);
xnor U3349 (N_3349,N_2559,N_2667);
xnor U3350 (N_3350,N_2335,N_2494);
xor U3351 (N_3351,N_2104,N_2085);
nand U3352 (N_3352,N_2067,N_2768);
or U3353 (N_3353,N_2479,N_2460);
nand U3354 (N_3354,N_2519,N_2127);
or U3355 (N_3355,N_2888,N_2867);
or U3356 (N_3356,N_2680,N_2149);
or U3357 (N_3357,N_2658,N_2327);
and U3358 (N_3358,N_2308,N_2571);
xnor U3359 (N_3359,N_2845,N_2168);
xnor U3360 (N_3360,N_2955,N_2303);
nand U3361 (N_3361,N_2627,N_2808);
nor U3362 (N_3362,N_2260,N_2991);
nor U3363 (N_3363,N_2670,N_2037);
or U3364 (N_3364,N_2279,N_2585);
nor U3365 (N_3365,N_2819,N_2886);
nor U3366 (N_3366,N_2077,N_2051);
or U3367 (N_3367,N_2893,N_2179);
nor U3368 (N_3368,N_2238,N_2005);
and U3369 (N_3369,N_2401,N_2317);
or U3370 (N_3370,N_2854,N_2199);
nor U3371 (N_3371,N_2950,N_2255);
or U3372 (N_3372,N_2881,N_2986);
xor U3373 (N_3373,N_2773,N_2432);
or U3374 (N_3374,N_2677,N_2353);
or U3375 (N_3375,N_2309,N_2732);
and U3376 (N_3376,N_2596,N_2235);
nand U3377 (N_3377,N_2873,N_2520);
or U3378 (N_3378,N_2564,N_2669);
or U3379 (N_3379,N_2421,N_2907);
xor U3380 (N_3380,N_2236,N_2417);
nor U3381 (N_3381,N_2202,N_2731);
nor U3382 (N_3382,N_2746,N_2165);
nand U3383 (N_3383,N_2340,N_2572);
or U3384 (N_3384,N_2468,N_2135);
and U3385 (N_3385,N_2574,N_2527);
and U3386 (N_3386,N_2289,N_2933);
xor U3387 (N_3387,N_2851,N_2291);
nand U3388 (N_3388,N_2311,N_2046);
or U3389 (N_3389,N_2586,N_2405);
and U3390 (N_3390,N_2030,N_2169);
or U3391 (N_3391,N_2446,N_2952);
xnor U3392 (N_3392,N_2318,N_2408);
or U3393 (N_3393,N_2799,N_2908);
or U3394 (N_3394,N_2515,N_2045);
nand U3395 (N_3395,N_2806,N_2936);
or U3396 (N_3396,N_2648,N_2048);
nor U3397 (N_3397,N_2467,N_2843);
or U3398 (N_3398,N_2101,N_2123);
nor U3399 (N_3399,N_2391,N_2240);
or U3400 (N_3400,N_2502,N_2758);
nand U3401 (N_3401,N_2770,N_2787);
nand U3402 (N_3402,N_2476,N_2116);
nor U3403 (N_3403,N_2622,N_2128);
and U3404 (N_3404,N_2964,N_2387);
or U3405 (N_3405,N_2518,N_2884);
or U3406 (N_3406,N_2956,N_2389);
and U3407 (N_3407,N_2871,N_2576);
nor U3408 (N_3408,N_2659,N_2995);
or U3409 (N_3409,N_2137,N_2322);
nor U3410 (N_3410,N_2992,N_2913);
nor U3411 (N_3411,N_2705,N_2556);
and U3412 (N_3412,N_2646,N_2336);
nand U3413 (N_3413,N_2761,N_2713);
or U3414 (N_3414,N_2754,N_2451);
nand U3415 (N_3415,N_2396,N_2071);
and U3416 (N_3416,N_2358,N_2896);
and U3417 (N_3417,N_2697,N_2909);
or U3418 (N_3418,N_2718,N_2158);
nor U3419 (N_3419,N_2439,N_2022);
nor U3420 (N_3420,N_2060,N_2982);
and U3421 (N_3421,N_2062,N_2016);
and U3422 (N_3422,N_2393,N_2593);
nand U3423 (N_3423,N_2195,N_2239);
nand U3424 (N_3424,N_2729,N_2810);
nand U3425 (N_3425,N_2115,N_2625);
and U3426 (N_3426,N_2994,N_2419);
or U3427 (N_3427,N_2390,N_2274);
and U3428 (N_3428,N_2200,N_2112);
nand U3429 (N_3429,N_2618,N_2192);
and U3430 (N_3430,N_2751,N_2134);
or U3431 (N_3431,N_2510,N_2383);
or U3432 (N_3432,N_2244,N_2091);
nor U3433 (N_3433,N_2694,N_2735);
or U3434 (N_3434,N_2268,N_2708);
or U3435 (N_3435,N_2412,N_2263);
nand U3436 (N_3436,N_2969,N_2575);
nand U3437 (N_3437,N_2805,N_2264);
or U3438 (N_3438,N_2591,N_2902);
or U3439 (N_3439,N_2271,N_2522);
xnor U3440 (N_3440,N_2105,N_2388);
nand U3441 (N_3441,N_2464,N_2452);
nor U3442 (N_3442,N_2878,N_2372);
nand U3443 (N_3443,N_2968,N_2321);
nor U3444 (N_3444,N_2064,N_2275);
nand U3445 (N_3445,N_2251,N_2078);
and U3446 (N_3446,N_2313,N_2036);
or U3447 (N_3447,N_2038,N_2426);
nor U3448 (N_3448,N_2310,N_2359);
or U3449 (N_3449,N_2047,N_2565);
nor U3450 (N_3450,N_2879,N_2928);
nand U3451 (N_3451,N_2911,N_2861);
and U3452 (N_3452,N_2999,N_2674);
and U3453 (N_3453,N_2707,N_2784);
and U3454 (N_3454,N_2750,N_2954);
and U3455 (N_3455,N_2828,N_2639);
nand U3456 (N_3456,N_2859,N_2076);
and U3457 (N_3457,N_2117,N_2156);
and U3458 (N_3458,N_2090,N_2711);
nand U3459 (N_3459,N_2350,N_2539);
xor U3460 (N_3460,N_2486,N_2970);
and U3461 (N_3461,N_2781,N_2427);
or U3462 (N_3462,N_2099,N_2481);
or U3463 (N_3463,N_2889,N_2924);
or U3464 (N_3464,N_2177,N_2395);
or U3465 (N_3465,N_2261,N_2465);
and U3466 (N_3466,N_2882,N_2506);
or U3467 (N_3467,N_2661,N_2948);
or U3468 (N_3468,N_2775,N_2589);
or U3469 (N_3469,N_2931,N_2500);
nor U3470 (N_3470,N_2857,N_2250);
and U3471 (N_3471,N_2416,N_2247);
nor U3472 (N_3472,N_2208,N_2210);
nand U3473 (N_3473,N_2725,N_2790);
nand U3474 (N_3474,N_2641,N_2131);
and U3475 (N_3475,N_2259,N_2927);
or U3476 (N_3476,N_2068,N_2897);
and U3477 (N_3477,N_2266,N_2997);
nor U3478 (N_3478,N_2934,N_2267);
and U3479 (N_3479,N_2606,N_2615);
and U3480 (N_3480,N_2172,N_2540);
nor U3481 (N_3481,N_2737,N_2380);
or U3482 (N_3482,N_2568,N_2290);
nand U3483 (N_3483,N_2147,N_2160);
nor U3484 (N_3484,N_2739,N_2645);
or U3485 (N_3485,N_2616,N_2217);
nand U3486 (N_3486,N_2042,N_2848);
nand U3487 (N_3487,N_2492,N_2779);
xor U3488 (N_3488,N_2702,N_2788);
nand U3489 (N_3489,N_2374,N_2887);
or U3490 (N_3490,N_2369,N_2366);
or U3491 (N_3491,N_2081,N_2671);
and U3492 (N_3492,N_2657,N_2642);
or U3493 (N_3493,N_2524,N_2965);
or U3494 (N_3494,N_2505,N_2114);
nand U3495 (N_3495,N_2602,N_2445);
and U3496 (N_3496,N_2577,N_2921);
xnor U3497 (N_3497,N_2007,N_2798);
and U3498 (N_3498,N_2015,N_2521);
nand U3499 (N_3499,N_2186,N_2919);
and U3500 (N_3500,N_2841,N_2193);
or U3501 (N_3501,N_2927,N_2773);
nor U3502 (N_3502,N_2213,N_2741);
or U3503 (N_3503,N_2823,N_2640);
and U3504 (N_3504,N_2386,N_2820);
nor U3505 (N_3505,N_2906,N_2419);
nand U3506 (N_3506,N_2958,N_2618);
or U3507 (N_3507,N_2909,N_2476);
xnor U3508 (N_3508,N_2434,N_2528);
nand U3509 (N_3509,N_2624,N_2617);
or U3510 (N_3510,N_2370,N_2818);
xor U3511 (N_3511,N_2604,N_2824);
nand U3512 (N_3512,N_2501,N_2329);
nand U3513 (N_3513,N_2999,N_2928);
nand U3514 (N_3514,N_2568,N_2553);
nand U3515 (N_3515,N_2435,N_2461);
xnor U3516 (N_3516,N_2227,N_2713);
nor U3517 (N_3517,N_2737,N_2492);
nand U3518 (N_3518,N_2426,N_2955);
nand U3519 (N_3519,N_2475,N_2533);
and U3520 (N_3520,N_2523,N_2240);
and U3521 (N_3521,N_2720,N_2786);
or U3522 (N_3522,N_2639,N_2181);
or U3523 (N_3523,N_2683,N_2383);
or U3524 (N_3524,N_2734,N_2133);
nor U3525 (N_3525,N_2785,N_2884);
nor U3526 (N_3526,N_2353,N_2044);
or U3527 (N_3527,N_2650,N_2761);
nand U3528 (N_3528,N_2974,N_2748);
nand U3529 (N_3529,N_2233,N_2511);
or U3530 (N_3530,N_2243,N_2126);
nand U3531 (N_3531,N_2261,N_2412);
nand U3532 (N_3532,N_2611,N_2438);
xnor U3533 (N_3533,N_2415,N_2328);
nor U3534 (N_3534,N_2248,N_2083);
and U3535 (N_3535,N_2849,N_2540);
or U3536 (N_3536,N_2562,N_2755);
nor U3537 (N_3537,N_2688,N_2419);
or U3538 (N_3538,N_2057,N_2386);
nand U3539 (N_3539,N_2351,N_2868);
nor U3540 (N_3540,N_2386,N_2750);
and U3541 (N_3541,N_2524,N_2443);
nand U3542 (N_3542,N_2342,N_2971);
nor U3543 (N_3543,N_2677,N_2393);
xnor U3544 (N_3544,N_2411,N_2661);
nand U3545 (N_3545,N_2196,N_2901);
or U3546 (N_3546,N_2294,N_2805);
xor U3547 (N_3547,N_2156,N_2073);
nor U3548 (N_3548,N_2559,N_2932);
nor U3549 (N_3549,N_2112,N_2970);
or U3550 (N_3550,N_2343,N_2475);
nor U3551 (N_3551,N_2317,N_2440);
xnor U3552 (N_3552,N_2347,N_2663);
nor U3553 (N_3553,N_2863,N_2342);
or U3554 (N_3554,N_2049,N_2268);
or U3555 (N_3555,N_2907,N_2773);
nor U3556 (N_3556,N_2425,N_2060);
nand U3557 (N_3557,N_2069,N_2263);
and U3558 (N_3558,N_2808,N_2259);
or U3559 (N_3559,N_2475,N_2238);
or U3560 (N_3560,N_2447,N_2243);
and U3561 (N_3561,N_2621,N_2972);
nand U3562 (N_3562,N_2234,N_2876);
nor U3563 (N_3563,N_2864,N_2375);
nand U3564 (N_3564,N_2049,N_2592);
and U3565 (N_3565,N_2302,N_2810);
or U3566 (N_3566,N_2336,N_2987);
nand U3567 (N_3567,N_2170,N_2964);
nor U3568 (N_3568,N_2175,N_2803);
nor U3569 (N_3569,N_2066,N_2642);
nand U3570 (N_3570,N_2002,N_2953);
or U3571 (N_3571,N_2425,N_2045);
nand U3572 (N_3572,N_2337,N_2491);
nor U3573 (N_3573,N_2781,N_2489);
nor U3574 (N_3574,N_2367,N_2091);
or U3575 (N_3575,N_2312,N_2376);
or U3576 (N_3576,N_2725,N_2413);
or U3577 (N_3577,N_2695,N_2311);
nand U3578 (N_3578,N_2908,N_2426);
nand U3579 (N_3579,N_2086,N_2541);
nor U3580 (N_3580,N_2056,N_2034);
xor U3581 (N_3581,N_2691,N_2867);
and U3582 (N_3582,N_2292,N_2318);
nor U3583 (N_3583,N_2226,N_2521);
and U3584 (N_3584,N_2448,N_2016);
nand U3585 (N_3585,N_2378,N_2850);
nand U3586 (N_3586,N_2861,N_2800);
nor U3587 (N_3587,N_2372,N_2903);
xnor U3588 (N_3588,N_2293,N_2929);
or U3589 (N_3589,N_2848,N_2683);
or U3590 (N_3590,N_2172,N_2344);
and U3591 (N_3591,N_2536,N_2156);
and U3592 (N_3592,N_2277,N_2378);
and U3593 (N_3593,N_2251,N_2973);
or U3594 (N_3594,N_2271,N_2689);
or U3595 (N_3595,N_2570,N_2257);
nand U3596 (N_3596,N_2904,N_2464);
nor U3597 (N_3597,N_2294,N_2991);
or U3598 (N_3598,N_2639,N_2106);
nor U3599 (N_3599,N_2373,N_2408);
and U3600 (N_3600,N_2281,N_2033);
xor U3601 (N_3601,N_2805,N_2293);
nor U3602 (N_3602,N_2530,N_2634);
nor U3603 (N_3603,N_2764,N_2534);
xnor U3604 (N_3604,N_2239,N_2196);
nand U3605 (N_3605,N_2394,N_2727);
xnor U3606 (N_3606,N_2534,N_2521);
nor U3607 (N_3607,N_2992,N_2033);
nand U3608 (N_3608,N_2894,N_2412);
or U3609 (N_3609,N_2940,N_2860);
or U3610 (N_3610,N_2461,N_2072);
and U3611 (N_3611,N_2399,N_2238);
xnor U3612 (N_3612,N_2066,N_2925);
nand U3613 (N_3613,N_2393,N_2585);
nand U3614 (N_3614,N_2959,N_2908);
nand U3615 (N_3615,N_2519,N_2997);
and U3616 (N_3616,N_2012,N_2077);
nor U3617 (N_3617,N_2871,N_2722);
and U3618 (N_3618,N_2416,N_2924);
or U3619 (N_3619,N_2779,N_2523);
and U3620 (N_3620,N_2982,N_2273);
or U3621 (N_3621,N_2036,N_2605);
xnor U3622 (N_3622,N_2408,N_2490);
nor U3623 (N_3623,N_2095,N_2045);
or U3624 (N_3624,N_2082,N_2809);
or U3625 (N_3625,N_2671,N_2311);
nand U3626 (N_3626,N_2074,N_2110);
or U3627 (N_3627,N_2727,N_2284);
nand U3628 (N_3628,N_2827,N_2096);
nand U3629 (N_3629,N_2146,N_2393);
nor U3630 (N_3630,N_2168,N_2859);
nor U3631 (N_3631,N_2189,N_2355);
nand U3632 (N_3632,N_2551,N_2027);
or U3633 (N_3633,N_2088,N_2816);
and U3634 (N_3634,N_2573,N_2038);
and U3635 (N_3635,N_2133,N_2104);
nor U3636 (N_3636,N_2932,N_2249);
nand U3637 (N_3637,N_2283,N_2403);
or U3638 (N_3638,N_2684,N_2206);
or U3639 (N_3639,N_2335,N_2334);
or U3640 (N_3640,N_2333,N_2566);
nand U3641 (N_3641,N_2561,N_2713);
nor U3642 (N_3642,N_2887,N_2481);
nand U3643 (N_3643,N_2522,N_2658);
nand U3644 (N_3644,N_2229,N_2218);
or U3645 (N_3645,N_2421,N_2049);
and U3646 (N_3646,N_2582,N_2827);
and U3647 (N_3647,N_2312,N_2478);
nor U3648 (N_3648,N_2075,N_2733);
or U3649 (N_3649,N_2264,N_2578);
nor U3650 (N_3650,N_2313,N_2912);
nand U3651 (N_3651,N_2174,N_2404);
nor U3652 (N_3652,N_2452,N_2947);
and U3653 (N_3653,N_2143,N_2137);
or U3654 (N_3654,N_2926,N_2482);
nand U3655 (N_3655,N_2523,N_2385);
and U3656 (N_3656,N_2756,N_2996);
or U3657 (N_3657,N_2777,N_2937);
nor U3658 (N_3658,N_2695,N_2595);
or U3659 (N_3659,N_2550,N_2955);
nor U3660 (N_3660,N_2554,N_2761);
nand U3661 (N_3661,N_2529,N_2309);
nand U3662 (N_3662,N_2831,N_2217);
xor U3663 (N_3663,N_2356,N_2581);
nor U3664 (N_3664,N_2334,N_2012);
or U3665 (N_3665,N_2652,N_2454);
or U3666 (N_3666,N_2370,N_2130);
nor U3667 (N_3667,N_2060,N_2751);
and U3668 (N_3668,N_2293,N_2300);
nand U3669 (N_3669,N_2636,N_2524);
nand U3670 (N_3670,N_2233,N_2246);
or U3671 (N_3671,N_2437,N_2332);
or U3672 (N_3672,N_2184,N_2707);
xor U3673 (N_3673,N_2062,N_2329);
nor U3674 (N_3674,N_2748,N_2040);
nor U3675 (N_3675,N_2745,N_2158);
or U3676 (N_3676,N_2723,N_2702);
nor U3677 (N_3677,N_2228,N_2877);
or U3678 (N_3678,N_2102,N_2681);
nor U3679 (N_3679,N_2722,N_2807);
nand U3680 (N_3680,N_2671,N_2503);
and U3681 (N_3681,N_2092,N_2602);
nor U3682 (N_3682,N_2956,N_2483);
or U3683 (N_3683,N_2959,N_2272);
nand U3684 (N_3684,N_2097,N_2943);
nor U3685 (N_3685,N_2883,N_2293);
nand U3686 (N_3686,N_2313,N_2316);
nor U3687 (N_3687,N_2817,N_2914);
nor U3688 (N_3688,N_2783,N_2425);
or U3689 (N_3689,N_2214,N_2368);
nand U3690 (N_3690,N_2626,N_2836);
nor U3691 (N_3691,N_2024,N_2077);
xnor U3692 (N_3692,N_2052,N_2575);
nand U3693 (N_3693,N_2371,N_2349);
nand U3694 (N_3694,N_2773,N_2279);
and U3695 (N_3695,N_2348,N_2541);
and U3696 (N_3696,N_2937,N_2985);
or U3697 (N_3697,N_2793,N_2051);
nor U3698 (N_3698,N_2659,N_2299);
or U3699 (N_3699,N_2615,N_2648);
nor U3700 (N_3700,N_2342,N_2258);
and U3701 (N_3701,N_2127,N_2452);
and U3702 (N_3702,N_2624,N_2754);
and U3703 (N_3703,N_2810,N_2131);
xor U3704 (N_3704,N_2735,N_2119);
or U3705 (N_3705,N_2464,N_2998);
or U3706 (N_3706,N_2251,N_2932);
and U3707 (N_3707,N_2579,N_2263);
nor U3708 (N_3708,N_2668,N_2930);
and U3709 (N_3709,N_2999,N_2719);
nand U3710 (N_3710,N_2128,N_2563);
nor U3711 (N_3711,N_2247,N_2571);
nor U3712 (N_3712,N_2337,N_2306);
or U3713 (N_3713,N_2660,N_2551);
nand U3714 (N_3714,N_2924,N_2079);
and U3715 (N_3715,N_2465,N_2963);
and U3716 (N_3716,N_2567,N_2930);
and U3717 (N_3717,N_2448,N_2618);
nand U3718 (N_3718,N_2480,N_2113);
nand U3719 (N_3719,N_2004,N_2297);
and U3720 (N_3720,N_2595,N_2846);
nor U3721 (N_3721,N_2917,N_2260);
or U3722 (N_3722,N_2140,N_2071);
and U3723 (N_3723,N_2766,N_2878);
and U3724 (N_3724,N_2942,N_2799);
and U3725 (N_3725,N_2241,N_2424);
xnor U3726 (N_3726,N_2838,N_2422);
or U3727 (N_3727,N_2472,N_2968);
nor U3728 (N_3728,N_2116,N_2166);
or U3729 (N_3729,N_2683,N_2914);
nand U3730 (N_3730,N_2396,N_2305);
and U3731 (N_3731,N_2474,N_2271);
or U3732 (N_3732,N_2007,N_2195);
nor U3733 (N_3733,N_2987,N_2114);
and U3734 (N_3734,N_2119,N_2342);
nand U3735 (N_3735,N_2101,N_2681);
or U3736 (N_3736,N_2891,N_2082);
nor U3737 (N_3737,N_2128,N_2815);
nand U3738 (N_3738,N_2577,N_2843);
and U3739 (N_3739,N_2785,N_2192);
or U3740 (N_3740,N_2979,N_2835);
nand U3741 (N_3741,N_2851,N_2354);
nand U3742 (N_3742,N_2266,N_2767);
and U3743 (N_3743,N_2945,N_2925);
or U3744 (N_3744,N_2702,N_2103);
nor U3745 (N_3745,N_2534,N_2399);
and U3746 (N_3746,N_2411,N_2544);
nor U3747 (N_3747,N_2197,N_2585);
or U3748 (N_3748,N_2387,N_2325);
xnor U3749 (N_3749,N_2713,N_2663);
xnor U3750 (N_3750,N_2506,N_2518);
and U3751 (N_3751,N_2312,N_2137);
or U3752 (N_3752,N_2635,N_2605);
nand U3753 (N_3753,N_2586,N_2166);
and U3754 (N_3754,N_2463,N_2275);
and U3755 (N_3755,N_2831,N_2287);
and U3756 (N_3756,N_2331,N_2978);
and U3757 (N_3757,N_2630,N_2633);
xnor U3758 (N_3758,N_2314,N_2378);
nor U3759 (N_3759,N_2766,N_2045);
nand U3760 (N_3760,N_2706,N_2609);
and U3761 (N_3761,N_2395,N_2726);
nor U3762 (N_3762,N_2380,N_2789);
nand U3763 (N_3763,N_2560,N_2084);
and U3764 (N_3764,N_2617,N_2444);
or U3765 (N_3765,N_2478,N_2855);
and U3766 (N_3766,N_2928,N_2516);
and U3767 (N_3767,N_2610,N_2225);
nand U3768 (N_3768,N_2581,N_2911);
and U3769 (N_3769,N_2827,N_2674);
nand U3770 (N_3770,N_2167,N_2028);
nand U3771 (N_3771,N_2389,N_2755);
xnor U3772 (N_3772,N_2767,N_2705);
xor U3773 (N_3773,N_2244,N_2624);
nor U3774 (N_3774,N_2930,N_2859);
or U3775 (N_3775,N_2071,N_2868);
nand U3776 (N_3776,N_2235,N_2569);
nand U3777 (N_3777,N_2742,N_2283);
and U3778 (N_3778,N_2812,N_2763);
and U3779 (N_3779,N_2879,N_2136);
and U3780 (N_3780,N_2651,N_2162);
and U3781 (N_3781,N_2040,N_2549);
and U3782 (N_3782,N_2134,N_2549);
nand U3783 (N_3783,N_2416,N_2454);
or U3784 (N_3784,N_2085,N_2428);
nor U3785 (N_3785,N_2549,N_2004);
or U3786 (N_3786,N_2053,N_2125);
or U3787 (N_3787,N_2211,N_2716);
nor U3788 (N_3788,N_2477,N_2591);
nand U3789 (N_3789,N_2309,N_2005);
nor U3790 (N_3790,N_2029,N_2800);
and U3791 (N_3791,N_2557,N_2496);
nor U3792 (N_3792,N_2644,N_2755);
or U3793 (N_3793,N_2452,N_2190);
xnor U3794 (N_3794,N_2642,N_2607);
and U3795 (N_3795,N_2384,N_2121);
nand U3796 (N_3796,N_2615,N_2620);
or U3797 (N_3797,N_2340,N_2719);
or U3798 (N_3798,N_2180,N_2966);
and U3799 (N_3799,N_2502,N_2509);
and U3800 (N_3800,N_2431,N_2180);
nand U3801 (N_3801,N_2580,N_2241);
and U3802 (N_3802,N_2778,N_2981);
nor U3803 (N_3803,N_2633,N_2689);
xor U3804 (N_3804,N_2684,N_2129);
or U3805 (N_3805,N_2213,N_2785);
or U3806 (N_3806,N_2174,N_2537);
or U3807 (N_3807,N_2884,N_2024);
and U3808 (N_3808,N_2141,N_2092);
or U3809 (N_3809,N_2000,N_2679);
or U3810 (N_3810,N_2461,N_2293);
nor U3811 (N_3811,N_2433,N_2036);
or U3812 (N_3812,N_2395,N_2426);
or U3813 (N_3813,N_2634,N_2175);
nand U3814 (N_3814,N_2903,N_2923);
and U3815 (N_3815,N_2069,N_2986);
and U3816 (N_3816,N_2053,N_2467);
nand U3817 (N_3817,N_2150,N_2594);
nand U3818 (N_3818,N_2787,N_2834);
xor U3819 (N_3819,N_2524,N_2816);
nor U3820 (N_3820,N_2272,N_2971);
and U3821 (N_3821,N_2769,N_2410);
and U3822 (N_3822,N_2508,N_2257);
nand U3823 (N_3823,N_2617,N_2284);
and U3824 (N_3824,N_2820,N_2168);
or U3825 (N_3825,N_2180,N_2247);
nor U3826 (N_3826,N_2552,N_2768);
nor U3827 (N_3827,N_2179,N_2922);
nor U3828 (N_3828,N_2479,N_2379);
nor U3829 (N_3829,N_2732,N_2407);
nand U3830 (N_3830,N_2127,N_2457);
nand U3831 (N_3831,N_2187,N_2540);
nand U3832 (N_3832,N_2644,N_2820);
nor U3833 (N_3833,N_2953,N_2092);
nor U3834 (N_3834,N_2873,N_2540);
or U3835 (N_3835,N_2003,N_2752);
or U3836 (N_3836,N_2076,N_2823);
nor U3837 (N_3837,N_2694,N_2919);
nand U3838 (N_3838,N_2987,N_2117);
and U3839 (N_3839,N_2102,N_2520);
xnor U3840 (N_3840,N_2476,N_2066);
nand U3841 (N_3841,N_2913,N_2609);
nand U3842 (N_3842,N_2203,N_2694);
nor U3843 (N_3843,N_2388,N_2398);
and U3844 (N_3844,N_2356,N_2600);
and U3845 (N_3845,N_2224,N_2872);
or U3846 (N_3846,N_2913,N_2917);
or U3847 (N_3847,N_2760,N_2146);
and U3848 (N_3848,N_2489,N_2349);
nor U3849 (N_3849,N_2419,N_2746);
and U3850 (N_3850,N_2845,N_2659);
nand U3851 (N_3851,N_2429,N_2500);
and U3852 (N_3852,N_2834,N_2323);
nand U3853 (N_3853,N_2736,N_2477);
nand U3854 (N_3854,N_2220,N_2690);
or U3855 (N_3855,N_2915,N_2469);
nand U3856 (N_3856,N_2314,N_2218);
or U3857 (N_3857,N_2821,N_2165);
nand U3858 (N_3858,N_2693,N_2724);
nor U3859 (N_3859,N_2531,N_2675);
or U3860 (N_3860,N_2875,N_2317);
nor U3861 (N_3861,N_2925,N_2196);
and U3862 (N_3862,N_2378,N_2146);
xnor U3863 (N_3863,N_2849,N_2212);
or U3864 (N_3864,N_2605,N_2787);
xnor U3865 (N_3865,N_2707,N_2531);
and U3866 (N_3866,N_2606,N_2504);
and U3867 (N_3867,N_2272,N_2127);
nand U3868 (N_3868,N_2812,N_2218);
nor U3869 (N_3869,N_2266,N_2839);
or U3870 (N_3870,N_2465,N_2472);
and U3871 (N_3871,N_2716,N_2220);
xor U3872 (N_3872,N_2082,N_2108);
and U3873 (N_3873,N_2540,N_2513);
nor U3874 (N_3874,N_2220,N_2167);
nor U3875 (N_3875,N_2094,N_2992);
nor U3876 (N_3876,N_2792,N_2042);
and U3877 (N_3877,N_2141,N_2734);
and U3878 (N_3878,N_2117,N_2326);
and U3879 (N_3879,N_2101,N_2391);
nand U3880 (N_3880,N_2727,N_2434);
nor U3881 (N_3881,N_2084,N_2775);
nor U3882 (N_3882,N_2223,N_2791);
and U3883 (N_3883,N_2629,N_2691);
nor U3884 (N_3884,N_2835,N_2602);
and U3885 (N_3885,N_2606,N_2428);
nor U3886 (N_3886,N_2938,N_2068);
nor U3887 (N_3887,N_2545,N_2817);
or U3888 (N_3888,N_2372,N_2094);
or U3889 (N_3889,N_2674,N_2277);
or U3890 (N_3890,N_2787,N_2937);
nand U3891 (N_3891,N_2678,N_2399);
nor U3892 (N_3892,N_2888,N_2114);
or U3893 (N_3893,N_2389,N_2522);
nand U3894 (N_3894,N_2149,N_2564);
or U3895 (N_3895,N_2718,N_2251);
and U3896 (N_3896,N_2464,N_2281);
nand U3897 (N_3897,N_2671,N_2448);
xnor U3898 (N_3898,N_2164,N_2552);
or U3899 (N_3899,N_2330,N_2630);
nor U3900 (N_3900,N_2676,N_2654);
and U3901 (N_3901,N_2268,N_2392);
or U3902 (N_3902,N_2264,N_2267);
and U3903 (N_3903,N_2437,N_2174);
nand U3904 (N_3904,N_2450,N_2000);
nor U3905 (N_3905,N_2342,N_2005);
and U3906 (N_3906,N_2356,N_2258);
nand U3907 (N_3907,N_2556,N_2245);
or U3908 (N_3908,N_2005,N_2297);
nor U3909 (N_3909,N_2566,N_2812);
nand U3910 (N_3910,N_2785,N_2118);
and U3911 (N_3911,N_2230,N_2314);
or U3912 (N_3912,N_2480,N_2763);
or U3913 (N_3913,N_2032,N_2787);
or U3914 (N_3914,N_2894,N_2626);
nand U3915 (N_3915,N_2671,N_2328);
or U3916 (N_3916,N_2084,N_2700);
or U3917 (N_3917,N_2641,N_2143);
or U3918 (N_3918,N_2163,N_2588);
nor U3919 (N_3919,N_2539,N_2995);
xnor U3920 (N_3920,N_2152,N_2417);
or U3921 (N_3921,N_2594,N_2454);
nor U3922 (N_3922,N_2762,N_2912);
nor U3923 (N_3923,N_2878,N_2992);
and U3924 (N_3924,N_2342,N_2424);
nand U3925 (N_3925,N_2230,N_2596);
nand U3926 (N_3926,N_2003,N_2823);
and U3927 (N_3927,N_2869,N_2622);
or U3928 (N_3928,N_2099,N_2436);
nor U3929 (N_3929,N_2156,N_2730);
nand U3930 (N_3930,N_2324,N_2243);
nand U3931 (N_3931,N_2132,N_2833);
or U3932 (N_3932,N_2812,N_2352);
xor U3933 (N_3933,N_2670,N_2305);
nor U3934 (N_3934,N_2272,N_2111);
nand U3935 (N_3935,N_2268,N_2731);
or U3936 (N_3936,N_2745,N_2012);
nand U3937 (N_3937,N_2966,N_2006);
nand U3938 (N_3938,N_2569,N_2589);
nor U3939 (N_3939,N_2778,N_2863);
nor U3940 (N_3940,N_2657,N_2031);
or U3941 (N_3941,N_2867,N_2566);
or U3942 (N_3942,N_2381,N_2652);
nor U3943 (N_3943,N_2633,N_2510);
nand U3944 (N_3944,N_2737,N_2383);
and U3945 (N_3945,N_2931,N_2175);
and U3946 (N_3946,N_2657,N_2306);
nand U3947 (N_3947,N_2463,N_2625);
nor U3948 (N_3948,N_2071,N_2985);
or U3949 (N_3949,N_2724,N_2594);
nor U3950 (N_3950,N_2064,N_2721);
nor U3951 (N_3951,N_2569,N_2779);
or U3952 (N_3952,N_2046,N_2407);
or U3953 (N_3953,N_2258,N_2047);
xnor U3954 (N_3954,N_2232,N_2488);
and U3955 (N_3955,N_2695,N_2191);
xnor U3956 (N_3956,N_2436,N_2293);
or U3957 (N_3957,N_2444,N_2574);
nor U3958 (N_3958,N_2037,N_2173);
or U3959 (N_3959,N_2932,N_2694);
or U3960 (N_3960,N_2649,N_2578);
and U3961 (N_3961,N_2032,N_2940);
or U3962 (N_3962,N_2171,N_2178);
nor U3963 (N_3963,N_2610,N_2727);
nor U3964 (N_3964,N_2502,N_2192);
nand U3965 (N_3965,N_2650,N_2323);
nor U3966 (N_3966,N_2351,N_2118);
xor U3967 (N_3967,N_2914,N_2690);
nand U3968 (N_3968,N_2492,N_2033);
and U3969 (N_3969,N_2291,N_2064);
and U3970 (N_3970,N_2917,N_2131);
nand U3971 (N_3971,N_2569,N_2138);
nor U3972 (N_3972,N_2171,N_2771);
nor U3973 (N_3973,N_2869,N_2349);
nor U3974 (N_3974,N_2097,N_2274);
or U3975 (N_3975,N_2153,N_2365);
and U3976 (N_3976,N_2003,N_2386);
and U3977 (N_3977,N_2851,N_2289);
nor U3978 (N_3978,N_2043,N_2824);
or U3979 (N_3979,N_2914,N_2262);
and U3980 (N_3980,N_2718,N_2309);
or U3981 (N_3981,N_2288,N_2954);
nand U3982 (N_3982,N_2937,N_2607);
nor U3983 (N_3983,N_2725,N_2977);
xnor U3984 (N_3984,N_2608,N_2775);
xor U3985 (N_3985,N_2428,N_2508);
or U3986 (N_3986,N_2439,N_2711);
or U3987 (N_3987,N_2329,N_2538);
and U3988 (N_3988,N_2383,N_2050);
nor U3989 (N_3989,N_2199,N_2990);
or U3990 (N_3990,N_2401,N_2171);
or U3991 (N_3991,N_2055,N_2477);
and U3992 (N_3992,N_2445,N_2028);
or U3993 (N_3993,N_2039,N_2933);
and U3994 (N_3994,N_2684,N_2078);
nand U3995 (N_3995,N_2952,N_2853);
nand U3996 (N_3996,N_2890,N_2595);
nand U3997 (N_3997,N_2350,N_2797);
nand U3998 (N_3998,N_2190,N_2163);
xnor U3999 (N_3999,N_2860,N_2589);
and U4000 (N_4000,N_3864,N_3525);
xnor U4001 (N_4001,N_3298,N_3980);
xor U4002 (N_4002,N_3183,N_3404);
xor U4003 (N_4003,N_3444,N_3038);
nor U4004 (N_4004,N_3308,N_3415);
nor U4005 (N_4005,N_3324,N_3730);
nand U4006 (N_4006,N_3982,N_3316);
and U4007 (N_4007,N_3584,N_3725);
nor U4008 (N_4008,N_3609,N_3485);
or U4009 (N_4009,N_3332,N_3520);
and U4010 (N_4010,N_3411,N_3868);
or U4011 (N_4011,N_3860,N_3495);
and U4012 (N_4012,N_3877,N_3243);
and U4013 (N_4013,N_3438,N_3381);
nand U4014 (N_4014,N_3744,N_3664);
nand U4015 (N_4015,N_3244,N_3674);
nand U4016 (N_4016,N_3505,N_3733);
nand U4017 (N_4017,N_3513,N_3543);
xnor U4018 (N_4018,N_3201,N_3550);
or U4019 (N_4019,N_3228,N_3130);
nand U4020 (N_4020,N_3254,N_3140);
nand U4021 (N_4021,N_3061,N_3171);
and U4022 (N_4022,N_3820,N_3494);
xor U4023 (N_4023,N_3185,N_3343);
nor U4024 (N_4024,N_3242,N_3050);
xnor U4025 (N_4025,N_3181,N_3263);
and U4026 (N_4026,N_3591,N_3321);
xor U4027 (N_4027,N_3335,N_3680);
nor U4028 (N_4028,N_3429,N_3519);
nor U4029 (N_4029,N_3743,N_3153);
or U4030 (N_4030,N_3663,N_3803);
nand U4031 (N_4031,N_3333,N_3425);
or U4032 (N_4032,N_3292,N_3043);
nor U4033 (N_4033,N_3857,N_3068);
nor U4034 (N_4034,N_3622,N_3654);
nand U4035 (N_4035,N_3675,N_3987);
and U4036 (N_4036,N_3122,N_3363);
nand U4037 (N_4037,N_3096,N_3671);
nor U4038 (N_4038,N_3349,N_3439);
or U4039 (N_4039,N_3512,N_3095);
or U4040 (N_4040,N_3466,N_3001);
or U4041 (N_4041,N_3112,N_3356);
nand U4042 (N_4042,N_3277,N_3510);
and U4043 (N_4043,N_3738,N_3881);
nor U4044 (N_4044,N_3880,N_3399);
nand U4045 (N_4045,N_3607,N_3567);
or U4046 (N_4046,N_3736,N_3257);
nor U4047 (N_4047,N_3037,N_3156);
and U4048 (N_4048,N_3986,N_3045);
nand U4049 (N_4049,N_3119,N_3817);
nand U4050 (N_4050,N_3295,N_3370);
or U4051 (N_4051,N_3081,N_3933);
or U4052 (N_4052,N_3760,N_3943);
and U4053 (N_4053,N_3827,N_3233);
or U4054 (N_4054,N_3237,N_3960);
nor U4055 (N_4055,N_3871,N_3692);
xor U4056 (N_4056,N_3268,N_3280);
and U4057 (N_4057,N_3379,N_3687);
nor U4058 (N_4058,N_3284,N_3646);
and U4059 (N_4059,N_3831,N_3899);
nor U4060 (N_4060,N_3144,N_3142);
and U4061 (N_4061,N_3287,N_3666);
or U4062 (N_4062,N_3884,N_3883);
and U4063 (N_4063,N_3610,N_3615);
and U4064 (N_4064,N_3063,N_3057);
xnor U4065 (N_4065,N_3524,N_3407);
or U4066 (N_4066,N_3894,N_3891);
nor U4067 (N_4067,N_3464,N_3098);
nor U4068 (N_4068,N_3107,N_3976);
and U4069 (N_4069,N_3361,N_3120);
xnor U4070 (N_4070,N_3317,N_3949);
nor U4071 (N_4071,N_3561,N_3583);
xor U4072 (N_4072,N_3420,N_3431);
and U4073 (N_4073,N_3806,N_3282);
and U4074 (N_4074,N_3461,N_3252);
nor U4075 (N_4075,N_3897,N_3065);
nand U4076 (N_4076,N_3636,N_3970);
nor U4077 (N_4077,N_3443,N_3025);
nor U4078 (N_4078,N_3787,N_3851);
nand U4079 (N_4079,N_3329,N_3101);
or U4080 (N_4080,N_3470,N_3482);
nand U4081 (N_4081,N_3704,N_3442);
nor U4082 (N_4082,N_3269,N_3149);
or U4083 (N_4083,N_3934,N_3367);
and U4084 (N_4084,N_3087,N_3216);
nor U4085 (N_4085,N_3385,N_3350);
and U4086 (N_4086,N_3932,N_3441);
or U4087 (N_4087,N_3376,N_3916);
nand U4088 (N_4088,N_3785,N_3476);
and U4089 (N_4089,N_3781,N_3498);
or U4090 (N_4090,N_3977,N_3716);
nor U4091 (N_4091,N_3215,N_3239);
nand U4092 (N_4092,N_3380,N_3993);
and U4093 (N_4093,N_3283,N_3508);
nor U4094 (N_4094,N_3305,N_3995);
xor U4095 (N_4095,N_3875,N_3223);
nor U4096 (N_4096,N_3770,N_3265);
or U4097 (N_4097,N_3445,N_3746);
nand U4098 (N_4098,N_3768,N_3569);
xnor U4099 (N_4099,N_3759,N_3762);
or U4100 (N_4100,N_3289,N_3401);
and U4101 (N_4101,N_3889,N_3752);
nand U4102 (N_4102,N_3334,N_3196);
nor U4103 (N_4103,N_3849,N_3089);
or U4104 (N_4104,N_3163,N_3413);
or U4105 (N_4105,N_3603,N_3031);
or U4106 (N_4106,N_3858,N_3491);
nor U4107 (N_4107,N_3094,N_3565);
nand U4108 (N_4108,N_3867,N_3225);
xor U4109 (N_4109,N_3967,N_3108);
nor U4110 (N_4110,N_3896,N_3805);
and U4111 (N_4111,N_3330,N_3191);
xnor U4112 (N_4112,N_3132,N_3497);
or U4113 (N_4113,N_3850,N_3104);
nor U4114 (N_4114,N_3926,N_3903);
and U4115 (N_4115,N_3146,N_3170);
nand U4116 (N_4116,N_3285,N_3209);
or U4117 (N_4117,N_3058,N_3315);
xor U4118 (N_4118,N_3255,N_3137);
nand U4119 (N_4119,N_3428,N_3595);
and U4120 (N_4120,N_3016,N_3804);
and U4121 (N_4121,N_3055,N_3973);
or U4122 (N_4122,N_3323,N_3007);
and U4123 (N_4123,N_3410,N_3500);
and U4124 (N_4124,N_3518,N_3408);
nand U4125 (N_4125,N_3168,N_3328);
nor U4126 (N_4126,N_3172,N_3480);
nand U4127 (N_4127,N_3731,N_3521);
nand U4128 (N_4128,N_3802,N_3366);
or U4129 (N_4129,N_3048,N_3763);
and U4130 (N_4130,N_3021,N_3325);
or U4131 (N_4131,N_3433,N_3530);
and U4132 (N_4132,N_3258,N_3248);
nand U4133 (N_4133,N_3430,N_3227);
xor U4134 (N_4134,N_3378,N_3475);
nand U4135 (N_4135,N_3639,N_3296);
nor U4136 (N_4136,N_3865,N_3992);
or U4137 (N_4137,N_3117,N_3126);
nor U4138 (N_4138,N_3737,N_3272);
or U4139 (N_4139,N_3651,N_3083);
and U4140 (N_4140,N_3326,N_3758);
nor U4141 (N_4141,N_3229,N_3649);
or U4142 (N_4142,N_3162,N_3199);
or U4143 (N_4143,N_3092,N_3869);
nand U4144 (N_4144,N_3592,N_3022);
nor U4145 (N_4145,N_3909,N_3054);
and U4146 (N_4146,N_3791,N_3825);
xor U4147 (N_4147,N_3003,N_3091);
nor U4148 (N_4148,N_3790,N_3940);
or U4149 (N_4149,N_3202,N_3560);
or U4150 (N_4150,N_3256,N_3632);
nor U4151 (N_4151,N_3585,N_3541);
nand U4152 (N_4152,N_3432,N_3630);
nand U4153 (N_4153,N_3732,N_3895);
nand U4154 (N_4154,N_3637,N_3856);
nor U4155 (N_4155,N_3965,N_3211);
xnor U4156 (N_4156,N_3067,N_3559);
or U4157 (N_4157,N_3734,N_3337);
nand U4158 (N_4158,N_3971,N_3205);
or U4159 (N_4159,N_3206,N_3693);
nand U4160 (N_4160,N_3611,N_3576);
or U4161 (N_4161,N_3819,N_3138);
nand U4162 (N_4162,N_3571,N_3617);
or U4163 (N_4163,N_3383,N_3810);
xnor U4164 (N_4164,N_3157,N_3818);
xnor U4165 (N_4165,N_3952,N_3673);
nand U4166 (N_4166,N_3241,N_3417);
nand U4167 (N_4167,N_3957,N_3483);
nor U4168 (N_4168,N_3536,N_3253);
nor U4169 (N_4169,N_3826,N_3465);
and U4170 (N_4170,N_3918,N_3930);
or U4171 (N_4171,N_3879,N_3658);
nand U4172 (N_4172,N_3474,N_3745);
xnor U4173 (N_4173,N_3062,N_3691);
nor U4174 (N_4174,N_3783,N_3319);
or U4175 (N_4175,N_3580,N_3177);
and U4176 (N_4176,N_3531,N_3369);
nor U4177 (N_4177,N_3772,N_3188);
nor U4178 (N_4178,N_3460,N_3719);
nand U4179 (N_4179,N_3700,N_3042);
xnor U4180 (N_4180,N_3017,N_3566);
nor U4181 (N_4181,N_3102,N_3391);
nor U4182 (N_4182,N_3564,N_3027);
or U4183 (N_4183,N_3780,N_3346);
and U4184 (N_4184,N_3695,N_3833);
nand U4185 (N_4185,N_3948,N_3912);
and U4186 (N_4186,N_3070,N_3481);
or U4187 (N_4187,N_3714,N_3900);
or U4188 (N_4188,N_3661,N_3240);
nor U4189 (N_4189,N_3558,N_3997);
nor U4190 (N_4190,N_3813,N_3080);
nand U4191 (N_4191,N_3046,N_3060);
nor U4192 (N_4192,N_3488,N_3499);
nand U4193 (N_4193,N_3423,N_3890);
xor U4194 (N_4194,N_3862,N_3832);
and U4195 (N_4195,N_3589,N_3047);
nor U4196 (N_4196,N_3836,N_3626);
nor U4197 (N_4197,N_3553,N_3472);
and U4198 (N_4198,N_3484,N_3886);
or U4199 (N_4199,N_3621,N_3917);
xor U4200 (N_4200,N_3642,N_3271);
nand U4201 (N_4201,N_3400,N_3434);
nor U4202 (N_4202,N_3563,N_3882);
and U4203 (N_4203,N_3000,N_3338);
nand U4204 (N_4204,N_3793,N_3808);
nor U4205 (N_4205,N_3624,N_3638);
nor U4206 (N_4206,N_3118,N_3774);
or U4207 (N_4207,N_3712,N_3134);
nand U4208 (N_4208,N_3812,N_3677);
and U4209 (N_4209,N_3606,N_3978);
nand U4210 (N_4210,N_3573,N_3359);
nand U4211 (N_4211,N_3164,N_3694);
or U4212 (N_4212,N_3623,N_3984);
nand U4213 (N_4213,N_3852,N_3259);
or U4214 (N_4214,N_3174,N_3371);
or U4215 (N_4215,N_3801,N_3396);
or U4216 (N_4216,N_3554,N_3535);
nand U4217 (N_4217,N_3028,N_3222);
or U4218 (N_4218,N_3347,N_3260);
nand U4219 (N_4219,N_3778,N_3750);
or U4220 (N_4220,N_3656,N_3516);
nor U4221 (N_4221,N_3853,N_3866);
or U4222 (N_4222,N_3150,N_3275);
nor U4223 (N_4223,N_3005,N_3526);
and U4224 (N_4224,N_3468,N_3436);
or U4225 (N_4225,N_3711,N_3614);
nand U4226 (N_4226,N_3198,N_3190);
xnor U4227 (N_4227,N_3990,N_3924);
and U4228 (N_4228,N_3527,N_3686);
and U4229 (N_4229,N_3395,N_3684);
nand U4230 (N_4230,N_3556,N_3032);
xor U4231 (N_4231,N_3139,N_3915);
nor U4232 (N_4232,N_3601,N_3155);
nand U4233 (N_4233,N_3872,N_3794);
or U4234 (N_4234,N_3988,N_3653);
or U4235 (N_4235,N_3847,N_3771);
or U4236 (N_4236,N_3898,N_3800);
and U4237 (N_4237,N_3085,N_3023);
and U4238 (N_4238,N_3471,N_3299);
or U4239 (N_4239,N_3451,N_3235);
and U4240 (N_4240,N_3368,N_3220);
or U4241 (N_4241,N_3715,N_3504);
nand U4242 (N_4242,N_3578,N_3297);
nand U4243 (N_4243,N_3302,N_3914);
nor U4244 (N_4244,N_3148,N_3355);
xor U4245 (N_4245,N_3238,N_3477);
or U4246 (N_4246,N_3014,N_3892);
xnor U4247 (N_4247,N_3147,N_3964);
or U4248 (N_4248,N_3840,N_3697);
xnor U4249 (N_4249,N_3403,N_3035);
nor U4250 (N_4250,N_3983,N_3821);
or U4251 (N_4251,N_3384,N_3717);
or U4252 (N_4252,N_3136,N_3309);
nor U4253 (N_4253,N_3887,N_3278);
xnor U4254 (N_4254,N_3718,N_3077);
and U4255 (N_4255,N_3469,N_3208);
or U4256 (N_4256,N_3293,N_3811);
xor U4257 (N_4257,N_3307,N_3904);
nand U4258 (N_4258,N_3757,N_3449);
and U4259 (N_4259,N_3360,N_3902);
xor U4260 (N_4260,N_3416,N_3270);
or U4261 (N_4261,N_3194,N_3019);
or U4262 (N_4262,N_3975,N_3339);
and U4263 (N_4263,N_3870,N_3012);
or U4264 (N_4264,N_3944,N_3179);
or U4265 (N_4265,N_3074,N_3753);
nand U4266 (N_4266,N_3006,N_3125);
nand U4267 (N_4267,N_3294,N_3863);
nand U4268 (N_4268,N_3121,N_3453);
and U4269 (N_4269,N_3231,N_3931);
or U4270 (N_4270,N_3795,N_3458);
nor U4271 (N_4271,N_3596,N_3486);
nand U4272 (N_4272,N_3167,N_3358);
and U4273 (N_4273,N_3577,N_3688);
nand U4274 (N_4274,N_3537,N_3011);
xor U4275 (N_4275,N_3600,N_3764);
nand U4276 (N_4276,N_3645,N_3389);
or U4277 (N_4277,N_3854,N_3503);
or U4278 (N_4278,N_3180,N_3552);
and U4279 (N_4279,N_3546,N_3088);
or U4280 (N_4280,N_3246,N_3217);
or U4281 (N_4281,N_3459,N_3901);
nor U4282 (N_4282,N_3311,N_3873);
nor U4283 (N_4283,N_3581,N_3844);
or U4284 (N_4284,N_3648,N_3517);
and U4285 (N_4285,N_3398,N_3212);
nand U4286 (N_4286,N_3816,N_3955);
xnor U4287 (N_4287,N_3506,N_3075);
nand U4288 (N_4288,N_3099,N_3644);
or U4289 (N_4289,N_3158,N_3628);
nand U4290 (N_4290,N_3701,N_3665);
nand U4291 (N_4291,N_3418,N_3913);
nor U4292 (N_4292,N_3613,N_3008);
and U4293 (N_4293,N_3002,N_3925);
xnor U4294 (N_4294,N_3799,N_3713);
and U4295 (N_4295,N_3775,N_3114);
nand U4296 (N_4296,N_3619,N_3348);
and U4297 (N_4297,N_3655,N_3166);
nand U4298 (N_4298,N_3123,N_3928);
or U4299 (N_4299,N_3030,N_3448);
nor U4300 (N_4300,N_3274,N_3652);
and U4301 (N_4301,N_3250,N_3698);
nor U4302 (N_4302,N_3026,N_3093);
xor U4303 (N_4303,N_3921,N_3226);
xor U4304 (N_4304,N_3210,N_3127);
xnor U4305 (N_4305,N_3557,N_3203);
and U4306 (N_4306,N_3236,N_3039);
and U4307 (N_4307,N_3247,N_3455);
nor U4308 (N_4308,N_3570,N_3186);
and U4309 (N_4309,N_3245,N_3192);
nand U4310 (N_4310,N_3009,N_3421);
nand U4311 (N_4311,N_3195,N_3962);
xnor U4312 (N_4312,N_3105,N_3357);
nor U4313 (N_4313,N_3702,N_3534);
and U4314 (N_4314,N_3013,N_3078);
nand U4315 (N_4315,N_3354,N_3669);
nand U4316 (N_4316,N_3647,N_3662);
and U4317 (N_4317,N_3788,N_3549);
and U4318 (N_4318,N_3532,N_3066);
nor U4319 (N_4319,N_3815,N_3740);
nand U4320 (N_4320,N_3100,N_3888);
and U4321 (N_4321,N_3659,N_3842);
and U4322 (N_4322,N_3773,N_3910);
nor U4323 (N_4323,N_3073,N_3291);
xnor U4324 (N_4324,N_3273,N_3193);
and U4325 (N_4325,N_3056,N_3705);
xnor U4326 (N_4326,N_3739,N_3036);
or U4327 (N_4327,N_3594,N_3160);
nand U4328 (N_4328,N_3044,N_3232);
nand U4329 (N_4329,N_3598,N_3103);
xnor U4330 (N_4330,N_3985,N_3110);
and U4331 (N_4331,N_3279,N_3414);
xor U4332 (N_4332,N_3843,N_3447);
nand U4333 (N_4333,N_3789,N_3939);
nor U4334 (N_4334,N_3069,N_3207);
nor U4335 (N_4335,N_3462,N_3841);
or U4336 (N_4336,N_3735,N_3511);
nor U4337 (N_4337,N_3076,N_3784);
or U4338 (N_4338,N_3911,N_3681);
and U4339 (N_4339,N_3457,N_3397);
nand U4340 (N_4340,N_3386,N_3523);
or U4341 (N_4341,N_3189,N_3450);
or U4342 (N_4342,N_3345,N_3135);
or U4343 (N_4343,N_3479,N_3290);
nor U4344 (N_4344,N_3961,N_3742);
and U4345 (N_4345,N_3582,N_3084);
or U4346 (N_4346,N_3452,N_3187);
nor U4347 (N_4347,N_3015,N_3922);
nor U4348 (N_4348,N_3340,N_3051);
and U4349 (N_4349,N_3830,N_3766);
or U4350 (N_4350,N_3824,N_3777);
nor U4351 (N_4351,N_3956,N_3456);
nor U4352 (N_4352,N_3489,N_3204);
nor U4353 (N_4353,N_3641,N_3169);
nor U4354 (N_4354,N_3959,N_3353);
nor U4355 (N_4355,N_3551,N_3446);
or U4356 (N_4356,N_3562,N_3539);
nor U4357 (N_4357,N_3176,N_3721);
xnor U4358 (N_4358,N_3676,N_3572);
and U4359 (N_4359,N_3786,N_3848);
xnor U4360 (N_4360,N_3540,N_3767);
nor U4361 (N_4361,N_3129,N_3152);
nor U4362 (N_4362,N_3953,N_3575);
xnor U4363 (N_4363,N_3966,N_3927);
and U4364 (N_4364,N_3998,N_3286);
nor U4365 (N_4365,N_3667,N_3920);
xor U4366 (N_4366,N_3951,N_3728);
nor U4367 (N_4367,N_3942,N_3234);
nand U4368 (N_4368,N_3706,N_3547);
nor U4369 (N_4369,N_3709,N_3175);
nand U4370 (N_4370,N_3586,N_3529);
nor U4371 (N_4371,N_3544,N_3463);
nand U4372 (N_4372,N_3336,N_3538);
nand U4373 (N_4373,N_3392,N_3839);
nor U4374 (N_4374,N_3427,N_3300);
nor U4375 (N_4375,N_3616,N_3221);
nor U4376 (N_4376,N_3230,N_3929);
nor U4377 (N_4377,N_3679,N_3116);
nor U4378 (N_4378,N_3327,N_3478);
xor U4379 (N_4379,N_3024,N_3635);
and U4380 (N_4380,N_3249,N_3542);
nand U4381 (N_4381,N_3859,N_3672);
or U4382 (N_4382,N_3304,N_3969);
nor U4383 (N_4383,N_3612,N_3440);
nand U4384 (N_4384,N_3905,N_3593);
or U4385 (N_4385,N_3200,N_3004);
or U4386 (N_4386,N_3958,N_3052);
nor U4387 (N_4387,N_3267,N_3141);
nor U4388 (N_4388,N_3303,N_3722);
xor U4389 (N_4389,N_3729,N_3133);
or U4390 (N_4390,N_3310,N_3143);
nand U4391 (N_4391,N_3213,N_3588);
and U4392 (N_4392,N_3314,N_3590);
nand U4393 (N_4393,N_3769,N_3487);
nor U4394 (N_4394,N_3473,N_3341);
and U4395 (N_4395,N_3604,N_3782);
nor U4396 (N_4396,N_3322,N_3393);
nand U4397 (N_4397,N_3251,N_3660);
nor U4398 (N_4398,N_3422,N_3545);
or U4399 (N_4399,N_3765,N_3587);
nor U4400 (N_4400,N_3219,N_3747);
and U4401 (N_4401,N_3097,N_3184);
and U4402 (N_4402,N_3128,N_3419);
xor U4403 (N_4403,N_3318,N_3115);
or U4404 (N_4404,N_3979,N_3726);
xor U4405 (N_4405,N_3568,N_3972);
and U4406 (N_4406,N_3375,N_3344);
nand U4407 (N_4407,N_3707,N_3878);
nor U4408 (N_4408,N_3390,N_3165);
nand U4409 (N_4409,N_3741,N_3426);
and U4410 (N_4410,N_3937,N_3829);
nor U4411 (N_4411,N_3313,N_3796);
nand U4412 (N_4412,N_3838,N_3145);
nand U4413 (N_4413,N_3634,N_3845);
or U4414 (N_4414,N_3352,N_3938);
nand U4415 (N_4415,N_3424,N_3608);
and U4416 (N_4416,N_3364,N_3668);
or U4417 (N_4417,N_3331,N_3779);
nor U4418 (N_4418,N_3797,N_3111);
nand U4419 (N_4419,N_3320,N_3749);
and U4420 (N_4420,N_3161,N_3633);
nand U4421 (N_4421,N_3574,N_3690);
nand U4422 (N_4422,N_3224,N_3454);
or U4423 (N_4423,N_3823,N_3412);
or U4424 (N_4424,N_3072,N_3034);
nor U4425 (N_4425,N_3994,N_3919);
and U4426 (N_4426,N_3281,N_3082);
nand U4427 (N_4427,N_3492,N_3178);
or U4428 (N_4428,N_3776,N_3602);
nand U4429 (N_4429,N_3493,N_3515);
nor U4430 (N_4430,N_3053,N_3533);
nand U4431 (N_4431,N_3388,N_3079);
xnor U4432 (N_4432,N_3113,N_3124);
nand U4433 (N_4433,N_3723,N_3214);
nand U4434 (N_4434,N_3620,N_3159);
and U4435 (N_4435,N_3792,N_3382);
nand U4436 (N_4436,N_3755,N_3814);
nand U4437 (N_4437,N_3276,N_3040);
or U4438 (N_4438,N_3683,N_3991);
nor U4439 (N_4439,N_3131,N_3365);
and U4440 (N_4440,N_3861,N_3650);
nand U4441 (N_4441,N_3059,N_3514);
and U4442 (N_4442,N_3855,N_3874);
nand U4443 (N_4443,N_3018,N_3923);
and U4444 (N_4444,N_3387,N_3885);
nand U4445 (N_4445,N_3710,N_3947);
or U4446 (N_4446,N_3809,N_3631);
and U4447 (N_4447,N_3798,N_3682);
and U4448 (N_4448,N_3989,N_3968);
nand U4449 (N_4449,N_3437,N_3696);
nand U4450 (N_4450,N_3579,N_3312);
nand U4451 (N_4451,N_3724,N_3509);
nand U4452 (N_4452,N_3467,N_3751);
nand U4453 (N_4453,N_3893,N_3049);
or U4454 (N_4454,N_3756,N_3605);
nor U4455 (N_4455,N_3218,N_3406);
or U4456 (N_4456,N_3377,N_3678);
nand U4457 (N_4457,N_3996,N_3748);
nor U4458 (N_4458,N_3109,N_3699);
nand U4459 (N_4459,N_3936,N_3496);
xor U4460 (N_4460,N_3490,N_3086);
and U4461 (N_4461,N_3981,N_3727);
xor U4462 (N_4462,N_3033,N_3154);
and U4463 (N_4463,N_3941,N_3950);
or U4464 (N_4464,N_3618,N_3522);
and U4465 (N_4465,N_3703,N_3197);
nand U4466 (N_4466,N_3071,N_3708);
and U4467 (N_4467,N_3528,N_3182);
nand U4468 (N_4468,N_3640,N_3945);
nor U4469 (N_4469,N_3908,N_3974);
or U4470 (N_4470,N_3627,N_3846);
and U4471 (N_4471,N_3507,N_3362);
and U4472 (N_4472,N_3090,N_3963);
nor U4473 (N_4473,N_3288,N_3548);
nand U4474 (N_4474,N_3834,N_3264);
nor U4475 (N_4475,N_3754,N_3837);
nand U4476 (N_4476,N_3685,N_3689);
nand U4477 (N_4477,N_3262,N_3010);
and U4478 (N_4478,N_3501,N_3405);
or U4479 (N_4479,N_3435,N_3402);
nand U4480 (N_4480,N_3409,N_3629);
and U4481 (N_4481,N_3173,N_3064);
or U4482 (N_4482,N_3807,N_3372);
xnor U4483 (N_4483,N_3351,N_3041);
and U4484 (N_4484,N_3029,N_3822);
nand U4485 (N_4485,N_3625,N_3954);
or U4486 (N_4486,N_3373,N_3907);
and U4487 (N_4487,N_3670,N_3597);
or U4488 (N_4488,N_3876,N_3720);
nor U4489 (N_4489,N_3761,N_3106);
or U4490 (N_4490,N_3835,N_3306);
or U4491 (N_4491,N_3266,N_3946);
nand U4492 (N_4492,N_3301,N_3906);
xor U4493 (N_4493,N_3657,N_3935);
or U4494 (N_4494,N_3342,N_3261);
or U4495 (N_4495,N_3828,N_3394);
nand U4496 (N_4496,N_3999,N_3151);
or U4497 (N_4497,N_3599,N_3643);
nor U4498 (N_4498,N_3555,N_3374);
or U4499 (N_4499,N_3020,N_3502);
or U4500 (N_4500,N_3331,N_3254);
nor U4501 (N_4501,N_3561,N_3250);
xor U4502 (N_4502,N_3743,N_3887);
nand U4503 (N_4503,N_3767,N_3979);
or U4504 (N_4504,N_3009,N_3724);
or U4505 (N_4505,N_3779,N_3854);
nand U4506 (N_4506,N_3167,N_3864);
and U4507 (N_4507,N_3938,N_3402);
or U4508 (N_4508,N_3312,N_3853);
nand U4509 (N_4509,N_3729,N_3628);
nand U4510 (N_4510,N_3933,N_3715);
nor U4511 (N_4511,N_3496,N_3863);
and U4512 (N_4512,N_3467,N_3794);
nand U4513 (N_4513,N_3037,N_3900);
xor U4514 (N_4514,N_3385,N_3941);
and U4515 (N_4515,N_3477,N_3321);
xor U4516 (N_4516,N_3631,N_3165);
nor U4517 (N_4517,N_3443,N_3173);
and U4518 (N_4518,N_3180,N_3495);
nor U4519 (N_4519,N_3810,N_3581);
nor U4520 (N_4520,N_3588,N_3828);
nand U4521 (N_4521,N_3475,N_3520);
and U4522 (N_4522,N_3135,N_3402);
or U4523 (N_4523,N_3338,N_3527);
xor U4524 (N_4524,N_3482,N_3758);
or U4525 (N_4525,N_3168,N_3439);
or U4526 (N_4526,N_3474,N_3542);
and U4527 (N_4527,N_3348,N_3423);
and U4528 (N_4528,N_3635,N_3403);
and U4529 (N_4529,N_3247,N_3477);
nand U4530 (N_4530,N_3978,N_3538);
nand U4531 (N_4531,N_3535,N_3889);
and U4532 (N_4532,N_3184,N_3276);
and U4533 (N_4533,N_3911,N_3878);
nand U4534 (N_4534,N_3182,N_3264);
nand U4535 (N_4535,N_3078,N_3649);
nand U4536 (N_4536,N_3921,N_3551);
nor U4537 (N_4537,N_3958,N_3740);
nor U4538 (N_4538,N_3777,N_3112);
nand U4539 (N_4539,N_3559,N_3473);
or U4540 (N_4540,N_3554,N_3809);
nor U4541 (N_4541,N_3595,N_3612);
xnor U4542 (N_4542,N_3497,N_3133);
and U4543 (N_4543,N_3344,N_3844);
nand U4544 (N_4544,N_3507,N_3987);
xor U4545 (N_4545,N_3200,N_3021);
nand U4546 (N_4546,N_3253,N_3405);
or U4547 (N_4547,N_3669,N_3487);
nand U4548 (N_4548,N_3931,N_3400);
or U4549 (N_4549,N_3276,N_3278);
or U4550 (N_4550,N_3495,N_3807);
and U4551 (N_4551,N_3598,N_3301);
and U4552 (N_4552,N_3248,N_3283);
nor U4553 (N_4553,N_3920,N_3441);
and U4554 (N_4554,N_3993,N_3593);
nand U4555 (N_4555,N_3955,N_3996);
nand U4556 (N_4556,N_3852,N_3144);
and U4557 (N_4557,N_3125,N_3482);
nand U4558 (N_4558,N_3559,N_3199);
nor U4559 (N_4559,N_3011,N_3694);
and U4560 (N_4560,N_3408,N_3015);
or U4561 (N_4561,N_3279,N_3327);
nand U4562 (N_4562,N_3062,N_3141);
nor U4563 (N_4563,N_3102,N_3553);
or U4564 (N_4564,N_3873,N_3738);
xor U4565 (N_4565,N_3393,N_3054);
and U4566 (N_4566,N_3550,N_3235);
nor U4567 (N_4567,N_3869,N_3155);
nand U4568 (N_4568,N_3266,N_3909);
and U4569 (N_4569,N_3016,N_3092);
and U4570 (N_4570,N_3105,N_3304);
nand U4571 (N_4571,N_3433,N_3329);
xor U4572 (N_4572,N_3242,N_3134);
nand U4573 (N_4573,N_3680,N_3017);
nor U4574 (N_4574,N_3202,N_3435);
or U4575 (N_4575,N_3436,N_3845);
and U4576 (N_4576,N_3044,N_3926);
xor U4577 (N_4577,N_3041,N_3834);
and U4578 (N_4578,N_3674,N_3361);
or U4579 (N_4579,N_3982,N_3061);
and U4580 (N_4580,N_3880,N_3509);
xor U4581 (N_4581,N_3563,N_3082);
nand U4582 (N_4582,N_3965,N_3347);
nand U4583 (N_4583,N_3753,N_3788);
or U4584 (N_4584,N_3198,N_3669);
nand U4585 (N_4585,N_3896,N_3412);
nor U4586 (N_4586,N_3675,N_3451);
nand U4587 (N_4587,N_3706,N_3804);
xnor U4588 (N_4588,N_3935,N_3045);
nand U4589 (N_4589,N_3861,N_3263);
and U4590 (N_4590,N_3365,N_3495);
nand U4591 (N_4591,N_3454,N_3046);
or U4592 (N_4592,N_3465,N_3671);
nor U4593 (N_4593,N_3267,N_3082);
and U4594 (N_4594,N_3503,N_3703);
nor U4595 (N_4595,N_3301,N_3953);
or U4596 (N_4596,N_3668,N_3940);
xnor U4597 (N_4597,N_3939,N_3852);
or U4598 (N_4598,N_3185,N_3238);
nor U4599 (N_4599,N_3249,N_3936);
nand U4600 (N_4600,N_3021,N_3192);
and U4601 (N_4601,N_3674,N_3604);
nor U4602 (N_4602,N_3108,N_3394);
or U4603 (N_4603,N_3565,N_3978);
and U4604 (N_4604,N_3566,N_3827);
xor U4605 (N_4605,N_3263,N_3202);
nand U4606 (N_4606,N_3317,N_3791);
xnor U4607 (N_4607,N_3323,N_3700);
nand U4608 (N_4608,N_3484,N_3668);
nand U4609 (N_4609,N_3522,N_3267);
xor U4610 (N_4610,N_3574,N_3280);
nand U4611 (N_4611,N_3465,N_3894);
or U4612 (N_4612,N_3171,N_3246);
or U4613 (N_4613,N_3812,N_3840);
or U4614 (N_4614,N_3351,N_3200);
and U4615 (N_4615,N_3922,N_3370);
xor U4616 (N_4616,N_3826,N_3845);
xor U4617 (N_4617,N_3813,N_3983);
and U4618 (N_4618,N_3010,N_3039);
nand U4619 (N_4619,N_3849,N_3525);
and U4620 (N_4620,N_3913,N_3550);
nor U4621 (N_4621,N_3504,N_3700);
nor U4622 (N_4622,N_3697,N_3991);
or U4623 (N_4623,N_3977,N_3918);
nand U4624 (N_4624,N_3233,N_3285);
nor U4625 (N_4625,N_3555,N_3292);
and U4626 (N_4626,N_3660,N_3526);
nand U4627 (N_4627,N_3056,N_3249);
or U4628 (N_4628,N_3357,N_3912);
xor U4629 (N_4629,N_3465,N_3346);
nor U4630 (N_4630,N_3335,N_3745);
xor U4631 (N_4631,N_3728,N_3298);
nor U4632 (N_4632,N_3218,N_3321);
or U4633 (N_4633,N_3918,N_3069);
nor U4634 (N_4634,N_3460,N_3345);
nand U4635 (N_4635,N_3756,N_3143);
and U4636 (N_4636,N_3363,N_3080);
nand U4637 (N_4637,N_3678,N_3247);
nor U4638 (N_4638,N_3238,N_3981);
nor U4639 (N_4639,N_3902,N_3502);
nor U4640 (N_4640,N_3696,N_3771);
nand U4641 (N_4641,N_3344,N_3974);
and U4642 (N_4642,N_3942,N_3617);
nand U4643 (N_4643,N_3074,N_3751);
nor U4644 (N_4644,N_3359,N_3253);
xor U4645 (N_4645,N_3299,N_3131);
nand U4646 (N_4646,N_3846,N_3962);
nor U4647 (N_4647,N_3923,N_3300);
nor U4648 (N_4648,N_3606,N_3528);
or U4649 (N_4649,N_3816,N_3944);
xor U4650 (N_4650,N_3813,N_3238);
or U4651 (N_4651,N_3347,N_3671);
or U4652 (N_4652,N_3244,N_3154);
nand U4653 (N_4653,N_3846,N_3777);
and U4654 (N_4654,N_3715,N_3103);
or U4655 (N_4655,N_3240,N_3333);
xor U4656 (N_4656,N_3265,N_3293);
nand U4657 (N_4657,N_3693,N_3714);
or U4658 (N_4658,N_3646,N_3240);
nand U4659 (N_4659,N_3572,N_3824);
nor U4660 (N_4660,N_3395,N_3339);
or U4661 (N_4661,N_3256,N_3478);
and U4662 (N_4662,N_3391,N_3516);
and U4663 (N_4663,N_3717,N_3958);
and U4664 (N_4664,N_3293,N_3307);
nand U4665 (N_4665,N_3607,N_3625);
xor U4666 (N_4666,N_3762,N_3025);
nor U4667 (N_4667,N_3800,N_3291);
nor U4668 (N_4668,N_3843,N_3605);
nand U4669 (N_4669,N_3068,N_3446);
nand U4670 (N_4670,N_3624,N_3516);
xnor U4671 (N_4671,N_3532,N_3438);
and U4672 (N_4672,N_3867,N_3576);
and U4673 (N_4673,N_3373,N_3854);
and U4674 (N_4674,N_3191,N_3238);
and U4675 (N_4675,N_3791,N_3183);
nand U4676 (N_4676,N_3999,N_3013);
nor U4677 (N_4677,N_3413,N_3346);
xor U4678 (N_4678,N_3583,N_3312);
nor U4679 (N_4679,N_3168,N_3833);
nand U4680 (N_4680,N_3442,N_3937);
nor U4681 (N_4681,N_3244,N_3226);
nor U4682 (N_4682,N_3642,N_3319);
and U4683 (N_4683,N_3554,N_3333);
or U4684 (N_4684,N_3958,N_3374);
or U4685 (N_4685,N_3687,N_3180);
or U4686 (N_4686,N_3388,N_3731);
or U4687 (N_4687,N_3561,N_3055);
xnor U4688 (N_4688,N_3776,N_3921);
or U4689 (N_4689,N_3393,N_3668);
nor U4690 (N_4690,N_3462,N_3992);
nor U4691 (N_4691,N_3777,N_3736);
nor U4692 (N_4692,N_3339,N_3691);
nand U4693 (N_4693,N_3127,N_3344);
and U4694 (N_4694,N_3835,N_3432);
or U4695 (N_4695,N_3886,N_3968);
nand U4696 (N_4696,N_3880,N_3749);
and U4697 (N_4697,N_3282,N_3447);
and U4698 (N_4698,N_3924,N_3070);
or U4699 (N_4699,N_3315,N_3909);
and U4700 (N_4700,N_3225,N_3701);
nand U4701 (N_4701,N_3565,N_3761);
or U4702 (N_4702,N_3279,N_3347);
and U4703 (N_4703,N_3638,N_3326);
and U4704 (N_4704,N_3002,N_3374);
nor U4705 (N_4705,N_3336,N_3334);
or U4706 (N_4706,N_3947,N_3728);
nand U4707 (N_4707,N_3848,N_3756);
or U4708 (N_4708,N_3893,N_3483);
nor U4709 (N_4709,N_3263,N_3741);
or U4710 (N_4710,N_3636,N_3957);
nor U4711 (N_4711,N_3820,N_3317);
xor U4712 (N_4712,N_3625,N_3835);
nand U4713 (N_4713,N_3475,N_3660);
or U4714 (N_4714,N_3213,N_3140);
xnor U4715 (N_4715,N_3542,N_3812);
or U4716 (N_4716,N_3544,N_3981);
or U4717 (N_4717,N_3856,N_3734);
and U4718 (N_4718,N_3629,N_3460);
or U4719 (N_4719,N_3929,N_3415);
and U4720 (N_4720,N_3494,N_3743);
or U4721 (N_4721,N_3901,N_3057);
xor U4722 (N_4722,N_3367,N_3558);
and U4723 (N_4723,N_3151,N_3808);
and U4724 (N_4724,N_3979,N_3439);
nor U4725 (N_4725,N_3633,N_3700);
xor U4726 (N_4726,N_3058,N_3255);
nand U4727 (N_4727,N_3422,N_3890);
nor U4728 (N_4728,N_3351,N_3655);
nand U4729 (N_4729,N_3732,N_3454);
and U4730 (N_4730,N_3114,N_3791);
or U4731 (N_4731,N_3508,N_3452);
nor U4732 (N_4732,N_3975,N_3205);
and U4733 (N_4733,N_3916,N_3005);
xnor U4734 (N_4734,N_3091,N_3897);
and U4735 (N_4735,N_3070,N_3455);
or U4736 (N_4736,N_3289,N_3637);
or U4737 (N_4737,N_3722,N_3872);
nor U4738 (N_4738,N_3178,N_3319);
or U4739 (N_4739,N_3490,N_3711);
or U4740 (N_4740,N_3749,N_3478);
and U4741 (N_4741,N_3035,N_3122);
or U4742 (N_4742,N_3715,N_3747);
nor U4743 (N_4743,N_3965,N_3093);
or U4744 (N_4744,N_3687,N_3411);
xnor U4745 (N_4745,N_3533,N_3552);
and U4746 (N_4746,N_3877,N_3473);
nand U4747 (N_4747,N_3586,N_3554);
and U4748 (N_4748,N_3381,N_3477);
nand U4749 (N_4749,N_3586,N_3521);
xnor U4750 (N_4750,N_3599,N_3937);
or U4751 (N_4751,N_3088,N_3983);
or U4752 (N_4752,N_3706,N_3401);
or U4753 (N_4753,N_3935,N_3199);
and U4754 (N_4754,N_3218,N_3869);
xor U4755 (N_4755,N_3281,N_3259);
nand U4756 (N_4756,N_3050,N_3195);
or U4757 (N_4757,N_3697,N_3410);
or U4758 (N_4758,N_3291,N_3201);
nor U4759 (N_4759,N_3409,N_3306);
and U4760 (N_4760,N_3193,N_3178);
and U4761 (N_4761,N_3210,N_3170);
and U4762 (N_4762,N_3555,N_3562);
xnor U4763 (N_4763,N_3101,N_3256);
or U4764 (N_4764,N_3352,N_3546);
nor U4765 (N_4765,N_3141,N_3166);
nand U4766 (N_4766,N_3465,N_3033);
nand U4767 (N_4767,N_3306,N_3673);
nor U4768 (N_4768,N_3109,N_3130);
nor U4769 (N_4769,N_3813,N_3217);
or U4770 (N_4770,N_3493,N_3926);
nand U4771 (N_4771,N_3636,N_3710);
xor U4772 (N_4772,N_3982,N_3896);
or U4773 (N_4773,N_3111,N_3497);
nor U4774 (N_4774,N_3240,N_3374);
nand U4775 (N_4775,N_3748,N_3962);
nand U4776 (N_4776,N_3822,N_3067);
and U4777 (N_4777,N_3874,N_3390);
and U4778 (N_4778,N_3963,N_3044);
nor U4779 (N_4779,N_3826,N_3888);
and U4780 (N_4780,N_3575,N_3589);
nor U4781 (N_4781,N_3113,N_3802);
xor U4782 (N_4782,N_3621,N_3294);
or U4783 (N_4783,N_3252,N_3931);
nor U4784 (N_4784,N_3702,N_3618);
nor U4785 (N_4785,N_3888,N_3274);
and U4786 (N_4786,N_3285,N_3576);
or U4787 (N_4787,N_3996,N_3295);
nand U4788 (N_4788,N_3984,N_3312);
or U4789 (N_4789,N_3973,N_3997);
or U4790 (N_4790,N_3453,N_3225);
nand U4791 (N_4791,N_3445,N_3707);
nor U4792 (N_4792,N_3307,N_3560);
or U4793 (N_4793,N_3923,N_3552);
and U4794 (N_4794,N_3154,N_3099);
and U4795 (N_4795,N_3271,N_3095);
or U4796 (N_4796,N_3699,N_3292);
nor U4797 (N_4797,N_3235,N_3583);
and U4798 (N_4798,N_3926,N_3628);
nand U4799 (N_4799,N_3803,N_3770);
and U4800 (N_4800,N_3502,N_3887);
or U4801 (N_4801,N_3937,N_3636);
and U4802 (N_4802,N_3411,N_3423);
and U4803 (N_4803,N_3812,N_3260);
or U4804 (N_4804,N_3588,N_3296);
nor U4805 (N_4805,N_3018,N_3186);
xnor U4806 (N_4806,N_3797,N_3611);
and U4807 (N_4807,N_3556,N_3943);
or U4808 (N_4808,N_3024,N_3338);
nor U4809 (N_4809,N_3579,N_3010);
nor U4810 (N_4810,N_3122,N_3570);
nor U4811 (N_4811,N_3346,N_3306);
and U4812 (N_4812,N_3508,N_3619);
or U4813 (N_4813,N_3004,N_3156);
or U4814 (N_4814,N_3038,N_3743);
and U4815 (N_4815,N_3813,N_3368);
or U4816 (N_4816,N_3118,N_3282);
nor U4817 (N_4817,N_3702,N_3748);
and U4818 (N_4818,N_3442,N_3008);
or U4819 (N_4819,N_3392,N_3397);
xor U4820 (N_4820,N_3869,N_3702);
nor U4821 (N_4821,N_3034,N_3971);
nor U4822 (N_4822,N_3594,N_3329);
and U4823 (N_4823,N_3261,N_3413);
or U4824 (N_4824,N_3337,N_3228);
or U4825 (N_4825,N_3061,N_3802);
nand U4826 (N_4826,N_3390,N_3345);
and U4827 (N_4827,N_3746,N_3204);
xor U4828 (N_4828,N_3764,N_3450);
nand U4829 (N_4829,N_3690,N_3447);
xnor U4830 (N_4830,N_3623,N_3774);
or U4831 (N_4831,N_3289,N_3367);
or U4832 (N_4832,N_3609,N_3649);
nand U4833 (N_4833,N_3693,N_3425);
nor U4834 (N_4834,N_3389,N_3783);
or U4835 (N_4835,N_3248,N_3157);
nand U4836 (N_4836,N_3199,N_3391);
or U4837 (N_4837,N_3053,N_3475);
or U4838 (N_4838,N_3412,N_3828);
and U4839 (N_4839,N_3929,N_3575);
nor U4840 (N_4840,N_3940,N_3255);
or U4841 (N_4841,N_3929,N_3391);
nor U4842 (N_4842,N_3972,N_3852);
xnor U4843 (N_4843,N_3475,N_3204);
xnor U4844 (N_4844,N_3907,N_3516);
nor U4845 (N_4845,N_3485,N_3040);
nor U4846 (N_4846,N_3218,N_3787);
nor U4847 (N_4847,N_3964,N_3828);
nand U4848 (N_4848,N_3918,N_3326);
and U4849 (N_4849,N_3963,N_3490);
nor U4850 (N_4850,N_3454,N_3107);
nor U4851 (N_4851,N_3441,N_3208);
and U4852 (N_4852,N_3224,N_3191);
nor U4853 (N_4853,N_3491,N_3932);
xor U4854 (N_4854,N_3994,N_3700);
or U4855 (N_4855,N_3639,N_3020);
nand U4856 (N_4856,N_3652,N_3670);
nand U4857 (N_4857,N_3743,N_3627);
and U4858 (N_4858,N_3673,N_3925);
or U4859 (N_4859,N_3546,N_3454);
nand U4860 (N_4860,N_3505,N_3050);
nor U4861 (N_4861,N_3403,N_3964);
and U4862 (N_4862,N_3385,N_3899);
xor U4863 (N_4863,N_3157,N_3718);
nor U4864 (N_4864,N_3786,N_3551);
and U4865 (N_4865,N_3270,N_3061);
or U4866 (N_4866,N_3464,N_3998);
xnor U4867 (N_4867,N_3996,N_3575);
and U4868 (N_4868,N_3452,N_3720);
nor U4869 (N_4869,N_3370,N_3595);
xnor U4870 (N_4870,N_3419,N_3982);
and U4871 (N_4871,N_3483,N_3900);
nor U4872 (N_4872,N_3980,N_3948);
or U4873 (N_4873,N_3883,N_3112);
and U4874 (N_4874,N_3534,N_3260);
and U4875 (N_4875,N_3570,N_3219);
and U4876 (N_4876,N_3907,N_3725);
nor U4877 (N_4877,N_3973,N_3628);
and U4878 (N_4878,N_3119,N_3492);
nand U4879 (N_4879,N_3569,N_3075);
or U4880 (N_4880,N_3674,N_3269);
nand U4881 (N_4881,N_3508,N_3923);
xor U4882 (N_4882,N_3475,N_3500);
or U4883 (N_4883,N_3820,N_3029);
nand U4884 (N_4884,N_3647,N_3512);
or U4885 (N_4885,N_3469,N_3906);
nor U4886 (N_4886,N_3852,N_3042);
or U4887 (N_4887,N_3082,N_3585);
nand U4888 (N_4888,N_3259,N_3534);
nand U4889 (N_4889,N_3700,N_3126);
and U4890 (N_4890,N_3026,N_3965);
nor U4891 (N_4891,N_3710,N_3200);
and U4892 (N_4892,N_3528,N_3889);
nand U4893 (N_4893,N_3562,N_3887);
nand U4894 (N_4894,N_3417,N_3045);
or U4895 (N_4895,N_3405,N_3629);
and U4896 (N_4896,N_3417,N_3879);
nand U4897 (N_4897,N_3127,N_3437);
and U4898 (N_4898,N_3969,N_3257);
nand U4899 (N_4899,N_3190,N_3715);
nor U4900 (N_4900,N_3640,N_3342);
and U4901 (N_4901,N_3996,N_3261);
and U4902 (N_4902,N_3384,N_3268);
or U4903 (N_4903,N_3034,N_3247);
and U4904 (N_4904,N_3019,N_3120);
nor U4905 (N_4905,N_3634,N_3749);
xnor U4906 (N_4906,N_3711,N_3088);
xor U4907 (N_4907,N_3504,N_3895);
nor U4908 (N_4908,N_3550,N_3535);
nand U4909 (N_4909,N_3453,N_3157);
nand U4910 (N_4910,N_3320,N_3271);
nand U4911 (N_4911,N_3537,N_3018);
nand U4912 (N_4912,N_3141,N_3847);
nand U4913 (N_4913,N_3890,N_3464);
nand U4914 (N_4914,N_3854,N_3299);
or U4915 (N_4915,N_3875,N_3471);
nand U4916 (N_4916,N_3058,N_3683);
and U4917 (N_4917,N_3531,N_3126);
or U4918 (N_4918,N_3423,N_3823);
and U4919 (N_4919,N_3944,N_3198);
nand U4920 (N_4920,N_3226,N_3158);
and U4921 (N_4921,N_3745,N_3994);
xor U4922 (N_4922,N_3619,N_3613);
or U4923 (N_4923,N_3706,N_3320);
nor U4924 (N_4924,N_3248,N_3709);
and U4925 (N_4925,N_3144,N_3764);
and U4926 (N_4926,N_3210,N_3686);
nor U4927 (N_4927,N_3785,N_3282);
or U4928 (N_4928,N_3308,N_3327);
nand U4929 (N_4929,N_3982,N_3791);
and U4930 (N_4930,N_3588,N_3227);
nand U4931 (N_4931,N_3854,N_3959);
nand U4932 (N_4932,N_3487,N_3546);
nand U4933 (N_4933,N_3502,N_3054);
and U4934 (N_4934,N_3435,N_3984);
nand U4935 (N_4935,N_3258,N_3846);
xor U4936 (N_4936,N_3356,N_3696);
nand U4937 (N_4937,N_3252,N_3235);
nor U4938 (N_4938,N_3400,N_3774);
nand U4939 (N_4939,N_3089,N_3486);
nor U4940 (N_4940,N_3161,N_3512);
or U4941 (N_4941,N_3130,N_3922);
or U4942 (N_4942,N_3077,N_3555);
nand U4943 (N_4943,N_3837,N_3359);
nor U4944 (N_4944,N_3733,N_3989);
nand U4945 (N_4945,N_3378,N_3631);
xnor U4946 (N_4946,N_3010,N_3339);
or U4947 (N_4947,N_3411,N_3672);
xnor U4948 (N_4948,N_3071,N_3886);
and U4949 (N_4949,N_3284,N_3810);
xor U4950 (N_4950,N_3587,N_3259);
nor U4951 (N_4951,N_3800,N_3905);
nand U4952 (N_4952,N_3503,N_3852);
or U4953 (N_4953,N_3045,N_3819);
or U4954 (N_4954,N_3422,N_3370);
and U4955 (N_4955,N_3051,N_3633);
xor U4956 (N_4956,N_3719,N_3639);
xor U4957 (N_4957,N_3091,N_3373);
or U4958 (N_4958,N_3136,N_3958);
xnor U4959 (N_4959,N_3122,N_3997);
nand U4960 (N_4960,N_3630,N_3900);
or U4961 (N_4961,N_3363,N_3550);
nor U4962 (N_4962,N_3472,N_3221);
or U4963 (N_4963,N_3405,N_3052);
xnor U4964 (N_4964,N_3416,N_3611);
or U4965 (N_4965,N_3024,N_3704);
nor U4966 (N_4966,N_3539,N_3235);
nand U4967 (N_4967,N_3514,N_3690);
xnor U4968 (N_4968,N_3803,N_3558);
and U4969 (N_4969,N_3363,N_3907);
nand U4970 (N_4970,N_3037,N_3317);
or U4971 (N_4971,N_3461,N_3448);
and U4972 (N_4972,N_3661,N_3231);
nand U4973 (N_4973,N_3950,N_3652);
or U4974 (N_4974,N_3587,N_3668);
nor U4975 (N_4975,N_3834,N_3666);
nor U4976 (N_4976,N_3781,N_3511);
nand U4977 (N_4977,N_3343,N_3427);
and U4978 (N_4978,N_3248,N_3129);
nand U4979 (N_4979,N_3177,N_3774);
nor U4980 (N_4980,N_3378,N_3517);
or U4981 (N_4981,N_3375,N_3091);
and U4982 (N_4982,N_3546,N_3839);
nor U4983 (N_4983,N_3885,N_3135);
nand U4984 (N_4984,N_3393,N_3020);
or U4985 (N_4985,N_3181,N_3423);
nor U4986 (N_4986,N_3156,N_3811);
and U4987 (N_4987,N_3976,N_3418);
nor U4988 (N_4988,N_3753,N_3633);
and U4989 (N_4989,N_3568,N_3737);
or U4990 (N_4990,N_3497,N_3828);
and U4991 (N_4991,N_3637,N_3065);
nor U4992 (N_4992,N_3073,N_3113);
or U4993 (N_4993,N_3072,N_3454);
nand U4994 (N_4994,N_3381,N_3780);
and U4995 (N_4995,N_3002,N_3138);
and U4996 (N_4996,N_3162,N_3441);
and U4997 (N_4997,N_3170,N_3434);
and U4998 (N_4998,N_3607,N_3691);
or U4999 (N_4999,N_3550,N_3898);
or U5000 (N_5000,N_4259,N_4159);
nor U5001 (N_5001,N_4086,N_4476);
and U5002 (N_5002,N_4134,N_4613);
nor U5003 (N_5003,N_4985,N_4514);
nor U5004 (N_5004,N_4633,N_4709);
or U5005 (N_5005,N_4933,N_4844);
and U5006 (N_5006,N_4503,N_4301);
nor U5007 (N_5007,N_4160,N_4698);
nand U5008 (N_5008,N_4750,N_4278);
and U5009 (N_5009,N_4625,N_4911);
or U5010 (N_5010,N_4900,N_4415);
nor U5011 (N_5011,N_4426,N_4334);
or U5012 (N_5012,N_4240,N_4832);
and U5013 (N_5013,N_4353,N_4117);
and U5014 (N_5014,N_4712,N_4345);
nor U5015 (N_5015,N_4688,N_4665);
nand U5016 (N_5016,N_4536,N_4286);
or U5017 (N_5017,N_4987,N_4223);
nand U5018 (N_5018,N_4372,N_4109);
nand U5019 (N_5019,N_4010,N_4733);
and U5020 (N_5020,N_4848,N_4738);
or U5021 (N_5021,N_4128,N_4899);
nor U5022 (N_5022,N_4910,N_4367);
nor U5023 (N_5023,N_4091,N_4041);
nand U5024 (N_5024,N_4178,N_4836);
xor U5025 (N_5025,N_4562,N_4168);
or U5026 (N_5026,N_4115,N_4690);
nor U5027 (N_5027,N_4611,N_4151);
nand U5028 (N_5028,N_4204,N_4771);
nor U5029 (N_5029,N_4138,N_4045);
nand U5030 (N_5030,N_4004,N_4057);
and U5031 (N_5031,N_4338,N_4608);
xor U5032 (N_5032,N_4953,N_4099);
or U5033 (N_5033,N_4837,N_4724);
nand U5034 (N_5034,N_4105,N_4454);
nand U5035 (N_5035,N_4304,N_4446);
nand U5036 (N_5036,N_4157,N_4827);
and U5037 (N_5037,N_4965,N_4671);
and U5038 (N_5038,N_4340,N_4731);
xor U5039 (N_5039,N_4834,N_4428);
or U5040 (N_5040,N_4918,N_4571);
or U5041 (N_5041,N_4579,N_4840);
or U5042 (N_5042,N_4002,N_4528);
and U5043 (N_5043,N_4743,N_4598);
and U5044 (N_5044,N_4084,N_4810);
xnor U5045 (N_5045,N_4211,N_4385);
nand U5046 (N_5046,N_4043,N_4470);
or U5047 (N_5047,N_4387,N_4683);
or U5048 (N_5048,N_4129,N_4904);
or U5049 (N_5049,N_4967,N_4107);
nand U5050 (N_5050,N_4144,N_4578);
and U5051 (N_5051,N_4461,N_4110);
or U5052 (N_5052,N_4568,N_4746);
or U5053 (N_5053,N_4540,N_4484);
nor U5054 (N_5054,N_4508,N_4612);
or U5055 (N_5055,N_4251,N_4245);
and U5056 (N_5056,N_4335,N_4298);
xor U5057 (N_5057,N_4591,N_4560);
nor U5058 (N_5058,N_4894,N_4203);
or U5059 (N_5059,N_4255,N_4890);
nand U5060 (N_5060,N_4457,N_4914);
and U5061 (N_5061,N_4843,N_4992);
xor U5062 (N_5062,N_4988,N_4627);
and U5063 (N_5063,N_4063,N_4352);
xor U5064 (N_5064,N_4552,N_4363);
nand U5065 (N_5065,N_4575,N_4088);
xor U5066 (N_5066,N_4893,N_4871);
nor U5067 (N_5067,N_4821,N_4408);
nor U5068 (N_5068,N_4268,N_4262);
xnor U5069 (N_5069,N_4137,N_4441);
and U5070 (N_5070,N_4563,N_4475);
nor U5071 (N_5071,N_4477,N_4153);
and U5072 (N_5072,N_4773,N_4456);
and U5073 (N_5073,N_4407,N_4977);
and U5074 (N_5074,N_4290,N_4735);
nor U5075 (N_5075,N_4649,N_4725);
nor U5076 (N_5076,N_4691,N_4819);
and U5077 (N_5077,N_4588,N_4865);
nor U5078 (N_5078,N_4806,N_4554);
nand U5079 (N_5079,N_4418,N_4142);
nor U5080 (N_5080,N_4346,N_4551);
or U5081 (N_5081,N_4845,N_4960);
and U5082 (N_5082,N_4609,N_4047);
nor U5083 (N_5083,N_4319,N_4523);
and U5084 (N_5084,N_4669,N_4077);
nand U5085 (N_5085,N_4677,N_4708);
and U5086 (N_5086,N_4530,N_4841);
nand U5087 (N_5087,N_4713,N_4616);
nand U5088 (N_5088,N_4235,N_4141);
or U5089 (N_5089,N_4417,N_4777);
nor U5090 (N_5090,N_4539,N_4440);
or U5091 (N_5091,N_4429,N_4519);
nand U5092 (N_5092,N_4732,N_4720);
nor U5093 (N_5093,N_4497,N_4792);
and U5094 (N_5094,N_4909,N_4023);
nand U5095 (N_5095,N_4557,N_4584);
xor U5096 (N_5096,N_4167,N_4413);
nand U5097 (N_5097,N_4747,N_4762);
and U5098 (N_5098,N_4220,N_4228);
and U5099 (N_5099,N_4550,N_4132);
nand U5100 (N_5100,N_4897,N_4814);
nor U5101 (N_5101,N_4863,N_4615);
nor U5102 (N_5102,N_4740,N_4222);
nor U5103 (N_5103,N_4487,N_4518);
and U5104 (N_5104,N_4087,N_4823);
nor U5105 (N_5105,N_4797,N_4788);
and U5106 (N_5106,N_4246,N_4486);
nor U5107 (N_5107,N_4573,N_4617);
or U5108 (N_5108,N_4705,N_4650);
and U5109 (N_5109,N_4076,N_4394);
xnor U5110 (N_5110,N_4504,N_4804);
nand U5111 (N_5111,N_4870,N_4012);
and U5112 (N_5112,N_4913,N_4005);
and U5113 (N_5113,N_4036,N_4420);
xnor U5114 (N_5114,N_4386,N_4316);
xor U5115 (N_5115,N_4040,N_4383);
nand U5116 (N_5116,N_4274,N_4603);
nand U5117 (N_5117,N_4405,N_4048);
nand U5118 (N_5118,N_4053,N_4793);
and U5119 (N_5119,N_4825,N_4474);
and U5120 (N_5120,N_4171,N_4473);
and U5121 (N_5121,N_4499,N_4604);
or U5122 (N_5122,N_4368,N_4051);
nor U5123 (N_5123,N_4139,N_4555);
and U5124 (N_5124,N_4674,N_4857);
and U5125 (N_5125,N_4585,N_4937);
nor U5126 (N_5126,N_4285,N_4449);
nand U5127 (N_5127,N_4196,N_4459);
and U5128 (N_5128,N_4136,N_4124);
nand U5129 (N_5129,N_4347,N_4730);
or U5130 (N_5130,N_4984,N_4064);
and U5131 (N_5131,N_4166,N_4719);
nand U5132 (N_5132,N_4920,N_4080);
and U5133 (N_5133,N_4995,N_4875);
and U5134 (N_5134,N_4097,N_4968);
and U5135 (N_5135,N_4974,N_4685);
nor U5136 (N_5136,N_4774,N_4619);
or U5137 (N_5137,N_4782,N_4791);
or U5138 (N_5138,N_4453,N_4780);
and U5139 (N_5139,N_4233,N_4243);
nand U5140 (N_5140,N_4739,N_4288);
nand U5141 (N_5141,N_4763,N_4325);
xnor U5142 (N_5142,N_4976,N_4775);
and U5143 (N_5143,N_4994,N_4496);
nand U5144 (N_5144,N_4905,N_4506);
nor U5145 (N_5145,N_4037,N_4670);
or U5146 (N_5146,N_4951,N_4143);
nor U5147 (N_5147,N_4833,N_4558);
or U5148 (N_5148,N_4637,N_4860);
or U5149 (N_5149,N_4892,N_4435);
nand U5150 (N_5150,N_4714,N_4851);
or U5151 (N_5151,N_4501,N_4807);
or U5152 (N_5152,N_4626,N_4458);
nor U5153 (N_5153,N_4513,N_4629);
nor U5154 (N_5154,N_4336,N_4675);
and U5155 (N_5155,N_4073,N_4831);
or U5156 (N_5156,N_4970,N_4483);
nor U5157 (N_5157,N_4582,N_4645);
and U5158 (N_5158,N_4013,N_4252);
or U5159 (N_5159,N_4277,N_4515);
nand U5160 (N_5160,N_4303,N_4718);
or U5161 (N_5161,N_4664,N_4172);
nor U5162 (N_5162,N_4083,N_4666);
nand U5163 (N_5163,N_4856,N_4266);
and U5164 (N_5164,N_4502,N_4812);
nor U5165 (N_5165,N_4924,N_4663);
or U5166 (N_5166,N_4225,N_4498);
nand U5167 (N_5167,N_4210,N_4442);
nor U5168 (N_5168,N_4853,N_4123);
nor U5169 (N_5169,N_4206,N_4755);
xor U5170 (N_5170,N_4727,N_4276);
and U5171 (N_5171,N_4500,N_4958);
nand U5172 (N_5172,N_4697,N_4672);
nor U5173 (N_5173,N_4706,N_4219);
nor U5174 (N_5174,N_4521,N_4309);
or U5175 (N_5175,N_4015,N_4054);
or U5176 (N_5176,N_4280,N_4642);
and U5177 (N_5177,N_4926,N_4902);
nor U5178 (N_5178,N_4018,N_4776);
nor U5179 (N_5179,N_4576,N_4945);
and U5180 (N_5180,N_4721,N_4438);
nand U5181 (N_5181,N_4399,N_4886);
or U5182 (N_5182,N_4574,N_4194);
nor U5183 (N_5183,N_4640,N_4195);
and U5184 (N_5184,N_4366,N_4361);
nor U5185 (N_5185,N_4180,N_4569);
xnor U5186 (N_5186,N_4990,N_4330);
or U5187 (N_5187,N_4027,N_4273);
and U5188 (N_5188,N_4207,N_4849);
nor U5189 (N_5189,N_4131,N_4261);
nand U5190 (N_5190,N_4895,N_4751);
and U5191 (N_5191,N_4090,N_4964);
xor U5192 (N_5192,N_4855,N_4781);
nor U5193 (N_5193,N_4177,N_4947);
or U5194 (N_5194,N_4511,N_4534);
nand U5195 (N_5195,N_4093,N_4601);
xnor U5196 (N_5196,N_4433,N_4232);
and U5197 (N_5197,N_4916,N_4049);
nor U5198 (N_5198,N_4050,N_4946);
nor U5199 (N_5199,N_4711,N_4737);
xor U5200 (N_5200,N_4770,N_4074);
or U5201 (N_5201,N_4314,N_4622);
or U5202 (N_5202,N_4798,N_4787);
nand U5203 (N_5203,N_4800,N_4492);
nor U5204 (N_5204,N_4891,N_4039);
nor U5205 (N_5205,N_4692,N_4313);
and U5206 (N_5206,N_4963,N_4779);
and U5207 (N_5207,N_4898,N_4029);
and U5208 (N_5208,N_4300,N_4120);
nor U5209 (N_5209,N_4809,N_4481);
xnor U5210 (N_5210,N_4969,N_4422);
nand U5211 (N_5211,N_4885,N_4795);
nor U5212 (N_5212,N_4308,N_4516);
and U5213 (N_5213,N_4305,N_4033);
nor U5214 (N_5214,N_4699,N_4021);
or U5215 (N_5215,N_4025,N_4962);
or U5216 (N_5216,N_4344,N_4238);
nand U5217 (N_5217,N_4289,N_4365);
or U5218 (N_5218,N_4936,N_4455);
or U5219 (N_5219,N_4643,N_4250);
nor U5220 (N_5220,N_4060,N_4148);
nor U5221 (N_5221,N_4269,N_4130);
or U5222 (N_5222,N_4906,N_4022);
or U5223 (N_5223,N_4864,N_4146);
and U5224 (N_5224,N_4191,N_4075);
nand U5225 (N_5225,N_4358,N_4348);
or U5226 (N_5226,N_4693,N_4009);
and U5227 (N_5227,N_4430,N_4955);
or U5228 (N_5228,N_4566,N_4876);
nor U5229 (N_5229,N_4260,N_4101);
nand U5230 (N_5230,N_4778,N_4597);
xor U5231 (N_5231,N_4371,N_4662);
or U5232 (N_5232,N_4785,N_4887);
and U5233 (N_5233,N_4654,N_4014);
nor U5234 (N_5234,N_4636,N_4034);
xnor U5235 (N_5235,N_4586,N_4212);
xnor U5236 (N_5236,N_4059,N_4676);
and U5237 (N_5237,N_4541,N_4623);
and U5238 (N_5238,N_4401,N_4479);
nand U5239 (N_5239,N_4001,N_4607);
nand U5240 (N_5240,N_4218,N_4509);
xnor U5241 (N_5241,N_4526,N_4024);
nand U5242 (N_5242,N_4265,N_4042);
nand U5243 (N_5243,N_4297,N_4412);
nor U5244 (N_5244,N_4802,N_4614);
nand U5245 (N_5245,N_4877,N_4700);
and U5246 (N_5246,N_4764,N_4769);
and U5247 (N_5247,N_4247,N_4306);
xor U5248 (N_5248,N_4606,N_4928);
nand U5249 (N_5249,N_4468,N_4444);
nand U5250 (N_5250,N_4324,N_4038);
or U5251 (N_5251,N_4374,N_4000);
and U5252 (N_5252,N_4436,N_4862);
and U5253 (N_5253,N_4017,N_4098);
nand U5254 (N_5254,N_4150,N_4103);
and U5255 (N_5255,N_4164,N_4230);
or U5256 (N_5256,N_4684,N_4535);
or U5257 (N_5257,N_4572,N_4801);
and U5258 (N_5258,N_4495,N_4320);
xnor U5259 (N_5259,N_4696,N_4198);
or U5260 (N_5260,N_4646,N_4941);
or U5261 (N_5261,N_4859,N_4370);
or U5262 (N_5262,N_4409,N_4618);
or U5263 (N_5263,N_4193,N_4874);
nand U5264 (N_5264,N_4227,N_4881);
or U5265 (N_5265,N_4332,N_4527);
nand U5266 (N_5266,N_4546,N_4307);
and U5267 (N_5267,N_4704,N_4111);
nand U5268 (N_5268,N_4201,N_4217);
xnor U5269 (N_5269,N_4263,N_4373);
xor U5270 (N_5270,N_4016,N_4469);
or U5271 (N_5271,N_4971,N_4478);
nor U5272 (N_5272,N_4961,N_4184);
xor U5273 (N_5273,N_4384,N_4872);
and U5274 (N_5274,N_4581,N_4085);
and U5275 (N_5275,N_4723,N_4765);
or U5276 (N_5276,N_4402,N_4679);
and U5277 (N_5277,N_4754,N_4125);
or U5278 (N_5278,N_4903,N_4322);
nand U5279 (N_5279,N_4998,N_4467);
xnor U5280 (N_5280,N_4364,N_4689);
and U5281 (N_5281,N_4295,N_4156);
nand U5282 (N_5282,N_4728,N_4078);
xnor U5283 (N_5283,N_4587,N_4861);
or U5284 (N_5284,N_4279,N_4517);
and U5285 (N_5285,N_4339,N_4231);
nand U5286 (N_5286,N_4326,N_4596);
nor U5287 (N_5287,N_4653,N_4826);
or U5288 (N_5288,N_4242,N_4427);
and U5289 (N_5289,N_4678,N_4152);
or U5290 (N_5290,N_4032,N_4377);
nor U5291 (N_5291,N_4185,N_4189);
xor U5292 (N_5292,N_4256,N_4561);
xor U5293 (N_5293,N_4452,N_4239);
nand U5294 (N_5294,N_4439,N_4652);
or U5295 (N_5295,N_4410,N_4659);
or U5296 (N_5296,N_4888,N_4957);
nand U5297 (N_5297,N_4866,N_4956);
nand U5298 (N_5298,N_4556,N_4434);
nand U5299 (N_5299,N_4174,N_4959);
xnor U5300 (N_5300,N_4443,N_4681);
nand U5301 (N_5301,N_4208,N_4342);
nand U5302 (N_5302,N_4717,N_4667);
and U5303 (N_5303,N_4533,N_4726);
and U5304 (N_5304,N_4736,N_4980);
xor U5305 (N_5305,N_4046,N_4828);
nor U5306 (N_5306,N_4628,N_4471);
nor U5307 (N_5307,N_4982,N_4082);
and U5308 (N_5308,N_4062,N_4624);
xnor U5309 (N_5309,N_4448,N_4829);
xor U5310 (N_5310,N_4026,N_4154);
xnor U5311 (N_5311,N_4553,N_4915);
nor U5312 (N_5312,N_4602,N_4466);
xor U5313 (N_5313,N_4337,N_4522);
nor U5314 (N_5314,N_4391,N_4068);
nand U5315 (N_5315,N_4701,N_4935);
or U5316 (N_5316,N_4999,N_4249);
nor U5317 (N_5317,N_4818,N_4419);
nor U5318 (N_5318,N_4752,N_4545);
nor U5319 (N_5319,N_4165,N_4388);
and U5320 (N_5320,N_4593,N_4100);
xnor U5321 (N_5321,N_4092,N_4954);
and U5322 (N_5322,N_4236,N_4912);
and U5323 (N_5323,N_4379,N_4925);
and U5324 (N_5324,N_4794,N_4096);
nand U5325 (N_5325,N_4395,N_4796);
or U5326 (N_5326,N_4271,N_4594);
or U5327 (N_5327,N_4710,N_4272);
or U5328 (N_5328,N_4199,N_4996);
nor U5329 (N_5329,N_4748,N_4917);
and U5330 (N_5330,N_4424,N_4600);
xnor U5331 (N_5331,N_4161,N_4943);
nand U5332 (N_5332,N_4291,N_4414);
or U5333 (N_5333,N_4835,N_4072);
and U5334 (N_5334,N_4565,N_4451);
nor U5335 (N_5335,N_4173,N_4820);
nand U5336 (N_5336,N_4425,N_4482);
and U5337 (N_5337,N_4396,N_4462);
and U5338 (N_5338,N_4922,N_4651);
nor U5339 (N_5339,N_4008,N_4112);
or U5340 (N_5340,N_4376,N_4020);
and U5341 (N_5341,N_4661,N_4753);
or U5342 (N_5342,N_4331,N_4544);
or U5343 (N_5343,N_4140,N_4067);
and U5344 (N_5344,N_4716,N_4981);
and U5345 (N_5345,N_4932,N_4393);
xor U5346 (N_5346,N_4284,N_4170);
or U5347 (N_5347,N_4879,N_4229);
and U5348 (N_5348,N_4382,N_4878);
nor U5349 (N_5349,N_4197,N_4816);
nand U5350 (N_5350,N_4842,N_4310);
and U5351 (N_5351,N_4254,N_4437);
and U5352 (N_5352,N_4610,N_4811);
or U5353 (N_5353,N_4592,N_4460);
nor U5354 (N_5354,N_4986,N_4445);
or U5355 (N_5355,N_4850,N_4595);
and U5356 (N_5356,N_4564,N_4119);
or U5357 (N_5357,N_4873,N_4491);
nand U5358 (N_5358,N_4525,N_4095);
or U5359 (N_5359,N_4464,N_4817);
xnor U5360 (N_5360,N_4880,N_4356);
nand U5361 (N_5361,N_4003,N_4357);
nor U5362 (N_5362,N_4923,N_4948);
or U5363 (N_5363,N_4241,N_4949);
nor U5364 (N_5364,N_4655,N_4056);
nand U5365 (N_5365,N_4432,N_4214);
nand U5366 (N_5366,N_4296,N_4884);
xor U5367 (N_5367,N_4416,N_4094);
or U5368 (N_5368,N_4397,N_4318);
xnor U5369 (N_5369,N_4846,N_4639);
and U5370 (N_5370,N_4389,N_4055);
or U5371 (N_5371,N_4852,N_4993);
nor U5372 (N_5372,N_4803,N_4934);
nor U5373 (N_5373,N_4179,N_4789);
xor U5374 (N_5374,N_4108,N_4605);
nor U5375 (N_5375,N_4169,N_4071);
or U5376 (N_5376,N_4808,N_4411);
nor U5377 (N_5377,N_4549,N_4343);
nor U5378 (N_5378,N_4749,N_4181);
nor U5379 (N_5379,N_4267,N_4813);
nand U5380 (N_5380,N_4707,N_4896);
nor U5381 (N_5381,N_4421,N_4767);
and U5382 (N_5382,N_4537,N_4830);
nor U5383 (N_5383,N_4044,N_4400);
nor U5384 (N_5384,N_4931,N_4673);
or U5385 (N_5385,N_4145,N_4938);
or U5386 (N_5386,N_4599,N_4360);
nand U5387 (N_5387,N_4989,N_4589);
or U5388 (N_5388,N_4490,N_4580);
nor U5389 (N_5389,N_4494,N_4973);
nand U5390 (N_5390,N_4761,N_4686);
nor U5391 (N_5391,N_4991,N_4529);
nand U5392 (N_5392,N_4327,N_4822);
nand U5393 (N_5393,N_4149,N_4312);
or U5394 (N_5394,N_4532,N_4919);
and U5395 (N_5395,N_4351,N_4950);
nand U5396 (N_5396,N_4321,N_4734);
or U5397 (N_5397,N_4634,N_4378);
nor U5398 (N_5398,N_4799,N_4641);
and U5399 (N_5399,N_4052,N_4703);
or U5400 (N_5400,N_4694,N_4258);
or U5401 (N_5401,N_4621,N_4742);
or U5402 (N_5402,N_4213,N_4889);
and U5403 (N_5403,N_4715,N_4507);
or U5404 (N_5404,N_4224,N_4404);
or U5405 (N_5405,N_4590,N_4398);
nor U5406 (N_5406,N_4907,N_4349);
xor U5407 (N_5407,N_4175,N_4768);
xnor U5408 (N_5408,N_4695,N_4390);
or U5409 (N_5409,N_4081,N_4786);
or U5410 (N_5410,N_4729,N_4680);
and U5411 (N_5411,N_4403,N_4485);
nand U5412 (N_5412,N_4510,N_4660);
or U5413 (N_5413,N_4237,N_4183);
and U5414 (N_5414,N_4538,N_4035);
and U5415 (N_5415,N_4293,N_4058);
or U5416 (N_5416,N_4952,N_4070);
or U5417 (N_5417,N_4186,N_4940);
nand U5418 (N_5418,N_4190,N_4983);
or U5419 (N_5419,N_4858,N_4647);
and U5420 (N_5420,N_4253,N_4784);
xnor U5421 (N_5421,N_4543,N_4317);
or U5422 (N_5422,N_4283,N_4908);
or U5423 (N_5423,N_4163,N_4011);
or U5424 (N_5424,N_4531,N_4202);
nand U5425 (N_5425,N_4282,N_4176);
and U5426 (N_5426,N_4979,N_4205);
nand U5427 (N_5427,N_4065,N_4463);
or U5428 (N_5428,N_4133,N_4121);
xor U5429 (N_5429,N_4216,N_4741);
or U5430 (N_5430,N_4069,N_4978);
nand U5431 (N_5431,N_4355,N_4362);
or U5432 (N_5432,N_4847,N_4155);
or U5433 (N_5433,N_4632,N_4323);
and U5434 (N_5434,N_4760,N_4548);
or U5435 (N_5435,N_4192,N_4375);
nor U5436 (N_5436,N_4577,N_4570);
nor U5437 (N_5437,N_4630,N_4854);
nor U5438 (N_5438,N_4089,N_4031);
nand U5439 (N_5439,N_4638,N_4722);
or U5440 (N_5440,N_4512,N_4480);
nand U5441 (N_5441,N_4028,N_4359);
nand U5442 (N_5442,N_4244,N_4315);
and U5443 (N_5443,N_4758,N_4583);
and U5444 (N_5444,N_4270,N_4868);
nor U5445 (N_5445,N_4209,N_4882);
nor U5446 (N_5446,N_4328,N_4187);
nand U5447 (N_5447,N_4182,N_4867);
nor U5448 (N_5448,N_4524,N_4423);
nand U5449 (N_5449,N_4972,N_4406);
nor U5450 (N_5450,N_4975,N_4921);
nand U5451 (N_5451,N_4215,N_4234);
nand U5452 (N_5452,N_4966,N_4431);
and U5453 (N_5453,N_4311,N_4380);
and U5454 (N_5454,N_4657,N_4489);
or U5455 (N_5455,N_4547,N_4901);
nand U5456 (N_5456,N_4354,N_4682);
nand U5457 (N_5457,N_4221,N_4226);
nand U5458 (N_5458,N_4162,N_4927);
xor U5459 (N_5459,N_4079,N_4635);
nor U5460 (N_5460,N_4006,N_4188);
nand U5461 (N_5461,N_4333,N_4007);
nor U5462 (N_5462,N_4116,N_4299);
and U5463 (N_5463,N_4930,N_4465);
nor U5464 (N_5464,N_4559,N_4381);
or U5465 (N_5465,N_4869,N_4944);
or U5466 (N_5466,N_4772,N_4104);
nand U5467 (N_5467,N_4350,N_4839);
and U5468 (N_5468,N_4147,N_4294);
xnor U5469 (N_5469,N_4113,N_4702);
nor U5470 (N_5470,N_4668,N_4493);
nand U5471 (N_5471,N_4805,N_4200);
nand U5472 (N_5472,N_4745,N_4275);
nand U5473 (N_5473,N_4102,N_4542);
nor U5474 (N_5474,N_4620,N_4790);
and U5475 (N_5475,N_4329,N_4472);
and U5476 (N_5476,N_4815,N_4341);
and U5477 (N_5477,N_4127,N_4118);
nand U5478 (N_5478,N_4257,N_4648);
nand U5479 (N_5479,N_4939,N_4766);
xnor U5480 (N_5480,N_4264,N_4135);
nand U5481 (N_5481,N_4997,N_4759);
nand U5482 (N_5482,N_4292,N_4488);
or U5483 (N_5483,N_4756,N_4126);
or U5484 (N_5484,N_4450,N_4122);
xor U5485 (N_5485,N_4929,N_4658);
and U5486 (N_5486,N_4656,N_4757);
or U5487 (N_5487,N_4392,N_4783);
nor U5488 (N_5488,N_4838,N_4520);
xor U5489 (N_5489,N_4505,N_4287);
or U5490 (N_5490,N_4066,N_4030);
xor U5491 (N_5491,N_4824,N_4106);
or U5492 (N_5492,N_4061,N_4019);
nor U5493 (N_5493,N_4158,N_4942);
nor U5494 (N_5494,N_4744,N_4248);
nand U5495 (N_5495,N_4644,N_4687);
xnor U5496 (N_5496,N_4302,N_4883);
nand U5497 (N_5497,N_4281,N_4631);
and U5498 (N_5498,N_4447,N_4369);
nand U5499 (N_5499,N_4567,N_4114);
or U5500 (N_5500,N_4111,N_4653);
nor U5501 (N_5501,N_4680,N_4089);
xor U5502 (N_5502,N_4302,N_4568);
nor U5503 (N_5503,N_4691,N_4114);
and U5504 (N_5504,N_4678,N_4564);
nand U5505 (N_5505,N_4828,N_4521);
or U5506 (N_5506,N_4421,N_4820);
nand U5507 (N_5507,N_4833,N_4750);
and U5508 (N_5508,N_4234,N_4555);
xor U5509 (N_5509,N_4810,N_4312);
xnor U5510 (N_5510,N_4929,N_4932);
nand U5511 (N_5511,N_4242,N_4603);
nand U5512 (N_5512,N_4766,N_4439);
xnor U5513 (N_5513,N_4892,N_4672);
nand U5514 (N_5514,N_4251,N_4454);
nor U5515 (N_5515,N_4811,N_4980);
nand U5516 (N_5516,N_4199,N_4769);
and U5517 (N_5517,N_4897,N_4683);
nor U5518 (N_5518,N_4246,N_4370);
or U5519 (N_5519,N_4914,N_4993);
and U5520 (N_5520,N_4342,N_4913);
and U5521 (N_5521,N_4868,N_4141);
and U5522 (N_5522,N_4728,N_4132);
or U5523 (N_5523,N_4117,N_4352);
nor U5524 (N_5524,N_4783,N_4843);
xnor U5525 (N_5525,N_4652,N_4094);
or U5526 (N_5526,N_4695,N_4795);
nand U5527 (N_5527,N_4440,N_4083);
and U5528 (N_5528,N_4063,N_4015);
or U5529 (N_5529,N_4387,N_4643);
nand U5530 (N_5530,N_4545,N_4886);
nor U5531 (N_5531,N_4746,N_4687);
nand U5532 (N_5532,N_4778,N_4504);
xnor U5533 (N_5533,N_4869,N_4225);
and U5534 (N_5534,N_4699,N_4057);
or U5535 (N_5535,N_4650,N_4691);
and U5536 (N_5536,N_4099,N_4392);
and U5537 (N_5537,N_4613,N_4263);
nor U5538 (N_5538,N_4093,N_4354);
nand U5539 (N_5539,N_4116,N_4960);
and U5540 (N_5540,N_4937,N_4060);
nand U5541 (N_5541,N_4743,N_4240);
nor U5542 (N_5542,N_4169,N_4288);
and U5543 (N_5543,N_4576,N_4640);
nand U5544 (N_5544,N_4501,N_4586);
or U5545 (N_5545,N_4652,N_4661);
nand U5546 (N_5546,N_4367,N_4600);
or U5547 (N_5547,N_4665,N_4545);
and U5548 (N_5548,N_4497,N_4326);
xnor U5549 (N_5549,N_4584,N_4953);
or U5550 (N_5550,N_4233,N_4058);
xor U5551 (N_5551,N_4082,N_4435);
and U5552 (N_5552,N_4994,N_4024);
nand U5553 (N_5553,N_4340,N_4788);
and U5554 (N_5554,N_4674,N_4792);
and U5555 (N_5555,N_4356,N_4122);
or U5556 (N_5556,N_4502,N_4307);
or U5557 (N_5557,N_4850,N_4752);
nor U5558 (N_5558,N_4764,N_4303);
nand U5559 (N_5559,N_4783,N_4517);
and U5560 (N_5560,N_4781,N_4440);
xnor U5561 (N_5561,N_4762,N_4481);
nand U5562 (N_5562,N_4297,N_4506);
xnor U5563 (N_5563,N_4196,N_4680);
nor U5564 (N_5564,N_4910,N_4968);
nand U5565 (N_5565,N_4391,N_4940);
xor U5566 (N_5566,N_4989,N_4055);
or U5567 (N_5567,N_4265,N_4790);
nand U5568 (N_5568,N_4128,N_4122);
nand U5569 (N_5569,N_4359,N_4865);
or U5570 (N_5570,N_4665,N_4888);
nor U5571 (N_5571,N_4437,N_4593);
nand U5572 (N_5572,N_4629,N_4055);
or U5573 (N_5573,N_4819,N_4789);
or U5574 (N_5574,N_4152,N_4492);
nand U5575 (N_5575,N_4881,N_4113);
xnor U5576 (N_5576,N_4643,N_4126);
or U5577 (N_5577,N_4419,N_4966);
nor U5578 (N_5578,N_4111,N_4073);
and U5579 (N_5579,N_4962,N_4292);
and U5580 (N_5580,N_4399,N_4691);
or U5581 (N_5581,N_4569,N_4117);
nor U5582 (N_5582,N_4705,N_4106);
and U5583 (N_5583,N_4016,N_4751);
nor U5584 (N_5584,N_4183,N_4315);
nand U5585 (N_5585,N_4493,N_4701);
or U5586 (N_5586,N_4496,N_4654);
or U5587 (N_5587,N_4609,N_4895);
nand U5588 (N_5588,N_4936,N_4241);
xnor U5589 (N_5589,N_4663,N_4209);
and U5590 (N_5590,N_4428,N_4469);
and U5591 (N_5591,N_4954,N_4369);
and U5592 (N_5592,N_4480,N_4429);
or U5593 (N_5593,N_4937,N_4691);
nor U5594 (N_5594,N_4587,N_4255);
or U5595 (N_5595,N_4181,N_4301);
or U5596 (N_5596,N_4896,N_4011);
and U5597 (N_5597,N_4603,N_4156);
or U5598 (N_5598,N_4125,N_4617);
and U5599 (N_5599,N_4309,N_4626);
and U5600 (N_5600,N_4944,N_4127);
nor U5601 (N_5601,N_4062,N_4090);
and U5602 (N_5602,N_4959,N_4526);
and U5603 (N_5603,N_4635,N_4898);
nand U5604 (N_5604,N_4199,N_4109);
and U5605 (N_5605,N_4350,N_4947);
nand U5606 (N_5606,N_4478,N_4185);
nand U5607 (N_5607,N_4858,N_4228);
nand U5608 (N_5608,N_4416,N_4943);
or U5609 (N_5609,N_4379,N_4777);
and U5610 (N_5610,N_4311,N_4257);
or U5611 (N_5611,N_4252,N_4985);
and U5612 (N_5612,N_4112,N_4017);
and U5613 (N_5613,N_4504,N_4233);
and U5614 (N_5614,N_4132,N_4643);
or U5615 (N_5615,N_4109,N_4981);
and U5616 (N_5616,N_4168,N_4594);
and U5617 (N_5617,N_4342,N_4473);
nand U5618 (N_5618,N_4713,N_4187);
and U5619 (N_5619,N_4051,N_4162);
or U5620 (N_5620,N_4027,N_4492);
and U5621 (N_5621,N_4490,N_4673);
xnor U5622 (N_5622,N_4089,N_4474);
nor U5623 (N_5623,N_4125,N_4882);
nand U5624 (N_5624,N_4052,N_4906);
xor U5625 (N_5625,N_4223,N_4641);
or U5626 (N_5626,N_4497,N_4675);
nand U5627 (N_5627,N_4606,N_4513);
or U5628 (N_5628,N_4245,N_4427);
nand U5629 (N_5629,N_4659,N_4344);
nor U5630 (N_5630,N_4816,N_4214);
nand U5631 (N_5631,N_4142,N_4051);
nor U5632 (N_5632,N_4522,N_4900);
and U5633 (N_5633,N_4413,N_4808);
nor U5634 (N_5634,N_4209,N_4232);
nand U5635 (N_5635,N_4404,N_4643);
or U5636 (N_5636,N_4894,N_4135);
or U5637 (N_5637,N_4256,N_4742);
nand U5638 (N_5638,N_4835,N_4232);
and U5639 (N_5639,N_4625,N_4180);
nand U5640 (N_5640,N_4056,N_4359);
nand U5641 (N_5641,N_4898,N_4781);
and U5642 (N_5642,N_4146,N_4006);
or U5643 (N_5643,N_4807,N_4598);
nand U5644 (N_5644,N_4724,N_4607);
nand U5645 (N_5645,N_4020,N_4923);
and U5646 (N_5646,N_4771,N_4295);
nor U5647 (N_5647,N_4635,N_4983);
nand U5648 (N_5648,N_4725,N_4773);
or U5649 (N_5649,N_4255,N_4347);
nor U5650 (N_5650,N_4597,N_4426);
nand U5651 (N_5651,N_4135,N_4430);
and U5652 (N_5652,N_4523,N_4778);
nor U5653 (N_5653,N_4163,N_4687);
or U5654 (N_5654,N_4846,N_4662);
nand U5655 (N_5655,N_4920,N_4292);
and U5656 (N_5656,N_4733,N_4311);
and U5657 (N_5657,N_4190,N_4379);
or U5658 (N_5658,N_4279,N_4005);
and U5659 (N_5659,N_4978,N_4020);
and U5660 (N_5660,N_4130,N_4475);
and U5661 (N_5661,N_4265,N_4551);
nor U5662 (N_5662,N_4959,N_4505);
and U5663 (N_5663,N_4688,N_4422);
or U5664 (N_5664,N_4942,N_4176);
or U5665 (N_5665,N_4486,N_4783);
and U5666 (N_5666,N_4506,N_4917);
or U5667 (N_5667,N_4626,N_4323);
nor U5668 (N_5668,N_4791,N_4536);
and U5669 (N_5669,N_4020,N_4953);
nand U5670 (N_5670,N_4616,N_4600);
nor U5671 (N_5671,N_4740,N_4852);
and U5672 (N_5672,N_4517,N_4162);
or U5673 (N_5673,N_4490,N_4482);
or U5674 (N_5674,N_4056,N_4673);
nand U5675 (N_5675,N_4461,N_4286);
and U5676 (N_5676,N_4586,N_4043);
and U5677 (N_5677,N_4911,N_4948);
and U5678 (N_5678,N_4467,N_4698);
and U5679 (N_5679,N_4086,N_4762);
nor U5680 (N_5680,N_4776,N_4066);
or U5681 (N_5681,N_4615,N_4976);
and U5682 (N_5682,N_4435,N_4462);
nand U5683 (N_5683,N_4277,N_4852);
and U5684 (N_5684,N_4778,N_4850);
or U5685 (N_5685,N_4520,N_4631);
nor U5686 (N_5686,N_4483,N_4094);
xnor U5687 (N_5687,N_4359,N_4463);
nor U5688 (N_5688,N_4099,N_4390);
nand U5689 (N_5689,N_4524,N_4157);
nand U5690 (N_5690,N_4574,N_4632);
nand U5691 (N_5691,N_4802,N_4370);
or U5692 (N_5692,N_4397,N_4298);
and U5693 (N_5693,N_4804,N_4302);
or U5694 (N_5694,N_4956,N_4188);
nand U5695 (N_5695,N_4671,N_4829);
nand U5696 (N_5696,N_4142,N_4863);
or U5697 (N_5697,N_4021,N_4984);
or U5698 (N_5698,N_4373,N_4094);
nand U5699 (N_5699,N_4725,N_4627);
nor U5700 (N_5700,N_4190,N_4201);
and U5701 (N_5701,N_4877,N_4348);
and U5702 (N_5702,N_4124,N_4145);
and U5703 (N_5703,N_4285,N_4481);
nand U5704 (N_5704,N_4870,N_4860);
nor U5705 (N_5705,N_4144,N_4255);
and U5706 (N_5706,N_4396,N_4067);
or U5707 (N_5707,N_4748,N_4975);
nand U5708 (N_5708,N_4354,N_4423);
nor U5709 (N_5709,N_4017,N_4146);
nor U5710 (N_5710,N_4469,N_4055);
or U5711 (N_5711,N_4634,N_4891);
nor U5712 (N_5712,N_4289,N_4855);
nor U5713 (N_5713,N_4000,N_4838);
or U5714 (N_5714,N_4865,N_4535);
xnor U5715 (N_5715,N_4953,N_4398);
nand U5716 (N_5716,N_4680,N_4117);
and U5717 (N_5717,N_4744,N_4422);
and U5718 (N_5718,N_4091,N_4759);
nor U5719 (N_5719,N_4901,N_4350);
or U5720 (N_5720,N_4635,N_4407);
and U5721 (N_5721,N_4014,N_4212);
nand U5722 (N_5722,N_4953,N_4208);
or U5723 (N_5723,N_4273,N_4766);
nand U5724 (N_5724,N_4433,N_4336);
or U5725 (N_5725,N_4150,N_4421);
nand U5726 (N_5726,N_4469,N_4771);
and U5727 (N_5727,N_4944,N_4270);
or U5728 (N_5728,N_4461,N_4570);
xnor U5729 (N_5729,N_4366,N_4896);
nand U5730 (N_5730,N_4562,N_4700);
or U5731 (N_5731,N_4339,N_4800);
nand U5732 (N_5732,N_4368,N_4161);
xnor U5733 (N_5733,N_4811,N_4301);
nor U5734 (N_5734,N_4427,N_4151);
or U5735 (N_5735,N_4908,N_4136);
nor U5736 (N_5736,N_4456,N_4384);
or U5737 (N_5737,N_4475,N_4372);
or U5738 (N_5738,N_4733,N_4652);
nand U5739 (N_5739,N_4399,N_4100);
nand U5740 (N_5740,N_4980,N_4668);
and U5741 (N_5741,N_4339,N_4910);
nor U5742 (N_5742,N_4415,N_4780);
xor U5743 (N_5743,N_4122,N_4640);
and U5744 (N_5744,N_4017,N_4258);
nand U5745 (N_5745,N_4386,N_4106);
and U5746 (N_5746,N_4095,N_4331);
and U5747 (N_5747,N_4128,N_4712);
xor U5748 (N_5748,N_4735,N_4612);
or U5749 (N_5749,N_4240,N_4626);
and U5750 (N_5750,N_4207,N_4569);
and U5751 (N_5751,N_4493,N_4835);
nand U5752 (N_5752,N_4995,N_4831);
or U5753 (N_5753,N_4260,N_4183);
nand U5754 (N_5754,N_4808,N_4691);
nor U5755 (N_5755,N_4522,N_4576);
or U5756 (N_5756,N_4472,N_4440);
or U5757 (N_5757,N_4748,N_4290);
and U5758 (N_5758,N_4404,N_4125);
xor U5759 (N_5759,N_4492,N_4907);
and U5760 (N_5760,N_4245,N_4270);
and U5761 (N_5761,N_4482,N_4733);
and U5762 (N_5762,N_4115,N_4183);
nor U5763 (N_5763,N_4814,N_4681);
nor U5764 (N_5764,N_4430,N_4355);
or U5765 (N_5765,N_4675,N_4251);
nand U5766 (N_5766,N_4816,N_4738);
and U5767 (N_5767,N_4555,N_4086);
or U5768 (N_5768,N_4407,N_4491);
nor U5769 (N_5769,N_4408,N_4376);
or U5770 (N_5770,N_4393,N_4157);
and U5771 (N_5771,N_4714,N_4391);
nand U5772 (N_5772,N_4107,N_4377);
and U5773 (N_5773,N_4125,N_4043);
xor U5774 (N_5774,N_4732,N_4077);
and U5775 (N_5775,N_4076,N_4360);
and U5776 (N_5776,N_4210,N_4076);
nand U5777 (N_5777,N_4873,N_4467);
and U5778 (N_5778,N_4532,N_4030);
or U5779 (N_5779,N_4175,N_4425);
nor U5780 (N_5780,N_4702,N_4746);
nor U5781 (N_5781,N_4539,N_4449);
and U5782 (N_5782,N_4103,N_4368);
nor U5783 (N_5783,N_4848,N_4980);
nor U5784 (N_5784,N_4339,N_4512);
nor U5785 (N_5785,N_4643,N_4355);
nand U5786 (N_5786,N_4517,N_4229);
nor U5787 (N_5787,N_4716,N_4872);
nor U5788 (N_5788,N_4574,N_4799);
nand U5789 (N_5789,N_4480,N_4462);
nand U5790 (N_5790,N_4441,N_4128);
nor U5791 (N_5791,N_4024,N_4318);
nor U5792 (N_5792,N_4060,N_4019);
and U5793 (N_5793,N_4599,N_4201);
xnor U5794 (N_5794,N_4177,N_4862);
and U5795 (N_5795,N_4695,N_4396);
nand U5796 (N_5796,N_4935,N_4343);
xnor U5797 (N_5797,N_4665,N_4741);
and U5798 (N_5798,N_4342,N_4607);
nand U5799 (N_5799,N_4505,N_4896);
nand U5800 (N_5800,N_4989,N_4908);
nand U5801 (N_5801,N_4955,N_4364);
nor U5802 (N_5802,N_4165,N_4213);
or U5803 (N_5803,N_4418,N_4388);
nor U5804 (N_5804,N_4939,N_4392);
and U5805 (N_5805,N_4108,N_4724);
and U5806 (N_5806,N_4123,N_4329);
nor U5807 (N_5807,N_4720,N_4885);
nor U5808 (N_5808,N_4089,N_4556);
or U5809 (N_5809,N_4764,N_4722);
or U5810 (N_5810,N_4772,N_4594);
nor U5811 (N_5811,N_4752,N_4737);
and U5812 (N_5812,N_4019,N_4360);
or U5813 (N_5813,N_4629,N_4517);
xor U5814 (N_5814,N_4760,N_4585);
or U5815 (N_5815,N_4986,N_4563);
or U5816 (N_5816,N_4174,N_4077);
or U5817 (N_5817,N_4180,N_4291);
xnor U5818 (N_5818,N_4173,N_4210);
nor U5819 (N_5819,N_4322,N_4835);
nor U5820 (N_5820,N_4751,N_4504);
nor U5821 (N_5821,N_4804,N_4444);
xor U5822 (N_5822,N_4429,N_4059);
nor U5823 (N_5823,N_4650,N_4428);
and U5824 (N_5824,N_4609,N_4361);
nand U5825 (N_5825,N_4947,N_4030);
and U5826 (N_5826,N_4095,N_4267);
nor U5827 (N_5827,N_4851,N_4239);
or U5828 (N_5828,N_4286,N_4070);
nand U5829 (N_5829,N_4996,N_4075);
and U5830 (N_5830,N_4014,N_4260);
nand U5831 (N_5831,N_4551,N_4959);
xnor U5832 (N_5832,N_4612,N_4174);
and U5833 (N_5833,N_4972,N_4535);
xor U5834 (N_5834,N_4755,N_4925);
and U5835 (N_5835,N_4250,N_4794);
or U5836 (N_5836,N_4250,N_4087);
and U5837 (N_5837,N_4971,N_4527);
nor U5838 (N_5838,N_4726,N_4623);
nor U5839 (N_5839,N_4254,N_4874);
or U5840 (N_5840,N_4132,N_4027);
nor U5841 (N_5841,N_4379,N_4497);
or U5842 (N_5842,N_4699,N_4837);
nor U5843 (N_5843,N_4464,N_4198);
or U5844 (N_5844,N_4019,N_4096);
or U5845 (N_5845,N_4147,N_4758);
nand U5846 (N_5846,N_4586,N_4987);
and U5847 (N_5847,N_4494,N_4555);
or U5848 (N_5848,N_4101,N_4352);
nand U5849 (N_5849,N_4647,N_4428);
nor U5850 (N_5850,N_4984,N_4652);
nor U5851 (N_5851,N_4089,N_4622);
or U5852 (N_5852,N_4896,N_4094);
and U5853 (N_5853,N_4392,N_4849);
nor U5854 (N_5854,N_4931,N_4336);
xor U5855 (N_5855,N_4957,N_4017);
nand U5856 (N_5856,N_4606,N_4945);
nor U5857 (N_5857,N_4380,N_4802);
or U5858 (N_5858,N_4707,N_4054);
nor U5859 (N_5859,N_4454,N_4683);
nand U5860 (N_5860,N_4244,N_4340);
and U5861 (N_5861,N_4093,N_4148);
or U5862 (N_5862,N_4697,N_4725);
nor U5863 (N_5863,N_4265,N_4997);
and U5864 (N_5864,N_4538,N_4435);
and U5865 (N_5865,N_4774,N_4484);
nor U5866 (N_5866,N_4576,N_4097);
nor U5867 (N_5867,N_4545,N_4167);
nor U5868 (N_5868,N_4881,N_4680);
or U5869 (N_5869,N_4933,N_4440);
nand U5870 (N_5870,N_4685,N_4936);
xnor U5871 (N_5871,N_4786,N_4195);
and U5872 (N_5872,N_4250,N_4974);
nand U5873 (N_5873,N_4815,N_4459);
and U5874 (N_5874,N_4998,N_4714);
and U5875 (N_5875,N_4227,N_4876);
xnor U5876 (N_5876,N_4499,N_4855);
xor U5877 (N_5877,N_4543,N_4367);
nand U5878 (N_5878,N_4862,N_4194);
and U5879 (N_5879,N_4298,N_4370);
nor U5880 (N_5880,N_4361,N_4455);
or U5881 (N_5881,N_4932,N_4484);
and U5882 (N_5882,N_4783,N_4488);
nor U5883 (N_5883,N_4283,N_4567);
nand U5884 (N_5884,N_4262,N_4198);
xor U5885 (N_5885,N_4709,N_4749);
nand U5886 (N_5886,N_4011,N_4467);
and U5887 (N_5887,N_4594,N_4190);
nor U5888 (N_5888,N_4239,N_4587);
nor U5889 (N_5889,N_4412,N_4975);
nand U5890 (N_5890,N_4307,N_4306);
and U5891 (N_5891,N_4583,N_4356);
nor U5892 (N_5892,N_4303,N_4605);
nand U5893 (N_5893,N_4672,N_4746);
xnor U5894 (N_5894,N_4068,N_4059);
xor U5895 (N_5895,N_4228,N_4160);
or U5896 (N_5896,N_4691,N_4594);
or U5897 (N_5897,N_4207,N_4508);
and U5898 (N_5898,N_4613,N_4731);
xor U5899 (N_5899,N_4167,N_4828);
nand U5900 (N_5900,N_4224,N_4154);
xor U5901 (N_5901,N_4157,N_4742);
nor U5902 (N_5902,N_4701,N_4619);
and U5903 (N_5903,N_4437,N_4170);
nor U5904 (N_5904,N_4918,N_4882);
nand U5905 (N_5905,N_4695,N_4274);
nor U5906 (N_5906,N_4656,N_4651);
nor U5907 (N_5907,N_4323,N_4253);
and U5908 (N_5908,N_4337,N_4202);
and U5909 (N_5909,N_4777,N_4649);
xor U5910 (N_5910,N_4560,N_4364);
nor U5911 (N_5911,N_4895,N_4001);
or U5912 (N_5912,N_4638,N_4002);
nand U5913 (N_5913,N_4869,N_4895);
and U5914 (N_5914,N_4087,N_4258);
or U5915 (N_5915,N_4588,N_4708);
and U5916 (N_5916,N_4372,N_4082);
nor U5917 (N_5917,N_4930,N_4803);
and U5918 (N_5918,N_4367,N_4098);
nand U5919 (N_5919,N_4049,N_4100);
nand U5920 (N_5920,N_4837,N_4392);
nand U5921 (N_5921,N_4305,N_4998);
or U5922 (N_5922,N_4797,N_4131);
nor U5923 (N_5923,N_4276,N_4004);
nor U5924 (N_5924,N_4737,N_4779);
xnor U5925 (N_5925,N_4877,N_4003);
xnor U5926 (N_5926,N_4289,N_4582);
or U5927 (N_5927,N_4250,N_4005);
or U5928 (N_5928,N_4950,N_4565);
nor U5929 (N_5929,N_4690,N_4457);
nand U5930 (N_5930,N_4152,N_4971);
and U5931 (N_5931,N_4578,N_4575);
or U5932 (N_5932,N_4263,N_4242);
nor U5933 (N_5933,N_4848,N_4206);
nand U5934 (N_5934,N_4435,N_4879);
nor U5935 (N_5935,N_4396,N_4325);
and U5936 (N_5936,N_4198,N_4946);
nor U5937 (N_5937,N_4940,N_4887);
and U5938 (N_5938,N_4400,N_4013);
nand U5939 (N_5939,N_4099,N_4349);
nor U5940 (N_5940,N_4641,N_4329);
and U5941 (N_5941,N_4219,N_4003);
or U5942 (N_5942,N_4178,N_4176);
nor U5943 (N_5943,N_4921,N_4150);
nor U5944 (N_5944,N_4208,N_4957);
or U5945 (N_5945,N_4306,N_4404);
nand U5946 (N_5946,N_4927,N_4524);
xnor U5947 (N_5947,N_4978,N_4265);
nor U5948 (N_5948,N_4143,N_4384);
and U5949 (N_5949,N_4893,N_4425);
nor U5950 (N_5950,N_4828,N_4496);
nand U5951 (N_5951,N_4217,N_4559);
or U5952 (N_5952,N_4081,N_4866);
and U5953 (N_5953,N_4261,N_4356);
or U5954 (N_5954,N_4730,N_4335);
xor U5955 (N_5955,N_4094,N_4183);
nor U5956 (N_5956,N_4990,N_4250);
and U5957 (N_5957,N_4750,N_4447);
or U5958 (N_5958,N_4285,N_4787);
xor U5959 (N_5959,N_4159,N_4519);
nand U5960 (N_5960,N_4835,N_4354);
xor U5961 (N_5961,N_4783,N_4051);
or U5962 (N_5962,N_4372,N_4440);
or U5963 (N_5963,N_4395,N_4280);
nor U5964 (N_5964,N_4183,N_4480);
and U5965 (N_5965,N_4108,N_4761);
nand U5966 (N_5966,N_4379,N_4805);
xnor U5967 (N_5967,N_4640,N_4860);
nor U5968 (N_5968,N_4222,N_4159);
and U5969 (N_5969,N_4105,N_4696);
or U5970 (N_5970,N_4473,N_4135);
nor U5971 (N_5971,N_4344,N_4005);
nor U5972 (N_5972,N_4662,N_4967);
or U5973 (N_5973,N_4896,N_4408);
and U5974 (N_5974,N_4308,N_4474);
nand U5975 (N_5975,N_4148,N_4114);
nand U5976 (N_5976,N_4810,N_4236);
nor U5977 (N_5977,N_4463,N_4245);
xor U5978 (N_5978,N_4894,N_4021);
nor U5979 (N_5979,N_4136,N_4827);
and U5980 (N_5980,N_4074,N_4273);
or U5981 (N_5981,N_4968,N_4387);
nor U5982 (N_5982,N_4526,N_4296);
or U5983 (N_5983,N_4814,N_4870);
or U5984 (N_5984,N_4986,N_4160);
or U5985 (N_5985,N_4485,N_4697);
or U5986 (N_5986,N_4288,N_4209);
and U5987 (N_5987,N_4027,N_4048);
or U5988 (N_5988,N_4872,N_4307);
or U5989 (N_5989,N_4696,N_4258);
nor U5990 (N_5990,N_4712,N_4555);
nand U5991 (N_5991,N_4698,N_4647);
and U5992 (N_5992,N_4185,N_4956);
or U5993 (N_5993,N_4223,N_4246);
or U5994 (N_5994,N_4482,N_4163);
nand U5995 (N_5995,N_4539,N_4973);
and U5996 (N_5996,N_4816,N_4508);
or U5997 (N_5997,N_4269,N_4231);
nand U5998 (N_5998,N_4601,N_4857);
nor U5999 (N_5999,N_4736,N_4310);
or U6000 (N_6000,N_5047,N_5026);
xnor U6001 (N_6001,N_5821,N_5570);
nor U6002 (N_6002,N_5660,N_5860);
and U6003 (N_6003,N_5842,N_5094);
or U6004 (N_6004,N_5087,N_5925);
and U6005 (N_6005,N_5033,N_5136);
and U6006 (N_6006,N_5484,N_5974);
nor U6007 (N_6007,N_5084,N_5099);
xnor U6008 (N_6008,N_5778,N_5269);
or U6009 (N_6009,N_5317,N_5984);
or U6010 (N_6010,N_5780,N_5729);
nand U6011 (N_6011,N_5332,N_5196);
and U6012 (N_6012,N_5478,N_5315);
nand U6013 (N_6013,N_5189,N_5472);
nor U6014 (N_6014,N_5384,N_5572);
nand U6015 (N_6015,N_5085,N_5641);
nand U6016 (N_6016,N_5093,N_5683);
and U6017 (N_6017,N_5951,N_5068);
and U6018 (N_6018,N_5468,N_5635);
and U6019 (N_6019,N_5993,N_5637);
and U6020 (N_6020,N_5413,N_5682);
or U6021 (N_6021,N_5278,N_5333);
nand U6022 (N_6022,N_5091,N_5724);
or U6023 (N_6023,N_5012,N_5175);
nor U6024 (N_6024,N_5814,N_5446);
or U6025 (N_6025,N_5098,N_5289);
xnor U6026 (N_6026,N_5751,N_5082);
nor U6027 (N_6027,N_5710,N_5545);
nor U6028 (N_6028,N_5907,N_5146);
nand U6029 (N_6029,N_5030,N_5688);
nor U6030 (N_6030,N_5133,N_5777);
or U6031 (N_6031,N_5941,N_5104);
nand U6032 (N_6032,N_5153,N_5251);
nor U6033 (N_6033,N_5743,N_5198);
or U6034 (N_6034,N_5161,N_5308);
nor U6035 (N_6035,N_5767,N_5071);
or U6036 (N_6036,N_5523,N_5281);
nor U6037 (N_6037,N_5915,N_5550);
xor U6038 (N_6038,N_5272,N_5488);
and U6039 (N_6039,N_5326,N_5676);
xor U6040 (N_6040,N_5638,N_5952);
nand U6041 (N_6041,N_5687,N_5748);
nor U6042 (N_6042,N_5843,N_5540);
nor U6043 (N_6043,N_5385,N_5311);
nor U6044 (N_6044,N_5874,N_5669);
nand U6045 (N_6045,N_5116,N_5790);
nor U6046 (N_6046,N_5896,N_5036);
and U6047 (N_6047,N_5018,N_5188);
nand U6048 (N_6048,N_5969,N_5256);
or U6049 (N_6049,N_5931,N_5728);
nor U6050 (N_6050,N_5906,N_5782);
nand U6051 (N_6051,N_5062,N_5788);
nor U6052 (N_6052,N_5159,N_5422);
nand U6053 (N_6053,N_5863,N_5578);
nor U6054 (N_6054,N_5861,N_5849);
nor U6055 (N_6055,N_5519,N_5636);
nand U6056 (N_6056,N_5648,N_5978);
xnor U6057 (N_6057,N_5869,N_5428);
nor U6058 (N_6058,N_5988,N_5998);
nor U6059 (N_6059,N_5194,N_5190);
and U6060 (N_6060,N_5866,N_5061);
nand U6061 (N_6061,N_5096,N_5742);
xor U6062 (N_6062,N_5327,N_5177);
nor U6063 (N_6063,N_5890,N_5054);
xor U6064 (N_6064,N_5912,N_5409);
and U6065 (N_6065,N_5297,N_5926);
and U6066 (N_6066,N_5427,N_5028);
nand U6067 (N_6067,N_5264,N_5608);
nor U6068 (N_6068,N_5110,N_5704);
and U6069 (N_6069,N_5548,N_5711);
and U6070 (N_6070,N_5368,N_5474);
xnor U6071 (N_6071,N_5496,N_5661);
nand U6072 (N_6072,N_5070,N_5822);
and U6073 (N_6073,N_5986,N_5838);
xnor U6074 (N_6074,N_5255,N_5049);
and U6075 (N_6075,N_5663,N_5835);
and U6076 (N_6076,N_5508,N_5217);
or U6077 (N_6077,N_5485,N_5078);
and U6078 (N_6078,N_5749,N_5574);
nor U6079 (N_6079,N_5832,N_5075);
nor U6080 (N_6080,N_5000,N_5817);
nor U6081 (N_6081,N_5740,N_5919);
xnor U6082 (N_6082,N_5666,N_5065);
and U6083 (N_6083,N_5122,N_5921);
or U6084 (N_6084,N_5802,N_5199);
or U6085 (N_6085,N_5873,N_5050);
and U6086 (N_6086,N_5219,N_5557);
or U6087 (N_6087,N_5195,N_5363);
and U6088 (N_6088,N_5418,N_5544);
or U6089 (N_6089,N_5909,N_5871);
nor U6090 (N_6090,N_5567,N_5505);
and U6091 (N_6091,N_5733,N_5492);
nand U6092 (N_6092,N_5744,N_5376);
nor U6093 (N_6093,N_5825,N_5481);
and U6094 (N_6094,N_5577,N_5373);
and U6095 (N_6095,N_5365,N_5980);
nor U6096 (N_6096,N_5059,N_5725);
nor U6097 (N_6097,N_5552,N_5690);
and U6098 (N_6098,N_5149,N_5214);
xor U6099 (N_6099,N_5207,N_5918);
and U6100 (N_6100,N_5282,N_5714);
and U6101 (N_6101,N_5223,N_5105);
nand U6102 (N_6102,N_5148,N_5715);
and U6103 (N_6103,N_5302,N_5312);
or U6104 (N_6104,N_5045,N_5003);
and U6105 (N_6105,N_5979,N_5722);
and U6106 (N_6106,N_5445,N_5417);
and U6107 (N_6107,N_5609,N_5304);
xor U6108 (N_6108,N_5820,N_5526);
or U6109 (N_6109,N_5250,N_5670);
nor U6110 (N_6110,N_5518,N_5364);
and U6111 (N_6111,N_5855,N_5181);
nor U6112 (N_6112,N_5348,N_5537);
and U6113 (N_6113,N_5447,N_5450);
nand U6114 (N_6114,N_5453,N_5610);
xor U6115 (N_6115,N_5144,N_5953);
xor U6116 (N_6116,N_5624,N_5513);
nor U6117 (N_6117,N_5593,N_5757);
or U6118 (N_6118,N_5386,N_5996);
nand U6119 (N_6119,N_5032,N_5463);
or U6120 (N_6120,N_5095,N_5007);
nor U6121 (N_6121,N_5631,N_5839);
xor U6122 (N_6122,N_5206,N_5827);
nand U6123 (N_6123,N_5170,N_5604);
nand U6124 (N_6124,N_5872,N_5039);
nor U6125 (N_6125,N_5657,N_5703);
xnor U6126 (N_6126,N_5948,N_5210);
and U6127 (N_6127,N_5625,N_5868);
nand U6128 (N_6128,N_5156,N_5423);
and U6129 (N_6129,N_5656,N_5237);
or U6130 (N_6130,N_5811,N_5647);
and U6131 (N_6131,N_5880,N_5718);
nand U6132 (N_6132,N_5720,N_5841);
nand U6133 (N_6133,N_5081,N_5727);
nor U6134 (N_6134,N_5960,N_5726);
nor U6135 (N_6135,N_5753,N_5784);
nor U6136 (N_6136,N_5112,N_5746);
nor U6137 (N_6137,N_5142,N_5069);
nor U6138 (N_6138,N_5213,N_5789);
nand U6139 (N_6139,N_5329,N_5247);
nor U6140 (N_6140,N_5920,N_5686);
or U6141 (N_6141,N_5245,N_5949);
and U6142 (N_6142,N_5419,N_5038);
or U6143 (N_6143,N_5296,N_5367);
xnor U6144 (N_6144,N_5435,N_5125);
and U6145 (N_6145,N_5933,N_5138);
nor U6146 (N_6146,N_5893,N_5056);
nand U6147 (N_6147,N_5566,N_5944);
and U6148 (N_6148,N_5897,N_5322);
nand U6149 (N_6149,N_5037,N_5774);
nor U6150 (N_6150,N_5318,N_5731);
nand U6151 (N_6151,N_5233,N_5950);
and U6152 (N_6152,N_5954,N_5225);
nand U6153 (N_6153,N_5180,N_5187);
nand U6154 (N_6154,N_5515,N_5712);
or U6155 (N_6155,N_5975,N_5354);
and U6156 (N_6156,N_5590,N_5168);
and U6157 (N_6157,N_5303,N_5917);
nand U6158 (N_6158,N_5380,N_5286);
or U6159 (N_6159,N_5027,N_5306);
xor U6160 (N_6160,N_5378,N_5414);
nor U6161 (N_6161,N_5004,N_5929);
nor U6162 (N_6162,N_5394,N_5623);
nand U6163 (N_6163,N_5211,N_5005);
or U6164 (N_6164,N_5534,N_5536);
xnor U6165 (N_6165,N_5891,N_5410);
or U6166 (N_6166,N_5645,N_5695);
nand U6167 (N_6167,N_5400,N_5372);
xor U6168 (N_6168,N_5227,N_5791);
or U6169 (N_6169,N_5330,N_5503);
and U6170 (N_6170,N_5852,N_5080);
or U6171 (N_6171,N_5582,N_5216);
and U6172 (N_6172,N_5800,N_5076);
nor U6173 (N_6173,N_5491,N_5309);
or U6174 (N_6174,N_5338,N_5232);
nand U6175 (N_6175,N_5618,N_5815);
and U6176 (N_6176,N_5416,N_5246);
or U6177 (N_6177,N_5430,N_5215);
nor U6178 (N_6178,N_5653,N_5809);
or U6179 (N_6179,N_5458,N_5983);
and U6180 (N_6180,N_5730,N_5797);
nand U6181 (N_6181,N_5597,N_5183);
or U6182 (N_6182,N_5339,N_5292);
xnor U6183 (N_6183,N_5875,N_5088);
or U6184 (N_6184,N_5139,N_5575);
nand U6185 (N_6185,N_5239,N_5259);
or U6186 (N_6186,N_5353,N_5429);
and U6187 (N_6187,N_5383,N_5600);
and U6188 (N_6188,N_5531,N_5114);
nand U6189 (N_6189,N_5379,N_5796);
or U6190 (N_6190,N_5799,N_5514);
and U6191 (N_6191,N_5109,N_5524);
and U6192 (N_6192,N_5019,N_5443);
or U6193 (N_6193,N_5222,N_5500);
and U6194 (N_6194,N_5375,N_5313);
nand U6195 (N_6195,N_5042,N_5763);
xor U6196 (N_6196,N_5958,N_5280);
nand U6197 (N_6197,N_5585,N_5164);
xor U6198 (N_6198,N_5197,N_5990);
and U6199 (N_6199,N_5620,N_5779);
nand U6200 (N_6200,N_5675,N_5671);
nor U6201 (N_6201,N_5111,N_5204);
nand U6202 (N_6202,N_5632,N_5684);
nand U6203 (N_6203,N_5209,N_5685);
nor U6204 (N_6204,N_5659,N_5846);
nor U6205 (N_6205,N_5619,N_5321);
nor U6206 (N_6206,N_5963,N_5977);
xnor U6207 (N_6207,N_5141,N_5258);
nand U6208 (N_6208,N_5421,N_5499);
or U6209 (N_6209,N_5399,N_5831);
nor U6210 (N_6210,N_5455,N_5626);
and U6211 (N_6211,N_5616,N_5323);
nor U6212 (N_6212,N_5016,N_5549);
nor U6213 (N_6213,N_5129,N_5274);
nand U6214 (N_6214,N_5760,N_5943);
or U6215 (N_6215,N_5457,N_5202);
nor U6216 (N_6216,N_5079,N_5127);
and U6217 (N_6217,N_5864,N_5178);
nor U6218 (N_6218,N_5436,N_5511);
nand U6219 (N_6219,N_5558,N_5654);
xor U6220 (N_6220,N_5271,N_5284);
nand U6221 (N_6221,N_5442,N_5693);
nor U6222 (N_6222,N_5203,N_5701);
nand U6223 (N_6223,N_5390,N_5449);
and U6224 (N_6224,N_5605,N_5762);
nor U6225 (N_6225,N_5073,N_5966);
nor U6226 (N_6226,N_5355,N_5147);
nor U6227 (N_6227,N_5781,N_5651);
and U6228 (N_6228,N_5089,N_5542);
nand U6229 (N_6229,N_5591,N_5432);
nor U6230 (N_6230,N_5930,N_5801);
nand U6231 (N_6231,N_5392,N_5408);
or U6232 (N_6232,N_5721,N_5658);
xor U6233 (N_6233,N_5291,N_5301);
nand U6234 (N_6234,N_5755,N_5900);
or U6235 (N_6235,N_5448,N_5561);
or U6236 (N_6236,N_5745,N_5667);
and U6237 (N_6237,N_5155,N_5451);
nor U6238 (N_6238,N_5962,N_5803);
or U6239 (N_6239,N_5100,N_5509);
and U6240 (N_6240,N_5220,N_5899);
and U6241 (N_6241,N_5381,N_5889);
or U6242 (N_6242,N_5571,N_5165);
nand U6243 (N_6243,N_5525,N_5783);
and U6244 (N_6244,N_5771,N_5504);
nor U6245 (N_6245,N_5342,N_5403);
and U6246 (N_6246,N_5169,N_5307);
nor U6247 (N_6247,N_5128,N_5288);
nand U6248 (N_6248,N_5924,N_5171);
nor U6249 (N_6249,N_5253,N_5847);
or U6250 (N_6250,N_5359,N_5927);
xor U6251 (N_6251,N_5011,N_5117);
and U6252 (N_6252,N_5521,N_5388);
xnor U6253 (N_6253,N_5260,N_5680);
nor U6254 (N_6254,N_5903,N_5193);
or U6255 (N_6255,N_5877,N_5241);
and U6256 (N_6256,N_5135,N_5738);
and U6257 (N_6257,N_5976,N_5614);
and U6258 (N_6258,N_5601,N_5853);
nand U6259 (N_6259,N_5512,N_5696);
and U6260 (N_6260,N_5476,N_5025);
nor U6261 (N_6261,N_5166,N_5997);
nand U6262 (N_6262,N_5101,N_5064);
and U6263 (N_6263,N_5287,N_5989);
nor U6264 (N_6264,N_5160,N_5218);
nand U6265 (N_6265,N_5603,N_5498);
nor U6266 (N_6266,N_5480,N_5533);
nand U6267 (N_6267,N_5756,N_5955);
xnor U6268 (N_6268,N_5629,N_5124);
or U6269 (N_6269,N_5857,N_5828);
xnor U6270 (N_6270,N_5946,N_5981);
nor U6271 (N_6271,N_5565,N_5358);
nand U6272 (N_6272,N_5140,N_5063);
nand U6273 (N_6273,N_5765,N_5876);
nor U6274 (N_6274,N_5794,N_5646);
nand U6275 (N_6275,N_5238,N_5606);
nor U6276 (N_6276,N_5664,N_5438);
or U6277 (N_6277,N_5973,N_5908);
or U6278 (N_6278,N_5581,N_5115);
or U6279 (N_6279,N_5126,N_5341);
nand U6280 (N_6280,N_5807,N_5810);
and U6281 (N_6281,N_5516,N_5477);
or U6282 (N_6282,N_5437,N_5460);
nand U6283 (N_6283,N_5034,N_5754);
nor U6284 (N_6284,N_5324,N_5404);
or U6285 (N_6285,N_5425,N_5356);
or U6286 (N_6286,N_5599,N_5957);
nand U6287 (N_6287,N_5834,N_5242);
or U6288 (N_6288,N_5556,N_5795);
nor U6289 (N_6289,N_5405,N_5072);
xor U6290 (N_6290,N_5895,N_5276);
and U6291 (N_6291,N_5885,N_5229);
and U6292 (N_6292,N_5490,N_5162);
and U6293 (N_6293,N_5475,N_5494);
and U6294 (N_6294,N_5179,N_5967);
nand U6295 (N_6295,N_5554,N_5299);
or U6296 (N_6296,N_5644,N_5887);
or U6297 (N_6297,N_5879,N_5888);
nor U6298 (N_6298,N_5634,N_5627);
and U6299 (N_6299,N_5611,N_5506);
xor U6300 (N_6300,N_5652,N_5560);
xnor U6301 (N_6301,N_5735,N_5569);
and U6302 (N_6302,N_5902,N_5649);
nor U6303 (N_6303,N_5923,N_5283);
nor U6304 (N_6304,N_5938,N_5439);
nor U6305 (N_6305,N_5267,N_5995);
nand U6306 (N_6306,N_5393,N_5830);
and U6307 (N_6307,N_5334,N_5639);
and U6308 (N_6308,N_5029,N_5497);
nand U6309 (N_6309,N_5699,N_5612);
and U6310 (N_6310,N_5357,N_5320);
nor U6311 (N_6311,N_5426,N_5185);
nand U6312 (N_6312,N_5407,N_5716);
or U6313 (N_6313,N_5679,N_5244);
or U6314 (N_6314,N_5462,N_5066);
and U6315 (N_6315,N_5633,N_5325);
and U6316 (N_6316,N_5243,N_5553);
nand U6317 (N_6317,N_5395,N_5910);
and U6318 (N_6318,N_5901,N_5048);
nand U6319 (N_6319,N_5013,N_5167);
nand U6320 (N_6320,N_5991,N_5184);
nand U6321 (N_6321,N_5719,N_5006);
or U6322 (N_6322,N_5773,N_5535);
or U6323 (N_6323,N_5502,N_5466);
or U6324 (N_6324,N_5522,N_5607);
nor U6325 (N_6325,N_5350,N_5904);
or U6326 (N_6326,N_5040,N_5401);
xnor U6327 (N_6327,N_5892,N_5086);
nand U6328 (N_6328,N_5792,N_5343);
nand U6329 (N_6329,N_5886,N_5495);
nand U6330 (N_6330,N_5798,N_5433);
or U6331 (N_6331,N_5236,N_5470);
nand U6332 (N_6332,N_5043,N_5362);
and U6333 (N_6333,N_5532,N_5444);
or U6334 (N_6334,N_5965,N_5224);
nand U6335 (N_6335,N_5833,N_5517);
or U6336 (N_6336,N_5226,N_5487);
xnor U6337 (N_6337,N_5389,N_5273);
and U6338 (N_6338,N_5878,N_5805);
and U6339 (N_6339,N_5120,N_5994);
and U6340 (N_6340,N_5482,N_5507);
and U6341 (N_6341,N_5622,N_5858);
or U6342 (N_6342,N_5102,N_5848);
nor U6343 (N_6343,N_5939,N_5415);
nor U6344 (N_6344,N_5583,N_5961);
and U6345 (N_6345,N_5576,N_5275);
xor U6346 (N_6346,N_5655,N_5052);
or U6347 (N_6347,N_5694,N_5008);
or U6348 (N_6348,N_5824,N_5461);
nand U6349 (N_6349,N_5192,N_5345);
or U6350 (N_6350,N_5741,N_5761);
nand U6351 (N_6351,N_5228,N_5999);
nand U6352 (N_6352,N_5083,N_5862);
and U6353 (N_6353,N_5440,N_5707);
nand U6354 (N_6354,N_5265,N_5884);
nor U6355 (N_6355,N_5713,N_5851);
nor U6356 (N_6356,N_5947,N_5022);
nand U6357 (N_6357,N_5053,N_5235);
xor U6358 (N_6358,N_5493,N_5739);
or U6359 (N_6359,N_5420,N_5252);
nor U6360 (N_6360,N_5382,N_5501);
nor U6361 (N_6361,N_5586,N_5617);
nor U6362 (N_6362,N_5592,N_5298);
or U6363 (N_6363,N_5881,N_5021);
and U6364 (N_6364,N_5650,N_5914);
and U6365 (N_6365,N_5543,N_5594);
and U6366 (N_6366,N_5369,N_5595);
nand U6367 (N_6367,N_5844,N_5826);
or U6368 (N_6368,N_5396,N_5121);
and U6369 (N_6369,N_5031,N_5257);
nor U6370 (N_6370,N_5674,N_5630);
nor U6371 (N_6371,N_5361,N_5691);
nor U6372 (N_6372,N_5060,N_5541);
or U6373 (N_6373,N_5922,N_5928);
xnor U6374 (N_6374,N_5151,N_5279);
nand U6375 (N_6375,N_5234,N_5563);
nand U6376 (N_6376,N_5568,N_5530);
or U6377 (N_6377,N_5935,N_5231);
xnor U6378 (N_6378,N_5732,N_5467);
nand U6379 (N_6379,N_5837,N_5208);
and U6380 (N_6380,N_5294,N_5240);
or U6381 (N_6381,N_5770,N_5551);
nand U6382 (N_6382,N_5854,N_5584);
and U6383 (N_6383,N_5776,N_5137);
and U6384 (N_6384,N_5894,N_5270);
xor U6385 (N_6385,N_5176,N_5046);
nand U6386 (N_6386,N_5559,N_5628);
and U6387 (N_6387,N_5263,N_5143);
nor U6388 (N_6388,N_5934,N_5845);
nand U6389 (N_6389,N_5248,N_5058);
nor U6390 (N_6390,N_5971,N_5035);
or U6391 (N_6391,N_5972,N_5009);
nor U6392 (N_6392,N_5806,N_5662);
and U6393 (N_6393,N_5057,N_5905);
nor U6394 (N_6394,N_5314,N_5692);
xor U6395 (N_6395,N_5898,N_5434);
or U6396 (N_6396,N_5172,N_5812);
nand U6397 (N_6397,N_5945,N_5374);
and U6398 (N_6398,N_5579,N_5793);
or U6399 (N_6399,N_5305,N_5103);
nor U6400 (N_6400,N_5402,N_5913);
or U6401 (N_6401,N_5459,N_5051);
nand U6402 (N_6402,N_5836,N_5829);
xnor U6403 (N_6403,N_5201,N_5107);
nand U6404 (N_6404,N_5883,N_5598);
nor U6405 (N_6405,N_5391,N_5668);
xor U6406 (N_6406,N_5564,N_5174);
and U6407 (N_6407,N_5527,N_5587);
xnor U6408 (N_6408,N_5775,N_5067);
xnor U6409 (N_6409,N_5336,N_5786);
nand U6410 (N_6410,N_5510,N_5615);
or U6411 (N_6411,N_5186,N_5596);
or U6412 (N_6412,N_5588,N_5677);
or U6413 (N_6413,N_5191,N_5131);
nor U6414 (N_6414,N_5772,N_5424);
xnor U6415 (N_6415,N_5766,N_5266);
and U6416 (N_6416,N_5486,N_5882);
or U6417 (N_6417,N_5471,N_5347);
or U6418 (N_6418,N_5473,N_5681);
or U6419 (N_6419,N_5759,N_5335);
nand U6420 (N_6420,N_5816,N_5818);
or U6421 (N_6421,N_5819,N_5340);
and U6422 (N_6422,N_5956,N_5200);
or U6423 (N_6423,N_5940,N_5916);
nand U6424 (N_6424,N_5001,N_5431);
nor U6425 (N_6425,N_5024,N_5539);
nor U6426 (N_6426,N_5665,N_5441);
and U6427 (N_6427,N_5709,N_5015);
nor U6428 (N_6428,N_5859,N_5787);
or U6429 (N_6429,N_5130,N_5092);
nand U6430 (N_6430,N_5483,N_5942);
and U6431 (N_6431,N_5736,N_5014);
xnor U6432 (N_6432,N_5708,N_5262);
or U6433 (N_6433,N_5173,N_5119);
and U6434 (N_6434,N_5589,N_5643);
nor U6435 (N_6435,N_5074,N_5529);
nand U6436 (N_6436,N_5163,N_5528);
or U6437 (N_6437,N_5157,N_5123);
xnor U6438 (N_6438,N_5813,N_5769);
and U6439 (N_6439,N_5454,N_5982);
xnor U6440 (N_6440,N_5573,N_5705);
or U6441 (N_6441,N_5700,N_5932);
nand U6442 (N_6442,N_5118,N_5752);
nor U6443 (N_6443,N_5268,N_5106);
or U6444 (N_6444,N_5642,N_5290);
xor U6445 (N_6445,N_5785,N_5959);
nand U6446 (N_6446,N_5808,N_5398);
nand U6447 (N_6447,N_5293,N_5987);
nand U6448 (N_6448,N_5717,N_5285);
or U6449 (N_6449,N_5737,N_5154);
nand U6450 (N_6450,N_5985,N_5602);
or U6451 (N_6451,N_5344,N_5230);
nor U6452 (N_6452,N_5865,N_5968);
and U6453 (N_6453,N_5352,N_5254);
or U6454 (N_6454,N_5337,N_5328);
nor U6455 (N_6455,N_5562,N_5758);
or U6456 (N_6456,N_5640,N_5412);
nand U6457 (N_6457,N_5547,N_5465);
or U6458 (N_6458,N_5366,N_5406);
nor U6459 (N_6459,N_5300,N_5371);
nand U6460 (N_6460,N_5840,N_5055);
nand U6461 (N_6461,N_5456,N_5698);
nor U6462 (N_6462,N_5360,N_5734);
nand U6463 (N_6463,N_5489,N_5621);
xnor U6464 (N_6464,N_5134,N_5132);
and U6465 (N_6465,N_5351,N_5182);
nand U6466 (N_6466,N_5804,N_5464);
and U6467 (N_6467,N_5020,N_5261);
and U6468 (N_6468,N_5002,N_5702);
nand U6469 (N_6469,N_5097,N_5723);
nor U6470 (N_6470,N_5689,N_5221);
and U6471 (N_6471,N_5277,N_5673);
or U6472 (N_6472,N_5747,N_5823);
nand U6473 (N_6473,N_5555,N_5387);
xor U6474 (N_6474,N_5346,N_5867);
and U6475 (N_6475,N_5349,N_5108);
nor U6476 (N_6476,N_5452,N_5469);
and U6477 (N_6477,N_5397,N_5113);
nand U6478 (N_6478,N_5613,N_5538);
and U6479 (N_6479,N_5090,N_5911);
and U6480 (N_6480,N_5017,N_5212);
or U6481 (N_6481,N_5158,N_5319);
nand U6482 (N_6482,N_5077,N_5706);
or U6483 (N_6483,N_5370,N_5479);
nor U6484 (N_6484,N_5316,N_5546);
and U6485 (N_6485,N_5970,N_5580);
nand U6486 (N_6486,N_5672,N_5992);
or U6487 (N_6487,N_5150,N_5520);
nor U6488 (N_6488,N_5041,N_5697);
xnor U6489 (N_6489,N_5044,N_5764);
nand U6490 (N_6490,N_5768,N_5249);
xor U6491 (N_6491,N_5145,N_5377);
nand U6492 (N_6492,N_5411,N_5750);
nand U6493 (N_6493,N_5870,N_5678);
xnor U6494 (N_6494,N_5850,N_5310);
nor U6495 (N_6495,N_5010,N_5023);
or U6496 (N_6496,N_5964,N_5856);
and U6497 (N_6497,N_5937,N_5936);
xor U6498 (N_6498,N_5331,N_5205);
or U6499 (N_6499,N_5295,N_5152);
nor U6500 (N_6500,N_5794,N_5704);
and U6501 (N_6501,N_5502,N_5683);
nand U6502 (N_6502,N_5274,N_5172);
or U6503 (N_6503,N_5629,N_5115);
xor U6504 (N_6504,N_5122,N_5023);
and U6505 (N_6505,N_5554,N_5930);
xnor U6506 (N_6506,N_5241,N_5105);
nor U6507 (N_6507,N_5580,N_5459);
nor U6508 (N_6508,N_5609,N_5597);
nand U6509 (N_6509,N_5401,N_5419);
nand U6510 (N_6510,N_5485,N_5252);
or U6511 (N_6511,N_5627,N_5118);
nor U6512 (N_6512,N_5404,N_5588);
and U6513 (N_6513,N_5801,N_5802);
and U6514 (N_6514,N_5226,N_5402);
xnor U6515 (N_6515,N_5126,N_5971);
or U6516 (N_6516,N_5695,N_5770);
and U6517 (N_6517,N_5967,N_5090);
nand U6518 (N_6518,N_5218,N_5272);
and U6519 (N_6519,N_5359,N_5021);
or U6520 (N_6520,N_5865,N_5126);
nand U6521 (N_6521,N_5833,N_5607);
nand U6522 (N_6522,N_5291,N_5064);
nand U6523 (N_6523,N_5184,N_5899);
nand U6524 (N_6524,N_5636,N_5848);
nor U6525 (N_6525,N_5006,N_5657);
nor U6526 (N_6526,N_5196,N_5903);
nand U6527 (N_6527,N_5093,N_5580);
nand U6528 (N_6528,N_5550,N_5861);
nor U6529 (N_6529,N_5750,N_5275);
or U6530 (N_6530,N_5627,N_5826);
or U6531 (N_6531,N_5004,N_5309);
or U6532 (N_6532,N_5933,N_5820);
and U6533 (N_6533,N_5568,N_5550);
and U6534 (N_6534,N_5716,N_5185);
or U6535 (N_6535,N_5057,N_5302);
nor U6536 (N_6536,N_5989,N_5561);
and U6537 (N_6537,N_5091,N_5056);
nor U6538 (N_6538,N_5858,N_5841);
nor U6539 (N_6539,N_5651,N_5010);
and U6540 (N_6540,N_5839,N_5330);
or U6541 (N_6541,N_5583,N_5811);
and U6542 (N_6542,N_5020,N_5427);
xor U6543 (N_6543,N_5704,N_5763);
nor U6544 (N_6544,N_5269,N_5085);
nor U6545 (N_6545,N_5023,N_5934);
and U6546 (N_6546,N_5951,N_5920);
xor U6547 (N_6547,N_5210,N_5259);
or U6548 (N_6548,N_5330,N_5731);
and U6549 (N_6549,N_5978,N_5356);
nor U6550 (N_6550,N_5735,N_5678);
xor U6551 (N_6551,N_5680,N_5306);
and U6552 (N_6552,N_5436,N_5216);
and U6553 (N_6553,N_5735,N_5958);
nand U6554 (N_6554,N_5100,N_5633);
or U6555 (N_6555,N_5411,N_5310);
or U6556 (N_6556,N_5264,N_5670);
nand U6557 (N_6557,N_5323,N_5069);
xnor U6558 (N_6558,N_5328,N_5088);
nand U6559 (N_6559,N_5529,N_5691);
or U6560 (N_6560,N_5562,N_5604);
or U6561 (N_6561,N_5997,N_5741);
nor U6562 (N_6562,N_5374,N_5888);
or U6563 (N_6563,N_5260,N_5356);
or U6564 (N_6564,N_5178,N_5878);
nand U6565 (N_6565,N_5835,N_5093);
and U6566 (N_6566,N_5474,N_5192);
nand U6567 (N_6567,N_5400,N_5321);
xnor U6568 (N_6568,N_5354,N_5660);
nor U6569 (N_6569,N_5947,N_5978);
xor U6570 (N_6570,N_5109,N_5237);
nand U6571 (N_6571,N_5221,N_5252);
nor U6572 (N_6572,N_5630,N_5036);
or U6573 (N_6573,N_5753,N_5660);
nor U6574 (N_6574,N_5673,N_5636);
xor U6575 (N_6575,N_5472,N_5266);
nor U6576 (N_6576,N_5350,N_5531);
nand U6577 (N_6577,N_5224,N_5557);
nand U6578 (N_6578,N_5523,N_5977);
nor U6579 (N_6579,N_5699,N_5998);
nor U6580 (N_6580,N_5900,N_5776);
and U6581 (N_6581,N_5802,N_5844);
xor U6582 (N_6582,N_5283,N_5814);
and U6583 (N_6583,N_5901,N_5441);
nand U6584 (N_6584,N_5003,N_5696);
nor U6585 (N_6585,N_5003,N_5888);
xor U6586 (N_6586,N_5224,N_5705);
nand U6587 (N_6587,N_5786,N_5371);
nor U6588 (N_6588,N_5686,N_5772);
nor U6589 (N_6589,N_5679,N_5004);
nor U6590 (N_6590,N_5834,N_5478);
nand U6591 (N_6591,N_5434,N_5435);
nor U6592 (N_6592,N_5390,N_5056);
nor U6593 (N_6593,N_5284,N_5709);
and U6594 (N_6594,N_5217,N_5872);
and U6595 (N_6595,N_5215,N_5842);
and U6596 (N_6596,N_5602,N_5924);
or U6597 (N_6597,N_5033,N_5149);
nor U6598 (N_6598,N_5785,N_5868);
nand U6599 (N_6599,N_5321,N_5972);
nand U6600 (N_6600,N_5487,N_5259);
or U6601 (N_6601,N_5447,N_5206);
nor U6602 (N_6602,N_5608,N_5229);
or U6603 (N_6603,N_5266,N_5105);
or U6604 (N_6604,N_5915,N_5392);
or U6605 (N_6605,N_5978,N_5509);
nand U6606 (N_6606,N_5330,N_5353);
and U6607 (N_6607,N_5770,N_5371);
and U6608 (N_6608,N_5198,N_5049);
nand U6609 (N_6609,N_5044,N_5299);
nor U6610 (N_6610,N_5447,N_5041);
nand U6611 (N_6611,N_5283,N_5445);
nand U6612 (N_6612,N_5299,N_5195);
xor U6613 (N_6613,N_5297,N_5390);
nor U6614 (N_6614,N_5287,N_5020);
xor U6615 (N_6615,N_5626,N_5689);
and U6616 (N_6616,N_5404,N_5950);
xor U6617 (N_6617,N_5077,N_5207);
nor U6618 (N_6618,N_5495,N_5241);
nand U6619 (N_6619,N_5842,N_5796);
nor U6620 (N_6620,N_5610,N_5357);
xnor U6621 (N_6621,N_5696,N_5410);
nand U6622 (N_6622,N_5552,N_5391);
nor U6623 (N_6623,N_5775,N_5755);
and U6624 (N_6624,N_5516,N_5792);
nor U6625 (N_6625,N_5548,N_5384);
nand U6626 (N_6626,N_5684,N_5523);
xnor U6627 (N_6627,N_5148,N_5784);
nand U6628 (N_6628,N_5357,N_5945);
nand U6629 (N_6629,N_5513,N_5552);
nand U6630 (N_6630,N_5715,N_5722);
nor U6631 (N_6631,N_5242,N_5162);
and U6632 (N_6632,N_5932,N_5325);
and U6633 (N_6633,N_5064,N_5780);
nand U6634 (N_6634,N_5226,N_5822);
or U6635 (N_6635,N_5999,N_5418);
xnor U6636 (N_6636,N_5834,N_5477);
nand U6637 (N_6637,N_5755,N_5125);
or U6638 (N_6638,N_5386,N_5375);
nor U6639 (N_6639,N_5383,N_5089);
nand U6640 (N_6640,N_5430,N_5502);
and U6641 (N_6641,N_5048,N_5733);
nor U6642 (N_6642,N_5361,N_5885);
or U6643 (N_6643,N_5130,N_5586);
or U6644 (N_6644,N_5878,N_5858);
xor U6645 (N_6645,N_5236,N_5925);
xor U6646 (N_6646,N_5383,N_5498);
nand U6647 (N_6647,N_5168,N_5600);
nand U6648 (N_6648,N_5231,N_5680);
or U6649 (N_6649,N_5350,N_5066);
and U6650 (N_6650,N_5565,N_5112);
and U6651 (N_6651,N_5399,N_5333);
nand U6652 (N_6652,N_5046,N_5825);
or U6653 (N_6653,N_5949,N_5067);
and U6654 (N_6654,N_5464,N_5541);
nand U6655 (N_6655,N_5079,N_5728);
nand U6656 (N_6656,N_5871,N_5959);
nand U6657 (N_6657,N_5801,N_5397);
and U6658 (N_6658,N_5504,N_5797);
xor U6659 (N_6659,N_5988,N_5045);
xnor U6660 (N_6660,N_5281,N_5113);
and U6661 (N_6661,N_5445,N_5864);
nor U6662 (N_6662,N_5281,N_5115);
xnor U6663 (N_6663,N_5355,N_5468);
nand U6664 (N_6664,N_5059,N_5533);
or U6665 (N_6665,N_5334,N_5976);
nor U6666 (N_6666,N_5468,N_5138);
and U6667 (N_6667,N_5651,N_5994);
nor U6668 (N_6668,N_5175,N_5265);
and U6669 (N_6669,N_5735,N_5998);
or U6670 (N_6670,N_5631,N_5804);
and U6671 (N_6671,N_5630,N_5366);
and U6672 (N_6672,N_5219,N_5875);
or U6673 (N_6673,N_5874,N_5343);
and U6674 (N_6674,N_5069,N_5101);
nand U6675 (N_6675,N_5925,N_5203);
nand U6676 (N_6676,N_5641,N_5658);
xnor U6677 (N_6677,N_5659,N_5918);
xnor U6678 (N_6678,N_5680,N_5111);
and U6679 (N_6679,N_5201,N_5907);
or U6680 (N_6680,N_5672,N_5427);
and U6681 (N_6681,N_5314,N_5306);
and U6682 (N_6682,N_5894,N_5922);
nor U6683 (N_6683,N_5578,N_5805);
or U6684 (N_6684,N_5794,N_5837);
and U6685 (N_6685,N_5861,N_5122);
nand U6686 (N_6686,N_5234,N_5475);
and U6687 (N_6687,N_5419,N_5711);
or U6688 (N_6688,N_5679,N_5258);
nor U6689 (N_6689,N_5035,N_5076);
and U6690 (N_6690,N_5012,N_5329);
or U6691 (N_6691,N_5308,N_5241);
nor U6692 (N_6692,N_5324,N_5007);
nor U6693 (N_6693,N_5604,N_5870);
xnor U6694 (N_6694,N_5408,N_5962);
or U6695 (N_6695,N_5559,N_5263);
nand U6696 (N_6696,N_5593,N_5207);
or U6697 (N_6697,N_5736,N_5234);
xor U6698 (N_6698,N_5117,N_5487);
and U6699 (N_6699,N_5043,N_5419);
and U6700 (N_6700,N_5520,N_5780);
and U6701 (N_6701,N_5440,N_5693);
nor U6702 (N_6702,N_5572,N_5687);
and U6703 (N_6703,N_5705,N_5271);
nor U6704 (N_6704,N_5581,N_5789);
or U6705 (N_6705,N_5517,N_5977);
and U6706 (N_6706,N_5512,N_5095);
nand U6707 (N_6707,N_5004,N_5757);
and U6708 (N_6708,N_5871,N_5924);
nand U6709 (N_6709,N_5845,N_5231);
and U6710 (N_6710,N_5291,N_5907);
nand U6711 (N_6711,N_5042,N_5163);
nand U6712 (N_6712,N_5052,N_5239);
and U6713 (N_6713,N_5729,N_5345);
nand U6714 (N_6714,N_5179,N_5199);
nand U6715 (N_6715,N_5853,N_5718);
or U6716 (N_6716,N_5626,N_5552);
and U6717 (N_6717,N_5151,N_5591);
or U6718 (N_6718,N_5716,N_5922);
and U6719 (N_6719,N_5528,N_5612);
and U6720 (N_6720,N_5023,N_5041);
nor U6721 (N_6721,N_5777,N_5599);
and U6722 (N_6722,N_5182,N_5998);
or U6723 (N_6723,N_5164,N_5482);
and U6724 (N_6724,N_5492,N_5659);
and U6725 (N_6725,N_5144,N_5483);
nor U6726 (N_6726,N_5166,N_5509);
xor U6727 (N_6727,N_5524,N_5242);
and U6728 (N_6728,N_5718,N_5904);
nor U6729 (N_6729,N_5437,N_5564);
and U6730 (N_6730,N_5463,N_5789);
or U6731 (N_6731,N_5060,N_5776);
xor U6732 (N_6732,N_5337,N_5068);
xor U6733 (N_6733,N_5405,N_5598);
nand U6734 (N_6734,N_5255,N_5895);
nor U6735 (N_6735,N_5307,N_5405);
nor U6736 (N_6736,N_5622,N_5561);
and U6737 (N_6737,N_5589,N_5708);
xnor U6738 (N_6738,N_5205,N_5564);
or U6739 (N_6739,N_5063,N_5288);
or U6740 (N_6740,N_5553,N_5005);
nor U6741 (N_6741,N_5400,N_5999);
nor U6742 (N_6742,N_5615,N_5233);
nand U6743 (N_6743,N_5950,N_5914);
and U6744 (N_6744,N_5750,N_5089);
nor U6745 (N_6745,N_5935,N_5107);
or U6746 (N_6746,N_5927,N_5991);
and U6747 (N_6747,N_5164,N_5682);
or U6748 (N_6748,N_5892,N_5275);
or U6749 (N_6749,N_5951,N_5495);
and U6750 (N_6750,N_5825,N_5030);
and U6751 (N_6751,N_5086,N_5882);
nor U6752 (N_6752,N_5431,N_5384);
nand U6753 (N_6753,N_5948,N_5196);
nand U6754 (N_6754,N_5472,N_5153);
nand U6755 (N_6755,N_5844,N_5361);
nor U6756 (N_6756,N_5273,N_5833);
or U6757 (N_6757,N_5324,N_5858);
xor U6758 (N_6758,N_5985,N_5756);
nand U6759 (N_6759,N_5839,N_5410);
or U6760 (N_6760,N_5358,N_5610);
nor U6761 (N_6761,N_5160,N_5873);
nand U6762 (N_6762,N_5810,N_5278);
nor U6763 (N_6763,N_5957,N_5670);
nand U6764 (N_6764,N_5708,N_5043);
nand U6765 (N_6765,N_5789,N_5029);
or U6766 (N_6766,N_5981,N_5675);
nor U6767 (N_6767,N_5067,N_5279);
or U6768 (N_6768,N_5021,N_5243);
or U6769 (N_6769,N_5683,N_5979);
nor U6770 (N_6770,N_5212,N_5046);
or U6771 (N_6771,N_5162,N_5416);
nor U6772 (N_6772,N_5439,N_5914);
nor U6773 (N_6773,N_5219,N_5384);
or U6774 (N_6774,N_5326,N_5896);
or U6775 (N_6775,N_5423,N_5171);
xor U6776 (N_6776,N_5807,N_5142);
nor U6777 (N_6777,N_5946,N_5250);
and U6778 (N_6778,N_5637,N_5947);
or U6779 (N_6779,N_5583,N_5169);
nor U6780 (N_6780,N_5050,N_5983);
xnor U6781 (N_6781,N_5201,N_5255);
or U6782 (N_6782,N_5470,N_5286);
nand U6783 (N_6783,N_5250,N_5004);
nand U6784 (N_6784,N_5382,N_5971);
or U6785 (N_6785,N_5900,N_5062);
and U6786 (N_6786,N_5474,N_5382);
xor U6787 (N_6787,N_5071,N_5427);
nor U6788 (N_6788,N_5597,N_5134);
nor U6789 (N_6789,N_5897,N_5429);
nand U6790 (N_6790,N_5792,N_5892);
or U6791 (N_6791,N_5630,N_5142);
nand U6792 (N_6792,N_5065,N_5646);
and U6793 (N_6793,N_5544,N_5329);
or U6794 (N_6794,N_5299,N_5545);
nand U6795 (N_6795,N_5330,N_5905);
nand U6796 (N_6796,N_5235,N_5909);
or U6797 (N_6797,N_5755,N_5578);
and U6798 (N_6798,N_5304,N_5651);
nand U6799 (N_6799,N_5245,N_5038);
or U6800 (N_6800,N_5561,N_5540);
nor U6801 (N_6801,N_5302,N_5158);
nor U6802 (N_6802,N_5532,N_5801);
and U6803 (N_6803,N_5938,N_5332);
or U6804 (N_6804,N_5088,N_5406);
or U6805 (N_6805,N_5074,N_5137);
and U6806 (N_6806,N_5994,N_5383);
nand U6807 (N_6807,N_5937,N_5835);
nor U6808 (N_6808,N_5650,N_5974);
and U6809 (N_6809,N_5867,N_5537);
nor U6810 (N_6810,N_5142,N_5867);
or U6811 (N_6811,N_5020,N_5751);
nand U6812 (N_6812,N_5699,N_5176);
and U6813 (N_6813,N_5911,N_5400);
nand U6814 (N_6814,N_5205,N_5726);
nor U6815 (N_6815,N_5200,N_5948);
and U6816 (N_6816,N_5457,N_5718);
xnor U6817 (N_6817,N_5327,N_5750);
nor U6818 (N_6818,N_5683,N_5876);
or U6819 (N_6819,N_5395,N_5101);
and U6820 (N_6820,N_5384,N_5938);
nor U6821 (N_6821,N_5208,N_5850);
and U6822 (N_6822,N_5878,N_5340);
nand U6823 (N_6823,N_5373,N_5489);
nand U6824 (N_6824,N_5514,N_5202);
nand U6825 (N_6825,N_5941,N_5614);
nand U6826 (N_6826,N_5743,N_5279);
and U6827 (N_6827,N_5302,N_5887);
or U6828 (N_6828,N_5866,N_5050);
and U6829 (N_6829,N_5967,N_5651);
and U6830 (N_6830,N_5601,N_5911);
and U6831 (N_6831,N_5839,N_5783);
nor U6832 (N_6832,N_5388,N_5506);
nor U6833 (N_6833,N_5403,N_5082);
or U6834 (N_6834,N_5558,N_5493);
or U6835 (N_6835,N_5780,N_5336);
and U6836 (N_6836,N_5347,N_5613);
nand U6837 (N_6837,N_5385,N_5001);
and U6838 (N_6838,N_5560,N_5002);
nand U6839 (N_6839,N_5819,N_5596);
nand U6840 (N_6840,N_5310,N_5988);
nor U6841 (N_6841,N_5679,N_5051);
nor U6842 (N_6842,N_5345,N_5517);
nand U6843 (N_6843,N_5301,N_5554);
and U6844 (N_6844,N_5274,N_5967);
nor U6845 (N_6845,N_5322,N_5381);
and U6846 (N_6846,N_5418,N_5519);
nor U6847 (N_6847,N_5053,N_5653);
or U6848 (N_6848,N_5258,N_5755);
nor U6849 (N_6849,N_5093,N_5757);
or U6850 (N_6850,N_5205,N_5809);
and U6851 (N_6851,N_5551,N_5753);
xor U6852 (N_6852,N_5941,N_5354);
or U6853 (N_6853,N_5717,N_5956);
nor U6854 (N_6854,N_5712,N_5485);
xor U6855 (N_6855,N_5328,N_5308);
nor U6856 (N_6856,N_5107,N_5374);
and U6857 (N_6857,N_5540,N_5767);
and U6858 (N_6858,N_5974,N_5122);
xor U6859 (N_6859,N_5494,N_5610);
or U6860 (N_6860,N_5852,N_5348);
or U6861 (N_6861,N_5935,N_5695);
or U6862 (N_6862,N_5031,N_5502);
and U6863 (N_6863,N_5918,N_5776);
and U6864 (N_6864,N_5456,N_5865);
nand U6865 (N_6865,N_5058,N_5274);
or U6866 (N_6866,N_5307,N_5861);
and U6867 (N_6867,N_5661,N_5673);
xor U6868 (N_6868,N_5594,N_5115);
or U6869 (N_6869,N_5081,N_5122);
or U6870 (N_6870,N_5719,N_5604);
and U6871 (N_6871,N_5862,N_5033);
nand U6872 (N_6872,N_5868,N_5370);
or U6873 (N_6873,N_5196,N_5176);
xor U6874 (N_6874,N_5811,N_5551);
nand U6875 (N_6875,N_5377,N_5675);
nand U6876 (N_6876,N_5752,N_5083);
or U6877 (N_6877,N_5624,N_5239);
nand U6878 (N_6878,N_5969,N_5338);
nand U6879 (N_6879,N_5392,N_5005);
nand U6880 (N_6880,N_5391,N_5985);
nand U6881 (N_6881,N_5997,N_5211);
and U6882 (N_6882,N_5765,N_5310);
nor U6883 (N_6883,N_5753,N_5654);
nand U6884 (N_6884,N_5061,N_5511);
nor U6885 (N_6885,N_5466,N_5987);
nand U6886 (N_6886,N_5189,N_5903);
or U6887 (N_6887,N_5989,N_5837);
nand U6888 (N_6888,N_5518,N_5430);
and U6889 (N_6889,N_5676,N_5764);
nand U6890 (N_6890,N_5337,N_5493);
nor U6891 (N_6891,N_5997,N_5620);
nor U6892 (N_6892,N_5327,N_5329);
or U6893 (N_6893,N_5752,N_5576);
or U6894 (N_6894,N_5460,N_5743);
or U6895 (N_6895,N_5912,N_5157);
nand U6896 (N_6896,N_5429,N_5798);
and U6897 (N_6897,N_5703,N_5210);
and U6898 (N_6898,N_5979,N_5408);
or U6899 (N_6899,N_5751,N_5093);
nor U6900 (N_6900,N_5170,N_5283);
and U6901 (N_6901,N_5654,N_5961);
and U6902 (N_6902,N_5383,N_5373);
nor U6903 (N_6903,N_5239,N_5097);
or U6904 (N_6904,N_5900,N_5516);
nand U6905 (N_6905,N_5060,N_5981);
nand U6906 (N_6906,N_5817,N_5670);
and U6907 (N_6907,N_5192,N_5715);
nor U6908 (N_6908,N_5333,N_5884);
xnor U6909 (N_6909,N_5301,N_5113);
nor U6910 (N_6910,N_5588,N_5205);
xnor U6911 (N_6911,N_5610,N_5393);
nand U6912 (N_6912,N_5198,N_5679);
nand U6913 (N_6913,N_5207,N_5738);
xor U6914 (N_6914,N_5593,N_5908);
and U6915 (N_6915,N_5064,N_5924);
and U6916 (N_6916,N_5840,N_5733);
or U6917 (N_6917,N_5285,N_5632);
or U6918 (N_6918,N_5309,N_5368);
nand U6919 (N_6919,N_5082,N_5590);
and U6920 (N_6920,N_5316,N_5989);
xnor U6921 (N_6921,N_5003,N_5143);
nor U6922 (N_6922,N_5967,N_5965);
nor U6923 (N_6923,N_5130,N_5002);
and U6924 (N_6924,N_5381,N_5574);
or U6925 (N_6925,N_5711,N_5080);
nor U6926 (N_6926,N_5504,N_5320);
nand U6927 (N_6927,N_5835,N_5354);
nor U6928 (N_6928,N_5748,N_5526);
nor U6929 (N_6929,N_5430,N_5976);
nand U6930 (N_6930,N_5227,N_5017);
and U6931 (N_6931,N_5119,N_5913);
nor U6932 (N_6932,N_5436,N_5867);
nor U6933 (N_6933,N_5456,N_5522);
xor U6934 (N_6934,N_5960,N_5445);
and U6935 (N_6935,N_5872,N_5126);
nand U6936 (N_6936,N_5678,N_5099);
and U6937 (N_6937,N_5654,N_5418);
nor U6938 (N_6938,N_5094,N_5443);
or U6939 (N_6939,N_5021,N_5014);
and U6940 (N_6940,N_5821,N_5122);
nor U6941 (N_6941,N_5467,N_5940);
nand U6942 (N_6942,N_5710,N_5847);
or U6943 (N_6943,N_5195,N_5568);
nand U6944 (N_6944,N_5031,N_5705);
or U6945 (N_6945,N_5654,N_5406);
xor U6946 (N_6946,N_5350,N_5283);
xor U6947 (N_6947,N_5035,N_5148);
and U6948 (N_6948,N_5502,N_5017);
nor U6949 (N_6949,N_5977,N_5783);
and U6950 (N_6950,N_5894,N_5398);
or U6951 (N_6951,N_5606,N_5503);
nand U6952 (N_6952,N_5639,N_5095);
xnor U6953 (N_6953,N_5455,N_5865);
and U6954 (N_6954,N_5267,N_5399);
or U6955 (N_6955,N_5827,N_5883);
xor U6956 (N_6956,N_5455,N_5322);
or U6957 (N_6957,N_5400,N_5196);
nor U6958 (N_6958,N_5891,N_5791);
and U6959 (N_6959,N_5446,N_5783);
or U6960 (N_6960,N_5479,N_5905);
xor U6961 (N_6961,N_5744,N_5957);
nand U6962 (N_6962,N_5285,N_5535);
xnor U6963 (N_6963,N_5114,N_5980);
xor U6964 (N_6964,N_5991,N_5054);
xor U6965 (N_6965,N_5090,N_5872);
nor U6966 (N_6966,N_5970,N_5227);
nand U6967 (N_6967,N_5309,N_5310);
nand U6968 (N_6968,N_5911,N_5214);
or U6969 (N_6969,N_5656,N_5161);
and U6970 (N_6970,N_5960,N_5708);
and U6971 (N_6971,N_5060,N_5037);
nand U6972 (N_6972,N_5190,N_5390);
nor U6973 (N_6973,N_5375,N_5853);
or U6974 (N_6974,N_5673,N_5981);
and U6975 (N_6975,N_5680,N_5576);
nor U6976 (N_6976,N_5885,N_5111);
nand U6977 (N_6977,N_5838,N_5441);
and U6978 (N_6978,N_5101,N_5208);
and U6979 (N_6979,N_5015,N_5090);
nand U6980 (N_6980,N_5105,N_5310);
or U6981 (N_6981,N_5796,N_5186);
and U6982 (N_6982,N_5255,N_5952);
nor U6983 (N_6983,N_5737,N_5918);
and U6984 (N_6984,N_5622,N_5486);
nor U6985 (N_6985,N_5908,N_5918);
nand U6986 (N_6986,N_5560,N_5745);
nand U6987 (N_6987,N_5032,N_5996);
nor U6988 (N_6988,N_5875,N_5674);
and U6989 (N_6989,N_5293,N_5456);
and U6990 (N_6990,N_5308,N_5279);
nand U6991 (N_6991,N_5450,N_5256);
and U6992 (N_6992,N_5781,N_5255);
nor U6993 (N_6993,N_5174,N_5220);
and U6994 (N_6994,N_5971,N_5918);
nor U6995 (N_6995,N_5742,N_5193);
or U6996 (N_6996,N_5537,N_5466);
and U6997 (N_6997,N_5462,N_5015);
nand U6998 (N_6998,N_5317,N_5077);
nand U6999 (N_6999,N_5266,N_5617);
and U7000 (N_7000,N_6516,N_6842);
and U7001 (N_7001,N_6670,N_6690);
xnor U7002 (N_7002,N_6780,N_6575);
xor U7003 (N_7003,N_6436,N_6165);
nor U7004 (N_7004,N_6904,N_6605);
nand U7005 (N_7005,N_6832,N_6583);
nor U7006 (N_7006,N_6430,N_6635);
or U7007 (N_7007,N_6547,N_6084);
and U7008 (N_7008,N_6132,N_6926);
and U7009 (N_7009,N_6879,N_6413);
and U7010 (N_7010,N_6660,N_6317);
and U7011 (N_7011,N_6481,N_6802);
and U7012 (N_7012,N_6141,N_6040);
nand U7013 (N_7013,N_6594,N_6743);
or U7014 (N_7014,N_6445,N_6927);
and U7015 (N_7015,N_6965,N_6088);
nand U7016 (N_7016,N_6607,N_6221);
nand U7017 (N_7017,N_6759,N_6433);
nand U7018 (N_7018,N_6910,N_6324);
or U7019 (N_7019,N_6036,N_6370);
or U7020 (N_7020,N_6891,N_6995);
nor U7021 (N_7021,N_6854,N_6111);
nor U7022 (N_7022,N_6341,N_6820);
nand U7023 (N_7023,N_6708,N_6488);
and U7024 (N_7024,N_6231,N_6022);
nand U7025 (N_7025,N_6963,N_6089);
and U7026 (N_7026,N_6086,N_6396);
nor U7027 (N_7027,N_6405,N_6801);
nand U7028 (N_7028,N_6588,N_6002);
nand U7029 (N_7029,N_6360,N_6951);
nand U7030 (N_7030,N_6090,N_6980);
and U7031 (N_7031,N_6447,N_6182);
xor U7032 (N_7032,N_6807,N_6905);
nor U7033 (N_7033,N_6848,N_6915);
nor U7034 (N_7034,N_6145,N_6792);
or U7035 (N_7035,N_6144,N_6730);
nand U7036 (N_7036,N_6301,N_6782);
nor U7037 (N_7037,N_6418,N_6282);
or U7038 (N_7038,N_6200,N_6471);
and U7039 (N_7039,N_6307,N_6810);
nor U7040 (N_7040,N_6299,N_6985);
and U7041 (N_7041,N_6202,N_6806);
nor U7042 (N_7042,N_6121,N_6937);
or U7043 (N_7043,N_6417,N_6161);
or U7044 (N_7044,N_6258,N_6816);
and U7045 (N_7045,N_6160,N_6343);
nor U7046 (N_7046,N_6817,N_6725);
and U7047 (N_7047,N_6813,N_6442);
nor U7048 (N_7048,N_6552,N_6726);
nor U7049 (N_7049,N_6909,N_6600);
nor U7050 (N_7050,N_6455,N_6305);
or U7051 (N_7051,N_6509,N_6123);
nand U7052 (N_7052,N_6033,N_6765);
or U7053 (N_7053,N_6784,N_6596);
and U7054 (N_7054,N_6535,N_6595);
or U7055 (N_7055,N_6793,N_6928);
nor U7056 (N_7056,N_6239,N_6653);
nand U7057 (N_7057,N_6811,N_6948);
or U7058 (N_7058,N_6008,N_6054);
nand U7059 (N_7059,N_6727,N_6391);
xor U7060 (N_7060,N_6917,N_6210);
nor U7061 (N_7061,N_6235,N_6987);
or U7062 (N_7062,N_6450,N_6183);
xnor U7063 (N_7063,N_6122,N_6911);
nor U7064 (N_7064,N_6335,N_6888);
or U7065 (N_7065,N_6023,N_6614);
or U7066 (N_7066,N_6511,N_6678);
or U7067 (N_7067,N_6869,N_6972);
nand U7068 (N_7068,N_6382,N_6626);
and U7069 (N_7069,N_6250,N_6613);
nand U7070 (N_7070,N_6698,N_6975);
nand U7071 (N_7071,N_6289,N_6380);
and U7072 (N_7072,N_6104,N_6032);
xnor U7073 (N_7073,N_6428,N_6761);
and U7074 (N_7074,N_6047,N_6066);
and U7075 (N_7075,N_6143,N_6974);
nand U7076 (N_7076,N_6188,N_6700);
and U7077 (N_7077,N_6618,N_6701);
and U7078 (N_7078,N_6003,N_6757);
and U7079 (N_7079,N_6611,N_6196);
nor U7080 (N_7080,N_6648,N_6679);
or U7081 (N_7081,N_6247,N_6006);
nand U7082 (N_7082,N_6402,N_6979);
nand U7083 (N_7083,N_6933,N_6174);
or U7084 (N_7084,N_6944,N_6156);
and U7085 (N_7085,N_6489,N_6860);
nor U7086 (N_7086,N_6691,N_6201);
nor U7087 (N_7087,N_6107,N_6186);
nor U7088 (N_7088,N_6293,N_6105);
and U7089 (N_7089,N_6898,N_6712);
and U7090 (N_7090,N_6046,N_6146);
or U7091 (N_7091,N_6866,N_6395);
nor U7092 (N_7092,N_6497,N_6986);
or U7093 (N_7093,N_6821,N_6052);
nand U7094 (N_7094,N_6722,N_6303);
and U7095 (N_7095,N_6955,N_6207);
nor U7096 (N_7096,N_6456,N_6276);
and U7097 (N_7097,N_6192,N_6110);
nor U7098 (N_7098,N_6525,N_6919);
or U7099 (N_7099,N_6199,N_6078);
xnor U7100 (N_7100,N_6732,N_6997);
and U7101 (N_7101,N_6030,N_6357);
or U7102 (N_7102,N_6119,N_6855);
or U7103 (N_7103,N_6018,N_6181);
nand U7104 (N_7104,N_6067,N_6234);
nand U7105 (N_7105,N_6443,N_6283);
and U7106 (N_7106,N_6735,N_6237);
and U7107 (N_7107,N_6561,N_6296);
and U7108 (N_7108,N_6387,N_6220);
nand U7109 (N_7109,N_6706,N_6072);
and U7110 (N_7110,N_6696,N_6559);
nor U7111 (N_7111,N_6758,N_6458);
or U7112 (N_7112,N_6826,N_6334);
or U7113 (N_7113,N_6913,N_6823);
or U7114 (N_7114,N_6211,N_6197);
xnor U7115 (N_7115,N_6562,N_6278);
xnor U7116 (N_7116,N_6604,N_6886);
xnor U7117 (N_7117,N_6486,N_6058);
and U7118 (N_7118,N_6134,N_6342);
and U7119 (N_7119,N_6924,N_6592);
nand U7120 (N_7120,N_6885,N_6464);
and U7121 (N_7121,N_6203,N_6271);
and U7122 (N_7122,N_6059,N_6615);
and U7123 (N_7123,N_6749,N_6045);
or U7124 (N_7124,N_6652,N_6640);
nand U7125 (N_7125,N_6410,N_6272);
nand U7126 (N_7126,N_6333,N_6275);
xor U7127 (N_7127,N_6063,N_6876);
nor U7128 (N_7128,N_6808,N_6889);
nor U7129 (N_7129,N_6795,N_6356);
or U7130 (N_7130,N_6835,N_6731);
nand U7131 (N_7131,N_6347,N_6365);
nand U7132 (N_7132,N_6208,N_6563);
and U7133 (N_7133,N_6338,N_6718);
nand U7134 (N_7134,N_6238,N_6620);
or U7135 (N_7135,N_6408,N_6873);
and U7136 (N_7136,N_6949,N_6853);
and U7137 (N_7137,N_6568,N_6457);
and U7138 (N_7138,N_6786,N_6300);
and U7139 (N_7139,N_6064,N_6262);
nor U7140 (N_7140,N_6688,N_6740);
and U7141 (N_7141,N_6709,N_6479);
or U7142 (N_7142,N_6976,N_6403);
nor U7143 (N_7143,N_6325,N_6222);
nand U7144 (N_7144,N_6263,N_6249);
nor U7145 (N_7145,N_6930,N_6109);
and U7146 (N_7146,N_6358,N_6112);
nor U7147 (N_7147,N_6268,N_6477);
or U7148 (N_7148,N_6093,N_6623);
or U7149 (N_7149,N_6796,N_6870);
and U7150 (N_7150,N_6541,N_6850);
and U7151 (N_7151,N_6680,N_6179);
nand U7152 (N_7152,N_6374,N_6857);
nor U7153 (N_7153,N_6935,N_6881);
nor U7154 (N_7154,N_6131,N_6633);
nor U7155 (N_7155,N_6591,N_6554);
nand U7156 (N_7156,N_6906,N_6460);
nand U7157 (N_7157,N_6280,N_6564);
or U7158 (N_7158,N_6232,N_6589);
nand U7159 (N_7159,N_6503,N_6474);
nand U7160 (N_7160,N_6116,N_6149);
xnor U7161 (N_7161,N_6557,N_6543);
nor U7162 (N_7162,N_6827,N_6065);
xnor U7163 (N_7163,N_6133,N_6159);
xor U7164 (N_7164,N_6839,N_6274);
or U7165 (N_7165,N_6713,N_6597);
and U7166 (N_7166,N_6969,N_6137);
or U7167 (N_7167,N_6916,N_6081);
and U7168 (N_7168,N_6669,N_6892);
or U7169 (N_7169,N_6261,N_6799);
or U7170 (N_7170,N_6327,N_6627);
nand U7171 (N_7171,N_6742,N_6931);
nand U7172 (N_7172,N_6377,N_6998);
or U7173 (N_7173,N_6630,N_6332);
and U7174 (N_7174,N_6354,N_6057);
nor U7175 (N_7175,N_6290,N_6896);
xnor U7176 (N_7176,N_6363,N_6245);
nor U7177 (N_7177,N_6230,N_6136);
and U7178 (N_7178,N_6170,N_6331);
nor U7179 (N_7179,N_6496,N_6053);
nor U7180 (N_7180,N_6942,N_6958);
or U7181 (N_7181,N_6493,N_6007);
and U7182 (N_7182,N_6120,N_6102);
nor U7183 (N_7183,N_6298,N_6426);
nor U7184 (N_7184,N_6394,N_6756);
nor U7185 (N_7185,N_6752,N_6233);
and U7186 (N_7186,N_6687,N_6828);
and U7187 (N_7187,N_6314,N_6152);
xnor U7188 (N_7188,N_6026,N_6567);
or U7189 (N_7189,N_6814,N_6637);
and U7190 (N_7190,N_6462,N_6406);
and U7191 (N_7191,N_6362,N_6427);
nor U7192 (N_7192,N_6809,N_6175);
or U7193 (N_7193,N_6527,N_6586);
nand U7194 (N_7194,N_6952,N_6621);
nor U7195 (N_7195,N_6649,N_6114);
and U7196 (N_7196,N_6555,N_6536);
nor U7197 (N_7197,N_6281,N_6168);
or U7198 (N_7198,N_6968,N_6862);
and U7199 (N_7199,N_6506,N_6704);
nand U7200 (N_7200,N_6566,N_6981);
and U7201 (N_7201,N_6724,N_6710);
and U7202 (N_7202,N_6060,N_6528);
nand U7203 (N_7203,N_6872,N_6517);
or U7204 (N_7204,N_6666,N_6939);
and U7205 (N_7205,N_6647,N_6225);
nand U7206 (N_7206,N_6316,N_6452);
nand U7207 (N_7207,N_6480,N_6505);
and U7208 (N_7208,N_6599,N_6602);
and U7209 (N_7209,N_6893,N_6800);
or U7210 (N_7210,N_6767,N_6882);
nand U7211 (N_7211,N_6849,N_6075);
nor U7212 (N_7212,N_6010,N_6651);
or U7213 (N_7213,N_6512,N_6073);
and U7214 (N_7214,N_6254,N_6750);
nand U7215 (N_7215,N_6490,N_6076);
nor U7216 (N_7216,N_6993,N_6843);
and U7217 (N_7217,N_6431,N_6071);
or U7218 (N_7218,N_6932,N_6962);
nor U7219 (N_7219,N_6585,N_6351);
nand U7220 (N_7220,N_6227,N_6265);
nand U7221 (N_7221,N_6988,N_6302);
or U7222 (N_7222,N_6689,N_6773);
and U7223 (N_7223,N_6309,N_6884);
nor U7224 (N_7224,N_6451,N_6631);
or U7225 (N_7225,N_6819,N_6542);
and U7226 (N_7226,N_6856,N_6950);
nand U7227 (N_7227,N_6330,N_6390);
nor U7228 (N_7228,N_6518,N_6492);
or U7229 (N_7229,N_6124,N_6521);
xnor U7230 (N_7230,N_6661,N_6617);
nand U7231 (N_7231,N_6646,N_6619);
or U7232 (N_7232,N_6092,N_6941);
xor U7233 (N_7233,N_6625,N_6794);
nor U7234 (N_7234,N_6297,N_6683);
or U7235 (N_7235,N_6744,N_6344);
or U7236 (N_7236,N_6781,N_6502);
and U7237 (N_7237,N_6665,N_6957);
xor U7238 (N_7238,N_6864,N_6508);
or U7239 (N_7239,N_6887,N_6004);
or U7240 (N_7240,N_6533,N_6553);
nor U7241 (N_7241,N_6548,N_6522);
nor U7242 (N_7242,N_6257,N_6106);
nor U7243 (N_7243,N_6108,N_6540);
or U7244 (N_7244,N_6013,N_6644);
nand U7245 (N_7245,N_6544,N_6478);
xnor U7246 (N_7246,N_6472,N_6778);
xnor U7247 (N_7247,N_6096,N_6947);
and U7248 (N_7248,N_6014,N_6598);
or U7249 (N_7249,N_6659,N_6984);
or U7250 (N_7250,N_6118,N_6438);
and U7251 (N_7251,N_6769,N_6654);
or U7252 (N_7252,N_6310,N_6774);
nor U7253 (N_7253,N_6736,N_6844);
xor U7254 (N_7254,N_6049,N_6601);
or U7255 (N_7255,N_6982,N_6579);
and U7256 (N_7256,N_6323,N_6270);
nor U7257 (N_7257,N_6142,N_6345);
nand U7258 (N_7258,N_6404,N_6476);
or U7259 (N_7259,N_6584,N_6677);
nor U7260 (N_7260,N_6000,N_6153);
xor U7261 (N_7261,N_6126,N_6244);
and U7262 (N_7262,N_6069,N_6087);
or U7263 (N_7263,N_6461,N_6815);
nand U7264 (N_7264,N_6024,N_6176);
xor U7265 (N_7265,N_6914,N_6966);
and U7266 (N_7266,N_6632,N_6499);
or U7267 (N_7267,N_6603,N_6895);
and U7268 (N_7268,N_6441,N_6240);
nand U7269 (N_7269,N_6009,N_6779);
nand U7270 (N_7270,N_6125,N_6838);
or U7271 (N_7271,N_6286,N_6279);
nand U7272 (N_7272,N_6100,N_6352);
or U7273 (N_7273,N_6373,N_6184);
nand U7274 (N_7274,N_6874,N_6812);
xnor U7275 (N_7275,N_6287,N_6349);
nor U7276 (N_7276,N_6346,N_6039);
nand U7277 (N_7277,N_6538,N_6042);
or U7278 (N_7278,N_6167,N_6117);
or U7279 (N_7279,N_6714,N_6675);
and U7280 (N_7280,N_6751,N_6241);
or U7281 (N_7281,N_6269,N_6050);
nor U7282 (N_7282,N_6861,N_6587);
nor U7283 (N_7283,N_6925,N_6673);
nand U7284 (N_7284,N_6135,N_6399);
nor U7285 (N_7285,N_6074,N_6482);
and U7286 (N_7286,N_6558,N_6498);
or U7287 (N_7287,N_6285,N_6775);
or U7288 (N_7288,N_6733,N_6771);
nand U7289 (N_7289,N_6051,N_6035);
and U7290 (N_7290,N_6804,N_6034);
nor U7291 (N_7291,N_6593,N_6140);
or U7292 (N_7292,N_6918,N_6858);
or U7293 (N_7293,N_6101,N_6546);
or U7294 (N_7294,N_6520,N_6384);
or U7295 (N_7295,N_6319,N_6791);
or U7296 (N_7296,N_6468,N_6663);
nor U7297 (N_7297,N_6897,N_6487);
and U7298 (N_7298,N_6529,N_6372);
or U7299 (N_7299,N_6788,N_6996);
nor U7300 (N_7300,N_6414,N_6868);
nand U7301 (N_7301,N_6429,N_6961);
nor U7302 (N_7302,N_6571,N_6212);
nand U7303 (N_7303,N_6890,N_6259);
and U7304 (N_7304,N_6005,N_6037);
nor U7305 (N_7305,N_6252,N_6485);
or U7306 (N_7306,N_6790,N_6639);
and U7307 (N_7307,N_6255,N_6163);
and U7308 (N_7308,N_6328,N_6943);
nor U7309 (N_7309,N_6320,N_6634);
xor U7310 (N_7310,N_6187,N_6524);
and U7311 (N_7311,N_6015,N_6157);
and U7312 (N_7312,N_6409,N_6574);
nand U7313 (N_7313,N_6971,N_6318);
and U7314 (N_7314,N_6416,N_6671);
and U7315 (N_7315,N_6940,N_6218);
nand U7316 (N_7316,N_6702,N_6251);
or U7317 (N_7317,N_6507,N_6178);
or U7318 (N_7318,N_6510,N_6491);
nand U7319 (N_7319,N_6348,N_6992);
xnor U7320 (N_7320,N_6851,N_6194);
nor U7321 (N_7321,N_6746,N_6745);
nor U7322 (N_7322,N_6267,N_6664);
or U7323 (N_7323,N_6171,N_6818);
nor U7324 (N_7324,N_6453,N_6500);
nor U7325 (N_7325,N_6763,N_6400);
nand U7326 (N_7326,N_6608,N_6643);
nand U7327 (N_7327,N_6900,N_6921);
or U7328 (N_7328,N_6019,N_6190);
nand U7329 (N_7329,N_6681,N_6741);
or U7330 (N_7330,N_6029,N_6154);
xor U7331 (N_7331,N_6908,N_6582);
and U7332 (N_7332,N_6385,N_6983);
or U7333 (N_7333,N_6193,N_6578);
or U7334 (N_7334,N_6959,N_6027);
xnor U7335 (N_7335,N_6312,N_6381);
and U7336 (N_7336,N_6720,N_6077);
or U7337 (N_7337,N_6228,N_6329);
nand U7338 (N_7338,N_6629,N_6217);
or U7339 (N_7339,N_6754,N_6923);
and U7340 (N_7340,N_6501,N_6304);
or U7341 (N_7341,N_6967,N_6871);
and U7342 (N_7342,N_6070,N_6376);
nand U7343 (N_7343,N_6266,N_6173);
nand U7344 (N_7344,N_6368,N_6805);
or U7345 (N_7345,N_6095,N_6655);
xnor U7346 (N_7346,N_6437,N_6638);
nor U7347 (N_7347,N_6662,N_6929);
nand U7348 (N_7348,N_6738,N_6021);
nor U7349 (N_7349,N_6115,N_6539);
nand U7350 (N_7350,N_6674,N_6565);
or U7351 (N_7351,N_6990,N_6766);
and U7352 (N_7352,N_6657,N_6797);
and U7353 (N_7353,N_6169,N_6094);
or U7354 (N_7354,N_6189,N_6798);
nor U7355 (N_7355,N_6353,N_6056);
and U7356 (N_7356,N_6676,N_6292);
and U7357 (N_7357,N_6459,N_6246);
and U7358 (N_7358,N_6534,N_6721);
or U7359 (N_7359,N_6658,N_6907);
and U7360 (N_7360,N_6446,N_6822);
and U7361 (N_7361,N_6569,N_6642);
or U7362 (N_7362,N_6705,N_6256);
xnor U7363 (N_7363,N_6734,N_6515);
or U7364 (N_7364,N_6610,N_6945);
and U7365 (N_7365,N_6011,N_6248);
or U7366 (N_7366,N_6716,N_6624);
and U7367 (N_7367,N_6964,N_6686);
nand U7368 (N_7368,N_6545,N_6361);
nand U7369 (N_7369,N_6313,N_6463);
nor U7370 (N_7370,N_6098,N_6530);
or U7371 (N_7371,N_6219,N_6158);
xnor U7372 (N_7372,N_6902,N_6423);
and U7373 (N_7373,N_6723,N_6172);
nand U7374 (N_7374,N_6466,N_6707);
or U7375 (N_7375,N_6355,N_6392);
xnor U7376 (N_7376,N_6475,N_6155);
nand U7377 (N_7377,N_6224,N_6867);
nor U7378 (N_7378,N_6830,N_6180);
xor U7379 (N_7379,N_6865,N_6747);
xor U7380 (N_7380,N_6837,N_6080);
or U7381 (N_7381,N_6883,N_6205);
nor U7382 (N_7382,N_6719,N_6787);
and U7383 (N_7383,N_6277,N_6762);
or U7384 (N_7384,N_6421,N_6079);
and U7385 (N_7385,N_6877,N_6411);
and U7386 (N_7386,N_6432,N_6048);
xor U7387 (N_7387,N_6785,N_6229);
and U7388 (N_7388,N_6209,N_6061);
nor U7389 (N_7389,N_6549,N_6936);
nor U7390 (N_7390,N_6020,N_6513);
or U7391 (N_7391,N_6609,N_6684);
nor U7392 (N_7392,N_6424,N_6448);
nand U7393 (N_7393,N_6859,N_6526);
nor U7394 (N_7394,N_6894,N_6306);
nor U7395 (N_7395,N_6612,N_6833);
or U7396 (N_7396,N_6028,N_6147);
and U7397 (N_7397,N_6001,N_6337);
nand U7398 (N_7398,N_6622,N_6519);
or U7399 (N_7399,N_6128,N_6204);
nor U7400 (N_7400,N_6473,N_6960);
nor U7401 (N_7401,N_6717,N_6590);
or U7402 (N_7402,N_6216,N_6692);
and U7403 (N_7403,N_6956,N_6166);
or U7404 (N_7404,N_6291,N_6770);
nand U7405 (N_7405,N_6494,N_6903);
or U7406 (N_7406,N_6339,N_6378);
or U7407 (N_7407,N_6215,N_6043);
or U7408 (N_7408,N_6836,N_6954);
xnor U7409 (N_7409,N_6322,N_6383);
or U7410 (N_7410,N_6369,N_6308);
nor U7411 (N_7411,N_6082,N_6777);
or U7412 (N_7412,N_6068,N_6573);
and U7413 (N_7413,N_6041,N_6863);
and U7414 (N_7414,N_6693,N_6444);
or U7415 (N_7415,N_6206,N_6099);
and U7416 (N_7416,N_6129,N_6017);
or U7417 (N_7417,N_6878,N_6946);
and U7418 (N_7418,N_6401,N_6127);
or U7419 (N_7419,N_6899,N_6697);
and U7420 (N_7420,N_6055,N_6336);
or U7421 (N_7421,N_6425,N_6550);
or U7422 (N_7422,N_6435,N_6748);
and U7423 (N_7423,N_6537,N_6148);
nand U7424 (N_7424,N_6572,N_6185);
and U7425 (N_7425,N_6420,N_6531);
nand U7426 (N_7426,N_6243,N_6953);
nand U7427 (N_7427,N_6668,N_6581);
nand U7428 (N_7428,N_6934,N_6514);
or U7429 (N_7429,N_6831,N_6164);
nor U7430 (N_7430,N_6650,N_6083);
nand U7431 (N_7431,N_6699,N_6834);
nand U7432 (N_7432,N_6407,N_6576);
or U7433 (N_7433,N_6577,N_6091);
nand U7434 (N_7434,N_6214,N_6776);
nand U7435 (N_7435,N_6920,N_6415);
or U7436 (N_7436,N_6580,N_6139);
nor U7437 (N_7437,N_6616,N_6412);
or U7438 (N_7438,N_6326,N_6570);
xor U7439 (N_7439,N_6440,N_6973);
nand U7440 (N_7440,N_6978,N_6845);
and U7441 (N_7441,N_6242,N_6560);
or U7442 (N_7442,N_6038,N_6991);
and U7443 (N_7443,N_6551,N_6768);
and U7444 (N_7444,N_6847,N_6150);
and U7445 (N_7445,N_6236,N_6350);
and U7446 (N_7446,N_6829,N_6025);
nor U7447 (N_7447,N_6467,N_6852);
and U7448 (N_7448,N_6226,N_6223);
xor U7449 (N_7449,N_6484,N_6875);
nand U7450 (N_7450,N_6311,N_6685);
and U7451 (N_7451,N_6044,N_6151);
xor U7452 (N_7452,N_6062,N_6371);
or U7453 (N_7453,N_6840,N_6532);
xor U7454 (N_7454,N_6162,N_6469);
or U7455 (N_7455,N_6288,N_6783);
or U7456 (N_7456,N_6523,N_6359);
nor U7457 (N_7457,N_6439,N_6999);
and U7458 (N_7458,N_6641,N_6977);
nor U7459 (N_7459,N_6273,N_6294);
xnor U7460 (N_7460,N_6989,N_6667);
or U7461 (N_7461,N_6449,N_6253);
nor U7462 (N_7462,N_6138,N_6824);
and U7463 (N_7463,N_6606,N_6970);
xnor U7464 (N_7464,N_6340,N_6880);
nand U7465 (N_7465,N_6315,N_6825);
and U7466 (N_7466,N_6483,N_6703);
xnor U7467 (N_7467,N_6113,N_6715);
and U7468 (N_7468,N_6470,N_6803);
and U7469 (N_7469,N_6656,N_6495);
or U7470 (N_7470,N_6389,N_6284);
xnor U7471 (N_7471,N_6386,N_6645);
xor U7472 (N_7472,N_6191,N_6760);
and U7473 (N_7473,N_6260,N_6682);
nand U7474 (N_7474,N_6419,N_6031);
and U7475 (N_7475,N_6295,N_6103);
nand U7476 (N_7476,N_6177,N_6366);
xnor U7477 (N_7477,N_6321,N_6016);
xor U7478 (N_7478,N_6213,N_6398);
and U7479 (N_7479,N_6711,N_6465);
nor U7480 (N_7480,N_6379,N_6737);
and U7481 (N_7481,N_6556,N_6994);
nand U7482 (N_7482,N_6739,N_6504);
nor U7483 (N_7483,N_6753,N_6422);
nand U7484 (N_7484,N_6922,N_6367);
or U7485 (N_7485,N_6672,N_6764);
nor U7486 (N_7486,N_6695,N_6846);
or U7487 (N_7487,N_6397,N_6841);
nor U7488 (N_7488,N_6085,N_6454);
nor U7489 (N_7489,N_6130,N_6628);
xnor U7490 (N_7490,N_6901,N_6364);
and U7491 (N_7491,N_6388,N_6198);
xor U7492 (N_7492,N_6729,N_6264);
and U7493 (N_7493,N_6694,N_6012);
nand U7494 (N_7494,N_6195,N_6772);
and U7495 (N_7495,N_6636,N_6393);
nor U7496 (N_7496,N_6097,N_6755);
nand U7497 (N_7497,N_6789,N_6912);
nand U7498 (N_7498,N_6434,N_6375);
nand U7499 (N_7499,N_6728,N_6938);
or U7500 (N_7500,N_6169,N_6120);
xor U7501 (N_7501,N_6951,N_6473);
nand U7502 (N_7502,N_6079,N_6254);
or U7503 (N_7503,N_6956,N_6445);
nor U7504 (N_7504,N_6560,N_6951);
or U7505 (N_7505,N_6755,N_6685);
nand U7506 (N_7506,N_6222,N_6690);
or U7507 (N_7507,N_6076,N_6128);
xnor U7508 (N_7508,N_6967,N_6045);
or U7509 (N_7509,N_6825,N_6520);
nand U7510 (N_7510,N_6413,N_6016);
xnor U7511 (N_7511,N_6090,N_6069);
and U7512 (N_7512,N_6631,N_6220);
nand U7513 (N_7513,N_6414,N_6312);
and U7514 (N_7514,N_6693,N_6210);
nand U7515 (N_7515,N_6465,N_6250);
and U7516 (N_7516,N_6727,N_6270);
nor U7517 (N_7517,N_6551,N_6117);
and U7518 (N_7518,N_6760,N_6376);
nor U7519 (N_7519,N_6303,N_6700);
xnor U7520 (N_7520,N_6090,N_6725);
nor U7521 (N_7521,N_6644,N_6075);
or U7522 (N_7522,N_6609,N_6419);
and U7523 (N_7523,N_6047,N_6296);
nand U7524 (N_7524,N_6375,N_6496);
xnor U7525 (N_7525,N_6659,N_6830);
xnor U7526 (N_7526,N_6026,N_6939);
or U7527 (N_7527,N_6882,N_6515);
or U7528 (N_7528,N_6759,N_6152);
and U7529 (N_7529,N_6123,N_6894);
nor U7530 (N_7530,N_6080,N_6345);
nor U7531 (N_7531,N_6679,N_6572);
and U7532 (N_7532,N_6451,N_6591);
or U7533 (N_7533,N_6879,N_6295);
nand U7534 (N_7534,N_6976,N_6166);
xnor U7535 (N_7535,N_6534,N_6553);
or U7536 (N_7536,N_6104,N_6396);
nand U7537 (N_7537,N_6869,N_6755);
xnor U7538 (N_7538,N_6481,N_6195);
nor U7539 (N_7539,N_6177,N_6191);
or U7540 (N_7540,N_6362,N_6517);
nand U7541 (N_7541,N_6546,N_6297);
nor U7542 (N_7542,N_6346,N_6155);
or U7543 (N_7543,N_6329,N_6078);
or U7544 (N_7544,N_6907,N_6568);
nor U7545 (N_7545,N_6246,N_6788);
nor U7546 (N_7546,N_6470,N_6366);
and U7547 (N_7547,N_6342,N_6408);
xnor U7548 (N_7548,N_6330,N_6933);
xnor U7549 (N_7549,N_6866,N_6730);
xnor U7550 (N_7550,N_6540,N_6518);
and U7551 (N_7551,N_6795,N_6225);
xnor U7552 (N_7552,N_6476,N_6676);
or U7553 (N_7553,N_6894,N_6791);
and U7554 (N_7554,N_6033,N_6692);
and U7555 (N_7555,N_6291,N_6250);
and U7556 (N_7556,N_6976,N_6581);
nand U7557 (N_7557,N_6295,N_6631);
and U7558 (N_7558,N_6337,N_6048);
nor U7559 (N_7559,N_6484,N_6981);
nor U7560 (N_7560,N_6668,N_6241);
or U7561 (N_7561,N_6780,N_6523);
and U7562 (N_7562,N_6974,N_6101);
and U7563 (N_7563,N_6764,N_6628);
and U7564 (N_7564,N_6501,N_6535);
nand U7565 (N_7565,N_6086,N_6615);
or U7566 (N_7566,N_6348,N_6210);
nor U7567 (N_7567,N_6030,N_6050);
nor U7568 (N_7568,N_6415,N_6043);
or U7569 (N_7569,N_6318,N_6895);
nand U7570 (N_7570,N_6586,N_6099);
xor U7571 (N_7571,N_6056,N_6075);
xor U7572 (N_7572,N_6876,N_6198);
and U7573 (N_7573,N_6132,N_6475);
nor U7574 (N_7574,N_6907,N_6962);
nor U7575 (N_7575,N_6977,N_6676);
nor U7576 (N_7576,N_6242,N_6665);
or U7577 (N_7577,N_6651,N_6292);
and U7578 (N_7578,N_6348,N_6512);
nor U7579 (N_7579,N_6606,N_6588);
nand U7580 (N_7580,N_6668,N_6917);
nand U7581 (N_7581,N_6322,N_6494);
nand U7582 (N_7582,N_6697,N_6039);
or U7583 (N_7583,N_6221,N_6629);
and U7584 (N_7584,N_6037,N_6878);
or U7585 (N_7585,N_6373,N_6458);
or U7586 (N_7586,N_6149,N_6031);
or U7587 (N_7587,N_6446,N_6282);
or U7588 (N_7588,N_6762,N_6596);
nand U7589 (N_7589,N_6768,N_6010);
and U7590 (N_7590,N_6130,N_6989);
or U7591 (N_7591,N_6392,N_6096);
nor U7592 (N_7592,N_6921,N_6400);
nand U7593 (N_7593,N_6456,N_6297);
nand U7594 (N_7594,N_6014,N_6231);
nand U7595 (N_7595,N_6922,N_6688);
or U7596 (N_7596,N_6296,N_6580);
xor U7597 (N_7597,N_6791,N_6897);
or U7598 (N_7598,N_6013,N_6429);
or U7599 (N_7599,N_6736,N_6290);
or U7600 (N_7600,N_6257,N_6312);
nand U7601 (N_7601,N_6847,N_6988);
nand U7602 (N_7602,N_6563,N_6032);
nand U7603 (N_7603,N_6446,N_6533);
nor U7604 (N_7604,N_6520,N_6864);
and U7605 (N_7605,N_6902,N_6226);
and U7606 (N_7606,N_6578,N_6367);
or U7607 (N_7607,N_6770,N_6848);
nor U7608 (N_7608,N_6406,N_6495);
nor U7609 (N_7609,N_6276,N_6894);
nor U7610 (N_7610,N_6331,N_6575);
and U7611 (N_7611,N_6929,N_6562);
and U7612 (N_7612,N_6750,N_6388);
nand U7613 (N_7613,N_6495,N_6231);
nand U7614 (N_7614,N_6227,N_6862);
nor U7615 (N_7615,N_6191,N_6907);
nor U7616 (N_7616,N_6819,N_6779);
or U7617 (N_7617,N_6483,N_6163);
nand U7618 (N_7618,N_6848,N_6481);
or U7619 (N_7619,N_6617,N_6988);
xor U7620 (N_7620,N_6976,N_6853);
and U7621 (N_7621,N_6660,N_6798);
nor U7622 (N_7622,N_6156,N_6259);
nand U7623 (N_7623,N_6045,N_6754);
nor U7624 (N_7624,N_6089,N_6711);
nor U7625 (N_7625,N_6839,N_6841);
nand U7626 (N_7626,N_6310,N_6735);
nand U7627 (N_7627,N_6585,N_6606);
nand U7628 (N_7628,N_6668,N_6606);
nand U7629 (N_7629,N_6471,N_6938);
nand U7630 (N_7630,N_6708,N_6799);
or U7631 (N_7631,N_6988,N_6829);
or U7632 (N_7632,N_6742,N_6208);
nand U7633 (N_7633,N_6052,N_6060);
or U7634 (N_7634,N_6436,N_6866);
nor U7635 (N_7635,N_6692,N_6578);
nand U7636 (N_7636,N_6874,N_6948);
and U7637 (N_7637,N_6755,N_6727);
nor U7638 (N_7638,N_6556,N_6986);
nor U7639 (N_7639,N_6408,N_6534);
nor U7640 (N_7640,N_6961,N_6677);
xor U7641 (N_7641,N_6931,N_6421);
or U7642 (N_7642,N_6474,N_6293);
nor U7643 (N_7643,N_6748,N_6759);
or U7644 (N_7644,N_6296,N_6585);
and U7645 (N_7645,N_6249,N_6295);
xnor U7646 (N_7646,N_6801,N_6642);
nand U7647 (N_7647,N_6556,N_6327);
or U7648 (N_7648,N_6952,N_6281);
and U7649 (N_7649,N_6302,N_6067);
nand U7650 (N_7650,N_6322,N_6792);
nor U7651 (N_7651,N_6344,N_6371);
nand U7652 (N_7652,N_6639,N_6046);
nand U7653 (N_7653,N_6492,N_6125);
or U7654 (N_7654,N_6066,N_6018);
and U7655 (N_7655,N_6402,N_6726);
or U7656 (N_7656,N_6416,N_6767);
and U7657 (N_7657,N_6923,N_6579);
nor U7658 (N_7658,N_6912,N_6330);
nor U7659 (N_7659,N_6077,N_6740);
nor U7660 (N_7660,N_6365,N_6013);
nor U7661 (N_7661,N_6344,N_6192);
nand U7662 (N_7662,N_6462,N_6912);
nor U7663 (N_7663,N_6507,N_6383);
nor U7664 (N_7664,N_6286,N_6627);
or U7665 (N_7665,N_6297,N_6651);
and U7666 (N_7666,N_6044,N_6069);
nand U7667 (N_7667,N_6414,N_6502);
nor U7668 (N_7668,N_6181,N_6148);
or U7669 (N_7669,N_6851,N_6702);
nor U7670 (N_7670,N_6626,N_6434);
nor U7671 (N_7671,N_6784,N_6539);
or U7672 (N_7672,N_6791,N_6026);
nor U7673 (N_7673,N_6986,N_6093);
nand U7674 (N_7674,N_6011,N_6597);
or U7675 (N_7675,N_6745,N_6638);
and U7676 (N_7676,N_6011,N_6948);
nor U7677 (N_7677,N_6732,N_6516);
nor U7678 (N_7678,N_6704,N_6095);
xnor U7679 (N_7679,N_6959,N_6197);
or U7680 (N_7680,N_6997,N_6559);
or U7681 (N_7681,N_6971,N_6093);
or U7682 (N_7682,N_6943,N_6550);
or U7683 (N_7683,N_6116,N_6281);
or U7684 (N_7684,N_6273,N_6309);
xor U7685 (N_7685,N_6718,N_6055);
nor U7686 (N_7686,N_6612,N_6307);
and U7687 (N_7687,N_6213,N_6223);
or U7688 (N_7688,N_6389,N_6611);
nor U7689 (N_7689,N_6435,N_6326);
and U7690 (N_7690,N_6931,N_6790);
nand U7691 (N_7691,N_6682,N_6350);
or U7692 (N_7692,N_6615,N_6472);
nand U7693 (N_7693,N_6777,N_6487);
or U7694 (N_7694,N_6055,N_6023);
or U7695 (N_7695,N_6964,N_6849);
nor U7696 (N_7696,N_6089,N_6709);
and U7697 (N_7697,N_6108,N_6702);
nand U7698 (N_7698,N_6732,N_6065);
xnor U7699 (N_7699,N_6070,N_6404);
and U7700 (N_7700,N_6300,N_6319);
and U7701 (N_7701,N_6535,N_6852);
and U7702 (N_7702,N_6541,N_6303);
or U7703 (N_7703,N_6365,N_6764);
or U7704 (N_7704,N_6962,N_6501);
nand U7705 (N_7705,N_6466,N_6802);
or U7706 (N_7706,N_6725,N_6386);
nand U7707 (N_7707,N_6485,N_6518);
nand U7708 (N_7708,N_6039,N_6650);
xor U7709 (N_7709,N_6434,N_6263);
nor U7710 (N_7710,N_6068,N_6535);
xnor U7711 (N_7711,N_6542,N_6965);
or U7712 (N_7712,N_6070,N_6652);
nor U7713 (N_7713,N_6004,N_6795);
nand U7714 (N_7714,N_6097,N_6050);
and U7715 (N_7715,N_6632,N_6040);
nand U7716 (N_7716,N_6818,N_6359);
or U7717 (N_7717,N_6084,N_6394);
nand U7718 (N_7718,N_6187,N_6168);
or U7719 (N_7719,N_6968,N_6840);
and U7720 (N_7720,N_6827,N_6949);
nor U7721 (N_7721,N_6269,N_6316);
nand U7722 (N_7722,N_6940,N_6030);
and U7723 (N_7723,N_6822,N_6526);
nor U7724 (N_7724,N_6038,N_6595);
or U7725 (N_7725,N_6865,N_6561);
or U7726 (N_7726,N_6820,N_6019);
nor U7727 (N_7727,N_6705,N_6767);
nor U7728 (N_7728,N_6932,N_6735);
nor U7729 (N_7729,N_6949,N_6952);
xor U7730 (N_7730,N_6610,N_6264);
nor U7731 (N_7731,N_6978,N_6352);
nand U7732 (N_7732,N_6204,N_6615);
or U7733 (N_7733,N_6264,N_6969);
or U7734 (N_7734,N_6261,N_6276);
or U7735 (N_7735,N_6545,N_6425);
or U7736 (N_7736,N_6705,N_6249);
nand U7737 (N_7737,N_6779,N_6247);
and U7738 (N_7738,N_6179,N_6229);
or U7739 (N_7739,N_6758,N_6793);
or U7740 (N_7740,N_6426,N_6097);
and U7741 (N_7741,N_6720,N_6887);
or U7742 (N_7742,N_6140,N_6080);
or U7743 (N_7743,N_6403,N_6604);
nor U7744 (N_7744,N_6603,N_6350);
nor U7745 (N_7745,N_6607,N_6238);
nor U7746 (N_7746,N_6882,N_6498);
or U7747 (N_7747,N_6002,N_6468);
nor U7748 (N_7748,N_6572,N_6189);
xor U7749 (N_7749,N_6307,N_6732);
and U7750 (N_7750,N_6753,N_6268);
xor U7751 (N_7751,N_6669,N_6234);
and U7752 (N_7752,N_6497,N_6654);
xnor U7753 (N_7753,N_6048,N_6029);
or U7754 (N_7754,N_6682,N_6851);
and U7755 (N_7755,N_6594,N_6287);
or U7756 (N_7756,N_6544,N_6625);
and U7757 (N_7757,N_6142,N_6550);
nor U7758 (N_7758,N_6760,N_6805);
or U7759 (N_7759,N_6191,N_6415);
or U7760 (N_7760,N_6996,N_6101);
or U7761 (N_7761,N_6818,N_6013);
and U7762 (N_7762,N_6963,N_6641);
and U7763 (N_7763,N_6677,N_6270);
and U7764 (N_7764,N_6048,N_6159);
or U7765 (N_7765,N_6633,N_6182);
and U7766 (N_7766,N_6153,N_6027);
and U7767 (N_7767,N_6382,N_6163);
and U7768 (N_7768,N_6091,N_6978);
nand U7769 (N_7769,N_6992,N_6262);
nor U7770 (N_7770,N_6656,N_6128);
nand U7771 (N_7771,N_6088,N_6813);
or U7772 (N_7772,N_6237,N_6522);
or U7773 (N_7773,N_6807,N_6997);
xor U7774 (N_7774,N_6671,N_6021);
nor U7775 (N_7775,N_6629,N_6396);
or U7776 (N_7776,N_6265,N_6449);
and U7777 (N_7777,N_6417,N_6250);
or U7778 (N_7778,N_6638,N_6109);
nor U7779 (N_7779,N_6904,N_6459);
nor U7780 (N_7780,N_6822,N_6631);
nand U7781 (N_7781,N_6942,N_6114);
and U7782 (N_7782,N_6387,N_6805);
xor U7783 (N_7783,N_6961,N_6728);
nand U7784 (N_7784,N_6813,N_6406);
nor U7785 (N_7785,N_6564,N_6572);
nand U7786 (N_7786,N_6004,N_6481);
or U7787 (N_7787,N_6641,N_6533);
nand U7788 (N_7788,N_6288,N_6753);
nor U7789 (N_7789,N_6383,N_6019);
nand U7790 (N_7790,N_6021,N_6989);
nor U7791 (N_7791,N_6362,N_6903);
nor U7792 (N_7792,N_6131,N_6533);
and U7793 (N_7793,N_6338,N_6159);
nand U7794 (N_7794,N_6410,N_6250);
and U7795 (N_7795,N_6111,N_6388);
nor U7796 (N_7796,N_6191,N_6113);
nor U7797 (N_7797,N_6724,N_6591);
or U7798 (N_7798,N_6568,N_6667);
or U7799 (N_7799,N_6176,N_6159);
and U7800 (N_7800,N_6578,N_6470);
or U7801 (N_7801,N_6811,N_6098);
or U7802 (N_7802,N_6422,N_6362);
and U7803 (N_7803,N_6291,N_6761);
nand U7804 (N_7804,N_6378,N_6523);
and U7805 (N_7805,N_6083,N_6907);
or U7806 (N_7806,N_6003,N_6793);
nor U7807 (N_7807,N_6276,N_6012);
nor U7808 (N_7808,N_6170,N_6957);
or U7809 (N_7809,N_6146,N_6489);
and U7810 (N_7810,N_6929,N_6925);
or U7811 (N_7811,N_6556,N_6069);
or U7812 (N_7812,N_6159,N_6653);
and U7813 (N_7813,N_6651,N_6097);
xor U7814 (N_7814,N_6935,N_6825);
nand U7815 (N_7815,N_6344,N_6504);
or U7816 (N_7816,N_6024,N_6193);
and U7817 (N_7817,N_6249,N_6957);
or U7818 (N_7818,N_6902,N_6442);
and U7819 (N_7819,N_6501,N_6842);
and U7820 (N_7820,N_6004,N_6003);
and U7821 (N_7821,N_6727,N_6707);
or U7822 (N_7822,N_6551,N_6401);
or U7823 (N_7823,N_6869,N_6611);
nor U7824 (N_7824,N_6767,N_6988);
nor U7825 (N_7825,N_6638,N_6353);
nor U7826 (N_7826,N_6905,N_6453);
nor U7827 (N_7827,N_6004,N_6335);
nor U7828 (N_7828,N_6156,N_6593);
and U7829 (N_7829,N_6945,N_6976);
and U7830 (N_7830,N_6648,N_6922);
nor U7831 (N_7831,N_6692,N_6370);
or U7832 (N_7832,N_6922,N_6601);
nand U7833 (N_7833,N_6789,N_6229);
nor U7834 (N_7834,N_6888,N_6127);
and U7835 (N_7835,N_6802,N_6636);
and U7836 (N_7836,N_6116,N_6887);
and U7837 (N_7837,N_6848,N_6492);
xor U7838 (N_7838,N_6570,N_6166);
nand U7839 (N_7839,N_6560,N_6083);
nand U7840 (N_7840,N_6832,N_6026);
xnor U7841 (N_7841,N_6753,N_6291);
nor U7842 (N_7842,N_6670,N_6918);
nand U7843 (N_7843,N_6564,N_6869);
and U7844 (N_7844,N_6068,N_6652);
xnor U7845 (N_7845,N_6192,N_6082);
nand U7846 (N_7846,N_6435,N_6430);
nand U7847 (N_7847,N_6704,N_6283);
nor U7848 (N_7848,N_6876,N_6067);
and U7849 (N_7849,N_6791,N_6263);
nand U7850 (N_7850,N_6435,N_6112);
nor U7851 (N_7851,N_6443,N_6391);
or U7852 (N_7852,N_6677,N_6855);
or U7853 (N_7853,N_6098,N_6689);
and U7854 (N_7854,N_6342,N_6354);
nand U7855 (N_7855,N_6093,N_6264);
and U7856 (N_7856,N_6077,N_6064);
xor U7857 (N_7857,N_6881,N_6639);
nand U7858 (N_7858,N_6974,N_6908);
nand U7859 (N_7859,N_6673,N_6824);
and U7860 (N_7860,N_6340,N_6515);
nor U7861 (N_7861,N_6698,N_6369);
xnor U7862 (N_7862,N_6723,N_6480);
or U7863 (N_7863,N_6314,N_6832);
or U7864 (N_7864,N_6790,N_6076);
nand U7865 (N_7865,N_6410,N_6097);
nor U7866 (N_7866,N_6135,N_6620);
nor U7867 (N_7867,N_6544,N_6060);
nand U7868 (N_7868,N_6357,N_6086);
or U7869 (N_7869,N_6042,N_6190);
or U7870 (N_7870,N_6136,N_6765);
nor U7871 (N_7871,N_6219,N_6686);
or U7872 (N_7872,N_6981,N_6143);
or U7873 (N_7873,N_6499,N_6824);
or U7874 (N_7874,N_6302,N_6458);
or U7875 (N_7875,N_6088,N_6810);
or U7876 (N_7876,N_6866,N_6940);
nor U7877 (N_7877,N_6775,N_6688);
xor U7878 (N_7878,N_6739,N_6612);
nand U7879 (N_7879,N_6959,N_6451);
and U7880 (N_7880,N_6616,N_6284);
and U7881 (N_7881,N_6019,N_6621);
nor U7882 (N_7882,N_6730,N_6774);
or U7883 (N_7883,N_6777,N_6224);
and U7884 (N_7884,N_6673,N_6591);
or U7885 (N_7885,N_6483,N_6093);
nor U7886 (N_7886,N_6652,N_6488);
xnor U7887 (N_7887,N_6339,N_6498);
xnor U7888 (N_7888,N_6638,N_6903);
and U7889 (N_7889,N_6038,N_6743);
or U7890 (N_7890,N_6268,N_6046);
nor U7891 (N_7891,N_6119,N_6908);
or U7892 (N_7892,N_6130,N_6798);
nand U7893 (N_7893,N_6710,N_6436);
or U7894 (N_7894,N_6507,N_6101);
and U7895 (N_7895,N_6563,N_6405);
nor U7896 (N_7896,N_6295,N_6999);
nand U7897 (N_7897,N_6201,N_6017);
and U7898 (N_7898,N_6157,N_6047);
nor U7899 (N_7899,N_6768,N_6578);
nand U7900 (N_7900,N_6581,N_6333);
nor U7901 (N_7901,N_6872,N_6797);
or U7902 (N_7902,N_6617,N_6236);
or U7903 (N_7903,N_6200,N_6162);
xor U7904 (N_7904,N_6553,N_6576);
or U7905 (N_7905,N_6567,N_6737);
nor U7906 (N_7906,N_6322,N_6605);
nand U7907 (N_7907,N_6750,N_6292);
or U7908 (N_7908,N_6280,N_6375);
nor U7909 (N_7909,N_6472,N_6518);
and U7910 (N_7910,N_6781,N_6903);
nand U7911 (N_7911,N_6670,N_6429);
nand U7912 (N_7912,N_6949,N_6283);
nor U7913 (N_7913,N_6856,N_6885);
nand U7914 (N_7914,N_6699,N_6503);
nor U7915 (N_7915,N_6170,N_6159);
and U7916 (N_7916,N_6607,N_6549);
nand U7917 (N_7917,N_6209,N_6066);
and U7918 (N_7918,N_6009,N_6023);
nor U7919 (N_7919,N_6148,N_6078);
and U7920 (N_7920,N_6012,N_6383);
or U7921 (N_7921,N_6345,N_6521);
or U7922 (N_7922,N_6429,N_6730);
or U7923 (N_7923,N_6423,N_6711);
or U7924 (N_7924,N_6624,N_6549);
and U7925 (N_7925,N_6977,N_6902);
and U7926 (N_7926,N_6797,N_6512);
or U7927 (N_7927,N_6713,N_6314);
nor U7928 (N_7928,N_6022,N_6569);
nand U7929 (N_7929,N_6485,N_6031);
nor U7930 (N_7930,N_6466,N_6353);
nand U7931 (N_7931,N_6246,N_6441);
xnor U7932 (N_7932,N_6244,N_6165);
xnor U7933 (N_7933,N_6127,N_6411);
nor U7934 (N_7934,N_6423,N_6552);
or U7935 (N_7935,N_6300,N_6113);
nor U7936 (N_7936,N_6682,N_6956);
xnor U7937 (N_7937,N_6708,N_6687);
nand U7938 (N_7938,N_6164,N_6418);
nand U7939 (N_7939,N_6550,N_6735);
nor U7940 (N_7940,N_6248,N_6536);
and U7941 (N_7941,N_6937,N_6936);
nand U7942 (N_7942,N_6562,N_6043);
nand U7943 (N_7943,N_6662,N_6410);
xor U7944 (N_7944,N_6194,N_6585);
and U7945 (N_7945,N_6179,N_6543);
nand U7946 (N_7946,N_6370,N_6192);
nand U7947 (N_7947,N_6884,N_6210);
nand U7948 (N_7948,N_6577,N_6131);
nand U7949 (N_7949,N_6964,N_6434);
xnor U7950 (N_7950,N_6178,N_6545);
nor U7951 (N_7951,N_6294,N_6692);
nand U7952 (N_7952,N_6795,N_6992);
and U7953 (N_7953,N_6454,N_6296);
xor U7954 (N_7954,N_6789,N_6327);
and U7955 (N_7955,N_6541,N_6312);
nor U7956 (N_7956,N_6728,N_6707);
nand U7957 (N_7957,N_6722,N_6349);
or U7958 (N_7958,N_6931,N_6814);
and U7959 (N_7959,N_6295,N_6543);
or U7960 (N_7960,N_6491,N_6162);
nand U7961 (N_7961,N_6458,N_6659);
nand U7962 (N_7962,N_6163,N_6685);
or U7963 (N_7963,N_6186,N_6936);
and U7964 (N_7964,N_6218,N_6848);
nor U7965 (N_7965,N_6196,N_6748);
or U7966 (N_7966,N_6248,N_6696);
or U7967 (N_7967,N_6909,N_6395);
nor U7968 (N_7968,N_6408,N_6720);
or U7969 (N_7969,N_6875,N_6966);
and U7970 (N_7970,N_6084,N_6876);
and U7971 (N_7971,N_6643,N_6753);
or U7972 (N_7972,N_6003,N_6001);
nor U7973 (N_7973,N_6920,N_6634);
and U7974 (N_7974,N_6972,N_6559);
nor U7975 (N_7975,N_6537,N_6399);
and U7976 (N_7976,N_6990,N_6941);
nor U7977 (N_7977,N_6248,N_6717);
nand U7978 (N_7978,N_6966,N_6458);
xnor U7979 (N_7979,N_6639,N_6364);
and U7980 (N_7980,N_6318,N_6938);
xor U7981 (N_7981,N_6525,N_6141);
and U7982 (N_7982,N_6288,N_6738);
nor U7983 (N_7983,N_6034,N_6781);
and U7984 (N_7984,N_6742,N_6617);
and U7985 (N_7985,N_6239,N_6476);
nor U7986 (N_7986,N_6320,N_6359);
and U7987 (N_7987,N_6313,N_6887);
and U7988 (N_7988,N_6472,N_6422);
or U7989 (N_7989,N_6685,N_6917);
nand U7990 (N_7990,N_6276,N_6247);
and U7991 (N_7991,N_6431,N_6267);
nand U7992 (N_7992,N_6605,N_6577);
and U7993 (N_7993,N_6307,N_6345);
xor U7994 (N_7994,N_6505,N_6767);
and U7995 (N_7995,N_6625,N_6665);
or U7996 (N_7996,N_6727,N_6316);
and U7997 (N_7997,N_6530,N_6169);
nor U7998 (N_7998,N_6150,N_6674);
or U7999 (N_7999,N_6997,N_6145);
or U8000 (N_8000,N_7071,N_7215);
or U8001 (N_8001,N_7683,N_7355);
nand U8002 (N_8002,N_7765,N_7196);
or U8003 (N_8003,N_7781,N_7570);
and U8004 (N_8004,N_7663,N_7508);
nand U8005 (N_8005,N_7477,N_7268);
nor U8006 (N_8006,N_7396,N_7918);
nand U8007 (N_8007,N_7757,N_7173);
nor U8008 (N_8008,N_7401,N_7271);
nand U8009 (N_8009,N_7133,N_7790);
nand U8010 (N_8010,N_7548,N_7564);
nand U8011 (N_8011,N_7599,N_7277);
nor U8012 (N_8012,N_7189,N_7245);
nor U8013 (N_8013,N_7398,N_7300);
xor U8014 (N_8014,N_7090,N_7574);
nand U8015 (N_8015,N_7719,N_7014);
and U8016 (N_8016,N_7280,N_7169);
nor U8017 (N_8017,N_7136,N_7659);
or U8018 (N_8018,N_7038,N_7550);
and U8019 (N_8019,N_7875,N_7655);
or U8020 (N_8020,N_7129,N_7710);
and U8021 (N_8021,N_7382,N_7160);
nand U8022 (N_8022,N_7664,N_7483);
nor U8023 (N_8023,N_7876,N_7638);
or U8024 (N_8024,N_7920,N_7461);
and U8025 (N_8025,N_7950,N_7510);
or U8026 (N_8026,N_7403,N_7054);
nor U8027 (N_8027,N_7528,N_7732);
nand U8028 (N_8028,N_7715,N_7122);
nand U8029 (N_8029,N_7837,N_7946);
nor U8030 (N_8030,N_7368,N_7824);
and U8031 (N_8031,N_7413,N_7163);
or U8032 (N_8032,N_7526,N_7421);
and U8033 (N_8033,N_7834,N_7285);
or U8034 (N_8034,N_7767,N_7417);
xnor U8035 (N_8035,N_7956,N_7456);
and U8036 (N_8036,N_7220,N_7546);
and U8037 (N_8037,N_7035,N_7385);
nand U8038 (N_8038,N_7282,N_7430);
and U8039 (N_8039,N_7606,N_7545);
nand U8040 (N_8040,N_7185,N_7935);
and U8041 (N_8041,N_7747,N_7411);
or U8042 (N_8042,N_7378,N_7549);
nor U8043 (N_8043,N_7206,N_7869);
or U8044 (N_8044,N_7472,N_7001);
nand U8045 (N_8045,N_7375,N_7340);
nor U8046 (N_8046,N_7441,N_7449);
nand U8047 (N_8047,N_7958,N_7697);
nor U8048 (N_8048,N_7119,N_7709);
and U8049 (N_8049,N_7429,N_7082);
or U8050 (N_8050,N_7888,N_7877);
nor U8051 (N_8051,N_7974,N_7825);
nor U8052 (N_8052,N_7476,N_7512);
nor U8053 (N_8053,N_7514,N_7819);
nor U8054 (N_8054,N_7543,N_7162);
nand U8055 (N_8055,N_7776,N_7165);
or U8056 (N_8056,N_7726,N_7433);
nand U8057 (N_8057,N_7644,N_7835);
nand U8058 (N_8058,N_7575,N_7089);
and U8059 (N_8059,N_7399,N_7467);
nand U8060 (N_8060,N_7903,N_7839);
nand U8061 (N_8061,N_7395,N_7681);
xnor U8062 (N_8062,N_7390,N_7147);
nor U8063 (N_8063,N_7808,N_7130);
xor U8064 (N_8064,N_7093,N_7642);
nand U8065 (N_8065,N_7507,N_7144);
or U8066 (N_8066,N_7931,N_7897);
and U8067 (N_8067,N_7474,N_7986);
nand U8068 (N_8068,N_7496,N_7034);
nor U8069 (N_8069,N_7198,N_7096);
or U8070 (N_8070,N_7112,N_7070);
nand U8071 (N_8071,N_7556,N_7813);
nor U8072 (N_8072,N_7088,N_7343);
nand U8073 (N_8073,N_7754,N_7000);
and U8074 (N_8074,N_7774,N_7454);
nor U8075 (N_8075,N_7468,N_7370);
and U8076 (N_8076,N_7745,N_7306);
and U8077 (N_8077,N_7730,N_7311);
nand U8078 (N_8078,N_7928,N_7424);
nor U8079 (N_8079,N_7572,N_7404);
or U8080 (N_8080,N_7565,N_7366);
nor U8081 (N_8081,N_7201,N_7797);
or U8082 (N_8082,N_7436,N_7979);
xor U8083 (N_8083,N_7077,N_7870);
nor U8084 (N_8084,N_7110,N_7019);
nor U8085 (N_8085,N_7566,N_7900);
nor U8086 (N_8086,N_7831,N_7039);
or U8087 (N_8087,N_7867,N_7651);
and U8088 (N_8088,N_7631,N_7209);
nor U8089 (N_8089,N_7256,N_7252);
and U8090 (N_8090,N_7041,N_7911);
nand U8091 (N_8091,N_7585,N_7624);
or U8092 (N_8092,N_7978,N_7955);
and U8093 (N_8093,N_7905,N_7637);
nand U8094 (N_8094,N_7324,N_7031);
nand U8095 (N_8095,N_7380,N_7455);
and U8096 (N_8096,N_7260,N_7348);
or U8097 (N_8097,N_7578,N_7587);
or U8098 (N_8098,N_7632,N_7591);
nand U8099 (N_8099,N_7061,N_7672);
nand U8100 (N_8100,N_7314,N_7316);
and U8101 (N_8101,N_7018,N_7191);
nor U8102 (N_8102,N_7742,N_7864);
or U8103 (N_8103,N_7750,N_7361);
and U8104 (N_8104,N_7751,N_7002);
nand U8105 (N_8105,N_7836,N_7749);
nand U8106 (N_8106,N_7713,N_7722);
nand U8107 (N_8107,N_7091,N_7502);
or U8108 (N_8108,N_7109,N_7301);
xor U8109 (N_8109,N_7878,N_7051);
and U8110 (N_8110,N_7278,N_7418);
nand U8111 (N_8111,N_7581,N_7064);
and U8112 (N_8112,N_7701,N_7434);
nor U8113 (N_8113,N_7953,N_7707);
and U8114 (N_8114,N_7970,N_7973);
or U8115 (N_8115,N_7297,N_7762);
nor U8116 (N_8116,N_7753,N_7580);
and U8117 (N_8117,N_7519,N_7919);
and U8118 (N_8118,N_7805,N_7120);
nor U8119 (N_8119,N_7597,N_7407);
or U8120 (N_8120,N_7717,N_7907);
nand U8121 (N_8121,N_7138,N_7636);
xnor U8122 (N_8122,N_7254,N_7296);
and U8123 (N_8123,N_7320,N_7352);
nor U8124 (N_8124,N_7678,N_7536);
or U8125 (N_8125,N_7617,N_7299);
nand U8126 (N_8126,N_7902,N_7858);
nand U8127 (N_8127,N_7972,N_7854);
or U8128 (N_8128,N_7230,N_7229);
nor U8129 (N_8129,N_7339,N_7036);
and U8130 (N_8130,N_7304,N_7076);
or U8131 (N_8131,N_7965,N_7557);
and U8132 (N_8132,N_7438,N_7537);
or U8133 (N_8133,N_7239,N_7298);
or U8134 (N_8134,N_7116,N_7621);
and U8135 (N_8135,N_7504,N_7139);
xnor U8136 (N_8136,N_7272,N_7576);
or U8137 (N_8137,N_7459,N_7097);
nand U8138 (N_8138,N_7987,N_7952);
and U8139 (N_8139,N_7111,N_7688);
or U8140 (N_8140,N_7086,N_7547);
nand U8141 (N_8141,N_7029,N_7971);
and U8142 (N_8142,N_7107,N_7243);
and U8143 (N_8143,N_7182,N_7552);
and U8144 (N_8144,N_7609,N_7143);
or U8145 (N_8145,N_7253,N_7698);
nand U8146 (N_8146,N_7703,N_7588);
xnor U8147 (N_8147,N_7479,N_7208);
nand U8148 (N_8148,N_7328,N_7675);
or U8149 (N_8149,N_7095,N_7889);
or U8150 (N_8150,N_7880,N_7326);
or U8151 (N_8151,N_7569,N_7851);
nor U8152 (N_8152,N_7553,N_7855);
and U8153 (N_8153,N_7170,N_7319);
or U8154 (N_8154,N_7440,N_7224);
and U8155 (N_8155,N_7665,N_7148);
and U8156 (N_8156,N_7234,N_7988);
or U8157 (N_8157,N_7737,N_7026);
nor U8158 (N_8158,N_7293,N_7981);
nor U8159 (N_8159,N_7168,N_7778);
and U8160 (N_8160,N_7210,N_7821);
and U8161 (N_8161,N_7481,N_7446);
or U8162 (N_8162,N_7108,N_7011);
and U8163 (N_8163,N_7786,N_7740);
and U8164 (N_8164,N_7735,N_7025);
xnor U8165 (N_8165,N_7693,N_7844);
and U8166 (N_8166,N_7099,N_7596);
and U8167 (N_8167,N_7893,N_7799);
or U8168 (N_8168,N_7012,N_7241);
xnor U8169 (N_8169,N_7680,N_7194);
nand U8170 (N_8170,N_7992,N_7305);
nand U8171 (N_8171,N_7323,N_7712);
nor U8172 (N_8172,N_7392,N_7998);
or U8173 (N_8173,N_7906,N_7346);
nand U8174 (N_8174,N_7419,N_7968);
and U8175 (N_8175,N_7336,N_7460);
or U8176 (N_8176,N_7167,N_7977);
nor U8177 (N_8177,N_7743,N_7338);
xor U8178 (N_8178,N_7330,N_7529);
or U8179 (N_8179,N_7866,N_7374);
nor U8180 (N_8180,N_7535,N_7629);
xor U8181 (N_8181,N_7333,N_7846);
and U8182 (N_8182,N_7444,N_7145);
nand U8183 (N_8183,N_7179,N_7830);
nand U8184 (N_8184,N_7691,N_7388);
nand U8185 (N_8185,N_7595,N_7868);
and U8186 (N_8186,N_7004,N_7222);
or U8187 (N_8187,N_7020,N_7945);
and U8188 (N_8188,N_7817,N_7639);
nor U8189 (N_8189,N_7544,N_7685);
nand U8190 (N_8190,N_7793,N_7727);
nand U8191 (N_8191,N_7066,N_7792);
nor U8192 (N_8192,N_7933,N_7290);
and U8193 (N_8193,N_7690,N_7416);
nor U8194 (N_8194,N_7258,N_7431);
xnor U8195 (N_8195,N_7190,N_7860);
nand U8196 (N_8196,N_7859,N_7376);
xor U8197 (N_8197,N_7197,N_7373);
and U8198 (N_8198,N_7627,N_7729);
nor U8199 (N_8199,N_7648,N_7003);
or U8200 (N_8200,N_7501,N_7497);
nand U8201 (N_8201,N_7708,N_7265);
nor U8202 (N_8202,N_7892,N_7980);
or U8203 (N_8203,N_7223,N_7493);
nor U8204 (N_8204,N_7957,N_7761);
nor U8205 (N_8205,N_7153,N_7882);
nor U8206 (N_8206,N_7775,N_7056);
nor U8207 (N_8207,N_7414,N_7803);
or U8208 (N_8208,N_7848,N_7563);
nor U8209 (N_8209,N_7159,N_7873);
nor U8210 (N_8210,N_7721,N_7006);
nor U8211 (N_8211,N_7983,N_7849);
or U8212 (N_8212,N_7723,N_7604);
nor U8213 (N_8213,N_7562,N_7826);
xor U8214 (N_8214,N_7852,N_7647);
and U8215 (N_8215,N_7755,N_7287);
xnor U8216 (N_8216,N_7068,N_7522);
xor U8217 (N_8217,N_7841,N_7871);
and U8218 (N_8218,N_7538,N_7515);
nand U8219 (N_8219,N_7270,N_7827);
xor U8220 (N_8220,N_7009,N_7353);
nand U8221 (N_8221,N_7505,N_7037);
and U8222 (N_8222,N_7807,N_7259);
nor U8223 (N_8223,N_7480,N_7427);
nand U8224 (N_8224,N_7042,N_7049);
nand U8225 (N_8225,N_7771,N_7023);
or U8226 (N_8226,N_7518,N_7887);
and U8227 (N_8227,N_7211,N_7541);
nor U8228 (N_8228,N_7227,N_7135);
or U8229 (N_8229,N_7065,N_7113);
xnor U8230 (N_8230,N_7787,N_7125);
and U8231 (N_8231,N_7796,N_7758);
or U8232 (N_8232,N_7250,N_7532);
and U8233 (N_8233,N_7117,N_7458);
and U8234 (N_8234,N_7509,N_7842);
or U8235 (N_8235,N_7612,N_7608);
and U8236 (N_8236,N_7325,N_7393);
xor U8237 (N_8237,N_7985,N_7628);
xor U8238 (N_8238,N_7815,N_7660);
and U8239 (N_8239,N_7534,N_7498);
xnor U8240 (N_8240,N_7262,N_7798);
nor U8241 (N_8241,N_7577,N_7816);
nand U8242 (N_8242,N_7982,N_7275);
or U8243 (N_8243,N_7804,N_7360);
or U8244 (N_8244,N_7976,N_7236);
nor U8245 (N_8245,N_7856,N_7890);
and U8246 (N_8246,N_7412,N_7752);
or U8247 (N_8247,N_7058,N_7074);
nor U8248 (N_8248,N_7073,N_7050);
nor U8249 (N_8249,N_7788,N_7590);
or U8250 (N_8250,N_7216,N_7668);
nand U8251 (N_8251,N_7200,N_7178);
xnor U8252 (N_8252,N_7760,N_7207);
nor U8253 (N_8253,N_7315,N_7674);
nand U8254 (N_8254,N_7212,N_7415);
and U8255 (N_8255,N_7769,N_7488);
nand U8256 (N_8256,N_7499,N_7180);
xnor U8257 (N_8257,N_7598,N_7266);
nor U8258 (N_8258,N_7643,N_7601);
and U8259 (N_8259,N_7923,N_7267);
and U8260 (N_8260,N_7115,N_7756);
and U8261 (N_8261,N_7202,N_7818);
nor U8262 (N_8262,N_7962,N_7341);
nor U8263 (N_8263,N_7473,N_7464);
and U8264 (N_8264,N_7630,N_7832);
nor U8265 (N_8265,N_7150,N_7308);
nand U8266 (N_8266,N_7137,N_7883);
xor U8267 (N_8267,N_7810,N_7937);
and U8268 (N_8268,N_7055,N_7925);
nor U8269 (N_8269,N_7913,N_7344);
nand U8270 (N_8270,N_7232,N_7914);
nand U8271 (N_8271,N_7533,N_7022);
nand U8272 (N_8272,N_7874,N_7641);
nand U8273 (N_8273,N_7432,N_7741);
xnor U8274 (N_8274,N_7045,N_7181);
nor U8275 (N_8275,N_7235,N_7838);
xor U8276 (N_8276,N_7205,N_7661);
or U8277 (N_8277,N_7166,N_7184);
and U8278 (N_8278,N_7284,N_7291);
nand U8279 (N_8279,N_7809,N_7782);
xor U8280 (N_8280,N_7695,N_7899);
nand U8281 (N_8281,N_7938,N_7586);
or U8282 (N_8282,N_7164,N_7583);
xor U8283 (N_8283,N_7731,N_7802);
or U8284 (N_8284,N_7635,N_7462);
nor U8285 (N_8285,N_7008,N_7611);
nand U8286 (N_8286,N_7240,N_7622);
nand U8287 (N_8287,N_7186,N_7062);
xnor U8288 (N_8288,N_7584,N_7289);
or U8289 (N_8289,N_7199,N_7482);
and U8290 (N_8290,N_7420,N_7218);
nor U8291 (N_8291,N_7397,N_7523);
and U8292 (N_8292,N_7244,N_7439);
nor U8293 (N_8293,N_7540,N_7142);
nor U8294 (N_8294,N_7724,N_7487);
xnor U8295 (N_8295,N_7384,N_7466);
nor U8296 (N_8296,N_7942,N_7669);
and U8297 (N_8297,N_7307,N_7996);
or U8298 (N_8298,N_7939,N_7383);
and U8299 (N_8299,N_7030,N_7356);
or U8300 (N_8300,N_7118,N_7806);
or U8301 (N_8301,N_7005,N_7963);
nor U8302 (N_8302,N_7387,N_7362);
and U8303 (N_8303,N_7673,N_7060);
nand U8304 (N_8304,N_7865,N_7936);
nand U8305 (N_8305,N_7885,N_7204);
xnor U8306 (N_8306,N_7657,N_7896);
or U8307 (N_8307,N_7171,N_7400);
or U8308 (N_8308,N_7850,N_7377);
xor U8309 (N_8309,N_7716,N_7350);
or U8310 (N_8310,N_7530,N_7469);
xnor U8311 (N_8311,N_7152,N_7554);
and U8312 (N_8312,N_7312,N_7491);
and U8313 (N_8313,N_7746,N_7379);
xnor U8314 (N_8314,N_7967,N_7531);
and U8315 (N_8315,N_7465,N_7520);
nand U8316 (N_8316,N_7475,N_7862);
nor U8317 (N_8317,N_7910,N_7149);
nor U8318 (N_8318,N_7525,N_7650);
and U8319 (N_8319,N_7898,N_7126);
nand U8320 (N_8320,N_7934,N_7155);
or U8321 (N_8321,N_7511,N_7335);
nand U8322 (N_8322,N_7524,N_7921);
and U8323 (N_8323,N_7052,N_7121);
and U8324 (N_8324,N_7784,N_7246);
nand U8325 (N_8325,N_7156,N_7561);
or U8326 (N_8326,N_7711,N_7895);
and U8327 (N_8327,N_7423,N_7221);
nor U8328 (N_8328,N_7013,N_7706);
nor U8329 (N_8329,N_7555,N_7948);
nor U8330 (N_8330,N_7408,N_7010);
nor U8331 (N_8331,N_7600,N_7264);
or U8332 (N_8332,N_7527,N_7733);
and U8333 (N_8333,N_7916,N_7046);
or U8334 (N_8334,N_7327,N_7302);
or U8335 (N_8335,N_7990,N_7684);
xor U8336 (N_8336,N_7559,N_7457);
nand U8337 (N_8337,N_7195,N_7947);
or U8338 (N_8338,N_7909,N_7357);
or U8339 (N_8339,N_7822,N_7364);
and U8340 (N_8340,N_7944,N_7917);
and U8341 (N_8341,N_7884,N_7800);
or U8342 (N_8342,N_7106,N_7174);
nand U8343 (N_8343,N_7791,N_7059);
nor U8344 (N_8344,N_7242,N_7228);
nor U8345 (N_8345,N_7394,N_7739);
nand U8346 (N_8346,N_7975,N_7941);
and U8347 (N_8347,N_7367,N_7331);
or U8348 (N_8348,N_7605,N_7078);
xnor U8349 (N_8349,N_7640,N_7063);
nand U8350 (N_8350,N_7853,N_7687);
nor U8351 (N_8351,N_7613,N_7248);
nor U8352 (N_8352,N_7620,N_7927);
and U8353 (N_8353,N_7484,N_7828);
or U8354 (N_8354,N_7705,N_7105);
nand U8355 (N_8355,N_7704,N_7615);
and U8356 (N_8356,N_7653,N_7676);
or U8357 (N_8357,N_7104,N_7682);
nand U8358 (N_8358,N_7463,N_7568);
or U8359 (N_8359,N_7677,N_7017);
nor U8360 (N_8360,N_7114,N_7351);
nand U8361 (N_8361,N_7292,N_7225);
or U8362 (N_8362,N_7214,N_7219);
nor U8363 (N_8363,N_7542,N_7551);
nand U8364 (N_8364,N_7579,N_7334);
or U8365 (N_8365,N_7666,N_7625);
and U8366 (N_8366,N_7649,N_7513);
or U8367 (N_8367,N_7177,N_7768);
or U8368 (N_8368,N_7217,N_7633);
nand U8369 (N_8369,N_7043,N_7671);
or U8370 (N_8370,N_7738,N_7226);
nor U8371 (N_8371,N_7007,N_7718);
or U8372 (N_8372,N_7273,N_7506);
nor U8373 (N_8373,N_7820,N_7833);
and U8374 (N_8374,N_7085,N_7053);
xor U8375 (N_8375,N_7485,N_7966);
or U8376 (N_8376,N_7881,N_7623);
nand U8377 (N_8377,N_7626,N_7363);
nor U8378 (N_8378,N_7069,N_7904);
xor U8379 (N_8379,N_7571,N_7961);
and U8380 (N_8380,N_7779,N_7686);
nor U8381 (N_8381,N_7098,N_7645);
or U8382 (N_8382,N_7389,N_7175);
nand U8383 (N_8383,N_7471,N_7470);
nor U8384 (N_8384,N_7132,N_7764);
and U8385 (N_8385,N_7080,N_7789);
and U8386 (N_8386,N_7829,N_7402);
or U8387 (N_8387,N_7773,N_7172);
xor U8388 (N_8388,N_7814,N_7453);
nand U8389 (N_8389,N_7193,N_7154);
and U8390 (N_8390,N_7894,N_7517);
and U8391 (N_8391,N_7692,N_7321);
or U8392 (N_8392,N_7322,N_7354);
and U8393 (N_8393,N_7616,N_7539);
nand U8394 (N_8394,N_7696,N_7081);
nor U8395 (N_8395,N_7728,N_7342);
nand U8396 (N_8396,N_7329,N_7734);
or U8397 (N_8397,N_7083,N_7263);
nand U8398 (N_8398,N_7161,N_7072);
nor U8399 (N_8399,N_7840,N_7103);
and U8400 (N_8400,N_7603,N_7087);
and U8401 (N_8401,N_7100,N_7646);
or U8402 (N_8402,N_7811,N_7075);
nand U8403 (N_8403,N_7593,N_7780);
nand U8404 (N_8404,N_7619,N_7192);
nand U8405 (N_8405,N_7028,N_7237);
xnor U8406 (N_8406,N_7954,N_7261);
xnor U8407 (N_8407,N_7024,N_7908);
nor U8408 (N_8408,N_7123,N_7255);
and U8409 (N_8409,N_7929,N_7067);
nor U8410 (N_8410,N_7592,N_7332);
xor U8411 (N_8411,N_7656,N_7614);
xnor U8412 (N_8412,N_7922,N_7251);
or U8413 (N_8413,N_7309,N_7924);
nor U8414 (N_8414,N_7318,N_7288);
nor U8415 (N_8415,N_7274,N_7079);
and U8416 (N_8416,N_7405,N_7140);
or U8417 (N_8417,N_7926,N_7618);
nor U8418 (N_8418,N_7092,N_7188);
nand U8419 (N_8419,N_7203,N_7759);
and U8420 (N_8420,N_7033,N_7406);
nor U8421 (N_8421,N_7032,N_7714);
or U8422 (N_8422,N_7447,N_7422);
nor U8423 (N_8423,N_7999,N_7901);
nand U8424 (N_8424,N_7516,N_7951);
and U8425 (N_8425,N_7993,N_7448);
nand U8426 (N_8426,N_7594,N_7879);
and U8427 (N_8427,N_7658,N_7128);
and U8428 (N_8428,N_7233,N_7286);
or U8429 (N_8429,N_7358,N_7748);
xnor U8430 (N_8430,N_7409,N_7964);
and U8431 (N_8431,N_7634,N_7694);
nand U8432 (N_8432,N_7847,N_7812);
nor U8433 (N_8433,N_7047,N_7744);
xor U8434 (N_8434,N_7146,N_7391);
and U8435 (N_8435,N_7369,N_7720);
nor U8436 (N_8436,N_7558,N_7699);
nor U8437 (N_8437,N_7560,N_7021);
nor U8438 (N_8438,N_7607,N_7969);
nand U8439 (N_8439,N_7127,N_7158);
and U8440 (N_8440,N_7213,N_7365);
nor U8441 (N_8441,N_7295,N_7777);
nor U8442 (N_8442,N_7176,N_7503);
and U8443 (N_8443,N_7281,N_7959);
nand U8444 (N_8444,N_7845,N_7231);
and U8445 (N_8445,N_7801,N_7303);
nand U8446 (N_8446,N_7861,N_7451);
or U8447 (N_8447,N_7843,N_7437);
nor U8448 (N_8448,N_7667,N_7700);
and U8449 (N_8449,N_7489,N_7371);
or U8450 (N_8450,N_7381,N_7763);
or U8451 (N_8451,N_7016,N_7442);
xor U8452 (N_8452,N_7101,N_7102);
and U8453 (N_8453,N_7766,N_7269);
nor U8454 (N_8454,N_7486,N_7991);
and U8455 (N_8455,N_7943,N_7567);
nor U8456 (N_8456,N_7347,N_7094);
xnor U8457 (N_8457,N_7725,N_7349);
and U8458 (N_8458,N_7187,N_7582);
and U8459 (N_8459,N_7932,N_7915);
and U8460 (N_8460,N_7772,N_7048);
and U8461 (N_8461,N_7151,N_7960);
nand U8462 (N_8462,N_7589,N_7997);
or U8463 (N_8463,N_7794,N_7426);
nor U8464 (N_8464,N_7317,N_7410);
or U8465 (N_8465,N_7652,N_7238);
xnor U8466 (N_8466,N_7602,N_7654);
xor U8467 (N_8467,N_7863,N_7823);
nand U8468 (N_8468,N_7891,N_7495);
and U8469 (N_8469,N_7134,N_7492);
or U8470 (N_8470,N_7500,N_7886);
or U8471 (N_8471,N_7027,N_7940);
or U8472 (N_8472,N_7872,N_7736);
and U8473 (N_8473,N_7279,N_7247);
and U8474 (N_8474,N_7450,N_7989);
nand U8475 (N_8475,N_7995,N_7057);
nand U8476 (N_8476,N_7702,N_7345);
and U8477 (N_8477,N_7478,N_7452);
or U8478 (N_8478,N_7679,N_7183);
and U8479 (N_8479,N_7044,N_7912);
or U8480 (N_8480,N_7015,N_7783);
nor U8481 (N_8481,N_7276,N_7662);
or U8482 (N_8482,N_7610,N_7573);
nor U8483 (N_8483,N_7372,N_7249);
nand U8484 (N_8484,N_7930,N_7443);
or U8485 (N_8485,N_7131,N_7984);
or U8486 (N_8486,N_7124,N_7157);
nor U8487 (N_8487,N_7040,N_7313);
nor U8488 (N_8488,N_7795,N_7257);
or U8489 (N_8489,N_7310,N_7386);
and U8490 (N_8490,N_7359,N_7141);
nor U8491 (N_8491,N_7283,N_7857);
nand U8492 (N_8492,N_7689,N_7428);
or U8493 (N_8493,N_7670,N_7994);
nor U8494 (N_8494,N_7337,N_7435);
xnor U8495 (N_8495,N_7785,N_7294);
nor U8496 (N_8496,N_7949,N_7521);
xor U8497 (N_8497,N_7770,N_7445);
or U8498 (N_8498,N_7084,N_7494);
nand U8499 (N_8499,N_7425,N_7490);
nand U8500 (N_8500,N_7591,N_7388);
or U8501 (N_8501,N_7432,N_7187);
and U8502 (N_8502,N_7772,N_7780);
nand U8503 (N_8503,N_7838,N_7001);
xnor U8504 (N_8504,N_7634,N_7656);
xnor U8505 (N_8505,N_7233,N_7570);
nor U8506 (N_8506,N_7902,N_7767);
nor U8507 (N_8507,N_7526,N_7410);
nor U8508 (N_8508,N_7414,N_7639);
and U8509 (N_8509,N_7715,N_7930);
nor U8510 (N_8510,N_7125,N_7448);
nand U8511 (N_8511,N_7581,N_7434);
nand U8512 (N_8512,N_7048,N_7246);
and U8513 (N_8513,N_7150,N_7143);
and U8514 (N_8514,N_7601,N_7067);
nand U8515 (N_8515,N_7018,N_7428);
or U8516 (N_8516,N_7921,N_7776);
and U8517 (N_8517,N_7268,N_7194);
nand U8518 (N_8518,N_7240,N_7806);
nand U8519 (N_8519,N_7655,N_7783);
nand U8520 (N_8520,N_7131,N_7633);
and U8521 (N_8521,N_7850,N_7021);
xor U8522 (N_8522,N_7084,N_7166);
xor U8523 (N_8523,N_7226,N_7419);
nand U8524 (N_8524,N_7738,N_7061);
and U8525 (N_8525,N_7251,N_7523);
nor U8526 (N_8526,N_7392,N_7359);
or U8527 (N_8527,N_7348,N_7493);
or U8528 (N_8528,N_7496,N_7129);
and U8529 (N_8529,N_7962,N_7183);
xnor U8530 (N_8530,N_7841,N_7886);
nor U8531 (N_8531,N_7368,N_7415);
nor U8532 (N_8532,N_7446,N_7867);
nor U8533 (N_8533,N_7965,N_7847);
xor U8534 (N_8534,N_7420,N_7707);
and U8535 (N_8535,N_7266,N_7995);
and U8536 (N_8536,N_7544,N_7215);
or U8537 (N_8537,N_7569,N_7173);
and U8538 (N_8538,N_7245,N_7151);
nand U8539 (N_8539,N_7579,N_7478);
xnor U8540 (N_8540,N_7808,N_7412);
nor U8541 (N_8541,N_7538,N_7384);
xor U8542 (N_8542,N_7741,N_7387);
xor U8543 (N_8543,N_7410,N_7580);
nand U8544 (N_8544,N_7580,N_7232);
and U8545 (N_8545,N_7416,N_7961);
or U8546 (N_8546,N_7945,N_7745);
or U8547 (N_8547,N_7976,N_7283);
or U8548 (N_8548,N_7348,N_7265);
nand U8549 (N_8549,N_7207,N_7900);
nand U8550 (N_8550,N_7938,N_7772);
and U8551 (N_8551,N_7105,N_7558);
nor U8552 (N_8552,N_7224,N_7347);
nor U8553 (N_8553,N_7026,N_7285);
and U8554 (N_8554,N_7697,N_7319);
and U8555 (N_8555,N_7093,N_7936);
and U8556 (N_8556,N_7838,N_7291);
nand U8557 (N_8557,N_7236,N_7536);
or U8558 (N_8558,N_7838,N_7121);
nand U8559 (N_8559,N_7762,N_7391);
and U8560 (N_8560,N_7512,N_7341);
nor U8561 (N_8561,N_7259,N_7306);
nand U8562 (N_8562,N_7838,N_7771);
and U8563 (N_8563,N_7434,N_7039);
nor U8564 (N_8564,N_7942,N_7620);
nor U8565 (N_8565,N_7223,N_7252);
nand U8566 (N_8566,N_7692,N_7320);
xor U8567 (N_8567,N_7755,N_7705);
or U8568 (N_8568,N_7828,N_7925);
nor U8569 (N_8569,N_7749,N_7676);
and U8570 (N_8570,N_7061,N_7384);
nand U8571 (N_8571,N_7890,N_7897);
or U8572 (N_8572,N_7591,N_7899);
nor U8573 (N_8573,N_7048,N_7867);
or U8574 (N_8574,N_7049,N_7512);
nor U8575 (N_8575,N_7630,N_7406);
nor U8576 (N_8576,N_7741,N_7635);
nor U8577 (N_8577,N_7350,N_7255);
or U8578 (N_8578,N_7059,N_7856);
or U8579 (N_8579,N_7046,N_7260);
nor U8580 (N_8580,N_7982,N_7890);
or U8581 (N_8581,N_7684,N_7450);
and U8582 (N_8582,N_7349,N_7313);
nor U8583 (N_8583,N_7237,N_7434);
and U8584 (N_8584,N_7161,N_7685);
nand U8585 (N_8585,N_7983,N_7001);
nor U8586 (N_8586,N_7372,N_7262);
or U8587 (N_8587,N_7231,N_7215);
xnor U8588 (N_8588,N_7939,N_7856);
nor U8589 (N_8589,N_7983,N_7614);
and U8590 (N_8590,N_7989,N_7582);
or U8591 (N_8591,N_7221,N_7524);
nand U8592 (N_8592,N_7613,N_7720);
xor U8593 (N_8593,N_7518,N_7408);
nor U8594 (N_8594,N_7791,N_7437);
nor U8595 (N_8595,N_7682,N_7585);
and U8596 (N_8596,N_7018,N_7165);
nand U8597 (N_8597,N_7476,N_7251);
or U8598 (N_8598,N_7693,N_7124);
xnor U8599 (N_8599,N_7729,N_7420);
nor U8600 (N_8600,N_7336,N_7298);
nand U8601 (N_8601,N_7177,N_7931);
or U8602 (N_8602,N_7648,N_7007);
nand U8603 (N_8603,N_7761,N_7986);
nor U8604 (N_8604,N_7593,N_7280);
nor U8605 (N_8605,N_7195,N_7187);
nand U8606 (N_8606,N_7324,N_7139);
nor U8607 (N_8607,N_7177,N_7953);
or U8608 (N_8608,N_7281,N_7606);
xnor U8609 (N_8609,N_7284,N_7498);
and U8610 (N_8610,N_7504,N_7422);
nand U8611 (N_8611,N_7861,N_7438);
nand U8612 (N_8612,N_7586,N_7983);
nor U8613 (N_8613,N_7109,N_7565);
nor U8614 (N_8614,N_7027,N_7199);
nor U8615 (N_8615,N_7996,N_7054);
nor U8616 (N_8616,N_7572,N_7627);
or U8617 (N_8617,N_7144,N_7061);
nand U8618 (N_8618,N_7753,N_7731);
nor U8619 (N_8619,N_7753,N_7136);
nand U8620 (N_8620,N_7104,N_7038);
and U8621 (N_8621,N_7637,N_7029);
nand U8622 (N_8622,N_7661,N_7362);
and U8623 (N_8623,N_7216,N_7330);
nor U8624 (N_8624,N_7849,N_7183);
or U8625 (N_8625,N_7009,N_7080);
and U8626 (N_8626,N_7747,N_7138);
nand U8627 (N_8627,N_7354,N_7829);
nor U8628 (N_8628,N_7375,N_7697);
xor U8629 (N_8629,N_7724,N_7145);
nor U8630 (N_8630,N_7001,N_7123);
nor U8631 (N_8631,N_7891,N_7339);
or U8632 (N_8632,N_7036,N_7713);
xnor U8633 (N_8633,N_7137,N_7404);
or U8634 (N_8634,N_7231,N_7145);
nand U8635 (N_8635,N_7011,N_7236);
nor U8636 (N_8636,N_7771,N_7184);
nand U8637 (N_8637,N_7478,N_7577);
nand U8638 (N_8638,N_7877,N_7635);
nor U8639 (N_8639,N_7465,N_7863);
nand U8640 (N_8640,N_7927,N_7982);
or U8641 (N_8641,N_7523,N_7303);
nor U8642 (N_8642,N_7901,N_7687);
nor U8643 (N_8643,N_7441,N_7059);
xor U8644 (N_8644,N_7955,N_7314);
nand U8645 (N_8645,N_7539,N_7427);
and U8646 (N_8646,N_7038,N_7545);
nor U8647 (N_8647,N_7675,N_7607);
or U8648 (N_8648,N_7265,N_7542);
and U8649 (N_8649,N_7880,N_7996);
and U8650 (N_8650,N_7562,N_7483);
and U8651 (N_8651,N_7711,N_7373);
or U8652 (N_8652,N_7632,N_7176);
nand U8653 (N_8653,N_7695,N_7673);
and U8654 (N_8654,N_7834,N_7926);
nand U8655 (N_8655,N_7256,N_7804);
nand U8656 (N_8656,N_7214,N_7907);
and U8657 (N_8657,N_7349,N_7923);
or U8658 (N_8658,N_7404,N_7564);
or U8659 (N_8659,N_7293,N_7561);
or U8660 (N_8660,N_7485,N_7331);
nand U8661 (N_8661,N_7498,N_7043);
or U8662 (N_8662,N_7796,N_7052);
and U8663 (N_8663,N_7233,N_7946);
or U8664 (N_8664,N_7718,N_7687);
and U8665 (N_8665,N_7017,N_7904);
nor U8666 (N_8666,N_7711,N_7346);
nor U8667 (N_8667,N_7355,N_7557);
or U8668 (N_8668,N_7021,N_7694);
nand U8669 (N_8669,N_7256,N_7626);
nor U8670 (N_8670,N_7483,N_7969);
nor U8671 (N_8671,N_7194,N_7157);
and U8672 (N_8672,N_7003,N_7211);
or U8673 (N_8673,N_7464,N_7828);
or U8674 (N_8674,N_7780,N_7113);
or U8675 (N_8675,N_7884,N_7279);
nor U8676 (N_8676,N_7513,N_7484);
nor U8677 (N_8677,N_7663,N_7459);
nand U8678 (N_8678,N_7330,N_7733);
or U8679 (N_8679,N_7934,N_7319);
nor U8680 (N_8680,N_7465,N_7856);
nor U8681 (N_8681,N_7855,N_7823);
nor U8682 (N_8682,N_7903,N_7477);
nand U8683 (N_8683,N_7968,N_7479);
xor U8684 (N_8684,N_7753,N_7687);
nand U8685 (N_8685,N_7558,N_7544);
nor U8686 (N_8686,N_7978,N_7817);
nand U8687 (N_8687,N_7937,N_7495);
or U8688 (N_8688,N_7095,N_7355);
nor U8689 (N_8689,N_7565,N_7032);
nand U8690 (N_8690,N_7445,N_7523);
xnor U8691 (N_8691,N_7322,N_7428);
xnor U8692 (N_8692,N_7873,N_7580);
xor U8693 (N_8693,N_7539,N_7954);
nor U8694 (N_8694,N_7307,N_7193);
nand U8695 (N_8695,N_7922,N_7768);
nor U8696 (N_8696,N_7745,N_7725);
or U8697 (N_8697,N_7658,N_7031);
nor U8698 (N_8698,N_7738,N_7322);
nor U8699 (N_8699,N_7836,N_7638);
and U8700 (N_8700,N_7197,N_7338);
xor U8701 (N_8701,N_7758,N_7562);
and U8702 (N_8702,N_7549,N_7520);
and U8703 (N_8703,N_7037,N_7680);
or U8704 (N_8704,N_7312,N_7796);
or U8705 (N_8705,N_7882,N_7795);
nand U8706 (N_8706,N_7018,N_7733);
nand U8707 (N_8707,N_7175,N_7274);
nand U8708 (N_8708,N_7015,N_7329);
nand U8709 (N_8709,N_7003,N_7495);
and U8710 (N_8710,N_7902,N_7822);
xor U8711 (N_8711,N_7173,N_7343);
and U8712 (N_8712,N_7688,N_7691);
nand U8713 (N_8713,N_7147,N_7144);
or U8714 (N_8714,N_7636,N_7584);
nand U8715 (N_8715,N_7650,N_7199);
nand U8716 (N_8716,N_7444,N_7757);
or U8717 (N_8717,N_7155,N_7364);
nor U8718 (N_8718,N_7500,N_7491);
nor U8719 (N_8719,N_7810,N_7749);
nor U8720 (N_8720,N_7089,N_7704);
or U8721 (N_8721,N_7049,N_7386);
nor U8722 (N_8722,N_7039,N_7719);
xor U8723 (N_8723,N_7560,N_7274);
nand U8724 (N_8724,N_7091,N_7049);
xor U8725 (N_8725,N_7751,N_7220);
xor U8726 (N_8726,N_7699,N_7899);
and U8727 (N_8727,N_7311,N_7726);
and U8728 (N_8728,N_7684,N_7706);
nor U8729 (N_8729,N_7693,N_7797);
nand U8730 (N_8730,N_7271,N_7280);
and U8731 (N_8731,N_7566,N_7876);
or U8732 (N_8732,N_7286,N_7946);
and U8733 (N_8733,N_7589,N_7868);
nand U8734 (N_8734,N_7362,N_7858);
nor U8735 (N_8735,N_7812,N_7565);
nor U8736 (N_8736,N_7101,N_7554);
or U8737 (N_8737,N_7111,N_7216);
and U8738 (N_8738,N_7754,N_7038);
nor U8739 (N_8739,N_7725,N_7120);
and U8740 (N_8740,N_7245,N_7208);
nand U8741 (N_8741,N_7996,N_7597);
xnor U8742 (N_8742,N_7680,N_7398);
nand U8743 (N_8743,N_7334,N_7938);
or U8744 (N_8744,N_7629,N_7105);
xnor U8745 (N_8745,N_7938,N_7497);
nor U8746 (N_8746,N_7380,N_7063);
or U8747 (N_8747,N_7875,N_7190);
nor U8748 (N_8748,N_7249,N_7459);
and U8749 (N_8749,N_7445,N_7490);
xor U8750 (N_8750,N_7747,N_7252);
or U8751 (N_8751,N_7222,N_7807);
xnor U8752 (N_8752,N_7543,N_7927);
nor U8753 (N_8753,N_7644,N_7155);
nand U8754 (N_8754,N_7609,N_7979);
xor U8755 (N_8755,N_7735,N_7380);
nand U8756 (N_8756,N_7792,N_7827);
nor U8757 (N_8757,N_7177,N_7324);
or U8758 (N_8758,N_7688,N_7245);
or U8759 (N_8759,N_7506,N_7201);
nand U8760 (N_8760,N_7510,N_7785);
xor U8761 (N_8761,N_7638,N_7526);
nor U8762 (N_8762,N_7206,N_7666);
xnor U8763 (N_8763,N_7880,N_7753);
nor U8764 (N_8764,N_7638,N_7820);
nand U8765 (N_8765,N_7022,N_7617);
or U8766 (N_8766,N_7501,N_7967);
and U8767 (N_8767,N_7002,N_7905);
and U8768 (N_8768,N_7589,N_7718);
nor U8769 (N_8769,N_7706,N_7014);
nor U8770 (N_8770,N_7242,N_7181);
and U8771 (N_8771,N_7539,N_7150);
nand U8772 (N_8772,N_7219,N_7391);
nand U8773 (N_8773,N_7844,N_7598);
nor U8774 (N_8774,N_7287,N_7268);
nand U8775 (N_8775,N_7774,N_7707);
xnor U8776 (N_8776,N_7128,N_7621);
nand U8777 (N_8777,N_7366,N_7064);
or U8778 (N_8778,N_7833,N_7801);
nand U8779 (N_8779,N_7549,N_7971);
nor U8780 (N_8780,N_7282,N_7399);
nand U8781 (N_8781,N_7235,N_7135);
nand U8782 (N_8782,N_7202,N_7816);
nor U8783 (N_8783,N_7271,N_7717);
nand U8784 (N_8784,N_7028,N_7214);
nand U8785 (N_8785,N_7095,N_7720);
nand U8786 (N_8786,N_7910,N_7909);
nor U8787 (N_8787,N_7894,N_7976);
xor U8788 (N_8788,N_7250,N_7379);
nor U8789 (N_8789,N_7720,N_7917);
and U8790 (N_8790,N_7760,N_7010);
nand U8791 (N_8791,N_7169,N_7365);
xnor U8792 (N_8792,N_7666,N_7897);
and U8793 (N_8793,N_7171,N_7407);
or U8794 (N_8794,N_7802,N_7269);
xnor U8795 (N_8795,N_7592,N_7040);
nand U8796 (N_8796,N_7116,N_7549);
nand U8797 (N_8797,N_7206,N_7005);
nand U8798 (N_8798,N_7586,N_7796);
nand U8799 (N_8799,N_7740,N_7639);
nand U8800 (N_8800,N_7305,N_7439);
nand U8801 (N_8801,N_7249,N_7818);
and U8802 (N_8802,N_7837,N_7957);
or U8803 (N_8803,N_7344,N_7873);
nor U8804 (N_8804,N_7690,N_7200);
xor U8805 (N_8805,N_7255,N_7287);
nand U8806 (N_8806,N_7822,N_7737);
nor U8807 (N_8807,N_7735,N_7748);
nand U8808 (N_8808,N_7186,N_7241);
nand U8809 (N_8809,N_7762,N_7733);
and U8810 (N_8810,N_7150,N_7770);
nand U8811 (N_8811,N_7098,N_7635);
or U8812 (N_8812,N_7554,N_7622);
and U8813 (N_8813,N_7149,N_7905);
or U8814 (N_8814,N_7165,N_7107);
xnor U8815 (N_8815,N_7967,N_7421);
nor U8816 (N_8816,N_7617,N_7053);
xor U8817 (N_8817,N_7402,N_7541);
and U8818 (N_8818,N_7926,N_7832);
and U8819 (N_8819,N_7362,N_7908);
nand U8820 (N_8820,N_7157,N_7083);
nor U8821 (N_8821,N_7218,N_7596);
or U8822 (N_8822,N_7151,N_7583);
and U8823 (N_8823,N_7621,N_7012);
nand U8824 (N_8824,N_7457,N_7619);
xor U8825 (N_8825,N_7339,N_7280);
xnor U8826 (N_8826,N_7391,N_7211);
and U8827 (N_8827,N_7050,N_7544);
or U8828 (N_8828,N_7692,N_7634);
nor U8829 (N_8829,N_7362,N_7057);
or U8830 (N_8830,N_7076,N_7238);
nor U8831 (N_8831,N_7242,N_7113);
nor U8832 (N_8832,N_7639,N_7298);
and U8833 (N_8833,N_7185,N_7060);
nand U8834 (N_8834,N_7453,N_7200);
or U8835 (N_8835,N_7070,N_7195);
or U8836 (N_8836,N_7298,N_7491);
xnor U8837 (N_8837,N_7873,N_7736);
or U8838 (N_8838,N_7095,N_7154);
nor U8839 (N_8839,N_7126,N_7662);
and U8840 (N_8840,N_7305,N_7647);
nand U8841 (N_8841,N_7218,N_7999);
or U8842 (N_8842,N_7790,N_7615);
nand U8843 (N_8843,N_7298,N_7396);
nor U8844 (N_8844,N_7647,N_7515);
and U8845 (N_8845,N_7801,N_7701);
nor U8846 (N_8846,N_7823,N_7711);
and U8847 (N_8847,N_7281,N_7150);
and U8848 (N_8848,N_7198,N_7124);
or U8849 (N_8849,N_7550,N_7155);
and U8850 (N_8850,N_7663,N_7612);
nor U8851 (N_8851,N_7762,N_7041);
nand U8852 (N_8852,N_7080,N_7481);
and U8853 (N_8853,N_7161,N_7032);
or U8854 (N_8854,N_7111,N_7632);
nand U8855 (N_8855,N_7219,N_7048);
nand U8856 (N_8856,N_7606,N_7888);
and U8857 (N_8857,N_7133,N_7318);
nand U8858 (N_8858,N_7209,N_7993);
xor U8859 (N_8859,N_7674,N_7056);
or U8860 (N_8860,N_7170,N_7158);
nand U8861 (N_8861,N_7272,N_7352);
and U8862 (N_8862,N_7346,N_7585);
or U8863 (N_8863,N_7293,N_7900);
and U8864 (N_8864,N_7013,N_7799);
nand U8865 (N_8865,N_7943,N_7520);
and U8866 (N_8866,N_7866,N_7874);
nor U8867 (N_8867,N_7275,N_7037);
xnor U8868 (N_8868,N_7934,N_7671);
nor U8869 (N_8869,N_7597,N_7585);
or U8870 (N_8870,N_7144,N_7499);
nand U8871 (N_8871,N_7075,N_7547);
nand U8872 (N_8872,N_7765,N_7607);
nor U8873 (N_8873,N_7019,N_7360);
or U8874 (N_8874,N_7776,N_7371);
nor U8875 (N_8875,N_7386,N_7812);
and U8876 (N_8876,N_7657,N_7323);
and U8877 (N_8877,N_7271,N_7085);
nand U8878 (N_8878,N_7815,N_7665);
nand U8879 (N_8879,N_7465,N_7091);
or U8880 (N_8880,N_7967,N_7066);
and U8881 (N_8881,N_7006,N_7581);
nand U8882 (N_8882,N_7322,N_7264);
or U8883 (N_8883,N_7118,N_7418);
or U8884 (N_8884,N_7366,N_7976);
nor U8885 (N_8885,N_7942,N_7407);
and U8886 (N_8886,N_7542,N_7935);
or U8887 (N_8887,N_7235,N_7054);
nor U8888 (N_8888,N_7211,N_7139);
nor U8889 (N_8889,N_7636,N_7987);
or U8890 (N_8890,N_7187,N_7537);
nand U8891 (N_8891,N_7446,N_7342);
or U8892 (N_8892,N_7656,N_7541);
nor U8893 (N_8893,N_7552,N_7303);
or U8894 (N_8894,N_7155,N_7274);
xnor U8895 (N_8895,N_7661,N_7235);
and U8896 (N_8896,N_7476,N_7283);
xor U8897 (N_8897,N_7715,N_7963);
and U8898 (N_8898,N_7852,N_7690);
nand U8899 (N_8899,N_7314,N_7523);
nor U8900 (N_8900,N_7250,N_7504);
or U8901 (N_8901,N_7955,N_7430);
nand U8902 (N_8902,N_7857,N_7766);
nand U8903 (N_8903,N_7033,N_7914);
xnor U8904 (N_8904,N_7169,N_7870);
or U8905 (N_8905,N_7590,N_7867);
and U8906 (N_8906,N_7236,N_7360);
nor U8907 (N_8907,N_7844,N_7117);
nand U8908 (N_8908,N_7397,N_7530);
and U8909 (N_8909,N_7525,N_7108);
or U8910 (N_8910,N_7861,N_7868);
or U8911 (N_8911,N_7304,N_7488);
nor U8912 (N_8912,N_7854,N_7030);
nand U8913 (N_8913,N_7129,N_7649);
nor U8914 (N_8914,N_7130,N_7945);
and U8915 (N_8915,N_7700,N_7346);
nor U8916 (N_8916,N_7008,N_7356);
nor U8917 (N_8917,N_7732,N_7216);
nand U8918 (N_8918,N_7842,N_7624);
or U8919 (N_8919,N_7026,N_7226);
and U8920 (N_8920,N_7437,N_7921);
or U8921 (N_8921,N_7558,N_7001);
nand U8922 (N_8922,N_7065,N_7509);
nor U8923 (N_8923,N_7413,N_7134);
or U8924 (N_8924,N_7618,N_7874);
or U8925 (N_8925,N_7228,N_7925);
xnor U8926 (N_8926,N_7376,N_7545);
nand U8927 (N_8927,N_7254,N_7891);
nand U8928 (N_8928,N_7215,N_7021);
nand U8929 (N_8929,N_7550,N_7743);
and U8930 (N_8930,N_7935,N_7648);
and U8931 (N_8931,N_7236,N_7902);
nand U8932 (N_8932,N_7253,N_7487);
nor U8933 (N_8933,N_7813,N_7070);
nor U8934 (N_8934,N_7283,N_7497);
xnor U8935 (N_8935,N_7262,N_7031);
nand U8936 (N_8936,N_7640,N_7546);
nand U8937 (N_8937,N_7383,N_7179);
or U8938 (N_8938,N_7048,N_7522);
or U8939 (N_8939,N_7894,N_7134);
or U8940 (N_8940,N_7197,N_7399);
and U8941 (N_8941,N_7369,N_7941);
xnor U8942 (N_8942,N_7544,N_7161);
or U8943 (N_8943,N_7634,N_7596);
nor U8944 (N_8944,N_7123,N_7237);
nand U8945 (N_8945,N_7934,N_7069);
and U8946 (N_8946,N_7988,N_7858);
nor U8947 (N_8947,N_7222,N_7166);
nand U8948 (N_8948,N_7616,N_7618);
nor U8949 (N_8949,N_7917,N_7432);
nand U8950 (N_8950,N_7423,N_7799);
nand U8951 (N_8951,N_7753,N_7056);
and U8952 (N_8952,N_7641,N_7553);
or U8953 (N_8953,N_7913,N_7495);
nor U8954 (N_8954,N_7213,N_7829);
nor U8955 (N_8955,N_7790,N_7407);
xnor U8956 (N_8956,N_7647,N_7395);
nand U8957 (N_8957,N_7849,N_7780);
nand U8958 (N_8958,N_7419,N_7495);
nand U8959 (N_8959,N_7781,N_7580);
or U8960 (N_8960,N_7793,N_7752);
nor U8961 (N_8961,N_7106,N_7158);
nand U8962 (N_8962,N_7589,N_7521);
nor U8963 (N_8963,N_7084,N_7736);
xnor U8964 (N_8964,N_7365,N_7455);
nor U8965 (N_8965,N_7646,N_7467);
nor U8966 (N_8966,N_7388,N_7507);
nor U8967 (N_8967,N_7338,N_7268);
or U8968 (N_8968,N_7665,N_7005);
nor U8969 (N_8969,N_7489,N_7321);
nor U8970 (N_8970,N_7845,N_7349);
nand U8971 (N_8971,N_7083,N_7089);
xor U8972 (N_8972,N_7742,N_7523);
or U8973 (N_8973,N_7297,N_7427);
or U8974 (N_8974,N_7869,N_7944);
nor U8975 (N_8975,N_7162,N_7120);
and U8976 (N_8976,N_7342,N_7327);
nor U8977 (N_8977,N_7021,N_7797);
or U8978 (N_8978,N_7907,N_7586);
nor U8979 (N_8979,N_7601,N_7806);
nor U8980 (N_8980,N_7284,N_7797);
nor U8981 (N_8981,N_7524,N_7460);
and U8982 (N_8982,N_7804,N_7750);
or U8983 (N_8983,N_7880,N_7906);
xnor U8984 (N_8984,N_7273,N_7269);
xnor U8985 (N_8985,N_7684,N_7296);
or U8986 (N_8986,N_7320,N_7294);
nand U8987 (N_8987,N_7285,N_7589);
and U8988 (N_8988,N_7123,N_7527);
nor U8989 (N_8989,N_7335,N_7093);
nor U8990 (N_8990,N_7698,N_7749);
or U8991 (N_8991,N_7345,N_7363);
or U8992 (N_8992,N_7048,N_7202);
nand U8993 (N_8993,N_7048,N_7681);
nor U8994 (N_8994,N_7354,N_7843);
xnor U8995 (N_8995,N_7069,N_7117);
or U8996 (N_8996,N_7052,N_7339);
and U8997 (N_8997,N_7234,N_7231);
nor U8998 (N_8998,N_7488,N_7943);
or U8999 (N_8999,N_7398,N_7810);
and U9000 (N_9000,N_8011,N_8859);
and U9001 (N_9001,N_8389,N_8662);
nand U9002 (N_9002,N_8818,N_8324);
nand U9003 (N_9003,N_8481,N_8686);
and U9004 (N_9004,N_8467,N_8938);
nor U9005 (N_9005,N_8320,N_8739);
nand U9006 (N_9006,N_8709,N_8723);
nand U9007 (N_9007,N_8963,N_8283);
nor U9008 (N_9008,N_8910,N_8230);
and U9009 (N_9009,N_8304,N_8051);
or U9010 (N_9010,N_8242,N_8484);
xnor U9011 (N_9011,N_8544,N_8599);
or U9012 (N_9012,N_8770,N_8347);
or U9013 (N_9013,N_8502,N_8372);
nand U9014 (N_9014,N_8329,N_8319);
or U9015 (N_9015,N_8003,N_8955);
or U9016 (N_9016,N_8618,N_8937);
xor U9017 (N_9017,N_8174,N_8430);
or U9018 (N_9018,N_8468,N_8398);
and U9019 (N_9019,N_8703,N_8844);
nand U9020 (N_9020,N_8078,N_8228);
xnor U9021 (N_9021,N_8914,N_8908);
nor U9022 (N_9022,N_8298,N_8753);
and U9023 (N_9023,N_8515,N_8269);
or U9024 (N_9024,N_8335,N_8868);
and U9025 (N_9025,N_8388,N_8953);
nand U9026 (N_9026,N_8040,N_8750);
or U9027 (N_9027,N_8704,N_8001);
and U9028 (N_9028,N_8728,N_8352);
and U9029 (N_9029,N_8710,N_8161);
nor U9030 (N_9030,N_8475,N_8521);
or U9031 (N_9031,N_8623,N_8035);
and U9032 (N_9032,N_8375,N_8511);
or U9033 (N_9033,N_8848,N_8672);
or U9034 (N_9034,N_8429,N_8217);
nand U9035 (N_9035,N_8474,N_8852);
xor U9036 (N_9036,N_8842,N_8622);
and U9037 (N_9037,N_8558,N_8266);
xnor U9038 (N_9038,N_8743,N_8680);
and U9039 (N_9039,N_8940,N_8000);
nor U9040 (N_9040,N_8446,N_8719);
xnor U9041 (N_9041,N_8082,N_8810);
or U9042 (N_9042,N_8769,N_8655);
or U9043 (N_9043,N_8529,N_8567);
or U9044 (N_9044,N_8221,N_8459);
and U9045 (N_9045,N_8886,N_8768);
nor U9046 (N_9046,N_8187,N_8302);
and U9047 (N_9047,N_8562,N_8516);
and U9048 (N_9048,N_8006,N_8321);
or U9049 (N_9049,N_8986,N_8184);
nor U9050 (N_9050,N_8913,N_8280);
or U9051 (N_9051,N_8873,N_8155);
or U9052 (N_9052,N_8846,N_8311);
nor U9053 (N_9053,N_8210,N_8564);
nor U9054 (N_9054,N_8636,N_8486);
and U9055 (N_9055,N_8954,N_8919);
xor U9056 (N_9056,N_8890,N_8050);
nor U9057 (N_9057,N_8104,N_8584);
nand U9058 (N_9058,N_8610,N_8393);
nand U9059 (N_9059,N_8142,N_8421);
nor U9060 (N_9060,N_8075,N_8668);
xnor U9061 (N_9061,N_8885,N_8355);
nor U9062 (N_9062,N_8721,N_8215);
or U9063 (N_9063,N_8649,N_8927);
nand U9064 (N_9064,N_8359,N_8935);
and U9065 (N_9065,N_8858,N_8904);
or U9066 (N_9066,N_8626,N_8160);
and U9067 (N_9067,N_8219,N_8088);
nand U9068 (N_9068,N_8089,N_8026);
nand U9069 (N_9069,N_8439,N_8235);
and U9070 (N_9070,N_8748,N_8362);
nor U9071 (N_9071,N_8381,N_8385);
and U9072 (N_9072,N_8682,N_8870);
or U9073 (N_9073,N_8609,N_8119);
or U9074 (N_9074,N_8985,N_8896);
nand U9075 (N_9075,N_8592,N_8106);
nor U9076 (N_9076,N_8772,N_8336);
nand U9077 (N_9077,N_8891,N_8037);
and U9078 (N_9078,N_8419,N_8978);
or U9079 (N_9079,N_8277,N_8493);
nor U9080 (N_9080,N_8416,N_8379);
xnor U9081 (N_9081,N_8476,N_8532);
nand U9082 (N_9082,N_8305,N_8783);
and U9083 (N_9083,N_8248,N_8345);
and U9084 (N_9084,N_8926,N_8237);
nor U9085 (N_9085,N_8295,N_8265);
or U9086 (N_9086,N_8877,N_8044);
nand U9087 (N_9087,N_8363,N_8767);
nor U9088 (N_9088,N_8547,N_8201);
nor U9089 (N_9089,N_8572,N_8069);
nor U9090 (N_9090,N_8025,N_8561);
or U9091 (N_9091,N_8101,N_8096);
or U9092 (N_9092,N_8100,N_8471);
or U9093 (N_9093,N_8951,N_8137);
nor U9094 (N_9094,N_8495,N_8538);
nor U9095 (N_9095,N_8800,N_8700);
and U9096 (N_9096,N_8679,N_8008);
nor U9097 (N_9097,N_8675,N_8845);
xor U9098 (N_9098,N_8880,N_8310);
nand U9099 (N_9099,N_8537,N_8929);
nand U9100 (N_9100,N_8799,N_8976);
or U9101 (N_9101,N_8965,N_8642);
or U9102 (N_9102,N_8226,N_8167);
nand U9103 (N_9103,N_8340,N_8997);
nand U9104 (N_9104,N_8604,N_8922);
or U9105 (N_9105,N_8854,N_8548);
or U9106 (N_9106,N_8202,N_8047);
nor U9107 (N_9107,N_8261,N_8673);
nand U9108 (N_9108,N_8331,N_8071);
nand U9109 (N_9109,N_8941,N_8199);
xor U9110 (N_9110,N_8090,N_8024);
xnor U9111 (N_9111,N_8092,N_8969);
nand U9112 (N_9112,N_8658,N_8125);
and U9113 (N_9113,N_8826,N_8166);
nor U9114 (N_9114,N_8346,N_8002);
or U9115 (N_9115,N_8897,N_8150);
nand U9116 (N_9116,N_8272,N_8395);
and U9117 (N_9117,N_8365,N_8020);
nor U9118 (N_9118,N_8061,N_8653);
nand U9119 (N_9119,N_8693,N_8225);
nand U9120 (N_9120,N_8654,N_8023);
xnor U9121 (N_9121,N_8569,N_8522);
and U9122 (N_9122,N_8670,N_8640);
and U9123 (N_9123,N_8987,N_8815);
or U9124 (N_9124,N_8696,N_8671);
and U9125 (N_9125,N_8557,N_8190);
and U9126 (N_9126,N_8134,N_8862);
nor U9127 (N_9127,N_8478,N_8426);
and U9128 (N_9128,N_8909,N_8053);
and U9129 (N_9129,N_8308,N_8126);
or U9130 (N_9130,N_8593,N_8041);
or U9131 (N_9131,N_8282,N_8921);
nand U9132 (N_9132,N_8930,N_8959);
and U9133 (N_9133,N_8369,N_8268);
nand U9134 (N_9134,N_8177,N_8578);
xnor U9135 (N_9135,N_8761,N_8249);
or U9136 (N_9136,N_8832,N_8875);
nor U9137 (N_9137,N_8813,N_8549);
nor U9138 (N_9138,N_8725,N_8583);
nor U9139 (N_9139,N_8232,N_8692);
nand U9140 (N_9140,N_8286,N_8573);
nand U9141 (N_9141,N_8776,N_8924);
and U9142 (N_9142,N_8131,N_8747);
nand U9143 (N_9143,N_8338,N_8974);
and U9144 (N_9144,N_8962,N_8669);
and U9145 (N_9145,N_8513,N_8588);
or U9146 (N_9146,N_8605,N_8076);
or U9147 (N_9147,N_8775,N_8932);
or U9148 (N_9148,N_8118,N_8254);
and U9149 (N_9149,N_8496,N_8713);
or U9150 (N_9150,N_8469,N_8330);
xor U9151 (N_9151,N_8087,N_8864);
nor U9152 (N_9152,N_8386,N_8146);
or U9153 (N_9153,N_8780,N_8115);
nor U9154 (N_9154,N_8508,N_8638);
xor U9155 (N_9155,N_8796,N_8505);
nor U9156 (N_9156,N_8449,N_8110);
and U9157 (N_9157,N_8808,N_8151);
and U9158 (N_9158,N_8480,N_8099);
or U9159 (N_9159,N_8968,N_8742);
and U9160 (N_9160,N_8267,N_8530);
or U9161 (N_9161,N_8033,N_8807);
xnor U9162 (N_9162,N_8227,N_8466);
and U9163 (N_9163,N_8400,N_8758);
xnor U9164 (N_9164,N_8433,N_8760);
nor U9165 (N_9165,N_8519,N_8062);
xnor U9166 (N_9166,N_8643,N_8863);
and U9167 (N_9167,N_8869,N_8133);
and U9168 (N_9168,N_8804,N_8209);
nor U9169 (N_9169,N_8039,N_8361);
and U9170 (N_9170,N_8180,N_8339);
or U9171 (N_9171,N_8902,N_8181);
nand U9172 (N_9172,N_8980,N_8022);
or U9173 (N_9173,N_8911,N_8958);
and U9174 (N_9174,N_8895,N_8198);
and U9175 (N_9175,N_8540,N_8881);
xnor U9176 (N_9176,N_8835,N_8491);
nor U9177 (N_9177,N_8646,N_8535);
and U9178 (N_9178,N_8317,N_8438);
or U9179 (N_9179,N_8787,N_8171);
or U9180 (N_9180,N_8417,N_8034);
or U9181 (N_9181,N_8425,N_8794);
nand U9182 (N_9182,N_8314,N_8829);
nor U9183 (N_9183,N_8326,N_8690);
and U9184 (N_9184,N_8664,N_8531);
and U9185 (N_9185,N_8387,N_8706);
or U9186 (N_9186,N_8916,N_8801);
and U9187 (N_9187,N_8652,N_8773);
xnor U9188 (N_9188,N_8485,N_8410);
nand U9189 (N_9189,N_8162,N_8506);
nand U9190 (N_9190,N_8114,N_8831);
or U9191 (N_9191,N_8503,N_8418);
nor U9192 (N_9192,N_8836,N_8175);
xor U9193 (N_9193,N_8934,N_8458);
nor U9194 (N_9194,N_8793,N_8716);
or U9195 (N_9195,N_8325,N_8192);
nand U9196 (N_9196,N_8143,N_8526);
and U9197 (N_9197,N_8729,N_8094);
or U9198 (N_9198,N_8018,N_8737);
nor U9199 (N_9199,N_8887,N_8463);
nand U9200 (N_9200,N_8312,N_8250);
and U9201 (N_9201,N_8782,N_8809);
nand U9202 (N_9202,N_8553,N_8205);
nand U9203 (N_9203,N_8698,N_8377);
nor U9204 (N_9204,N_8197,N_8855);
and U9205 (N_9205,N_8098,N_8689);
and U9206 (N_9206,N_8193,N_8477);
or U9207 (N_9207,N_8371,N_8580);
or U9208 (N_9208,N_8045,N_8453);
nand U9209 (N_9209,N_8762,N_8194);
nand U9210 (N_9210,N_8163,N_8582);
nand U9211 (N_9211,N_8255,N_8333);
nor U9212 (N_9212,N_8273,N_8617);
nor U9213 (N_9213,N_8517,N_8647);
or U9214 (N_9214,N_8139,N_8661);
nor U9215 (N_9215,N_8074,N_8472);
nand U9216 (N_9216,N_8204,N_8399);
nand U9217 (N_9217,N_8473,N_8883);
nand U9218 (N_9218,N_8173,N_8032);
xnor U9219 (N_9219,N_8394,N_8296);
or U9220 (N_9220,N_8214,N_8176);
or U9221 (N_9221,N_8406,N_8754);
nand U9222 (N_9222,N_8520,N_8523);
nor U9223 (N_9223,N_8281,N_8252);
xor U9224 (N_9224,N_8946,N_8920);
nand U9225 (N_9225,N_8405,N_8524);
nor U9226 (N_9226,N_8591,N_8939);
and U9227 (N_9227,N_8085,N_8639);
nor U9228 (N_9228,N_8504,N_8067);
xnor U9229 (N_9229,N_8510,N_8917);
or U9230 (N_9230,N_8309,N_8634);
or U9231 (N_9231,N_8574,N_8964);
and U9232 (N_9232,N_8840,N_8595);
nand U9233 (N_9233,N_8103,N_8853);
nor U9234 (N_9234,N_8158,N_8996);
and U9235 (N_9235,N_8683,N_8132);
nand U9236 (N_9236,N_8494,N_8749);
nor U9237 (N_9237,N_8284,N_8925);
nor U9238 (N_9238,N_8814,N_8373);
and U9239 (N_9239,N_8983,N_8489);
and U9240 (N_9240,N_8454,N_8822);
nor U9241 (N_9241,N_8536,N_8534);
nand U9242 (N_9242,N_8243,N_8995);
and U9243 (N_9243,N_8083,N_8397);
nor U9244 (N_9244,N_8961,N_8650);
xor U9245 (N_9245,N_8148,N_8641);
nand U9246 (N_9246,N_8744,N_8354);
nand U9247 (N_9247,N_8712,N_8726);
nand U9248 (N_9248,N_8200,N_8428);
or U9249 (N_9249,N_8292,N_8931);
and U9250 (N_9250,N_8060,N_8460);
nor U9251 (N_9251,N_8152,N_8701);
or U9252 (N_9252,N_8518,N_8630);
or U9253 (N_9253,N_8789,N_8492);
nand U9254 (N_9254,N_8483,N_8031);
or U9255 (N_9255,N_8656,N_8404);
and U9256 (N_9256,N_8236,N_8420);
xor U9257 (N_9257,N_8186,N_8833);
nor U9258 (N_9258,N_8203,N_8563);
and U9259 (N_9259,N_8279,N_8994);
and U9260 (N_9260,N_8967,N_8358);
and U9261 (N_9261,N_8154,N_8241);
and U9262 (N_9262,N_8752,N_8797);
or U9263 (N_9263,N_8102,N_8111);
nand U9264 (N_9264,N_8733,N_8621);
and U9265 (N_9265,N_8790,N_8966);
xor U9266 (N_9266,N_8651,N_8447);
xor U9267 (N_9267,N_8356,N_8565);
nand U9268 (N_9268,N_8688,N_8571);
and U9269 (N_9269,N_8570,N_8830);
nand U9270 (N_9270,N_8707,N_8351);
or U9271 (N_9271,N_8608,N_8612);
or U9272 (N_9272,N_8512,N_8253);
and U9273 (N_9273,N_8258,N_8063);
nand U9274 (N_9274,N_8973,N_8942);
nand U9275 (N_9275,N_8556,N_8015);
nor U9276 (N_9276,N_8322,N_8884);
nor U9277 (N_9277,N_8287,N_8348);
nor U9278 (N_9278,N_8834,N_8380);
or U9279 (N_9279,N_8587,N_8819);
and U9280 (N_9280,N_8285,N_8016);
nor U9281 (N_9281,N_8216,N_8042);
nor U9282 (N_9282,N_8189,N_8527);
nand U9283 (N_9283,N_8212,N_8576);
nand U9284 (N_9284,N_8828,N_8817);
nor U9285 (N_9285,N_8977,N_8313);
and U9286 (N_9286,N_8350,N_8368);
nand U9287 (N_9287,N_8756,N_8208);
or U9288 (N_9288,N_8005,N_8989);
and U9289 (N_9289,N_8635,N_8093);
nor U9290 (N_9290,N_8038,N_8971);
nand U9291 (N_9291,N_8164,N_8271);
or U9292 (N_9292,N_8383,N_8297);
nor U9293 (N_9293,N_8147,N_8220);
nand U9294 (N_9294,N_8718,N_8191);
and U9295 (N_9295,N_8247,N_8620);
nand U9296 (N_9296,N_8603,N_8676);
or U9297 (N_9297,N_8207,N_8849);
or U9298 (N_9298,N_8708,N_8695);
or U9299 (N_9299,N_8434,N_8879);
or U9300 (N_9300,N_8856,N_8455);
nand U9301 (N_9301,N_8301,N_8169);
nor U9302 (N_9302,N_8123,N_8751);
nand U9303 (N_9303,N_8012,N_8509);
or U9304 (N_9304,N_8555,N_8949);
or U9305 (N_9305,N_8999,N_8898);
or U9306 (N_9306,N_8256,N_8805);
nor U9307 (N_9307,N_8627,N_8239);
and U9308 (N_9308,N_8763,N_8857);
nand U9309 (N_9309,N_8979,N_8874);
or U9310 (N_9310,N_8841,N_8928);
or U9311 (N_9311,N_8488,N_8278);
and U9312 (N_9312,N_8262,N_8129);
nand U9313 (N_9313,N_8436,N_8888);
nand U9314 (N_9314,N_8081,N_8121);
nand U9315 (N_9315,N_8059,N_8543);
nand U9316 (N_9316,N_8140,N_8407);
nor U9317 (N_9317,N_8990,N_8843);
or U9318 (N_9318,N_8264,N_8795);
or U9319 (N_9319,N_8936,N_8982);
and U9320 (N_9320,N_8188,N_8528);
nand U9321 (N_9321,N_8316,N_8464);
nor U9322 (N_9322,N_8364,N_8714);
and U9323 (N_9323,N_8401,N_8112);
nand U9324 (N_9324,N_8777,N_8745);
or U9325 (N_9325,N_8440,N_8616);
nor U9326 (N_9326,N_8409,N_8900);
nor U9327 (N_9327,N_8457,N_8798);
and U9328 (N_9328,N_8396,N_8731);
xnor U9329 (N_9329,N_8514,N_8392);
and U9330 (N_9330,N_8288,N_8274);
xnor U9331 (N_9331,N_8168,N_8550);
or U9332 (N_9332,N_8452,N_8443);
nand U9333 (N_9333,N_8165,N_8705);
and U9334 (N_9334,N_8947,N_8499);
and U9335 (N_9335,N_8108,N_8577);
or U9336 (N_9336,N_8678,N_8657);
xnor U9337 (N_9337,N_8086,N_8736);
and U9338 (N_9338,N_8299,N_8231);
nand U9339 (N_9339,N_8195,N_8027);
and U9340 (N_9340,N_8575,N_8233);
and U9341 (N_9341,N_8507,N_8560);
nand U9342 (N_9342,N_8130,N_8244);
nor U9343 (N_9343,N_8357,N_8812);
nand U9344 (N_9344,N_8013,N_8975);
and U9345 (N_9345,N_8402,N_8960);
nor U9346 (N_9346,N_8988,N_8213);
nor U9347 (N_9347,N_8554,N_8991);
and U9348 (N_9348,N_8732,N_8117);
nand U9349 (N_9349,N_8431,N_8702);
and U9350 (N_9350,N_8791,N_8172);
nand U9351 (N_9351,N_8289,N_8501);
nand U9352 (N_9352,N_8290,N_8923);
nor U9353 (N_9353,N_8145,N_8028);
and U9354 (N_9354,N_8327,N_8633);
and U9355 (N_9355,N_8907,N_8590);
nor U9356 (N_9356,N_8120,N_8972);
or U9357 (N_9357,N_8334,N_8614);
and U9358 (N_9358,N_8811,N_8624);
nand U9359 (N_9359,N_8912,N_8533);
nand U9360 (N_9360,N_8918,N_8344);
and U9361 (N_9361,N_8066,N_8224);
nor U9362 (N_9362,N_8802,N_8435);
and U9363 (N_9363,N_8784,N_8222);
xor U9364 (N_9364,N_8437,N_8771);
or U9365 (N_9365,N_8602,N_8043);
or U9366 (N_9366,N_8091,N_8957);
and U9367 (N_9367,N_8867,N_8337);
or U9368 (N_9368,N_8122,N_8984);
nor U9369 (N_9369,N_8470,N_8291);
or U9370 (N_9370,N_8838,N_8981);
and U9371 (N_9371,N_8303,N_8036);
or U9372 (N_9372,N_8792,N_8185);
nor U9373 (N_9373,N_8645,N_8766);
nor U9374 (N_9374,N_8779,N_8077);
and U9375 (N_9375,N_8611,N_8052);
and U9376 (N_9376,N_8153,N_8684);
or U9377 (N_9377,N_8084,N_8539);
or U9378 (N_9378,N_8422,N_8411);
nor U9379 (N_9379,N_8442,N_8097);
nor U9380 (N_9380,N_8229,N_8915);
or U9381 (N_9381,N_8821,N_8542);
nand U9382 (N_9382,N_8004,N_8579);
nand U9383 (N_9383,N_8566,N_8223);
and U9384 (N_9384,N_8666,N_8992);
xnor U9385 (N_9385,N_8781,N_8765);
and U9386 (N_9386,N_8674,N_8029);
xnor U9387 (N_9387,N_8159,N_8057);
or U9388 (N_9388,N_8601,N_8851);
or U9389 (N_9389,N_8054,N_8816);
and U9390 (N_9390,N_8376,N_8600);
nand U9391 (N_9391,N_8183,N_8391);
xnor U9392 (N_9392,N_8774,N_8541);
nand U9393 (N_9393,N_8720,N_8559);
nand U9394 (N_9394,N_8245,N_8157);
nand U9395 (N_9395,N_8615,N_8257);
nor U9396 (N_9396,N_8586,N_8839);
nand U9397 (N_9397,N_8384,N_8487);
nor U9398 (N_9398,N_8741,N_8070);
and U9399 (N_9399,N_8196,N_8901);
nand U9400 (N_9400,N_8850,N_8056);
nor U9401 (N_9401,N_8307,N_8755);
nor U9402 (N_9402,N_8724,N_8894);
or U9403 (N_9403,N_8500,N_8049);
xor U9404 (N_9404,N_8251,N_8105);
nand U9405 (N_9405,N_8892,N_8080);
nor U9406 (N_9406,N_8759,N_8068);
nor U9407 (N_9407,N_8631,N_8677);
nand U9408 (N_9408,N_8367,N_8525);
xor U9409 (N_9409,N_8594,N_8149);
and U9410 (N_9410,N_8107,N_8246);
nand U9411 (N_9411,N_8551,N_8156);
and U9412 (N_9412,N_8497,N_8903);
and U9413 (N_9413,N_8135,N_8598);
and U9414 (N_9414,N_8697,N_8432);
and U9415 (N_9415,N_8803,N_8374);
nand U9416 (N_9416,N_8717,N_8889);
xnor U9417 (N_9417,N_8342,N_8625);
and U9418 (N_9418,N_8872,N_8825);
nand U9419 (N_9419,N_8568,N_8451);
nor U9420 (N_9420,N_8055,N_8427);
and U9421 (N_9421,N_8546,N_8127);
nor U9422 (N_9422,N_8370,N_8735);
nor U9423 (N_9423,N_8685,N_8138);
and U9424 (N_9424,N_8727,N_8993);
xor U9425 (N_9425,N_8589,N_8619);
nor U9426 (N_9426,N_8667,N_8847);
nor U9427 (N_9427,N_8058,N_8360);
nand U9428 (N_9428,N_8017,N_8412);
and U9429 (N_9429,N_8699,N_8906);
nand U9430 (N_9430,N_8585,N_8628);
xnor U9431 (N_9431,N_8009,N_8182);
xnor U9432 (N_9432,N_8490,N_8141);
nand U9433 (N_9433,N_8461,N_8136);
and U9434 (N_9434,N_8046,N_8240);
or U9435 (N_9435,N_8206,N_8823);
nand U9436 (N_9436,N_8933,N_8456);
nor U9437 (N_9437,N_8637,N_8450);
and U9438 (N_9438,N_8413,N_8865);
and U9439 (N_9439,N_8238,N_8415);
or U9440 (N_9440,N_8970,N_8332);
nor U9441 (N_9441,N_8144,N_8366);
and U9442 (N_9442,N_8956,N_8871);
nand U9443 (N_9443,N_8820,N_8079);
or U9444 (N_9444,N_8660,N_8806);
or U9445 (N_9445,N_8876,N_8293);
nor U9446 (N_9446,N_8275,N_8234);
or U9447 (N_9447,N_8014,N_8270);
and U9448 (N_9448,N_8306,N_8545);
nor U9449 (N_9449,N_8764,N_8691);
and U9450 (N_9450,N_8659,N_8952);
nor U9451 (N_9451,N_8482,N_8294);
xor U9452 (N_9452,N_8738,N_8866);
and U9453 (N_9453,N_8109,N_8178);
and U9454 (N_9454,N_8613,N_8943);
or U9455 (N_9455,N_8893,N_8606);
nor U9456 (N_9456,N_8378,N_8341);
or U9457 (N_9457,N_8581,N_8423);
nor U9458 (N_9458,N_8552,N_8179);
or U9459 (N_9459,N_8073,N_8128);
and U9460 (N_9460,N_8632,N_8607);
or U9461 (N_9461,N_8064,N_8837);
nor U9462 (N_9462,N_8785,N_8328);
nor U9463 (N_9463,N_8259,N_8382);
nand U9464 (N_9464,N_8072,N_8681);
nor U9465 (N_9465,N_8629,N_8408);
or U9466 (N_9466,N_8030,N_8878);
nor U9467 (N_9467,N_8065,N_8444);
nor U9468 (N_9468,N_8882,N_8711);
nor U9469 (N_9469,N_8263,N_8300);
nand U9470 (N_9470,N_8860,N_8462);
or U9471 (N_9471,N_8124,N_8390);
and U9472 (N_9472,N_8663,N_8276);
and U9473 (N_9473,N_8343,N_8424);
nor U9474 (N_9474,N_8441,N_8757);
and U9475 (N_9475,N_8746,N_8445);
and U9476 (N_9476,N_8403,N_8414);
nor U9477 (N_9477,N_8944,N_8824);
nor U9478 (N_9478,N_8113,N_8665);
nand U9479 (N_9479,N_8095,N_8715);
nor U9480 (N_9480,N_8007,N_8644);
nand U9481 (N_9481,N_8722,N_8734);
nand U9482 (N_9482,N_8465,N_8448);
and U9483 (N_9483,N_8899,N_8948);
nand U9484 (N_9484,N_8786,N_8170);
and U9485 (N_9485,N_8498,N_8479);
nand U9486 (N_9486,N_8694,N_8687);
nor U9487 (N_9487,N_8218,N_8827);
nand U9488 (N_9488,N_8596,N_8740);
or U9489 (N_9489,N_8730,N_8905);
xor U9490 (N_9490,N_8788,N_8648);
nor U9491 (N_9491,N_8998,N_8778);
and U9492 (N_9492,N_8021,N_8048);
xor U9493 (N_9493,N_8211,N_8353);
nand U9494 (N_9494,N_8861,N_8950);
nor U9495 (N_9495,N_8010,N_8260);
nand U9496 (N_9496,N_8945,N_8019);
nor U9497 (N_9497,N_8349,N_8318);
nor U9498 (N_9498,N_8315,N_8116);
or U9499 (N_9499,N_8323,N_8597);
nand U9500 (N_9500,N_8897,N_8985);
nor U9501 (N_9501,N_8527,N_8178);
nor U9502 (N_9502,N_8445,N_8429);
and U9503 (N_9503,N_8584,N_8393);
nor U9504 (N_9504,N_8767,N_8987);
nor U9505 (N_9505,N_8209,N_8034);
nand U9506 (N_9506,N_8626,N_8232);
and U9507 (N_9507,N_8752,N_8696);
and U9508 (N_9508,N_8086,N_8815);
xor U9509 (N_9509,N_8038,N_8582);
or U9510 (N_9510,N_8014,N_8614);
nor U9511 (N_9511,N_8101,N_8183);
and U9512 (N_9512,N_8499,N_8636);
or U9513 (N_9513,N_8786,N_8611);
and U9514 (N_9514,N_8606,N_8437);
and U9515 (N_9515,N_8080,N_8188);
or U9516 (N_9516,N_8895,N_8111);
and U9517 (N_9517,N_8686,N_8897);
nand U9518 (N_9518,N_8602,N_8425);
and U9519 (N_9519,N_8123,N_8174);
nor U9520 (N_9520,N_8129,N_8351);
nor U9521 (N_9521,N_8111,N_8268);
nand U9522 (N_9522,N_8426,N_8095);
nand U9523 (N_9523,N_8206,N_8545);
nor U9524 (N_9524,N_8189,N_8481);
or U9525 (N_9525,N_8930,N_8908);
nand U9526 (N_9526,N_8726,N_8156);
nand U9527 (N_9527,N_8194,N_8737);
or U9528 (N_9528,N_8960,N_8704);
nor U9529 (N_9529,N_8663,N_8316);
and U9530 (N_9530,N_8443,N_8602);
and U9531 (N_9531,N_8590,N_8135);
nor U9532 (N_9532,N_8059,N_8855);
or U9533 (N_9533,N_8518,N_8345);
xor U9534 (N_9534,N_8055,N_8181);
nor U9535 (N_9535,N_8884,N_8589);
or U9536 (N_9536,N_8785,N_8530);
or U9537 (N_9537,N_8013,N_8619);
nand U9538 (N_9538,N_8969,N_8197);
or U9539 (N_9539,N_8703,N_8327);
or U9540 (N_9540,N_8002,N_8579);
nor U9541 (N_9541,N_8089,N_8972);
xnor U9542 (N_9542,N_8181,N_8218);
and U9543 (N_9543,N_8167,N_8248);
nand U9544 (N_9544,N_8395,N_8227);
or U9545 (N_9545,N_8137,N_8388);
xnor U9546 (N_9546,N_8992,N_8092);
nor U9547 (N_9547,N_8419,N_8251);
or U9548 (N_9548,N_8056,N_8184);
nand U9549 (N_9549,N_8188,N_8543);
nand U9550 (N_9550,N_8454,N_8947);
or U9551 (N_9551,N_8151,N_8658);
and U9552 (N_9552,N_8941,N_8620);
nor U9553 (N_9553,N_8201,N_8988);
nor U9554 (N_9554,N_8492,N_8029);
and U9555 (N_9555,N_8757,N_8761);
and U9556 (N_9556,N_8958,N_8909);
nor U9557 (N_9557,N_8778,N_8624);
nand U9558 (N_9558,N_8379,N_8613);
or U9559 (N_9559,N_8563,N_8753);
nand U9560 (N_9560,N_8733,N_8368);
nand U9561 (N_9561,N_8247,N_8830);
and U9562 (N_9562,N_8222,N_8101);
nor U9563 (N_9563,N_8039,N_8980);
nand U9564 (N_9564,N_8016,N_8597);
or U9565 (N_9565,N_8696,N_8703);
or U9566 (N_9566,N_8845,N_8293);
and U9567 (N_9567,N_8713,N_8447);
and U9568 (N_9568,N_8086,N_8909);
xnor U9569 (N_9569,N_8355,N_8445);
nor U9570 (N_9570,N_8963,N_8749);
nand U9571 (N_9571,N_8898,N_8677);
nor U9572 (N_9572,N_8415,N_8266);
nand U9573 (N_9573,N_8929,N_8556);
and U9574 (N_9574,N_8194,N_8078);
or U9575 (N_9575,N_8808,N_8471);
and U9576 (N_9576,N_8691,N_8283);
and U9577 (N_9577,N_8494,N_8530);
or U9578 (N_9578,N_8246,N_8854);
xnor U9579 (N_9579,N_8195,N_8429);
or U9580 (N_9580,N_8451,N_8115);
xnor U9581 (N_9581,N_8960,N_8000);
nor U9582 (N_9582,N_8251,N_8106);
nand U9583 (N_9583,N_8922,N_8981);
nor U9584 (N_9584,N_8636,N_8150);
nor U9585 (N_9585,N_8902,N_8059);
nand U9586 (N_9586,N_8590,N_8442);
xor U9587 (N_9587,N_8788,N_8726);
or U9588 (N_9588,N_8673,N_8823);
and U9589 (N_9589,N_8254,N_8278);
nor U9590 (N_9590,N_8157,N_8877);
nor U9591 (N_9591,N_8786,N_8788);
xnor U9592 (N_9592,N_8113,N_8508);
and U9593 (N_9593,N_8776,N_8085);
or U9594 (N_9594,N_8751,N_8325);
or U9595 (N_9595,N_8647,N_8165);
and U9596 (N_9596,N_8568,N_8316);
or U9597 (N_9597,N_8578,N_8843);
and U9598 (N_9598,N_8333,N_8410);
and U9599 (N_9599,N_8182,N_8978);
and U9600 (N_9600,N_8916,N_8596);
nor U9601 (N_9601,N_8040,N_8688);
nor U9602 (N_9602,N_8401,N_8615);
or U9603 (N_9603,N_8303,N_8617);
nor U9604 (N_9604,N_8015,N_8407);
nor U9605 (N_9605,N_8351,N_8451);
or U9606 (N_9606,N_8353,N_8157);
or U9607 (N_9607,N_8344,N_8175);
nor U9608 (N_9608,N_8164,N_8155);
and U9609 (N_9609,N_8052,N_8029);
nor U9610 (N_9610,N_8619,N_8428);
nor U9611 (N_9611,N_8557,N_8431);
and U9612 (N_9612,N_8082,N_8289);
and U9613 (N_9613,N_8114,N_8748);
nor U9614 (N_9614,N_8403,N_8375);
xnor U9615 (N_9615,N_8737,N_8831);
or U9616 (N_9616,N_8364,N_8578);
or U9617 (N_9617,N_8559,N_8761);
nor U9618 (N_9618,N_8504,N_8190);
or U9619 (N_9619,N_8072,N_8706);
nor U9620 (N_9620,N_8717,N_8745);
xor U9621 (N_9621,N_8516,N_8960);
xor U9622 (N_9622,N_8191,N_8804);
or U9623 (N_9623,N_8237,N_8281);
and U9624 (N_9624,N_8022,N_8458);
nor U9625 (N_9625,N_8594,N_8556);
xnor U9626 (N_9626,N_8811,N_8261);
nor U9627 (N_9627,N_8871,N_8286);
xor U9628 (N_9628,N_8661,N_8282);
and U9629 (N_9629,N_8473,N_8727);
xor U9630 (N_9630,N_8716,N_8680);
nand U9631 (N_9631,N_8376,N_8285);
nor U9632 (N_9632,N_8759,N_8310);
xnor U9633 (N_9633,N_8897,N_8002);
nand U9634 (N_9634,N_8148,N_8543);
nand U9635 (N_9635,N_8880,N_8411);
and U9636 (N_9636,N_8565,N_8782);
and U9637 (N_9637,N_8127,N_8688);
and U9638 (N_9638,N_8485,N_8858);
and U9639 (N_9639,N_8463,N_8836);
nand U9640 (N_9640,N_8985,N_8720);
or U9641 (N_9641,N_8654,N_8831);
xor U9642 (N_9642,N_8203,N_8689);
and U9643 (N_9643,N_8262,N_8955);
nor U9644 (N_9644,N_8035,N_8973);
and U9645 (N_9645,N_8540,N_8019);
nand U9646 (N_9646,N_8037,N_8763);
xnor U9647 (N_9647,N_8269,N_8852);
and U9648 (N_9648,N_8538,N_8911);
xor U9649 (N_9649,N_8470,N_8301);
and U9650 (N_9650,N_8902,N_8912);
or U9651 (N_9651,N_8811,N_8843);
nand U9652 (N_9652,N_8048,N_8764);
or U9653 (N_9653,N_8401,N_8703);
nand U9654 (N_9654,N_8017,N_8875);
nand U9655 (N_9655,N_8209,N_8339);
nand U9656 (N_9656,N_8292,N_8324);
and U9657 (N_9657,N_8463,N_8403);
nor U9658 (N_9658,N_8071,N_8020);
nand U9659 (N_9659,N_8566,N_8160);
and U9660 (N_9660,N_8775,N_8809);
or U9661 (N_9661,N_8762,N_8513);
or U9662 (N_9662,N_8200,N_8182);
xor U9663 (N_9663,N_8890,N_8463);
or U9664 (N_9664,N_8393,N_8476);
and U9665 (N_9665,N_8553,N_8128);
or U9666 (N_9666,N_8713,N_8360);
xnor U9667 (N_9667,N_8619,N_8695);
or U9668 (N_9668,N_8637,N_8362);
nand U9669 (N_9669,N_8900,N_8931);
and U9670 (N_9670,N_8177,N_8000);
nor U9671 (N_9671,N_8425,N_8319);
or U9672 (N_9672,N_8340,N_8220);
and U9673 (N_9673,N_8508,N_8087);
or U9674 (N_9674,N_8737,N_8849);
nor U9675 (N_9675,N_8196,N_8600);
nor U9676 (N_9676,N_8911,N_8675);
or U9677 (N_9677,N_8068,N_8560);
nor U9678 (N_9678,N_8109,N_8742);
nor U9679 (N_9679,N_8257,N_8096);
nand U9680 (N_9680,N_8271,N_8364);
nor U9681 (N_9681,N_8245,N_8359);
nor U9682 (N_9682,N_8866,N_8895);
or U9683 (N_9683,N_8337,N_8957);
and U9684 (N_9684,N_8505,N_8281);
or U9685 (N_9685,N_8515,N_8017);
nor U9686 (N_9686,N_8541,N_8820);
or U9687 (N_9687,N_8456,N_8828);
nor U9688 (N_9688,N_8582,N_8233);
and U9689 (N_9689,N_8565,N_8700);
xnor U9690 (N_9690,N_8020,N_8602);
nor U9691 (N_9691,N_8012,N_8785);
xnor U9692 (N_9692,N_8564,N_8130);
xnor U9693 (N_9693,N_8182,N_8305);
and U9694 (N_9694,N_8433,N_8261);
nand U9695 (N_9695,N_8796,N_8992);
or U9696 (N_9696,N_8926,N_8645);
or U9697 (N_9697,N_8198,N_8156);
or U9698 (N_9698,N_8392,N_8063);
nand U9699 (N_9699,N_8420,N_8644);
or U9700 (N_9700,N_8520,N_8743);
or U9701 (N_9701,N_8043,N_8646);
xor U9702 (N_9702,N_8723,N_8830);
nand U9703 (N_9703,N_8772,N_8202);
nand U9704 (N_9704,N_8253,N_8838);
xnor U9705 (N_9705,N_8160,N_8831);
xnor U9706 (N_9706,N_8039,N_8801);
or U9707 (N_9707,N_8137,N_8086);
nand U9708 (N_9708,N_8530,N_8919);
nand U9709 (N_9709,N_8324,N_8497);
nor U9710 (N_9710,N_8087,N_8011);
nand U9711 (N_9711,N_8449,N_8533);
or U9712 (N_9712,N_8539,N_8688);
or U9713 (N_9713,N_8244,N_8496);
or U9714 (N_9714,N_8580,N_8327);
nor U9715 (N_9715,N_8474,N_8283);
nor U9716 (N_9716,N_8089,N_8171);
and U9717 (N_9717,N_8736,N_8314);
or U9718 (N_9718,N_8607,N_8163);
and U9719 (N_9719,N_8600,N_8565);
or U9720 (N_9720,N_8226,N_8039);
and U9721 (N_9721,N_8625,N_8853);
xnor U9722 (N_9722,N_8149,N_8168);
and U9723 (N_9723,N_8473,N_8017);
nand U9724 (N_9724,N_8288,N_8167);
nor U9725 (N_9725,N_8697,N_8582);
or U9726 (N_9726,N_8192,N_8491);
nor U9727 (N_9727,N_8438,N_8156);
and U9728 (N_9728,N_8070,N_8807);
and U9729 (N_9729,N_8858,N_8078);
or U9730 (N_9730,N_8451,N_8036);
nand U9731 (N_9731,N_8130,N_8625);
and U9732 (N_9732,N_8056,N_8552);
nor U9733 (N_9733,N_8402,N_8500);
nand U9734 (N_9734,N_8098,N_8298);
nor U9735 (N_9735,N_8014,N_8902);
or U9736 (N_9736,N_8045,N_8049);
and U9737 (N_9737,N_8809,N_8108);
nand U9738 (N_9738,N_8461,N_8722);
and U9739 (N_9739,N_8882,N_8864);
and U9740 (N_9740,N_8562,N_8161);
or U9741 (N_9741,N_8017,N_8191);
nand U9742 (N_9742,N_8342,N_8979);
nand U9743 (N_9743,N_8556,N_8805);
or U9744 (N_9744,N_8824,N_8466);
or U9745 (N_9745,N_8277,N_8308);
nor U9746 (N_9746,N_8648,N_8284);
and U9747 (N_9747,N_8778,N_8712);
and U9748 (N_9748,N_8668,N_8713);
and U9749 (N_9749,N_8558,N_8985);
nor U9750 (N_9750,N_8915,N_8445);
nor U9751 (N_9751,N_8600,N_8465);
and U9752 (N_9752,N_8638,N_8681);
and U9753 (N_9753,N_8354,N_8970);
and U9754 (N_9754,N_8027,N_8554);
nor U9755 (N_9755,N_8476,N_8186);
nand U9756 (N_9756,N_8567,N_8842);
and U9757 (N_9757,N_8901,N_8475);
nor U9758 (N_9758,N_8359,N_8889);
or U9759 (N_9759,N_8214,N_8242);
nand U9760 (N_9760,N_8946,N_8917);
xor U9761 (N_9761,N_8227,N_8305);
nand U9762 (N_9762,N_8271,N_8527);
nor U9763 (N_9763,N_8583,N_8154);
nand U9764 (N_9764,N_8274,N_8255);
nor U9765 (N_9765,N_8885,N_8371);
and U9766 (N_9766,N_8484,N_8572);
or U9767 (N_9767,N_8183,N_8473);
and U9768 (N_9768,N_8173,N_8408);
nor U9769 (N_9769,N_8072,N_8598);
nor U9770 (N_9770,N_8897,N_8499);
nand U9771 (N_9771,N_8962,N_8744);
or U9772 (N_9772,N_8937,N_8914);
nand U9773 (N_9773,N_8557,N_8290);
or U9774 (N_9774,N_8941,N_8926);
nand U9775 (N_9775,N_8884,N_8541);
or U9776 (N_9776,N_8367,N_8965);
xnor U9777 (N_9777,N_8611,N_8505);
or U9778 (N_9778,N_8013,N_8633);
nor U9779 (N_9779,N_8519,N_8734);
and U9780 (N_9780,N_8289,N_8587);
and U9781 (N_9781,N_8780,N_8156);
nand U9782 (N_9782,N_8244,N_8994);
or U9783 (N_9783,N_8436,N_8829);
and U9784 (N_9784,N_8841,N_8629);
and U9785 (N_9785,N_8899,N_8833);
and U9786 (N_9786,N_8239,N_8699);
nand U9787 (N_9787,N_8968,N_8160);
and U9788 (N_9788,N_8956,N_8625);
and U9789 (N_9789,N_8299,N_8141);
xor U9790 (N_9790,N_8568,N_8206);
or U9791 (N_9791,N_8167,N_8644);
xor U9792 (N_9792,N_8188,N_8006);
nor U9793 (N_9793,N_8273,N_8314);
nor U9794 (N_9794,N_8488,N_8339);
nand U9795 (N_9795,N_8799,N_8135);
xor U9796 (N_9796,N_8605,N_8059);
nand U9797 (N_9797,N_8575,N_8056);
and U9798 (N_9798,N_8201,N_8512);
nor U9799 (N_9799,N_8594,N_8624);
nor U9800 (N_9800,N_8922,N_8082);
or U9801 (N_9801,N_8166,N_8404);
nor U9802 (N_9802,N_8052,N_8075);
nor U9803 (N_9803,N_8078,N_8587);
and U9804 (N_9804,N_8901,N_8354);
or U9805 (N_9805,N_8338,N_8538);
nor U9806 (N_9806,N_8955,N_8426);
nand U9807 (N_9807,N_8058,N_8527);
or U9808 (N_9808,N_8660,N_8114);
and U9809 (N_9809,N_8154,N_8964);
or U9810 (N_9810,N_8006,N_8480);
nand U9811 (N_9811,N_8674,N_8239);
or U9812 (N_9812,N_8309,N_8242);
and U9813 (N_9813,N_8493,N_8050);
or U9814 (N_9814,N_8150,N_8830);
and U9815 (N_9815,N_8121,N_8104);
and U9816 (N_9816,N_8962,N_8376);
nor U9817 (N_9817,N_8276,N_8234);
or U9818 (N_9818,N_8085,N_8928);
nand U9819 (N_9819,N_8291,N_8467);
or U9820 (N_9820,N_8185,N_8191);
or U9821 (N_9821,N_8378,N_8470);
and U9822 (N_9822,N_8854,N_8306);
nand U9823 (N_9823,N_8163,N_8116);
nand U9824 (N_9824,N_8423,N_8720);
nand U9825 (N_9825,N_8409,N_8739);
xnor U9826 (N_9826,N_8807,N_8831);
nand U9827 (N_9827,N_8253,N_8478);
nand U9828 (N_9828,N_8727,N_8040);
xor U9829 (N_9829,N_8210,N_8743);
nor U9830 (N_9830,N_8645,N_8585);
xnor U9831 (N_9831,N_8034,N_8140);
or U9832 (N_9832,N_8551,N_8085);
nand U9833 (N_9833,N_8613,N_8132);
xnor U9834 (N_9834,N_8724,N_8974);
and U9835 (N_9835,N_8271,N_8336);
nand U9836 (N_9836,N_8652,N_8668);
nor U9837 (N_9837,N_8540,N_8753);
nor U9838 (N_9838,N_8158,N_8166);
nand U9839 (N_9839,N_8971,N_8214);
xnor U9840 (N_9840,N_8141,N_8575);
xor U9841 (N_9841,N_8160,N_8112);
and U9842 (N_9842,N_8068,N_8999);
or U9843 (N_9843,N_8923,N_8822);
nor U9844 (N_9844,N_8917,N_8325);
nor U9845 (N_9845,N_8082,N_8248);
and U9846 (N_9846,N_8657,N_8562);
or U9847 (N_9847,N_8840,N_8504);
or U9848 (N_9848,N_8373,N_8552);
nor U9849 (N_9849,N_8874,N_8998);
and U9850 (N_9850,N_8126,N_8715);
and U9851 (N_9851,N_8011,N_8977);
nor U9852 (N_9852,N_8496,N_8326);
or U9853 (N_9853,N_8374,N_8691);
and U9854 (N_9854,N_8890,N_8483);
nor U9855 (N_9855,N_8582,N_8802);
nor U9856 (N_9856,N_8478,N_8291);
and U9857 (N_9857,N_8170,N_8573);
xor U9858 (N_9858,N_8198,N_8382);
xor U9859 (N_9859,N_8882,N_8855);
or U9860 (N_9860,N_8180,N_8098);
and U9861 (N_9861,N_8664,N_8694);
and U9862 (N_9862,N_8626,N_8544);
and U9863 (N_9863,N_8049,N_8496);
or U9864 (N_9864,N_8292,N_8781);
nand U9865 (N_9865,N_8352,N_8881);
xor U9866 (N_9866,N_8988,N_8493);
xor U9867 (N_9867,N_8668,N_8969);
nor U9868 (N_9868,N_8588,N_8771);
xnor U9869 (N_9869,N_8083,N_8638);
and U9870 (N_9870,N_8262,N_8292);
or U9871 (N_9871,N_8087,N_8771);
or U9872 (N_9872,N_8652,N_8584);
and U9873 (N_9873,N_8867,N_8941);
or U9874 (N_9874,N_8697,N_8957);
nor U9875 (N_9875,N_8020,N_8529);
or U9876 (N_9876,N_8777,N_8533);
or U9877 (N_9877,N_8586,N_8681);
nor U9878 (N_9878,N_8923,N_8143);
nand U9879 (N_9879,N_8158,N_8569);
nor U9880 (N_9880,N_8877,N_8194);
nand U9881 (N_9881,N_8070,N_8582);
nor U9882 (N_9882,N_8985,N_8356);
or U9883 (N_9883,N_8639,N_8250);
nor U9884 (N_9884,N_8757,N_8616);
nor U9885 (N_9885,N_8725,N_8802);
and U9886 (N_9886,N_8502,N_8818);
nand U9887 (N_9887,N_8571,N_8531);
or U9888 (N_9888,N_8396,N_8666);
or U9889 (N_9889,N_8418,N_8586);
nor U9890 (N_9890,N_8070,N_8889);
nor U9891 (N_9891,N_8431,N_8818);
nand U9892 (N_9892,N_8812,N_8076);
or U9893 (N_9893,N_8997,N_8549);
nor U9894 (N_9894,N_8175,N_8358);
nor U9895 (N_9895,N_8907,N_8961);
nor U9896 (N_9896,N_8257,N_8002);
xnor U9897 (N_9897,N_8447,N_8995);
nor U9898 (N_9898,N_8753,N_8998);
and U9899 (N_9899,N_8110,N_8697);
nand U9900 (N_9900,N_8427,N_8725);
nor U9901 (N_9901,N_8065,N_8834);
or U9902 (N_9902,N_8708,N_8153);
nand U9903 (N_9903,N_8253,N_8345);
or U9904 (N_9904,N_8798,N_8097);
and U9905 (N_9905,N_8229,N_8618);
or U9906 (N_9906,N_8013,N_8854);
nor U9907 (N_9907,N_8179,N_8747);
or U9908 (N_9908,N_8900,N_8088);
and U9909 (N_9909,N_8790,N_8405);
nor U9910 (N_9910,N_8319,N_8776);
nand U9911 (N_9911,N_8514,N_8027);
nor U9912 (N_9912,N_8227,N_8792);
xor U9913 (N_9913,N_8377,N_8074);
or U9914 (N_9914,N_8278,N_8974);
and U9915 (N_9915,N_8195,N_8654);
or U9916 (N_9916,N_8728,N_8569);
or U9917 (N_9917,N_8205,N_8889);
and U9918 (N_9918,N_8832,N_8797);
nand U9919 (N_9919,N_8494,N_8104);
nand U9920 (N_9920,N_8574,N_8108);
or U9921 (N_9921,N_8052,N_8427);
and U9922 (N_9922,N_8698,N_8736);
and U9923 (N_9923,N_8559,N_8884);
or U9924 (N_9924,N_8738,N_8254);
xnor U9925 (N_9925,N_8489,N_8861);
nand U9926 (N_9926,N_8096,N_8600);
nor U9927 (N_9927,N_8213,N_8309);
nor U9928 (N_9928,N_8863,N_8016);
xor U9929 (N_9929,N_8396,N_8279);
nand U9930 (N_9930,N_8627,N_8866);
nand U9931 (N_9931,N_8001,N_8919);
or U9932 (N_9932,N_8425,N_8530);
nor U9933 (N_9933,N_8535,N_8047);
and U9934 (N_9934,N_8754,N_8924);
nand U9935 (N_9935,N_8088,N_8503);
and U9936 (N_9936,N_8880,N_8597);
nor U9937 (N_9937,N_8449,N_8221);
nand U9938 (N_9938,N_8227,N_8729);
nor U9939 (N_9939,N_8370,N_8180);
and U9940 (N_9940,N_8390,N_8681);
nand U9941 (N_9941,N_8576,N_8452);
and U9942 (N_9942,N_8166,N_8927);
nor U9943 (N_9943,N_8216,N_8985);
and U9944 (N_9944,N_8326,N_8065);
nand U9945 (N_9945,N_8110,N_8579);
or U9946 (N_9946,N_8444,N_8372);
nor U9947 (N_9947,N_8697,N_8278);
or U9948 (N_9948,N_8101,N_8767);
nand U9949 (N_9949,N_8292,N_8014);
nand U9950 (N_9950,N_8999,N_8928);
nand U9951 (N_9951,N_8983,N_8158);
nor U9952 (N_9952,N_8790,N_8850);
and U9953 (N_9953,N_8667,N_8230);
and U9954 (N_9954,N_8158,N_8788);
nand U9955 (N_9955,N_8107,N_8880);
or U9956 (N_9956,N_8536,N_8783);
or U9957 (N_9957,N_8258,N_8530);
nand U9958 (N_9958,N_8302,N_8706);
and U9959 (N_9959,N_8471,N_8810);
or U9960 (N_9960,N_8917,N_8773);
and U9961 (N_9961,N_8369,N_8780);
xnor U9962 (N_9962,N_8932,N_8181);
or U9963 (N_9963,N_8754,N_8884);
and U9964 (N_9964,N_8167,N_8752);
or U9965 (N_9965,N_8211,N_8294);
and U9966 (N_9966,N_8339,N_8059);
or U9967 (N_9967,N_8755,N_8992);
nand U9968 (N_9968,N_8410,N_8576);
nor U9969 (N_9969,N_8950,N_8689);
or U9970 (N_9970,N_8059,N_8703);
and U9971 (N_9971,N_8199,N_8545);
xor U9972 (N_9972,N_8644,N_8139);
or U9973 (N_9973,N_8091,N_8305);
xor U9974 (N_9974,N_8988,N_8925);
or U9975 (N_9975,N_8362,N_8316);
xnor U9976 (N_9976,N_8679,N_8905);
and U9977 (N_9977,N_8025,N_8385);
nand U9978 (N_9978,N_8839,N_8808);
nor U9979 (N_9979,N_8562,N_8196);
nand U9980 (N_9980,N_8094,N_8262);
and U9981 (N_9981,N_8616,N_8593);
nor U9982 (N_9982,N_8524,N_8174);
nand U9983 (N_9983,N_8540,N_8284);
nor U9984 (N_9984,N_8078,N_8701);
nand U9985 (N_9985,N_8681,N_8271);
nand U9986 (N_9986,N_8570,N_8950);
nor U9987 (N_9987,N_8628,N_8857);
nand U9988 (N_9988,N_8930,N_8833);
or U9989 (N_9989,N_8640,N_8812);
nand U9990 (N_9990,N_8388,N_8035);
nand U9991 (N_9991,N_8067,N_8742);
or U9992 (N_9992,N_8700,N_8205);
and U9993 (N_9993,N_8179,N_8723);
and U9994 (N_9994,N_8835,N_8519);
or U9995 (N_9995,N_8400,N_8481);
xnor U9996 (N_9996,N_8364,N_8223);
nand U9997 (N_9997,N_8858,N_8955);
or U9998 (N_9998,N_8886,N_8636);
nand U9999 (N_9999,N_8467,N_8875);
or U10000 (N_10000,N_9458,N_9820);
nor U10001 (N_10001,N_9270,N_9715);
nand U10002 (N_10002,N_9767,N_9823);
nor U10003 (N_10003,N_9911,N_9514);
xor U10004 (N_10004,N_9214,N_9080);
nand U10005 (N_10005,N_9440,N_9895);
or U10006 (N_10006,N_9757,N_9240);
and U10007 (N_10007,N_9495,N_9184);
or U10008 (N_10008,N_9225,N_9663);
and U10009 (N_10009,N_9671,N_9811);
or U10010 (N_10010,N_9208,N_9108);
and U10011 (N_10011,N_9350,N_9325);
or U10012 (N_10012,N_9993,N_9346);
or U10013 (N_10013,N_9349,N_9500);
or U10014 (N_10014,N_9436,N_9309);
and U10015 (N_10015,N_9157,N_9571);
nor U10016 (N_10016,N_9907,N_9683);
nor U10017 (N_10017,N_9211,N_9931);
or U10018 (N_10018,N_9394,N_9796);
or U10019 (N_10019,N_9024,N_9424);
or U10020 (N_10020,N_9432,N_9611);
xor U10021 (N_10021,N_9568,N_9827);
nor U10022 (N_10022,N_9178,N_9520);
or U10023 (N_10023,N_9244,N_9552);
or U10024 (N_10024,N_9737,N_9076);
or U10025 (N_10025,N_9430,N_9065);
and U10026 (N_10026,N_9973,N_9173);
or U10027 (N_10027,N_9885,N_9170);
xnor U10028 (N_10028,N_9083,N_9402);
nor U10029 (N_10029,N_9762,N_9978);
and U10030 (N_10030,N_9097,N_9861);
nand U10031 (N_10031,N_9155,N_9620);
xnor U10032 (N_10032,N_9171,N_9860);
and U10033 (N_10033,N_9769,N_9738);
xnor U10034 (N_10034,N_9238,N_9412);
nand U10035 (N_10035,N_9179,N_9467);
and U10036 (N_10036,N_9853,N_9073);
nand U10037 (N_10037,N_9233,N_9708);
nand U10038 (N_10038,N_9582,N_9988);
and U10039 (N_10039,N_9169,N_9718);
nand U10040 (N_10040,N_9049,N_9797);
nand U10041 (N_10041,N_9360,N_9926);
and U10042 (N_10042,N_9289,N_9351);
and U10043 (N_10043,N_9296,N_9857);
nand U10044 (N_10044,N_9743,N_9254);
and U10045 (N_10045,N_9121,N_9417);
nand U10046 (N_10046,N_9995,N_9116);
or U10047 (N_10047,N_9471,N_9426);
xnor U10048 (N_10048,N_9947,N_9256);
nor U10049 (N_10049,N_9129,N_9835);
nor U10050 (N_10050,N_9992,N_9069);
and U10051 (N_10051,N_9052,N_9475);
nor U10052 (N_10052,N_9186,N_9175);
xnor U10053 (N_10053,N_9508,N_9604);
xnor U10054 (N_10054,N_9450,N_9519);
xor U10055 (N_10055,N_9927,N_9493);
or U10056 (N_10056,N_9573,N_9026);
nand U10057 (N_10057,N_9451,N_9834);
nor U10058 (N_10058,N_9567,N_9779);
nand U10059 (N_10059,N_9209,N_9333);
nand U10060 (N_10060,N_9729,N_9785);
and U10061 (N_10061,N_9628,N_9373);
and U10062 (N_10062,N_9643,N_9269);
and U10063 (N_10063,N_9122,N_9196);
or U10064 (N_10064,N_9848,N_9476);
xnor U10065 (N_10065,N_9282,N_9151);
and U10066 (N_10066,N_9093,N_9913);
or U10067 (N_10067,N_9422,N_9599);
nor U10068 (N_10068,N_9691,N_9572);
nor U10069 (N_10069,N_9974,N_9938);
or U10070 (N_10070,N_9388,N_9539);
nor U10071 (N_10071,N_9301,N_9286);
and U10072 (N_10072,N_9385,N_9403);
nor U10073 (N_10073,N_9665,N_9112);
nand U10074 (N_10074,N_9940,N_9361);
and U10075 (N_10075,N_9088,N_9057);
xnor U10076 (N_10076,N_9427,N_9871);
xor U10077 (N_10077,N_9874,N_9198);
nor U10078 (N_10078,N_9676,N_9644);
nand U10079 (N_10079,N_9159,N_9594);
or U10080 (N_10080,N_9949,N_9210);
and U10081 (N_10081,N_9692,N_9919);
or U10082 (N_10082,N_9852,N_9790);
and U10083 (N_10083,N_9677,N_9841);
nor U10084 (N_10084,N_9405,N_9952);
nor U10085 (N_10085,N_9353,N_9425);
nand U10086 (N_10086,N_9845,N_9008);
nor U10087 (N_10087,N_9660,N_9124);
and U10088 (N_10088,N_9344,N_9058);
or U10089 (N_10089,N_9487,N_9929);
and U10090 (N_10090,N_9684,N_9123);
nand U10091 (N_10091,N_9858,N_9043);
nor U10092 (N_10092,N_9367,N_9750);
and U10093 (N_10093,N_9255,N_9366);
nand U10094 (N_10094,N_9051,N_9881);
nor U10095 (N_10095,N_9386,N_9113);
nand U10096 (N_10096,N_9951,N_9488);
nor U10097 (N_10097,N_9066,N_9085);
and U10098 (N_10098,N_9987,N_9530);
nor U10099 (N_10099,N_9923,N_9239);
nor U10100 (N_10100,N_9261,N_9017);
or U10101 (N_10101,N_9001,N_9358);
nor U10102 (N_10102,N_9106,N_9616);
nor U10103 (N_10103,N_9580,N_9204);
nor U10104 (N_10104,N_9730,N_9783);
xnor U10105 (N_10105,N_9401,N_9545);
or U10106 (N_10106,N_9292,N_9777);
xnor U10107 (N_10107,N_9236,N_9682);
nand U10108 (N_10108,N_9936,N_9110);
and U10109 (N_10109,N_9512,N_9321);
or U10110 (N_10110,N_9842,N_9521);
nor U10111 (N_10111,N_9818,N_9452);
xnor U10112 (N_10112,N_9142,N_9964);
nor U10113 (N_10113,N_9966,N_9391);
nor U10114 (N_10114,N_9011,N_9335);
or U10115 (N_10115,N_9562,N_9320);
xnor U10116 (N_10116,N_9633,N_9074);
or U10117 (N_10117,N_9924,N_9435);
or U10118 (N_10118,N_9522,N_9235);
xnor U10119 (N_10119,N_9429,N_9681);
nand U10120 (N_10120,N_9679,N_9339);
or U10121 (N_10121,N_9503,N_9946);
xor U10122 (N_10122,N_9190,N_9816);
and U10123 (N_10123,N_9498,N_9578);
nor U10124 (N_10124,N_9393,N_9880);
or U10125 (N_10125,N_9221,N_9437);
or U10126 (N_10126,N_9200,N_9598);
and U10127 (N_10127,N_9315,N_9004);
or U10128 (N_10128,N_9433,N_9119);
nor U10129 (N_10129,N_9457,N_9095);
nand U10130 (N_10130,N_9741,N_9478);
and U10131 (N_10131,N_9227,N_9185);
and U10132 (N_10132,N_9591,N_9299);
nand U10133 (N_10133,N_9833,N_9197);
and U10134 (N_10134,N_9039,N_9998);
or U10135 (N_10135,N_9021,N_9710);
or U10136 (N_10136,N_9831,N_9070);
nor U10137 (N_10137,N_9768,N_9917);
or U10138 (N_10138,N_9442,N_9517);
and U10139 (N_10139,N_9048,N_9593);
and U10140 (N_10140,N_9002,N_9559);
nor U10141 (N_10141,N_9300,N_9023);
nor U10142 (N_10142,N_9844,N_9318);
nand U10143 (N_10143,N_9400,N_9824);
or U10144 (N_10144,N_9370,N_9601);
or U10145 (N_10145,N_9975,N_9307);
nor U10146 (N_10146,N_9415,N_9870);
nand U10147 (N_10147,N_9647,N_9212);
nor U10148 (N_10148,N_9690,N_9053);
nor U10149 (N_10149,N_9584,N_9484);
or U10150 (N_10150,N_9480,N_9075);
nand U10151 (N_10151,N_9543,N_9202);
nand U10152 (N_10152,N_9609,N_9094);
nand U10153 (N_10153,N_9701,N_9772);
or U10154 (N_10154,N_9986,N_9306);
and U10155 (N_10155,N_9461,N_9996);
or U10156 (N_10156,N_9516,N_9983);
and U10157 (N_10157,N_9194,N_9656);
and U10158 (N_10158,N_9213,N_9629);
or U10159 (N_10159,N_9332,N_9859);
xor U10160 (N_10160,N_9133,N_9152);
and U10161 (N_10161,N_9589,N_9968);
and U10162 (N_10162,N_9161,N_9542);
nor U10163 (N_10163,N_9406,N_9943);
nor U10164 (N_10164,N_9587,N_9937);
nor U10165 (N_10165,N_9727,N_9970);
nor U10166 (N_10166,N_9253,N_9003);
xnor U10167 (N_10167,N_9932,N_9814);
nand U10168 (N_10168,N_9680,N_9265);
and U10169 (N_10169,N_9341,N_9794);
nand U10170 (N_10170,N_9696,N_9409);
nand U10171 (N_10171,N_9600,N_9804);
and U10172 (N_10172,N_9028,N_9810);
xor U10173 (N_10173,N_9398,N_9780);
or U10174 (N_10174,N_9303,N_9372);
or U10175 (N_10175,N_9061,N_9836);
xnor U10176 (N_10176,N_9808,N_9613);
nand U10177 (N_10177,N_9063,N_9231);
nor U10178 (N_10178,N_9109,N_9379);
nor U10179 (N_10179,N_9087,N_9215);
nand U10180 (N_10180,N_9150,N_9532);
nand U10181 (N_10181,N_9511,N_9251);
or U10182 (N_10182,N_9592,N_9954);
and U10183 (N_10183,N_9447,N_9483);
nand U10184 (N_10184,N_9252,N_9877);
nor U10185 (N_10185,N_9693,N_9506);
and U10186 (N_10186,N_9275,N_9368);
nor U10187 (N_10187,N_9298,N_9470);
or U10188 (N_10188,N_9149,N_9217);
and U10189 (N_10189,N_9637,N_9618);
nor U10190 (N_10190,N_9807,N_9421);
xor U10191 (N_10191,N_9297,N_9581);
nor U10192 (N_10192,N_9898,N_9548);
nor U10193 (N_10193,N_9362,N_9262);
nor U10194 (N_10194,N_9802,N_9799);
xor U10195 (N_10195,N_9268,N_9359);
nand U10196 (N_10196,N_9771,N_9625);
xor U10197 (N_10197,N_9101,N_9466);
or U10198 (N_10198,N_9164,N_9384);
and U10199 (N_10199,N_9634,N_9441);
nand U10200 (N_10200,N_9626,N_9603);
or U10201 (N_10201,N_9704,N_9977);
nand U10202 (N_10202,N_9688,N_9364);
and U10203 (N_10203,N_9960,N_9719);
or U10204 (N_10204,N_9781,N_9886);
and U10205 (N_10205,N_9419,N_9279);
xor U10206 (N_10206,N_9764,N_9355);
nor U10207 (N_10207,N_9033,N_9846);
and U10208 (N_10208,N_9013,N_9672);
nand U10209 (N_10209,N_9906,N_9955);
or U10210 (N_10210,N_9959,N_9020);
nand U10211 (N_10211,N_9939,N_9830);
or U10212 (N_10212,N_9163,N_9192);
or U10213 (N_10213,N_9272,N_9027);
or U10214 (N_10214,N_9037,N_9237);
and U10215 (N_10215,N_9733,N_9042);
xnor U10216 (N_10216,N_9759,N_9153);
and U10217 (N_10217,N_9761,N_9915);
nand U10218 (N_10218,N_9904,N_9054);
and U10219 (N_10219,N_9854,N_9099);
or U10220 (N_10220,N_9553,N_9188);
and U10221 (N_10221,N_9675,N_9100);
nand U10222 (N_10222,N_9742,N_9642);
or U10223 (N_10223,N_9181,N_9882);
nor U10224 (N_10224,N_9577,N_9566);
nor U10225 (N_10225,N_9574,N_9728);
nand U10226 (N_10226,N_9563,N_9492);
xor U10227 (N_10227,N_9795,N_9472);
xor U10228 (N_10228,N_9617,N_9380);
nor U10229 (N_10229,N_9815,N_9878);
and U10230 (N_10230,N_9961,N_9407);
nor U10231 (N_10231,N_9850,N_9312);
or U10232 (N_10232,N_9868,N_9136);
or U10233 (N_10233,N_9006,N_9029);
nor U10234 (N_10234,N_9131,N_9957);
and U10235 (N_10235,N_9867,N_9336);
and U10236 (N_10236,N_9132,N_9050);
nand U10237 (N_10237,N_9847,N_9126);
nand U10238 (N_10238,N_9597,N_9328);
nor U10239 (N_10239,N_9605,N_9277);
nor U10240 (N_10240,N_9242,N_9507);
and U10241 (N_10241,N_9007,N_9338);
nand U10242 (N_10242,N_9148,N_9486);
nor U10243 (N_10243,N_9956,N_9645);
and U10244 (N_10244,N_9736,N_9014);
and U10245 (N_10245,N_9334,N_9851);
and U10246 (N_10246,N_9707,N_9792);
xnor U10247 (N_10247,N_9144,N_9305);
nand U10248 (N_10248,N_9176,N_9260);
xnor U10249 (N_10249,N_9428,N_9524);
or U10250 (N_10250,N_9285,N_9245);
nor U10251 (N_10251,N_9224,N_9758);
nand U10252 (N_10252,N_9979,N_9264);
and U10253 (N_10253,N_9474,N_9127);
or U10254 (N_10254,N_9230,N_9313);
nand U10255 (N_10255,N_9935,N_9473);
nor U10256 (N_10256,N_9031,N_9342);
and U10257 (N_10257,N_9056,N_9627);
xor U10258 (N_10258,N_9655,N_9716);
xnor U10259 (N_10259,N_9047,N_9523);
xnor U10260 (N_10260,N_9717,N_9304);
xnor U10261 (N_10261,N_9840,N_9195);
or U10262 (N_10262,N_9653,N_9894);
nand U10263 (N_10263,N_9032,N_9250);
nand U10264 (N_10264,N_9963,N_9143);
nand U10265 (N_10265,N_9773,N_9182);
or U10266 (N_10266,N_9377,N_9751);
nand U10267 (N_10267,N_9259,N_9431);
nand U10268 (N_10268,N_9748,N_9310);
nand U10269 (N_10269,N_9501,N_9639);
or U10270 (N_10270,N_9739,N_9942);
nand U10271 (N_10271,N_9413,N_9535);
xnor U10272 (N_10272,N_9775,N_9283);
or U10273 (N_10273,N_9725,N_9763);
nor U10274 (N_10274,N_9243,N_9103);
nand U10275 (N_10275,N_9754,N_9079);
nand U10276 (N_10276,N_9348,N_9928);
and U10277 (N_10277,N_9482,N_9547);
or U10278 (N_10278,N_9137,N_9722);
nand U10279 (N_10279,N_9753,N_9345);
nand U10280 (N_10280,N_9068,N_9549);
nor U10281 (N_10281,N_9558,N_9546);
xor U10282 (N_10282,N_9019,N_9135);
nor U10283 (N_10283,N_9219,N_9976);
nor U10284 (N_10284,N_9000,N_9766);
nor U10285 (N_10285,N_9223,N_9865);
or U10286 (N_10286,N_9557,N_9776);
nand U10287 (N_10287,N_9381,N_9104);
nor U10288 (N_10288,N_9491,N_9788);
and U10289 (N_10289,N_9556,N_9371);
and U10290 (N_10290,N_9167,N_9276);
or U10291 (N_10291,N_9570,N_9651);
and U10292 (N_10292,N_9241,N_9347);
and U10293 (N_10293,N_9891,N_9786);
nor U10294 (N_10294,N_9658,N_9396);
and U10295 (N_10295,N_9327,N_9839);
nor U10296 (N_10296,N_9463,N_9791);
and U10297 (N_10297,N_9699,N_9669);
xor U10298 (N_10298,N_9843,N_9034);
nand U10299 (N_10299,N_9632,N_9879);
and U10300 (N_10300,N_9485,N_9141);
nor U10301 (N_10301,N_9005,N_9443);
nor U10302 (N_10302,N_9555,N_9612);
xor U10303 (N_10303,N_9838,N_9117);
nand U10304 (N_10304,N_9295,N_9308);
nor U10305 (N_10305,N_9703,N_9528);
or U10306 (N_10306,N_9965,N_9569);
nand U10307 (N_10307,N_9908,N_9071);
nor U10308 (N_10308,N_9046,N_9218);
and U10309 (N_10309,N_9969,N_9229);
and U10310 (N_10310,N_9468,N_9293);
nand U10311 (N_10311,N_9111,N_9872);
or U10312 (N_10312,N_9608,N_9652);
nand U10313 (N_10313,N_9529,N_9925);
nor U10314 (N_10314,N_9944,N_9331);
or U10315 (N_10315,N_9661,N_9010);
and U10316 (N_10316,N_9294,N_9274);
and U10317 (N_10317,N_9089,N_9096);
or U10318 (N_10318,N_9686,N_9774);
nor U10319 (N_10319,N_9726,N_9174);
or U10320 (N_10320,N_9712,N_9025);
or U10321 (N_10321,N_9374,N_9948);
and U10322 (N_10322,N_9564,N_9438);
or U10323 (N_10323,N_9550,N_9525);
xnor U10324 (N_10324,N_9869,N_9165);
nand U10325 (N_10325,N_9356,N_9551);
nand U10326 (N_10326,N_9921,N_9803);
nand U10327 (N_10327,N_9410,N_9787);
and U10328 (N_10328,N_9752,N_9317);
xnor U10329 (N_10329,N_9271,N_9278);
nand U10330 (N_10330,N_9694,N_9950);
nor U10331 (N_10331,N_9756,N_9984);
or U10332 (N_10332,N_9670,N_9418);
or U10333 (N_10333,N_9674,N_9041);
xor U10334 (N_10334,N_9631,N_9232);
xor U10335 (N_10335,N_9228,N_9082);
nor U10336 (N_10336,N_9392,N_9090);
or U10337 (N_10337,N_9990,N_9630);
nor U10338 (N_10338,N_9395,N_9586);
and U10339 (N_10339,N_9258,N_9622);
nand U10340 (N_10340,N_9449,N_9565);
or U10341 (N_10341,N_9453,N_9343);
or U10342 (N_10342,N_9247,N_9903);
and U10343 (N_10343,N_9900,N_9092);
and U10344 (N_10344,N_9585,N_9896);
and U10345 (N_10345,N_9249,N_9806);
or U10346 (N_10346,N_9789,N_9575);
nor U10347 (N_10347,N_9504,N_9376);
nor U10348 (N_10348,N_9291,N_9825);
nand U10349 (N_10349,N_9664,N_9765);
nor U10350 (N_10350,N_9183,N_9914);
and U10351 (N_10351,N_9352,N_9724);
or U10352 (N_10352,N_9387,N_9160);
or U10353 (N_10353,N_9454,N_9784);
nand U10354 (N_10354,N_9828,N_9060);
or U10355 (N_10355,N_9246,N_9641);
nand U10356 (N_10356,N_9740,N_9981);
xnor U10357 (N_10357,N_9972,N_9624);
nor U10358 (N_10358,N_9561,N_9234);
and U10359 (N_10359,N_9105,N_9832);
and U10360 (N_10360,N_9875,N_9505);
nand U10361 (N_10361,N_9445,N_9448);
or U10362 (N_10362,N_9280,N_9798);
nor U10363 (N_10363,N_9678,N_9770);
and U10364 (N_10364,N_9540,N_9420);
nor U10365 (N_10365,N_9337,N_9809);
nor U10366 (N_10366,N_9905,N_9864);
or U10367 (N_10367,N_9889,N_9311);
and U10368 (N_10368,N_9813,N_9078);
xnor U10369 (N_10369,N_9615,N_9702);
xor U10370 (N_10370,N_9901,N_9330);
nor U10371 (N_10371,N_9933,N_9720);
xnor U10372 (N_10372,N_9140,N_9967);
and U10373 (N_10373,N_9460,N_9399);
or U10374 (N_10374,N_9554,N_9817);
nand U10375 (N_10375,N_9888,N_9316);
nor U10376 (N_10376,N_9201,N_9579);
and U10377 (N_10377,N_9668,N_9700);
or U10378 (N_10378,N_9156,N_9375);
and U10379 (N_10379,N_9172,N_9793);
or U10380 (N_10380,N_9389,N_9267);
nor U10381 (N_10381,N_9538,N_9821);
xnor U10382 (N_10382,N_9439,N_9610);
nand U10383 (N_10383,N_9829,N_9583);
and U10384 (N_10384,N_9685,N_9128);
nor U10385 (N_10385,N_9494,N_9866);
or U10386 (N_10386,N_9994,N_9837);
or U10387 (N_10387,N_9062,N_9499);
and U10388 (N_10388,N_9084,N_9030);
or U10389 (N_10389,N_9953,N_9745);
nand U10390 (N_10390,N_9576,N_9513);
xnor U10391 (N_10391,N_9216,N_9081);
nor U10392 (N_10392,N_9098,N_9180);
nor U10393 (N_10393,N_9302,N_9248);
nand U10394 (N_10394,N_9281,N_9922);
and U10395 (N_10395,N_9411,N_9654);
nor U10396 (N_10396,N_9456,N_9623);
and U10397 (N_10397,N_9640,N_9365);
or U10398 (N_10398,N_9731,N_9910);
and U10399 (N_10399,N_9502,N_9962);
xor U10400 (N_10400,N_9036,N_9273);
nand U10401 (N_10401,N_9012,N_9897);
nor U10402 (N_10402,N_9189,N_9490);
or U10403 (N_10403,N_9035,N_9287);
nor U10404 (N_10404,N_9390,N_9714);
and U10405 (N_10405,N_9314,N_9383);
nor U10406 (N_10406,N_9022,N_9746);
nor U10407 (N_10407,N_9607,N_9177);
nor U10408 (N_10408,N_9689,N_9469);
nor U10409 (N_10409,N_9744,N_9920);
and U10410 (N_10410,N_9883,N_9414);
and U10411 (N_10411,N_9755,N_9462);
nor U10412 (N_10412,N_9226,N_9635);
nor U10413 (N_10413,N_9064,N_9510);
or U10414 (N_10414,N_9222,N_9544);
nor U10415 (N_10415,N_9697,N_9077);
and U10416 (N_10416,N_9166,N_9114);
nor U10417 (N_10417,N_9091,N_9489);
xnor U10418 (N_10418,N_9072,N_9408);
nor U10419 (N_10419,N_9340,N_9884);
or U10420 (N_10420,N_9369,N_9941);
nand U10421 (N_10421,N_9638,N_9536);
and U10422 (N_10422,N_9997,N_9706);
nor U10423 (N_10423,N_9203,N_9560);
nand U10424 (N_10424,N_9596,N_9404);
nand U10425 (N_10425,N_9760,N_9782);
nor U10426 (N_10426,N_9687,N_9481);
nand U10427 (N_10427,N_9899,N_9902);
nand U10428 (N_10428,N_9734,N_9735);
or U10429 (N_10429,N_9059,N_9323);
nor U10430 (N_10430,N_9606,N_9162);
xnor U10431 (N_10431,N_9206,N_9541);
xnor U10432 (N_10432,N_9588,N_9397);
or U10433 (N_10433,N_9934,N_9705);
nand U10434 (N_10434,N_9115,N_9916);
nand U10435 (N_10435,N_9518,N_9444);
xor U10436 (N_10436,N_9354,N_9434);
nand U10437 (N_10437,N_9721,N_9288);
nor U10438 (N_10438,N_9357,N_9199);
nor U10439 (N_10439,N_9120,N_9045);
and U10440 (N_10440,N_9863,N_9892);
and U10441 (N_10441,N_9319,N_9455);
nand U10442 (N_10442,N_9220,N_9849);
nand U10443 (N_10443,N_9855,N_9732);
nand U10444 (N_10444,N_9650,N_9266);
nand U10445 (N_10445,N_9477,N_9146);
nand U10446 (N_10446,N_9497,N_9018);
xor U10447 (N_10447,N_9107,N_9086);
and U10448 (N_10448,N_9648,N_9909);
xor U10449 (N_10449,N_9531,N_9659);
or U10450 (N_10450,N_9749,N_9912);
nand U10451 (N_10451,N_9322,N_9464);
or U10452 (N_10452,N_9055,N_9038);
or U10453 (N_10453,N_9595,N_9812);
nor U10454 (N_10454,N_9856,N_9695);
nor U10455 (N_10455,N_9980,N_9709);
nand U10456 (N_10456,N_9590,N_9329);
nor U10457 (N_10457,N_9147,N_9805);
and U10458 (N_10458,N_9971,N_9862);
or U10459 (N_10459,N_9991,N_9711);
nand U10460 (N_10460,N_9667,N_9636);
nand U10461 (N_10461,N_9154,N_9040);
or U10462 (N_10462,N_9930,N_9999);
and U10463 (N_10463,N_9778,N_9819);
nand U10464 (N_10464,N_9826,N_9290);
nor U10465 (N_10465,N_9465,N_9324);
and U10466 (N_10466,N_9191,N_9459);
and U10467 (N_10467,N_9378,N_9193);
nand U10468 (N_10468,N_9662,N_9666);
nand U10469 (N_10469,N_9534,N_9257);
or U10470 (N_10470,N_9893,N_9982);
nand U10471 (N_10471,N_9800,N_9207);
nor U10472 (N_10472,N_9887,N_9145);
or U10473 (N_10473,N_9723,N_9890);
nand U10474 (N_10474,N_9263,N_9158);
or U10475 (N_10475,N_9918,N_9713);
xnor U10476 (N_10476,N_9284,N_9958);
nor U10477 (N_10477,N_9118,N_9168);
nand U10478 (N_10478,N_9646,N_9125);
or U10479 (N_10479,N_9363,N_9326);
nand U10480 (N_10480,N_9602,N_9945);
or U10481 (N_10481,N_9446,N_9673);
nand U10482 (N_10482,N_9649,N_9423);
or U10483 (N_10483,N_9130,N_9016);
and U10484 (N_10484,N_9015,N_9496);
nand U10485 (N_10485,N_9985,N_9537);
nor U10486 (N_10486,N_9009,N_9382);
nand U10487 (N_10487,N_9134,N_9526);
nor U10488 (N_10488,N_9657,N_9989);
nor U10489 (N_10489,N_9527,N_9533);
nor U10490 (N_10490,N_9416,N_9614);
nor U10491 (N_10491,N_9044,N_9619);
nand U10492 (N_10492,N_9509,N_9515);
nand U10493 (N_10493,N_9102,N_9873);
and U10494 (N_10494,N_9479,N_9801);
nor U10495 (N_10495,N_9747,N_9698);
nor U10496 (N_10496,N_9876,N_9067);
and U10497 (N_10497,N_9139,N_9138);
and U10498 (N_10498,N_9822,N_9205);
nand U10499 (N_10499,N_9621,N_9187);
nand U10500 (N_10500,N_9897,N_9678);
nand U10501 (N_10501,N_9708,N_9707);
nand U10502 (N_10502,N_9952,N_9023);
and U10503 (N_10503,N_9243,N_9454);
and U10504 (N_10504,N_9756,N_9325);
and U10505 (N_10505,N_9755,N_9240);
xnor U10506 (N_10506,N_9694,N_9851);
nor U10507 (N_10507,N_9598,N_9013);
nand U10508 (N_10508,N_9349,N_9246);
nor U10509 (N_10509,N_9888,N_9522);
nand U10510 (N_10510,N_9196,N_9070);
and U10511 (N_10511,N_9406,N_9693);
and U10512 (N_10512,N_9175,N_9540);
nor U10513 (N_10513,N_9835,N_9989);
or U10514 (N_10514,N_9665,N_9174);
nand U10515 (N_10515,N_9048,N_9024);
nor U10516 (N_10516,N_9087,N_9280);
or U10517 (N_10517,N_9537,N_9271);
and U10518 (N_10518,N_9230,N_9562);
xnor U10519 (N_10519,N_9365,N_9653);
nand U10520 (N_10520,N_9887,N_9594);
nand U10521 (N_10521,N_9420,N_9929);
nor U10522 (N_10522,N_9162,N_9421);
nor U10523 (N_10523,N_9783,N_9633);
xnor U10524 (N_10524,N_9085,N_9872);
nor U10525 (N_10525,N_9414,N_9261);
nor U10526 (N_10526,N_9459,N_9176);
or U10527 (N_10527,N_9999,N_9685);
xor U10528 (N_10528,N_9592,N_9975);
nand U10529 (N_10529,N_9328,N_9385);
nand U10530 (N_10530,N_9709,N_9454);
nor U10531 (N_10531,N_9783,N_9263);
nand U10532 (N_10532,N_9184,N_9774);
and U10533 (N_10533,N_9449,N_9099);
or U10534 (N_10534,N_9668,N_9735);
or U10535 (N_10535,N_9611,N_9081);
or U10536 (N_10536,N_9422,N_9374);
and U10537 (N_10537,N_9898,N_9539);
xnor U10538 (N_10538,N_9789,N_9034);
and U10539 (N_10539,N_9315,N_9798);
nor U10540 (N_10540,N_9969,N_9464);
or U10541 (N_10541,N_9287,N_9697);
nand U10542 (N_10542,N_9749,N_9250);
nor U10543 (N_10543,N_9911,N_9321);
or U10544 (N_10544,N_9644,N_9099);
nand U10545 (N_10545,N_9741,N_9760);
xor U10546 (N_10546,N_9183,N_9610);
and U10547 (N_10547,N_9833,N_9754);
nand U10548 (N_10548,N_9476,N_9022);
and U10549 (N_10549,N_9704,N_9301);
nand U10550 (N_10550,N_9734,N_9251);
or U10551 (N_10551,N_9943,N_9172);
xnor U10552 (N_10552,N_9785,N_9608);
and U10553 (N_10553,N_9826,N_9300);
nand U10554 (N_10554,N_9533,N_9088);
nor U10555 (N_10555,N_9908,N_9848);
xor U10556 (N_10556,N_9079,N_9812);
nand U10557 (N_10557,N_9395,N_9858);
and U10558 (N_10558,N_9221,N_9051);
and U10559 (N_10559,N_9089,N_9775);
nand U10560 (N_10560,N_9398,N_9142);
or U10561 (N_10561,N_9346,N_9975);
or U10562 (N_10562,N_9007,N_9633);
or U10563 (N_10563,N_9555,N_9297);
nand U10564 (N_10564,N_9476,N_9935);
or U10565 (N_10565,N_9055,N_9917);
or U10566 (N_10566,N_9436,N_9580);
and U10567 (N_10567,N_9707,N_9718);
nand U10568 (N_10568,N_9199,N_9482);
nand U10569 (N_10569,N_9321,N_9408);
or U10570 (N_10570,N_9783,N_9493);
xor U10571 (N_10571,N_9639,N_9148);
nand U10572 (N_10572,N_9360,N_9668);
xnor U10573 (N_10573,N_9928,N_9462);
or U10574 (N_10574,N_9512,N_9247);
or U10575 (N_10575,N_9607,N_9962);
nor U10576 (N_10576,N_9584,N_9416);
xor U10577 (N_10577,N_9495,N_9920);
and U10578 (N_10578,N_9925,N_9776);
or U10579 (N_10579,N_9351,N_9573);
nor U10580 (N_10580,N_9761,N_9610);
nand U10581 (N_10581,N_9732,N_9355);
and U10582 (N_10582,N_9941,N_9655);
or U10583 (N_10583,N_9895,N_9395);
nand U10584 (N_10584,N_9373,N_9086);
and U10585 (N_10585,N_9259,N_9950);
and U10586 (N_10586,N_9025,N_9686);
nand U10587 (N_10587,N_9732,N_9492);
nand U10588 (N_10588,N_9325,N_9592);
nand U10589 (N_10589,N_9658,N_9035);
xor U10590 (N_10590,N_9579,N_9407);
and U10591 (N_10591,N_9700,N_9795);
or U10592 (N_10592,N_9578,N_9942);
and U10593 (N_10593,N_9214,N_9440);
nor U10594 (N_10594,N_9723,N_9783);
nor U10595 (N_10595,N_9864,N_9669);
nor U10596 (N_10596,N_9744,N_9424);
or U10597 (N_10597,N_9135,N_9416);
nand U10598 (N_10598,N_9427,N_9691);
nand U10599 (N_10599,N_9947,N_9136);
or U10600 (N_10600,N_9766,N_9812);
or U10601 (N_10601,N_9730,N_9737);
or U10602 (N_10602,N_9467,N_9351);
nor U10603 (N_10603,N_9287,N_9786);
nand U10604 (N_10604,N_9820,N_9123);
nor U10605 (N_10605,N_9945,N_9898);
or U10606 (N_10606,N_9910,N_9848);
and U10607 (N_10607,N_9622,N_9507);
nor U10608 (N_10608,N_9411,N_9681);
nor U10609 (N_10609,N_9081,N_9778);
and U10610 (N_10610,N_9755,N_9320);
and U10611 (N_10611,N_9556,N_9061);
or U10612 (N_10612,N_9525,N_9886);
or U10613 (N_10613,N_9738,N_9964);
or U10614 (N_10614,N_9133,N_9798);
nor U10615 (N_10615,N_9054,N_9079);
nand U10616 (N_10616,N_9063,N_9504);
and U10617 (N_10617,N_9195,N_9841);
or U10618 (N_10618,N_9680,N_9407);
or U10619 (N_10619,N_9419,N_9614);
or U10620 (N_10620,N_9094,N_9117);
nand U10621 (N_10621,N_9328,N_9432);
xnor U10622 (N_10622,N_9609,N_9566);
and U10623 (N_10623,N_9881,N_9366);
nand U10624 (N_10624,N_9017,N_9403);
or U10625 (N_10625,N_9501,N_9083);
nor U10626 (N_10626,N_9744,N_9104);
or U10627 (N_10627,N_9932,N_9498);
nand U10628 (N_10628,N_9514,N_9042);
or U10629 (N_10629,N_9930,N_9597);
and U10630 (N_10630,N_9551,N_9355);
or U10631 (N_10631,N_9109,N_9356);
or U10632 (N_10632,N_9219,N_9398);
or U10633 (N_10633,N_9151,N_9798);
nand U10634 (N_10634,N_9718,N_9620);
or U10635 (N_10635,N_9398,N_9611);
and U10636 (N_10636,N_9651,N_9905);
nor U10637 (N_10637,N_9225,N_9834);
nor U10638 (N_10638,N_9298,N_9742);
or U10639 (N_10639,N_9958,N_9896);
or U10640 (N_10640,N_9877,N_9225);
nand U10641 (N_10641,N_9726,N_9830);
xnor U10642 (N_10642,N_9830,N_9626);
and U10643 (N_10643,N_9910,N_9324);
or U10644 (N_10644,N_9642,N_9329);
or U10645 (N_10645,N_9006,N_9429);
or U10646 (N_10646,N_9969,N_9483);
nand U10647 (N_10647,N_9781,N_9026);
xnor U10648 (N_10648,N_9650,N_9365);
and U10649 (N_10649,N_9861,N_9144);
nand U10650 (N_10650,N_9314,N_9127);
nand U10651 (N_10651,N_9321,N_9690);
nor U10652 (N_10652,N_9842,N_9907);
or U10653 (N_10653,N_9759,N_9605);
nand U10654 (N_10654,N_9847,N_9556);
and U10655 (N_10655,N_9997,N_9553);
or U10656 (N_10656,N_9319,N_9116);
and U10657 (N_10657,N_9688,N_9124);
nor U10658 (N_10658,N_9466,N_9647);
or U10659 (N_10659,N_9279,N_9111);
nor U10660 (N_10660,N_9312,N_9069);
and U10661 (N_10661,N_9746,N_9179);
nor U10662 (N_10662,N_9048,N_9580);
and U10663 (N_10663,N_9056,N_9024);
nor U10664 (N_10664,N_9861,N_9757);
nor U10665 (N_10665,N_9155,N_9446);
xnor U10666 (N_10666,N_9677,N_9049);
nand U10667 (N_10667,N_9601,N_9627);
and U10668 (N_10668,N_9955,N_9799);
nor U10669 (N_10669,N_9515,N_9506);
nor U10670 (N_10670,N_9714,N_9873);
nor U10671 (N_10671,N_9763,N_9829);
nor U10672 (N_10672,N_9824,N_9065);
xor U10673 (N_10673,N_9547,N_9065);
or U10674 (N_10674,N_9085,N_9723);
and U10675 (N_10675,N_9226,N_9673);
nand U10676 (N_10676,N_9938,N_9779);
or U10677 (N_10677,N_9779,N_9538);
nor U10678 (N_10678,N_9805,N_9298);
xnor U10679 (N_10679,N_9963,N_9382);
nand U10680 (N_10680,N_9453,N_9814);
nand U10681 (N_10681,N_9875,N_9229);
or U10682 (N_10682,N_9984,N_9966);
xor U10683 (N_10683,N_9682,N_9885);
or U10684 (N_10684,N_9440,N_9515);
or U10685 (N_10685,N_9507,N_9496);
nand U10686 (N_10686,N_9982,N_9089);
nand U10687 (N_10687,N_9938,N_9337);
or U10688 (N_10688,N_9760,N_9080);
nor U10689 (N_10689,N_9641,N_9391);
xnor U10690 (N_10690,N_9594,N_9033);
nand U10691 (N_10691,N_9269,N_9386);
or U10692 (N_10692,N_9102,N_9198);
nor U10693 (N_10693,N_9123,N_9882);
nor U10694 (N_10694,N_9229,N_9395);
xnor U10695 (N_10695,N_9654,N_9746);
and U10696 (N_10696,N_9243,N_9053);
xnor U10697 (N_10697,N_9555,N_9217);
nor U10698 (N_10698,N_9091,N_9275);
nor U10699 (N_10699,N_9844,N_9679);
or U10700 (N_10700,N_9212,N_9576);
and U10701 (N_10701,N_9961,N_9353);
nand U10702 (N_10702,N_9684,N_9292);
or U10703 (N_10703,N_9126,N_9596);
nand U10704 (N_10704,N_9631,N_9332);
and U10705 (N_10705,N_9223,N_9946);
nand U10706 (N_10706,N_9920,N_9958);
xnor U10707 (N_10707,N_9848,N_9778);
nor U10708 (N_10708,N_9167,N_9757);
nand U10709 (N_10709,N_9542,N_9723);
nand U10710 (N_10710,N_9937,N_9992);
nand U10711 (N_10711,N_9406,N_9851);
nor U10712 (N_10712,N_9021,N_9781);
nor U10713 (N_10713,N_9085,N_9888);
nand U10714 (N_10714,N_9189,N_9745);
nand U10715 (N_10715,N_9787,N_9030);
nand U10716 (N_10716,N_9137,N_9951);
xor U10717 (N_10717,N_9084,N_9867);
nand U10718 (N_10718,N_9645,N_9606);
xnor U10719 (N_10719,N_9940,N_9732);
and U10720 (N_10720,N_9514,N_9531);
and U10721 (N_10721,N_9303,N_9803);
and U10722 (N_10722,N_9647,N_9500);
nor U10723 (N_10723,N_9409,N_9276);
xor U10724 (N_10724,N_9826,N_9314);
and U10725 (N_10725,N_9456,N_9132);
nor U10726 (N_10726,N_9346,N_9333);
nand U10727 (N_10727,N_9617,N_9314);
xnor U10728 (N_10728,N_9250,N_9996);
nand U10729 (N_10729,N_9042,N_9725);
nand U10730 (N_10730,N_9502,N_9013);
and U10731 (N_10731,N_9030,N_9488);
nand U10732 (N_10732,N_9514,N_9841);
nor U10733 (N_10733,N_9143,N_9676);
nand U10734 (N_10734,N_9483,N_9272);
or U10735 (N_10735,N_9095,N_9427);
or U10736 (N_10736,N_9319,N_9355);
and U10737 (N_10737,N_9153,N_9808);
nand U10738 (N_10738,N_9870,N_9775);
nor U10739 (N_10739,N_9476,N_9497);
or U10740 (N_10740,N_9064,N_9735);
and U10741 (N_10741,N_9840,N_9002);
and U10742 (N_10742,N_9330,N_9789);
nand U10743 (N_10743,N_9344,N_9015);
nand U10744 (N_10744,N_9597,N_9693);
nand U10745 (N_10745,N_9091,N_9805);
nand U10746 (N_10746,N_9056,N_9166);
nand U10747 (N_10747,N_9230,N_9290);
and U10748 (N_10748,N_9702,N_9200);
nor U10749 (N_10749,N_9615,N_9551);
nand U10750 (N_10750,N_9605,N_9280);
nor U10751 (N_10751,N_9680,N_9627);
and U10752 (N_10752,N_9825,N_9863);
or U10753 (N_10753,N_9637,N_9365);
and U10754 (N_10754,N_9230,N_9451);
nor U10755 (N_10755,N_9362,N_9680);
or U10756 (N_10756,N_9227,N_9100);
nand U10757 (N_10757,N_9979,N_9309);
xor U10758 (N_10758,N_9857,N_9400);
or U10759 (N_10759,N_9490,N_9295);
nor U10760 (N_10760,N_9129,N_9974);
and U10761 (N_10761,N_9890,N_9530);
nand U10762 (N_10762,N_9536,N_9242);
nand U10763 (N_10763,N_9821,N_9837);
nor U10764 (N_10764,N_9016,N_9236);
or U10765 (N_10765,N_9727,N_9157);
xnor U10766 (N_10766,N_9252,N_9683);
or U10767 (N_10767,N_9065,N_9279);
and U10768 (N_10768,N_9097,N_9910);
nor U10769 (N_10769,N_9021,N_9780);
nor U10770 (N_10770,N_9832,N_9141);
nand U10771 (N_10771,N_9220,N_9500);
nand U10772 (N_10772,N_9767,N_9554);
nand U10773 (N_10773,N_9697,N_9680);
and U10774 (N_10774,N_9150,N_9278);
or U10775 (N_10775,N_9093,N_9903);
nor U10776 (N_10776,N_9403,N_9257);
nor U10777 (N_10777,N_9629,N_9188);
nand U10778 (N_10778,N_9371,N_9792);
or U10779 (N_10779,N_9275,N_9599);
and U10780 (N_10780,N_9562,N_9268);
xor U10781 (N_10781,N_9962,N_9281);
nor U10782 (N_10782,N_9168,N_9841);
and U10783 (N_10783,N_9372,N_9220);
or U10784 (N_10784,N_9427,N_9250);
nand U10785 (N_10785,N_9653,N_9275);
and U10786 (N_10786,N_9340,N_9533);
or U10787 (N_10787,N_9356,N_9298);
nor U10788 (N_10788,N_9732,N_9352);
nor U10789 (N_10789,N_9578,N_9168);
nor U10790 (N_10790,N_9697,N_9406);
nand U10791 (N_10791,N_9538,N_9376);
nand U10792 (N_10792,N_9285,N_9314);
xor U10793 (N_10793,N_9689,N_9886);
or U10794 (N_10794,N_9319,N_9216);
nor U10795 (N_10795,N_9794,N_9889);
and U10796 (N_10796,N_9190,N_9939);
xnor U10797 (N_10797,N_9960,N_9614);
and U10798 (N_10798,N_9964,N_9251);
nor U10799 (N_10799,N_9424,N_9402);
nor U10800 (N_10800,N_9232,N_9484);
or U10801 (N_10801,N_9661,N_9313);
or U10802 (N_10802,N_9008,N_9450);
or U10803 (N_10803,N_9627,N_9330);
or U10804 (N_10804,N_9823,N_9533);
nor U10805 (N_10805,N_9446,N_9766);
and U10806 (N_10806,N_9766,N_9773);
or U10807 (N_10807,N_9480,N_9563);
or U10808 (N_10808,N_9576,N_9902);
or U10809 (N_10809,N_9118,N_9406);
nor U10810 (N_10810,N_9829,N_9476);
nor U10811 (N_10811,N_9964,N_9678);
nor U10812 (N_10812,N_9401,N_9414);
and U10813 (N_10813,N_9580,N_9673);
or U10814 (N_10814,N_9730,N_9455);
or U10815 (N_10815,N_9691,N_9466);
nor U10816 (N_10816,N_9592,N_9448);
and U10817 (N_10817,N_9856,N_9677);
and U10818 (N_10818,N_9382,N_9299);
nand U10819 (N_10819,N_9467,N_9263);
nor U10820 (N_10820,N_9939,N_9998);
nor U10821 (N_10821,N_9839,N_9539);
xnor U10822 (N_10822,N_9805,N_9936);
xnor U10823 (N_10823,N_9801,N_9033);
nor U10824 (N_10824,N_9113,N_9699);
nor U10825 (N_10825,N_9452,N_9174);
nand U10826 (N_10826,N_9820,N_9550);
or U10827 (N_10827,N_9924,N_9326);
nor U10828 (N_10828,N_9744,N_9260);
nand U10829 (N_10829,N_9351,N_9353);
and U10830 (N_10830,N_9855,N_9309);
and U10831 (N_10831,N_9619,N_9268);
nor U10832 (N_10832,N_9956,N_9425);
nand U10833 (N_10833,N_9063,N_9925);
or U10834 (N_10834,N_9424,N_9598);
or U10835 (N_10835,N_9271,N_9140);
or U10836 (N_10836,N_9677,N_9125);
nand U10837 (N_10837,N_9186,N_9403);
nand U10838 (N_10838,N_9514,N_9701);
nor U10839 (N_10839,N_9846,N_9895);
and U10840 (N_10840,N_9282,N_9919);
and U10841 (N_10841,N_9860,N_9004);
nand U10842 (N_10842,N_9845,N_9345);
nor U10843 (N_10843,N_9235,N_9462);
nor U10844 (N_10844,N_9240,N_9196);
and U10845 (N_10845,N_9950,N_9292);
or U10846 (N_10846,N_9474,N_9791);
nand U10847 (N_10847,N_9784,N_9444);
or U10848 (N_10848,N_9731,N_9162);
and U10849 (N_10849,N_9325,N_9596);
or U10850 (N_10850,N_9732,N_9041);
and U10851 (N_10851,N_9611,N_9378);
or U10852 (N_10852,N_9684,N_9824);
nor U10853 (N_10853,N_9965,N_9957);
xor U10854 (N_10854,N_9371,N_9921);
or U10855 (N_10855,N_9324,N_9088);
nand U10856 (N_10856,N_9970,N_9700);
nand U10857 (N_10857,N_9197,N_9731);
or U10858 (N_10858,N_9883,N_9069);
xor U10859 (N_10859,N_9337,N_9482);
nand U10860 (N_10860,N_9645,N_9898);
and U10861 (N_10861,N_9017,N_9137);
or U10862 (N_10862,N_9049,N_9675);
nand U10863 (N_10863,N_9591,N_9854);
or U10864 (N_10864,N_9267,N_9117);
nand U10865 (N_10865,N_9775,N_9930);
nand U10866 (N_10866,N_9827,N_9660);
or U10867 (N_10867,N_9755,N_9348);
nor U10868 (N_10868,N_9147,N_9857);
nand U10869 (N_10869,N_9904,N_9088);
and U10870 (N_10870,N_9501,N_9488);
nand U10871 (N_10871,N_9193,N_9576);
nor U10872 (N_10872,N_9672,N_9559);
nor U10873 (N_10873,N_9863,N_9805);
nor U10874 (N_10874,N_9472,N_9674);
and U10875 (N_10875,N_9384,N_9583);
and U10876 (N_10876,N_9197,N_9750);
nand U10877 (N_10877,N_9983,N_9929);
or U10878 (N_10878,N_9484,N_9186);
nor U10879 (N_10879,N_9763,N_9994);
nand U10880 (N_10880,N_9251,N_9086);
xor U10881 (N_10881,N_9038,N_9240);
or U10882 (N_10882,N_9111,N_9800);
nand U10883 (N_10883,N_9683,N_9856);
or U10884 (N_10884,N_9401,N_9462);
and U10885 (N_10885,N_9271,N_9748);
and U10886 (N_10886,N_9947,N_9073);
or U10887 (N_10887,N_9086,N_9199);
or U10888 (N_10888,N_9528,N_9967);
xor U10889 (N_10889,N_9073,N_9136);
nand U10890 (N_10890,N_9896,N_9175);
nand U10891 (N_10891,N_9875,N_9111);
nand U10892 (N_10892,N_9242,N_9804);
and U10893 (N_10893,N_9395,N_9259);
or U10894 (N_10894,N_9481,N_9095);
nor U10895 (N_10895,N_9433,N_9976);
and U10896 (N_10896,N_9603,N_9557);
nand U10897 (N_10897,N_9697,N_9395);
and U10898 (N_10898,N_9895,N_9506);
and U10899 (N_10899,N_9455,N_9769);
and U10900 (N_10900,N_9723,N_9822);
and U10901 (N_10901,N_9563,N_9443);
and U10902 (N_10902,N_9819,N_9761);
nand U10903 (N_10903,N_9301,N_9672);
nor U10904 (N_10904,N_9436,N_9069);
nand U10905 (N_10905,N_9370,N_9083);
nand U10906 (N_10906,N_9561,N_9403);
nand U10907 (N_10907,N_9389,N_9162);
and U10908 (N_10908,N_9257,N_9904);
or U10909 (N_10909,N_9473,N_9126);
nor U10910 (N_10910,N_9325,N_9215);
and U10911 (N_10911,N_9841,N_9780);
and U10912 (N_10912,N_9210,N_9673);
xor U10913 (N_10913,N_9562,N_9598);
or U10914 (N_10914,N_9752,N_9629);
nand U10915 (N_10915,N_9087,N_9641);
or U10916 (N_10916,N_9204,N_9507);
and U10917 (N_10917,N_9791,N_9472);
or U10918 (N_10918,N_9149,N_9048);
xnor U10919 (N_10919,N_9222,N_9918);
nand U10920 (N_10920,N_9424,N_9433);
or U10921 (N_10921,N_9169,N_9357);
nor U10922 (N_10922,N_9830,N_9116);
or U10923 (N_10923,N_9990,N_9046);
nand U10924 (N_10924,N_9438,N_9510);
nor U10925 (N_10925,N_9297,N_9271);
nand U10926 (N_10926,N_9732,N_9886);
xor U10927 (N_10927,N_9601,N_9881);
nand U10928 (N_10928,N_9725,N_9537);
nand U10929 (N_10929,N_9497,N_9413);
and U10930 (N_10930,N_9133,N_9681);
nor U10931 (N_10931,N_9775,N_9246);
and U10932 (N_10932,N_9972,N_9641);
xor U10933 (N_10933,N_9383,N_9005);
xor U10934 (N_10934,N_9585,N_9310);
and U10935 (N_10935,N_9423,N_9567);
and U10936 (N_10936,N_9066,N_9012);
nand U10937 (N_10937,N_9658,N_9335);
nand U10938 (N_10938,N_9463,N_9801);
xor U10939 (N_10939,N_9899,N_9831);
nand U10940 (N_10940,N_9278,N_9507);
and U10941 (N_10941,N_9376,N_9902);
or U10942 (N_10942,N_9592,N_9284);
xor U10943 (N_10943,N_9254,N_9656);
nand U10944 (N_10944,N_9635,N_9076);
and U10945 (N_10945,N_9011,N_9458);
or U10946 (N_10946,N_9584,N_9525);
nor U10947 (N_10947,N_9781,N_9442);
and U10948 (N_10948,N_9313,N_9684);
nand U10949 (N_10949,N_9456,N_9683);
and U10950 (N_10950,N_9787,N_9317);
nand U10951 (N_10951,N_9051,N_9333);
and U10952 (N_10952,N_9727,N_9452);
xnor U10953 (N_10953,N_9970,N_9186);
and U10954 (N_10954,N_9060,N_9759);
or U10955 (N_10955,N_9698,N_9313);
xor U10956 (N_10956,N_9542,N_9071);
or U10957 (N_10957,N_9712,N_9626);
xor U10958 (N_10958,N_9691,N_9902);
and U10959 (N_10959,N_9867,N_9357);
or U10960 (N_10960,N_9746,N_9360);
and U10961 (N_10961,N_9989,N_9951);
and U10962 (N_10962,N_9537,N_9634);
nand U10963 (N_10963,N_9085,N_9383);
nor U10964 (N_10964,N_9576,N_9003);
nor U10965 (N_10965,N_9621,N_9373);
nor U10966 (N_10966,N_9071,N_9145);
nand U10967 (N_10967,N_9335,N_9710);
or U10968 (N_10968,N_9139,N_9375);
nand U10969 (N_10969,N_9941,N_9548);
xnor U10970 (N_10970,N_9843,N_9141);
nor U10971 (N_10971,N_9061,N_9393);
nor U10972 (N_10972,N_9041,N_9117);
nand U10973 (N_10973,N_9067,N_9159);
and U10974 (N_10974,N_9973,N_9277);
nand U10975 (N_10975,N_9188,N_9939);
and U10976 (N_10976,N_9817,N_9193);
and U10977 (N_10977,N_9949,N_9025);
and U10978 (N_10978,N_9092,N_9216);
nor U10979 (N_10979,N_9395,N_9628);
and U10980 (N_10980,N_9587,N_9028);
and U10981 (N_10981,N_9701,N_9828);
xnor U10982 (N_10982,N_9136,N_9850);
and U10983 (N_10983,N_9196,N_9646);
and U10984 (N_10984,N_9091,N_9802);
and U10985 (N_10985,N_9911,N_9028);
or U10986 (N_10986,N_9861,N_9278);
nor U10987 (N_10987,N_9355,N_9199);
nand U10988 (N_10988,N_9303,N_9130);
and U10989 (N_10989,N_9390,N_9776);
nor U10990 (N_10990,N_9003,N_9674);
nand U10991 (N_10991,N_9572,N_9370);
nand U10992 (N_10992,N_9540,N_9040);
and U10993 (N_10993,N_9253,N_9153);
or U10994 (N_10994,N_9594,N_9172);
or U10995 (N_10995,N_9403,N_9657);
or U10996 (N_10996,N_9756,N_9879);
xor U10997 (N_10997,N_9687,N_9505);
and U10998 (N_10998,N_9052,N_9650);
and U10999 (N_10999,N_9646,N_9426);
nand U11000 (N_11000,N_10506,N_10042);
nand U11001 (N_11001,N_10673,N_10767);
nor U11002 (N_11002,N_10843,N_10408);
nor U11003 (N_11003,N_10264,N_10133);
nor U11004 (N_11004,N_10790,N_10505);
nand U11005 (N_11005,N_10924,N_10130);
nand U11006 (N_11006,N_10309,N_10791);
nor U11007 (N_11007,N_10737,N_10804);
nor U11008 (N_11008,N_10648,N_10836);
nand U11009 (N_11009,N_10046,N_10813);
and U11010 (N_11010,N_10221,N_10271);
nand U11011 (N_11011,N_10554,N_10805);
and U11012 (N_11012,N_10128,N_10519);
and U11013 (N_11013,N_10972,N_10549);
xor U11014 (N_11014,N_10329,N_10674);
nor U11015 (N_11015,N_10663,N_10390);
nand U11016 (N_11016,N_10706,N_10454);
or U11017 (N_11017,N_10644,N_10884);
or U11018 (N_11018,N_10085,N_10107);
xor U11019 (N_11019,N_10571,N_10212);
or U11020 (N_11020,N_10950,N_10341);
and U11021 (N_11021,N_10520,N_10470);
nand U11022 (N_11022,N_10627,N_10353);
nand U11023 (N_11023,N_10598,N_10686);
nor U11024 (N_11024,N_10382,N_10602);
nand U11025 (N_11025,N_10227,N_10536);
and U11026 (N_11026,N_10177,N_10297);
nor U11027 (N_11027,N_10287,N_10176);
nor U11028 (N_11028,N_10963,N_10181);
nor U11029 (N_11029,N_10149,N_10175);
nor U11030 (N_11030,N_10491,N_10040);
nand U11031 (N_11031,N_10858,N_10882);
and U11032 (N_11032,N_10386,N_10835);
nand U11033 (N_11033,N_10510,N_10546);
nor U11034 (N_11034,N_10240,N_10122);
nor U11035 (N_11035,N_10577,N_10684);
nor U11036 (N_11036,N_10490,N_10263);
or U11037 (N_11037,N_10411,N_10863);
and U11038 (N_11038,N_10944,N_10982);
nand U11039 (N_11039,N_10065,N_10051);
nor U11040 (N_11040,N_10129,N_10912);
nor U11041 (N_11041,N_10859,N_10292);
xor U11042 (N_11042,N_10529,N_10480);
and U11043 (N_11043,N_10504,N_10066);
and U11044 (N_11044,N_10985,N_10942);
nor U11045 (N_11045,N_10072,N_10270);
and U11046 (N_11046,N_10570,N_10330);
nor U11047 (N_11047,N_10855,N_10693);
or U11048 (N_11048,N_10245,N_10739);
and U11049 (N_11049,N_10731,N_10907);
nand U11050 (N_11050,N_10567,N_10643);
and U11051 (N_11051,N_10339,N_10239);
and U11052 (N_11052,N_10825,N_10032);
and U11053 (N_11053,N_10485,N_10868);
nor U11054 (N_11054,N_10679,N_10797);
nor U11055 (N_11055,N_10153,N_10180);
or U11056 (N_11056,N_10395,N_10246);
nor U11057 (N_11057,N_10438,N_10163);
nand U11058 (N_11058,N_10495,N_10310);
or U11059 (N_11059,N_10185,N_10012);
nor U11060 (N_11060,N_10487,N_10050);
and U11061 (N_11061,N_10917,N_10315);
and U11062 (N_11062,N_10933,N_10704);
nand U11063 (N_11063,N_10213,N_10318);
xor U11064 (N_11064,N_10630,N_10916);
nor U11065 (N_11065,N_10764,N_10187);
nor U11066 (N_11066,N_10286,N_10726);
or U11067 (N_11067,N_10594,N_10407);
nor U11068 (N_11068,N_10134,N_10711);
xnor U11069 (N_11069,N_10559,N_10344);
or U11070 (N_11070,N_10957,N_10492);
nand U11071 (N_11071,N_10342,N_10874);
xnor U11072 (N_11072,N_10174,N_10735);
or U11073 (N_11073,N_10477,N_10161);
and U11074 (N_11074,N_10325,N_10850);
and U11075 (N_11075,N_10038,N_10199);
nor U11076 (N_11076,N_10777,N_10540);
or U11077 (N_11077,N_10603,N_10772);
or U11078 (N_11078,N_10784,N_10381);
and U11079 (N_11079,N_10126,N_10494);
or U11080 (N_11080,N_10482,N_10727);
or U11081 (N_11081,N_10866,N_10336);
nand U11082 (N_11082,N_10771,N_10064);
or U11083 (N_11083,N_10593,N_10662);
or U11084 (N_11084,N_10834,N_10432);
nor U11085 (N_11085,N_10366,N_10397);
nor U11086 (N_11086,N_10458,N_10501);
and U11087 (N_11087,N_10139,N_10101);
and U11088 (N_11088,N_10111,N_10869);
nor U11089 (N_11089,N_10750,N_10734);
nor U11090 (N_11090,N_10160,N_10808);
nor U11091 (N_11091,N_10232,N_10707);
xor U11092 (N_11092,N_10024,N_10668);
xor U11093 (N_11093,N_10521,N_10523);
nor U11094 (N_11094,N_10682,N_10440);
nand U11095 (N_11095,N_10766,N_10569);
nor U11096 (N_11096,N_10090,N_10945);
nand U11097 (N_11097,N_10518,N_10483);
or U11098 (N_11098,N_10370,N_10465);
nand U11099 (N_11099,N_10178,N_10842);
nor U11100 (N_11100,N_10118,N_10755);
nand U11101 (N_11101,N_10113,N_10965);
and U11102 (N_11102,N_10345,N_10563);
and U11103 (N_11103,N_10304,N_10312);
nand U11104 (N_11104,N_10936,N_10335);
or U11105 (N_11105,N_10299,N_10967);
nand U11106 (N_11106,N_10516,N_10189);
nor U11107 (N_11107,N_10925,N_10851);
nor U11108 (N_11108,N_10200,N_10242);
nand U11109 (N_11109,N_10875,N_10588);
nand U11110 (N_11110,N_10419,N_10296);
nand U11111 (N_11111,N_10383,N_10496);
and U11112 (N_11112,N_10956,N_10452);
or U11113 (N_11113,N_10717,N_10226);
nand U11114 (N_11114,N_10604,N_10430);
nor U11115 (N_11115,N_10334,N_10898);
or U11116 (N_11116,N_10670,N_10459);
nand U11117 (N_11117,N_10481,N_10449);
nor U11118 (N_11118,N_10198,N_10098);
nand U11119 (N_11119,N_10471,N_10261);
or U11120 (N_11120,N_10574,N_10484);
or U11121 (N_11121,N_10014,N_10966);
xnor U11122 (N_11122,N_10436,N_10517);
and U11123 (N_11123,N_10155,N_10365);
nand U11124 (N_11124,N_10412,N_10154);
and U11125 (N_11125,N_10787,N_10624);
and U11126 (N_11126,N_10939,N_10416);
or U11127 (N_11127,N_10091,N_10252);
nor U11128 (N_11128,N_10020,N_10428);
and U11129 (N_11129,N_10317,N_10368);
nand U11130 (N_11130,N_10188,N_10075);
and U11131 (N_11131,N_10260,N_10691);
and U11132 (N_11132,N_10099,N_10741);
nor U11133 (N_11133,N_10981,N_10757);
nand U11134 (N_11134,N_10262,N_10337);
or U11135 (N_11135,N_10222,N_10887);
nor U11136 (N_11136,N_10530,N_10687);
nor U11137 (N_11137,N_10067,N_10142);
or U11138 (N_11138,N_10398,N_10970);
or U11139 (N_11139,N_10938,N_10906);
or U11140 (N_11140,N_10553,N_10612);
nor U11141 (N_11141,N_10675,N_10980);
nand U11142 (N_11142,N_10027,N_10993);
and U11143 (N_11143,N_10323,N_10632);
or U11144 (N_11144,N_10460,N_10307);
nor U11145 (N_11145,N_10247,N_10531);
xor U11146 (N_11146,N_10406,N_10558);
nor U11147 (N_11147,N_10902,N_10223);
or U11148 (N_11148,N_10838,N_10457);
and U11149 (N_11149,N_10280,N_10828);
and U11150 (N_11150,N_10584,N_10742);
nor U11151 (N_11151,N_10431,N_10006);
nand U11152 (N_11152,N_10702,N_10657);
nand U11153 (N_11153,N_10525,N_10217);
nor U11154 (N_11154,N_10231,N_10683);
or U11155 (N_11155,N_10900,N_10467);
nand U11156 (N_11156,N_10203,N_10968);
or U11157 (N_11157,N_10044,N_10388);
nor U11158 (N_11158,N_10953,N_10059);
or U11159 (N_11159,N_10782,N_10697);
and U11160 (N_11160,N_10753,N_10685);
xnor U11161 (N_11161,N_10745,N_10660);
or U11162 (N_11162,N_10705,N_10359);
and U11163 (N_11163,N_10442,N_10798);
xnor U11164 (N_11164,N_10961,N_10620);
nor U11165 (N_11165,N_10369,N_10417);
nor U11166 (N_11166,N_10669,N_10688);
or U11167 (N_11167,N_10761,N_10826);
nor U11168 (N_11168,N_10392,N_10427);
nor U11169 (N_11169,N_10690,N_10818);
or U11170 (N_11170,N_10311,N_10008);
or U11171 (N_11171,N_10303,N_10897);
nand U11172 (N_11172,N_10827,N_10197);
xor U11173 (N_11173,N_10255,N_10135);
or U11174 (N_11174,N_10182,N_10347);
nor U11175 (N_11175,N_10236,N_10638);
xor U11176 (N_11176,N_10049,N_10931);
nand U11177 (N_11177,N_10300,N_10812);
or U11178 (N_11178,N_10581,N_10057);
or U11179 (N_11179,N_10807,N_10324);
nand U11180 (N_11180,N_10783,N_10003);
or U11181 (N_11181,N_10589,N_10551);
nor U11182 (N_11182,N_10780,N_10533);
nor U11183 (N_11183,N_10733,N_10087);
nand U11184 (N_11184,N_10977,N_10082);
nor U11185 (N_11185,N_10201,N_10418);
nand U11186 (N_11186,N_10526,N_10384);
nor U11187 (N_11187,N_10606,N_10173);
nor U11188 (N_11188,N_10448,N_10909);
nor U11189 (N_11189,N_10940,N_10946);
nand U11190 (N_11190,N_10768,N_10656);
nor U11191 (N_11191,N_10722,N_10026);
and U11192 (N_11192,N_10959,N_10964);
nor U11193 (N_11193,N_10877,N_10441);
or U11194 (N_11194,N_10011,N_10932);
and U11195 (N_11195,N_10241,N_10018);
nand U11196 (N_11196,N_10935,N_10860);
and U11197 (N_11197,N_10746,N_10689);
or U11198 (N_11198,N_10796,N_10186);
or U11199 (N_11199,N_10566,N_10852);
nand U11200 (N_11200,N_10209,N_10385);
xor U11201 (N_11201,N_10695,N_10216);
xnor U11202 (N_11202,N_10387,N_10105);
nor U11203 (N_11203,N_10379,N_10327);
nand U11204 (N_11204,N_10081,N_10910);
and U11205 (N_11205,N_10234,N_10035);
nand U11206 (N_11206,N_10775,N_10166);
and U11207 (N_11207,N_10016,N_10502);
nor U11208 (N_11208,N_10019,N_10658);
nor U11209 (N_11209,N_10439,N_10524);
or U11210 (N_11210,N_10819,N_10845);
xnor U11211 (N_11211,N_10522,N_10774);
nor U11212 (N_11212,N_10595,N_10815);
or U11213 (N_11213,N_10928,N_10844);
nor U11214 (N_11214,N_10269,N_10478);
and U11215 (N_11215,N_10760,N_10713);
or U11216 (N_11216,N_10360,N_10219);
nor U11217 (N_11217,N_10076,N_10915);
nor U11218 (N_11218,N_10943,N_10306);
xor U11219 (N_11219,N_10565,N_10375);
and U11220 (N_11220,N_10374,N_10641);
xor U11221 (N_11221,N_10749,N_10393);
nor U11222 (N_11222,N_10556,N_10279);
nand U11223 (N_11223,N_10389,N_10779);
and U11224 (N_11224,N_10747,N_10272);
nand U11225 (N_11225,N_10572,N_10196);
nand U11226 (N_11226,N_10476,N_10308);
and U11227 (N_11227,N_10194,N_10031);
nor U11228 (N_11228,N_10541,N_10116);
nand U11229 (N_11229,N_10718,N_10251);
or U11230 (N_11230,N_10999,N_10290);
or U11231 (N_11231,N_10616,N_10429);
and U11232 (N_11232,N_10396,N_10672);
nand U11233 (N_11233,N_10990,N_10028);
or U11234 (N_11234,N_10853,N_10547);
and U11235 (N_11235,N_10973,N_10215);
or U11236 (N_11236,N_10088,N_10888);
or U11237 (N_11237,N_10880,N_10424);
or U11238 (N_11238,N_10168,N_10824);
nor U11239 (N_11239,N_10507,N_10350);
and U11240 (N_11240,N_10991,N_10047);
nand U11241 (N_11241,N_10921,N_10948);
and U11242 (N_11242,N_10511,N_10413);
xor U11243 (N_11243,N_10822,N_10840);
and U11244 (N_11244,N_10409,N_10354);
nor U11245 (N_11245,N_10585,N_10754);
nand U11246 (N_11246,N_10738,N_10445);
nand U11247 (N_11247,N_10109,N_10839);
nor U11248 (N_11248,N_10282,N_10022);
nand U11249 (N_11249,N_10911,N_10238);
nand U11250 (N_11250,N_10205,N_10351);
and U11251 (N_11251,N_10810,N_10821);
and U11252 (N_11252,N_10462,N_10415);
nor U11253 (N_11253,N_10146,N_10137);
or U11254 (N_11254,N_10361,N_10293);
or U11255 (N_11255,N_10914,N_10131);
or U11256 (N_11256,N_10534,N_10343);
and U11257 (N_11257,N_10895,N_10710);
or U11258 (N_11258,N_10614,N_10698);
nand U11259 (N_11259,N_10642,N_10358);
xor U11260 (N_11260,N_10106,N_10714);
nand U11261 (N_11261,N_10002,N_10979);
and U11262 (N_11262,N_10623,N_10652);
or U11263 (N_11263,N_10041,N_10294);
or U11264 (N_11264,N_10070,N_10218);
nor U11265 (N_11265,N_10628,N_10951);
or U11266 (N_11266,N_10878,N_10110);
and U11267 (N_11267,N_10364,N_10756);
nor U11268 (N_11268,N_10865,N_10856);
nand U11269 (N_11269,N_10591,N_10677);
or U11270 (N_11270,N_10681,N_10605);
nor U11271 (N_11271,N_10876,N_10962);
and U11272 (N_11272,N_10039,N_10561);
nor U11273 (N_11273,N_10645,N_10947);
or U11274 (N_11274,N_10348,N_10538);
nand U11275 (N_11275,N_10191,N_10486);
and U11276 (N_11276,N_10000,N_10077);
or U11277 (N_11277,N_10514,N_10785);
nor U11278 (N_11278,N_10671,N_10873);
xor U11279 (N_11279,N_10033,N_10362);
xor U11280 (N_11280,N_10224,N_10352);
or U11281 (N_11281,N_10905,N_10404);
nor U11282 (N_11282,N_10125,N_10794);
and U11283 (N_11283,N_10237,N_10862);
or U11284 (N_11284,N_10007,N_10736);
nand U11285 (N_11285,N_10879,N_10474);
or U11286 (N_11286,N_10037,N_10512);
or U11287 (N_11287,N_10367,N_10629);
nor U11288 (N_11288,N_10208,N_10610);
or U11289 (N_11289,N_10720,N_10184);
nor U11290 (N_11290,N_10127,N_10061);
and U11291 (N_11291,N_10103,N_10568);
or U11292 (N_11292,N_10752,N_10871);
nor U11293 (N_11293,N_10665,N_10093);
or U11294 (N_11294,N_10254,N_10883);
or U11295 (N_11295,N_10192,N_10094);
nor U11296 (N_11296,N_10573,N_10901);
and U11297 (N_11297,N_10017,N_10618);
xor U11298 (N_11298,N_10164,N_10841);
nor U11299 (N_11299,N_10983,N_10600);
nor U11300 (N_11300,N_10437,N_10446);
xor U11301 (N_11301,N_10326,N_10560);
nand U11302 (N_11302,N_10770,N_10580);
nor U11303 (N_11303,N_10653,N_10958);
or U11304 (N_11304,N_10617,N_10823);
nor U11305 (N_11305,N_10758,N_10056);
xor U11306 (N_11306,N_10423,N_10190);
and U11307 (N_11307,N_10316,N_10892);
nand U11308 (N_11308,N_10357,N_10709);
and U11309 (N_11309,N_10214,N_10500);
nor U11310 (N_11310,N_10058,N_10954);
nor U11311 (N_11311,N_10976,N_10071);
or U11312 (N_11312,N_10619,N_10147);
and U11313 (N_11313,N_10700,N_10301);
xor U11314 (N_11314,N_10273,N_10918);
xor U11315 (N_11315,N_10115,N_10377);
or U11316 (N_11316,N_10952,N_10576);
or U11317 (N_11317,N_10244,N_10055);
or U11318 (N_11318,N_10340,N_10372);
and U11319 (N_11319,N_10613,N_10586);
nand U11320 (N_11320,N_10258,N_10170);
and U11321 (N_11321,N_10829,N_10941);
nand U11322 (N_11322,N_10582,N_10403);
nand U11323 (N_11323,N_10207,N_10699);
and U11324 (N_11324,N_10814,N_10193);
or U11325 (N_11325,N_10289,N_10664);
nor U11326 (N_11326,N_10759,N_10926);
nor U11327 (N_11327,N_10371,N_10179);
nor U11328 (N_11328,N_10453,N_10692);
or U11329 (N_11329,N_10036,N_10854);
and U11330 (N_11330,N_10890,N_10053);
nand U11331 (N_11331,N_10248,N_10243);
nor U11332 (N_11332,N_10074,N_10984);
nor U11333 (N_11333,N_10083,N_10661);
nor U11334 (N_11334,N_10528,N_10268);
and U11335 (N_11335,N_10535,N_10277);
nor U11336 (N_11336,N_10647,N_10724);
xnor U11337 (N_11337,N_10183,N_10527);
and U11338 (N_11338,N_10729,N_10275);
nor U11339 (N_11339,N_10886,N_10092);
and U11340 (N_11340,N_10550,N_10144);
xnor U11341 (N_11341,N_10143,N_10847);
nand U11342 (N_11342,N_10156,N_10048);
nand U11343 (N_11343,N_10363,N_10479);
nand U11344 (N_11344,N_10635,N_10167);
and U11345 (N_11345,N_10278,N_10744);
and U11346 (N_11346,N_10728,N_10579);
and U11347 (N_11347,N_10313,N_10920);
xnor U11348 (N_11348,N_10678,N_10778);
nor U11349 (N_11349,N_10537,N_10062);
nor U11350 (N_11350,N_10443,N_10426);
nor U11351 (N_11351,N_10743,N_10634);
or U11352 (N_11352,N_10667,N_10493);
nor U11353 (N_11353,N_10762,N_10010);
nor U11354 (N_11354,N_10599,N_10539);
nand U11355 (N_11355,N_10434,N_10009);
nor U11356 (N_11356,N_10861,N_10461);
or U11357 (N_11357,N_10253,N_10013);
nand U11358 (N_11358,N_10832,N_10305);
nand U11359 (N_11359,N_10195,N_10848);
nand U11360 (N_11360,N_10148,N_10857);
and U11361 (N_11361,N_10562,N_10158);
or U11362 (N_11362,N_10622,N_10896);
and U11363 (N_11363,N_10488,N_10456);
xor U11364 (N_11364,N_10157,N_10811);
and U11365 (N_11365,N_10543,N_10751);
and U11366 (N_11366,N_10291,N_10475);
nand U11367 (N_11367,N_10285,N_10373);
nand U11368 (N_11368,N_10596,N_10575);
and U11369 (N_11369,N_10302,N_10108);
nand U11370 (N_11370,N_10054,N_10152);
nand U11371 (N_11371,N_10060,N_10637);
or U11372 (N_11372,N_10402,N_10004);
nor U11373 (N_11373,N_10444,N_10640);
or U11374 (N_11374,N_10078,N_10626);
and U11375 (N_11375,N_10872,N_10124);
xor U11376 (N_11376,N_10765,N_10295);
or U11377 (N_11377,N_10532,N_10079);
or U11378 (N_11378,N_10120,N_10583);
or U11379 (N_11379,N_10096,N_10422);
nand U11380 (N_11380,N_10816,N_10712);
nor U11381 (N_11381,N_10346,N_10229);
nand U11382 (N_11382,N_10281,N_10328);
xnor U11383 (N_11383,N_10889,N_10903);
nand U11384 (N_11384,N_10498,N_10225);
or U11385 (N_11385,N_10447,N_10894);
nand U11386 (N_11386,N_10202,N_10468);
or U11387 (N_11387,N_10870,N_10646);
and U11388 (N_11388,N_10102,N_10833);
xnor U11389 (N_11389,N_10151,N_10650);
xnor U11390 (N_11390,N_10971,N_10117);
and U11391 (N_11391,N_10320,N_10676);
xor U11392 (N_11392,N_10321,N_10420);
nor U11393 (N_11393,N_10450,N_10809);
nand U11394 (N_11394,N_10654,N_10314);
and U11395 (N_11395,N_10989,N_10159);
nand U11396 (N_11396,N_10846,N_10069);
nor U11397 (N_11397,N_10376,N_10803);
nor U11398 (N_11398,N_10548,N_10503);
and U11399 (N_11399,N_10414,N_10927);
nand U11400 (N_11400,N_10045,N_10138);
nor U11401 (N_11401,N_10721,N_10084);
xor U11402 (N_11402,N_10788,N_10233);
nand U11403 (N_11403,N_10235,N_10121);
and U11404 (N_11404,N_10930,N_10908);
and U11405 (N_11405,N_10680,N_10433);
xor U11406 (N_11406,N_10349,N_10095);
nand U11407 (N_11407,N_10464,N_10463);
or U11408 (N_11408,N_10659,N_10904);
nand U11409 (N_11409,N_10725,N_10881);
nand U11410 (N_11410,N_10030,N_10922);
or U11411 (N_11411,N_10849,N_10472);
nor U11412 (N_11412,N_10696,N_10994);
xor U11413 (N_11413,N_10817,N_10043);
nand U11414 (N_11414,N_10800,N_10391);
nand U11415 (N_11415,N_10781,N_10666);
or U11416 (N_11416,N_10021,N_10978);
xor U11417 (N_11417,N_10799,N_10283);
nor U11418 (N_11418,N_10631,N_10104);
or U11419 (N_11419,N_10969,N_10140);
nand U11420 (N_11420,N_10730,N_10332);
and U11421 (N_11421,N_10701,N_10732);
nor U11422 (N_11422,N_10988,N_10748);
nand U11423 (N_11423,N_10867,N_10162);
or U11424 (N_11424,N_10410,N_10259);
nand U11425 (N_11425,N_10975,N_10001);
or U11426 (N_11426,N_10331,N_10996);
and U11427 (N_11427,N_10987,N_10802);
and U11428 (N_11428,N_10986,N_10399);
and U11429 (N_11429,N_10298,N_10716);
nand U11430 (N_11430,N_10793,N_10608);
nor U11431 (N_11431,N_10937,N_10929);
xor U11432 (N_11432,N_10786,N_10469);
or U11433 (N_11433,N_10497,N_10545);
nand U11434 (N_11434,N_10992,N_10034);
nand U11435 (N_11435,N_10831,N_10489);
or U11436 (N_11436,N_10322,N_10592);
xnor U11437 (N_11437,N_10333,N_10145);
or U11438 (N_11438,N_10338,N_10806);
nand U11439 (N_11439,N_10288,N_10923);
and U11440 (N_11440,N_10249,N_10473);
or U11441 (N_11441,N_10997,N_10891);
and U11442 (N_11442,N_10708,N_10172);
nand U11443 (N_11443,N_10089,N_10451);
nor U11444 (N_11444,N_10960,N_10068);
nand U11445 (N_11445,N_10763,N_10421);
or U11446 (N_11446,N_10703,N_10740);
and U11447 (N_11447,N_10995,N_10005);
nor U11448 (N_11448,N_10080,N_10210);
nand U11449 (N_11449,N_10590,N_10356);
nand U11450 (N_11450,N_10220,N_10425);
nor U11451 (N_11451,N_10150,N_10204);
nand U11452 (N_11452,N_10400,N_10893);
xnor U11453 (N_11453,N_10974,N_10837);
nand U11454 (N_11454,N_10114,N_10792);
and U11455 (N_11455,N_10601,N_10276);
and U11456 (N_11456,N_10649,N_10609);
and U11457 (N_11457,N_10607,N_10557);
nand U11458 (N_11458,N_10769,N_10625);
nand U11459 (N_11459,N_10633,N_10564);
and U11460 (N_11460,N_10949,N_10509);
xor U11461 (N_11461,N_10211,N_10455);
and U11462 (N_11462,N_10265,N_10955);
and U11463 (N_11463,N_10132,N_10141);
nand U11464 (N_11464,N_10256,N_10394);
and U11465 (N_11465,N_10513,N_10715);
nor U11466 (N_11466,N_10401,N_10820);
nand U11467 (N_11467,N_10266,N_10206);
or U11468 (N_11468,N_10015,N_10380);
nand U11469 (N_11469,N_10029,N_10655);
nand U11470 (N_11470,N_10073,N_10611);
and U11471 (N_11471,N_10169,N_10165);
or U11472 (N_11472,N_10899,N_10998);
nor U11473 (N_11473,N_10405,N_10123);
xor U11474 (N_11474,N_10119,N_10555);
xnor U11475 (N_11475,N_10597,N_10136);
nand U11476 (N_11476,N_10885,N_10587);
nand U11477 (N_11477,N_10795,N_10542);
nand U11478 (N_11478,N_10100,N_10515);
nand U11479 (N_11479,N_10319,N_10052);
xor U11480 (N_11480,N_10719,N_10544);
nand U11481 (N_11481,N_10257,N_10801);
and U11482 (N_11482,N_10578,N_10789);
xnor U11483 (N_11483,N_10023,N_10508);
xor U11484 (N_11484,N_10267,N_10913);
and U11485 (N_11485,N_10499,N_10615);
or U11486 (N_11486,N_10694,N_10621);
nor U11487 (N_11487,N_10636,N_10086);
and U11488 (N_11488,N_10723,N_10250);
or U11489 (N_11489,N_10466,N_10378);
nor U11490 (N_11490,N_10639,N_10651);
and U11491 (N_11491,N_10435,N_10230);
and U11492 (N_11492,N_10552,N_10097);
and U11493 (N_11493,N_10830,N_10934);
nor U11494 (N_11494,N_10025,N_10776);
nand U11495 (N_11495,N_10274,N_10171);
xor U11496 (N_11496,N_10284,N_10864);
or U11497 (N_11497,N_10112,N_10063);
and U11498 (N_11498,N_10919,N_10773);
or U11499 (N_11499,N_10355,N_10228);
and U11500 (N_11500,N_10423,N_10755);
nor U11501 (N_11501,N_10880,N_10639);
and U11502 (N_11502,N_10574,N_10351);
nand U11503 (N_11503,N_10099,N_10421);
and U11504 (N_11504,N_10706,N_10830);
nor U11505 (N_11505,N_10671,N_10425);
or U11506 (N_11506,N_10750,N_10803);
nor U11507 (N_11507,N_10863,N_10999);
nor U11508 (N_11508,N_10574,N_10522);
or U11509 (N_11509,N_10631,N_10124);
or U11510 (N_11510,N_10510,N_10680);
nand U11511 (N_11511,N_10491,N_10292);
or U11512 (N_11512,N_10675,N_10207);
nand U11513 (N_11513,N_10664,N_10954);
and U11514 (N_11514,N_10830,N_10397);
or U11515 (N_11515,N_10622,N_10972);
nor U11516 (N_11516,N_10286,N_10887);
or U11517 (N_11517,N_10457,N_10430);
xor U11518 (N_11518,N_10898,N_10542);
nand U11519 (N_11519,N_10755,N_10483);
or U11520 (N_11520,N_10395,N_10818);
and U11521 (N_11521,N_10742,N_10427);
or U11522 (N_11522,N_10099,N_10461);
nor U11523 (N_11523,N_10754,N_10524);
xor U11524 (N_11524,N_10836,N_10940);
xnor U11525 (N_11525,N_10017,N_10811);
nor U11526 (N_11526,N_10729,N_10443);
and U11527 (N_11527,N_10536,N_10535);
and U11528 (N_11528,N_10313,N_10316);
nand U11529 (N_11529,N_10262,N_10459);
nor U11530 (N_11530,N_10312,N_10664);
nand U11531 (N_11531,N_10095,N_10955);
nand U11532 (N_11532,N_10073,N_10647);
and U11533 (N_11533,N_10214,N_10022);
and U11534 (N_11534,N_10644,N_10471);
and U11535 (N_11535,N_10310,N_10017);
and U11536 (N_11536,N_10348,N_10059);
and U11537 (N_11537,N_10074,N_10365);
or U11538 (N_11538,N_10935,N_10487);
nor U11539 (N_11539,N_10741,N_10098);
or U11540 (N_11540,N_10171,N_10954);
nand U11541 (N_11541,N_10773,N_10627);
and U11542 (N_11542,N_10016,N_10172);
and U11543 (N_11543,N_10154,N_10380);
and U11544 (N_11544,N_10761,N_10057);
or U11545 (N_11545,N_10841,N_10851);
nand U11546 (N_11546,N_10925,N_10250);
xnor U11547 (N_11547,N_10992,N_10216);
nor U11548 (N_11548,N_10328,N_10683);
and U11549 (N_11549,N_10144,N_10055);
xor U11550 (N_11550,N_10606,N_10292);
xnor U11551 (N_11551,N_10444,N_10903);
nand U11552 (N_11552,N_10539,N_10538);
or U11553 (N_11553,N_10033,N_10804);
nor U11554 (N_11554,N_10356,N_10850);
or U11555 (N_11555,N_10627,N_10780);
and U11556 (N_11556,N_10744,N_10054);
nand U11557 (N_11557,N_10258,N_10213);
nor U11558 (N_11558,N_10243,N_10506);
or U11559 (N_11559,N_10482,N_10035);
nand U11560 (N_11560,N_10927,N_10581);
nand U11561 (N_11561,N_10587,N_10651);
nand U11562 (N_11562,N_10644,N_10626);
and U11563 (N_11563,N_10472,N_10166);
and U11564 (N_11564,N_10625,N_10708);
nand U11565 (N_11565,N_10310,N_10907);
nand U11566 (N_11566,N_10143,N_10275);
and U11567 (N_11567,N_10745,N_10274);
nor U11568 (N_11568,N_10687,N_10942);
nor U11569 (N_11569,N_10443,N_10928);
nor U11570 (N_11570,N_10323,N_10300);
nand U11571 (N_11571,N_10999,N_10490);
nor U11572 (N_11572,N_10654,N_10853);
and U11573 (N_11573,N_10647,N_10324);
and U11574 (N_11574,N_10233,N_10815);
nor U11575 (N_11575,N_10920,N_10517);
xor U11576 (N_11576,N_10361,N_10735);
or U11577 (N_11577,N_10757,N_10612);
xnor U11578 (N_11578,N_10201,N_10125);
nand U11579 (N_11579,N_10178,N_10415);
nor U11580 (N_11580,N_10070,N_10362);
or U11581 (N_11581,N_10555,N_10416);
nand U11582 (N_11582,N_10186,N_10419);
and U11583 (N_11583,N_10691,N_10740);
and U11584 (N_11584,N_10561,N_10237);
or U11585 (N_11585,N_10578,N_10281);
xor U11586 (N_11586,N_10706,N_10897);
and U11587 (N_11587,N_10543,N_10252);
nor U11588 (N_11588,N_10376,N_10114);
nor U11589 (N_11589,N_10470,N_10953);
or U11590 (N_11590,N_10466,N_10815);
nand U11591 (N_11591,N_10310,N_10854);
nand U11592 (N_11592,N_10726,N_10717);
or U11593 (N_11593,N_10723,N_10789);
and U11594 (N_11594,N_10627,N_10741);
nor U11595 (N_11595,N_10112,N_10886);
nand U11596 (N_11596,N_10142,N_10694);
xor U11597 (N_11597,N_10235,N_10880);
nand U11598 (N_11598,N_10108,N_10092);
and U11599 (N_11599,N_10178,N_10132);
and U11600 (N_11600,N_10548,N_10099);
or U11601 (N_11601,N_10893,N_10742);
nand U11602 (N_11602,N_10248,N_10705);
nand U11603 (N_11603,N_10848,N_10045);
and U11604 (N_11604,N_10975,N_10854);
nand U11605 (N_11605,N_10349,N_10864);
nand U11606 (N_11606,N_10807,N_10403);
and U11607 (N_11607,N_10531,N_10825);
and U11608 (N_11608,N_10061,N_10896);
nor U11609 (N_11609,N_10718,N_10144);
nand U11610 (N_11610,N_10295,N_10539);
nand U11611 (N_11611,N_10837,N_10242);
nand U11612 (N_11612,N_10595,N_10311);
xor U11613 (N_11613,N_10423,N_10416);
nand U11614 (N_11614,N_10376,N_10195);
nor U11615 (N_11615,N_10729,N_10422);
nand U11616 (N_11616,N_10406,N_10668);
nand U11617 (N_11617,N_10737,N_10808);
nand U11618 (N_11618,N_10006,N_10067);
or U11619 (N_11619,N_10866,N_10248);
and U11620 (N_11620,N_10726,N_10462);
nor U11621 (N_11621,N_10906,N_10483);
and U11622 (N_11622,N_10840,N_10987);
and U11623 (N_11623,N_10311,N_10972);
or U11624 (N_11624,N_10725,N_10006);
nand U11625 (N_11625,N_10995,N_10598);
or U11626 (N_11626,N_10891,N_10905);
or U11627 (N_11627,N_10141,N_10470);
or U11628 (N_11628,N_10230,N_10366);
or U11629 (N_11629,N_10817,N_10821);
nor U11630 (N_11630,N_10103,N_10724);
nor U11631 (N_11631,N_10996,N_10385);
and U11632 (N_11632,N_10527,N_10950);
xnor U11633 (N_11633,N_10166,N_10319);
xnor U11634 (N_11634,N_10362,N_10824);
and U11635 (N_11635,N_10779,N_10081);
xnor U11636 (N_11636,N_10105,N_10395);
and U11637 (N_11637,N_10250,N_10556);
nand U11638 (N_11638,N_10589,N_10964);
nor U11639 (N_11639,N_10904,N_10532);
nand U11640 (N_11640,N_10487,N_10035);
xnor U11641 (N_11641,N_10487,N_10791);
and U11642 (N_11642,N_10379,N_10839);
and U11643 (N_11643,N_10685,N_10332);
and U11644 (N_11644,N_10681,N_10994);
nor U11645 (N_11645,N_10278,N_10445);
nand U11646 (N_11646,N_10451,N_10540);
and U11647 (N_11647,N_10901,N_10980);
or U11648 (N_11648,N_10057,N_10530);
nor U11649 (N_11649,N_10000,N_10621);
and U11650 (N_11650,N_10922,N_10449);
nor U11651 (N_11651,N_10466,N_10593);
or U11652 (N_11652,N_10771,N_10388);
or U11653 (N_11653,N_10328,N_10906);
nand U11654 (N_11654,N_10680,N_10665);
nor U11655 (N_11655,N_10581,N_10393);
nand U11656 (N_11656,N_10868,N_10730);
and U11657 (N_11657,N_10957,N_10553);
and U11658 (N_11658,N_10668,N_10524);
nand U11659 (N_11659,N_10562,N_10186);
and U11660 (N_11660,N_10235,N_10558);
nand U11661 (N_11661,N_10376,N_10805);
nand U11662 (N_11662,N_10899,N_10486);
nand U11663 (N_11663,N_10429,N_10233);
and U11664 (N_11664,N_10897,N_10508);
nand U11665 (N_11665,N_10942,N_10800);
nand U11666 (N_11666,N_10429,N_10633);
xor U11667 (N_11667,N_10542,N_10384);
or U11668 (N_11668,N_10645,N_10567);
nand U11669 (N_11669,N_10837,N_10570);
nor U11670 (N_11670,N_10873,N_10060);
nand U11671 (N_11671,N_10008,N_10411);
xnor U11672 (N_11672,N_10181,N_10118);
nand U11673 (N_11673,N_10712,N_10860);
nand U11674 (N_11674,N_10764,N_10813);
nor U11675 (N_11675,N_10426,N_10378);
nand U11676 (N_11676,N_10339,N_10712);
and U11677 (N_11677,N_10329,N_10320);
nand U11678 (N_11678,N_10958,N_10472);
xor U11679 (N_11679,N_10817,N_10249);
nand U11680 (N_11680,N_10221,N_10053);
or U11681 (N_11681,N_10300,N_10011);
and U11682 (N_11682,N_10831,N_10625);
and U11683 (N_11683,N_10686,N_10254);
nand U11684 (N_11684,N_10967,N_10179);
and U11685 (N_11685,N_10527,N_10126);
nor U11686 (N_11686,N_10760,N_10202);
xor U11687 (N_11687,N_10413,N_10927);
nor U11688 (N_11688,N_10981,N_10713);
nand U11689 (N_11689,N_10778,N_10560);
nor U11690 (N_11690,N_10848,N_10473);
and U11691 (N_11691,N_10418,N_10317);
xnor U11692 (N_11692,N_10614,N_10958);
and U11693 (N_11693,N_10306,N_10340);
or U11694 (N_11694,N_10536,N_10546);
nor U11695 (N_11695,N_10342,N_10870);
nand U11696 (N_11696,N_10865,N_10738);
and U11697 (N_11697,N_10798,N_10695);
or U11698 (N_11698,N_10406,N_10153);
nand U11699 (N_11699,N_10770,N_10164);
nor U11700 (N_11700,N_10595,N_10181);
nor U11701 (N_11701,N_10876,N_10956);
nand U11702 (N_11702,N_10187,N_10238);
or U11703 (N_11703,N_10722,N_10062);
or U11704 (N_11704,N_10396,N_10883);
or U11705 (N_11705,N_10948,N_10692);
and U11706 (N_11706,N_10679,N_10240);
nand U11707 (N_11707,N_10384,N_10355);
nor U11708 (N_11708,N_10264,N_10809);
xor U11709 (N_11709,N_10311,N_10689);
and U11710 (N_11710,N_10902,N_10533);
xor U11711 (N_11711,N_10084,N_10458);
and U11712 (N_11712,N_10350,N_10757);
or U11713 (N_11713,N_10198,N_10160);
or U11714 (N_11714,N_10796,N_10732);
nor U11715 (N_11715,N_10599,N_10304);
and U11716 (N_11716,N_10976,N_10740);
xnor U11717 (N_11717,N_10715,N_10771);
or U11718 (N_11718,N_10686,N_10197);
and U11719 (N_11719,N_10961,N_10058);
and U11720 (N_11720,N_10917,N_10101);
xor U11721 (N_11721,N_10316,N_10053);
or U11722 (N_11722,N_10239,N_10692);
or U11723 (N_11723,N_10721,N_10975);
nor U11724 (N_11724,N_10432,N_10039);
nor U11725 (N_11725,N_10858,N_10049);
nor U11726 (N_11726,N_10626,N_10109);
xnor U11727 (N_11727,N_10104,N_10571);
xnor U11728 (N_11728,N_10946,N_10857);
and U11729 (N_11729,N_10196,N_10006);
nor U11730 (N_11730,N_10485,N_10810);
nand U11731 (N_11731,N_10253,N_10961);
or U11732 (N_11732,N_10979,N_10375);
and U11733 (N_11733,N_10431,N_10674);
and U11734 (N_11734,N_10588,N_10371);
nor U11735 (N_11735,N_10305,N_10970);
or U11736 (N_11736,N_10443,N_10149);
nor U11737 (N_11737,N_10828,N_10379);
or U11738 (N_11738,N_10331,N_10007);
nand U11739 (N_11739,N_10520,N_10553);
and U11740 (N_11740,N_10598,N_10606);
or U11741 (N_11741,N_10020,N_10446);
or U11742 (N_11742,N_10199,N_10991);
and U11743 (N_11743,N_10109,N_10547);
or U11744 (N_11744,N_10215,N_10075);
nor U11745 (N_11745,N_10118,N_10981);
nor U11746 (N_11746,N_10359,N_10197);
and U11747 (N_11747,N_10994,N_10930);
xor U11748 (N_11748,N_10170,N_10495);
nor U11749 (N_11749,N_10603,N_10055);
nand U11750 (N_11750,N_10042,N_10715);
nand U11751 (N_11751,N_10531,N_10485);
xor U11752 (N_11752,N_10775,N_10697);
nand U11753 (N_11753,N_10658,N_10180);
and U11754 (N_11754,N_10883,N_10214);
nand U11755 (N_11755,N_10157,N_10215);
and U11756 (N_11756,N_10651,N_10314);
xor U11757 (N_11757,N_10287,N_10057);
nor U11758 (N_11758,N_10182,N_10763);
nor U11759 (N_11759,N_10078,N_10143);
and U11760 (N_11760,N_10600,N_10745);
or U11761 (N_11761,N_10374,N_10944);
nand U11762 (N_11762,N_10347,N_10438);
and U11763 (N_11763,N_10073,N_10461);
and U11764 (N_11764,N_10598,N_10760);
and U11765 (N_11765,N_10775,N_10291);
nand U11766 (N_11766,N_10313,N_10468);
nand U11767 (N_11767,N_10044,N_10342);
nor U11768 (N_11768,N_10231,N_10220);
nor U11769 (N_11769,N_10154,N_10697);
and U11770 (N_11770,N_10423,N_10318);
nor U11771 (N_11771,N_10229,N_10055);
xor U11772 (N_11772,N_10221,N_10880);
or U11773 (N_11773,N_10623,N_10195);
and U11774 (N_11774,N_10758,N_10587);
or U11775 (N_11775,N_10840,N_10266);
xor U11776 (N_11776,N_10171,N_10726);
and U11777 (N_11777,N_10923,N_10859);
xor U11778 (N_11778,N_10694,N_10297);
or U11779 (N_11779,N_10208,N_10500);
xnor U11780 (N_11780,N_10723,N_10037);
and U11781 (N_11781,N_10133,N_10517);
xnor U11782 (N_11782,N_10070,N_10598);
nand U11783 (N_11783,N_10415,N_10065);
nor U11784 (N_11784,N_10650,N_10689);
xor U11785 (N_11785,N_10473,N_10494);
or U11786 (N_11786,N_10908,N_10457);
nand U11787 (N_11787,N_10309,N_10111);
nor U11788 (N_11788,N_10854,N_10453);
nand U11789 (N_11789,N_10801,N_10100);
nand U11790 (N_11790,N_10870,N_10274);
and U11791 (N_11791,N_10758,N_10299);
or U11792 (N_11792,N_10025,N_10136);
nand U11793 (N_11793,N_10718,N_10896);
xor U11794 (N_11794,N_10096,N_10498);
or U11795 (N_11795,N_10689,N_10699);
nor U11796 (N_11796,N_10469,N_10100);
nor U11797 (N_11797,N_10074,N_10644);
nor U11798 (N_11798,N_10035,N_10811);
nand U11799 (N_11799,N_10339,N_10959);
nand U11800 (N_11800,N_10073,N_10510);
nor U11801 (N_11801,N_10168,N_10578);
or U11802 (N_11802,N_10884,N_10015);
nor U11803 (N_11803,N_10799,N_10576);
nor U11804 (N_11804,N_10883,N_10167);
nor U11805 (N_11805,N_10124,N_10675);
xnor U11806 (N_11806,N_10543,N_10995);
or U11807 (N_11807,N_10855,N_10890);
nor U11808 (N_11808,N_10715,N_10329);
and U11809 (N_11809,N_10585,N_10206);
or U11810 (N_11810,N_10957,N_10803);
and U11811 (N_11811,N_10989,N_10126);
nand U11812 (N_11812,N_10361,N_10850);
nor U11813 (N_11813,N_10189,N_10982);
nor U11814 (N_11814,N_10013,N_10164);
and U11815 (N_11815,N_10819,N_10066);
xor U11816 (N_11816,N_10567,N_10443);
nand U11817 (N_11817,N_10601,N_10068);
nand U11818 (N_11818,N_10649,N_10767);
nand U11819 (N_11819,N_10709,N_10315);
xor U11820 (N_11820,N_10213,N_10399);
and U11821 (N_11821,N_10931,N_10550);
xor U11822 (N_11822,N_10414,N_10539);
or U11823 (N_11823,N_10363,N_10984);
and U11824 (N_11824,N_10973,N_10026);
and U11825 (N_11825,N_10606,N_10424);
nand U11826 (N_11826,N_10201,N_10231);
nor U11827 (N_11827,N_10557,N_10406);
nand U11828 (N_11828,N_10204,N_10425);
xnor U11829 (N_11829,N_10174,N_10350);
xnor U11830 (N_11830,N_10565,N_10348);
and U11831 (N_11831,N_10264,N_10042);
nand U11832 (N_11832,N_10668,N_10007);
nor U11833 (N_11833,N_10797,N_10961);
and U11834 (N_11834,N_10761,N_10836);
and U11835 (N_11835,N_10004,N_10745);
and U11836 (N_11836,N_10070,N_10379);
and U11837 (N_11837,N_10108,N_10261);
nor U11838 (N_11838,N_10613,N_10571);
and U11839 (N_11839,N_10548,N_10328);
or U11840 (N_11840,N_10450,N_10631);
and U11841 (N_11841,N_10416,N_10916);
nand U11842 (N_11842,N_10815,N_10281);
nor U11843 (N_11843,N_10268,N_10237);
or U11844 (N_11844,N_10155,N_10740);
nor U11845 (N_11845,N_10947,N_10007);
nor U11846 (N_11846,N_10951,N_10347);
or U11847 (N_11847,N_10343,N_10707);
xor U11848 (N_11848,N_10005,N_10206);
nor U11849 (N_11849,N_10362,N_10344);
or U11850 (N_11850,N_10346,N_10480);
or U11851 (N_11851,N_10548,N_10403);
and U11852 (N_11852,N_10405,N_10853);
or U11853 (N_11853,N_10792,N_10404);
or U11854 (N_11854,N_10771,N_10628);
nand U11855 (N_11855,N_10861,N_10662);
nor U11856 (N_11856,N_10634,N_10872);
nor U11857 (N_11857,N_10738,N_10227);
or U11858 (N_11858,N_10744,N_10232);
and U11859 (N_11859,N_10918,N_10338);
and U11860 (N_11860,N_10804,N_10843);
and U11861 (N_11861,N_10893,N_10203);
nand U11862 (N_11862,N_10128,N_10748);
and U11863 (N_11863,N_10236,N_10513);
or U11864 (N_11864,N_10209,N_10973);
nor U11865 (N_11865,N_10300,N_10478);
nand U11866 (N_11866,N_10938,N_10771);
nor U11867 (N_11867,N_10229,N_10279);
and U11868 (N_11868,N_10505,N_10623);
xor U11869 (N_11869,N_10380,N_10832);
nor U11870 (N_11870,N_10729,N_10845);
xor U11871 (N_11871,N_10988,N_10158);
nand U11872 (N_11872,N_10582,N_10103);
or U11873 (N_11873,N_10767,N_10598);
nor U11874 (N_11874,N_10047,N_10584);
nand U11875 (N_11875,N_10802,N_10953);
nor U11876 (N_11876,N_10797,N_10578);
nand U11877 (N_11877,N_10212,N_10279);
xor U11878 (N_11878,N_10499,N_10272);
nand U11879 (N_11879,N_10777,N_10049);
and U11880 (N_11880,N_10793,N_10972);
and U11881 (N_11881,N_10921,N_10243);
and U11882 (N_11882,N_10691,N_10412);
nand U11883 (N_11883,N_10148,N_10412);
xnor U11884 (N_11884,N_10313,N_10259);
nor U11885 (N_11885,N_10858,N_10790);
or U11886 (N_11886,N_10625,N_10402);
nor U11887 (N_11887,N_10896,N_10060);
or U11888 (N_11888,N_10054,N_10121);
and U11889 (N_11889,N_10891,N_10099);
and U11890 (N_11890,N_10147,N_10450);
nor U11891 (N_11891,N_10311,N_10498);
or U11892 (N_11892,N_10171,N_10767);
xnor U11893 (N_11893,N_10939,N_10181);
and U11894 (N_11894,N_10490,N_10334);
and U11895 (N_11895,N_10144,N_10360);
nand U11896 (N_11896,N_10531,N_10250);
nand U11897 (N_11897,N_10179,N_10562);
nand U11898 (N_11898,N_10761,N_10672);
and U11899 (N_11899,N_10440,N_10893);
and U11900 (N_11900,N_10091,N_10118);
nor U11901 (N_11901,N_10356,N_10602);
nand U11902 (N_11902,N_10351,N_10582);
and U11903 (N_11903,N_10360,N_10886);
nand U11904 (N_11904,N_10000,N_10196);
nand U11905 (N_11905,N_10162,N_10539);
or U11906 (N_11906,N_10587,N_10865);
and U11907 (N_11907,N_10506,N_10397);
and U11908 (N_11908,N_10823,N_10211);
and U11909 (N_11909,N_10841,N_10527);
and U11910 (N_11910,N_10435,N_10538);
or U11911 (N_11911,N_10649,N_10732);
and U11912 (N_11912,N_10373,N_10915);
nand U11913 (N_11913,N_10313,N_10229);
and U11914 (N_11914,N_10975,N_10882);
or U11915 (N_11915,N_10622,N_10950);
or U11916 (N_11916,N_10623,N_10577);
xnor U11917 (N_11917,N_10669,N_10907);
nand U11918 (N_11918,N_10022,N_10312);
nor U11919 (N_11919,N_10083,N_10185);
nor U11920 (N_11920,N_10939,N_10599);
nand U11921 (N_11921,N_10647,N_10148);
xnor U11922 (N_11922,N_10575,N_10188);
nand U11923 (N_11923,N_10336,N_10775);
xnor U11924 (N_11924,N_10885,N_10065);
xnor U11925 (N_11925,N_10510,N_10675);
nor U11926 (N_11926,N_10470,N_10264);
nand U11927 (N_11927,N_10558,N_10031);
nand U11928 (N_11928,N_10270,N_10417);
xor U11929 (N_11929,N_10425,N_10991);
and U11930 (N_11930,N_10302,N_10801);
or U11931 (N_11931,N_10322,N_10188);
or U11932 (N_11932,N_10834,N_10029);
or U11933 (N_11933,N_10274,N_10851);
or U11934 (N_11934,N_10324,N_10300);
or U11935 (N_11935,N_10345,N_10318);
and U11936 (N_11936,N_10488,N_10965);
or U11937 (N_11937,N_10173,N_10161);
nand U11938 (N_11938,N_10322,N_10562);
nor U11939 (N_11939,N_10930,N_10890);
xnor U11940 (N_11940,N_10656,N_10947);
nor U11941 (N_11941,N_10404,N_10628);
and U11942 (N_11942,N_10230,N_10599);
nand U11943 (N_11943,N_10748,N_10023);
or U11944 (N_11944,N_10480,N_10409);
nor U11945 (N_11945,N_10024,N_10997);
nor U11946 (N_11946,N_10227,N_10306);
xor U11947 (N_11947,N_10882,N_10358);
xnor U11948 (N_11948,N_10745,N_10684);
or U11949 (N_11949,N_10849,N_10317);
nor U11950 (N_11950,N_10251,N_10157);
nor U11951 (N_11951,N_10470,N_10895);
nor U11952 (N_11952,N_10171,N_10836);
nand U11953 (N_11953,N_10736,N_10671);
nor U11954 (N_11954,N_10411,N_10271);
nand U11955 (N_11955,N_10227,N_10534);
and U11956 (N_11956,N_10727,N_10225);
nor U11957 (N_11957,N_10581,N_10786);
and U11958 (N_11958,N_10983,N_10528);
and U11959 (N_11959,N_10441,N_10299);
nand U11960 (N_11960,N_10372,N_10400);
xor U11961 (N_11961,N_10147,N_10036);
and U11962 (N_11962,N_10650,N_10242);
and U11963 (N_11963,N_10604,N_10831);
nand U11964 (N_11964,N_10244,N_10425);
or U11965 (N_11965,N_10160,N_10035);
nor U11966 (N_11966,N_10965,N_10348);
nor U11967 (N_11967,N_10481,N_10269);
or U11968 (N_11968,N_10104,N_10211);
and U11969 (N_11969,N_10866,N_10284);
nor U11970 (N_11970,N_10934,N_10273);
nor U11971 (N_11971,N_10466,N_10631);
or U11972 (N_11972,N_10842,N_10697);
nand U11973 (N_11973,N_10720,N_10264);
or U11974 (N_11974,N_10803,N_10392);
and U11975 (N_11975,N_10491,N_10755);
nand U11976 (N_11976,N_10953,N_10678);
and U11977 (N_11977,N_10734,N_10971);
or U11978 (N_11978,N_10940,N_10674);
nand U11979 (N_11979,N_10055,N_10931);
nor U11980 (N_11980,N_10574,N_10874);
and U11981 (N_11981,N_10999,N_10829);
or U11982 (N_11982,N_10364,N_10551);
or U11983 (N_11983,N_10079,N_10796);
nand U11984 (N_11984,N_10688,N_10115);
or U11985 (N_11985,N_10979,N_10569);
nand U11986 (N_11986,N_10938,N_10265);
nand U11987 (N_11987,N_10346,N_10762);
xor U11988 (N_11988,N_10826,N_10121);
nand U11989 (N_11989,N_10411,N_10323);
nand U11990 (N_11990,N_10179,N_10747);
and U11991 (N_11991,N_10884,N_10043);
nor U11992 (N_11992,N_10120,N_10476);
nor U11993 (N_11993,N_10619,N_10793);
or U11994 (N_11994,N_10532,N_10461);
nor U11995 (N_11995,N_10991,N_10158);
or U11996 (N_11996,N_10998,N_10494);
nor U11997 (N_11997,N_10945,N_10836);
and U11998 (N_11998,N_10525,N_10823);
or U11999 (N_11999,N_10889,N_10039);
xor U12000 (N_12000,N_11757,N_11383);
nor U12001 (N_12001,N_11909,N_11474);
xnor U12002 (N_12002,N_11290,N_11895);
or U12003 (N_12003,N_11178,N_11982);
xnor U12004 (N_12004,N_11174,N_11994);
xnor U12005 (N_12005,N_11812,N_11544);
and U12006 (N_12006,N_11580,N_11542);
nor U12007 (N_12007,N_11855,N_11839);
nor U12008 (N_12008,N_11509,N_11700);
nand U12009 (N_12009,N_11936,N_11680);
nor U12010 (N_12010,N_11167,N_11521);
or U12011 (N_12011,N_11473,N_11179);
or U12012 (N_12012,N_11803,N_11486);
xor U12013 (N_12013,N_11183,N_11977);
nand U12014 (N_12014,N_11616,N_11748);
nor U12015 (N_12015,N_11975,N_11300);
or U12016 (N_12016,N_11349,N_11976);
or U12017 (N_12017,N_11273,N_11711);
or U12018 (N_12018,N_11854,N_11328);
nor U12019 (N_12019,N_11076,N_11106);
nand U12020 (N_12020,N_11518,N_11279);
or U12021 (N_12021,N_11283,N_11872);
nand U12022 (N_12022,N_11114,N_11520);
nand U12023 (N_12023,N_11718,N_11494);
and U12024 (N_12024,N_11479,N_11480);
nor U12025 (N_12025,N_11564,N_11928);
and U12026 (N_12026,N_11029,N_11066);
or U12027 (N_12027,N_11438,N_11829);
or U12028 (N_12028,N_11792,N_11350);
or U12029 (N_12029,N_11362,N_11697);
and U12030 (N_12030,N_11151,N_11651);
or U12031 (N_12031,N_11033,N_11756);
nor U12032 (N_12032,N_11160,N_11950);
nor U12033 (N_12033,N_11638,N_11239);
or U12034 (N_12034,N_11660,N_11456);
and U12035 (N_12035,N_11560,N_11182);
nor U12036 (N_12036,N_11082,N_11095);
and U12037 (N_12037,N_11240,N_11497);
nor U12038 (N_12038,N_11437,N_11387);
or U12039 (N_12039,N_11695,N_11775);
or U12040 (N_12040,N_11003,N_11997);
or U12041 (N_12041,N_11611,N_11738);
and U12042 (N_12042,N_11750,N_11529);
nor U12043 (N_12043,N_11644,N_11837);
and U12044 (N_12044,N_11511,N_11315);
nor U12045 (N_12045,N_11797,N_11249);
and U12046 (N_12046,N_11716,N_11866);
nor U12047 (N_12047,N_11523,N_11094);
nand U12048 (N_12048,N_11203,N_11000);
or U12049 (N_12049,N_11134,N_11039);
nand U12050 (N_12050,N_11730,N_11578);
nand U12051 (N_12051,N_11368,N_11219);
and U12052 (N_12052,N_11342,N_11831);
nand U12053 (N_12053,N_11296,N_11954);
xnor U12054 (N_12054,N_11843,N_11195);
or U12055 (N_12055,N_11963,N_11250);
or U12056 (N_12056,N_11351,N_11031);
and U12057 (N_12057,N_11679,N_11386);
xnor U12058 (N_12058,N_11927,N_11026);
and U12059 (N_12059,N_11432,N_11339);
xnor U12060 (N_12060,N_11510,N_11728);
nand U12061 (N_12061,N_11876,N_11883);
nand U12062 (N_12062,N_11955,N_11708);
or U12063 (N_12063,N_11276,N_11689);
xnor U12064 (N_12064,N_11614,N_11329);
or U12065 (N_12065,N_11070,N_11487);
nor U12066 (N_12066,N_11304,N_11281);
and U12067 (N_12067,N_11528,N_11454);
or U12068 (N_12068,N_11779,N_11020);
or U12069 (N_12069,N_11147,N_11069);
nor U12070 (N_12070,N_11036,N_11531);
and U12071 (N_12071,N_11923,N_11533);
nor U12072 (N_12072,N_11972,N_11613);
or U12073 (N_12073,N_11159,N_11749);
xor U12074 (N_12074,N_11628,N_11598);
nor U12075 (N_12075,N_11277,N_11018);
and U12076 (N_12076,N_11796,N_11785);
or U12077 (N_12077,N_11085,N_11187);
nand U12078 (N_12078,N_11394,N_11781);
nor U12079 (N_12079,N_11687,N_11435);
and U12080 (N_12080,N_11222,N_11924);
and U12081 (N_12081,N_11333,N_11693);
and U12082 (N_12082,N_11419,N_11422);
and U12083 (N_12083,N_11633,N_11403);
nand U12084 (N_12084,N_11482,N_11395);
nor U12085 (N_12085,N_11554,N_11519);
or U12086 (N_12086,N_11625,N_11801);
nor U12087 (N_12087,N_11525,N_11710);
and U12088 (N_12088,N_11545,N_11649);
and U12089 (N_12089,N_11115,N_11794);
xor U12090 (N_12090,N_11524,N_11946);
and U12091 (N_12091,N_11251,N_11213);
or U12092 (N_12092,N_11062,N_11526);
or U12093 (N_12093,N_11705,N_11264);
or U12094 (N_12094,N_11814,N_11285);
or U12095 (N_12095,N_11173,N_11739);
and U12096 (N_12096,N_11925,N_11464);
and U12097 (N_12097,N_11458,N_11894);
or U12098 (N_12098,N_11821,N_11744);
nand U12099 (N_12099,N_11849,N_11120);
and U12100 (N_12100,N_11840,N_11408);
or U12101 (N_12101,N_11303,N_11742);
or U12102 (N_12102,N_11153,N_11323);
or U12103 (N_12103,N_11248,N_11216);
nor U12104 (N_12104,N_11162,N_11713);
and U12105 (N_12105,N_11129,N_11081);
and U12106 (N_12106,N_11788,N_11846);
and U12107 (N_12107,N_11990,N_11951);
or U12108 (N_12108,N_11973,N_11851);
xor U12109 (N_12109,N_11428,N_11916);
nand U12110 (N_12110,N_11127,N_11933);
and U12111 (N_12111,N_11067,N_11468);
nand U12112 (N_12112,N_11648,N_11238);
nand U12113 (N_12113,N_11343,N_11253);
or U12114 (N_12114,N_11671,N_11455);
nor U12115 (N_12115,N_11318,N_11833);
nor U12116 (N_12116,N_11536,N_11993);
xnor U12117 (N_12117,N_11449,N_11217);
nand U12118 (N_12118,N_11199,N_11181);
or U12119 (N_12119,N_11409,N_11360);
xnor U12120 (N_12120,N_11604,N_11286);
or U12121 (N_12121,N_11476,N_11607);
nand U12122 (N_12122,N_11722,N_11899);
or U12123 (N_12123,N_11763,N_11411);
xnor U12124 (N_12124,N_11672,N_11758);
or U12125 (N_12125,N_11201,N_11615);
nor U12126 (N_12126,N_11381,N_11211);
and U12127 (N_12127,N_11190,N_11887);
nor U12128 (N_12128,N_11294,N_11566);
nor U12129 (N_12129,N_11818,N_11208);
or U12130 (N_12130,N_11046,N_11502);
and U12131 (N_12131,N_11668,N_11112);
nand U12132 (N_12132,N_11929,N_11767);
nor U12133 (N_12133,N_11652,N_11466);
or U12134 (N_12134,N_11297,N_11926);
nor U12135 (N_12135,N_11786,N_11433);
or U12136 (N_12136,N_11275,N_11072);
nand U12137 (N_12137,N_11484,N_11049);
nand U12138 (N_12138,N_11724,N_11460);
or U12139 (N_12139,N_11501,N_11641);
or U12140 (N_12140,N_11327,N_11084);
xnor U12141 (N_12141,N_11577,N_11356);
or U12142 (N_12142,N_11569,N_11867);
and U12143 (N_12143,N_11585,N_11517);
or U12144 (N_12144,N_11077,N_11252);
nand U12145 (N_12145,N_11042,N_11374);
nand U12146 (N_12146,N_11143,N_11690);
nand U12147 (N_12147,N_11734,N_11787);
or U12148 (N_12148,N_11881,N_11389);
or U12149 (N_12149,N_11500,N_11844);
nand U12150 (N_12150,N_11175,N_11490);
or U12151 (N_12151,N_11956,N_11747);
and U12152 (N_12152,N_11241,N_11903);
or U12153 (N_12153,N_11061,N_11407);
nand U12154 (N_12154,N_11659,N_11393);
nand U12155 (N_12155,N_11759,N_11657);
nor U12156 (N_12156,N_11908,N_11311);
or U12157 (N_12157,N_11893,N_11558);
xnor U12158 (N_12158,N_11981,N_11047);
nor U12159 (N_12159,N_11282,N_11459);
xnor U12160 (N_12160,N_11359,N_11268);
and U12161 (N_12161,N_11793,N_11783);
nand U12162 (N_12162,N_11670,N_11807);
nand U12163 (N_12163,N_11637,N_11305);
nor U12164 (N_12164,N_11736,N_11961);
xor U12165 (N_12165,N_11421,N_11841);
or U12166 (N_12166,N_11231,N_11326);
nand U12167 (N_12167,N_11507,N_11301);
nand U12168 (N_12168,N_11574,N_11442);
xnor U12169 (N_12169,N_11567,N_11940);
nor U12170 (N_12170,N_11962,N_11847);
xnor U12171 (N_12171,N_11737,N_11683);
or U12172 (N_12172,N_11225,N_11891);
and U12173 (N_12173,N_11808,N_11462);
or U12174 (N_12174,N_11605,N_11367);
or U12175 (N_12175,N_11372,N_11256);
xor U12176 (N_12176,N_11774,N_11040);
xor U12177 (N_12177,N_11205,N_11157);
xor U12178 (N_12178,N_11423,N_11960);
nand U12179 (N_12179,N_11874,N_11025);
or U12180 (N_12180,N_11001,N_11864);
or U12181 (N_12181,N_11922,N_11071);
or U12182 (N_12182,N_11930,N_11862);
nand U12183 (N_12183,N_11901,N_11417);
nor U12184 (N_12184,N_11298,N_11243);
nand U12185 (N_12185,N_11498,N_11357);
and U12186 (N_12186,N_11481,N_11754);
and U12187 (N_12187,N_11373,N_11185);
nand U12188 (N_12188,N_11172,N_11152);
or U12189 (N_12189,N_11365,N_11802);
or U12190 (N_12190,N_11133,N_11232);
and U12191 (N_12191,N_11007,N_11642);
nand U12192 (N_12192,N_11865,N_11810);
nor U12193 (N_12193,N_11496,N_11773);
and U12194 (N_12194,N_11552,N_11137);
xor U12195 (N_12195,N_11986,N_11966);
nand U12196 (N_12196,N_11985,N_11132);
and U12197 (N_12197,N_11546,N_11154);
and U12198 (N_12198,N_11751,N_11572);
nand U12199 (N_12199,N_11341,N_11663);
nand U12200 (N_12200,N_11896,N_11809);
and U12201 (N_12201,N_11244,N_11043);
and U12202 (N_12202,N_11811,N_11609);
or U12203 (N_12203,N_11146,N_11242);
nand U12204 (N_12204,N_11145,N_11910);
nand U12205 (N_12205,N_11287,N_11694);
or U12206 (N_12206,N_11404,N_11983);
or U12207 (N_12207,N_11079,N_11828);
and U12208 (N_12208,N_11667,N_11092);
nand U12209 (N_12209,N_11547,N_11131);
nor U12210 (N_12210,N_11688,N_11380);
or U12211 (N_12211,N_11885,N_11931);
nor U12212 (N_12212,N_11942,N_11037);
and U12213 (N_12213,N_11588,N_11902);
nand U12214 (N_12214,N_11753,N_11587);
xnor U12215 (N_12215,N_11581,N_11714);
nand U12216 (N_12216,N_11379,N_11136);
nor U12217 (N_12217,N_11804,N_11645);
or U12218 (N_12218,N_11859,N_11553);
or U12219 (N_12219,N_11265,N_11508);
nor U12220 (N_12220,N_11745,N_11412);
nor U12221 (N_12221,N_11996,N_11712);
xor U12222 (N_12222,N_11845,N_11030);
or U12223 (N_12223,N_11623,N_11441);
nor U12224 (N_12224,N_11196,N_11912);
and U12225 (N_12225,N_11452,N_11014);
or U12226 (N_12226,N_11943,N_11051);
nor U12227 (N_12227,N_11512,N_11522);
and U12228 (N_12228,N_11023,N_11953);
nor U12229 (N_12229,N_11126,N_11974);
nor U12230 (N_12230,N_11543,N_11200);
or U12231 (N_12231,N_11110,N_11733);
nor U12232 (N_12232,N_11527,N_11675);
or U12233 (N_12233,N_11436,N_11410);
or U12234 (N_12234,N_11309,N_11875);
nand U12235 (N_12235,N_11321,N_11414);
xnor U12236 (N_12236,N_11332,N_11624);
nor U12237 (N_12237,N_11704,N_11948);
nor U12238 (N_12238,N_11168,N_11619);
nand U12239 (N_12239,N_11457,N_11465);
and U12240 (N_12240,N_11907,N_11059);
or U12241 (N_12241,N_11338,N_11590);
or U12242 (N_12242,N_11391,N_11906);
or U12243 (N_12243,N_11795,N_11093);
xnor U12244 (N_12244,N_11764,N_11686);
nor U12245 (N_12245,N_11706,N_11677);
and U12246 (N_12246,N_11871,N_11194);
or U12247 (N_12247,N_11832,N_11556);
nor U12248 (N_12248,N_11233,N_11453);
and U12249 (N_12249,N_11086,N_11723);
or U12250 (N_12250,N_11088,N_11778);
and U12251 (N_12251,N_11882,N_11691);
nand U12252 (N_12252,N_11878,N_11824);
nand U12253 (N_12253,N_11246,N_11731);
nor U12254 (N_12254,N_11149,N_11772);
nand U12255 (N_12255,N_11270,N_11354);
and U12256 (N_12256,N_11426,N_11259);
nor U12257 (N_12257,N_11941,N_11271);
or U12258 (N_12258,N_11424,N_11164);
and U12259 (N_12259,N_11877,N_11606);
or U12260 (N_12260,N_11445,N_11396);
xnor U12261 (N_12261,N_11382,N_11535);
or U12262 (N_12262,N_11563,N_11010);
or U12263 (N_12263,N_11293,N_11016);
and U12264 (N_12264,N_11299,N_11376);
nor U12265 (N_12265,N_11116,N_11852);
nor U12266 (N_12266,N_11888,N_11696);
nor U12267 (N_12267,N_11532,N_11212);
nor U12268 (N_12268,N_11215,N_11223);
xor U12269 (N_12269,N_11443,N_11234);
or U12270 (N_12270,N_11701,N_11289);
or U12271 (N_12271,N_11214,N_11087);
xnor U12272 (N_12272,N_11471,N_11467);
or U12273 (N_12273,N_11204,N_11335);
nor U12274 (N_12274,N_11057,N_11188);
or U12275 (N_12275,N_11889,N_11235);
nor U12276 (N_12276,N_11805,N_11819);
or U12277 (N_12277,N_11334,N_11541);
xor U12278 (N_12278,N_11207,N_11430);
or U12279 (N_12279,N_11169,N_11784);
nand U12280 (N_12280,N_11639,N_11261);
xor U12281 (N_12281,N_11970,N_11935);
nand U12282 (N_12282,N_11634,N_11483);
nand U12283 (N_12283,N_11097,N_11416);
nor U12284 (N_12284,N_11392,N_11390);
nor U12285 (N_12285,N_11197,N_11703);
xor U12286 (N_12286,N_11448,N_11073);
or U12287 (N_12287,N_11142,N_11269);
and U12288 (N_12288,N_11952,N_11038);
and U12289 (N_12289,N_11306,N_11555);
nor U12290 (N_12290,N_11375,N_11266);
and U12291 (N_12291,N_11180,N_11124);
nand U12292 (N_12292,N_11503,N_11743);
or U12293 (N_12293,N_11344,N_11969);
or U12294 (N_12294,N_11054,N_11944);
and U12295 (N_12295,N_11735,N_11017);
and U12296 (N_12296,N_11836,N_11592);
nand U12297 (N_12297,N_11107,N_11622);
xnor U12298 (N_12298,N_11939,N_11937);
or U12299 (N_12299,N_11766,N_11485);
xnor U12300 (N_12300,N_11488,N_11770);
and U12301 (N_12301,N_11582,N_11163);
or U12302 (N_12302,N_11074,N_11820);
or U12303 (N_12303,N_11674,N_11053);
and U12304 (N_12304,N_11415,N_11193);
nor U12305 (N_12305,N_11141,N_11626);
nor U12306 (N_12306,N_11715,N_11361);
nand U12307 (N_12307,N_11658,N_11440);
or U12308 (N_12308,N_11537,N_11980);
xor U12309 (N_12309,N_11665,N_11434);
nand U12310 (N_12310,N_11589,N_11089);
or U12311 (N_12311,N_11352,N_11913);
or U12312 (N_12312,N_11880,N_11539);
nand U12313 (N_12313,N_11230,N_11388);
and U12314 (N_12314,N_11959,N_11202);
nand U12315 (N_12315,N_11075,N_11186);
and U12316 (N_12316,N_11798,N_11761);
nand U12317 (N_12317,N_11358,N_11402);
xnor U12318 (N_12318,N_11478,N_11021);
nor U12319 (N_12319,N_11288,N_11769);
xnor U12320 (N_12320,N_11610,N_11005);
or U12321 (N_12321,N_11052,N_11009);
or U12322 (N_12322,N_11002,N_11041);
nand U12323 (N_12323,N_11726,N_11312);
nor U12324 (N_12324,N_11013,N_11965);
or U12325 (N_12325,N_11967,N_11596);
and U12326 (N_12326,N_11472,N_11601);
or U12327 (N_12327,N_11267,N_11104);
or U12328 (N_12328,N_11060,N_11091);
nor U12329 (N_12329,N_11884,N_11822);
or U12330 (N_12330,N_11121,N_11347);
or U12331 (N_12331,N_11138,N_11262);
and U12332 (N_12332,N_11184,N_11022);
nor U12333 (N_12333,N_11979,N_11024);
or U12334 (N_12334,N_11128,N_11559);
nor U12335 (N_12335,N_11918,N_11561);
xor U12336 (N_12336,N_11765,N_11111);
nor U12337 (N_12337,N_11673,N_11034);
xor U12338 (N_12338,N_11019,N_11105);
and U12339 (N_12339,N_11209,N_11274);
and U12340 (N_12340,N_11571,N_11117);
nand U12341 (N_12341,N_11676,N_11400);
and U12342 (N_12342,N_11932,N_11171);
nand U12343 (N_12343,N_11984,N_11938);
and U12344 (N_12344,N_11272,N_11661);
nor U12345 (N_12345,N_11055,N_11904);
or U12346 (N_12346,N_11919,N_11964);
and U12347 (N_12347,N_11450,N_11800);
or U12348 (N_12348,N_11284,N_11879);
and U12349 (N_12349,N_11848,N_11135);
and U12350 (N_12350,N_11322,N_11177);
or U12351 (N_12351,N_11860,N_11439);
and U12352 (N_12352,N_11406,N_11857);
or U12353 (N_12353,N_11618,N_11755);
and U12354 (N_12354,N_11399,N_11886);
xnor U12355 (N_12355,N_11863,N_11220);
or U12356 (N_12356,N_11015,N_11224);
and U12357 (N_12357,N_11870,N_11869);
and U12358 (N_12358,N_11709,N_11905);
and U12359 (N_12359,N_11385,N_11850);
nand U12360 (N_12360,N_11656,N_11418);
nor U12361 (N_12361,N_11155,N_11319);
or U12362 (N_12362,N_11254,N_11444);
nand U12363 (N_12363,N_11068,N_11446);
or U12364 (N_12364,N_11405,N_11065);
xor U12365 (N_12365,N_11762,N_11591);
xor U12366 (N_12366,N_11345,N_11505);
and U12367 (N_12367,N_11258,N_11325);
and U12368 (N_12368,N_11096,N_11534);
nor U12369 (N_12369,N_11122,N_11148);
and U12370 (N_12370,N_11586,N_11314);
or U12371 (N_12371,N_11429,N_11842);
xnor U12372 (N_12372,N_11346,N_11090);
nand U12373 (N_12373,N_11568,N_11506);
nand U12374 (N_12374,N_11237,N_11499);
nor U12375 (N_12375,N_11998,N_11741);
and U12376 (N_12376,N_11868,N_11492);
or U12377 (N_12377,N_11978,N_11100);
nand U12378 (N_12378,N_11247,N_11602);
and U12379 (N_12379,N_11698,N_11158);
nor U12380 (N_12380,N_11632,N_11856);
or U12381 (N_12381,N_11078,N_11720);
and U12382 (N_12382,N_11945,N_11210);
nor U12383 (N_12383,N_11370,N_11353);
nor U12384 (N_12384,N_11630,N_11384);
nand U12385 (N_12385,N_11469,N_11218);
xor U12386 (N_12386,N_11320,N_11401);
and U12387 (N_12387,N_11119,N_11915);
nand U12388 (N_12388,N_11640,N_11108);
nand U12389 (N_12389,N_11636,N_11830);
nor U12390 (N_12390,N_11617,N_11861);
nor U12391 (N_12391,N_11629,N_11892);
nor U12392 (N_12392,N_11717,N_11729);
or U12393 (N_12393,N_11364,N_11176);
nand U12394 (N_12394,N_11838,N_11548);
nor U12395 (N_12395,N_11777,N_11858);
nor U12396 (N_12396,N_11725,N_11198);
nand U12397 (N_12397,N_11227,N_11557);
nor U12398 (N_12398,N_11782,N_11123);
and U12399 (N_12399,N_11064,N_11958);
or U12400 (N_12400,N_11063,N_11643);
and U12401 (N_12401,N_11292,N_11427);
nor U12402 (N_12402,N_11681,N_11330);
and U12403 (N_12403,N_11991,N_11813);
or U12404 (N_12404,N_11011,N_11056);
or U12405 (N_12405,N_11477,N_11044);
nand U12406 (N_12406,N_11530,N_11635);
and U12407 (N_12407,N_11825,N_11228);
and U12408 (N_12408,N_11413,N_11257);
and U12409 (N_12409,N_11608,N_11504);
or U12410 (N_12410,N_11584,N_11835);
or U12411 (N_12411,N_11995,N_11150);
nor U12412 (N_12412,N_11118,N_11514);
and U12413 (N_12413,N_11166,N_11790);
and U12414 (N_12414,N_11650,N_11732);
xor U12415 (N_12415,N_11080,N_11226);
nor U12416 (N_12416,N_11971,N_11707);
or U12417 (N_12417,N_11035,N_11791);
nor U12418 (N_12418,N_11684,N_11570);
nand U12419 (N_12419,N_11806,N_11662);
nand U12420 (N_12420,N_11799,N_11463);
nor U12421 (N_12421,N_11475,N_11917);
nor U12422 (N_12422,N_11768,N_11398);
nand U12423 (N_12423,N_11594,N_11451);
and U12424 (N_12424,N_11826,N_11562);
or U12425 (N_12425,N_11006,N_11045);
nand U12426 (N_12426,N_11307,N_11620);
and U12427 (N_12427,N_11447,N_11316);
and U12428 (N_12428,N_11576,N_11947);
nor U12429 (N_12429,N_11170,N_11911);
and U12430 (N_12430,N_11914,N_11513);
xnor U12431 (N_12431,N_11083,N_11102);
nor U12432 (N_12432,N_11313,N_11776);
and U12433 (N_12433,N_11550,N_11666);
or U12434 (N_12434,N_11245,N_11600);
and U12435 (N_12435,N_11012,N_11898);
nand U12436 (N_12436,N_11310,N_11595);
and U12437 (N_12437,N_11760,N_11631);
nand U12438 (N_12438,N_11921,N_11109);
and U12439 (N_12439,N_11331,N_11890);
and U12440 (N_12440,N_11740,N_11692);
nand U12441 (N_12441,N_11058,N_11317);
and U12442 (N_12442,N_11495,N_11817);
nor U12443 (N_12443,N_11789,N_11161);
or U12444 (N_12444,N_11999,N_11655);
nor U12445 (N_12445,N_11551,N_11229);
nand U12446 (N_12446,N_11989,N_11008);
nor U12447 (N_12447,N_11719,N_11156);
nor U12448 (N_12448,N_11263,N_11255);
nand U12449 (N_12449,N_11278,N_11621);
nand U12450 (N_12450,N_11827,N_11125);
or U12451 (N_12451,N_11583,N_11627);
nand U12452 (N_12452,N_11988,N_11934);
or U12453 (N_12453,N_11165,N_11378);
xnor U12454 (N_12454,N_11032,N_11579);
and U12455 (N_12455,N_11593,N_11699);
nand U12456 (N_12456,N_11050,N_11669);
nand U12457 (N_12457,N_11144,N_11113);
nor U12458 (N_12458,N_11470,N_11302);
or U12459 (N_12459,N_11538,N_11004);
and U12460 (N_12460,N_11280,N_11992);
and U12461 (N_12461,N_11461,N_11140);
and U12462 (N_12462,N_11873,N_11491);
and U12463 (N_12463,N_11702,N_11816);
nand U12464 (N_12464,N_11130,N_11028);
and U12465 (N_12465,N_11540,N_11236);
and U12466 (N_12466,N_11420,N_11599);
nand U12467 (N_12467,N_11549,N_11957);
nand U12468 (N_12468,N_11295,N_11260);
and U12469 (N_12469,N_11612,N_11371);
nand U12470 (N_12470,N_11823,N_11348);
nand U12471 (N_12471,N_11746,N_11653);
nor U12472 (N_12472,N_11189,N_11685);
and U12473 (N_12473,N_11897,N_11366);
or U12474 (N_12474,N_11654,N_11493);
nand U12475 (N_12475,N_11324,N_11987);
nand U12476 (N_12476,N_11815,N_11647);
or U12477 (N_12477,N_11337,N_11099);
and U12478 (N_12478,N_11291,N_11489);
or U12479 (N_12479,N_11308,N_11103);
or U12480 (N_12480,N_11682,N_11949);
nor U12481 (N_12481,N_11516,N_11780);
or U12482 (N_12482,N_11575,N_11206);
and U12483 (N_12483,N_11369,N_11597);
and U12484 (N_12484,N_11900,N_11721);
or U12485 (N_12485,N_11573,N_11221);
nand U12486 (N_12486,N_11664,N_11565);
nor U12487 (N_12487,N_11397,N_11603);
nand U12488 (N_12488,N_11678,N_11752);
and U12489 (N_12489,N_11027,N_11853);
or U12490 (N_12490,N_11355,N_11646);
nand U12491 (N_12491,N_11101,N_11377);
nor U12492 (N_12492,N_11340,N_11425);
xor U12493 (N_12493,N_11363,N_11727);
xnor U12494 (N_12494,N_11191,N_11098);
nor U12495 (N_12495,N_11048,N_11920);
or U12496 (N_12496,N_11968,N_11431);
or U12497 (N_12497,N_11139,N_11336);
or U12498 (N_12498,N_11834,N_11515);
nor U12499 (N_12499,N_11192,N_11771);
or U12500 (N_12500,N_11662,N_11594);
xor U12501 (N_12501,N_11102,N_11681);
nand U12502 (N_12502,N_11410,N_11876);
and U12503 (N_12503,N_11786,N_11853);
or U12504 (N_12504,N_11747,N_11492);
or U12505 (N_12505,N_11734,N_11660);
xor U12506 (N_12506,N_11029,N_11775);
nand U12507 (N_12507,N_11872,N_11619);
nand U12508 (N_12508,N_11548,N_11755);
nand U12509 (N_12509,N_11407,N_11952);
xnor U12510 (N_12510,N_11556,N_11207);
nand U12511 (N_12511,N_11915,N_11619);
and U12512 (N_12512,N_11299,N_11009);
nor U12513 (N_12513,N_11910,N_11250);
and U12514 (N_12514,N_11089,N_11830);
and U12515 (N_12515,N_11763,N_11094);
or U12516 (N_12516,N_11161,N_11753);
nand U12517 (N_12517,N_11178,N_11121);
nor U12518 (N_12518,N_11624,N_11152);
nand U12519 (N_12519,N_11399,N_11269);
nor U12520 (N_12520,N_11627,N_11559);
or U12521 (N_12521,N_11488,N_11896);
and U12522 (N_12522,N_11307,N_11793);
nor U12523 (N_12523,N_11010,N_11299);
or U12524 (N_12524,N_11323,N_11025);
nor U12525 (N_12525,N_11347,N_11698);
nor U12526 (N_12526,N_11695,N_11380);
or U12527 (N_12527,N_11158,N_11565);
nand U12528 (N_12528,N_11057,N_11962);
or U12529 (N_12529,N_11523,N_11420);
nor U12530 (N_12530,N_11100,N_11686);
xor U12531 (N_12531,N_11422,N_11210);
nor U12532 (N_12532,N_11583,N_11955);
xor U12533 (N_12533,N_11199,N_11917);
nand U12534 (N_12534,N_11665,N_11921);
and U12535 (N_12535,N_11057,N_11856);
nor U12536 (N_12536,N_11639,N_11101);
or U12537 (N_12537,N_11402,N_11320);
or U12538 (N_12538,N_11943,N_11827);
nor U12539 (N_12539,N_11863,N_11914);
nor U12540 (N_12540,N_11012,N_11291);
nor U12541 (N_12541,N_11475,N_11902);
nor U12542 (N_12542,N_11658,N_11973);
or U12543 (N_12543,N_11883,N_11952);
or U12544 (N_12544,N_11173,N_11309);
xor U12545 (N_12545,N_11137,N_11484);
and U12546 (N_12546,N_11983,N_11780);
nor U12547 (N_12547,N_11589,N_11695);
nand U12548 (N_12548,N_11194,N_11235);
nor U12549 (N_12549,N_11686,N_11463);
nor U12550 (N_12550,N_11130,N_11963);
or U12551 (N_12551,N_11036,N_11932);
nand U12552 (N_12552,N_11344,N_11576);
nor U12553 (N_12553,N_11095,N_11493);
or U12554 (N_12554,N_11536,N_11228);
or U12555 (N_12555,N_11221,N_11356);
or U12556 (N_12556,N_11734,N_11771);
or U12557 (N_12557,N_11999,N_11523);
nor U12558 (N_12558,N_11955,N_11734);
and U12559 (N_12559,N_11727,N_11708);
nand U12560 (N_12560,N_11361,N_11403);
nand U12561 (N_12561,N_11639,N_11393);
nand U12562 (N_12562,N_11244,N_11000);
nor U12563 (N_12563,N_11521,N_11485);
or U12564 (N_12564,N_11453,N_11912);
or U12565 (N_12565,N_11566,N_11355);
nand U12566 (N_12566,N_11456,N_11100);
and U12567 (N_12567,N_11255,N_11393);
nand U12568 (N_12568,N_11000,N_11732);
and U12569 (N_12569,N_11314,N_11466);
nand U12570 (N_12570,N_11109,N_11833);
nand U12571 (N_12571,N_11626,N_11347);
nand U12572 (N_12572,N_11437,N_11585);
and U12573 (N_12573,N_11588,N_11855);
nand U12574 (N_12574,N_11480,N_11388);
nor U12575 (N_12575,N_11132,N_11803);
or U12576 (N_12576,N_11683,N_11293);
or U12577 (N_12577,N_11976,N_11713);
or U12578 (N_12578,N_11848,N_11626);
nand U12579 (N_12579,N_11243,N_11877);
nor U12580 (N_12580,N_11816,N_11254);
or U12581 (N_12581,N_11227,N_11125);
or U12582 (N_12582,N_11212,N_11193);
or U12583 (N_12583,N_11694,N_11440);
or U12584 (N_12584,N_11048,N_11268);
nor U12585 (N_12585,N_11242,N_11708);
nor U12586 (N_12586,N_11167,N_11175);
and U12587 (N_12587,N_11638,N_11731);
nor U12588 (N_12588,N_11501,N_11967);
nand U12589 (N_12589,N_11774,N_11656);
and U12590 (N_12590,N_11091,N_11002);
nor U12591 (N_12591,N_11632,N_11652);
nand U12592 (N_12592,N_11498,N_11042);
xor U12593 (N_12593,N_11754,N_11158);
nor U12594 (N_12594,N_11695,N_11666);
nor U12595 (N_12595,N_11093,N_11448);
or U12596 (N_12596,N_11192,N_11127);
and U12597 (N_12597,N_11190,N_11306);
or U12598 (N_12598,N_11160,N_11110);
nand U12599 (N_12599,N_11579,N_11061);
nand U12600 (N_12600,N_11683,N_11668);
xnor U12601 (N_12601,N_11534,N_11698);
and U12602 (N_12602,N_11804,N_11971);
or U12603 (N_12603,N_11356,N_11401);
nand U12604 (N_12604,N_11791,N_11559);
xnor U12605 (N_12605,N_11189,N_11705);
nand U12606 (N_12606,N_11285,N_11891);
and U12607 (N_12607,N_11203,N_11042);
nand U12608 (N_12608,N_11272,N_11213);
and U12609 (N_12609,N_11327,N_11044);
xnor U12610 (N_12610,N_11776,N_11273);
and U12611 (N_12611,N_11735,N_11406);
xnor U12612 (N_12612,N_11548,N_11907);
or U12613 (N_12613,N_11549,N_11427);
nor U12614 (N_12614,N_11561,N_11576);
or U12615 (N_12615,N_11326,N_11451);
nor U12616 (N_12616,N_11371,N_11645);
or U12617 (N_12617,N_11555,N_11616);
or U12618 (N_12618,N_11266,N_11335);
or U12619 (N_12619,N_11161,N_11771);
or U12620 (N_12620,N_11428,N_11197);
or U12621 (N_12621,N_11397,N_11245);
or U12622 (N_12622,N_11282,N_11395);
nand U12623 (N_12623,N_11791,N_11248);
or U12624 (N_12624,N_11399,N_11286);
and U12625 (N_12625,N_11533,N_11420);
nand U12626 (N_12626,N_11200,N_11974);
nor U12627 (N_12627,N_11991,N_11392);
or U12628 (N_12628,N_11604,N_11512);
xnor U12629 (N_12629,N_11587,N_11476);
nand U12630 (N_12630,N_11722,N_11426);
nor U12631 (N_12631,N_11492,N_11914);
nand U12632 (N_12632,N_11611,N_11641);
or U12633 (N_12633,N_11594,N_11493);
or U12634 (N_12634,N_11422,N_11068);
nand U12635 (N_12635,N_11820,N_11472);
or U12636 (N_12636,N_11057,N_11748);
xnor U12637 (N_12637,N_11576,N_11825);
and U12638 (N_12638,N_11640,N_11445);
or U12639 (N_12639,N_11389,N_11899);
xor U12640 (N_12640,N_11771,N_11363);
nor U12641 (N_12641,N_11086,N_11107);
nor U12642 (N_12642,N_11413,N_11880);
or U12643 (N_12643,N_11142,N_11075);
nor U12644 (N_12644,N_11140,N_11474);
nand U12645 (N_12645,N_11475,N_11911);
nor U12646 (N_12646,N_11891,N_11057);
or U12647 (N_12647,N_11370,N_11398);
or U12648 (N_12648,N_11205,N_11998);
xnor U12649 (N_12649,N_11406,N_11961);
nor U12650 (N_12650,N_11592,N_11933);
or U12651 (N_12651,N_11560,N_11654);
or U12652 (N_12652,N_11420,N_11563);
nand U12653 (N_12653,N_11321,N_11730);
nand U12654 (N_12654,N_11896,N_11548);
xnor U12655 (N_12655,N_11004,N_11872);
nand U12656 (N_12656,N_11286,N_11753);
nor U12657 (N_12657,N_11756,N_11594);
nor U12658 (N_12658,N_11499,N_11213);
xor U12659 (N_12659,N_11050,N_11612);
nor U12660 (N_12660,N_11202,N_11382);
nand U12661 (N_12661,N_11785,N_11803);
and U12662 (N_12662,N_11929,N_11683);
and U12663 (N_12663,N_11924,N_11298);
and U12664 (N_12664,N_11282,N_11349);
or U12665 (N_12665,N_11004,N_11701);
and U12666 (N_12666,N_11924,N_11043);
nor U12667 (N_12667,N_11721,N_11028);
and U12668 (N_12668,N_11970,N_11070);
nor U12669 (N_12669,N_11943,N_11337);
nor U12670 (N_12670,N_11257,N_11955);
and U12671 (N_12671,N_11481,N_11570);
nand U12672 (N_12672,N_11717,N_11642);
nor U12673 (N_12673,N_11929,N_11775);
and U12674 (N_12674,N_11940,N_11248);
nand U12675 (N_12675,N_11498,N_11472);
nand U12676 (N_12676,N_11787,N_11761);
and U12677 (N_12677,N_11268,N_11567);
nor U12678 (N_12678,N_11536,N_11257);
or U12679 (N_12679,N_11121,N_11884);
nand U12680 (N_12680,N_11069,N_11498);
or U12681 (N_12681,N_11798,N_11680);
or U12682 (N_12682,N_11869,N_11554);
or U12683 (N_12683,N_11596,N_11619);
or U12684 (N_12684,N_11398,N_11626);
nor U12685 (N_12685,N_11574,N_11789);
nor U12686 (N_12686,N_11575,N_11638);
or U12687 (N_12687,N_11792,N_11411);
or U12688 (N_12688,N_11115,N_11455);
nand U12689 (N_12689,N_11683,N_11512);
nand U12690 (N_12690,N_11944,N_11475);
nand U12691 (N_12691,N_11036,N_11313);
or U12692 (N_12692,N_11268,N_11942);
nor U12693 (N_12693,N_11319,N_11912);
or U12694 (N_12694,N_11484,N_11682);
nand U12695 (N_12695,N_11452,N_11358);
nand U12696 (N_12696,N_11804,N_11485);
nand U12697 (N_12697,N_11618,N_11551);
nor U12698 (N_12698,N_11737,N_11661);
nand U12699 (N_12699,N_11302,N_11117);
nand U12700 (N_12700,N_11044,N_11002);
nand U12701 (N_12701,N_11548,N_11159);
and U12702 (N_12702,N_11282,N_11714);
nand U12703 (N_12703,N_11221,N_11359);
xor U12704 (N_12704,N_11518,N_11827);
or U12705 (N_12705,N_11781,N_11761);
or U12706 (N_12706,N_11353,N_11880);
nor U12707 (N_12707,N_11500,N_11660);
and U12708 (N_12708,N_11517,N_11557);
or U12709 (N_12709,N_11843,N_11245);
and U12710 (N_12710,N_11263,N_11349);
or U12711 (N_12711,N_11781,N_11231);
and U12712 (N_12712,N_11333,N_11564);
xnor U12713 (N_12713,N_11596,N_11652);
and U12714 (N_12714,N_11399,N_11991);
nor U12715 (N_12715,N_11087,N_11900);
nor U12716 (N_12716,N_11752,N_11320);
or U12717 (N_12717,N_11150,N_11964);
nand U12718 (N_12718,N_11811,N_11979);
nor U12719 (N_12719,N_11352,N_11456);
nand U12720 (N_12720,N_11209,N_11858);
nor U12721 (N_12721,N_11417,N_11422);
or U12722 (N_12722,N_11627,N_11012);
or U12723 (N_12723,N_11584,N_11950);
nand U12724 (N_12724,N_11181,N_11718);
or U12725 (N_12725,N_11586,N_11744);
and U12726 (N_12726,N_11076,N_11856);
and U12727 (N_12727,N_11913,N_11396);
or U12728 (N_12728,N_11787,N_11722);
xnor U12729 (N_12729,N_11219,N_11227);
nor U12730 (N_12730,N_11717,N_11657);
or U12731 (N_12731,N_11321,N_11998);
and U12732 (N_12732,N_11231,N_11833);
nor U12733 (N_12733,N_11238,N_11646);
or U12734 (N_12734,N_11283,N_11434);
nor U12735 (N_12735,N_11407,N_11715);
xnor U12736 (N_12736,N_11599,N_11976);
nand U12737 (N_12737,N_11861,N_11106);
nor U12738 (N_12738,N_11345,N_11921);
or U12739 (N_12739,N_11914,N_11472);
and U12740 (N_12740,N_11279,N_11592);
nor U12741 (N_12741,N_11250,N_11641);
and U12742 (N_12742,N_11822,N_11940);
and U12743 (N_12743,N_11023,N_11689);
and U12744 (N_12744,N_11119,N_11654);
nand U12745 (N_12745,N_11999,N_11216);
nor U12746 (N_12746,N_11402,N_11711);
or U12747 (N_12747,N_11922,N_11969);
and U12748 (N_12748,N_11909,N_11926);
nor U12749 (N_12749,N_11331,N_11727);
or U12750 (N_12750,N_11957,N_11907);
and U12751 (N_12751,N_11704,N_11384);
nor U12752 (N_12752,N_11609,N_11080);
xnor U12753 (N_12753,N_11667,N_11105);
nor U12754 (N_12754,N_11819,N_11292);
nand U12755 (N_12755,N_11149,N_11169);
nand U12756 (N_12756,N_11695,N_11447);
and U12757 (N_12757,N_11111,N_11549);
and U12758 (N_12758,N_11281,N_11356);
or U12759 (N_12759,N_11615,N_11537);
xor U12760 (N_12760,N_11409,N_11063);
and U12761 (N_12761,N_11139,N_11100);
or U12762 (N_12762,N_11630,N_11237);
nor U12763 (N_12763,N_11167,N_11734);
and U12764 (N_12764,N_11731,N_11783);
nand U12765 (N_12765,N_11593,N_11022);
nor U12766 (N_12766,N_11769,N_11528);
and U12767 (N_12767,N_11377,N_11470);
nor U12768 (N_12768,N_11728,N_11653);
nor U12769 (N_12769,N_11970,N_11417);
or U12770 (N_12770,N_11602,N_11348);
nand U12771 (N_12771,N_11599,N_11325);
nor U12772 (N_12772,N_11357,N_11859);
nand U12773 (N_12773,N_11502,N_11024);
or U12774 (N_12774,N_11663,N_11800);
xor U12775 (N_12775,N_11616,N_11997);
nand U12776 (N_12776,N_11190,N_11201);
nor U12777 (N_12777,N_11072,N_11211);
xor U12778 (N_12778,N_11908,N_11826);
and U12779 (N_12779,N_11880,N_11627);
xor U12780 (N_12780,N_11087,N_11959);
nand U12781 (N_12781,N_11263,N_11759);
or U12782 (N_12782,N_11378,N_11137);
nand U12783 (N_12783,N_11336,N_11679);
nand U12784 (N_12784,N_11312,N_11531);
xor U12785 (N_12785,N_11770,N_11086);
nand U12786 (N_12786,N_11109,N_11444);
nor U12787 (N_12787,N_11713,N_11207);
nor U12788 (N_12788,N_11158,N_11718);
nand U12789 (N_12789,N_11154,N_11687);
and U12790 (N_12790,N_11551,N_11909);
and U12791 (N_12791,N_11892,N_11814);
and U12792 (N_12792,N_11660,N_11018);
nor U12793 (N_12793,N_11524,N_11237);
or U12794 (N_12794,N_11238,N_11212);
nor U12795 (N_12795,N_11463,N_11048);
nor U12796 (N_12796,N_11059,N_11278);
or U12797 (N_12797,N_11235,N_11056);
nor U12798 (N_12798,N_11044,N_11694);
xnor U12799 (N_12799,N_11561,N_11279);
nand U12800 (N_12800,N_11504,N_11689);
or U12801 (N_12801,N_11650,N_11448);
xnor U12802 (N_12802,N_11909,N_11427);
nor U12803 (N_12803,N_11837,N_11831);
xor U12804 (N_12804,N_11394,N_11608);
nand U12805 (N_12805,N_11092,N_11339);
nor U12806 (N_12806,N_11832,N_11686);
nor U12807 (N_12807,N_11000,N_11050);
nand U12808 (N_12808,N_11664,N_11466);
and U12809 (N_12809,N_11853,N_11206);
nor U12810 (N_12810,N_11833,N_11759);
nor U12811 (N_12811,N_11765,N_11767);
nor U12812 (N_12812,N_11276,N_11000);
nand U12813 (N_12813,N_11443,N_11926);
nand U12814 (N_12814,N_11266,N_11001);
nand U12815 (N_12815,N_11523,N_11341);
nand U12816 (N_12816,N_11221,N_11787);
nor U12817 (N_12817,N_11952,N_11071);
or U12818 (N_12818,N_11827,N_11420);
and U12819 (N_12819,N_11147,N_11629);
nand U12820 (N_12820,N_11672,N_11951);
and U12821 (N_12821,N_11463,N_11304);
nor U12822 (N_12822,N_11900,N_11266);
nand U12823 (N_12823,N_11553,N_11828);
and U12824 (N_12824,N_11569,N_11393);
nand U12825 (N_12825,N_11275,N_11875);
or U12826 (N_12826,N_11248,N_11741);
nor U12827 (N_12827,N_11248,N_11745);
and U12828 (N_12828,N_11455,N_11435);
and U12829 (N_12829,N_11711,N_11142);
or U12830 (N_12830,N_11544,N_11700);
or U12831 (N_12831,N_11568,N_11195);
xor U12832 (N_12832,N_11087,N_11349);
nor U12833 (N_12833,N_11294,N_11627);
or U12834 (N_12834,N_11636,N_11938);
or U12835 (N_12835,N_11128,N_11250);
and U12836 (N_12836,N_11641,N_11920);
or U12837 (N_12837,N_11860,N_11145);
xnor U12838 (N_12838,N_11126,N_11934);
or U12839 (N_12839,N_11230,N_11409);
nor U12840 (N_12840,N_11569,N_11769);
nor U12841 (N_12841,N_11081,N_11009);
nand U12842 (N_12842,N_11206,N_11048);
or U12843 (N_12843,N_11247,N_11409);
xnor U12844 (N_12844,N_11289,N_11851);
and U12845 (N_12845,N_11841,N_11569);
xnor U12846 (N_12846,N_11558,N_11935);
nand U12847 (N_12847,N_11236,N_11981);
nand U12848 (N_12848,N_11428,N_11583);
nand U12849 (N_12849,N_11425,N_11471);
and U12850 (N_12850,N_11740,N_11183);
nor U12851 (N_12851,N_11425,N_11370);
nor U12852 (N_12852,N_11766,N_11802);
or U12853 (N_12853,N_11052,N_11175);
xnor U12854 (N_12854,N_11399,N_11264);
nand U12855 (N_12855,N_11590,N_11726);
or U12856 (N_12856,N_11949,N_11232);
or U12857 (N_12857,N_11765,N_11566);
or U12858 (N_12858,N_11921,N_11484);
nor U12859 (N_12859,N_11799,N_11422);
xor U12860 (N_12860,N_11973,N_11764);
and U12861 (N_12861,N_11503,N_11332);
and U12862 (N_12862,N_11715,N_11781);
xor U12863 (N_12863,N_11571,N_11417);
nor U12864 (N_12864,N_11625,N_11376);
nor U12865 (N_12865,N_11701,N_11827);
nor U12866 (N_12866,N_11297,N_11063);
or U12867 (N_12867,N_11625,N_11654);
and U12868 (N_12868,N_11673,N_11710);
nand U12869 (N_12869,N_11545,N_11760);
and U12870 (N_12870,N_11063,N_11113);
nand U12871 (N_12871,N_11054,N_11836);
nand U12872 (N_12872,N_11781,N_11066);
and U12873 (N_12873,N_11525,N_11963);
nor U12874 (N_12874,N_11014,N_11350);
nand U12875 (N_12875,N_11399,N_11420);
and U12876 (N_12876,N_11816,N_11541);
nand U12877 (N_12877,N_11361,N_11614);
nor U12878 (N_12878,N_11609,N_11603);
and U12879 (N_12879,N_11034,N_11401);
or U12880 (N_12880,N_11721,N_11072);
or U12881 (N_12881,N_11093,N_11095);
nand U12882 (N_12882,N_11155,N_11686);
and U12883 (N_12883,N_11238,N_11180);
or U12884 (N_12884,N_11922,N_11615);
nor U12885 (N_12885,N_11517,N_11531);
nand U12886 (N_12886,N_11580,N_11004);
xor U12887 (N_12887,N_11120,N_11638);
xnor U12888 (N_12888,N_11249,N_11711);
or U12889 (N_12889,N_11609,N_11496);
and U12890 (N_12890,N_11143,N_11572);
and U12891 (N_12891,N_11973,N_11496);
or U12892 (N_12892,N_11025,N_11041);
or U12893 (N_12893,N_11166,N_11235);
and U12894 (N_12894,N_11985,N_11564);
nand U12895 (N_12895,N_11134,N_11507);
xor U12896 (N_12896,N_11789,N_11241);
nand U12897 (N_12897,N_11631,N_11179);
or U12898 (N_12898,N_11017,N_11036);
xnor U12899 (N_12899,N_11872,N_11366);
or U12900 (N_12900,N_11246,N_11307);
nor U12901 (N_12901,N_11474,N_11550);
xnor U12902 (N_12902,N_11675,N_11299);
xor U12903 (N_12903,N_11265,N_11598);
nand U12904 (N_12904,N_11998,N_11994);
xor U12905 (N_12905,N_11489,N_11064);
nand U12906 (N_12906,N_11900,N_11993);
nand U12907 (N_12907,N_11319,N_11698);
and U12908 (N_12908,N_11351,N_11454);
nand U12909 (N_12909,N_11999,N_11997);
xor U12910 (N_12910,N_11927,N_11531);
nor U12911 (N_12911,N_11105,N_11098);
nand U12912 (N_12912,N_11993,N_11446);
nor U12913 (N_12913,N_11472,N_11204);
nor U12914 (N_12914,N_11116,N_11542);
xor U12915 (N_12915,N_11200,N_11111);
or U12916 (N_12916,N_11703,N_11746);
and U12917 (N_12917,N_11333,N_11586);
or U12918 (N_12918,N_11053,N_11637);
nand U12919 (N_12919,N_11566,N_11808);
nand U12920 (N_12920,N_11472,N_11049);
nand U12921 (N_12921,N_11932,N_11142);
and U12922 (N_12922,N_11374,N_11935);
or U12923 (N_12923,N_11400,N_11823);
nand U12924 (N_12924,N_11723,N_11020);
and U12925 (N_12925,N_11778,N_11788);
nand U12926 (N_12926,N_11485,N_11482);
nor U12927 (N_12927,N_11632,N_11165);
nor U12928 (N_12928,N_11388,N_11688);
and U12929 (N_12929,N_11306,N_11225);
and U12930 (N_12930,N_11334,N_11480);
nand U12931 (N_12931,N_11838,N_11717);
nand U12932 (N_12932,N_11050,N_11963);
or U12933 (N_12933,N_11005,N_11002);
or U12934 (N_12934,N_11200,N_11674);
or U12935 (N_12935,N_11406,N_11356);
nor U12936 (N_12936,N_11442,N_11239);
xor U12937 (N_12937,N_11038,N_11231);
or U12938 (N_12938,N_11692,N_11345);
nand U12939 (N_12939,N_11989,N_11689);
nor U12940 (N_12940,N_11918,N_11994);
or U12941 (N_12941,N_11010,N_11513);
nand U12942 (N_12942,N_11969,N_11914);
and U12943 (N_12943,N_11737,N_11324);
or U12944 (N_12944,N_11161,N_11830);
and U12945 (N_12945,N_11798,N_11845);
and U12946 (N_12946,N_11030,N_11041);
or U12947 (N_12947,N_11250,N_11284);
nand U12948 (N_12948,N_11614,N_11120);
or U12949 (N_12949,N_11276,N_11289);
nand U12950 (N_12950,N_11174,N_11175);
xor U12951 (N_12951,N_11540,N_11526);
and U12952 (N_12952,N_11057,N_11238);
nand U12953 (N_12953,N_11597,N_11382);
and U12954 (N_12954,N_11243,N_11426);
and U12955 (N_12955,N_11316,N_11782);
xnor U12956 (N_12956,N_11299,N_11954);
nor U12957 (N_12957,N_11221,N_11884);
or U12958 (N_12958,N_11358,N_11604);
nor U12959 (N_12959,N_11230,N_11654);
and U12960 (N_12960,N_11982,N_11943);
nand U12961 (N_12961,N_11420,N_11761);
or U12962 (N_12962,N_11179,N_11817);
xor U12963 (N_12963,N_11992,N_11634);
nand U12964 (N_12964,N_11022,N_11115);
nand U12965 (N_12965,N_11525,N_11061);
nor U12966 (N_12966,N_11656,N_11800);
or U12967 (N_12967,N_11369,N_11878);
xor U12968 (N_12968,N_11666,N_11382);
or U12969 (N_12969,N_11513,N_11678);
nand U12970 (N_12970,N_11789,N_11183);
and U12971 (N_12971,N_11993,N_11597);
nand U12972 (N_12972,N_11714,N_11983);
or U12973 (N_12973,N_11564,N_11089);
nand U12974 (N_12974,N_11653,N_11439);
xnor U12975 (N_12975,N_11388,N_11826);
nor U12976 (N_12976,N_11837,N_11020);
and U12977 (N_12977,N_11532,N_11464);
nand U12978 (N_12978,N_11504,N_11371);
nand U12979 (N_12979,N_11497,N_11234);
xor U12980 (N_12980,N_11361,N_11245);
xnor U12981 (N_12981,N_11224,N_11989);
or U12982 (N_12982,N_11156,N_11191);
nand U12983 (N_12983,N_11119,N_11921);
or U12984 (N_12984,N_11533,N_11557);
and U12985 (N_12985,N_11016,N_11320);
or U12986 (N_12986,N_11491,N_11275);
nand U12987 (N_12987,N_11005,N_11590);
or U12988 (N_12988,N_11301,N_11085);
and U12989 (N_12989,N_11554,N_11144);
or U12990 (N_12990,N_11468,N_11646);
nor U12991 (N_12991,N_11184,N_11649);
nor U12992 (N_12992,N_11074,N_11251);
or U12993 (N_12993,N_11137,N_11079);
and U12994 (N_12994,N_11087,N_11027);
and U12995 (N_12995,N_11078,N_11922);
nand U12996 (N_12996,N_11024,N_11149);
nor U12997 (N_12997,N_11878,N_11424);
and U12998 (N_12998,N_11130,N_11701);
and U12999 (N_12999,N_11402,N_11113);
nor U13000 (N_13000,N_12265,N_12378);
nor U13001 (N_13001,N_12286,N_12898);
or U13002 (N_13002,N_12244,N_12587);
or U13003 (N_13003,N_12875,N_12781);
and U13004 (N_13004,N_12185,N_12803);
nand U13005 (N_13005,N_12178,N_12609);
nand U13006 (N_13006,N_12353,N_12094);
nand U13007 (N_13007,N_12801,N_12374);
and U13008 (N_13008,N_12261,N_12923);
or U13009 (N_13009,N_12561,N_12562);
nor U13010 (N_13010,N_12419,N_12070);
nor U13011 (N_13011,N_12922,N_12861);
nand U13012 (N_13012,N_12677,N_12766);
and U13013 (N_13013,N_12678,N_12951);
nand U13014 (N_13014,N_12571,N_12614);
or U13015 (N_13015,N_12332,N_12251);
nor U13016 (N_13016,N_12313,N_12514);
xnor U13017 (N_13017,N_12119,N_12640);
xor U13018 (N_13018,N_12664,N_12838);
nand U13019 (N_13019,N_12279,N_12130);
nand U13020 (N_13020,N_12260,N_12969);
and U13021 (N_13021,N_12051,N_12168);
xor U13022 (N_13022,N_12596,N_12320);
nor U13023 (N_13023,N_12852,N_12179);
nand U13024 (N_13024,N_12991,N_12149);
and U13025 (N_13025,N_12809,N_12485);
nand U13026 (N_13026,N_12800,N_12533);
nand U13027 (N_13027,N_12856,N_12772);
and U13028 (N_13028,N_12398,N_12407);
xor U13029 (N_13029,N_12518,N_12140);
or U13030 (N_13030,N_12906,N_12421);
and U13031 (N_13031,N_12019,N_12034);
nor U13032 (N_13032,N_12209,N_12584);
and U13033 (N_13033,N_12931,N_12732);
nand U13034 (N_13034,N_12045,N_12524);
nor U13035 (N_13035,N_12655,N_12764);
and U13036 (N_13036,N_12065,N_12462);
nor U13037 (N_13037,N_12897,N_12097);
nand U13038 (N_13038,N_12768,N_12158);
or U13039 (N_13039,N_12641,N_12101);
and U13040 (N_13040,N_12373,N_12709);
or U13041 (N_13041,N_12563,N_12936);
nor U13042 (N_13042,N_12984,N_12187);
and U13043 (N_13043,N_12659,N_12361);
or U13044 (N_13044,N_12352,N_12108);
nand U13045 (N_13045,N_12685,N_12282);
and U13046 (N_13046,N_12952,N_12267);
nand U13047 (N_13047,N_12109,N_12935);
or U13048 (N_13048,N_12157,N_12970);
nor U13049 (N_13049,N_12876,N_12203);
or U13050 (N_13050,N_12274,N_12428);
and U13051 (N_13051,N_12152,N_12191);
or U13052 (N_13052,N_12711,N_12560);
xor U13053 (N_13053,N_12002,N_12750);
or U13054 (N_13054,N_12758,N_12473);
or U13055 (N_13055,N_12722,N_12183);
xnor U13056 (N_13056,N_12981,N_12067);
nor U13057 (N_13057,N_12248,N_12872);
and U13058 (N_13058,N_12280,N_12502);
and U13059 (N_13059,N_12674,N_12782);
nor U13060 (N_13060,N_12276,N_12322);
nor U13061 (N_13061,N_12698,N_12375);
or U13062 (N_13062,N_12258,N_12504);
and U13063 (N_13063,N_12371,N_12586);
nand U13064 (N_13064,N_12329,N_12048);
nor U13065 (N_13065,N_12337,N_12864);
nand U13066 (N_13066,N_12488,N_12028);
nand U13067 (N_13067,N_12040,N_12061);
nand U13068 (N_13068,N_12435,N_12813);
or U13069 (N_13069,N_12619,N_12249);
xor U13070 (N_13070,N_12930,N_12990);
or U13071 (N_13071,N_12620,N_12921);
nand U13072 (N_13072,N_12779,N_12233);
xor U13073 (N_13073,N_12348,N_12475);
or U13074 (N_13074,N_12114,N_12938);
and U13075 (N_13075,N_12113,N_12683);
xor U13076 (N_13076,N_12010,N_12622);
nand U13077 (N_13077,N_12243,N_12252);
nor U13078 (N_13078,N_12066,N_12994);
or U13079 (N_13079,N_12013,N_12845);
nand U13080 (N_13080,N_12769,N_12391);
nor U13081 (N_13081,N_12738,N_12112);
nand U13082 (N_13082,N_12492,N_12886);
nand U13083 (N_13083,N_12083,N_12552);
and U13084 (N_13084,N_12023,N_12174);
and U13085 (N_13085,N_12145,N_12694);
nor U13086 (N_13086,N_12650,N_12041);
or U13087 (N_13087,N_12059,N_12491);
and U13088 (N_13088,N_12874,N_12626);
and U13089 (N_13089,N_12601,N_12850);
or U13090 (N_13090,N_12617,N_12849);
and U13091 (N_13091,N_12461,N_12530);
nand U13092 (N_13092,N_12494,N_12645);
nand U13093 (N_13093,N_12841,N_12554);
xnor U13094 (N_13094,N_12383,N_12965);
or U13095 (N_13095,N_12298,N_12259);
nor U13096 (N_13096,N_12172,N_12885);
nor U13097 (N_13097,N_12076,N_12700);
nand U13098 (N_13098,N_12791,N_12237);
nor U13099 (N_13099,N_12442,N_12519);
or U13100 (N_13100,N_12806,N_12598);
and U13101 (N_13101,N_12281,N_12808);
nor U13102 (N_13102,N_12205,N_12765);
nand U13103 (N_13103,N_12301,N_12451);
and U13104 (N_13104,N_12777,N_12229);
and U13105 (N_13105,N_12574,N_12448);
nand U13106 (N_13106,N_12250,N_12216);
or U13107 (N_13107,N_12624,N_12141);
and U13108 (N_13108,N_12033,N_12543);
and U13109 (N_13109,N_12816,N_12426);
and U13110 (N_13110,N_12135,N_12427);
nand U13111 (N_13111,N_12042,N_12465);
and U13112 (N_13112,N_12523,N_12107);
and U13113 (N_13113,N_12230,N_12939);
nand U13114 (N_13114,N_12382,N_12314);
nor U13115 (N_13115,N_12908,N_12745);
and U13116 (N_13116,N_12170,N_12054);
or U13117 (N_13117,N_12565,N_12629);
xor U13118 (N_13118,N_12416,N_12328);
nor U13119 (N_13119,N_12794,N_12495);
nand U13120 (N_13120,N_12522,N_12792);
or U13121 (N_13121,N_12163,N_12331);
or U13122 (N_13122,N_12394,N_12103);
or U13123 (N_13123,N_12245,N_12253);
and U13124 (N_13124,N_12049,N_12892);
nand U13125 (N_13125,N_12759,N_12775);
and U13126 (N_13126,N_12651,N_12521);
nand U13127 (N_13127,N_12275,N_12729);
nand U13128 (N_13128,N_12310,N_12973);
and U13129 (N_13129,N_12068,N_12071);
xor U13130 (N_13130,N_12096,N_12150);
and U13131 (N_13131,N_12215,N_12305);
or U13132 (N_13132,N_12404,N_12544);
and U13133 (N_13133,N_12551,N_12408);
or U13134 (N_13134,N_12716,N_12138);
and U13135 (N_13135,N_12901,N_12866);
nand U13136 (N_13136,N_12920,N_12463);
and U13137 (N_13137,N_12880,N_12480);
nand U13138 (N_13138,N_12748,N_12038);
xor U13139 (N_13139,N_12757,N_12628);
or U13140 (N_13140,N_12860,N_12293);
nand U13141 (N_13141,N_12025,N_12667);
or U13142 (N_13142,N_12985,N_12316);
or U13143 (N_13143,N_12290,N_12754);
or U13144 (N_13144,N_12919,N_12625);
or U13145 (N_13145,N_12032,N_12988);
nand U13146 (N_13146,N_12827,N_12616);
or U13147 (N_13147,N_12865,N_12610);
nor U13148 (N_13148,N_12199,N_12273);
xnor U13149 (N_13149,N_12003,N_12085);
or U13150 (N_13150,N_12099,N_12266);
nand U13151 (N_13151,N_12893,N_12555);
nand U13152 (N_13152,N_12749,N_12847);
nor U13153 (N_13153,N_12161,N_12029);
nor U13154 (N_13154,N_12569,N_12978);
nor U13155 (N_13155,N_12821,N_12081);
or U13156 (N_13156,N_12929,N_12499);
xor U13157 (N_13157,N_12330,N_12830);
nand U13158 (N_13158,N_12545,N_12341);
and U13159 (N_13159,N_12882,N_12899);
nor U13160 (N_13160,N_12136,N_12501);
nor U13161 (N_13161,N_12770,N_12190);
and U13162 (N_13162,N_12222,N_12660);
xnor U13163 (N_13163,N_12902,N_12015);
nor U13164 (N_13164,N_12840,N_12944);
nor U13165 (N_13165,N_12110,N_12911);
nand U13166 (N_13166,N_12868,N_12834);
and U13167 (N_13167,N_12934,N_12916);
or U13168 (N_13168,N_12043,N_12401);
nand U13169 (N_13169,N_12134,N_12747);
or U13170 (N_13170,N_12125,N_12637);
xnor U13171 (N_13171,N_12481,N_12387);
nand U13172 (N_13172,N_12546,N_12143);
nand U13173 (N_13173,N_12206,N_12208);
or U13174 (N_13174,N_12318,N_12513);
xor U13175 (N_13175,N_12195,N_12837);
nor U13176 (N_13176,N_12184,N_12350);
xor U13177 (N_13177,N_12011,N_12009);
and U13178 (N_13178,N_12117,N_12527);
or U13179 (N_13179,N_12839,N_12675);
and U13180 (N_13180,N_12086,N_12780);
nand U13181 (N_13181,N_12345,N_12133);
nor U13182 (N_13182,N_12520,N_12169);
or U13183 (N_13183,N_12851,N_12867);
xor U13184 (N_13184,N_12436,N_12805);
nor U13185 (N_13185,N_12662,N_12787);
or U13186 (N_13186,N_12347,N_12746);
nor U13187 (N_13187,N_12017,N_12654);
or U13188 (N_13188,N_12257,N_12093);
nand U13189 (N_13189,N_12665,N_12763);
and U13190 (N_13190,N_12294,N_12171);
or U13191 (N_13191,N_12949,N_12269);
or U13192 (N_13192,N_12734,N_12004);
xnor U13193 (N_13193,N_12497,N_12606);
or U13194 (N_13194,N_12723,N_12611);
or U13195 (N_13195,N_12046,N_12104);
and U13196 (N_13196,N_12486,N_12728);
nor U13197 (N_13197,N_12340,N_12388);
or U13198 (N_13198,N_12795,N_12317);
nand U13199 (N_13199,N_12210,N_12470);
nor U13200 (N_13200,N_12559,N_12026);
and U13201 (N_13201,N_12997,N_12979);
nand U13202 (N_13202,N_12177,N_12558);
nor U13203 (N_13203,N_12307,N_12213);
and U13204 (N_13204,N_12537,N_12115);
or U13205 (N_13205,N_12579,N_12553);
or U13206 (N_13206,N_12682,N_12464);
and U13207 (N_13207,N_12376,N_12385);
nand U13208 (N_13208,N_12365,N_12162);
nand U13209 (N_13209,N_12087,N_12724);
and U13210 (N_13210,N_12439,N_12164);
and U13211 (N_13211,N_12466,N_12272);
or U13212 (N_13212,N_12928,N_12599);
and U13213 (N_13213,N_12189,N_12308);
nand U13214 (N_13214,N_12594,N_12453);
and U13215 (N_13215,N_12820,N_12968);
nor U13216 (N_13216,N_12336,N_12590);
nor U13217 (N_13217,N_12062,N_12894);
nor U13218 (N_13218,N_12855,N_12566);
or U13219 (N_13219,N_12315,N_12440);
or U13220 (N_13220,N_12604,N_12680);
or U13221 (N_13221,N_12570,N_12532);
nand U13222 (N_13222,N_12511,N_12409);
nand U13223 (N_13223,N_12550,N_12073);
nand U13224 (N_13224,N_12681,N_12263);
xor U13225 (N_13225,N_12719,N_12088);
or U13226 (N_13226,N_12648,N_12151);
nor U13227 (N_13227,N_12679,N_12832);
or U13228 (N_13228,N_12612,N_12891);
nor U13229 (N_13229,N_12129,N_12717);
nor U13230 (N_13230,N_12535,N_12600);
and U13231 (N_13231,N_12471,N_12585);
nor U13232 (N_13232,N_12959,N_12016);
or U13233 (N_13233,N_12507,N_12863);
or U13234 (N_13234,N_12581,N_12656);
and U13235 (N_13235,N_12718,N_12676);
and U13236 (N_13236,N_12720,N_12159);
nor U13237 (N_13237,N_12778,N_12074);
xnor U13238 (N_13238,N_12057,N_12506);
or U13239 (N_13239,N_12418,N_12262);
xor U13240 (N_13240,N_12726,N_12657);
nand U13241 (N_13241,N_12767,N_12549);
and U13242 (N_13242,N_12669,N_12696);
or U13243 (N_13243,N_12181,N_12793);
or U13244 (N_13244,N_12338,N_12605);
xnor U13245 (N_13245,N_12105,N_12744);
nor U13246 (N_13246,N_12202,N_12536);
and U13247 (N_13247,N_12366,N_12241);
and U13248 (N_13248,N_12166,N_12644);
nand U13249 (N_13249,N_12354,N_12895);
and U13250 (N_13250,N_12888,N_12390);
or U13251 (N_13251,N_12214,N_12814);
nand U13252 (N_13252,N_12455,N_12001);
nand U13253 (N_13253,N_12077,N_12924);
and U13254 (N_13254,N_12092,N_12053);
or U13255 (N_13255,N_12913,N_12483);
nor U13256 (N_13256,N_12635,N_12634);
or U13257 (N_13257,N_12235,N_12627);
or U13258 (N_13258,N_12992,N_12283);
or U13259 (N_13259,N_12384,N_12608);
nor U13260 (N_13260,N_12417,N_12231);
or U13261 (N_13261,N_12413,N_12498);
nor U13262 (N_13262,N_12907,N_12349);
nor U13263 (N_13263,N_12014,N_12836);
nand U13264 (N_13264,N_12783,N_12446);
or U13265 (N_13265,N_12410,N_12264);
nor U13266 (N_13266,N_12091,N_12713);
xor U13267 (N_13267,N_12246,N_12126);
and U13268 (N_13268,N_12324,N_12437);
and U13269 (N_13269,N_12226,N_12429);
or U13270 (N_13270,N_12363,N_12842);
nand U13271 (N_13271,N_12695,N_12510);
and U13272 (N_13272,N_12423,N_12459);
xor U13273 (N_13273,N_12714,N_12996);
nor U13274 (N_13274,N_12873,N_12771);
nand U13275 (N_13275,N_12295,N_12344);
nor U13276 (N_13276,N_12036,N_12961);
xnor U13277 (N_13277,N_12478,N_12567);
nor U13278 (N_13278,N_12291,N_12197);
xor U13279 (N_13279,N_12623,N_12173);
and U13280 (N_13280,N_12127,N_12207);
nor U13281 (N_13281,N_12904,N_12037);
nor U13282 (N_13282,N_12686,N_12304);
and U13283 (N_13283,N_12831,N_12706);
and U13284 (N_13284,N_12699,N_12572);
and U13285 (N_13285,N_12854,N_12217);
or U13286 (N_13286,N_12303,N_12346);
nand U13287 (N_13287,N_12693,N_12937);
or U13288 (N_13288,N_12727,N_12517);
and U13289 (N_13289,N_12691,N_12646);
nand U13290 (N_13290,N_12548,N_12684);
nand U13291 (N_13291,N_12432,N_12639);
nand U13292 (N_13292,N_12529,N_12377);
nand U13293 (N_13293,N_12721,N_12974);
and U13294 (N_13294,N_12224,N_12080);
or U13295 (N_13295,N_12687,N_12121);
nor U13296 (N_13296,N_12386,N_12064);
nand U13297 (N_13297,N_12602,N_12180);
or U13298 (N_13298,N_12773,N_12397);
and U13299 (N_13299,N_12415,N_12167);
nor U13300 (N_13300,N_12542,N_12756);
nand U13301 (N_13301,N_12306,N_12058);
nand U13302 (N_13302,N_12673,N_12024);
and U13303 (N_13303,N_12035,N_12467);
or U13304 (N_13304,N_12829,N_12367);
nand U13305 (N_13305,N_12582,N_12192);
and U13306 (N_13306,N_12148,N_12633);
xor U13307 (N_13307,N_12896,N_12325);
and U13308 (N_13308,N_12578,N_12342);
nor U13309 (N_13309,N_12503,N_12715);
nor U13310 (N_13310,N_12790,N_12457);
nand U13311 (N_13311,N_12999,N_12116);
nand U13312 (N_13312,N_12881,N_12577);
nand U13313 (N_13313,N_12326,N_12406);
xnor U13314 (N_13314,N_12701,N_12603);
or U13315 (N_13315,N_12508,N_12368);
or U13316 (N_13316,N_12364,N_12884);
and U13317 (N_13317,N_12786,N_12903);
and U13318 (N_13318,N_12630,N_12947);
xor U13319 (N_13319,N_12468,N_12381);
and U13320 (N_13320,N_12573,N_12512);
nor U13321 (N_13321,N_12444,N_12731);
nand U13322 (N_13322,N_12255,N_12636);
nand U13323 (N_13323,N_12039,N_12556);
and U13324 (N_13324,N_12302,N_12232);
and U13325 (N_13325,N_12647,N_12500);
nand U13326 (N_13326,N_12487,N_12238);
nor U13327 (N_13327,N_12211,N_12964);
nor U13328 (N_13328,N_12846,N_12539);
or U13329 (N_13329,N_12201,N_12557);
or U13330 (N_13330,N_12186,N_12915);
xnor U13331 (N_13331,N_12917,N_12564);
nand U13332 (N_13332,N_12060,N_12589);
or U13333 (N_13333,N_12420,N_12431);
or U13334 (N_13334,N_12712,N_12661);
and U13335 (N_13335,N_12541,N_12963);
and U13336 (N_13336,N_12146,N_12493);
or U13337 (N_13337,N_12983,N_12752);
or U13338 (N_13338,N_12689,N_12405);
and U13339 (N_13339,N_12870,N_12853);
or U13340 (N_13340,N_12339,N_12818);
nand U13341 (N_13341,N_12312,N_12515);
nand U13342 (N_13342,N_12447,N_12730);
and U13343 (N_13343,N_12914,N_12194);
nor U13344 (N_13344,N_12069,N_12953);
nor U13345 (N_13345,N_12942,N_12595);
nand U13346 (N_13346,N_12670,N_12607);
nand U13347 (N_13347,N_12358,N_12547);
nor U13348 (N_13348,N_12490,N_12671);
nor U13349 (N_13349,N_12319,N_12030);
nor U13350 (N_13350,N_12132,N_12900);
xor U13351 (N_13351,N_12592,N_12425);
nor U13352 (N_13352,N_12271,N_12534);
or U13353 (N_13353,N_12335,N_12971);
nand U13354 (N_13354,N_12948,N_12621);
or U13355 (N_13355,N_12743,N_12707);
nor U13356 (N_13356,N_12247,N_12482);
or U13357 (N_13357,N_12343,N_12967);
and U13358 (N_13358,N_12323,N_12277);
nor U13359 (N_13359,N_12221,N_12018);
nand U13360 (N_13360,N_12739,N_12196);
nand U13361 (N_13361,N_12489,N_12445);
nand U13362 (N_13362,N_12688,N_12433);
or U13363 (N_13363,N_12084,N_12443);
or U13364 (N_13364,N_12441,N_12458);
and U13365 (N_13365,N_12956,N_12926);
nor U13366 (N_13366,N_12392,N_12154);
or U13367 (N_13367,N_12020,N_12424);
or U13368 (N_13368,N_12980,N_12869);
nor U13369 (N_13369,N_12859,N_12090);
nand U13370 (N_13370,N_12697,N_12089);
or U13371 (N_13371,N_12334,N_12153);
xnor U13372 (N_13372,N_12826,N_12666);
nand U13373 (N_13373,N_12509,N_12989);
or U13374 (N_13374,N_12742,N_12456);
or U13375 (N_13375,N_12147,N_12526);
nand U13376 (N_13376,N_12583,N_12102);
nor U13377 (N_13377,N_12848,N_12242);
or U13378 (N_13378,N_12450,N_12165);
and U13379 (N_13379,N_12198,N_12883);
nor U13380 (N_13380,N_12422,N_12652);
nor U13381 (N_13381,N_12360,N_12618);
nor U13382 (N_13382,N_12735,N_12580);
or U13383 (N_13383,N_12156,N_12844);
and U13384 (N_13384,N_12212,N_12710);
nor U13385 (N_13385,N_12160,N_12403);
nand U13386 (N_13386,N_12106,N_12395);
nor U13387 (N_13387,N_12995,N_12740);
xnor U13388 (N_13388,N_12288,N_12430);
nor U13389 (N_13389,N_12359,N_12007);
nand U13390 (N_13390,N_12741,N_12372);
nand U13391 (N_13391,N_12804,N_12796);
or U13392 (N_13392,N_12311,N_12005);
nor U13393 (N_13393,N_12857,N_12823);
nand U13394 (N_13394,N_12987,N_12824);
nand U13395 (N_13395,N_12668,N_12663);
nor U13396 (N_13396,N_12055,N_12950);
nand U13397 (N_13397,N_12516,N_12297);
and U13398 (N_13398,N_12412,N_12943);
or U13399 (N_13399,N_12692,N_12643);
or U13400 (N_13400,N_12708,N_12797);
nand U13401 (N_13401,N_12774,N_12972);
or U13402 (N_13402,N_12975,N_12131);
or U13403 (N_13403,N_12021,N_12672);
and U13404 (N_13404,N_12278,N_12393);
and U13405 (N_13405,N_12822,N_12270);
nand U13406 (N_13406,N_12932,N_12593);
nand U13407 (N_13407,N_12124,N_12568);
or U13408 (N_13408,N_12933,N_12998);
nor U13409 (N_13409,N_12176,N_12472);
and U13410 (N_13410,N_12878,N_12120);
nor U13411 (N_13411,N_12905,N_12063);
and U13412 (N_13412,N_12031,N_12910);
nand U13413 (N_13413,N_12219,N_12225);
or U13414 (N_13414,N_12438,N_12862);
and U13415 (N_13415,N_12380,N_12182);
or U13416 (N_13416,N_12044,N_12142);
and U13417 (N_13417,N_12940,N_12434);
or U13418 (N_13418,N_12528,N_12050);
or U13419 (N_13419,N_12414,N_12890);
and U13420 (N_13420,N_12236,N_12075);
nor U13421 (N_13421,N_12843,N_12296);
nor U13422 (N_13422,N_12505,N_12946);
and U13423 (N_13423,N_12144,N_12762);
xnor U13424 (N_13424,N_12538,N_12649);
or U13425 (N_13425,N_12725,N_12788);
and U13426 (N_13426,N_12653,N_12909);
and U13427 (N_13427,N_12828,N_12022);
or U13428 (N_13428,N_12576,N_12982);
nand U13429 (N_13429,N_12399,N_12299);
or U13430 (N_13430,N_12204,N_12760);
nand U13431 (N_13431,N_12012,N_12977);
and U13432 (N_13432,N_12155,N_12268);
and U13433 (N_13433,N_12702,N_12137);
or U13434 (N_13434,N_12098,N_12966);
nand U13435 (N_13435,N_12811,N_12289);
or U13436 (N_13436,N_12962,N_12469);
and U13437 (N_13437,N_12704,N_12887);
nand U13438 (N_13438,N_12784,N_12690);
nand U13439 (N_13439,N_12449,N_12100);
or U13440 (N_13440,N_12761,N_12474);
nand U13441 (N_13441,N_12175,N_12460);
nand U13442 (N_13442,N_12889,N_12402);
and U13443 (N_13443,N_12755,N_12751);
or U13444 (N_13444,N_12955,N_12642);
nand U13445 (N_13445,N_12082,N_12986);
nand U13446 (N_13446,N_12789,N_12810);
or U13447 (N_13447,N_12597,N_12912);
or U13448 (N_13448,N_12825,N_12078);
nor U13449 (N_13449,N_12123,N_12228);
nand U13450 (N_13450,N_12370,N_12812);
and U13451 (N_13451,N_12484,N_12240);
nand U13452 (N_13452,N_12351,N_12927);
nor U13453 (N_13453,N_12705,N_12591);
or U13454 (N_13454,N_12540,N_12118);
nand U13455 (N_13455,N_12632,N_12918);
xnor U13456 (N_13456,N_12193,N_12285);
nor U13457 (N_13457,N_12879,N_12223);
nand U13458 (N_13458,N_12128,N_12993);
or U13459 (N_13459,N_12817,N_12958);
nand U13460 (N_13460,N_12256,N_12389);
and U13461 (N_13461,N_12072,N_12333);
nor U13462 (N_13462,N_12321,N_12227);
or U13463 (N_13463,N_12052,N_12008);
nand U13464 (N_13464,N_12362,N_12833);
and U13465 (N_13465,N_12957,N_12976);
nand U13466 (N_13466,N_12284,N_12737);
nor U13467 (N_13467,N_12925,N_12819);
xnor U13468 (N_13468,N_12188,N_12200);
nor U13469 (N_13469,N_12400,N_12292);
nand U13470 (N_13470,N_12000,N_12815);
and U13471 (N_13471,N_12615,N_12411);
nor U13472 (N_13472,N_12379,N_12218);
or U13473 (N_13473,N_12799,N_12006);
nor U13474 (N_13474,N_12027,N_12369);
nor U13475 (N_13475,N_12785,N_12941);
and U13476 (N_13476,N_12807,N_12960);
or U13477 (N_13477,N_12798,N_12733);
and U13478 (N_13478,N_12356,N_12638);
and U13479 (N_13479,N_12871,N_12139);
or U13480 (N_13480,N_12954,N_12776);
and U13481 (N_13481,N_12254,N_12095);
nand U13482 (N_13482,N_12357,N_12234);
and U13483 (N_13483,N_12477,N_12703);
and U13484 (N_13484,N_12877,N_12452);
nand U13485 (N_13485,N_12122,N_12396);
or U13486 (N_13486,N_12588,N_12531);
and U13487 (N_13487,N_12300,N_12753);
or U13488 (N_13488,N_12355,N_12525);
nand U13489 (N_13489,N_12327,N_12613);
xnor U13490 (N_13490,N_12047,N_12658);
nor U13491 (N_13491,N_12111,N_12309);
and U13492 (N_13492,N_12056,N_12239);
or U13493 (N_13493,N_12496,N_12802);
or U13494 (N_13494,N_12287,N_12079);
xnor U13495 (N_13495,N_12945,N_12736);
nand U13496 (N_13496,N_12835,N_12631);
and U13497 (N_13497,N_12858,N_12476);
nand U13498 (N_13498,N_12220,N_12575);
and U13499 (N_13499,N_12454,N_12479);
and U13500 (N_13500,N_12344,N_12590);
and U13501 (N_13501,N_12900,N_12423);
xnor U13502 (N_13502,N_12474,N_12635);
nand U13503 (N_13503,N_12642,N_12640);
nor U13504 (N_13504,N_12664,N_12599);
nand U13505 (N_13505,N_12982,N_12892);
nor U13506 (N_13506,N_12892,N_12920);
and U13507 (N_13507,N_12079,N_12532);
nor U13508 (N_13508,N_12603,N_12721);
nor U13509 (N_13509,N_12726,N_12226);
nor U13510 (N_13510,N_12076,N_12297);
nor U13511 (N_13511,N_12339,N_12077);
nand U13512 (N_13512,N_12843,N_12090);
nand U13513 (N_13513,N_12585,N_12545);
or U13514 (N_13514,N_12910,N_12458);
or U13515 (N_13515,N_12094,N_12849);
nor U13516 (N_13516,N_12608,N_12023);
or U13517 (N_13517,N_12906,N_12871);
or U13518 (N_13518,N_12420,N_12097);
nand U13519 (N_13519,N_12250,N_12566);
or U13520 (N_13520,N_12396,N_12704);
and U13521 (N_13521,N_12391,N_12315);
nor U13522 (N_13522,N_12338,N_12427);
and U13523 (N_13523,N_12252,N_12834);
nor U13524 (N_13524,N_12008,N_12312);
and U13525 (N_13525,N_12147,N_12291);
nor U13526 (N_13526,N_12948,N_12683);
nand U13527 (N_13527,N_12276,N_12895);
and U13528 (N_13528,N_12015,N_12672);
nand U13529 (N_13529,N_12153,N_12690);
nor U13530 (N_13530,N_12542,N_12858);
or U13531 (N_13531,N_12946,N_12174);
nand U13532 (N_13532,N_12971,N_12375);
and U13533 (N_13533,N_12272,N_12643);
or U13534 (N_13534,N_12732,N_12644);
and U13535 (N_13535,N_12382,N_12800);
and U13536 (N_13536,N_12549,N_12037);
or U13537 (N_13537,N_12960,N_12127);
nor U13538 (N_13538,N_12864,N_12715);
and U13539 (N_13539,N_12131,N_12958);
and U13540 (N_13540,N_12742,N_12079);
nor U13541 (N_13541,N_12981,N_12839);
or U13542 (N_13542,N_12764,N_12218);
and U13543 (N_13543,N_12893,N_12937);
or U13544 (N_13544,N_12851,N_12439);
xnor U13545 (N_13545,N_12285,N_12713);
nand U13546 (N_13546,N_12457,N_12034);
nand U13547 (N_13547,N_12780,N_12351);
or U13548 (N_13548,N_12935,N_12076);
or U13549 (N_13549,N_12011,N_12889);
or U13550 (N_13550,N_12055,N_12045);
and U13551 (N_13551,N_12935,N_12093);
or U13552 (N_13552,N_12332,N_12047);
and U13553 (N_13553,N_12023,N_12155);
and U13554 (N_13554,N_12415,N_12471);
nor U13555 (N_13555,N_12489,N_12881);
and U13556 (N_13556,N_12215,N_12535);
nor U13557 (N_13557,N_12167,N_12071);
nor U13558 (N_13558,N_12492,N_12948);
or U13559 (N_13559,N_12208,N_12165);
xor U13560 (N_13560,N_12770,N_12171);
nand U13561 (N_13561,N_12296,N_12020);
nand U13562 (N_13562,N_12461,N_12146);
xor U13563 (N_13563,N_12397,N_12765);
and U13564 (N_13564,N_12393,N_12312);
nand U13565 (N_13565,N_12036,N_12460);
nor U13566 (N_13566,N_12362,N_12280);
nand U13567 (N_13567,N_12741,N_12661);
nand U13568 (N_13568,N_12489,N_12141);
and U13569 (N_13569,N_12257,N_12406);
nand U13570 (N_13570,N_12745,N_12244);
and U13571 (N_13571,N_12822,N_12725);
xnor U13572 (N_13572,N_12212,N_12253);
and U13573 (N_13573,N_12129,N_12498);
nor U13574 (N_13574,N_12197,N_12190);
xor U13575 (N_13575,N_12683,N_12254);
or U13576 (N_13576,N_12944,N_12213);
nand U13577 (N_13577,N_12376,N_12206);
or U13578 (N_13578,N_12886,N_12725);
xor U13579 (N_13579,N_12867,N_12593);
nand U13580 (N_13580,N_12377,N_12753);
nand U13581 (N_13581,N_12177,N_12741);
nand U13582 (N_13582,N_12908,N_12817);
nor U13583 (N_13583,N_12543,N_12404);
and U13584 (N_13584,N_12407,N_12011);
xor U13585 (N_13585,N_12996,N_12859);
nand U13586 (N_13586,N_12176,N_12213);
nand U13587 (N_13587,N_12023,N_12379);
or U13588 (N_13588,N_12830,N_12227);
and U13589 (N_13589,N_12012,N_12127);
xnor U13590 (N_13590,N_12261,N_12500);
nor U13591 (N_13591,N_12910,N_12836);
and U13592 (N_13592,N_12710,N_12656);
and U13593 (N_13593,N_12367,N_12501);
or U13594 (N_13594,N_12049,N_12803);
and U13595 (N_13595,N_12011,N_12079);
nand U13596 (N_13596,N_12474,N_12969);
nor U13597 (N_13597,N_12277,N_12081);
nor U13598 (N_13598,N_12894,N_12572);
and U13599 (N_13599,N_12555,N_12380);
nor U13600 (N_13600,N_12855,N_12012);
nor U13601 (N_13601,N_12978,N_12001);
or U13602 (N_13602,N_12754,N_12382);
and U13603 (N_13603,N_12890,N_12816);
or U13604 (N_13604,N_12378,N_12505);
nand U13605 (N_13605,N_12185,N_12166);
nor U13606 (N_13606,N_12965,N_12614);
or U13607 (N_13607,N_12596,N_12186);
nand U13608 (N_13608,N_12262,N_12781);
xnor U13609 (N_13609,N_12577,N_12614);
nand U13610 (N_13610,N_12537,N_12237);
or U13611 (N_13611,N_12912,N_12583);
and U13612 (N_13612,N_12278,N_12114);
xnor U13613 (N_13613,N_12092,N_12367);
nor U13614 (N_13614,N_12287,N_12604);
or U13615 (N_13615,N_12559,N_12950);
nand U13616 (N_13616,N_12814,N_12671);
and U13617 (N_13617,N_12127,N_12278);
nand U13618 (N_13618,N_12309,N_12672);
nor U13619 (N_13619,N_12347,N_12665);
and U13620 (N_13620,N_12452,N_12747);
and U13621 (N_13621,N_12614,N_12362);
or U13622 (N_13622,N_12895,N_12903);
or U13623 (N_13623,N_12229,N_12659);
and U13624 (N_13624,N_12754,N_12787);
nand U13625 (N_13625,N_12430,N_12829);
nand U13626 (N_13626,N_12859,N_12620);
nor U13627 (N_13627,N_12462,N_12068);
xor U13628 (N_13628,N_12356,N_12333);
nand U13629 (N_13629,N_12599,N_12340);
nand U13630 (N_13630,N_12246,N_12830);
or U13631 (N_13631,N_12961,N_12552);
nor U13632 (N_13632,N_12286,N_12108);
nand U13633 (N_13633,N_12433,N_12845);
nand U13634 (N_13634,N_12388,N_12439);
nand U13635 (N_13635,N_12204,N_12692);
xor U13636 (N_13636,N_12421,N_12997);
and U13637 (N_13637,N_12409,N_12431);
xor U13638 (N_13638,N_12464,N_12881);
and U13639 (N_13639,N_12337,N_12359);
or U13640 (N_13640,N_12369,N_12097);
nand U13641 (N_13641,N_12170,N_12364);
nor U13642 (N_13642,N_12920,N_12709);
and U13643 (N_13643,N_12806,N_12688);
nor U13644 (N_13644,N_12252,N_12268);
nor U13645 (N_13645,N_12527,N_12954);
nor U13646 (N_13646,N_12168,N_12580);
and U13647 (N_13647,N_12086,N_12704);
or U13648 (N_13648,N_12163,N_12383);
nand U13649 (N_13649,N_12115,N_12475);
and U13650 (N_13650,N_12141,N_12568);
or U13651 (N_13651,N_12256,N_12281);
or U13652 (N_13652,N_12243,N_12830);
nand U13653 (N_13653,N_12231,N_12057);
and U13654 (N_13654,N_12980,N_12711);
or U13655 (N_13655,N_12761,N_12905);
nand U13656 (N_13656,N_12098,N_12007);
or U13657 (N_13657,N_12559,N_12845);
nand U13658 (N_13658,N_12560,N_12805);
or U13659 (N_13659,N_12974,N_12571);
or U13660 (N_13660,N_12119,N_12665);
or U13661 (N_13661,N_12360,N_12565);
nand U13662 (N_13662,N_12765,N_12023);
and U13663 (N_13663,N_12230,N_12592);
nand U13664 (N_13664,N_12254,N_12473);
nand U13665 (N_13665,N_12584,N_12297);
nor U13666 (N_13666,N_12870,N_12129);
and U13667 (N_13667,N_12504,N_12850);
nand U13668 (N_13668,N_12109,N_12323);
nand U13669 (N_13669,N_12284,N_12670);
and U13670 (N_13670,N_12398,N_12513);
or U13671 (N_13671,N_12566,N_12141);
or U13672 (N_13672,N_12732,N_12808);
nor U13673 (N_13673,N_12936,N_12931);
or U13674 (N_13674,N_12031,N_12129);
or U13675 (N_13675,N_12363,N_12591);
nand U13676 (N_13676,N_12274,N_12691);
or U13677 (N_13677,N_12182,N_12073);
and U13678 (N_13678,N_12115,N_12436);
nand U13679 (N_13679,N_12210,N_12848);
and U13680 (N_13680,N_12780,N_12309);
nand U13681 (N_13681,N_12825,N_12989);
and U13682 (N_13682,N_12192,N_12446);
or U13683 (N_13683,N_12705,N_12209);
and U13684 (N_13684,N_12800,N_12774);
or U13685 (N_13685,N_12936,N_12532);
or U13686 (N_13686,N_12646,N_12832);
nand U13687 (N_13687,N_12312,N_12699);
and U13688 (N_13688,N_12309,N_12698);
nor U13689 (N_13689,N_12555,N_12092);
nor U13690 (N_13690,N_12949,N_12358);
nand U13691 (N_13691,N_12288,N_12274);
or U13692 (N_13692,N_12430,N_12109);
nor U13693 (N_13693,N_12509,N_12065);
or U13694 (N_13694,N_12985,N_12476);
or U13695 (N_13695,N_12960,N_12652);
nand U13696 (N_13696,N_12737,N_12170);
nor U13697 (N_13697,N_12209,N_12902);
nand U13698 (N_13698,N_12897,N_12492);
nand U13699 (N_13699,N_12879,N_12374);
nor U13700 (N_13700,N_12963,N_12095);
or U13701 (N_13701,N_12047,N_12049);
nor U13702 (N_13702,N_12092,N_12554);
nor U13703 (N_13703,N_12927,N_12263);
nand U13704 (N_13704,N_12171,N_12472);
nand U13705 (N_13705,N_12727,N_12836);
nor U13706 (N_13706,N_12699,N_12494);
and U13707 (N_13707,N_12030,N_12908);
nand U13708 (N_13708,N_12606,N_12930);
nand U13709 (N_13709,N_12504,N_12806);
and U13710 (N_13710,N_12761,N_12096);
or U13711 (N_13711,N_12381,N_12782);
or U13712 (N_13712,N_12419,N_12277);
xor U13713 (N_13713,N_12788,N_12870);
or U13714 (N_13714,N_12002,N_12359);
and U13715 (N_13715,N_12724,N_12932);
nand U13716 (N_13716,N_12030,N_12845);
nor U13717 (N_13717,N_12760,N_12730);
or U13718 (N_13718,N_12279,N_12016);
nand U13719 (N_13719,N_12091,N_12362);
xnor U13720 (N_13720,N_12953,N_12229);
or U13721 (N_13721,N_12242,N_12860);
nor U13722 (N_13722,N_12673,N_12568);
and U13723 (N_13723,N_12110,N_12938);
and U13724 (N_13724,N_12414,N_12352);
nand U13725 (N_13725,N_12177,N_12232);
and U13726 (N_13726,N_12779,N_12116);
nand U13727 (N_13727,N_12703,N_12990);
nand U13728 (N_13728,N_12388,N_12921);
nor U13729 (N_13729,N_12229,N_12818);
or U13730 (N_13730,N_12461,N_12642);
or U13731 (N_13731,N_12153,N_12702);
and U13732 (N_13732,N_12758,N_12310);
nor U13733 (N_13733,N_12115,N_12533);
nor U13734 (N_13734,N_12409,N_12226);
and U13735 (N_13735,N_12137,N_12493);
or U13736 (N_13736,N_12806,N_12844);
or U13737 (N_13737,N_12815,N_12066);
nor U13738 (N_13738,N_12725,N_12438);
and U13739 (N_13739,N_12370,N_12012);
and U13740 (N_13740,N_12173,N_12392);
and U13741 (N_13741,N_12500,N_12481);
or U13742 (N_13742,N_12454,N_12079);
or U13743 (N_13743,N_12798,N_12709);
nor U13744 (N_13744,N_12755,N_12564);
nand U13745 (N_13745,N_12546,N_12236);
or U13746 (N_13746,N_12203,N_12534);
or U13747 (N_13747,N_12909,N_12384);
and U13748 (N_13748,N_12386,N_12494);
xor U13749 (N_13749,N_12781,N_12275);
and U13750 (N_13750,N_12740,N_12405);
or U13751 (N_13751,N_12213,N_12836);
nand U13752 (N_13752,N_12536,N_12341);
or U13753 (N_13753,N_12869,N_12222);
xor U13754 (N_13754,N_12606,N_12783);
nand U13755 (N_13755,N_12946,N_12362);
and U13756 (N_13756,N_12245,N_12406);
nand U13757 (N_13757,N_12824,N_12042);
nor U13758 (N_13758,N_12838,N_12411);
xor U13759 (N_13759,N_12474,N_12657);
nand U13760 (N_13760,N_12022,N_12519);
nor U13761 (N_13761,N_12687,N_12843);
xor U13762 (N_13762,N_12310,N_12922);
or U13763 (N_13763,N_12007,N_12866);
and U13764 (N_13764,N_12117,N_12281);
and U13765 (N_13765,N_12034,N_12531);
or U13766 (N_13766,N_12016,N_12213);
nand U13767 (N_13767,N_12925,N_12437);
and U13768 (N_13768,N_12683,N_12646);
nor U13769 (N_13769,N_12005,N_12331);
nor U13770 (N_13770,N_12090,N_12296);
or U13771 (N_13771,N_12525,N_12646);
nor U13772 (N_13772,N_12489,N_12058);
nor U13773 (N_13773,N_12752,N_12878);
or U13774 (N_13774,N_12594,N_12878);
xor U13775 (N_13775,N_12302,N_12398);
and U13776 (N_13776,N_12208,N_12925);
nor U13777 (N_13777,N_12464,N_12792);
or U13778 (N_13778,N_12899,N_12593);
nand U13779 (N_13779,N_12899,N_12809);
nand U13780 (N_13780,N_12278,N_12475);
xnor U13781 (N_13781,N_12381,N_12813);
xnor U13782 (N_13782,N_12625,N_12797);
or U13783 (N_13783,N_12827,N_12537);
or U13784 (N_13784,N_12752,N_12774);
and U13785 (N_13785,N_12141,N_12859);
nor U13786 (N_13786,N_12634,N_12749);
or U13787 (N_13787,N_12727,N_12445);
nand U13788 (N_13788,N_12296,N_12340);
or U13789 (N_13789,N_12812,N_12085);
nor U13790 (N_13790,N_12496,N_12965);
and U13791 (N_13791,N_12835,N_12716);
xor U13792 (N_13792,N_12639,N_12987);
or U13793 (N_13793,N_12872,N_12909);
xnor U13794 (N_13794,N_12466,N_12170);
nand U13795 (N_13795,N_12611,N_12330);
xor U13796 (N_13796,N_12656,N_12022);
and U13797 (N_13797,N_12001,N_12950);
or U13798 (N_13798,N_12160,N_12279);
or U13799 (N_13799,N_12581,N_12224);
nand U13800 (N_13800,N_12163,N_12002);
nand U13801 (N_13801,N_12063,N_12642);
nand U13802 (N_13802,N_12706,N_12457);
or U13803 (N_13803,N_12405,N_12706);
and U13804 (N_13804,N_12718,N_12265);
nand U13805 (N_13805,N_12093,N_12183);
nor U13806 (N_13806,N_12037,N_12334);
and U13807 (N_13807,N_12309,N_12372);
and U13808 (N_13808,N_12626,N_12446);
nor U13809 (N_13809,N_12719,N_12677);
and U13810 (N_13810,N_12653,N_12941);
nand U13811 (N_13811,N_12604,N_12936);
or U13812 (N_13812,N_12491,N_12489);
and U13813 (N_13813,N_12241,N_12059);
or U13814 (N_13814,N_12809,N_12215);
nand U13815 (N_13815,N_12415,N_12467);
xor U13816 (N_13816,N_12699,N_12803);
and U13817 (N_13817,N_12490,N_12721);
and U13818 (N_13818,N_12517,N_12181);
nand U13819 (N_13819,N_12904,N_12691);
nand U13820 (N_13820,N_12790,N_12163);
nor U13821 (N_13821,N_12836,N_12934);
xnor U13822 (N_13822,N_12118,N_12765);
and U13823 (N_13823,N_12895,N_12142);
and U13824 (N_13824,N_12346,N_12022);
xor U13825 (N_13825,N_12474,N_12992);
nand U13826 (N_13826,N_12453,N_12432);
nand U13827 (N_13827,N_12766,N_12857);
nand U13828 (N_13828,N_12968,N_12322);
nand U13829 (N_13829,N_12213,N_12362);
or U13830 (N_13830,N_12536,N_12882);
nand U13831 (N_13831,N_12505,N_12208);
or U13832 (N_13832,N_12899,N_12559);
nand U13833 (N_13833,N_12798,N_12037);
or U13834 (N_13834,N_12818,N_12630);
or U13835 (N_13835,N_12318,N_12802);
nand U13836 (N_13836,N_12225,N_12402);
or U13837 (N_13837,N_12681,N_12876);
nor U13838 (N_13838,N_12740,N_12071);
and U13839 (N_13839,N_12989,N_12503);
and U13840 (N_13840,N_12170,N_12234);
xor U13841 (N_13841,N_12073,N_12751);
nand U13842 (N_13842,N_12352,N_12612);
nor U13843 (N_13843,N_12852,N_12116);
or U13844 (N_13844,N_12732,N_12395);
xnor U13845 (N_13845,N_12697,N_12894);
nor U13846 (N_13846,N_12996,N_12736);
nor U13847 (N_13847,N_12912,N_12511);
and U13848 (N_13848,N_12723,N_12456);
and U13849 (N_13849,N_12437,N_12711);
xnor U13850 (N_13850,N_12728,N_12837);
nor U13851 (N_13851,N_12637,N_12126);
nor U13852 (N_13852,N_12952,N_12690);
and U13853 (N_13853,N_12645,N_12189);
and U13854 (N_13854,N_12712,N_12903);
nand U13855 (N_13855,N_12590,N_12467);
and U13856 (N_13856,N_12278,N_12656);
nor U13857 (N_13857,N_12435,N_12473);
nand U13858 (N_13858,N_12437,N_12061);
or U13859 (N_13859,N_12601,N_12376);
nand U13860 (N_13860,N_12219,N_12091);
nand U13861 (N_13861,N_12806,N_12217);
xnor U13862 (N_13862,N_12289,N_12850);
or U13863 (N_13863,N_12407,N_12908);
and U13864 (N_13864,N_12290,N_12202);
nand U13865 (N_13865,N_12617,N_12647);
nor U13866 (N_13866,N_12306,N_12689);
nand U13867 (N_13867,N_12227,N_12057);
nand U13868 (N_13868,N_12924,N_12322);
and U13869 (N_13869,N_12034,N_12250);
xnor U13870 (N_13870,N_12254,N_12503);
and U13871 (N_13871,N_12397,N_12756);
and U13872 (N_13872,N_12235,N_12200);
nor U13873 (N_13873,N_12986,N_12074);
and U13874 (N_13874,N_12361,N_12868);
and U13875 (N_13875,N_12541,N_12248);
or U13876 (N_13876,N_12240,N_12110);
or U13877 (N_13877,N_12983,N_12137);
and U13878 (N_13878,N_12365,N_12569);
and U13879 (N_13879,N_12570,N_12286);
or U13880 (N_13880,N_12648,N_12764);
xor U13881 (N_13881,N_12952,N_12851);
or U13882 (N_13882,N_12053,N_12343);
and U13883 (N_13883,N_12468,N_12607);
and U13884 (N_13884,N_12677,N_12665);
or U13885 (N_13885,N_12124,N_12370);
nand U13886 (N_13886,N_12177,N_12878);
nor U13887 (N_13887,N_12182,N_12726);
or U13888 (N_13888,N_12812,N_12545);
or U13889 (N_13889,N_12731,N_12168);
or U13890 (N_13890,N_12068,N_12378);
and U13891 (N_13891,N_12792,N_12065);
and U13892 (N_13892,N_12351,N_12397);
nand U13893 (N_13893,N_12132,N_12971);
nor U13894 (N_13894,N_12896,N_12740);
nand U13895 (N_13895,N_12064,N_12546);
xnor U13896 (N_13896,N_12557,N_12273);
or U13897 (N_13897,N_12839,N_12062);
nor U13898 (N_13898,N_12789,N_12418);
and U13899 (N_13899,N_12549,N_12586);
or U13900 (N_13900,N_12674,N_12224);
nor U13901 (N_13901,N_12109,N_12741);
or U13902 (N_13902,N_12465,N_12670);
or U13903 (N_13903,N_12554,N_12809);
and U13904 (N_13904,N_12777,N_12127);
nor U13905 (N_13905,N_12037,N_12165);
nand U13906 (N_13906,N_12259,N_12942);
and U13907 (N_13907,N_12095,N_12056);
nand U13908 (N_13908,N_12796,N_12440);
nor U13909 (N_13909,N_12298,N_12025);
and U13910 (N_13910,N_12804,N_12061);
or U13911 (N_13911,N_12322,N_12175);
nor U13912 (N_13912,N_12644,N_12363);
and U13913 (N_13913,N_12524,N_12403);
nor U13914 (N_13914,N_12243,N_12604);
nor U13915 (N_13915,N_12979,N_12327);
or U13916 (N_13916,N_12704,N_12345);
nor U13917 (N_13917,N_12119,N_12993);
nand U13918 (N_13918,N_12695,N_12491);
and U13919 (N_13919,N_12150,N_12147);
and U13920 (N_13920,N_12565,N_12812);
nand U13921 (N_13921,N_12028,N_12224);
xnor U13922 (N_13922,N_12701,N_12168);
and U13923 (N_13923,N_12097,N_12712);
nand U13924 (N_13924,N_12481,N_12600);
nand U13925 (N_13925,N_12077,N_12491);
or U13926 (N_13926,N_12861,N_12211);
or U13927 (N_13927,N_12677,N_12968);
or U13928 (N_13928,N_12702,N_12956);
and U13929 (N_13929,N_12938,N_12102);
and U13930 (N_13930,N_12423,N_12868);
or U13931 (N_13931,N_12476,N_12411);
nor U13932 (N_13932,N_12418,N_12130);
or U13933 (N_13933,N_12480,N_12611);
nand U13934 (N_13934,N_12729,N_12393);
nand U13935 (N_13935,N_12726,N_12225);
or U13936 (N_13936,N_12704,N_12190);
and U13937 (N_13937,N_12071,N_12066);
or U13938 (N_13938,N_12890,N_12470);
or U13939 (N_13939,N_12407,N_12464);
nor U13940 (N_13940,N_12266,N_12529);
nand U13941 (N_13941,N_12285,N_12249);
xor U13942 (N_13942,N_12932,N_12805);
and U13943 (N_13943,N_12389,N_12671);
nand U13944 (N_13944,N_12173,N_12156);
or U13945 (N_13945,N_12401,N_12171);
or U13946 (N_13946,N_12453,N_12981);
nor U13947 (N_13947,N_12666,N_12231);
or U13948 (N_13948,N_12348,N_12151);
xnor U13949 (N_13949,N_12687,N_12464);
and U13950 (N_13950,N_12789,N_12142);
nor U13951 (N_13951,N_12178,N_12526);
nor U13952 (N_13952,N_12877,N_12769);
nor U13953 (N_13953,N_12170,N_12007);
and U13954 (N_13954,N_12989,N_12984);
and U13955 (N_13955,N_12361,N_12492);
nor U13956 (N_13956,N_12091,N_12636);
or U13957 (N_13957,N_12306,N_12261);
and U13958 (N_13958,N_12611,N_12936);
and U13959 (N_13959,N_12173,N_12760);
nand U13960 (N_13960,N_12863,N_12633);
and U13961 (N_13961,N_12706,N_12509);
nor U13962 (N_13962,N_12884,N_12939);
nand U13963 (N_13963,N_12284,N_12666);
or U13964 (N_13964,N_12598,N_12367);
or U13965 (N_13965,N_12640,N_12889);
or U13966 (N_13966,N_12379,N_12104);
nand U13967 (N_13967,N_12718,N_12140);
and U13968 (N_13968,N_12524,N_12834);
or U13969 (N_13969,N_12593,N_12836);
nand U13970 (N_13970,N_12120,N_12693);
nor U13971 (N_13971,N_12266,N_12556);
or U13972 (N_13972,N_12119,N_12541);
or U13973 (N_13973,N_12256,N_12483);
xnor U13974 (N_13974,N_12425,N_12431);
nand U13975 (N_13975,N_12536,N_12234);
nor U13976 (N_13976,N_12236,N_12793);
nand U13977 (N_13977,N_12989,N_12215);
and U13978 (N_13978,N_12004,N_12637);
and U13979 (N_13979,N_12789,N_12176);
nand U13980 (N_13980,N_12485,N_12300);
nor U13981 (N_13981,N_12336,N_12106);
or U13982 (N_13982,N_12842,N_12102);
and U13983 (N_13983,N_12868,N_12258);
and U13984 (N_13984,N_12533,N_12638);
nor U13985 (N_13985,N_12489,N_12512);
or U13986 (N_13986,N_12243,N_12162);
or U13987 (N_13987,N_12277,N_12175);
nor U13988 (N_13988,N_12606,N_12293);
and U13989 (N_13989,N_12741,N_12013);
nor U13990 (N_13990,N_12577,N_12344);
nor U13991 (N_13991,N_12082,N_12414);
nor U13992 (N_13992,N_12453,N_12015);
or U13993 (N_13993,N_12059,N_12462);
or U13994 (N_13994,N_12973,N_12558);
nand U13995 (N_13995,N_12589,N_12500);
and U13996 (N_13996,N_12231,N_12329);
xnor U13997 (N_13997,N_12020,N_12208);
or U13998 (N_13998,N_12908,N_12343);
or U13999 (N_13999,N_12216,N_12368);
nand U14000 (N_14000,N_13062,N_13154);
or U14001 (N_14001,N_13014,N_13173);
nand U14002 (N_14002,N_13262,N_13452);
nor U14003 (N_14003,N_13304,N_13879);
nand U14004 (N_14004,N_13116,N_13810);
nor U14005 (N_14005,N_13323,N_13573);
and U14006 (N_14006,N_13436,N_13309);
nor U14007 (N_14007,N_13583,N_13391);
nor U14008 (N_14008,N_13441,N_13887);
nand U14009 (N_14009,N_13222,N_13318);
nor U14010 (N_14010,N_13461,N_13494);
nand U14011 (N_14011,N_13900,N_13946);
and U14012 (N_14012,N_13083,N_13801);
nand U14013 (N_14013,N_13215,N_13413);
nand U14014 (N_14014,N_13431,N_13739);
nor U14015 (N_14015,N_13163,N_13827);
nor U14016 (N_14016,N_13148,N_13196);
nand U14017 (N_14017,N_13368,N_13866);
or U14018 (N_14018,N_13473,N_13036);
nor U14019 (N_14019,N_13904,N_13923);
xnor U14020 (N_14020,N_13940,N_13700);
nor U14021 (N_14021,N_13214,N_13080);
nand U14022 (N_14022,N_13628,N_13307);
nor U14023 (N_14023,N_13225,N_13563);
nand U14024 (N_14024,N_13634,N_13272);
xnor U14025 (N_14025,N_13791,N_13780);
nor U14026 (N_14026,N_13584,N_13803);
and U14027 (N_14027,N_13139,N_13496);
nor U14028 (N_14028,N_13103,N_13466);
nor U14029 (N_14029,N_13786,N_13953);
nand U14030 (N_14030,N_13269,N_13770);
nand U14031 (N_14031,N_13088,N_13102);
or U14032 (N_14032,N_13429,N_13699);
xnor U14033 (N_14033,N_13541,N_13186);
nand U14034 (N_14034,N_13144,N_13051);
nor U14035 (N_14035,N_13629,N_13329);
or U14036 (N_14036,N_13571,N_13868);
nor U14037 (N_14037,N_13426,N_13973);
nand U14038 (N_14038,N_13792,N_13212);
nand U14039 (N_14039,N_13798,N_13941);
nor U14040 (N_14040,N_13774,N_13185);
nor U14041 (N_14041,N_13005,N_13888);
nand U14042 (N_14042,N_13859,N_13901);
and U14043 (N_14043,N_13676,N_13395);
nand U14044 (N_14044,N_13048,N_13503);
or U14045 (N_14045,N_13776,N_13008);
nor U14046 (N_14046,N_13752,N_13182);
or U14047 (N_14047,N_13504,N_13680);
nor U14048 (N_14048,N_13971,N_13266);
nor U14049 (N_14049,N_13455,N_13058);
nand U14050 (N_14050,N_13811,N_13221);
and U14051 (N_14051,N_13002,N_13969);
and U14052 (N_14052,N_13821,N_13393);
or U14053 (N_14053,N_13617,N_13773);
xnor U14054 (N_14054,N_13932,N_13759);
nand U14055 (N_14055,N_13890,N_13268);
and U14056 (N_14056,N_13006,N_13814);
and U14057 (N_14057,N_13264,N_13877);
or U14058 (N_14058,N_13068,N_13790);
and U14059 (N_14059,N_13578,N_13779);
nand U14060 (N_14060,N_13709,N_13978);
xnor U14061 (N_14061,N_13302,N_13015);
and U14062 (N_14062,N_13483,N_13126);
nor U14063 (N_14063,N_13001,N_13618);
or U14064 (N_14064,N_13147,N_13647);
nor U14065 (N_14065,N_13606,N_13013);
and U14066 (N_14066,N_13576,N_13493);
xor U14067 (N_14067,N_13520,N_13511);
xor U14068 (N_14068,N_13101,N_13330);
or U14069 (N_14069,N_13097,N_13620);
nand U14070 (N_14070,N_13855,N_13374);
or U14071 (N_14071,N_13743,N_13316);
and U14072 (N_14072,N_13351,N_13366);
and U14073 (N_14073,N_13507,N_13470);
nand U14074 (N_14074,N_13767,N_13271);
and U14075 (N_14075,N_13482,N_13156);
nor U14076 (N_14076,N_13854,N_13995);
nand U14077 (N_14077,N_13254,N_13248);
xor U14078 (N_14078,N_13064,N_13050);
nor U14079 (N_14079,N_13621,N_13590);
and U14080 (N_14080,N_13771,N_13255);
or U14081 (N_14081,N_13392,N_13347);
and U14082 (N_14082,N_13909,N_13986);
nor U14083 (N_14083,N_13072,N_13108);
and U14084 (N_14084,N_13733,N_13469);
nor U14085 (N_14085,N_13242,N_13731);
or U14086 (N_14086,N_13265,N_13593);
nand U14087 (N_14087,N_13459,N_13761);
nand U14088 (N_14088,N_13555,N_13298);
nand U14089 (N_14089,N_13847,N_13554);
nor U14090 (N_14090,N_13447,N_13448);
nor U14091 (N_14091,N_13542,N_13484);
nor U14092 (N_14092,N_13105,N_13635);
and U14093 (N_14093,N_13550,N_13582);
nor U14094 (N_14094,N_13071,N_13875);
nand U14095 (N_14095,N_13960,N_13812);
nor U14096 (N_14096,N_13545,N_13913);
and U14097 (N_14097,N_13357,N_13365);
nand U14098 (N_14098,N_13870,N_13602);
nand U14099 (N_14099,N_13692,N_13694);
or U14100 (N_14100,N_13543,N_13742);
nand U14101 (N_14101,N_13894,N_13052);
xor U14102 (N_14102,N_13927,N_13527);
or U14103 (N_14103,N_13454,N_13658);
and U14104 (N_14104,N_13753,N_13586);
nand U14105 (N_14105,N_13158,N_13208);
or U14106 (N_14106,N_13976,N_13043);
nand U14107 (N_14107,N_13450,N_13518);
and U14108 (N_14108,N_13639,N_13107);
and U14109 (N_14109,N_13693,N_13853);
and U14110 (N_14110,N_13880,N_13125);
nand U14111 (N_14111,N_13138,N_13465);
and U14112 (N_14112,N_13641,N_13274);
nor U14113 (N_14113,N_13648,N_13111);
and U14114 (N_14114,N_13599,N_13835);
nand U14115 (N_14115,N_13134,N_13155);
nor U14116 (N_14116,N_13513,N_13179);
nand U14117 (N_14117,N_13200,N_13301);
nor U14118 (N_14118,N_13239,N_13028);
or U14119 (N_14119,N_13427,N_13010);
nand U14120 (N_14120,N_13980,N_13669);
or U14121 (N_14121,N_13865,N_13966);
nand U14122 (N_14122,N_13406,N_13443);
and U14123 (N_14123,N_13009,N_13831);
nor U14124 (N_14124,N_13569,N_13294);
or U14125 (N_14125,N_13460,N_13813);
and U14126 (N_14126,N_13589,N_13689);
and U14127 (N_14127,N_13420,N_13415);
or U14128 (N_14128,N_13505,N_13701);
nand U14129 (N_14129,N_13886,N_13799);
nor U14130 (N_14130,N_13174,N_13486);
nor U14131 (N_14131,N_13600,N_13964);
nand U14132 (N_14132,N_13388,N_13217);
or U14133 (N_14133,N_13491,N_13816);
or U14134 (N_14134,N_13640,N_13679);
nand U14135 (N_14135,N_13403,N_13033);
or U14136 (N_14136,N_13558,N_13710);
and U14137 (N_14137,N_13492,N_13547);
or U14138 (N_14138,N_13642,N_13345);
and U14139 (N_14139,N_13252,N_13842);
and U14140 (N_14140,N_13487,N_13556);
or U14141 (N_14141,N_13249,N_13231);
and U14142 (N_14142,N_13418,N_13416);
nand U14143 (N_14143,N_13595,N_13223);
or U14144 (N_14144,N_13777,N_13007);
nor U14145 (N_14145,N_13952,N_13588);
and U14146 (N_14146,N_13405,N_13178);
or U14147 (N_14147,N_13795,N_13757);
nand U14148 (N_14148,N_13848,N_13972);
and U14149 (N_14149,N_13346,N_13819);
nand U14150 (N_14150,N_13682,N_13018);
or U14151 (N_14151,N_13899,N_13306);
or U14152 (N_14152,N_13315,N_13678);
xor U14153 (N_14153,N_13830,N_13651);
nand U14154 (N_14154,N_13335,N_13945);
nor U14155 (N_14155,N_13142,N_13457);
or U14156 (N_14156,N_13096,N_13396);
and U14157 (N_14157,N_13871,N_13653);
nand U14158 (N_14158,N_13860,N_13191);
and U14159 (N_14159,N_13061,N_13381);
or U14160 (N_14160,N_13662,N_13749);
and U14161 (N_14161,N_13424,N_13806);
and U14162 (N_14162,N_13153,N_13261);
or U14163 (N_14163,N_13352,N_13775);
or U14164 (N_14164,N_13011,N_13224);
and U14165 (N_14165,N_13311,N_13074);
or U14166 (N_14166,N_13643,N_13611);
xnor U14167 (N_14167,N_13696,N_13402);
xnor U14168 (N_14168,N_13276,N_13688);
or U14169 (N_14169,N_13754,N_13997);
nor U14170 (N_14170,N_13082,N_13905);
nand U14171 (N_14171,N_13060,N_13591);
and U14172 (N_14172,N_13867,N_13296);
nand U14173 (N_14173,N_13442,N_13376);
xor U14174 (N_14174,N_13895,N_13979);
nor U14175 (N_14175,N_13260,N_13091);
nand U14176 (N_14176,N_13100,N_13747);
nand U14177 (N_14177,N_13146,N_13437);
or U14178 (N_14178,N_13110,N_13025);
or U14179 (N_14179,N_13862,N_13162);
and U14180 (N_14180,N_13331,N_13181);
or U14181 (N_14181,N_13516,N_13858);
nor U14182 (N_14182,N_13089,N_13120);
or U14183 (N_14183,N_13227,N_13587);
or U14184 (N_14184,N_13937,N_13884);
nor U14185 (N_14185,N_13788,N_13872);
and U14186 (N_14186,N_13857,N_13610);
nor U14187 (N_14187,N_13695,N_13324);
or U14188 (N_14188,N_13263,N_13425);
nor U14189 (N_14189,N_13724,N_13711);
and U14190 (N_14190,N_13336,N_13471);
and U14191 (N_14191,N_13526,N_13820);
and U14192 (N_14192,N_13697,N_13495);
nand U14193 (N_14193,N_13920,N_13644);
or U14194 (N_14194,N_13660,N_13737);
nor U14195 (N_14195,N_13290,N_13017);
nor U14196 (N_14196,N_13809,N_13197);
nand U14197 (N_14197,N_13565,N_13204);
or U14198 (N_14198,N_13687,N_13375);
nand U14199 (N_14199,N_13916,N_13203);
nor U14200 (N_14200,N_13029,N_13023);
and U14201 (N_14201,N_13581,N_13350);
nand U14202 (N_14202,N_13575,N_13159);
nor U14203 (N_14203,N_13671,N_13703);
nand U14204 (N_14204,N_13232,N_13519);
and U14205 (N_14205,N_13035,N_13921);
or U14206 (N_14206,N_13736,N_13444);
nand U14207 (N_14207,N_13422,N_13849);
xor U14208 (N_14208,N_13794,N_13746);
nand U14209 (N_14209,N_13414,N_13965);
xnor U14210 (N_14210,N_13480,N_13192);
xor U14211 (N_14211,N_13093,N_13510);
or U14212 (N_14212,N_13180,N_13283);
nor U14213 (N_14213,N_13822,N_13706);
or U14214 (N_14214,N_13279,N_13630);
nand U14215 (N_14215,N_13808,N_13509);
nand U14216 (N_14216,N_13579,N_13187);
nor U14217 (N_14217,N_13280,N_13213);
and U14218 (N_14218,N_13451,N_13387);
nor U14219 (N_14219,N_13053,N_13124);
nor U14220 (N_14220,N_13327,N_13299);
nor U14221 (N_14221,N_13157,N_13607);
and U14222 (N_14222,N_13218,N_13168);
xnor U14223 (N_14223,N_13852,N_13205);
or U14224 (N_14224,N_13019,N_13769);
nor U14225 (N_14225,N_13993,N_13615);
nor U14226 (N_14226,N_13656,N_13768);
nand U14227 (N_14227,N_13340,N_13065);
nand U14228 (N_14228,N_13207,N_13477);
nand U14229 (N_14229,N_13524,N_13604);
nor U14230 (N_14230,N_13004,N_13652);
xnor U14231 (N_14231,N_13898,N_13194);
or U14232 (N_14232,N_13423,N_13325);
nor U14233 (N_14233,N_13804,N_13281);
nand U14234 (N_14234,N_13650,N_13538);
nand U14235 (N_14235,N_13319,N_13490);
nor U14236 (N_14236,N_13850,N_13970);
and U14237 (N_14237,N_13807,N_13000);
and U14238 (N_14238,N_13359,N_13649);
and U14239 (N_14239,N_13531,N_13291);
xor U14240 (N_14240,N_13106,N_13975);
nand U14241 (N_14241,N_13367,N_13528);
nand U14242 (N_14242,N_13702,N_13958);
nor U14243 (N_14243,N_13672,N_13760);
or U14244 (N_14244,N_13338,N_13293);
nand U14245 (N_14245,N_13118,N_13614);
or U14246 (N_14246,N_13145,N_13715);
nand U14247 (N_14247,N_13435,N_13934);
nor U14248 (N_14248,N_13419,N_13991);
nor U14249 (N_14249,N_13836,N_13384);
or U14250 (N_14250,N_13841,N_13832);
and U14251 (N_14251,N_13383,N_13489);
nor U14252 (N_14252,N_13075,N_13161);
nand U14253 (N_14253,N_13561,N_13394);
nor U14254 (N_14254,N_13228,N_13633);
nand U14255 (N_14255,N_13517,N_13244);
and U14256 (N_14256,N_13099,N_13996);
nor U14257 (N_14257,N_13636,N_13034);
nand U14258 (N_14258,N_13627,N_13240);
nor U14259 (N_14259,N_13143,N_13479);
nand U14260 (N_14260,N_13974,N_13539);
nor U14261 (N_14261,N_13149,N_13951);
nor U14262 (N_14262,N_13674,N_13289);
nand U14263 (N_14263,N_13445,N_13499);
nor U14264 (N_14264,N_13881,N_13918);
or U14265 (N_14265,N_13559,N_13818);
or U14266 (N_14266,N_13675,N_13903);
nand U14267 (N_14267,N_13956,N_13778);
nand U14268 (N_14268,N_13401,N_13562);
nand U14269 (N_14269,N_13288,N_13536);
xor U14270 (N_14270,N_13421,N_13373);
or U14271 (N_14271,N_13341,N_13202);
xnor U14272 (N_14272,N_13121,N_13681);
and U14273 (N_14273,N_13598,N_13514);
nor U14274 (N_14274,N_13882,N_13968);
xor U14275 (N_14275,N_13521,N_13184);
or U14276 (N_14276,N_13597,N_13363);
nor U14277 (N_14277,N_13092,N_13762);
or U14278 (N_14278,N_13129,N_13928);
nand U14279 (N_14279,N_13726,N_13152);
xor U14280 (N_14280,N_13508,N_13472);
or U14281 (N_14281,N_13303,N_13123);
nor U14282 (N_14282,N_13719,N_13962);
xnor U14283 (N_14283,N_13137,N_13313);
and U14284 (N_14284,N_13988,N_13892);
xor U14285 (N_14285,N_13891,N_13021);
and U14286 (N_14286,N_13908,N_13332);
or U14287 (N_14287,N_13430,N_13532);
xnor U14288 (N_14288,N_13497,N_13704);
nor U14289 (N_14289,N_13377,N_13567);
or U14290 (N_14290,N_13580,N_13763);
and U14291 (N_14291,N_13044,N_13382);
and U14292 (N_14292,N_13308,N_13781);
xnor U14293 (N_14293,N_13128,N_13632);
and U14294 (N_14294,N_13949,N_13931);
nor U14295 (N_14295,N_13188,N_13464);
or U14296 (N_14296,N_13412,N_13049);
nor U14297 (N_14297,N_13135,N_13141);
nor U14298 (N_14298,N_13987,N_13721);
and U14299 (N_14299,N_13122,N_13467);
nor U14300 (N_14300,N_13863,N_13546);
nor U14301 (N_14301,N_13933,N_13233);
or U14302 (N_14302,N_13440,N_13716);
and U14303 (N_14303,N_13924,N_13079);
nand U14304 (N_14304,N_13344,N_13356);
or U14305 (N_14305,N_13164,N_13273);
xnor U14306 (N_14306,N_13989,N_13198);
and U14307 (N_14307,N_13646,N_13705);
and U14308 (N_14308,N_13544,N_13169);
or U14309 (N_14309,N_13055,N_13041);
and U14310 (N_14310,N_13553,N_13758);
and U14311 (N_14311,N_13284,N_13287);
xnor U14312 (N_14312,N_13312,N_13040);
or U14313 (N_14313,N_13596,N_13063);
nor U14314 (N_14314,N_13638,N_13084);
nand U14315 (N_14315,N_13211,N_13787);
and U14316 (N_14316,N_13655,N_13113);
or U14317 (N_14317,N_13201,N_13712);
nand U14318 (N_14318,N_13140,N_13399);
xnor U14319 (N_14319,N_13277,N_13684);
nand U14320 (N_14320,N_13081,N_13229);
nor U14321 (N_14321,N_13458,N_13410);
nor U14322 (N_14322,N_13119,N_13115);
nor U14323 (N_14323,N_13358,N_13286);
nand U14324 (N_14324,N_13797,N_13039);
or U14325 (N_14325,N_13474,N_13077);
nor U14326 (N_14326,N_13730,N_13557);
and U14327 (N_14327,N_13026,N_13506);
xor U14328 (N_14328,N_13906,N_13219);
nor U14329 (N_14329,N_13434,N_13237);
nor U14330 (N_14330,N_13800,N_13815);
nor U14331 (N_14331,N_13059,N_13664);
or U14332 (N_14332,N_13389,N_13167);
nor U14333 (N_14333,N_13605,N_13572);
nand U14334 (N_14334,N_13109,N_13372);
or U14335 (N_14335,N_13476,N_13755);
or U14336 (N_14336,N_13170,N_13564);
or U14337 (N_14337,N_13073,N_13723);
nor U14338 (N_14338,N_13817,N_13734);
or U14339 (N_14339,N_13825,N_13433);
nor U14340 (N_14340,N_13165,N_13275);
and U14341 (N_14341,N_13823,N_13525);
nand U14342 (N_14342,N_13210,N_13361);
nand U14343 (N_14343,N_13782,N_13612);
nor U14344 (N_14344,N_13127,N_13834);
and U14345 (N_14345,N_13876,N_13670);
nand U14346 (N_14346,N_13475,N_13560);
and U14347 (N_14347,N_13175,N_13328);
or U14348 (N_14348,N_13677,N_13744);
nor U14349 (N_14349,N_13577,N_13189);
nand U14350 (N_14350,N_13333,N_13270);
or U14351 (N_14351,N_13939,N_13177);
nand U14352 (N_14352,N_13959,N_13843);
and U14353 (N_14353,N_13257,N_13098);
xnor U14354 (N_14354,N_13585,N_13038);
or U14355 (N_14355,N_13845,N_13907);
or U14356 (N_14356,N_13086,N_13623);
and U14357 (N_14357,N_13826,N_13016);
or U14358 (N_14358,N_13805,N_13022);
xnor U14359 (N_14359,N_13378,N_13943);
nor U14360 (N_14360,N_13246,N_13666);
nand U14361 (N_14361,N_13522,N_13056);
or U14362 (N_14362,N_13343,N_13833);
and U14363 (N_14363,N_13030,N_13957);
nor U14364 (N_14364,N_13047,N_13305);
or U14365 (N_14365,N_13999,N_13603);
nand U14366 (N_14366,N_13529,N_13235);
nor U14367 (N_14367,N_13784,N_13789);
nand U14368 (N_14368,N_13369,N_13955);
or U14369 (N_14369,N_13861,N_13278);
and U14370 (N_14370,N_13717,N_13453);
nor U14371 (N_14371,N_13828,N_13171);
nand U14372 (N_14372,N_13718,N_13209);
or U14373 (N_14373,N_13772,N_13027);
nor U14374 (N_14374,N_13961,N_13873);
and U14375 (N_14375,N_13851,N_13947);
nand U14376 (N_14376,N_13117,N_13982);
nand U14377 (N_14377,N_13722,N_13824);
nand U14378 (N_14378,N_13183,N_13950);
nor U14379 (N_14379,N_13690,N_13708);
or U14380 (N_14380,N_13355,N_13478);
nor U14381 (N_14381,N_13463,N_13057);
nand U14382 (N_14382,N_13714,N_13616);
nand U14383 (N_14383,N_13728,N_13206);
nand U14384 (N_14384,N_13802,N_13915);
nand U14385 (N_14385,N_13750,N_13837);
nand U14386 (N_14386,N_13914,N_13066);
or U14387 (N_14387,N_13078,N_13929);
or U14388 (N_14388,N_13132,N_13994);
and U14389 (N_14389,N_13796,N_13902);
nor U14390 (N_14390,N_13364,N_13738);
nand U14391 (N_14391,N_13745,N_13922);
and U14392 (N_14392,N_13535,N_13613);
and U14393 (N_14393,N_13707,N_13594);
nor U14394 (N_14394,N_13321,N_13838);
nor U14395 (N_14395,N_13985,N_13253);
and U14396 (N_14396,N_13785,N_13337);
or U14397 (N_14397,N_13930,N_13151);
nand U14398 (N_14398,N_13500,N_13740);
and U14399 (N_14399,N_13216,N_13735);
or U14400 (N_14400,N_13411,N_13720);
nor U14401 (N_14401,N_13984,N_13727);
or U14402 (N_14402,N_13935,N_13530);
nor U14403 (N_14403,N_13371,N_13741);
or U14404 (N_14404,N_13574,N_13637);
and U14405 (N_14405,N_13668,N_13748);
and U14406 (N_14406,N_13462,N_13844);
and U14407 (N_14407,N_13090,N_13386);
and U14408 (N_14408,N_13468,N_13360);
nor U14409 (N_14409,N_13878,N_13896);
xor U14410 (N_14410,N_13609,N_13285);
or U14411 (N_14411,N_13258,N_13942);
nor U14412 (N_14412,N_13397,N_13334);
nand U14413 (N_14413,N_13549,N_13783);
xor U14414 (N_14414,N_13245,N_13295);
nand U14415 (N_14415,N_13267,N_13608);
or U14416 (N_14416,N_13085,N_13766);
and U14417 (N_14417,N_13398,N_13160);
nor U14418 (N_14418,N_13136,N_13874);
nor U14419 (N_14419,N_13326,N_13502);
nor U14420 (N_14420,N_13247,N_13897);
or U14421 (N_14421,N_13310,N_13515);
nor U14422 (N_14422,N_13917,N_13020);
or U14423 (N_14423,N_13626,N_13765);
or U14424 (N_14424,N_13657,N_13983);
nor U14425 (N_14425,N_13936,N_13076);
or U14426 (N_14426,N_13220,N_13501);
or U14427 (N_14427,N_13354,N_13446);
xnor U14428 (N_14428,N_13370,N_13481);
xor U14429 (N_14429,N_13300,N_13926);
nor U14430 (N_14430,N_13193,N_13869);
or U14431 (N_14431,N_13251,N_13297);
nand U14432 (N_14432,N_13534,N_13069);
xnor U14433 (N_14433,N_13981,N_13840);
or U14434 (N_14434,N_13439,N_13938);
nand U14435 (N_14435,N_13348,N_13732);
and U14436 (N_14436,N_13320,N_13856);
nor U14437 (N_14437,N_13911,N_13764);
xnor U14438 (N_14438,N_13967,N_13150);
and U14439 (N_14439,N_13087,N_13665);
xnor U14440 (N_14440,N_13339,N_13130);
or U14441 (N_14441,N_13977,N_13889);
nand U14442 (N_14442,N_13686,N_13659);
nor U14443 (N_14443,N_13751,N_13551);
or U14444 (N_14444,N_13417,N_13012);
and U14445 (N_14445,N_13485,N_13238);
nor U14446 (N_14446,N_13408,N_13654);
or U14447 (N_14447,N_13166,N_13725);
or U14448 (N_14448,N_13864,N_13176);
nand U14449 (N_14449,N_13380,N_13133);
or U14450 (N_14450,N_13404,N_13432);
nand U14451 (N_14451,N_13568,N_13846);
nand U14452 (N_14452,N_13428,N_13488);
and U14453 (N_14453,N_13910,N_13456);
and U14454 (N_14454,N_13954,N_13046);
or U14455 (N_14455,N_13661,N_13234);
xor U14456 (N_14456,N_13282,N_13362);
nor U14457 (N_14457,N_13031,N_13314);
or U14458 (N_14458,N_13195,N_13512);
nor U14459 (N_14459,N_13552,N_13230);
nand U14460 (N_14460,N_13292,N_13990);
nor U14461 (N_14461,N_13243,N_13112);
or U14462 (N_14462,N_13683,N_13925);
xnor U14463 (N_14463,N_13349,N_13131);
and U14464 (N_14464,N_13172,N_13685);
nor U14465 (N_14465,N_13663,N_13948);
and U14466 (N_14466,N_13645,N_13998);
xnor U14467 (N_14467,N_13400,N_13003);
nor U14468 (N_14468,N_13523,N_13793);
nor U14469 (N_14469,N_13094,N_13624);
nand U14470 (N_14470,N_13104,N_13631);
nand U14471 (N_14471,N_13037,N_13667);
nor U14472 (N_14472,N_13095,N_13409);
or U14473 (N_14473,N_13045,N_13673);
and U14474 (N_14474,N_13619,N_13498);
nor U14475 (N_14475,N_13625,N_13548);
nor U14476 (N_14476,N_13829,N_13407);
nor U14477 (N_14477,N_13067,N_13566);
nand U14478 (N_14478,N_13114,N_13944);
or U14479 (N_14479,N_13912,N_13893);
and U14480 (N_14480,N_13601,N_13317);
or U14481 (N_14481,N_13024,N_13390);
nand U14482 (N_14482,N_13226,N_13713);
or U14483 (N_14483,N_13592,N_13729);
or U14484 (N_14484,N_13241,N_13698);
or U14485 (N_14485,N_13622,N_13438);
nor U14486 (N_14486,N_13199,N_13054);
and U14487 (N_14487,N_13236,N_13883);
and U14488 (N_14488,N_13919,N_13070);
nor U14489 (N_14489,N_13533,N_13385);
and U14490 (N_14490,N_13042,N_13256);
nand U14491 (N_14491,N_13540,N_13570);
nand U14492 (N_14492,N_13379,N_13190);
nand U14493 (N_14493,N_13250,N_13885);
nand U14494 (N_14494,N_13537,N_13449);
nor U14495 (N_14495,N_13032,N_13259);
xnor U14496 (N_14496,N_13342,N_13322);
nand U14497 (N_14497,N_13992,N_13839);
or U14498 (N_14498,N_13963,N_13756);
nor U14499 (N_14499,N_13691,N_13353);
nand U14500 (N_14500,N_13767,N_13233);
nor U14501 (N_14501,N_13993,N_13837);
and U14502 (N_14502,N_13021,N_13289);
nor U14503 (N_14503,N_13428,N_13517);
and U14504 (N_14504,N_13466,N_13606);
xor U14505 (N_14505,N_13830,N_13088);
nand U14506 (N_14506,N_13383,N_13499);
and U14507 (N_14507,N_13464,N_13240);
nand U14508 (N_14508,N_13294,N_13394);
or U14509 (N_14509,N_13631,N_13126);
xor U14510 (N_14510,N_13833,N_13557);
nand U14511 (N_14511,N_13089,N_13719);
and U14512 (N_14512,N_13070,N_13218);
nand U14513 (N_14513,N_13211,N_13621);
nand U14514 (N_14514,N_13844,N_13930);
and U14515 (N_14515,N_13545,N_13992);
nor U14516 (N_14516,N_13314,N_13391);
or U14517 (N_14517,N_13045,N_13718);
or U14518 (N_14518,N_13212,N_13065);
and U14519 (N_14519,N_13211,N_13055);
nand U14520 (N_14520,N_13527,N_13529);
nand U14521 (N_14521,N_13454,N_13697);
or U14522 (N_14522,N_13080,N_13497);
nand U14523 (N_14523,N_13206,N_13140);
nor U14524 (N_14524,N_13876,N_13258);
or U14525 (N_14525,N_13864,N_13642);
nor U14526 (N_14526,N_13989,N_13431);
or U14527 (N_14527,N_13729,N_13388);
nand U14528 (N_14528,N_13488,N_13318);
or U14529 (N_14529,N_13743,N_13239);
or U14530 (N_14530,N_13579,N_13359);
and U14531 (N_14531,N_13991,N_13754);
nor U14532 (N_14532,N_13522,N_13726);
nand U14533 (N_14533,N_13396,N_13246);
nand U14534 (N_14534,N_13601,N_13120);
or U14535 (N_14535,N_13172,N_13800);
nor U14536 (N_14536,N_13036,N_13414);
nand U14537 (N_14537,N_13709,N_13710);
or U14538 (N_14538,N_13927,N_13238);
xnor U14539 (N_14539,N_13482,N_13580);
and U14540 (N_14540,N_13160,N_13144);
nor U14541 (N_14541,N_13168,N_13599);
nand U14542 (N_14542,N_13423,N_13076);
nor U14543 (N_14543,N_13339,N_13321);
or U14544 (N_14544,N_13498,N_13394);
and U14545 (N_14545,N_13450,N_13220);
and U14546 (N_14546,N_13087,N_13041);
and U14547 (N_14547,N_13687,N_13103);
nor U14548 (N_14548,N_13890,N_13373);
xnor U14549 (N_14549,N_13676,N_13944);
nand U14550 (N_14550,N_13040,N_13916);
nand U14551 (N_14551,N_13867,N_13670);
nand U14552 (N_14552,N_13403,N_13035);
nand U14553 (N_14553,N_13053,N_13890);
nor U14554 (N_14554,N_13696,N_13350);
nand U14555 (N_14555,N_13003,N_13601);
nand U14556 (N_14556,N_13015,N_13489);
nor U14557 (N_14557,N_13229,N_13862);
and U14558 (N_14558,N_13164,N_13430);
or U14559 (N_14559,N_13974,N_13858);
nand U14560 (N_14560,N_13912,N_13131);
or U14561 (N_14561,N_13125,N_13138);
nand U14562 (N_14562,N_13926,N_13058);
nand U14563 (N_14563,N_13956,N_13570);
and U14564 (N_14564,N_13626,N_13685);
nand U14565 (N_14565,N_13037,N_13677);
and U14566 (N_14566,N_13006,N_13261);
and U14567 (N_14567,N_13895,N_13337);
nand U14568 (N_14568,N_13749,N_13049);
nor U14569 (N_14569,N_13303,N_13592);
nor U14570 (N_14570,N_13349,N_13330);
or U14571 (N_14571,N_13814,N_13433);
nor U14572 (N_14572,N_13968,N_13698);
xnor U14573 (N_14573,N_13807,N_13405);
and U14574 (N_14574,N_13373,N_13338);
nor U14575 (N_14575,N_13818,N_13683);
nand U14576 (N_14576,N_13298,N_13263);
xor U14577 (N_14577,N_13737,N_13259);
or U14578 (N_14578,N_13642,N_13363);
and U14579 (N_14579,N_13481,N_13570);
and U14580 (N_14580,N_13416,N_13062);
xor U14581 (N_14581,N_13880,N_13129);
nor U14582 (N_14582,N_13940,N_13552);
or U14583 (N_14583,N_13305,N_13624);
and U14584 (N_14584,N_13662,N_13654);
or U14585 (N_14585,N_13614,N_13324);
or U14586 (N_14586,N_13741,N_13222);
or U14587 (N_14587,N_13827,N_13502);
or U14588 (N_14588,N_13132,N_13504);
or U14589 (N_14589,N_13892,N_13202);
and U14590 (N_14590,N_13440,N_13206);
and U14591 (N_14591,N_13874,N_13788);
nor U14592 (N_14592,N_13279,N_13893);
nand U14593 (N_14593,N_13827,N_13275);
or U14594 (N_14594,N_13928,N_13983);
or U14595 (N_14595,N_13061,N_13885);
nand U14596 (N_14596,N_13540,N_13991);
nor U14597 (N_14597,N_13028,N_13490);
and U14598 (N_14598,N_13478,N_13259);
and U14599 (N_14599,N_13623,N_13388);
nor U14600 (N_14600,N_13732,N_13629);
and U14601 (N_14601,N_13927,N_13098);
nand U14602 (N_14602,N_13162,N_13547);
and U14603 (N_14603,N_13729,N_13688);
and U14604 (N_14604,N_13811,N_13403);
and U14605 (N_14605,N_13812,N_13538);
and U14606 (N_14606,N_13013,N_13371);
nor U14607 (N_14607,N_13827,N_13073);
xnor U14608 (N_14608,N_13807,N_13363);
nand U14609 (N_14609,N_13090,N_13273);
nor U14610 (N_14610,N_13388,N_13133);
nand U14611 (N_14611,N_13352,N_13320);
or U14612 (N_14612,N_13297,N_13418);
and U14613 (N_14613,N_13919,N_13953);
and U14614 (N_14614,N_13924,N_13212);
and U14615 (N_14615,N_13435,N_13806);
and U14616 (N_14616,N_13089,N_13724);
nand U14617 (N_14617,N_13859,N_13237);
nor U14618 (N_14618,N_13669,N_13301);
nand U14619 (N_14619,N_13483,N_13982);
xnor U14620 (N_14620,N_13807,N_13732);
and U14621 (N_14621,N_13450,N_13183);
nand U14622 (N_14622,N_13900,N_13698);
and U14623 (N_14623,N_13184,N_13277);
and U14624 (N_14624,N_13895,N_13753);
or U14625 (N_14625,N_13923,N_13449);
nor U14626 (N_14626,N_13057,N_13654);
or U14627 (N_14627,N_13684,N_13337);
nand U14628 (N_14628,N_13149,N_13051);
or U14629 (N_14629,N_13755,N_13799);
nand U14630 (N_14630,N_13406,N_13123);
or U14631 (N_14631,N_13907,N_13486);
nand U14632 (N_14632,N_13525,N_13796);
nand U14633 (N_14633,N_13101,N_13739);
nand U14634 (N_14634,N_13338,N_13190);
nor U14635 (N_14635,N_13435,N_13614);
or U14636 (N_14636,N_13354,N_13184);
or U14637 (N_14637,N_13562,N_13812);
nor U14638 (N_14638,N_13931,N_13440);
and U14639 (N_14639,N_13195,N_13638);
and U14640 (N_14640,N_13809,N_13912);
nand U14641 (N_14641,N_13745,N_13619);
nor U14642 (N_14642,N_13892,N_13217);
nand U14643 (N_14643,N_13252,N_13717);
nand U14644 (N_14644,N_13718,N_13497);
nor U14645 (N_14645,N_13271,N_13811);
and U14646 (N_14646,N_13395,N_13819);
nand U14647 (N_14647,N_13027,N_13300);
nand U14648 (N_14648,N_13739,N_13982);
nand U14649 (N_14649,N_13182,N_13572);
nor U14650 (N_14650,N_13320,N_13802);
nor U14651 (N_14651,N_13247,N_13916);
and U14652 (N_14652,N_13798,N_13851);
xnor U14653 (N_14653,N_13239,N_13094);
and U14654 (N_14654,N_13719,N_13677);
nor U14655 (N_14655,N_13351,N_13824);
or U14656 (N_14656,N_13060,N_13803);
nand U14657 (N_14657,N_13989,N_13367);
or U14658 (N_14658,N_13966,N_13717);
or U14659 (N_14659,N_13309,N_13932);
nand U14660 (N_14660,N_13468,N_13142);
nor U14661 (N_14661,N_13666,N_13655);
xnor U14662 (N_14662,N_13355,N_13269);
or U14663 (N_14663,N_13064,N_13808);
nand U14664 (N_14664,N_13807,N_13960);
or U14665 (N_14665,N_13254,N_13766);
and U14666 (N_14666,N_13840,N_13399);
and U14667 (N_14667,N_13528,N_13771);
nor U14668 (N_14668,N_13809,N_13244);
nand U14669 (N_14669,N_13553,N_13497);
and U14670 (N_14670,N_13472,N_13242);
nand U14671 (N_14671,N_13648,N_13645);
or U14672 (N_14672,N_13177,N_13417);
xor U14673 (N_14673,N_13624,N_13602);
nand U14674 (N_14674,N_13402,N_13631);
nand U14675 (N_14675,N_13254,N_13128);
nand U14676 (N_14676,N_13556,N_13069);
nand U14677 (N_14677,N_13157,N_13187);
xor U14678 (N_14678,N_13367,N_13761);
nor U14679 (N_14679,N_13547,N_13643);
nand U14680 (N_14680,N_13760,N_13036);
and U14681 (N_14681,N_13734,N_13246);
or U14682 (N_14682,N_13684,N_13863);
xnor U14683 (N_14683,N_13671,N_13168);
nand U14684 (N_14684,N_13084,N_13096);
nor U14685 (N_14685,N_13259,N_13847);
or U14686 (N_14686,N_13907,N_13853);
nand U14687 (N_14687,N_13525,N_13499);
nor U14688 (N_14688,N_13527,N_13896);
and U14689 (N_14689,N_13866,N_13708);
nand U14690 (N_14690,N_13776,N_13608);
nor U14691 (N_14691,N_13395,N_13582);
nor U14692 (N_14692,N_13491,N_13897);
or U14693 (N_14693,N_13950,N_13547);
or U14694 (N_14694,N_13833,N_13945);
nor U14695 (N_14695,N_13350,N_13795);
and U14696 (N_14696,N_13378,N_13851);
nor U14697 (N_14697,N_13698,N_13532);
nand U14698 (N_14698,N_13054,N_13183);
nand U14699 (N_14699,N_13887,N_13122);
or U14700 (N_14700,N_13671,N_13487);
or U14701 (N_14701,N_13727,N_13667);
or U14702 (N_14702,N_13201,N_13865);
or U14703 (N_14703,N_13506,N_13926);
and U14704 (N_14704,N_13021,N_13151);
and U14705 (N_14705,N_13962,N_13929);
nand U14706 (N_14706,N_13629,N_13206);
nor U14707 (N_14707,N_13536,N_13427);
and U14708 (N_14708,N_13764,N_13363);
nor U14709 (N_14709,N_13480,N_13457);
or U14710 (N_14710,N_13696,N_13361);
and U14711 (N_14711,N_13749,N_13982);
or U14712 (N_14712,N_13533,N_13686);
nor U14713 (N_14713,N_13548,N_13493);
and U14714 (N_14714,N_13708,N_13864);
nand U14715 (N_14715,N_13533,N_13461);
and U14716 (N_14716,N_13235,N_13988);
nand U14717 (N_14717,N_13516,N_13865);
or U14718 (N_14718,N_13485,N_13775);
xor U14719 (N_14719,N_13973,N_13182);
nor U14720 (N_14720,N_13755,N_13426);
nand U14721 (N_14721,N_13100,N_13329);
xor U14722 (N_14722,N_13923,N_13520);
xor U14723 (N_14723,N_13602,N_13557);
nand U14724 (N_14724,N_13183,N_13319);
nand U14725 (N_14725,N_13621,N_13406);
nor U14726 (N_14726,N_13776,N_13313);
or U14727 (N_14727,N_13779,N_13387);
and U14728 (N_14728,N_13120,N_13776);
or U14729 (N_14729,N_13064,N_13364);
or U14730 (N_14730,N_13587,N_13412);
nor U14731 (N_14731,N_13497,N_13402);
or U14732 (N_14732,N_13436,N_13637);
nor U14733 (N_14733,N_13632,N_13689);
xor U14734 (N_14734,N_13086,N_13376);
nand U14735 (N_14735,N_13070,N_13006);
nor U14736 (N_14736,N_13206,N_13247);
or U14737 (N_14737,N_13387,N_13839);
and U14738 (N_14738,N_13275,N_13693);
xnor U14739 (N_14739,N_13638,N_13025);
and U14740 (N_14740,N_13006,N_13930);
and U14741 (N_14741,N_13143,N_13991);
or U14742 (N_14742,N_13174,N_13655);
nand U14743 (N_14743,N_13986,N_13499);
nand U14744 (N_14744,N_13155,N_13036);
nor U14745 (N_14745,N_13985,N_13771);
nor U14746 (N_14746,N_13096,N_13115);
or U14747 (N_14747,N_13165,N_13375);
or U14748 (N_14748,N_13517,N_13022);
and U14749 (N_14749,N_13654,N_13449);
and U14750 (N_14750,N_13646,N_13916);
nor U14751 (N_14751,N_13852,N_13183);
and U14752 (N_14752,N_13840,N_13930);
and U14753 (N_14753,N_13326,N_13784);
xor U14754 (N_14754,N_13691,N_13201);
or U14755 (N_14755,N_13736,N_13239);
nor U14756 (N_14756,N_13806,N_13782);
nor U14757 (N_14757,N_13427,N_13090);
nor U14758 (N_14758,N_13772,N_13195);
nand U14759 (N_14759,N_13099,N_13024);
and U14760 (N_14760,N_13335,N_13495);
nor U14761 (N_14761,N_13645,N_13159);
or U14762 (N_14762,N_13634,N_13642);
or U14763 (N_14763,N_13403,N_13952);
and U14764 (N_14764,N_13153,N_13133);
or U14765 (N_14765,N_13382,N_13734);
and U14766 (N_14766,N_13527,N_13847);
nor U14767 (N_14767,N_13596,N_13135);
nor U14768 (N_14768,N_13749,N_13657);
or U14769 (N_14769,N_13689,N_13713);
nor U14770 (N_14770,N_13564,N_13729);
nand U14771 (N_14771,N_13328,N_13894);
nor U14772 (N_14772,N_13614,N_13905);
or U14773 (N_14773,N_13684,N_13560);
and U14774 (N_14774,N_13750,N_13255);
nand U14775 (N_14775,N_13923,N_13946);
nor U14776 (N_14776,N_13010,N_13557);
nor U14777 (N_14777,N_13519,N_13937);
nand U14778 (N_14778,N_13908,N_13115);
nand U14779 (N_14779,N_13096,N_13438);
nand U14780 (N_14780,N_13629,N_13170);
and U14781 (N_14781,N_13502,N_13012);
or U14782 (N_14782,N_13896,N_13700);
and U14783 (N_14783,N_13267,N_13176);
and U14784 (N_14784,N_13447,N_13496);
nor U14785 (N_14785,N_13155,N_13945);
and U14786 (N_14786,N_13320,N_13873);
nor U14787 (N_14787,N_13163,N_13053);
nor U14788 (N_14788,N_13656,N_13702);
nor U14789 (N_14789,N_13493,N_13420);
nor U14790 (N_14790,N_13835,N_13688);
nand U14791 (N_14791,N_13614,N_13813);
nor U14792 (N_14792,N_13676,N_13250);
nand U14793 (N_14793,N_13694,N_13401);
nor U14794 (N_14794,N_13934,N_13361);
nand U14795 (N_14795,N_13590,N_13486);
nor U14796 (N_14796,N_13331,N_13875);
nor U14797 (N_14797,N_13779,N_13691);
xnor U14798 (N_14798,N_13313,N_13038);
and U14799 (N_14799,N_13849,N_13035);
nand U14800 (N_14800,N_13120,N_13187);
nor U14801 (N_14801,N_13057,N_13019);
nor U14802 (N_14802,N_13280,N_13171);
nand U14803 (N_14803,N_13409,N_13452);
or U14804 (N_14804,N_13951,N_13032);
and U14805 (N_14805,N_13747,N_13833);
nor U14806 (N_14806,N_13413,N_13840);
or U14807 (N_14807,N_13131,N_13104);
and U14808 (N_14808,N_13903,N_13546);
nor U14809 (N_14809,N_13250,N_13539);
or U14810 (N_14810,N_13355,N_13343);
xor U14811 (N_14811,N_13242,N_13250);
nand U14812 (N_14812,N_13809,N_13037);
nor U14813 (N_14813,N_13654,N_13530);
or U14814 (N_14814,N_13486,N_13257);
nor U14815 (N_14815,N_13972,N_13756);
nand U14816 (N_14816,N_13825,N_13954);
nor U14817 (N_14817,N_13087,N_13291);
and U14818 (N_14818,N_13989,N_13008);
or U14819 (N_14819,N_13247,N_13554);
or U14820 (N_14820,N_13609,N_13690);
nor U14821 (N_14821,N_13429,N_13016);
and U14822 (N_14822,N_13870,N_13871);
nand U14823 (N_14823,N_13539,N_13948);
and U14824 (N_14824,N_13522,N_13996);
nor U14825 (N_14825,N_13017,N_13563);
nor U14826 (N_14826,N_13845,N_13860);
and U14827 (N_14827,N_13017,N_13577);
or U14828 (N_14828,N_13483,N_13523);
and U14829 (N_14829,N_13622,N_13985);
and U14830 (N_14830,N_13737,N_13745);
and U14831 (N_14831,N_13203,N_13162);
nand U14832 (N_14832,N_13814,N_13660);
nor U14833 (N_14833,N_13648,N_13049);
or U14834 (N_14834,N_13301,N_13558);
nor U14835 (N_14835,N_13185,N_13750);
xor U14836 (N_14836,N_13796,N_13800);
nor U14837 (N_14837,N_13239,N_13559);
or U14838 (N_14838,N_13377,N_13770);
and U14839 (N_14839,N_13205,N_13347);
nor U14840 (N_14840,N_13282,N_13657);
xnor U14841 (N_14841,N_13629,N_13676);
nor U14842 (N_14842,N_13436,N_13178);
xor U14843 (N_14843,N_13219,N_13895);
nor U14844 (N_14844,N_13805,N_13742);
and U14845 (N_14845,N_13965,N_13855);
or U14846 (N_14846,N_13841,N_13213);
and U14847 (N_14847,N_13791,N_13072);
nand U14848 (N_14848,N_13020,N_13016);
nor U14849 (N_14849,N_13501,N_13265);
xor U14850 (N_14850,N_13188,N_13265);
and U14851 (N_14851,N_13229,N_13453);
nand U14852 (N_14852,N_13914,N_13434);
xor U14853 (N_14853,N_13141,N_13527);
nor U14854 (N_14854,N_13214,N_13408);
nor U14855 (N_14855,N_13979,N_13090);
and U14856 (N_14856,N_13747,N_13712);
nor U14857 (N_14857,N_13195,N_13321);
nand U14858 (N_14858,N_13587,N_13318);
nor U14859 (N_14859,N_13080,N_13377);
nor U14860 (N_14860,N_13254,N_13461);
nand U14861 (N_14861,N_13238,N_13477);
nor U14862 (N_14862,N_13338,N_13861);
nand U14863 (N_14863,N_13626,N_13133);
and U14864 (N_14864,N_13052,N_13896);
and U14865 (N_14865,N_13480,N_13516);
nor U14866 (N_14866,N_13198,N_13220);
nor U14867 (N_14867,N_13857,N_13453);
nor U14868 (N_14868,N_13408,N_13052);
xor U14869 (N_14869,N_13728,N_13649);
nand U14870 (N_14870,N_13523,N_13184);
or U14871 (N_14871,N_13966,N_13344);
or U14872 (N_14872,N_13979,N_13980);
and U14873 (N_14873,N_13177,N_13193);
nand U14874 (N_14874,N_13096,N_13599);
and U14875 (N_14875,N_13639,N_13965);
nor U14876 (N_14876,N_13062,N_13137);
and U14877 (N_14877,N_13790,N_13317);
nand U14878 (N_14878,N_13297,N_13151);
nor U14879 (N_14879,N_13238,N_13922);
xor U14880 (N_14880,N_13695,N_13851);
nor U14881 (N_14881,N_13222,N_13402);
or U14882 (N_14882,N_13559,N_13002);
nand U14883 (N_14883,N_13161,N_13467);
nor U14884 (N_14884,N_13309,N_13197);
nand U14885 (N_14885,N_13129,N_13194);
nand U14886 (N_14886,N_13293,N_13622);
nor U14887 (N_14887,N_13260,N_13129);
nor U14888 (N_14888,N_13513,N_13664);
nor U14889 (N_14889,N_13500,N_13371);
or U14890 (N_14890,N_13659,N_13523);
or U14891 (N_14891,N_13589,N_13215);
nor U14892 (N_14892,N_13468,N_13209);
xor U14893 (N_14893,N_13160,N_13068);
nor U14894 (N_14894,N_13470,N_13671);
nand U14895 (N_14895,N_13495,N_13524);
and U14896 (N_14896,N_13627,N_13704);
and U14897 (N_14897,N_13288,N_13654);
nand U14898 (N_14898,N_13123,N_13687);
or U14899 (N_14899,N_13026,N_13978);
nand U14900 (N_14900,N_13129,N_13384);
or U14901 (N_14901,N_13313,N_13957);
nand U14902 (N_14902,N_13252,N_13297);
xnor U14903 (N_14903,N_13293,N_13802);
nand U14904 (N_14904,N_13081,N_13087);
or U14905 (N_14905,N_13948,N_13203);
nor U14906 (N_14906,N_13818,N_13061);
xnor U14907 (N_14907,N_13506,N_13240);
and U14908 (N_14908,N_13943,N_13287);
nor U14909 (N_14909,N_13838,N_13729);
nor U14910 (N_14910,N_13243,N_13584);
nor U14911 (N_14911,N_13273,N_13142);
nor U14912 (N_14912,N_13692,N_13453);
and U14913 (N_14913,N_13766,N_13776);
or U14914 (N_14914,N_13167,N_13845);
nand U14915 (N_14915,N_13087,N_13403);
or U14916 (N_14916,N_13055,N_13062);
nor U14917 (N_14917,N_13500,N_13289);
or U14918 (N_14918,N_13022,N_13688);
nand U14919 (N_14919,N_13228,N_13672);
xnor U14920 (N_14920,N_13529,N_13836);
or U14921 (N_14921,N_13300,N_13430);
nand U14922 (N_14922,N_13056,N_13250);
nor U14923 (N_14923,N_13240,N_13964);
and U14924 (N_14924,N_13877,N_13856);
nand U14925 (N_14925,N_13046,N_13030);
and U14926 (N_14926,N_13214,N_13632);
nand U14927 (N_14927,N_13597,N_13474);
nor U14928 (N_14928,N_13122,N_13587);
nor U14929 (N_14929,N_13219,N_13622);
nor U14930 (N_14930,N_13107,N_13759);
and U14931 (N_14931,N_13859,N_13962);
or U14932 (N_14932,N_13522,N_13304);
or U14933 (N_14933,N_13477,N_13235);
and U14934 (N_14934,N_13900,N_13982);
or U14935 (N_14935,N_13908,N_13117);
and U14936 (N_14936,N_13678,N_13036);
and U14937 (N_14937,N_13773,N_13304);
and U14938 (N_14938,N_13441,N_13256);
nand U14939 (N_14939,N_13217,N_13882);
or U14940 (N_14940,N_13258,N_13571);
nand U14941 (N_14941,N_13690,N_13041);
xor U14942 (N_14942,N_13555,N_13981);
and U14943 (N_14943,N_13976,N_13574);
or U14944 (N_14944,N_13219,N_13368);
xnor U14945 (N_14945,N_13166,N_13883);
nor U14946 (N_14946,N_13159,N_13670);
nand U14947 (N_14947,N_13812,N_13141);
nand U14948 (N_14948,N_13303,N_13158);
nand U14949 (N_14949,N_13396,N_13461);
and U14950 (N_14950,N_13034,N_13728);
or U14951 (N_14951,N_13790,N_13156);
and U14952 (N_14952,N_13197,N_13649);
or U14953 (N_14953,N_13808,N_13957);
nor U14954 (N_14954,N_13360,N_13568);
nor U14955 (N_14955,N_13229,N_13806);
nor U14956 (N_14956,N_13578,N_13477);
nor U14957 (N_14957,N_13934,N_13338);
nor U14958 (N_14958,N_13507,N_13258);
nor U14959 (N_14959,N_13563,N_13804);
and U14960 (N_14960,N_13353,N_13103);
xor U14961 (N_14961,N_13266,N_13687);
or U14962 (N_14962,N_13184,N_13716);
nand U14963 (N_14963,N_13877,N_13610);
nor U14964 (N_14964,N_13678,N_13467);
or U14965 (N_14965,N_13327,N_13511);
or U14966 (N_14966,N_13757,N_13698);
nor U14967 (N_14967,N_13547,N_13757);
nor U14968 (N_14968,N_13855,N_13666);
nor U14969 (N_14969,N_13796,N_13264);
and U14970 (N_14970,N_13021,N_13545);
and U14971 (N_14971,N_13453,N_13845);
nor U14972 (N_14972,N_13394,N_13976);
nor U14973 (N_14973,N_13974,N_13274);
and U14974 (N_14974,N_13824,N_13831);
xor U14975 (N_14975,N_13242,N_13982);
nor U14976 (N_14976,N_13036,N_13270);
nand U14977 (N_14977,N_13536,N_13552);
nor U14978 (N_14978,N_13623,N_13129);
nand U14979 (N_14979,N_13893,N_13435);
or U14980 (N_14980,N_13835,N_13108);
xnor U14981 (N_14981,N_13935,N_13618);
and U14982 (N_14982,N_13878,N_13581);
nand U14983 (N_14983,N_13690,N_13499);
nand U14984 (N_14984,N_13250,N_13483);
xnor U14985 (N_14985,N_13768,N_13157);
nand U14986 (N_14986,N_13863,N_13196);
and U14987 (N_14987,N_13191,N_13128);
nor U14988 (N_14988,N_13611,N_13293);
nor U14989 (N_14989,N_13357,N_13400);
nand U14990 (N_14990,N_13885,N_13781);
and U14991 (N_14991,N_13741,N_13505);
xor U14992 (N_14992,N_13975,N_13581);
and U14993 (N_14993,N_13602,N_13913);
nand U14994 (N_14994,N_13709,N_13605);
or U14995 (N_14995,N_13862,N_13859);
nor U14996 (N_14996,N_13095,N_13871);
and U14997 (N_14997,N_13198,N_13037);
nor U14998 (N_14998,N_13953,N_13599);
or U14999 (N_14999,N_13507,N_13745);
nand UO_0 (O_0,N_14341,N_14254);
xor UO_1 (O_1,N_14389,N_14233);
nor UO_2 (O_2,N_14805,N_14049);
nand UO_3 (O_3,N_14068,N_14033);
nor UO_4 (O_4,N_14931,N_14729);
nand UO_5 (O_5,N_14234,N_14079);
or UO_6 (O_6,N_14764,N_14130);
or UO_7 (O_7,N_14983,N_14451);
or UO_8 (O_8,N_14149,N_14510);
or UO_9 (O_9,N_14560,N_14175);
nor UO_10 (O_10,N_14865,N_14089);
nand UO_11 (O_11,N_14830,N_14531);
nor UO_12 (O_12,N_14737,N_14487);
and UO_13 (O_13,N_14042,N_14210);
and UO_14 (O_14,N_14190,N_14620);
and UO_15 (O_15,N_14375,N_14230);
or UO_16 (O_16,N_14193,N_14488);
or UO_17 (O_17,N_14436,N_14144);
and UO_18 (O_18,N_14929,N_14432);
or UO_19 (O_19,N_14602,N_14008);
or UO_20 (O_20,N_14109,N_14904);
or UO_21 (O_21,N_14847,N_14031);
nand UO_22 (O_22,N_14697,N_14960);
nor UO_23 (O_23,N_14530,N_14124);
or UO_24 (O_24,N_14051,N_14666);
and UO_25 (O_25,N_14761,N_14744);
or UO_26 (O_26,N_14368,N_14677);
and UO_27 (O_27,N_14526,N_14102);
and UO_28 (O_28,N_14594,N_14395);
nand UO_29 (O_29,N_14854,N_14947);
nand UO_30 (O_30,N_14552,N_14428);
or UO_31 (O_31,N_14152,N_14514);
or UO_32 (O_32,N_14192,N_14353);
nor UO_33 (O_33,N_14544,N_14586);
nand UO_34 (O_34,N_14335,N_14166);
nor UO_35 (O_35,N_14386,N_14182);
and UO_36 (O_36,N_14610,N_14917);
or UO_37 (O_37,N_14021,N_14674);
nand UO_38 (O_38,N_14468,N_14229);
nor UO_39 (O_39,N_14748,N_14427);
xnor UO_40 (O_40,N_14665,N_14735);
nand UO_41 (O_41,N_14794,N_14287);
and UO_42 (O_42,N_14683,N_14529);
or UO_43 (O_43,N_14592,N_14481);
nand UO_44 (O_44,N_14754,N_14534);
nand UO_45 (O_45,N_14621,N_14453);
and UO_46 (O_46,N_14284,N_14298);
nand UO_47 (O_47,N_14088,N_14222);
nand UO_48 (O_48,N_14450,N_14694);
or UO_49 (O_49,N_14227,N_14826);
and UO_50 (O_50,N_14212,N_14155);
xnor UO_51 (O_51,N_14199,N_14743);
or UO_52 (O_52,N_14306,N_14009);
and UO_53 (O_53,N_14523,N_14404);
nand UO_54 (O_54,N_14954,N_14897);
and UO_55 (O_55,N_14377,N_14799);
nor UO_56 (O_56,N_14739,N_14116);
and UO_57 (O_57,N_14161,N_14725);
nand UO_58 (O_58,N_14583,N_14036);
xnor UO_59 (O_59,N_14658,N_14422);
nor UO_60 (O_60,N_14562,N_14397);
or UO_61 (O_61,N_14168,N_14862);
nor UO_62 (O_62,N_14218,N_14567);
nor UO_63 (O_63,N_14028,N_14221);
nor UO_64 (O_64,N_14507,N_14880);
nor UO_65 (O_65,N_14364,N_14480);
nor UO_66 (O_66,N_14123,N_14500);
nor UO_67 (O_67,N_14457,N_14357);
or UO_68 (O_68,N_14924,N_14374);
and UO_69 (O_69,N_14540,N_14173);
nand UO_70 (O_70,N_14614,N_14656);
or UO_71 (O_71,N_14188,N_14812);
xor UO_72 (O_72,N_14977,N_14626);
and UO_73 (O_73,N_14103,N_14231);
and UO_74 (O_74,N_14454,N_14623);
nand UO_75 (O_75,N_14069,N_14025);
nor UO_76 (O_76,N_14919,N_14803);
or UO_77 (O_77,N_14804,N_14435);
nand UO_78 (O_78,N_14420,N_14169);
and UO_79 (O_79,N_14934,N_14871);
xnor UO_80 (O_80,N_14249,N_14712);
xor UO_81 (O_81,N_14956,N_14825);
and UO_82 (O_82,N_14732,N_14047);
and UO_83 (O_83,N_14925,N_14545);
nor UO_84 (O_84,N_14408,N_14177);
nor UO_85 (O_85,N_14228,N_14020);
or UO_86 (O_86,N_14660,N_14708);
or UO_87 (O_87,N_14581,N_14914);
and UO_88 (O_88,N_14533,N_14074);
nor UO_89 (O_89,N_14553,N_14277);
nand UO_90 (O_90,N_14394,N_14446);
nor UO_91 (O_91,N_14183,N_14414);
nand UO_92 (O_92,N_14752,N_14490);
xor UO_93 (O_93,N_14981,N_14775);
or UO_94 (O_94,N_14477,N_14860);
and UO_95 (O_95,N_14097,N_14844);
xor UO_96 (O_96,N_14524,N_14519);
or UO_97 (O_97,N_14585,N_14271);
xor UO_98 (O_98,N_14355,N_14894);
nor UO_99 (O_99,N_14757,N_14441);
or UO_100 (O_100,N_14122,N_14841);
and UO_101 (O_101,N_14755,N_14989);
or UO_102 (O_102,N_14527,N_14098);
and UO_103 (O_103,N_14384,N_14834);
nand UO_104 (O_104,N_14232,N_14083);
and UO_105 (O_105,N_14588,N_14037);
or UO_106 (O_106,N_14817,N_14299);
and UO_107 (O_107,N_14644,N_14948);
or UO_108 (O_108,N_14348,N_14134);
or UO_109 (O_109,N_14317,N_14164);
and UO_110 (O_110,N_14387,N_14113);
nor UO_111 (O_111,N_14696,N_14986);
or UO_112 (O_112,N_14250,N_14849);
and UO_113 (O_113,N_14314,N_14738);
and UO_114 (O_114,N_14807,N_14253);
nor UO_115 (O_115,N_14520,N_14516);
or UO_116 (O_116,N_14591,N_14793);
or UO_117 (O_117,N_14749,N_14861);
nand UO_118 (O_118,N_14885,N_14874);
or UO_119 (O_119,N_14845,N_14979);
or UO_120 (O_120,N_14970,N_14247);
nand UO_121 (O_121,N_14165,N_14542);
and UO_122 (O_122,N_14310,N_14781);
and UO_123 (O_123,N_14902,N_14730);
and UO_124 (O_124,N_14506,N_14601);
or UO_125 (O_125,N_14637,N_14288);
and UO_126 (O_126,N_14908,N_14699);
nor UO_127 (O_127,N_14439,N_14121);
and UO_128 (O_128,N_14101,N_14686);
and UO_129 (O_129,N_14114,N_14731);
or UO_130 (O_130,N_14964,N_14443);
or UO_131 (O_131,N_14640,N_14330);
nand UO_132 (O_132,N_14401,N_14460);
xnor UO_133 (O_133,N_14779,N_14044);
and UO_134 (O_134,N_14638,N_14476);
or UO_135 (O_135,N_14590,N_14266);
nand UO_136 (O_136,N_14281,N_14302);
and UO_137 (O_137,N_14344,N_14503);
nand UO_138 (O_138,N_14001,N_14667);
nand UO_139 (O_139,N_14184,N_14492);
nor UO_140 (O_140,N_14099,N_14556);
nor UO_141 (O_141,N_14126,N_14251);
nor UO_142 (O_142,N_14559,N_14868);
nand UO_143 (O_143,N_14691,N_14709);
nor UO_144 (O_144,N_14572,N_14974);
nor UO_145 (O_145,N_14521,N_14379);
nor UO_146 (O_146,N_14551,N_14073);
nor UO_147 (O_147,N_14027,N_14693);
xor UO_148 (O_148,N_14574,N_14063);
nand UO_149 (O_149,N_14575,N_14426);
and UO_150 (O_150,N_14056,N_14349);
or UO_151 (O_151,N_14362,N_14313);
or UO_152 (O_152,N_14207,N_14046);
or UO_153 (O_153,N_14167,N_14373);
and UO_154 (O_154,N_14901,N_14273);
nor UO_155 (O_155,N_14787,N_14999);
or UO_156 (O_156,N_14054,N_14041);
nor UO_157 (O_157,N_14957,N_14608);
nand UO_158 (O_158,N_14189,N_14053);
nor UO_159 (O_159,N_14923,N_14953);
xor UO_160 (O_160,N_14040,N_14652);
xnor UO_161 (O_161,N_14061,N_14815);
nor UO_162 (O_162,N_14208,N_14331);
nor UO_163 (O_163,N_14518,N_14140);
or UO_164 (O_164,N_14390,N_14528);
and UO_165 (O_165,N_14186,N_14104);
nand UO_166 (O_166,N_14625,N_14196);
nor UO_167 (O_167,N_14760,N_14203);
nand UO_168 (O_168,N_14918,N_14776);
and UO_169 (O_169,N_14415,N_14241);
or UO_170 (O_170,N_14216,N_14367);
and UO_171 (O_171,N_14292,N_14052);
or UO_172 (O_172,N_14745,N_14998);
or UO_173 (O_173,N_14090,N_14796);
and UO_174 (O_174,N_14472,N_14498);
nand UO_175 (O_175,N_14238,N_14549);
nand UO_176 (O_176,N_14502,N_14452);
and UO_177 (O_177,N_14671,N_14151);
or UO_178 (O_178,N_14906,N_14370);
and UO_179 (O_179,N_14990,N_14176);
or UO_180 (O_180,N_14806,N_14034);
xor UO_181 (O_181,N_14282,N_14758);
nor UO_182 (O_182,N_14159,N_14064);
or UO_183 (O_183,N_14657,N_14710);
or UO_184 (O_184,N_14846,N_14645);
or UO_185 (O_185,N_14138,N_14599);
nor UO_186 (O_186,N_14486,N_14474);
nand UO_187 (O_187,N_14078,N_14339);
or UO_188 (O_188,N_14703,N_14820);
and UO_189 (O_189,N_14267,N_14418);
nor UO_190 (O_190,N_14162,N_14920);
or UO_191 (O_191,N_14410,N_14359);
nand UO_192 (O_192,N_14909,N_14067);
and UO_193 (O_193,N_14568,N_14839);
nand UO_194 (O_194,N_14726,N_14289);
and UO_195 (O_195,N_14765,N_14791);
nor UO_196 (O_196,N_14855,N_14566);
and UO_197 (O_197,N_14810,N_14782);
nor UO_198 (O_198,N_14360,N_14680);
nor UO_199 (O_199,N_14080,N_14322);
nor UO_200 (O_200,N_14900,N_14022);
or UO_201 (O_201,N_14940,N_14442);
nor UO_202 (O_202,N_14848,N_14185);
or UO_203 (O_203,N_14718,N_14783);
or UO_204 (O_204,N_14023,N_14741);
or UO_205 (O_205,N_14961,N_14984);
and UO_206 (O_206,N_14993,N_14043);
or UO_207 (O_207,N_14985,N_14600);
nor UO_208 (O_208,N_14096,N_14818);
or UO_209 (O_209,N_14076,N_14148);
nor UO_210 (O_210,N_14938,N_14639);
xor UO_211 (O_211,N_14136,N_14676);
and UO_212 (O_212,N_14011,N_14946);
xor UO_213 (O_213,N_14072,N_14747);
xor UO_214 (O_214,N_14728,N_14262);
nand UO_215 (O_215,N_14935,N_14944);
or UO_216 (O_216,N_14107,N_14388);
nor UO_217 (O_217,N_14672,N_14777);
and UO_218 (O_218,N_14899,N_14139);
or UO_219 (O_219,N_14685,N_14337);
nor UO_220 (O_220,N_14170,N_14504);
nor UO_221 (O_221,N_14641,N_14204);
and UO_222 (O_222,N_14091,N_14878);
xor UO_223 (O_223,N_14881,N_14770);
nor UO_224 (O_224,N_14603,N_14509);
and UO_225 (O_225,N_14424,N_14734);
nand UO_226 (O_226,N_14324,N_14886);
nand UO_227 (O_227,N_14835,N_14485);
nor UO_228 (O_228,N_14336,N_14987);
xnor UO_229 (O_229,N_14030,N_14154);
and UO_230 (O_230,N_14279,N_14045);
or UO_231 (O_231,N_14704,N_14700);
nor UO_232 (O_232,N_14129,N_14505);
and UO_233 (O_233,N_14746,N_14543);
xnor UO_234 (O_234,N_14320,N_14333);
and UO_235 (O_235,N_14921,N_14873);
and UO_236 (O_236,N_14851,N_14235);
nor UO_237 (O_237,N_14215,N_14882);
nand UO_238 (O_238,N_14692,N_14604);
or UO_239 (O_239,N_14634,N_14866);
and UO_240 (O_240,N_14967,N_14681);
nand UO_241 (O_241,N_14237,N_14365);
or UO_242 (O_242,N_14955,N_14135);
xor UO_243 (O_243,N_14483,N_14301);
or UO_244 (O_244,N_14513,N_14831);
or UO_245 (O_245,N_14890,N_14399);
xnor UO_246 (O_246,N_14363,N_14822);
nand UO_247 (O_247,N_14912,N_14576);
nor UO_248 (O_248,N_14720,N_14012);
xor UO_249 (O_249,N_14891,N_14265);
nand UO_250 (O_250,N_14112,N_14417);
nor UO_251 (O_251,N_14774,N_14589);
or UO_252 (O_252,N_14653,N_14536);
or UO_253 (O_253,N_14382,N_14870);
nand UO_254 (O_254,N_14716,N_14690);
nor UO_255 (O_255,N_14872,N_14558);
and UO_256 (O_256,N_14115,N_14577);
nand UO_257 (O_257,N_14085,N_14013);
and UO_258 (O_258,N_14778,N_14297);
or UO_259 (O_259,N_14461,N_14682);
xor UO_260 (O_260,N_14662,N_14290);
or UO_261 (O_261,N_14376,N_14580);
xor UO_262 (O_262,N_14338,N_14467);
or UO_263 (O_263,N_14879,N_14120);
nand UO_264 (O_264,N_14242,N_14635);
nand UO_265 (O_265,N_14828,N_14888);
nand UO_266 (O_266,N_14618,N_14717);
nor UO_267 (O_267,N_14911,N_14372);
xnor UO_268 (O_268,N_14315,N_14383);
nand UO_269 (O_269,N_14100,N_14156);
nand UO_270 (O_270,N_14187,N_14018);
or UO_271 (O_271,N_14833,N_14201);
nand UO_272 (O_272,N_14272,N_14239);
or UO_273 (O_273,N_14323,N_14615);
or UO_274 (O_274,N_14470,N_14016);
xnor UO_275 (O_275,N_14670,N_14128);
nor UO_276 (O_276,N_14412,N_14922);
xor UO_277 (O_277,N_14525,N_14191);
and UO_278 (O_278,N_14174,N_14260);
nor UO_279 (O_279,N_14800,N_14889);
xnor UO_280 (O_280,N_14555,N_14026);
xnor UO_281 (O_281,N_14892,N_14606);
or UO_282 (O_282,N_14393,N_14565);
nand UO_283 (O_283,N_14180,N_14941);
nand UO_284 (O_284,N_14569,N_14798);
nor UO_285 (O_285,N_14980,N_14263);
nand UO_286 (O_286,N_14226,N_14869);
nor UO_287 (O_287,N_14877,N_14198);
and UO_288 (O_288,N_14029,N_14449);
and UO_289 (O_289,N_14343,N_14719);
and UO_290 (O_290,N_14522,N_14243);
nand UO_291 (O_291,N_14887,N_14497);
or UO_292 (O_292,N_14548,N_14724);
and UO_293 (O_293,N_14236,N_14403);
or UO_294 (O_294,N_14907,N_14809);
and UO_295 (O_295,N_14132,N_14111);
nor UO_296 (O_296,N_14264,N_14982);
and UO_297 (O_297,N_14727,N_14780);
or UO_298 (O_298,N_14421,N_14311);
or UO_299 (O_299,N_14062,N_14274);
nand UO_300 (O_300,N_14673,N_14378);
nand UO_301 (O_301,N_14535,N_14932);
and UO_302 (O_302,N_14075,N_14973);
nor UO_303 (O_303,N_14352,N_14400);
nand UO_304 (O_304,N_14048,N_14547);
or UO_305 (O_305,N_14391,N_14679);
nand UO_306 (O_306,N_14145,N_14269);
nor UO_307 (O_307,N_14214,N_14814);
nand UO_308 (O_308,N_14707,N_14795);
and UO_309 (O_309,N_14392,N_14223);
or UO_310 (O_310,N_14605,N_14642);
and UO_311 (O_311,N_14711,N_14479);
nor UO_312 (O_312,N_14157,N_14444);
or UO_313 (O_313,N_14131,N_14596);
nand UO_314 (O_314,N_14629,N_14327);
nand UO_315 (O_315,N_14402,N_14915);
or UO_316 (O_316,N_14722,N_14296);
and UO_317 (O_317,N_14687,N_14092);
nor UO_318 (O_318,N_14786,N_14675);
nand UO_319 (O_319,N_14039,N_14936);
xor UO_320 (O_320,N_14276,N_14584);
and UO_321 (O_321,N_14661,N_14651);
nand UO_322 (O_322,N_14876,N_14325);
or UO_323 (O_323,N_14893,N_14838);
and UO_324 (O_324,N_14240,N_14705);
and UO_325 (O_325,N_14991,N_14319);
or UO_326 (O_326,N_14557,N_14756);
and UO_327 (O_327,N_14491,N_14930);
nor UO_328 (O_328,N_14406,N_14723);
nand UO_329 (O_329,N_14206,N_14702);
and UO_330 (O_330,N_14246,N_14416);
xor UO_331 (O_331,N_14050,N_14578);
or UO_332 (O_332,N_14994,N_14958);
nand UO_333 (O_333,N_14972,N_14750);
and UO_334 (O_334,N_14329,N_14407);
nor UO_335 (O_335,N_14385,N_14094);
or UO_336 (O_336,N_14773,N_14701);
or UO_337 (O_337,N_14005,N_14598);
or UO_338 (O_338,N_14494,N_14105);
and UO_339 (O_339,N_14294,N_14740);
or UO_340 (O_340,N_14867,N_14883);
and UO_341 (O_341,N_14976,N_14762);
and UO_342 (O_342,N_14733,N_14648);
nand UO_343 (O_343,N_14462,N_14573);
xor UO_344 (O_344,N_14633,N_14995);
or UO_345 (O_345,N_14181,N_14110);
nor UO_346 (O_346,N_14537,N_14484);
nand UO_347 (O_347,N_14448,N_14541);
nor UO_348 (O_348,N_14678,N_14624);
nand UO_349 (O_349,N_14579,N_14561);
nor UO_350 (O_350,N_14347,N_14926);
and UO_351 (O_351,N_14607,N_14646);
and UO_352 (O_352,N_14736,N_14808);
nand UO_353 (O_353,N_14664,N_14650);
nor UO_354 (O_354,N_14202,N_14000);
and UO_355 (O_355,N_14437,N_14975);
xor UO_356 (O_356,N_14963,N_14200);
nor UO_357 (O_357,N_14706,N_14086);
nor UO_358 (O_358,N_14714,N_14351);
nor UO_359 (O_359,N_14859,N_14065);
nand UO_360 (O_360,N_14419,N_14396);
nor UO_361 (O_361,N_14059,N_14007);
nand UO_362 (O_362,N_14832,N_14695);
nand UO_363 (O_363,N_14595,N_14689);
or UO_364 (O_364,N_14823,N_14827);
and UO_365 (O_365,N_14597,N_14413);
or UO_366 (O_366,N_14459,N_14160);
nor UO_367 (O_367,N_14628,N_14158);
or UO_368 (O_368,N_14721,N_14071);
nand UO_369 (O_369,N_14582,N_14627);
or UO_370 (O_370,N_14147,N_14270);
or UO_371 (O_371,N_14655,N_14713);
and UO_372 (O_372,N_14996,N_14913);
and UO_373 (O_373,N_14211,N_14636);
and UO_374 (O_374,N_14366,N_14261);
or UO_375 (O_375,N_14308,N_14496);
nand UO_376 (O_376,N_14884,N_14684);
and UO_377 (O_377,N_14127,N_14669);
nand UO_378 (O_378,N_14429,N_14334);
and UO_379 (O_379,N_14843,N_14482);
and UO_380 (O_380,N_14445,N_14440);
nor UO_381 (O_381,N_14268,N_14829);
nor UO_382 (O_382,N_14058,N_14649);
xor UO_383 (O_383,N_14035,N_14951);
nor UO_384 (O_384,N_14280,N_14788);
and UO_385 (O_385,N_14286,N_14587);
or UO_386 (O_386,N_14742,N_14434);
and UO_387 (O_387,N_14019,N_14864);
nand UO_388 (O_388,N_14093,N_14409);
nand UO_389 (O_389,N_14769,N_14593);
nor UO_390 (O_390,N_14398,N_14220);
or UO_391 (O_391,N_14501,N_14927);
and UO_392 (O_392,N_14789,N_14784);
nand UO_393 (O_393,N_14217,N_14117);
nor UO_394 (O_394,N_14178,N_14084);
or UO_395 (O_395,N_14458,N_14563);
or UO_396 (O_396,N_14082,N_14611);
xor UO_397 (O_397,N_14802,N_14455);
and UO_398 (O_398,N_14195,N_14354);
nand UO_399 (O_399,N_14617,N_14381);
or UO_400 (O_400,N_14425,N_14356);
xnor UO_401 (O_401,N_14546,N_14340);
xor UO_402 (O_402,N_14463,N_14225);
and UO_403 (O_403,N_14055,N_14856);
or UO_404 (O_404,N_14316,N_14332);
nand UO_405 (O_405,N_14002,N_14209);
nor UO_406 (O_406,N_14345,N_14473);
and UO_407 (O_407,N_14017,N_14006);
nand UO_408 (O_408,N_14863,N_14350);
or UO_409 (O_409,N_14309,N_14772);
and UO_410 (O_410,N_14060,N_14813);
nor UO_411 (O_411,N_14928,N_14303);
nor UO_412 (O_412,N_14875,N_14997);
and UO_413 (O_413,N_14465,N_14937);
nor UO_414 (O_414,N_14643,N_14371);
nand UO_415 (O_415,N_14137,N_14853);
nor UO_416 (O_416,N_14898,N_14971);
xor UO_417 (O_417,N_14307,N_14816);
xnor UO_418 (O_418,N_14038,N_14143);
and UO_419 (O_419,N_14179,N_14003);
or UO_420 (O_420,N_14125,N_14654);
nor UO_421 (O_421,N_14493,N_14171);
xnor UO_422 (O_422,N_14962,N_14087);
nand UO_423 (O_423,N_14939,N_14194);
or UO_424 (O_424,N_14213,N_14057);
and UO_425 (O_425,N_14118,N_14153);
and UO_426 (O_426,N_14751,N_14619);
or UO_427 (O_427,N_14508,N_14106);
and UO_428 (O_428,N_14571,N_14630);
xnor UO_429 (O_429,N_14609,N_14933);
and UO_430 (O_430,N_14968,N_14346);
or UO_431 (O_431,N_14688,N_14616);
and UO_432 (O_432,N_14108,N_14466);
nand UO_433 (O_433,N_14024,N_14857);
nor UO_434 (O_434,N_14768,N_14423);
nor UO_435 (O_435,N_14258,N_14300);
and UO_436 (O_436,N_14515,N_14430);
and UO_437 (O_437,N_14550,N_14992);
nor UO_438 (O_438,N_14622,N_14197);
xor UO_439 (O_439,N_14647,N_14405);
nor UO_440 (O_440,N_14369,N_14464);
or UO_441 (O_441,N_14245,N_14852);
nor UO_442 (O_442,N_14469,N_14959);
nand UO_443 (O_443,N_14753,N_14478);
nand UO_444 (O_444,N_14305,N_14517);
or UO_445 (O_445,N_14321,N_14819);
nand UO_446 (O_446,N_14766,N_14612);
or UO_447 (O_447,N_14163,N_14014);
nand UO_448 (O_448,N_14836,N_14942);
and UO_449 (O_449,N_14066,N_14797);
xor UO_450 (O_450,N_14431,N_14837);
and UO_451 (O_451,N_14133,N_14988);
nor UO_452 (O_452,N_14312,N_14293);
or UO_453 (O_453,N_14256,N_14965);
xor UO_454 (O_454,N_14141,N_14004);
or UO_455 (O_455,N_14248,N_14811);
nor UO_456 (O_456,N_14824,N_14790);
or UO_457 (O_457,N_14275,N_14257);
nor UO_458 (O_458,N_14255,N_14570);
nor UO_459 (O_459,N_14978,N_14081);
nand UO_460 (O_460,N_14146,N_14896);
and UO_461 (O_461,N_14304,N_14244);
nor UO_462 (O_462,N_14969,N_14792);
or UO_463 (O_463,N_14015,N_14291);
and UO_464 (O_464,N_14538,N_14966);
and UO_465 (O_465,N_14895,N_14905);
and UO_466 (O_466,N_14850,N_14219);
and UO_467 (O_467,N_14495,N_14438);
or UO_468 (O_468,N_14070,N_14489);
xor UO_469 (O_469,N_14142,N_14916);
and UO_470 (O_470,N_14278,N_14613);
xor UO_471 (O_471,N_14342,N_14318);
and UO_472 (O_472,N_14512,N_14943);
nor UO_473 (O_473,N_14858,N_14952);
and UO_474 (O_474,N_14759,N_14172);
and UO_475 (O_475,N_14539,N_14949);
nor UO_476 (O_476,N_14285,N_14767);
nand UO_477 (O_477,N_14554,N_14564);
xnor UO_478 (O_478,N_14259,N_14224);
and UO_479 (O_479,N_14821,N_14411);
and UO_480 (O_480,N_14499,N_14659);
and UO_481 (O_481,N_14842,N_14785);
and UO_482 (O_482,N_14840,N_14328);
nand UO_483 (O_483,N_14095,N_14771);
nand UO_484 (O_484,N_14380,N_14715);
nand UO_485 (O_485,N_14632,N_14150);
nor UO_486 (O_486,N_14205,N_14698);
nand UO_487 (O_487,N_14801,N_14252);
nor UO_488 (O_488,N_14631,N_14950);
nand UO_489 (O_489,N_14326,N_14077);
or UO_490 (O_490,N_14663,N_14119);
and UO_491 (O_491,N_14456,N_14295);
and UO_492 (O_492,N_14447,N_14668);
nand UO_493 (O_493,N_14433,N_14471);
nor UO_494 (O_494,N_14532,N_14283);
or UO_495 (O_495,N_14511,N_14945);
nor UO_496 (O_496,N_14475,N_14358);
or UO_497 (O_497,N_14763,N_14910);
or UO_498 (O_498,N_14032,N_14010);
or UO_499 (O_499,N_14361,N_14903);
nor UO_500 (O_500,N_14902,N_14325);
or UO_501 (O_501,N_14122,N_14977);
or UO_502 (O_502,N_14683,N_14024);
nor UO_503 (O_503,N_14079,N_14011);
nand UO_504 (O_504,N_14497,N_14412);
or UO_505 (O_505,N_14540,N_14387);
xnor UO_506 (O_506,N_14886,N_14074);
or UO_507 (O_507,N_14921,N_14107);
and UO_508 (O_508,N_14634,N_14284);
nor UO_509 (O_509,N_14236,N_14081);
or UO_510 (O_510,N_14966,N_14273);
and UO_511 (O_511,N_14789,N_14731);
and UO_512 (O_512,N_14160,N_14274);
and UO_513 (O_513,N_14488,N_14327);
xor UO_514 (O_514,N_14801,N_14896);
nor UO_515 (O_515,N_14623,N_14917);
nor UO_516 (O_516,N_14559,N_14855);
or UO_517 (O_517,N_14960,N_14909);
and UO_518 (O_518,N_14790,N_14213);
xnor UO_519 (O_519,N_14035,N_14994);
or UO_520 (O_520,N_14803,N_14133);
and UO_521 (O_521,N_14483,N_14861);
nor UO_522 (O_522,N_14650,N_14048);
and UO_523 (O_523,N_14843,N_14960);
nand UO_524 (O_524,N_14098,N_14265);
and UO_525 (O_525,N_14937,N_14666);
nor UO_526 (O_526,N_14455,N_14388);
or UO_527 (O_527,N_14274,N_14173);
and UO_528 (O_528,N_14178,N_14320);
or UO_529 (O_529,N_14609,N_14573);
or UO_530 (O_530,N_14412,N_14014);
nand UO_531 (O_531,N_14092,N_14134);
or UO_532 (O_532,N_14258,N_14866);
and UO_533 (O_533,N_14629,N_14465);
xnor UO_534 (O_534,N_14554,N_14415);
nor UO_535 (O_535,N_14751,N_14320);
nor UO_536 (O_536,N_14052,N_14520);
nand UO_537 (O_537,N_14879,N_14741);
xnor UO_538 (O_538,N_14077,N_14661);
nand UO_539 (O_539,N_14264,N_14301);
nor UO_540 (O_540,N_14408,N_14578);
or UO_541 (O_541,N_14141,N_14355);
nor UO_542 (O_542,N_14333,N_14908);
or UO_543 (O_543,N_14793,N_14616);
nor UO_544 (O_544,N_14417,N_14298);
and UO_545 (O_545,N_14778,N_14142);
nor UO_546 (O_546,N_14866,N_14203);
and UO_547 (O_547,N_14731,N_14526);
nand UO_548 (O_548,N_14974,N_14096);
nor UO_549 (O_549,N_14647,N_14883);
nor UO_550 (O_550,N_14099,N_14334);
xnor UO_551 (O_551,N_14641,N_14953);
and UO_552 (O_552,N_14333,N_14351);
nor UO_553 (O_553,N_14377,N_14644);
nor UO_554 (O_554,N_14088,N_14987);
nor UO_555 (O_555,N_14057,N_14340);
nand UO_556 (O_556,N_14120,N_14482);
or UO_557 (O_557,N_14980,N_14544);
or UO_558 (O_558,N_14708,N_14374);
nor UO_559 (O_559,N_14129,N_14539);
and UO_560 (O_560,N_14810,N_14311);
nand UO_561 (O_561,N_14609,N_14478);
xnor UO_562 (O_562,N_14335,N_14771);
nand UO_563 (O_563,N_14732,N_14197);
nand UO_564 (O_564,N_14951,N_14574);
or UO_565 (O_565,N_14352,N_14869);
or UO_566 (O_566,N_14620,N_14167);
nand UO_567 (O_567,N_14063,N_14415);
or UO_568 (O_568,N_14061,N_14510);
and UO_569 (O_569,N_14905,N_14002);
or UO_570 (O_570,N_14685,N_14785);
and UO_571 (O_571,N_14218,N_14796);
nor UO_572 (O_572,N_14226,N_14060);
nor UO_573 (O_573,N_14067,N_14263);
nor UO_574 (O_574,N_14757,N_14345);
nor UO_575 (O_575,N_14114,N_14929);
or UO_576 (O_576,N_14611,N_14857);
or UO_577 (O_577,N_14640,N_14639);
and UO_578 (O_578,N_14096,N_14584);
nor UO_579 (O_579,N_14141,N_14292);
and UO_580 (O_580,N_14910,N_14681);
or UO_581 (O_581,N_14083,N_14354);
and UO_582 (O_582,N_14336,N_14716);
nand UO_583 (O_583,N_14952,N_14839);
and UO_584 (O_584,N_14757,N_14973);
nor UO_585 (O_585,N_14565,N_14356);
xor UO_586 (O_586,N_14802,N_14280);
nand UO_587 (O_587,N_14385,N_14985);
xnor UO_588 (O_588,N_14593,N_14898);
nand UO_589 (O_589,N_14213,N_14443);
xor UO_590 (O_590,N_14922,N_14850);
nor UO_591 (O_591,N_14626,N_14301);
nor UO_592 (O_592,N_14920,N_14117);
nand UO_593 (O_593,N_14733,N_14553);
nand UO_594 (O_594,N_14195,N_14342);
or UO_595 (O_595,N_14378,N_14790);
nor UO_596 (O_596,N_14336,N_14963);
or UO_597 (O_597,N_14353,N_14670);
nand UO_598 (O_598,N_14848,N_14567);
and UO_599 (O_599,N_14372,N_14210);
nand UO_600 (O_600,N_14398,N_14858);
nor UO_601 (O_601,N_14964,N_14213);
and UO_602 (O_602,N_14306,N_14603);
nand UO_603 (O_603,N_14389,N_14250);
nor UO_604 (O_604,N_14195,N_14393);
xnor UO_605 (O_605,N_14281,N_14525);
and UO_606 (O_606,N_14282,N_14418);
nand UO_607 (O_607,N_14566,N_14251);
nand UO_608 (O_608,N_14264,N_14335);
nor UO_609 (O_609,N_14658,N_14184);
nor UO_610 (O_610,N_14093,N_14405);
and UO_611 (O_611,N_14802,N_14966);
or UO_612 (O_612,N_14200,N_14049);
or UO_613 (O_613,N_14239,N_14648);
xnor UO_614 (O_614,N_14166,N_14790);
nand UO_615 (O_615,N_14909,N_14776);
and UO_616 (O_616,N_14821,N_14880);
or UO_617 (O_617,N_14981,N_14259);
xnor UO_618 (O_618,N_14051,N_14818);
nor UO_619 (O_619,N_14306,N_14749);
nand UO_620 (O_620,N_14849,N_14230);
or UO_621 (O_621,N_14712,N_14597);
nor UO_622 (O_622,N_14013,N_14708);
nand UO_623 (O_623,N_14186,N_14313);
and UO_624 (O_624,N_14748,N_14960);
and UO_625 (O_625,N_14226,N_14327);
nor UO_626 (O_626,N_14738,N_14159);
nand UO_627 (O_627,N_14013,N_14875);
and UO_628 (O_628,N_14617,N_14294);
or UO_629 (O_629,N_14516,N_14030);
and UO_630 (O_630,N_14713,N_14683);
nand UO_631 (O_631,N_14384,N_14984);
xor UO_632 (O_632,N_14169,N_14019);
or UO_633 (O_633,N_14175,N_14643);
nand UO_634 (O_634,N_14183,N_14655);
nand UO_635 (O_635,N_14524,N_14319);
or UO_636 (O_636,N_14920,N_14062);
nor UO_637 (O_637,N_14163,N_14046);
nor UO_638 (O_638,N_14881,N_14365);
nor UO_639 (O_639,N_14859,N_14511);
nor UO_640 (O_640,N_14846,N_14506);
nand UO_641 (O_641,N_14114,N_14735);
nand UO_642 (O_642,N_14878,N_14995);
nor UO_643 (O_643,N_14231,N_14353);
xnor UO_644 (O_644,N_14738,N_14724);
nor UO_645 (O_645,N_14394,N_14005);
nand UO_646 (O_646,N_14229,N_14676);
nand UO_647 (O_647,N_14681,N_14141);
and UO_648 (O_648,N_14434,N_14075);
and UO_649 (O_649,N_14981,N_14929);
nand UO_650 (O_650,N_14556,N_14074);
nand UO_651 (O_651,N_14423,N_14245);
or UO_652 (O_652,N_14305,N_14368);
nand UO_653 (O_653,N_14245,N_14350);
xnor UO_654 (O_654,N_14132,N_14149);
or UO_655 (O_655,N_14004,N_14875);
and UO_656 (O_656,N_14534,N_14948);
and UO_657 (O_657,N_14640,N_14012);
or UO_658 (O_658,N_14153,N_14341);
nor UO_659 (O_659,N_14335,N_14821);
nor UO_660 (O_660,N_14010,N_14290);
and UO_661 (O_661,N_14266,N_14332);
nand UO_662 (O_662,N_14561,N_14709);
and UO_663 (O_663,N_14886,N_14674);
xnor UO_664 (O_664,N_14766,N_14671);
and UO_665 (O_665,N_14898,N_14618);
and UO_666 (O_666,N_14712,N_14856);
nand UO_667 (O_667,N_14233,N_14381);
and UO_668 (O_668,N_14841,N_14883);
nand UO_669 (O_669,N_14969,N_14993);
or UO_670 (O_670,N_14620,N_14729);
or UO_671 (O_671,N_14126,N_14046);
xnor UO_672 (O_672,N_14058,N_14245);
and UO_673 (O_673,N_14249,N_14220);
and UO_674 (O_674,N_14535,N_14569);
nand UO_675 (O_675,N_14821,N_14378);
nand UO_676 (O_676,N_14886,N_14063);
nand UO_677 (O_677,N_14166,N_14151);
and UO_678 (O_678,N_14564,N_14342);
or UO_679 (O_679,N_14809,N_14675);
and UO_680 (O_680,N_14255,N_14665);
nand UO_681 (O_681,N_14006,N_14409);
or UO_682 (O_682,N_14325,N_14334);
or UO_683 (O_683,N_14513,N_14168);
xnor UO_684 (O_684,N_14249,N_14040);
nand UO_685 (O_685,N_14970,N_14927);
or UO_686 (O_686,N_14184,N_14513);
nor UO_687 (O_687,N_14171,N_14721);
or UO_688 (O_688,N_14419,N_14341);
and UO_689 (O_689,N_14907,N_14566);
xnor UO_690 (O_690,N_14412,N_14125);
nor UO_691 (O_691,N_14346,N_14156);
nor UO_692 (O_692,N_14720,N_14321);
or UO_693 (O_693,N_14875,N_14989);
nor UO_694 (O_694,N_14360,N_14653);
and UO_695 (O_695,N_14681,N_14215);
nor UO_696 (O_696,N_14305,N_14147);
nand UO_697 (O_697,N_14348,N_14166);
and UO_698 (O_698,N_14944,N_14149);
nand UO_699 (O_699,N_14051,N_14813);
or UO_700 (O_700,N_14056,N_14657);
or UO_701 (O_701,N_14239,N_14232);
nand UO_702 (O_702,N_14113,N_14696);
xnor UO_703 (O_703,N_14790,N_14579);
nand UO_704 (O_704,N_14976,N_14963);
nand UO_705 (O_705,N_14747,N_14362);
and UO_706 (O_706,N_14652,N_14889);
or UO_707 (O_707,N_14532,N_14878);
nand UO_708 (O_708,N_14217,N_14259);
nand UO_709 (O_709,N_14872,N_14318);
and UO_710 (O_710,N_14751,N_14241);
nor UO_711 (O_711,N_14090,N_14831);
nand UO_712 (O_712,N_14074,N_14068);
and UO_713 (O_713,N_14162,N_14429);
xnor UO_714 (O_714,N_14899,N_14173);
xnor UO_715 (O_715,N_14266,N_14130);
xor UO_716 (O_716,N_14988,N_14004);
xor UO_717 (O_717,N_14790,N_14184);
nand UO_718 (O_718,N_14316,N_14313);
and UO_719 (O_719,N_14846,N_14106);
nand UO_720 (O_720,N_14517,N_14798);
nand UO_721 (O_721,N_14516,N_14765);
and UO_722 (O_722,N_14568,N_14871);
nand UO_723 (O_723,N_14393,N_14450);
or UO_724 (O_724,N_14966,N_14201);
or UO_725 (O_725,N_14394,N_14978);
nand UO_726 (O_726,N_14126,N_14837);
nand UO_727 (O_727,N_14255,N_14356);
nand UO_728 (O_728,N_14059,N_14924);
and UO_729 (O_729,N_14300,N_14530);
nand UO_730 (O_730,N_14849,N_14020);
and UO_731 (O_731,N_14842,N_14454);
nand UO_732 (O_732,N_14550,N_14760);
nor UO_733 (O_733,N_14184,N_14683);
nor UO_734 (O_734,N_14896,N_14846);
or UO_735 (O_735,N_14531,N_14692);
and UO_736 (O_736,N_14060,N_14559);
nor UO_737 (O_737,N_14183,N_14582);
or UO_738 (O_738,N_14836,N_14626);
nand UO_739 (O_739,N_14813,N_14780);
and UO_740 (O_740,N_14815,N_14874);
or UO_741 (O_741,N_14693,N_14086);
xnor UO_742 (O_742,N_14416,N_14013);
or UO_743 (O_743,N_14661,N_14668);
nor UO_744 (O_744,N_14111,N_14363);
or UO_745 (O_745,N_14922,N_14796);
and UO_746 (O_746,N_14190,N_14210);
nand UO_747 (O_747,N_14621,N_14530);
and UO_748 (O_748,N_14627,N_14275);
xnor UO_749 (O_749,N_14849,N_14381);
nand UO_750 (O_750,N_14735,N_14006);
nand UO_751 (O_751,N_14589,N_14930);
xnor UO_752 (O_752,N_14862,N_14607);
nand UO_753 (O_753,N_14429,N_14133);
or UO_754 (O_754,N_14703,N_14334);
nor UO_755 (O_755,N_14303,N_14328);
nor UO_756 (O_756,N_14769,N_14478);
nand UO_757 (O_757,N_14284,N_14034);
nor UO_758 (O_758,N_14285,N_14370);
or UO_759 (O_759,N_14815,N_14576);
nor UO_760 (O_760,N_14776,N_14088);
nor UO_761 (O_761,N_14226,N_14312);
xnor UO_762 (O_762,N_14661,N_14275);
and UO_763 (O_763,N_14986,N_14512);
nor UO_764 (O_764,N_14340,N_14735);
or UO_765 (O_765,N_14434,N_14448);
nor UO_766 (O_766,N_14123,N_14600);
nand UO_767 (O_767,N_14973,N_14544);
nor UO_768 (O_768,N_14035,N_14379);
or UO_769 (O_769,N_14283,N_14717);
and UO_770 (O_770,N_14914,N_14692);
nand UO_771 (O_771,N_14067,N_14052);
nand UO_772 (O_772,N_14198,N_14735);
nor UO_773 (O_773,N_14263,N_14098);
nor UO_774 (O_774,N_14359,N_14409);
nand UO_775 (O_775,N_14857,N_14840);
or UO_776 (O_776,N_14339,N_14425);
nor UO_777 (O_777,N_14770,N_14380);
nor UO_778 (O_778,N_14722,N_14069);
nand UO_779 (O_779,N_14130,N_14572);
nor UO_780 (O_780,N_14985,N_14139);
nor UO_781 (O_781,N_14489,N_14283);
and UO_782 (O_782,N_14665,N_14208);
or UO_783 (O_783,N_14056,N_14604);
or UO_784 (O_784,N_14548,N_14868);
or UO_785 (O_785,N_14339,N_14383);
nand UO_786 (O_786,N_14564,N_14212);
nor UO_787 (O_787,N_14823,N_14167);
xnor UO_788 (O_788,N_14518,N_14199);
nor UO_789 (O_789,N_14709,N_14654);
nand UO_790 (O_790,N_14109,N_14295);
nor UO_791 (O_791,N_14605,N_14698);
and UO_792 (O_792,N_14387,N_14749);
and UO_793 (O_793,N_14540,N_14843);
or UO_794 (O_794,N_14725,N_14255);
and UO_795 (O_795,N_14746,N_14318);
nor UO_796 (O_796,N_14677,N_14555);
nand UO_797 (O_797,N_14739,N_14132);
nor UO_798 (O_798,N_14635,N_14259);
and UO_799 (O_799,N_14812,N_14889);
nor UO_800 (O_800,N_14943,N_14035);
or UO_801 (O_801,N_14241,N_14547);
nor UO_802 (O_802,N_14026,N_14244);
and UO_803 (O_803,N_14518,N_14840);
xnor UO_804 (O_804,N_14842,N_14739);
or UO_805 (O_805,N_14075,N_14788);
or UO_806 (O_806,N_14542,N_14698);
nor UO_807 (O_807,N_14658,N_14274);
xor UO_808 (O_808,N_14980,N_14130);
nor UO_809 (O_809,N_14313,N_14015);
nor UO_810 (O_810,N_14476,N_14478);
nor UO_811 (O_811,N_14773,N_14612);
and UO_812 (O_812,N_14656,N_14577);
nor UO_813 (O_813,N_14933,N_14231);
and UO_814 (O_814,N_14688,N_14408);
and UO_815 (O_815,N_14709,N_14097);
xnor UO_816 (O_816,N_14702,N_14890);
nand UO_817 (O_817,N_14306,N_14530);
nor UO_818 (O_818,N_14816,N_14046);
or UO_819 (O_819,N_14485,N_14271);
nand UO_820 (O_820,N_14174,N_14068);
xor UO_821 (O_821,N_14530,N_14645);
nor UO_822 (O_822,N_14442,N_14414);
nor UO_823 (O_823,N_14686,N_14170);
xnor UO_824 (O_824,N_14372,N_14826);
nand UO_825 (O_825,N_14382,N_14637);
nor UO_826 (O_826,N_14895,N_14250);
or UO_827 (O_827,N_14365,N_14874);
and UO_828 (O_828,N_14998,N_14528);
and UO_829 (O_829,N_14708,N_14639);
nor UO_830 (O_830,N_14614,N_14854);
nor UO_831 (O_831,N_14336,N_14913);
nor UO_832 (O_832,N_14489,N_14364);
nand UO_833 (O_833,N_14675,N_14310);
xnor UO_834 (O_834,N_14449,N_14194);
and UO_835 (O_835,N_14755,N_14691);
xnor UO_836 (O_836,N_14784,N_14968);
nand UO_837 (O_837,N_14535,N_14320);
nand UO_838 (O_838,N_14241,N_14951);
nand UO_839 (O_839,N_14037,N_14172);
or UO_840 (O_840,N_14428,N_14988);
and UO_841 (O_841,N_14504,N_14218);
or UO_842 (O_842,N_14126,N_14867);
or UO_843 (O_843,N_14418,N_14962);
or UO_844 (O_844,N_14487,N_14026);
and UO_845 (O_845,N_14785,N_14631);
and UO_846 (O_846,N_14374,N_14443);
nor UO_847 (O_847,N_14456,N_14188);
and UO_848 (O_848,N_14651,N_14529);
nor UO_849 (O_849,N_14256,N_14026);
and UO_850 (O_850,N_14785,N_14246);
or UO_851 (O_851,N_14625,N_14611);
nand UO_852 (O_852,N_14140,N_14359);
nor UO_853 (O_853,N_14797,N_14996);
or UO_854 (O_854,N_14534,N_14994);
xor UO_855 (O_855,N_14168,N_14378);
or UO_856 (O_856,N_14005,N_14287);
nand UO_857 (O_857,N_14594,N_14145);
or UO_858 (O_858,N_14876,N_14463);
or UO_859 (O_859,N_14238,N_14913);
and UO_860 (O_860,N_14995,N_14833);
or UO_861 (O_861,N_14588,N_14124);
and UO_862 (O_862,N_14816,N_14776);
nand UO_863 (O_863,N_14920,N_14334);
and UO_864 (O_864,N_14134,N_14248);
xnor UO_865 (O_865,N_14847,N_14503);
and UO_866 (O_866,N_14599,N_14034);
nand UO_867 (O_867,N_14202,N_14435);
nand UO_868 (O_868,N_14631,N_14474);
and UO_869 (O_869,N_14860,N_14561);
or UO_870 (O_870,N_14285,N_14553);
and UO_871 (O_871,N_14931,N_14960);
nand UO_872 (O_872,N_14609,N_14486);
nand UO_873 (O_873,N_14584,N_14800);
or UO_874 (O_874,N_14467,N_14206);
nand UO_875 (O_875,N_14374,N_14603);
nor UO_876 (O_876,N_14253,N_14805);
or UO_877 (O_877,N_14938,N_14386);
or UO_878 (O_878,N_14598,N_14668);
xnor UO_879 (O_879,N_14950,N_14505);
and UO_880 (O_880,N_14015,N_14390);
nor UO_881 (O_881,N_14079,N_14908);
nor UO_882 (O_882,N_14746,N_14760);
nor UO_883 (O_883,N_14132,N_14384);
or UO_884 (O_884,N_14242,N_14496);
and UO_885 (O_885,N_14719,N_14989);
nor UO_886 (O_886,N_14473,N_14468);
or UO_887 (O_887,N_14360,N_14176);
or UO_888 (O_888,N_14785,N_14709);
nand UO_889 (O_889,N_14773,N_14053);
or UO_890 (O_890,N_14083,N_14203);
or UO_891 (O_891,N_14467,N_14639);
nand UO_892 (O_892,N_14119,N_14842);
nor UO_893 (O_893,N_14283,N_14093);
nor UO_894 (O_894,N_14374,N_14503);
xor UO_895 (O_895,N_14535,N_14001);
nor UO_896 (O_896,N_14325,N_14065);
nand UO_897 (O_897,N_14964,N_14896);
nand UO_898 (O_898,N_14051,N_14018);
and UO_899 (O_899,N_14198,N_14184);
nor UO_900 (O_900,N_14465,N_14003);
or UO_901 (O_901,N_14211,N_14279);
nand UO_902 (O_902,N_14072,N_14589);
nand UO_903 (O_903,N_14421,N_14578);
xnor UO_904 (O_904,N_14466,N_14526);
nor UO_905 (O_905,N_14027,N_14579);
nand UO_906 (O_906,N_14184,N_14544);
and UO_907 (O_907,N_14107,N_14544);
or UO_908 (O_908,N_14769,N_14669);
and UO_909 (O_909,N_14119,N_14733);
and UO_910 (O_910,N_14268,N_14350);
and UO_911 (O_911,N_14905,N_14945);
or UO_912 (O_912,N_14639,N_14392);
xor UO_913 (O_913,N_14039,N_14978);
and UO_914 (O_914,N_14916,N_14502);
and UO_915 (O_915,N_14384,N_14262);
or UO_916 (O_916,N_14198,N_14988);
xor UO_917 (O_917,N_14775,N_14048);
nand UO_918 (O_918,N_14344,N_14338);
or UO_919 (O_919,N_14561,N_14386);
nand UO_920 (O_920,N_14249,N_14651);
and UO_921 (O_921,N_14082,N_14042);
xor UO_922 (O_922,N_14666,N_14801);
and UO_923 (O_923,N_14015,N_14336);
and UO_924 (O_924,N_14153,N_14798);
and UO_925 (O_925,N_14383,N_14848);
nor UO_926 (O_926,N_14351,N_14061);
xnor UO_927 (O_927,N_14745,N_14376);
nand UO_928 (O_928,N_14296,N_14454);
nand UO_929 (O_929,N_14708,N_14690);
nor UO_930 (O_930,N_14686,N_14899);
and UO_931 (O_931,N_14579,N_14656);
and UO_932 (O_932,N_14459,N_14912);
nor UO_933 (O_933,N_14633,N_14154);
nor UO_934 (O_934,N_14080,N_14998);
or UO_935 (O_935,N_14926,N_14627);
xnor UO_936 (O_936,N_14199,N_14615);
nor UO_937 (O_937,N_14944,N_14203);
and UO_938 (O_938,N_14641,N_14223);
nor UO_939 (O_939,N_14258,N_14750);
or UO_940 (O_940,N_14589,N_14822);
or UO_941 (O_941,N_14497,N_14597);
nand UO_942 (O_942,N_14328,N_14825);
or UO_943 (O_943,N_14628,N_14292);
nor UO_944 (O_944,N_14232,N_14450);
nand UO_945 (O_945,N_14370,N_14337);
nand UO_946 (O_946,N_14856,N_14010);
xnor UO_947 (O_947,N_14072,N_14521);
nand UO_948 (O_948,N_14378,N_14883);
nand UO_949 (O_949,N_14480,N_14743);
xor UO_950 (O_950,N_14964,N_14180);
nand UO_951 (O_951,N_14181,N_14335);
nand UO_952 (O_952,N_14321,N_14826);
or UO_953 (O_953,N_14636,N_14595);
nand UO_954 (O_954,N_14313,N_14554);
xnor UO_955 (O_955,N_14671,N_14328);
or UO_956 (O_956,N_14574,N_14358);
and UO_957 (O_957,N_14145,N_14118);
xor UO_958 (O_958,N_14225,N_14083);
nor UO_959 (O_959,N_14657,N_14633);
or UO_960 (O_960,N_14694,N_14189);
or UO_961 (O_961,N_14534,N_14561);
nor UO_962 (O_962,N_14396,N_14607);
or UO_963 (O_963,N_14753,N_14915);
and UO_964 (O_964,N_14348,N_14735);
nor UO_965 (O_965,N_14845,N_14302);
or UO_966 (O_966,N_14776,N_14631);
nand UO_967 (O_967,N_14165,N_14670);
nor UO_968 (O_968,N_14347,N_14993);
nor UO_969 (O_969,N_14541,N_14594);
nand UO_970 (O_970,N_14522,N_14334);
nand UO_971 (O_971,N_14953,N_14599);
or UO_972 (O_972,N_14570,N_14480);
nor UO_973 (O_973,N_14963,N_14190);
nand UO_974 (O_974,N_14901,N_14063);
or UO_975 (O_975,N_14615,N_14045);
xor UO_976 (O_976,N_14432,N_14222);
and UO_977 (O_977,N_14690,N_14903);
nand UO_978 (O_978,N_14519,N_14857);
or UO_979 (O_979,N_14293,N_14895);
nor UO_980 (O_980,N_14468,N_14425);
xor UO_981 (O_981,N_14054,N_14479);
and UO_982 (O_982,N_14833,N_14944);
and UO_983 (O_983,N_14428,N_14883);
nand UO_984 (O_984,N_14514,N_14304);
and UO_985 (O_985,N_14093,N_14412);
or UO_986 (O_986,N_14490,N_14706);
and UO_987 (O_987,N_14257,N_14470);
and UO_988 (O_988,N_14255,N_14690);
nand UO_989 (O_989,N_14733,N_14463);
nor UO_990 (O_990,N_14600,N_14284);
nor UO_991 (O_991,N_14677,N_14521);
and UO_992 (O_992,N_14463,N_14272);
nand UO_993 (O_993,N_14577,N_14242);
nor UO_994 (O_994,N_14497,N_14421);
or UO_995 (O_995,N_14315,N_14296);
and UO_996 (O_996,N_14447,N_14272);
and UO_997 (O_997,N_14472,N_14781);
and UO_998 (O_998,N_14588,N_14755);
and UO_999 (O_999,N_14118,N_14401);
or UO_1000 (O_1000,N_14901,N_14622);
nor UO_1001 (O_1001,N_14291,N_14073);
nor UO_1002 (O_1002,N_14053,N_14094);
or UO_1003 (O_1003,N_14789,N_14716);
nand UO_1004 (O_1004,N_14000,N_14806);
nand UO_1005 (O_1005,N_14319,N_14204);
nor UO_1006 (O_1006,N_14190,N_14745);
or UO_1007 (O_1007,N_14778,N_14190);
or UO_1008 (O_1008,N_14371,N_14157);
nand UO_1009 (O_1009,N_14054,N_14160);
and UO_1010 (O_1010,N_14727,N_14943);
nand UO_1011 (O_1011,N_14315,N_14425);
or UO_1012 (O_1012,N_14533,N_14578);
or UO_1013 (O_1013,N_14101,N_14548);
nor UO_1014 (O_1014,N_14447,N_14945);
nand UO_1015 (O_1015,N_14431,N_14824);
xnor UO_1016 (O_1016,N_14013,N_14561);
and UO_1017 (O_1017,N_14271,N_14967);
nand UO_1018 (O_1018,N_14475,N_14827);
and UO_1019 (O_1019,N_14369,N_14923);
nand UO_1020 (O_1020,N_14628,N_14742);
nand UO_1021 (O_1021,N_14990,N_14147);
nand UO_1022 (O_1022,N_14748,N_14184);
and UO_1023 (O_1023,N_14522,N_14787);
or UO_1024 (O_1024,N_14929,N_14138);
nor UO_1025 (O_1025,N_14548,N_14669);
or UO_1026 (O_1026,N_14173,N_14176);
or UO_1027 (O_1027,N_14140,N_14130);
nor UO_1028 (O_1028,N_14903,N_14221);
nand UO_1029 (O_1029,N_14116,N_14619);
nor UO_1030 (O_1030,N_14633,N_14286);
and UO_1031 (O_1031,N_14915,N_14127);
nand UO_1032 (O_1032,N_14457,N_14110);
or UO_1033 (O_1033,N_14282,N_14912);
nand UO_1034 (O_1034,N_14801,N_14631);
nand UO_1035 (O_1035,N_14769,N_14771);
nand UO_1036 (O_1036,N_14320,N_14793);
or UO_1037 (O_1037,N_14531,N_14429);
nand UO_1038 (O_1038,N_14302,N_14957);
nor UO_1039 (O_1039,N_14268,N_14652);
and UO_1040 (O_1040,N_14795,N_14018);
nand UO_1041 (O_1041,N_14038,N_14576);
nand UO_1042 (O_1042,N_14403,N_14814);
nand UO_1043 (O_1043,N_14893,N_14343);
nor UO_1044 (O_1044,N_14523,N_14834);
and UO_1045 (O_1045,N_14155,N_14441);
xnor UO_1046 (O_1046,N_14920,N_14765);
nand UO_1047 (O_1047,N_14899,N_14514);
nor UO_1048 (O_1048,N_14873,N_14892);
nor UO_1049 (O_1049,N_14884,N_14549);
or UO_1050 (O_1050,N_14662,N_14557);
and UO_1051 (O_1051,N_14993,N_14056);
nor UO_1052 (O_1052,N_14716,N_14951);
or UO_1053 (O_1053,N_14259,N_14928);
or UO_1054 (O_1054,N_14767,N_14077);
and UO_1055 (O_1055,N_14094,N_14266);
xnor UO_1056 (O_1056,N_14789,N_14462);
xnor UO_1057 (O_1057,N_14505,N_14641);
and UO_1058 (O_1058,N_14082,N_14580);
nor UO_1059 (O_1059,N_14966,N_14102);
or UO_1060 (O_1060,N_14157,N_14690);
or UO_1061 (O_1061,N_14247,N_14530);
nand UO_1062 (O_1062,N_14982,N_14658);
xnor UO_1063 (O_1063,N_14416,N_14692);
and UO_1064 (O_1064,N_14801,N_14507);
or UO_1065 (O_1065,N_14085,N_14867);
or UO_1066 (O_1066,N_14860,N_14785);
nor UO_1067 (O_1067,N_14140,N_14351);
nor UO_1068 (O_1068,N_14571,N_14520);
or UO_1069 (O_1069,N_14442,N_14739);
nor UO_1070 (O_1070,N_14249,N_14297);
nor UO_1071 (O_1071,N_14931,N_14634);
or UO_1072 (O_1072,N_14050,N_14013);
or UO_1073 (O_1073,N_14402,N_14123);
nand UO_1074 (O_1074,N_14404,N_14429);
or UO_1075 (O_1075,N_14982,N_14200);
nor UO_1076 (O_1076,N_14025,N_14304);
and UO_1077 (O_1077,N_14024,N_14444);
nor UO_1078 (O_1078,N_14787,N_14405);
and UO_1079 (O_1079,N_14427,N_14029);
nand UO_1080 (O_1080,N_14527,N_14397);
nor UO_1081 (O_1081,N_14639,N_14191);
or UO_1082 (O_1082,N_14998,N_14855);
or UO_1083 (O_1083,N_14710,N_14186);
xnor UO_1084 (O_1084,N_14817,N_14372);
nor UO_1085 (O_1085,N_14829,N_14975);
nand UO_1086 (O_1086,N_14838,N_14196);
or UO_1087 (O_1087,N_14506,N_14341);
nor UO_1088 (O_1088,N_14299,N_14440);
and UO_1089 (O_1089,N_14322,N_14564);
nand UO_1090 (O_1090,N_14056,N_14723);
and UO_1091 (O_1091,N_14425,N_14967);
nand UO_1092 (O_1092,N_14952,N_14678);
and UO_1093 (O_1093,N_14308,N_14171);
and UO_1094 (O_1094,N_14992,N_14680);
or UO_1095 (O_1095,N_14429,N_14292);
xor UO_1096 (O_1096,N_14683,N_14213);
and UO_1097 (O_1097,N_14621,N_14544);
nor UO_1098 (O_1098,N_14992,N_14651);
and UO_1099 (O_1099,N_14186,N_14930);
or UO_1100 (O_1100,N_14826,N_14863);
and UO_1101 (O_1101,N_14316,N_14181);
nor UO_1102 (O_1102,N_14213,N_14233);
or UO_1103 (O_1103,N_14403,N_14359);
nand UO_1104 (O_1104,N_14773,N_14704);
or UO_1105 (O_1105,N_14595,N_14195);
nand UO_1106 (O_1106,N_14190,N_14612);
nor UO_1107 (O_1107,N_14483,N_14119);
or UO_1108 (O_1108,N_14080,N_14694);
nor UO_1109 (O_1109,N_14985,N_14405);
nor UO_1110 (O_1110,N_14271,N_14331);
nand UO_1111 (O_1111,N_14936,N_14947);
and UO_1112 (O_1112,N_14748,N_14454);
nor UO_1113 (O_1113,N_14102,N_14164);
and UO_1114 (O_1114,N_14200,N_14501);
nand UO_1115 (O_1115,N_14197,N_14234);
and UO_1116 (O_1116,N_14737,N_14499);
and UO_1117 (O_1117,N_14871,N_14862);
or UO_1118 (O_1118,N_14495,N_14386);
and UO_1119 (O_1119,N_14476,N_14330);
or UO_1120 (O_1120,N_14856,N_14431);
or UO_1121 (O_1121,N_14355,N_14318);
and UO_1122 (O_1122,N_14713,N_14059);
and UO_1123 (O_1123,N_14428,N_14348);
and UO_1124 (O_1124,N_14640,N_14868);
nor UO_1125 (O_1125,N_14658,N_14444);
nand UO_1126 (O_1126,N_14405,N_14077);
or UO_1127 (O_1127,N_14140,N_14343);
nor UO_1128 (O_1128,N_14815,N_14991);
or UO_1129 (O_1129,N_14846,N_14166);
nor UO_1130 (O_1130,N_14368,N_14714);
or UO_1131 (O_1131,N_14423,N_14925);
xnor UO_1132 (O_1132,N_14697,N_14689);
xor UO_1133 (O_1133,N_14743,N_14183);
and UO_1134 (O_1134,N_14167,N_14614);
or UO_1135 (O_1135,N_14326,N_14445);
nand UO_1136 (O_1136,N_14010,N_14621);
or UO_1137 (O_1137,N_14135,N_14058);
xor UO_1138 (O_1138,N_14355,N_14298);
nand UO_1139 (O_1139,N_14851,N_14642);
or UO_1140 (O_1140,N_14948,N_14044);
xor UO_1141 (O_1141,N_14291,N_14565);
or UO_1142 (O_1142,N_14218,N_14097);
nor UO_1143 (O_1143,N_14478,N_14879);
nor UO_1144 (O_1144,N_14320,N_14013);
or UO_1145 (O_1145,N_14406,N_14204);
nand UO_1146 (O_1146,N_14738,N_14801);
and UO_1147 (O_1147,N_14391,N_14064);
and UO_1148 (O_1148,N_14548,N_14966);
nand UO_1149 (O_1149,N_14300,N_14808);
nor UO_1150 (O_1150,N_14975,N_14024);
nand UO_1151 (O_1151,N_14197,N_14965);
nor UO_1152 (O_1152,N_14925,N_14354);
nand UO_1153 (O_1153,N_14821,N_14178);
and UO_1154 (O_1154,N_14072,N_14453);
nand UO_1155 (O_1155,N_14447,N_14644);
nand UO_1156 (O_1156,N_14956,N_14341);
nand UO_1157 (O_1157,N_14348,N_14303);
nor UO_1158 (O_1158,N_14302,N_14664);
and UO_1159 (O_1159,N_14275,N_14023);
or UO_1160 (O_1160,N_14871,N_14906);
or UO_1161 (O_1161,N_14189,N_14079);
nand UO_1162 (O_1162,N_14562,N_14997);
or UO_1163 (O_1163,N_14002,N_14507);
nand UO_1164 (O_1164,N_14226,N_14029);
or UO_1165 (O_1165,N_14187,N_14007);
or UO_1166 (O_1166,N_14599,N_14617);
nand UO_1167 (O_1167,N_14594,N_14472);
or UO_1168 (O_1168,N_14387,N_14550);
nand UO_1169 (O_1169,N_14346,N_14937);
xnor UO_1170 (O_1170,N_14682,N_14697);
xor UO_1171 (O_1171,N_14973,N_14721);
nand UO_1172 (O_1172,N_14593,N_14962);
or UO_1173 (O_1173,N_14597,N_14209);
or UO_1174 (O_1174,N_14126,N_14739);
nand UO_1175 (O_1175,N_14499,N_14601);
xnor UO_1176 (O_1176,N_14524,N_14832);
and UO_1177 (O_1177,N_14952,N_14634);
nor UO_1178 (O_1178,N_14148,N_14237);
and UO_1179 (O_1179,N_14982,N_14831);
or UO_1180 (O_1180,N_14197,N_14536);
and UO_1181 (O_1181,N_14912,N_14321);
and UO_1182 (O_1182,N_14145,N_14752);
or UO_1183 (O_1183,N_14869,N_14620);
xor UO_1184 (O_1184,N_14227,N_14232);
nand UO_1185 (O_1185,N_14014,N_14820);
nand UO_1186 (O_1186,N_14718,N_14770);
xor UO_1187 (O_1187,N_14255,N_14525);
or UO_1188 (O_1188,N_14469,N_14769);
or UO_1189 (O_1189,N_14267,N_14652);
nor UO_1190 (O_1190,N_14535,N_14396);
nor UO_1191 (O_1191,N_14136,N_14282);
and UO_1192 (O_1192,N_14861,N_14201);
xor UO_1193 (O_1193,N_14158,N_14381);
nor UO_1194 (O_1194,N_14946,N_14053);
xnor UO_1195 (O_1195,N_14073,N_14598);
and UO_1196 (O_1196,N_14346,N_14362);
or UO_1197 (O_1197,N_14020,N_14156);
and UO_1198 (O_1198,N_14220,N_14676);
nand UO_1199 (O_1199,N_14021,N_14470);
nand UO_1200 (O_1200,N_14225,N_14541);
nand UO_1201 (O_1201,N_14832,N_14713);
nand UO_1202 (O_1202,N_14826,N_14563);
xor UO_1203 (O_1203,N_14109,N_14256);
and UO_1204 (O_1204,N_14507,N_14373);
xnor UO_1205 (O_1205,N_14850,N_14046);
nor UO_1206 (O_1206,N_14416,N_14588);
nand UO_1207 (O_1207,N_14230,N_14125);
or UO_1208 (O_1208,N_14777,N_14006);
and UO_1209 (O_1209,N_14842,N_14976);
nor UO_1210 (O_1210,N_14206,N_14529);
xor UO_1211 (O_1211,N_14348,N_14001);
xnor UO_1212 (O_1212,N_14763,N_14801);
or UO_1213 (O_1213,N_14422,N_14420);
nand UO_1214 (O_1214,N_14464,N_14351);
nor UO_1215 (O_1215,N_14484,N_14968);
nand UO_1216 (O_1216,N_14223,N_14464);
nand UO_1217 (O_1217,N_14783,N_14313);
and UO_1218 (O_1218,N_14398,N_14391);
or UO_1219 (O_1219,N_14685,N_14361);
nor UO_1220 (O_1220,N_14233,N_14875);
nand UO_1221 (O_1221,N_14735,N_14657);
and UO_1222 (O_1222,N_14723,N_14716);
nand UO_1223 (O_1223,N_14140,N_14119);
and UO_1224 (O_1224,N_14687,N_14364);
or UO_1225 (O_1225,N_14057,N_14147);
and UO_1226 (O_1226,N_14230,N_14280);
xnor UO_1227 (O_1227,N_14695,N_14820);
nand UO_1228 (O_1228,N_14969,N_14477);
or UO_1229 (O_1229,N_14099,N_14962);
and UO_1230 (O_1230,N_14888,N_14547);
nor UO_1231 (O_1231,N_14952,N_14723);
and UO_1232 (O_1232,N_14787,N_14696);
nor UO_1233 (O_1233,N_14629,N_14020);
nor UO_1234 (O_1234,N_14129,N_14664);
xnor UO_1235 (O_1235,N_14818,N_14761);
and UO_1236 (O_1236,N_14992,N_14006);
or UO_1237 (O_1237,N_14501,N_14926);
and UO_1238 (O_1238,N_14492,N_14870);
and UO_1239 (O_1239,N_14003,N_14405);
and UO_1240 (O_1240,N_14616,N_14596);
and UO_1241 (O_1241,N_14039,N_14999);
xor UO_1242 (O_1242,N_14951,N_14769);
nand UO_1243 (O_1243,N_14028,N_14763);
nand UO_1244 (O_1244,N_14928,N_14026);
or UO_1245 (O_1245,N_14389,N_14308);
or UO_1246 (O_1246,N_14367,N_14094);
or UO_1247 (O_1247,N_14633,N_14617);
and UO_1248 (O_1248,N_14661,N_14925);
nand UO_1249 (O_1249,N_14103,N_14239);
xnor UO_1250 (O_1250,N_14255,N_14608);
nand UO_1251 (O_1251,N_14316,N_14421);
nor UO_1252 (O_1252,N_14892,N_14070);
and UO_1253 (O_1253,N_14251,N_14337);
or UO_1254 (O_1254,N_14496,N_14870);
and UO_1255 (O_1255,N_14767,N_14453);
nand UO_1256 (O_1256,N_14722,N_14619);
or UO_1257 (O_1257,N_14116,N_14682);
and UO_1258 (O_1258,N_14992,N_14930);
nor UO_1259 (O_1259,N_14899,N_14561);
xor UO_1260 (O_1260,N_14369,N_14843);
nor UO_1261 (O_1261,N_14302,N_14192);
nor UO_1262 (O_1262,N_14701,N_14660);
or UO_1263 (O_1263,N_14652,N_14522);
or UO_1264 (O_1264,N_14614,N_14607);
and UO_1265 (O_1265,N_14908,N_14009);
nand UO_1266 (O_1266,N_14185,N_14380);
xnor UO_1267 (O_1267,N_14147,N_14966);
and UO_1268 (O_1268,N_14988,N_14213);
and UO_1269 (O_1269,N_14726,N_14126);
nand UO_1270 (O_1270,N_14682,N_14932);
nand UO_1271 (O_1271,N_14319,N_14695);
and UO_1272 (O_1272,N_14502,N_14074);
xnor UO_1273 (O_1273,N_14029,N_14538);
nand UO_1274 (O_1274,N_14884,N_14546);
nor UO_1275 (O_1275,N_14953,N_14249);
or UO_1276 (O_1276,N_14079,N_14285);
and UO_1277 (O_1277,N_14830,N_14357);
and UO_1278 (O_1278,N_14771,N_14652);
xnor UO_1279 (O_1279,N_14110,N_14451);
and UO_1280 (O_1280,N_14678,N_14129);
or UO_1281 (O_1281,N_14939,N_14125);
nor UO_1282 (O_1282,N_14948,N_14685);
or UO_1283 (O_1283,N_14703,N_14199);
nand UO_1284 (O_1284,N_14644,N_14587);
xor UO_1285 (O_1285,N_14970,N_14155);
nor UO_1286 (O_1286,N_14767,N_14700);
xor UO_1287 (O_1287,N_14217,N_14347);
nand UO_1288 (O_1288,N_14336,N_14587);
nor UO_1289 (O_1289,N_14346,N_14171);
nor UO_1290 (O_1290,N_14643,N_14635);
and UO_1291 (O_1291,N_14640,N_14556);
nand UO_1292 (O_1292,N_14940,N_14115);
and UO_1293 (O_1293,N_14963,N_14825);
nor UO_1294 (O_1294,N_14595,N_14156);
nor UO_1295 (O_1295,N_14773,N_14321);
or UO_1296 (O_1296,N_14857,N_14448);
nand UO_1297 (O_1297,N_14468,N_14947);
and UO_1298 (O_1298,N_14407,N_14348);
and UO_1299 (O_1299,N_14676,N_14751);
and UO_1300 (O_1300,N_14689,N_14596);
and UO_1301 (O_1301,N_14838,N_14482);
nand UO_1302 (O_1302,N_14219,N_14941);
nor UO_1303 (O_1303,N_14472,N_14748);
nor UO_1304 (O_1304,N_14040,N_14861);
or UO_1305 (O_1305,N_14590,N_14293);
nand UO_1306 (O_1306,N_14110,N_14194);
and UO_1307 (O_1307,N_14934,N_14815);
and UO_1308 (O_1308,N_14534,N_14010);
and UO_1309 (O_1309,N_14192,N_14350);
nor UO_1310 (O_1310,N_14822,N_14350);
and UO_1311 (O_1311,N_14715,N_14547);
nor UO_1312 (O_1312,N_14645,N_14135);
nand UO_1313 (O_1313,N_14192,N_14029);
or UO_1314 (O_1314,N_14596,N_14344);
nor UO_1315 (O_1315,N_14914,N_14856);
nand UO_1316 (O_1316,N_14328,N_14370);
nand UO_1317 (O_1317,N_14382,N_14782);
and UO_1318 (O_1318,N_14836,N_14164);
nand UO_1319 (O_1319,N_14091,N_14906);
and UO_1320 (O_1320,N_14040,N_14507);
and UO_1321 (O_1321,N_14044,N_14000);
nor UO_1322 (O_1322,N_14068,N_14564);
or UO_1323 (O_1323,N_14368,N_14613);
nor UO_1324 (O_1324,N_14158,N_14512);
nor UO_1325 (O_1325,N_14192,N_14565);
nand UO_1326 (O_1326,N_14449,N_14723);
xnor UO_1327 (O_1327,N_14335,N_14733);
xor UO_1328 (O_1328,N_14098,N_14624);
nand UO_1329 (O_1329,N_14825,N_14199);
or UO_1330 (O_1330,N_14686,N_14492);
or UO_1331 (O_1331,N_14311,N_14612);
nand UO_1332 (O_1332,N_14268,N_14968);
and UO_1333 (O_1333,N_14542,N_14459);
nor UO_1334 (O_1334,N_14844,N_14222);
and UO_1335 (O_1335,N_14977,N_14203);
nor UO_1336 (O_1336,N_14763,N_14792);
and UO_1337 (O_1337,N_14578,N_14422);
or UO_1338 (O_1338,N_14841,N_14725);
and UO_1339 (O_1339,N_14460,N_14016);
xnor UO_1340 (O_1340,N_14206,N_14808);
and UO_1341 (O_1341,N_14948,N_14765);
nor UO_1342 (O_1342,N_14651,N_14234);
and UO_1343 (O_1343,N_14291,N_14101);
nand UO_1344 (O_1344,N_14402,N_14172);
nor UO_1345 (O_1345,N_14765,N_14837);
and UO_1346 (O_1346,N_14381,N_14577);
nand UO_1347 (O_1347,N_14437,N_14343);
and UO_1348 (O_1348,N_14132,N_14194);
xor UO_1349 (O_1349,N_14038,N_14202);
xor UO_1350 (O_1350,N_14347,N_14152);
and UO_1351 (O_1351,N_14430,N_14681);
xor UO_1352 (O_1352,N_14287,N_14850);
and UO_1353 (O_1353,N_14173,N_14606);
and UO_1354 (O_1354,N_14152,N_14708);
nor UO_1355 (O_1355,N_14186,N_14168);
and UO_1356 (O_1356,N_14350,N_14808);
and UO_1357 (O_1357,N_14053,N_14406);
nand UO_1358 (O_1358,N_14207,N_14885);
nor UO_1359 (O_1359,N_14924,N_14952);
xnor UO_1360 (O_1360,N_14911,N_14179);
and UO_1361 (O_1361,N_14078,N_14222);
nor UO_1362 (O_1362,N_14098,N_14327);
nand UO_1363 (O_1363,N_14919,N_14791);
and UO_1364 (O_1364,N_14771,N_14789);
or UO_1365 (O_1365,N_14922,N_14051);
nor UO_1366 (O_1366,N_14556,N_14180);
nand UO_1367 (O_1367,N_14132,N_14038);
or UO_1368 (O_1368,N_14576,N_14789);
nor UO_1369 (O_1369,N_14045,N_14180);
and UO_1370 (O_1370,N_14121,N_14932);
nor UO_1371 (O_1371,N_14470,N_14666);
nand UO_1372 (O_1372,N_14571,N_14093);
and UO_1373 (O_1373,N_14507,N_14985);
xnor UO_1374 (O_1374,N_14053,N_14222);
or UO_1375 (O_1375,N_14101,N_14583);
nand UO_1376 (O_1376,N_14197,N_14938);
xnor UO_1377 (O_1377,N_14840,N_14105);
xor UO_1378 (O_1378,N_14859,N_14246);
nand UO_1379 (O_1379,N_14767,N_14617);
nor UO_1380 (O_1380,N_14260,N_14418);
nand UO_1381 (O_1381,N_14311,N_14076);
nand UO_1382 (O_1382,N_14883,N_14551);
and UO_1383 (O_1383,N_14060,N_14010);
xor UO_1384 (O_1384,N_14202,N_14928);
or UO_1385 (O_1385,N_14078,N_14375);
nor UO_1386 (O_1386,N_14586,N_14349);
or UO_1387 (O_1387,N_14992,N_14214);
nand UO_1388 (O_1388,N_14768,N_14109);
nand UO_1389 (O_1389,N_14193,N_14756);
nand UO_1390 (O_1390,N_14909,N_14302);
or UO_1391 (O_1391,N_14056,N_14028);
or UO_1392 (O_1392,N_14195,N_14969);
or UO_1393 (O_1393,N_14470,N_14828);
and UO_1394 (O_1394,N_14221,N_14037);
xnor UO_1395 (O_1395,N_14035,N_14785);
nor UO_1396 (O_1396,N_14163,N_14122);
or UO_1397 (O_1397,N_14987,N_14392);
and UO_1398 (O_1398,N_14301,N_14635);
nand UO_1399 (O_1399,N_14481,N_14363);
xor UO_1400 (O_1400,N_14223,N_14937);
nor UO_1401 (O_1401,N_14864,N_14497);
or UO_1402 (O_1402,N_14553,N_14363);
or UO_1403 (O_1403,N_14200,N_14202);
nand UO_1404 (O_1404,N_14830,N_14679);
and UO_1405 (O_1405,N_14277,N_14842);
and UO_1406 (O_1406,N_14299,N_14983);
and UO_1407 (O_1407,N_14777,N_14621);
nor UO_1408 (O_1408,N_14408,N_14449);
xnor UO_1409 (O_1409,N_14500,N_14975);
nand UO_1410 (O_1410,N_14812,N_14390);
nor UO_1411 (O_1411,N_14098,N_14964);
or UO_1412 (O_1412,N_14145,N_14518);
nand UO_1413 (O_1413,N_14558,N_14494);
or UO_1414 (O_1414,N_14171,N_14871);
nand UO_1415 (O_1415,N_14145,N_14655);
and UO_1416 (O_1416,N_14866,N_14385);
nand UO_1417 (O_1417,N_14111,N_14516);
nand UO_1418 (O_1418,N_14825,N_14275);
nor UO_1419 (O_1419,N_14697,N_14772);
nor UO_1420 (O_1420,N_14400,N_14624);
nand UO_1421 (O_1421,N_14210,N_14140);
and UO_1422 (O_1422,N_14072,N_14937);
nor UO_1423 (O_1423,N_14721,N_14822);
or UO_1424 (O_1424,N_14663,N_14060);
nand UO_1425 (O_1425,N_14037,N_14734);
nor UO_1426 (O_1426,N_14439,N_14330);
nor UO_1427 (O_1427,N_14748,N_14544);
or UO_1428 (O_1428,N_14226,N_14339);
xnor UO_1429 (O_1429,N_14401,N_14551);
or UO_1430 (O_1430,N_14428,N_14696);
xnor UO_1431 (O_1431,N_14609,N_14763);
nor UO_1432 (O_1432,N_14447,N_14710);
and UO_1433 (O_1433,N_14176,N_14128);
nor UO_1434 (O_1434,N_14833,N_14819);
or UO_1435 (O_1435,N_14267,N_14629);
nand UO_1436 (O_1436,N_14947,N_14651);
nor UO_1437 (O_1437,N_14721,N_14291);
nand UO_1438 (O_1438,N_14193,N_14724);
and UO_1439 (O_1439,N_14348,N_14696);
or UO_1440 (O_1440,N_14055,N_14355);
xnor UO_1441 (O_1441,N_14614,N_14550);
or UO_1442 (O_1442,N_14317,N_14878);
or UO_1443 (O_1443,N_14660,N_14781);
nor UO_1444 (O_1444,N_14032,N_14212);
and UO_1445 (O_1445,N_14894,N_14444);
nand UO_1446 (O_1446,N_14231,N_14021);
nand UO_1447 (O_1447,N_14908,N_14514);
or UO_1448 (O_1448,N_14903,N_14508);
nand UO_1449 (O_1449,N_14015,N_14131);
nor UO_1450 (O_1450,N_14925,N_14511);
or UO_1451 (O_1451,N_14749,N_14326);
nand UO_1452 (O_1452,N_14310,N_14084);
or UO_1453 (O_1453,N_14747,N_14665);
or UO_1454 (O_1454,N_14066,N_14275);
and UO_1455 (O_1455,N_14296,N_14527);
and UO_1456 (O_1456,N_14483,N_14354);
or UO_1457 (O_1457,N_14506,N_14858);
nand UO_1458 (O_1458,N_14648,N_14392);
and UO_1459 (O_1459,N_14013,N_14686);
nand UO_1460 (O_1460,N_14916,N_14267);
nand UO_1461 (O_1461,N_14293,N_14819);
nand UO_1462 (O_1462,N_14087,N_14163);
xor UO_1463 (O_1463,N_14169,N_14154);
nor UO_1464 (O_1464,N_14038,N_14480);
or UO_1465 (O_1465,N_14627,N_14788);
and UO_1466 (O_1466,N_14289,N_14627);
nand UO_1467 (O_1467,N_14344,N_14536);
and UO_1468 (O_1468,N_14949,N_14804);
or UO_1469 (O_1469,N_14605,N_14551);
or UO_1470 (O_1470,N_14370,N_14645);
nand UO_1471 (O_1471,N_14459,N_14616);
nor UO_1472 (O_1472,N_14156,N_14250);
nor UO_1473 (O_1473,N_14134,N_14581);
nor UO_1474 (O_1474,N_14617,N_14818);
and UO_1475 (O_1475,N_14066,N_14761);
and UO_1476 (O_1476,N_14364,N_14699);
nand UO_1477 (O_1477,N_14063,N_14167);
nand UO_1478 (O_1478,N_14745,N_14736);
xnor UO_1479 (O_1479,N_14457,N_14518);
or UO_1480 (O_1480,N_14594,N_14828);
or UO_1481 (O_1481,N_14873,N_14030);
nor UO_1482 (O_1482,N_14527,N_14766);
nor UO_1483 (O_1483,N_14073,N_14145);
or UO_1484 (O_1484,N_14457,N_14487);
nor UO_1485 (O_1485,N_14628,N_14001);
and UO_1486 (O_1486,N_14365,N_14207);
or UO_1487 (O_1487,N_14219,N_14900);
and UO_1488 (O_1488,N_14380,N_14062);
and UO_1489 (O_1489,N_14349,N_14654);
xnor UO_1490 (O_1490,N_14932,N_14870);
or UO_1491 (O_1491,N_14237,N_14475);
or UO_1492 (O_1492,N_14877,N_14374);
and UO_1493 (O_1493,N_14120,N_14671);
nand UO_1494 (O_1494,N_14288,N_14783);
or UO_1495 (O_1495,N_14570,N_14308);
and UO_1496 (O_1496,N_14101,N_14451);
nor UO_1497 (O_1497,N_14950,N_14031);
nor UO_1498 (O_1498,N_14160,N_14268);
nor UO_1499 (O_1499,N_14519,N_14647);
or UO_1500 (O_1500,N_14927,N_14035);
and UO_1501 (O_1501,N_14356,N_14499);
or UO_1502 (O_1502,N_14205,N_14021);
and UO_1503 (O_1503,N_14252,N_14464);
nor UO_1504 (O_1504,N_14523,N_14356);
xor UO_1505 (O_1505,N_14788,N_14223);
nor UO_1506 (O_1506,N_14246,N_14022);
nor UO_1507 (O_1507,N_14221,N_14665);
and UO_1508 (O_1508,N_14875,N_14247);
nor UO_1509 (O_1509,N_14616,N_14590);
and UO_1510 (O_1510,N_14816,N_14763);
and UO_1511 (O_1511,N_14343,N_14641);
or UO_1512 (O_1512,N_14383,N_14238);
and UO_1513 (O_1513,N_14693,N_14590);
or UO_1514 (O_1514,N_14580,N_14826);
or UO_1515 (O_1515,N_14053,N_14399);
nor UO_1516 (O_1516,N_14020,N_14869);
and UO_1517 (O_1517,N_14005,N_14668);
and UO_1518 (O_1518,N_14027,N_14765);
nand UO_1519 (O_1519,N_14953,N_14768);
and UO_1520 (O_1520,N_14423,N_14555);
xnor UO_1521 (O_1521,N_14484,N_14368);
or UO_1522 (O_1522,N_14034,N_14906);
xnor UO_1523 (O_1523,N_14272,N_14163);
or UO_1524 (O_1524,N_14102,N_14194);
nor UO_1525 (O_1525,N_14761,N_14190);
nor UO_1526 (O_1526,N_14917,N_14082);
nand UO_1527 (O_1527,N_14259,N_14160);
and UO_1528 (O_1528,N_14974,N_14487);
nand UO_1529 (O_1529,N_14434,N_14594);
and UO_1530 (O_1530,N_14494,N_14533);
and UO_1531 (O_1531,N_14898,N_14613);
xnor UO_1532 (O_1532,N_14199,N_14831);
or UO_1533 (O_1533,N_14726,N_14749);
xnor UO_1534 (O_1534,N_14524,N_14163);
nor UO_1535 (O_1535,N_14312,N_14958);
nor UO_1536 (O_1536,N_14912,N_14447);
and UO_1537 (O_1537,N_14045,N_14235);
or UO_1538 (O_1538,N_14058,N_14059);
nor UO_1539 (O_1539,N_14103,N_14853);
nor UO_1540 (O_1540,N_14052,N_14670);
and UO_1541 (O_1541,N_14457,N_14059);
nor UO_1542 (O_1542,N_14719,N_14980);
and UO_1543 (O_1543,N_14262,N_14069);
nor UO_1544 (O_1544,N_14408,N_14192);
or UO_1545 (O_1545,N_14957,N_14391);
xor UO_1546 (O_1546,N_14904,N_14536);
nor UO_1547 (O_1547,N_14668,N_14307);
nand UO_1548 (O_1548,N_14429,N_14718);
and UO_1549 (O_1549,N_14006,N_14872);
nand UO_1550 (O_1550,N_14928,N_14801);
xor UO_1551 (O_1551,N_14781,N_14507);
and UO_1552 (O_1552,N_14811,N_14153);
nand UO_1553 (O_1553,N_14696,N_14037);
and UO_1554 (O_1554,N_14471,N_14889);
or UO_1555 (O_1555,N_14712,N_14287);
or UO_1556 (O_1556,N_14327,N_14160);
nor UO_1557 (O_1557,N_14608,N_14207);
nand UO_1558 (O_1558,N_14120,N_14816);
and UO_1559 (O_1559,N_14707,N_14959);
nor UO_1560 (O_1560,N_14246,N_14937);
and UO_1561 (O_1561,N_14820,N_14412);
nor UO_1562 (O_1562,N_14783,N_14480);
nor UO_1563 (O_1563,N_14586,N_14915);
and UO_1564 (O_1564,N_14362,N_14518);
nand UO_1565 (O_1565,N_14675,N_14559);
nand UO_1566 (O_1566,N_14640,N_14605);
nand UO_1567 (O_1567,N_14495,N_14550);
or UO_1568 (O_1568,N_14830,N_14285);
nor UO_1569 (O_1569,N_14969,N_14683);
nor UO_1570 (O_1570,N_14673,N_14310);
or UO_1571 (O_1571,N_14793,N_14154);
and UO_1572 (O_1572,N_14929,N_14671);
nand UO_1573 (O_1573,N_14886,N_14251);
or UO_1574 (O_1574,N_14082,N_14777);
or UO_1575 (O_1575,N_14050,N_14875);
and UO_1576 (O_1576,N_14655,N_14079);
and UO_1577 (O_1577,N_14579,N_14751);
and UO_1578 (O_1578,N_14578,N_14961);
or UO_1579 (O_1579,N_14353,N_14672);
nand UO_1580 (O_1580,N_14810,N_14384);
and UO_1581 (O_1581,N_14069,N_14753);
or UO_1582 (O_1582,N_14804,N_14587);
nor UO_1583 (O_1583,N_14668,N_14366);
or UO_1584 (O_1584,N_14471,N_14344);
xor UO_1585 (O_1585,N_14889,N_14552);
nand UO_1586 (O_1586,N_14228,N_14093);
nand UO_1587 (O_1587,N_14077,N_14703);
or UO_1588 (O_1588,N_14515,N_14084);
xor UO_1589 (O_1589,N_14539,N_14503);
or UO_1590 (O_1590,N_14656,N_14506);
nand UO_1591 (O_1591,N_14503,N_14246);
and UO_1592 (O_1592,N_14656,N_14859);
nor UO_1593 (O_1593,N_14462,N_14228);
nand UO_1594 (O_1594,N_14170,N_14210);
nor UO_1595 (O_1595,N_14367,N_14852);
and UO_1596 (O_1596,N_14693,N_14192);
and UO_1597 (O_1597,N_14682,N_14920);
and UO_1598 (O_1598,N_14805,N_14503);
xor UO_1599 (O_1599,N_14263,N_14736);
or UO_1600 (O_1600,N_14314,N_14512);
nand UO_1601 (O_1601,N_14184,N_14101);
and UO_1602 (O_1602,N_14956,N_14353);
and UO_1603 (O_1603,N_14780,N_14716);
nand UO_1604 (O_1604,N_14618,N_14488);
or UO_1605 (O_1605,N_14185,N_14776);
nor UO_1606 (O_1606,N_14065,N_14669);
nor UO_1607 (O_1607,N_14735,N_14677);
nor UO_1608 (O_1608,N_14436,N_14497);
xor UO_1609 (O_1609,N_14167,N_14396);
and UO_1610 (O_1610,N_14817,N_14115);
or UO_1611 (O_1611,N_14884,N_14911);
or UO_1612 (O_1612,N_14731,N_14335);
nor UO_1613 (O_1613,N_14009,N_14491);
nor UO_1614 (O_1614,N_14596,N_14186);
or UO_1615 (O_1615,N_14316,N_14021);
nand UO_1616 (O_1616,N_14714,N_14230);
nor UO_1617 (O_1617,N_14429,N_14901);
or UO_1618 (O_1618,N_14748,N_14609);
or UO_1619 (O_1619,N_14144,N_14877);
and UO_1620 (O_1620,N_14077,N_14712);
nand UO_1621 (O_1621,N_14035,N_14353);
and UO_1622 (O_1622,N_14907,N_14459);
or UO_1623 (O_1623,N_14336,N_14000);
nor UO_1624 (O_1624,N_14379,N_14960);
nor UO_1625 (O_1625,N_14824,N_14123);
and UO_1626 (O_1626,N_14087,N_14492);
nand UO_1627 (O_1627,N_14879,N_14530);
or UO_1628 (O_1628,N_14047,N_14669);
or UO_1629 (O_1629,N_14202,N_14934);
nor UO_1630 (O_1630,N_14666,N_14037);
nand UO_1631 (O_1631,N_14754,N_14500);
nand UO_1632 (O_1632,N_14678,N_14797);
nor UO_1633 (O_1633,N_14008,N_14741);
or UO_1634 (O_1634,N_14296,N_14281);
or UO_1635 (O_1635,N_14869,N_14032);
nor UO_1636 (O_1636,N_14895,N_14121);
or UO_1637 (O_1637,N_14450,N_14623);
nor UO_1638 (O_1638,N_14047,N_14837);
and UO_1639 (O_1639,N_14219,N_14705);
nor UO_1640 (O_1640,N_14165,N_14414);
xnor UO_1641 (O_1641,N_14266,N_14357);
nand UO_1642 (O_1642,N_14837,N_14543);
nor UO_1643 (O_1643,N_14202,N_14870);
and UO_1644 (O_1644,N_14100,N_14982);
or UO_1645 (O_1645,N_14536,N_14160);
nand UO_1646 (O_1646,N_14621,N_14172);
nand UO_1647 (O_1647,N_14355,N_14907);
nor UO_1648 (O_1648,N_14288,N_14486);
nand UO_1649 (O_1649,N_14912,N_14119);
and UO_1650 (O_1650,N_14479,N_14093);
or UO_1651 (O_1651,N_14723,N_14266);
and UO_1652 (O_1652,N_14219,N_14772);
nand UO_1653 (O_1653,N_14401,N_14868);
and UO_1654 (O_1654,N_14027,N_14732);
and UO_1655 (O_1655,N_14554,N_14826);
or UO_1656 (O_1656,N_14086,N_14421);
nor UO_1657 (O_1657,N_14868,N_14538);
nand UO_1658 (O_1658,N_14097,N_14963);
and UO_1659 (O_1659,N_14104,N_14968);
xnor UO_1660 (O_1660,N_14875,N_14824);
or UO_1661 (O_1661,N_14476,N_14752);
or UO_1662 (O_1662,N_14570,N_14541);
and UO_1663 (O_1663,N_14895,N_14866);
or UO_1664 (O_1664,N_14658,N_14390);
and UO_1665 (O_1665,N_14418,N_14052);
nor UO_1666 (O_1666,N_14044,N_14201);
and UO_1667 (O_1667,N_14186,N_14883);
or UO_1668 (O_1668,N_14421,N_14445);
or UO_1669 (O_1669,N_14885,N_14866);
nand UO_1670 (O_1670,N_14719,N_14743);
nand UO_1671 (O_1671,N_14909,N_14407);
nor UO_1672 (O_1672,N_14335,N_14751);
and UO_1673 (O_1673,N_14081,N_14293);
nand UO_1674 (O_1674,N_14961,N_14916);
nand UO_1675 (O_1675,N_14233,N_14782);
and UO_1676 (O_1676,N_14715,N_14622);
and UO_1677 (O_1677,N_14679,N_14538);
and UO_1678 (O_1678,N_14692,N_14346);
or UO_1679 (O_1679,N_14021,N_14105);
nand UO_1680 (O_1680,N_14320,N_14991);
nor UO_1681 (O_1681,N_14292,N_14256);
nand UO_1682 (O_1682,N_14788,N_14570);
or UO_1683 (O_1683,N_14799,N_14707);
xor UO_1684 (O_1684,N_14668,N_14956);
nand UO_1685 (O_1685,N_14272,N_14804);
or UO_1686 (O_1686,N_14775,N_14363);
or UO_1687 (O_1687,N_14255,N_14254);
nor UO_1688 (O_1688,N_14137,N_14960);
or UO_1689 (O_1689,N_14367,N_14189);
xnor UO_1690 (O_1690,N_14780,N_14098);
nand UO_1691 (O_1691,N_14463,N_14228);
or UO_1692 (O_1692,N_14953,N_14555);
nand UO_1693 (O_1693,N_14940,N_14017);
nand UO_1694 (O_1694,N_14746,N_14055);
nor UO_1695 (O_1695,N_14404,N_14449);
or UO_1696 (O_1696,N_14134,N_14395);
nand UO_1697 (O_1697,N_14074,N_14470);
xnor UO_1698 (O_1698,N_14108,N_14614);
or UO_1699 (O_1699,N_14039,N_14532);
and UO_1700 (O_1700,N_14607,N_14452);
nor UO_1701 (O_1701,N_14196,N_14544);
and UO_1702 (O_1702,N_14881,N_14961);
and UO_1703 (O_1703,N_14036,N_14321);
nor UO_1704 (O_1704,N_14674,N_14481);
and UO_1705 (O_1705,N_14970,N_14164);
nor UO_1706 (O_1706,N_14865,N_14652);
and UO_1707 (O_1707,N_14852,N_14029);
or UO_1708 (O_1708,N_14851,N_14938);
and UO_1709 (O_1709,N_14464,N_14140);
nand UO_1710 (O_1710,N_14259,N_14805);
nand UO_1711 (O_1711,N_14804,N_14982);
nand UO_1712 (O_1712,N_14240,N_14050);
nor UO_1713 (O_1713,N_14473,N_14942);
or UO_1714 (O_1714,N_14796,N_14817);
nor UO_1715 (O_1715,N_14076,N_14276);
or UO_1716 (O_1716,N_14811,N_14082);
and UO_1717 (O_1717,N_14969,N_14048);
or UO_1718 (O_1718,N_14955,N_14450);
nor UO_1719 (O_1719,N_14433,N_14000);
or UO_1720 (O_1720,N_14698,N_14604);
and UO_1721 (O_1721,N_14154,N_14291);
nand UO_1722 (O_1722,N_14169,N_14385);
and UO_1723 (O_1723,N_14642,N_14546);
nand UO_1724 (O_1724,N_14033,N_14298);
nand UO_1725 (O_1725,N_14959,N_14883);
nor UO_1726 (O_1726,N_14886,N_14006);
nand UO_1727 (O_1727,N_14847,N_14947);
or UO_1728 (O_1728,N_14396,N_14492);
nand UO_1729 (O_1729,N_14990,N_14605);
or UO_1730 (O_1730,N_14351,N_14282);
nor UO_1731 (O_1731,N_14037,N_14201);
and UO_1732 (O_1732,N_14814,N_14969);
nand UO_1733 (O_1733,N_14307,N_14462);
or UO_1734 (O_1734,N_14531,N_14191);
xor UO_1735 (O_1735,N_14892,N_14961);
nand UO_1736 (O_1736,N_14570,N_14272);
nor UO_1737 (O_1737,N_14762,N_14291);
xor UO_1738 (O_1738,N_14411,N_14593);
and UO_1739 (O_1739,N_14882,N_14454);
and UO_1740 (O_1740,N_14773,N_14730);
or UO_1741 (O_1741,N_14643,N_14488);
xor UO_1742 (O_1742,N_14075,N_14370);
nor UO_1743 (O_1743,N_14579,N_14360);
nor UO_1744 (O_1744,N_14398,N_14898);
or UO_1745 (O_1745,N_14343,N_14073);
xor UO_1746 (O_1746,N_14948,N_14775);
nor UO_1747 (O_1747,N_14195,N_14801);
nor UO_1748 (O_1748,N_14163,N_14120);
nor UO_1749 (O_1749,N_14847,N_14784);
or UO_1750 (O_1750,N_14805,N_14171);
nand UO_1751 (O_1751,N_14204,N_14930);
nor UO_1752 (O_1752,N_14718,N_14579);
and UO_1753 (O_1753,N_14146,N_14477);
xor UO_1754 (O_1754,N_14578,N_14214);
xor UO_1755 (O_1755,N_14957,N_14774);
nor UO_1756 (O_1756,N_14390,N_14436);
nand UO_1757 (O_1757,N_14454,N_14180);
or UO_1758 (O_1758,N_14811,N_14699);
or UO_1759 (O_1759,N_14452,N_14002);
or UO_1760 (O_1760,N_14128,N_14881);
xnor UO_1761 (O_1761,N_14528,N_14374);
nand UO_1762 (O_1762,N_14964,N_14749);
nand UO_1763 (O_1763,N_14239,N_14058);
nand UO_1764 (O_1764,N_14621,N_14340);
nor UO_1765 (O_1765,N_14640,N_14917);
nor UO_1766 (O_1766,N_14193,N_14942);
nor UO_1767 (O_1767,N_14618,N_14794);
and UO_1768 (O_1768,N_14472,N_14735);
nor UO_1769 (O_1769,N_14089,N_14083);
nor UO_1770 (O_1770,N_14546,N_14563);
or UO_1771 (O_1771,N_14948,N_14262);
nand UO_1772 (O_1772,N_14602,N_14985);
nor UO_1773 (O_1773,N_14667,N_14698);
nor UO_1774 (O_1774,N_14404,N_14023);
or UO_1775 (O_1775,N_14654,N_14176);
and UO_1776 (O_1776,N_14741,N_14798);
nor UO_1777 (O_1777,N_14704,N_14970);
or UO_1778 (O_1778,N_14557,N_14180);
nor UO_1779 (O_1779,N_14715,N_14402);
or UO_1780 (O_1780,N_14136,N_14763);
or UO_1781 (O_1781,N_14094,N_14560);
nand UO_1782 (O_1782,N_14256,N_14891);
or UO_1783 (O_1783,N_14030,N_14945);
or UO_1784 (O_1784,N_14975,N_14740);
or UO_1785 (O_1785,N_14896,N_14080);
and UO_1786 (O_1786,N_14522,N_14200);
or UO_1787 (O_1787,N_14120,N_14219);
nor UO_1788 (O_1788,N_14272,N_14243);
nor UO_1789 (O_1789,N_14719,N_14944);
nor UO_1790 (O_1790,N_14649,N_14070);
and UO_1791 (O_1791,N_14069,N_14338);
nand UO_1792 (O_1792,N_14656,N_14222);
nor UO_1793 (O_1793,N_14651,N_14775);
nand UO_1794 (O_1794,N_14944,N_14034);
nor UO_1795 (O_1795,N_14728,N_14174);
nand UO_1796 (O_1796,N_14240,N_14350);
nor UO_1797 (O_1797,N_14128,N_14527);
nand UO_1798 (O_1798,N_14341,N_14529);
or UO_1799 (O_1799,N_14623,N_14014);
or UO_1800 (O_1800,N_14754,N_14538);
nor UO_1801 (O_1801,N_14750,N_14865);
xnor UO_1802 (O_1802,N_14193,N_14899);
and UO_1803 (O_1803,N_14272,N_14645);
and UO_1804 (O_1804,N_14894,N_14060);
or UO_1805 (O_1805,N_14166,N_14154);
or UO_1806 (O_1806,N_14393,N_14128);
or UO_1807 (O_1807,N_14784,N_14878);
nor UO_1808 (O_1808,N_14765,N_14064);
nor UO_1809 (O_1809,N_14548,N_14918);
nor UO_1810 (O_1810,N_14703,N_14491);
nor UO_1811 (O_1811,N_14022,N_14745);
nor UO_1812 (O_1812,N_14457,N_14189);
or UO_1813 (O_1813,N_14091,N_14102);
nor UO_1814 (O_1814,N_14382,N_14336);
nand UO_1815 (O_1815,N_14118,N_14847);
nor UO_1816 (O_1816,N_14162,N_14776);
and UO_1817 (O_1817,N_14960,N_14224);
nor UO_1818 (O_1818,N_14112,N_14488);
or UO_1819 (O_1819,N_14886,N_14329);
xor UO_1820 (O_1820,N_14206,N_14653);
or UO_1821 (O_1821,N_14952,N_14877);
or UO_1822 (O_1822,N_14288,N_14861);
or UO_1823 (O_1823,N_14230,N_14672);
nand UO_1824 (O_1824,N_14657,N_14250);
nand UO_1825 (O_1825,N_14756,N_14511);
or UO_1826 (O_1826,N_14596,N_14483);
nand UO_1827 (O_1827,N_14379,N_14147);
nand UO_1828 (O_1828,N_14459,N_14800);
and UO_1829 (O_1829,N_14665,N_14982);
nand UO_1830 (O_1830,N_14694,N_14324);
nand UO_1831 (O_1831,N_14684,N_14353);
nand UO_1832 (O_1832,N_14823,N_14794);
or UO_1833 (O_1833,N_14908,N_14542);
nand UO_1834 (O_1834,N_14305,N_14643);
or UO_1835 (O_1835,N_14016,N_14911);
and UO_1836 (O_1836,N_14941,N_14417);
and UO_1837 (O_1837,N_14876,N_14759);
or UO_1838 (O_1838,N_14940,N_14437);
nor UO_1839 (O_1839,N_14513,N_14795);
xnor UO_1840 (O_1840,N_14024,N_14850);
or UO_1841 (O_1841,N_14832,N_14137);
or UO_1842 (O_1842,N_14739,N_14639);
nand UO_1843 (O_1843,N_14748,N_14829);
and UO_1844 (O_1844,N_14728,N_14812);
nor UO_1845 (O_1845,N_14487,N_14103);
or UO_1846 (O_1846,N_14739,N_14726);
nand UO_1847 (O_1847,N_14795,N_14827);
nand UO_1848 (O_1848,N_14932,N_14400);
nand UO_1849 (O_1849,N_14661,N_14791);
nand UO_1850 (O_1850,N_14500,N_14441);
or UO_1851 (O_1851,N_14334,N_14888);
and UO_1852 (O_1852,N_14198,N_14618);
and UO_1853 (O_1853,N_14601,N_14480);
or UO_1854 (O_1854,N_14686,N_14558);
nand UO_1855 (O_1855,N_14664,N_14643);
or UO_1856 (O_1856,N_14375,N_14194);
xnor UO_1857 (O_1857,N_14299,N_14395);
or UO_1858 (O_1858,N_14153,N_14886);
nand UO_1859 (O_1859,N_14968,N_14622);
or UO_1860 (O_1860,N_14086,N_14419);
nand UO_1861 (O_1861,N_14859,N_14926);
xnor UO_1862 (O_1862,N_14210,N_14656);
or UO_1863 (O_1863,N_14627,N_14448);
nor UO_1864 (O_1864,N_14114,N_14722);
nand UO_1865 (O_1865,N_14162,N_14784);
nor UO_1866 (O_1866,N_14819,N_14336);
and UO_1867 (O_1867,N_14485,N_14968);
or UO_1868 (O_1868,N_14300,N_14541);
or UO_1869 (O_1869,N_14417,N_14584);
and UO_1870 (O_1870,N_14838,N_14438);
nor UO_1871 (O_1871,N_14676,N_14417);
or UO_1872 (O_1872,N_14127,N_14460);
nand UO_1873 (O_1873,N_14187,N_14254);
or UO_1874 (O_1874,N_14250,N_14897);
nor UO_1875 (O_1875,N_14417,N_14276);
and UO_1876 (O_1876,N_14938,N_14392);
nand UO_1877 (O_1877,N_14243,N_14749);
nor UO_1878 (O_1878,N_14434,N_14032);
nor UO_1879 (O_1879,N_14883,N_14298);
xor UO_1880 (O_1880,N_14165,N_14662);
and UO_1881 (O_1881,N_14101,N_14940);
nor UO_1882 (O_1882,N_14009,N_14499);
nand UO_1883 (O_1883,N_14410,N_14592);
nand UO_1884 (O_1884,N_14513,N_14284);
nand UO_1885 (O_1885,N_14223,N_14288);
and UO_1886 (O_1886,N_14211,N_14722);
nor UO_1887 (O_1887,N_14267,N_14247);
xor UO_1888 (O_1888,N_14995,N_14432);
nor UO_1889 (O_1889,N_14107,N_14105);
nand UO_1890 (O_1890,N_14075,N_14681);
nand UO_1891 (O_1891,N_14526,N_14447);
nor UO_1892 (O_1892,N_14740,N_14397);
nand UO_1893 (O_1893,N_14852,N_14699);
nor UO_1894 (O_1894,N_14536,N_14551);
nand UO_1895 (O_1895,N_14457,N_14690);
and UO_1896 (O_1896,N_14786,N_14638);
nor UO_1897 (O_1897,N_14602,N_14895);
or UO_1898 (O_1898,N_14012,N_14255);
and UO_1899 (O_1899,N_14730,N_14132);
nand UO_1900 (O_1900,N_14085,N_14617);
nor UO_1901 (O_1901,N_14107,N_14543);
xnor UO_1902 (O_1902,N_14044,N_14871);
and UO_1903 (O_1903,N_14643,N_14346);
and UO_1904 (O_1904,N_14036,N_14581);
nand UO_1905 (O_1905,N_14471,N_14664);
nand UO_1906 (O_1906,N_14400,N_14698);
and UO_1907 (O_1907,N_14428,N_14026);
and UO_1908 (O_1908,N_14358,N_14711);
nand UO_1909 (O_1909,N_14128,N_14110);
nand UO_1910 (O_1910,N_14871,N_14306);
or UO_1911 (O_1911,N_14713,N_14113);
nor UO_1912 (O_1912,N_14595,N_14009);
or UO_1913 (O_1913,N_14350,N_14080);
nand UO_1914 (O_1914,N_14832,N_14667);
nand UO_1915 (O_1915,N_14520,N_14877);
and UO_1916 (O_1916,N_14782,N_14290);
nand UO_1917 (O_1917,N_14525,N_14606);
and UO_1918 (O_1918,N_14690,N_14331);
or UO_1919 (O_1919,N_14902,N_14201);
and UO_1920 (O_1920,N_14920,N_14669);
and UO_1921 (O_1921,N_14206,N_14450);
or UO_1922 (O_1922,N_14795,N_14477);
or UO_1923 (O_1923,N_14938,N_14148);
nand UO_1924 (O_1924,N_14527,N_14772);
and UO_1925 (O_1925,N_14941,N_14565);
nand UO_1926 (O_1926,N_14765,N_14364);
nor UO_1927 (O_1927,N_14678,N_14871);
or UO_1928 (O_1928,N_14871,N_14128);
or UO_1929 (O_1929,N_14050,N_14867);
or UO_1930 (O_1930,N_14608,N_14619);
nor UO_1931 (O_1931,N_14371,N_14013);
or UO_1932 (O_1932,N_14589,N_14724);
and UO_1933 (O_1933,N_14367,N_14898);
nor UO_1934 (O_1934,N_14500,N_14949);
nor UO_1935 (O_1935,N_14436,N_14467);
nand UO_1936 (O_1936,N_14236,N_14178);
and UO_1937 (O_1937,N_14447,N_14399);
xor UO_1938 (O_1938,N_14341,N_14536);
or UO_1939 (O_1939,N_14927,N_14339);
or UO_1940 (O_1940,N_14235,N_14181);
and UO_1941 (O_1941,N_14332,N_14082);
xor UO_1942 (O_1942,N_14984,N_14321);
or UO_1943 (O_1943,N_14154,N_14764);
nand UO_1944 (O_1944,N_14036,N_14833);
or UO_1945 (O_1945,N_14060,N_14141);
nor UO_1946 (O_1946,N_14675,N_14863);
and UO_1947 (O_1947,N_14759,N_14290);
nand UO_1948 (O_1948,N_14033,N_14335);
nand UO_1949 (O_1949,N_14159,N_14319);
nor UO_1950 (O_1950,N_14934,N_14584);
nor UO_1951 (O_1951,N_14298,N_14058);
nor UO_1952 (O_1952,N_14793,N_14328);
xnor UO_1953 (O_1953,N_14352,N_14604);
nand UO_1954 (O_1954,N_14176,N_14297);
nand UO_1955 (O_1955,N_14518,N_14246);
xor UO_1956 (O_1956,N_14317,N_14700);
nor UO_1957 (O_1957,N_14936,N_14314);
nand UO_1958 (O_1958,N_14746,N_14218);
nand UO_1959 (O_1959,N_14171,N_14470);
or UO_1960 (O_1960,N_14685,N_14052);
xnor UO_1961 (O_1961,N_14651,N_14917);
and UO_1962 (O_1962,N_14552,N_14203);
and UO_1963 (O_1963,N_14406,N_14692);
nand UO_1964 (O_1964,N_14328,N_14724);
or UO_1965 (O_1965,N_14661,N_14753);
or UO_1966 (O_1966,N_14187,N_14506);
or UO_1967 (O_1967,N_14513,N_14868);
or UO_1968 (O_1968,N_14182,N_14401);
nor UO_1969 (O_1969,N_14792,N_14114);
and UO_1970 (O_1970,N_14297,N_14037);
and UO_1971 (O_1971,N_14016,N_14084);
and UO_1972 (O_1972,N_14694,N_14274);
nor UO_1973 (O_1973,N_14056,N_14675);
or UO_1974 (O_1974,N_14623,N_14469);
or UO_1975 (O_1975,N_14298,N_14084);
xnor UO_1976 (O_1976,N_14820,N_14190);
xor UO_1977 (O_1977,N_14041,N_14660);
or UO_1978 (O_1978,N_14335,N_14225);
nand UO_1979 (O_1979,N_14260,N_14632);
nand UO_1980 (O_1980,N_14893,N_14903);
or UO_1981 (O_1981,N_14060,N_14602);
nand UO_1982 (O_1982,N_14221,N_14921);
xor UO_1983 (O_1983,N_14811,N_14761);
nor UO_1984 (O_1984,N_14487,N_14560);
nand UO_1985 (O_1985,N_14902,N_14364);
nor UO_1986 (O_1986,N_14175,N_14716);
nor UO_1987 (O_1987,N_14979,N_14088);
xnor UO_1988 (O_1988,N_14656,N_14268);
xor UO_1989 (O_1989,N_14419,N_14974);
or UO_1990 (O_1990,N_14287,N_14364);
nor UO_1991 (O_1991,N_14290,N_14941);
and UO_1992 (O_1992,N_14633,N_14415);
or UO_1993 (O_1993,N_14205,N_14590);
nand UO_1994 (O_1994,N_14336,N_14503);
nand UO_1995 (O_1995,N_14292,N_14305);
nand UO_1996 (O_1996,N_14163,N_14365);
xor UO_1997 (O_1997,N_14149,N_14514);
nor UO_1998 (O_1998,N_14728,N_14744);
or UO_1999 (O_1999,N_14819,N_14937);
endmodule