module basic_1000_10000_1500_2_levels_1xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5003,N_5004,N_5005,N_5006,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5017,N_5018,N_5022,N_5023,N_5026,N_5027,N_5029,N_5030,N_5032,N_5033,N_5035,N_5036,N_5037,N_5039,N_5041,N_5044,N_5046,N_5049,N_5051,N_5052,N_5055,N_5056,N_5058,N_5059,N_5062,N_5063,N_5064,N_5068,N_5069,N_5072,N_5073,N_5074,N_5076,N_5078,N_5080,N_5085,N_5086,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5099,N_5101,N_5102,N_5103,N_5104,N_5108,N_5109,N_5110,N_5113,N_5115,N_5116,N_5117,N_5118,N_5119,N_5121,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5142,N_5145,N_5149,N_5151,N_5152,N_5153,N_5155,N_5156,N_5158,N_5159,N_5160,N_5161,N_5163,N_5165,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5177,N_5182,N_5183,N_5186,N_5189,N_5190,N_5191,N_5193,N_5194,N_5195,N_5200,N_5202,N_5207,N_5209,N_5210,N_5211,N_5218,N_5219,N_5224,N_5225,N_5227,N_5228,N_5229,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5241,N_5243,N_5245,N_5247,N_5248,N_5249,N_5252,N_5253,N_5254,N_5255,N_5259,N_5261,N_5262,N_5266,N_5267,N_5268,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5289,N_5293,N_5295,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5304,N_5308,N_5310,N_5311,N_5312,N_5313,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5337,N_5338,N_5344,N_5348,N_5349,N_5350,N_5352,N_5354,N_5355,N_5356,N_5358,N_5359,N_5360,N_5361,N_5362,N_5364,N_5366,N_5367,N_5368,N_5369,N_5373,N_5374,N_5376,N_5377,N_5378,N_5379,N_5380,N_5384,N_5385,N_5386,N_5387,N_5389,N_5393,N_5396,N_5399,N_5400,N_5401,N_5402,N_5403,N_5406,N_5408,N_5410,N_5411,N_5412,N_5413,N_5417,N_5420,N_5422,N_5423,N_5424,N_5426,N_5427,N_5428,N_5433,N_5435,N_5437,N_5441,N_5442,N_5443,N_5445,N_5447,N_5448,N_5449,N_5450,N_5452,N_5453,N_5456,N_5460,N_5462,N_5463,N_5464,N_5467,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5484,N_5485,N_5488,N_5489,N_5491,N_5492,N_5494,N_5497,N_5499,N_5500,N_5501,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5511,N_5513,N_5514,N_5515,N_5516,N_5519,N_5520,N_5521,N_5522,N_5523,N_5525,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5536,N_5537,N_5539,N_5540,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5551,N_5553,N_5556,N_5558,N_5559,N_5560,N_5562,N_5563,N_5564,N_5565,N_5568,N_5569,N_5571,N_5572,N_5573,N_5576,N_5578,N_5579,N_5580,N_5583,N_5585,N_5586,N_5588,N_5589,N_5591,N_5593,N_5597,N_5599,N_5600,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5610,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5619,N_5620,N_5621,N_5622,N_5623,N_5625,N_5626,N_5627,N_5630,N_5634,N_5636,N_5637,N_5638,N_5640,N_5642,N_5643,N_5645,N_5646,N_5647,N_5648,N_5650,N_5653,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5680,N_5682,N_5683,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5695,N_5696,N_5697,N_5699,N_5700,N_5701,N_5702,N_5705,N_5706,N_5707,N_5710,N_5712,N_5713,N_5714,N_5715,N_5716,N_5720,N_5722,N_5723,N_5724,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5733,N_5734,N_5735,N_5737,N_5738,N_5739,N_5741,N_5742,N_5743,N_5746,N_5749,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5765,N_5768,N_5770,N_5772,N_5775,N_5776,N_5777,N_5779,N_5780,N_5781,N_5785,N_5786,N_5787,N_5788,N_5791,N_5795,N_5796,N_5799,N_5801,N_5802,N_5803,N_5805,N_5806,N_5807,N_5810,N_5812,N_5814,N_5815,N_5817,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5838,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5855,N_5857,N_5859,N_5860,N_5861,N_5862,N_5863,N_5867,N_5871,N_5872,N_5874,N_5875,N_5877,N_5879,N_5880,N_5881,N_5884,N_5888,N_5891,N_5894,N_5897,N_5899,N_5903,N_5904,N_5905,N_5906,N_5908,N_5909,N_5910,N_5911,N_5913,N_5914,N_5916,N_5918,N_5919,N_5920,N_5921,N_5922,N_5924,N_5926,N_5929,N_5930,N_5932,N_5933,N_5934,N_5935,N_5936,N_5938,N_5939,N_5942,N_5945,N_5946,N_5947,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5956,N_5957,N_5962,N_5963,N_5965,N_5968,N_5969,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5982,N_5984,N_5986,N_5987,N_5990,N_5991,N_5992,N_5993,N_5996,N_5998,N_5999,N_6000,N_6001,N_6002,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6013,N_6016,N_6017,N_6019,N_6020,N_6021,N_6022,N_6023,N_6026,N_6027,N_6028,N_6029,N_6031,N_6032,N_6033,N_6034,N_6036,N_6037,N_6040,N_6041,N_6043,N_6044,N_6049,N_6050,N_6053,N_6054,N_6055,N_6057,N_6060,N_6062,N_6068,N_6071,N_6075,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6087,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6101,N_6103,N_6104,N_6105,N_6108,N_6109,N_6110,N_6113,N_6114,N_6116,N_6120,N_6122,N_6123,N_6124,N_6125,N_6129,N_6130,N_6132,N_6133,N_6135,N_6137,N_6138,N_6139,N_6141,N_6142,N_6143,N_6144,N_6147,N_6148,N_6149,N_6150,N_6151,N_6153,N_6154,N_6155,N_6158,N_6159,N_6160,N_6161,N_6162,N_6164,N_6165,N_6166,N_6168,N_6171,N_6172,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6183,N_6184,N_6185,N_6186,N_6188,N_6189,N_6190,N_6192,N_6194,N_6195,N_6197,N_6198,N_6200,N_6202,N_6203,N_6204,N_6206,N_6207,N_6208,N_6209,N_6212,N_6213,N_6215,N_6218,N_6219,N_6220,N_6221,N_6222,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6238,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6248,N_6252,N_6254,N_6255,N_6256,N_6259,N_6260,N_6262,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6283,N_6284,N_6286,N_6287,N_6288,N_6292,N_6293,N_6294,N_6297,N_6299,N_6303,N_6307,N_6311,N_6312,N_6315,N_6317,N_6318,N_6320,N_6322,N_6323,N_6326,N_6327,N_6328,N_6329,N_6330,N_6332,N_6333,N_6334,N_6335,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6345,N_6347,N_6348,N_6349,N_6351,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6364,N_6365,N_6367,N_6368,N_6370,N_6371,N_6374,N_6379,N_6380,N_6381,N_6382,N_6383,N_6385,N_6387,N_6391,N_6393,N_6395,N_6396,N_6400,N_6401,N_6404,N_6407,N_6408,N_6409,N_6411,N_6412,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6434,N_6435,N_6437,N_6438,N_6441,N_6443,N_6444,N_6445,N_6446,N_6447,N_6450,N_6451,N_6454,N_6456,N_6458,N_6459,N_6460,N_6461,N_6464,N_6465,N_6466,N_6467,N_6468,N_6471,N_6475,N_6476,N_6477,N_6479,N_6481,N_6482,N_6484,N_6486,N_6487,N_6489,N_6490,N_6491,N_6492,N_6494,N_6497,N_6500,N_6502,N_6503,N_6505,N_6506,N_6509,N_6510,N_6513,N_6515,N_6517,N_6520,N_6523,N_6526,N_6527,N_6528,N_6530,N_6531,N_6533,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6543,N_6544,N_6545,N_6549,N_6550,N_6552,N_6554,N_6555,N_6557,N_6559,N_6561,N_6562,N_6564,N_6565,N_6569,N_6570,N_6572,N_6573,N_6575,N_6579,N_6580,N_6581,N_6582,N_6583,N_6585,N_6586,N_6588,N_6590,N_6591,N_6592,N_6595,N_6596,N_6598,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6610,N_6612,N_6614,N_6615,N_6617,N_6619,N_6620,N_6621,N_6622,N_6624,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6638,N_6640,N_6642,N_6644,N_6645,N_6646,N_6649,N_6650,N_6653,N_6654,N_6657,N_6658,N_6659,N_6661,N_6664,N_6666,N_6667,N_6668,N_6670,N_6671,N_6673,N_6674,N_6675,N_6677,N_6678,N_6683,N_6684,N_6685,N_6688,N_6690,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6707,N_6710,N_6711,N_6712,N_6714,N_6716,N_6717,N_6718,N_6719,N_6720,N_6722,N_6723,N_6725,N_6726,N_6727,N_6729,N_6730,N_6734,N_6735,N_6736,N_6737,N_6739,N_6740,N_6747,N_6749,N_6752,N_6754,N_6756,N_6758,N_6761,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6771,N_6774,N_6778,N_6781,N_6783,N_6786,N_6787,N_6790,N_6792,N_6793,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6808,N_6810,N_6811,N_6813,N_6817,N_6818,N_6820,N_6821,N_6822,N_6824,N_6826,N_6827,N_6828,N_6831,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6842,N_6843,N_6844,N_6848,N_6849,N_6850,N_6851,N_6854,N_6856,N_6857,N_6859,N_6862,N_6864,N_6867,N_6868,N_6870,N_6871,N_6874,N_6876,N_6877,N_6878,N_6880,N_6882,N_6884,N_6885,N_6886,N_6889,N_6891,N_6892,N_6893,N_6895,N_6899,N_6900,N_6901,N_6902,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6913,N_6914,N_6915,N_6916,N_6917,N_6919,N_6920,N_6921,N_6923,N_6924,N_6925,N_6926,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6938,N_6939,N_6940,N_6943,N_6944,N_6945,N_6949,N_6950,N_6953,N_6955,N_6960,N_6961,N_6962,N_6963,N_6964,N_6966,N_6967,N_6968,N_6969,N_6971,N_6972,N_6974,N_6977,N_6978,N_6979,N_6981,N_6983,N_6986,N_6988,N_6989,N_6991,N_6992,N_6995,N_6998,N_7000,N_7001,N_7003,N_7004,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7014,N_7015,N_7016,N_7018,N_7019,N_7020,N_7022,N_7025,N_7027,N_7028,N_7029,N_7031,N_7032,N_7033,N_7037,N_7038,N_7039,N_7041,N_7045,N_7046,N_7048,N_7049,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7060,N_7061,N_7062,N_7064,N_7066,N_7067,N_7068,N_7070,N_7072,N_7073,N_7075,N_7078,N_7079,N_7080,N_7085,N_7086,N_7088,N_7089,N_7090,N_7093,N_7095,N_7096,N_7097,N_7098,N_7099,N_7101,N_7103,N_7105,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7120,N_7121,N_7122,N_7125,N_7126,N_7128,N_7129,N_7130,N_7131,N_7133,N_7134,N_7137,N_7138,N_7140,N_7141,N_7142,N_7143,N_7145,N_7150,N_7151,N_7152,N_7155,N_7157,N_7158,N_7159,N_7160,N_7161,N_7165,N_7166,N_7169,N_7171,N_7172,N_7173,N_7176,N_7178,N_7179,N_7181,N_7184,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7194,N_7199,N_7200,N_7205,N_7206,N_7208,N_7211,N_7212,N_7213,N_7215,N_7217,N_7218,N_7219,N_7220,N_7222,N_7224,N_7225,N_7226,N_7227,N_7229,N_7230,N_7232,N_7233,N_7234,N_7235,N_7238,N_7239,N_7240,N_7241,N_7242,N_7246,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7257,N_7258,N_7259,N_7260,N_7261,N_7265,N_7267,N_7270,N_7271,N_7275,N_7278,N_7279,N_7281,N_7282,N_7283,N_7284,N_7285,N_7288,N_7290,N_7291,N_7292,N_7294,N_7297,N_7300,N_7301,N_7303,N_7304,N_7307,N_7308,N_7309,N_7311,N_7312,N_7313,N_7318,N_7319,N_7320,N_7321,N_7323,N_7324,N_7325,N_7328,N_7330,N_7332,N_7333,N_7334,N_7336,N_7337,N_7339,N_7341,N_7342,N_7343,N_7345,N_7346,N_7347,N_7348,N_7349,N_7351,N_7352,N_7353,N_7355,N_7356,N_7358,N_7359,N_7360,N_7361,N_7362,N_7364,N_7365,N_7368,N_7370,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7383,N_7385,N_7387,N_7388,N_7389,N_7391,N_7392,N_7393,N_7394,N_7397,N_7398,N_7400,N_7401,N_7402,N_7403,N_7405,N_7406,N_7407,N_7408,N_7410,N_7411,N_7413,N_7416,N_7417,N_7422,N_7423,N_7424,N_7427,N_7428,N_7429,N_7431,N_7432,N_7433,N_7435,N_7437,N_7442,N_7445,N_7446,N_7447,N_7448,N_7451,N_7452,N_7453,N_7454,N_7456,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7467,N_7470,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7479,N_7480,N_7482,N_7486,N_7487,N_7489,N_7492,N_7495,N_7496,N_7498,N_7500,N_7501,N_7503,N_7504,N_7505,N_7506,N_7509,N_7511,N_7514,N_7515,N_7519,N_7521,N_7522,N_7523,N_7526,N_7527,N_7528,N_7529,N_7530,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7546,N_7548,N_7550,N_7552,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7562,N_7563,N_7566,N_7567,N_7568,N_7571,N_7573,N_7574,N_7576,N_7578,N_7579,N_7581,N_7583,N_7584,N_7586,N_7587,N_7588,N_7589,N_7590,N_7593,N_7595,N_7597,N_7598,N_7600,N_7601,N_7602,N_7603,N_7605,N_7608,N_7609,N_7610,N_7611,N_7614,N_7618,N_7624,N_7625,N_7626,N_7627,N_7629,N_7630,N_7631,N_7634,N_7635,N_7638,N_7640,N_7641,N_7642,N_7644,N_7647,N_7648,N_7650,N_7651,N_7653,N_7656,N_7657,N_7659,N_7660,N_7661,N_7662,N_7666,N_7668,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7678,N_7679,N_7680,N_7681,N_7682,N_7684,N_7686,N_7687,N_7688,N_7690,N_7691,N_7692,N_7693,N_7695,N_7696,N_7697,N_7698,N_7701,N_7702,N_7705,N_7706,N_7709,N_7710,N_7712,N_7713,N_7716,N_7717,N_7719,N_7720,N_7721,N_7726,N_7728,N_7729,N_7730,N_7733,N_7736,N_7737,N_7738,N_7743,N_7744,N_7745,N_7746,N_7748,N_7750,N_7754,N_7756,N_7758,N_7760,N_7761,N_7762,N_7763,N_7764,N_7767,N_7768,N_7769,N_7771,N_7772,N_7774,N_7776,N_7777,N_7780,N_7781,N_7782,N_7784,N_7785,N_7786,N_7787,N_7791,N_7792,N_7793,N_7794,N_7799,N_7800,N_7803,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7813,N_7814,N_7816,N_7817,N_7819,N_7823,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7839,N_7842,N_7844,N_7845,N_7846,N_7850,N_7851,N_7852,N_7853,N_7854,N_7857,N_7859,N_7860,N_7861,N_7862,N_7865,N_7867,N_7869,N_7870,N_7872,N_7874,N_7875,N_7876,N_7879,N_7882,N_7883,N_7884,N_7888,N_7891,N_7893,N_7894,N_7895,N_7896,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7905,N_7906,N_7907,N_7910,N_7911,N_7912,N_7914,N_7919,N_7920,N_7922,N_7923,N_7924,N_7926,N_7927,N_7929,N_7930,N_7933,N_7934,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7945,N_7947,N_7950,N_7951,N_7953,N_7954,N_7955,N_7957,N_7959,N_7960,N_7967,N_7970,N_7973,N_7974,N_7976,N_7979,N_7980,N_7981,N_7982,N_7983,N_7986,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8003,N_8004,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8021,N_8023,N_8024,N_8027,N_8029,N_8030,N_8032,N_8034,N_8035,N_8036,N_8038,N_8039,N_8041,N_8042,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8067,N_8068,N_8069,N_8072,N_8073,N_8076,N_8077,N_8078,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8101,N_8102,N_8103,N_8104,N_8105,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8114,N_8116,N_8117,N_8118,N_8119,N_8122,N_8123,N_8125,N_8127,N_8128,N_8130,N_8134,N_8135,N_8136,N_8137,N_8138,N_8140,N_8146,N_8148,N_8149,N_8151,N_8152,N_8153,N_8154,N_8156,N_8157,N_8158,N_8159,N_8161,N_8162,N_8163,N_8164,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8179,N_8180,N_8181,N_8182,N_8184,N_8186,N_8187,N_8189,N_8190,N_8192,N_8194,N_8195,N_8196,N_8200,N_8202,N_8204,N_8206,N_8207,N_8209,N_8210,N_8211,N_8213,N_8215,N_8216,N_8220,N_8221,N_8226,N_8227,N_8229,N_8230,N_8233,N_8235,N_8236,N_8240,N_8241,N_8242,N_8243,N_8244,N_8248,N_8249,N_8251,N_8252,N_8254,N_8255,N_8258,N_8259,N_8260,N_8261,N_8263,N_8266,N_8267,N_8268,N_8271,N_8272,N_8274,N_8276,N_8277,N_8278,N_8279,N_8283,N_8284,N_8285,N_8286,N_8288,N_8289,N_8291,N_8292,N_8293,N_8294,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8304,N_8305,N_8307,N_8310,N_8313,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8325,N_8326,N_8328,N_8329,N_8334,N_8335,N_8336,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8345,N_8347,N_8348,N_8349,N_8350,N_8351,N_8353,N_8355,N_8356,N_8359,N_8360,N_8361,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8374,N_8375,N_8376,N_8377,N_8379,N_8380,N_8383,N_8386,N_8388,N_8389,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8401,N_8402,N_8403,N_8409,N_8410,N_8411,N_8415,N_8419,N_8420,N_8421,N_8422,N_8423,N_8426,N_8428,N_8432,N_8435,N_8436,N_8437,N_8438,N_8439,N_8441,N_8442,N_8443,N_8445,N_8446,N_8447,N_8450,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8461,N_8462,N_8463,N_8464,N_8466,N_8468,N_8469,N_8471,N_8472,N_8474,N_8477,N_8478,N_8479,N_8481,N_8482,N_8483,N_8486,N_8488,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8502,N_8503,N_8507,N_8508,N_8510,N_8514,N_8515,N_8516,N_8519,N_8520,N_8526,N_8528,N_8531,N_8532,N_8534,N_8536,N_8537,N_8538,N_8542,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8555,N_8556,N_8558,N_8560,N_8561,N_8563,N_8564,N_8566,N_8567,N_8569,N_8570,N_8571,N_8573,N_8575,N_8576,N_8577,N_8579,N_8580,N_8581,N_8582,N_8583,N_8585,N_8586,N_8589,N_8592,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8609,N_8610,N_8611,N_8612,N_8613,N_8620,N_8623,N_8626,N_8627,N_8629,N_8632,N_8633,N_8634,N_8636,N_8637,N_8639,N_8640,N_8642,N_8649,N_8650,N_8652,N_8653,N_8655,N_8656,N_8657,N_8661,N_8662,N_8663,N_8665,N_8666,N_8669,N_8670,N_8671,N_8672,N_8674,N_8675,N_8676,N_8678,N_8681,N_8682,N_8685,N_8686,N_8687,N_8688,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8698,N_8700,N_8701,N_8702,N_8704,N_8707,N_8711,N_8715,N_8716,N_8718,N_8719,N_8720,N_8721,N_8725,N_8726,N_8728,N_8729,N_8730,N_8731,N_8733,N_8738,N_8740,N_8743,N_8745,N_8747,N_8750,N_8751,N_8754,N_8756,N_8759,N_8760,N_8761,N_8763,N_8765,N_8767,N_8770,N_8771,N_8773,N_8774,N_8778,N_8779,N_8780,N_8781,N_8783,N_8785,N_8786,N_8787,N_8788,N_8789,N_8791,N_8792,N_8795,N_8797,N_8799,N_8800,N_8801,N_8802,N_8803,N_8805,N_8806,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8823,N_8826,N_8827,N_8830,N_8834,N_8835,N_8836,N_8840,N_8842,N_8844,N_8845,N_8847,N_8848,N_8849,N_8850,N_8851,N_8853,N_8855,N_8856,N_8857,N_8858,N_8859,N_8862,N_8864,N_8866,N_8867,N_8868,N_8870,N_8871,N_8872,N_8873,N_8876,N_8878,N_8881,N_8882,N_8885,N_8887,N_8892,N_8894,N_8897,N_8899,N_8900,N_8902,N_8904,N_8906,N_8909,N_8910,N_8911,N_8912,N_8914,N_8915,N_8917,N_8918,N_8924,N_8925,N_8926,N_8928,N_8929,N_8930,N_8931,N_8934,N_8937,N_8939,N_8940,N_8946,N_8947,N_8948,N_8952,N_8953,N_8955,N_8956,N_8957,N_8959,N_8960,N_8961,N_8965,N_8966,N_8967,N_8968,N_8972,N_8973,N_8976,N_8977,N_8978,N_8980,N_8981,N_8982,N_8985,N_8986,N_8987,N_8989,N_8990,N_8991,N_8992,N_8993,N_8996,N_8997,N_8998,N_9001,N_9002,N_9003,N_9004,N_9006,N_9008,N_9009,N_9010,N_9011,N_9013,N_9015,N_9016,N_9017,N_9018,N_9019,N_9022,N_9024,N_9025,N_9027,N_9028,N_9030,N_9031,N_9033,N_9034,N_9036,N_9037,N_9038,N_9041,N_9043,N_9047,N_9048,N_9049,N_9050,N_9051,N_9053,N_9054,N_9055,N_9056,N_9058,N_9059,N_9060,N_9061,N_9062,N_9064,N_9065,N_9066,N_9067,N_9070,N_9071,N_9073,N_9074,N_9075,N_9077,N_9078,N_9079,N_9081,N_9084,N_9085,N_9086,N_9087,N_9089,N_9090,N_9092,N_9093,N_9099,N_9101,N_9104,N_9105,N_9106,N_9108,N_9109,N_9110,N_9112,N_9116,N_9117,N_9118,N_9121,N_9122,N_9123,N_9125,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9138,N_9141,N_9142,N_9143,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9152,N_9155,N_9157,N_9158,N_9159,N_9162,N_9168,N_9169,N_9170,N_9171,N_9174,N_9178,N_9183,N_9186,N_9189,N_9190,N_9193,N_9196,N_9197,N_9204,N_9208,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9230,N_9232,N_9237,N_9238,N_9241,N_9242,N_9245,N_9247,N_9248,N_9251,N_9253,N_9254,N_9256,N_9261,N_9263,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9275,N_9276,N_9277,N_9279,N_9282,N_9283,N_9284,N_9285,N_9286,N_9288,N_9289,N_9290,N_9293,N_9294,N_9295,N_9297,N_9298,N_9299,N_9301,N_9302,N_9303,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9314,N_9315,N_9318,N_9319,N_9321,N_9322,N_9324,N_9325,N_9327,N_9328,N_9330,N_9331,N_9336,N_9337,N_9338,N_9340,N_9342,N_9343,N_9347,N_9348,N_9350,N_9352,N_9353,N_9354,N_9356,N_9360,N_9362,N_9363,N_9365,N_9366,N_9367,N_9368,N_9370,N_9374,N_9375,N_9376,N_9379,N_9380,N_9381,N_9382,N_9384,N_9387,N_9388,N_9389,N_9390,N_9393,N_9396,N_9400,N_9401,N_9403,N_9404,N_9405,N_9406,N_9407,N_9409,N_9411,N_9412,N_9414,N_9415,N_9416,N_9417,N_9418,N_9421,N_9423,N_9425,N_9427,N_9429,N_9435,N_9437,N_9438,N_9439,N_9441,N_9443,N_9444,N_9445,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9454,N_9456,N_9459,N_9460,N_9461,N_9464,N_9467,N_9468,N_9470,N_9472,N_9474,N_9475,N_9476,N_9477,N_9479,N_9480,N_9481,N_9483,N_9485,N_9486,N_9487,N_9489,N_9492,N_9493,N_9494,N_9496,N_9497,N_9500,N_9506,N_9507,N_9512,N_9513,N_9515,N_9516,N_9519,N_9521,N_9525,N_9527,N_9528,N_9530,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9541,N_9544,N_9545,N_9546,N_9547,N_9549,N_9551,N_9552,N_9553,N_9554,N_9555,N_9558,N_9564,N_9566,N_9568,N_9571,N_9574,N_9575,N_9578,N_9579,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9590,N_9591,N_9592,N_9596,N_9597,N_9599,N_9600,N_9603,N_9605,N_9606,N_9607,N_9608,N_9610,N_9611,N_9612,N_9613,N_9614,N_9617,N_9618,N_9620,N_9621,N_9623,N_9625,N_9626,N_9627,N_9630,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9651,N_9653,N_9655,N_9657,N_9658,N_9659,N_9661,N_9666,N_9669,N_9670,N_9671,N_9672,N_9673,N_9677,N_9679,N_9680,N_9681,N_9682,N_9683,N_9686,N_9687,N_9690,N_9691,N_9695,N_9696,N_9697,N_9699,N_9700,N_9703,N_9704,N_9705,N_9706,N_9708,N_9710,N_9711,N_9713,N_9715,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9729,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9757,N_9759,N_9761,N_9762,N_9763,N_9765,N_9766,N_9767,N_9770,N_9771,N_9772,N_9773,N_9774,N_9777,N_9778,N_9783,N_9784,N_9787,N_9788,N_9789,N_9790,N_9792,N_9793,N_9794,N_9795,N_9796,N_9799,N_9800,N_9803,N_9805,N_9807,N_9809,N_9810,N_9813,N_9814,N_9816,N_9818,N_9820,N_9821,N_9823,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9836,N_9839,N_9842,N_9843,N_9844,N_9845,N_9846,N_9854,N_9855,N_9856,N_9858,N_9859,N_9860,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9873,N_9876,N_9878,N_9879,N_9880,N_9882,N_9884,N_9886,N_9887,N_9893,N_9894,N_9895,N_9896,N_9899,N_9900,N_9902,N_9903,N_9908,N_9910,N_9911,N_9914,N_9915,N_9917,N_9918,N_9920,N_9928,N_9930,N_9934,N_9936,N_9937,N_9938,N_9939,N_9940,N_9943,N_9944,N_9945,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9964,N_9965,N_9968,N_9969,N_9976,N_9977,N_9978,N_9979,N_9981,N_9984,N_9986,N_9988,N_9992,N_9996,N_9999;
or U0 (N_0,In_502,In_257);
nor U1 (N_1,In_61,In_735);
nand U2 (N_2,In_270,In_599);
nand U3 (N_3,In_408,In_225);
nor U4 (N_4,In_439,In_963);
nor U5 (N_5,In_271,In_54);
nor U6 (N_6,In_552,In_495);
or U7 (N_7,In_337,In_978);
and U8 (N_8,In_340,In_618);
and U9 (N_9,In_78,In_349);
nor U10 (N_10,In_508,In_258);
or U11 (N_11,In_249,In_716);
and U12 (N_12,In_260,In_747);
nand U13 (N_13,In_646,In_840);
nand U14 (N_14,In_804,In_566);
and U15 (N_15,In_455,In_917);
nor U16 (N_16,In_347,In_129);
or U17 (N_17,In_720,In_724);
or U18 (N_18,In_119,In_703);
or U19 (N_19,In_571,In_158);
nand U20 (N_20,In_490,In_313);
nand U21 (N_21,In_3,In_197);
nand U22 (N_22,In_932,In_544);
and U23 (N_23,In_302,In_244);
or U24 (N_24,In_76,In_996);
and U25 (N_25,In_280,In_708);
nor U26 (N_26,In_900,In_780);
nor U27 (N_27,In_564,In_940);
or U28 (N_28,In_562,In_391);
or U29 (N_29,In_558,In_984);
and U30 (N_30,In_626,In_224);
nand U31 (N_31,In_176,In_367);
or U32 (N_32,In_550,In_142);
or U33 (N_33,In_605,In_8);
nand U34 (N_34,In_885,In_489);
nand U35 (N_35,In_476,In_306);
nor U36 (N_36,In_382,In_120);
or U37 (N_37,In_348,In_103);
nand U38 (N_38,In_240,In_210);
or U39 (N_39,In_288,In_737);
nor U40 (N_40,In_925,In_739);
and U41 (N_41,In_662,In_557);
nor U42 (N_42,In_146,In_664);
nand U43 (N_43,In_933,In_354);
and U44 (N_44,In_203,In_725);
and U45 (N_45,In_853,In_310);
nand U46 (N_46,In_364,In_635);
nor U47 (N_47,In_561,In_111);
nor U48 (N_48,In_128,In_897);
and U49 (N_49,In_682,In_384);
and U50 (N_50,In_190,In_356);
nand U51 (N_51,In_184,In_761);
nor U52 (N_52,In_623,In_164);
and U53 (N_53,In_469,In_463);
and U54 (N_54,In_654,In_785);
or U55 (N_55,In_15,In_899);
and U56 (N_56,In_707,In_715);
and U57 (N_57,In_729,In_631);
and U58 (N_58,In_868,In_907);
or U59 (N_59,In_771,In_393);
or U60 (N_60,In_808,In_714);
nand U61 (N_61,In_882,In_377);
and U62 (N_62,In_753,In_437);
and U63 (N_63,In_549,In_903);
nor U64 (N_64,In_48,In_829);
or U65 (N_65,In_308,In_777);
nand U66 (N_66,In_740,In_207);
nand U67 (N_67,In_28,In_137);
nor U68 (N_68,In_718,In_997);
nand U69 (N_69,In_500,In_236);
and U70 (N_70,In_583,In_171);
and U71 (N_71,In_669,In_973);
or U72 (N_72,In_417,In_923);
and U73 (N_73,In_191,In_212);
and U74 (N_74,In_974,In_162);
or U75 (N_75,In_374,In_969);
and U76 (N_76,In_10,In_649);
or U77 (N_77,In_172,In_185);
or U78 (N_78,In_67,In_757);
and U79 (N_79,In_555,In_49);
nand U80 (N_80,In_65,In_820);
nand U81 (N_81,In_956,In_234);
nand U82 (N_82,In_135,In_692);
and U83 (N_83,In_542,In_376);
and U84 (N_84,In_769,In_746);
and U85 (N_85,In_426,In_442);
nor U86 (N_86,In_4,In_767);
nand U87 (N_87,In_610,In_863);
or U88 (N_88,In_5,In_800);
or U89 (N_89,In_873,In_102);
or U90 (N_90,In_929,In_383);
or U91 (N_91,In_369,In_513);
xnor U92 (N_92,In_30,In_365);
nor U93 (N_93,In_309,In_99);
nor U94 (N_94,In_711,In_547);
xnor U95 (N_95,In_104,In_361);
and U96 (N_96,In_194,In_593);
and U97 (N_97,In_961,In_914);
and U98 (N_98,In_242,In_88);
and U99 (N_99,In_94,In_138);
xor U100 (N_100,In_401,In_663);
nand U101 (N_101,In_352,In_824);
nand U102 (N_102,In_188,In_399);
nor U103 (N_103,In_486,In_726);
xor U104 (N_104,In_642,In_857);
nand U105 (N_105,In_118,In_485);
or U106 (N_106,In_957,In_698);
nand U107 (N_107,In_226,In_545);
nor U108 (N_108,In_864,In_991);
nand U109 (N_109,In_670,In_748);
nand U110 (N_110,In_239,In_155);
and U111 (N_111,In_0,In_839);
nor U112 (N_112,In_784,In_216);
or U113 (N_113,In_228,In_717);
and U114 (N_114,In_533,In_499);
nor U115 (N_115,In_632,In_854);
nor U116 (N_116,In_315,In_628);
nand U117 (N_117,In_893,In_683);
xnor U118 (N_118,In_805,In_386);
nand U119 (N_119,In_27,In_659);
nor U120 (N_120,In_712,In_152);
and U121 (N_121,In_568,In_360);
or U122 (N_122,In_318,In_809);
or U123 (N_123,In_810,In_418);
nand U124 (N_124,In_336,In_275);
nand U125 (N_125,In_861,In_491);
and U126 (N_126,In_807,In_180);
and U127 (N_127,In_456,In_567);
nand U128 (N_128,In_330,In_208);
nor U129 (N_129,In_641,In_452);
and U130 (N_130,In_988,In_291);
and U131 (N_131,In_450,In_471);
nand U132 (N_132,In_372,In_968);
and U133 (N_133,In_189,In_107);
nand U134 (N_134,In_177,In_529);
nor U135 (N_135,In_967,In_749);
and U136 (N_136,In_532,In_939);
and U137 (N_137,In_287,In_582);
or U138 (N_138,In_205,In_920);
and U139 (N_139,In_601,In_994);
nor U140 (N_140,In_9,In_396);
or U141 (N_141,In_924,In_366);
or U142 (N_142,In_395,In_888);
nand U143 (N_143,In_802,In_523);
nor U144 (N_144,In_371,In_289);
nand U145 (N_145,In_458,In_701);
nor U146 (N_146,In_574,In_702);
and U147 (N_147,In_64,In_419);
or U148 (N_148,In_851,In_23);
or U149 (N_149,In_229,In_918);
nor U150 (N_150,In_121,In_744);
and U151 (N_151,In_141,In_167);
and U152 (N_152,In_355,In_422);
nand U153 (N_153,In_57,In_273);
nor U154 (N_154,In_584,In_930);
nor U155 (N_155,In_448,In_759);
or U156 (N_156,In_938,In_743);
nand U157 (N_157,In_53,In_675);
nand U158 (N_158,In_301,In_877);
nor U159 (N_159,In_390,In_551);
nand U160 (N_160,In_438,In_522);
nand U161 (N_161,In_43,In_342);
xnor U162 (N_162,In_541,In_353);
or U163 (N_163,In_592,In_344);
nor U164 (N_164,In_962,In_373);
or U165 (N_165,In_507,In_505);
xor U166 (N_166,In_136,In_254);
or U167 (N_167,In_145,In_81);
nand U168 (N_168,In_843,In_734);
nand U169 (N_169,In_612,In_1);
and U170 (N_170,In_790,In_83);
and U171 (N_171,In_462,In_274);
nand U172 (N_172,In_891,In_117);
and U173 (N_173,In_206,In_398);
nand U174 (N_174,In_90,In_878);
nand U175 (N_175,In_684,In_272);
xnor U176 (N_176,In_183,In_578);
and U177 (N_177,In_845,In_420);
nand U178 (N_178,In_453,In_527);
nor U179 (N_179,In_345,In_251);
or U180 (N_180,In_115,In_70);
nand U181 (N_181,In_50,In_440);
nand U182 (N_182,In_638,In_97);
xnor U183 (N_183,In_114,In_534);
and U184 (N_184,In_989,In_728);
and U185 (N_185,In_908,In_572);
or U186 (N_186,In_844,In_905);
nor U187 (N_187,In_143,In_656);
or U188 (N_188,In_85,In_588);
or U189 (N_189,In_585,In_82);
nor U190 (N_190,In_794,In_329);
nand U191 (N_191,In_37,In_444);
nand U192 (N_192,In_268,In_798);
nor U193 (N_193,In_697,In_652);
nand U194 (N_194,In_427,In_60);
and U195 (N_195,In_317,In_346);
nor U196 (N_196,In_441,In_327);
xor U197 (N_197,In_693,In_130);
nor U198 (N_198,In_106,In_783);
nor U199 (N_199,In_799,In_960);
nand U200 (N_200,In_482,In_326);
nand U201 (N_201,In_704,In_483);
xor U202 (N_202,In_409,In_887);
or U203 (N_203,In_546,In_919);
or U204 (N_204,In_846,In_341);
nand U205 (N_205,In_763,In_668);
nor U206 (N_206,In_525,In_665);
nor U207 (N_207,In_511,In_339);
and U208 (N_208,In_881,In_904);
nand U209 (N_209,In_316,In_223);
nand U210 (N_210,In_575,In_673);
nand U211 (N_211,In_245,In_633);
xnor U212 (N_212,In_402,In_620);
and U213 (N_213,In_359,In_524);
or U214 (N_214,In_435,In_168);
nand U215 (N_215,In_464,In_862);
or U216 (N_216,In_576,In_993);
nor U217 (N_217,In_101,In_613);
or U218 (N_218,In_110,In_46);
nor U219 (N_219,In_691,In_847);
nor U220 (N_220,In_506,In_445);
and U221 (N_221,In_296,In_209);
nor U222 (N_222,In_512,In_539);
nand U223 (N_223,In_977,In_222);
nor U224 (N_224,In_14,In_58);
and U225 (N_225,In_403,In_221);
and U226 (N_226,In_331,In_89);
nand U227 (N_227,In_127,In_335);
nor U228 (N_228,In_793,In_7);
and U229 (N_229,In_916,In_910);
or U230 (N_230,In_733,In_604);
nand U231 (N_231,In_986,In_741);
nor U232 (N_232,In_834,In_248);
or U233 (N_233,In_253,In_819);
or U234 (N_234,In_526,In_577);
and U235 (N_235,In_762,In_425);
or U236 (N_236,In_151,In_621);
and U237 (N_237,In_405,In_277);
nand U238 (N_238,In_745,In_952);
nor U239 (N_239,In_52,In_55);
and U240 (N_240,In_806,In_150);
or U241 (N_241,In_876,In_895);
nand U242 (N_242,In_695,In_123);
nand U243 (N_243,In_515,In_338);
nand U244 (N_244,In_134,In_560);
nor U245 (N_245,In_392,In_436);
or U246 (N_246,In_47,In_407);
nor U247 (N_247,In_414,In_657);
nand U248 (N_248,In_982,In_232);
nand U249 (N_249,In_990,In_39);
or U250 (N_250,In_487,In_661);
nor U251 (N_251,In_922,In_768);
or U252 (N_252,In_323,In_31);
and U253 (N_253,In_639,In_688);
or U254 (N_254,In_125,In_328);
nor U255 (N_255,In_278,In_159);
nand U256 (N_256,In_35,In_595);
and U257 (N_257,In_312,In_282);
xnor U258 (N_258,In_77,In_19);
and U259 (N_259,In_950,In_243);
nand U260 (N_260,In_264,In_321);
or U261 (N_261,In_473,In_368);
nor U262 (N_262,In_796,In_607);
nor U263 (N_263,In_211,In_433);
nand U264 (N_264,In_889,In_666);
nor U265 (N_265,In_214,In_926);
nor U266 (N_266,In_186,In_609);
and U267 (N_267,In_517,In_394);
and U268 (N_268,In_727,In_826);
and U269 (N_269,In_325,In_901);
nand U270 (N_270,In_149,In_970);
nand U271 (N_271,In_965,In_379);
nor U272 (N_272,In_400,In_459);
and U273 (N_273,In_596,In_852);
or U274 (N_274,In_559,In_730);
xnor U275 (N_275,In_333,In_816);
nand U276 (N_276,In_343,In_13);
nor U277 (N_277,In_856,In_421);
nand U278 (N_278,In_227,In_21);
and U279 (N_279,In_815,In_915);
or U280 (N_280,In_279,In_713);
and U281 (N_281,In_565,In_467);
nand U282 (N_282,In_71,In_87);
nor U283 (N_283,In_758,In_213);
and U284 (N_284,In_705,In_789);
or U285 (N_285,In_493,In_634);
nand U286 (N_286,In_432,In_516);
nand U287 (N_287,In_447,In_163);
nor U288 (N_288,In_6,In_685);
or U289 (N_289,In_590,In_812);
and U290 (N_290,In_230,In_774);
or U291 (N_291,In_267,In_643);
and U292 (N_292,In_797,In_11);
nor U293 (N_293,In_518,In_964);
nor U294 (N_294,In_837,In_801);
or U295 (N_295,In_286,In_126);
or U296 (N_296,In_497,In_26);
nor U297 (N_297,In_498,In_538);
nor U298 (N_298,In_283,In_756);
or U299 (N_299,In_896,In_200);
nor U300 (N_300,In_627,In_91);
nand U301 (N_301,In_776,In_937);
nor U302 (N_302,In_250,In_676);
or U303 (N_303,In_945,In_658);
or U304 (N_304,In_284,In_314);
and U305 (N_305,In_842,In_696);
and U306 (N_306,In_589,In_33);
nand U307 (N_307,In_667,In_298);
nand U308 (N_308,In_410,In_218);
nor U309 (N_309,In_17,In_514);
nor U310 (N_310,In_817,In_736);
nand U311 (N_311,In_468,In_912);
and U312 (N_312,In_98,In_237);
or U313 (N_313,In_597,In_570);
and U314 (N_314,In_179,In_803);
nand U315 (N_315,In_600,In_295);
nand U316 (N_316,In_474,In_18);
and U317 (N_317,In_201,In_966);
nor U318 (N_318,In_457,In_461);
or U319 (N_319,In_778,In_269);
nor U320 (N_320,In_528,In_319);
or U321 (N_321,In_59,In_690);
nand U322 (N_322,In_874,In_109);
and U323 (N_323,In_116,In_883);
and U324 (N_324,In_650,In_927);
nand U325 (N_325,In_165,In_220);
and U326 (N_326,In_255,In_169);
or U327 (N_327,In_446,In_217);
nand U328 (N_328,In_699,In_95);
or U329 (N_329,In_686,In_96);
nor U330 (N_330,In_680,In_449);
or U331 (N_331,In_174,In_36);
or U332 (N_332,In_20,In_363);
nand U333 (N_333,In_34,In_751);
nand U334 (N_334,In_781,In_504);
xnor U335 (N_335,In_981,In_870);
nor U336 (N_336,In_563,In_460);
nand U337 (N_337,In_995,In_569);
nor U338 (N_338,In_760,In_959);
and U339 (N_339,In_80,In_958);
or U340 (N_340,In_51,In_931);
nor U341 (N_341,In_16,In_503);
or U342 (N_342,In_178,In_246);
xnor U343 (N_343,In_509,In_488);
and U344 (N_344,In_955,In_241);
nand U345 (N_345,In_413,In_292);
or U346 (N_346,In_510,In_133);
or U347 (N_347,In_62,In_173);
nor U348 (N_348,In_651,In_865);
and U349 (N_349,In_548,In_928);
or U350 (N_350,In_521,In_540);
or U351 (N_351,In_247,In_478);
and U352 (N_352,In_719,In_351);
nand U353 (N_353,In_92,In_276);
nor U354 (N_354,In_535,In_775);
or U355 (N_355,In_943,In_266);
nand U356 (N_356,In_153,In_387);
or U357 (N_357,In_948,In_299);
or U358 (N_358,In_710,In_644);
and U359 (N_359,In_113,In_786);
nand U360 (N_360,In_231,In_378);
or U361 (N_361,In_941,In_764);
nand U362 (N_362,In_84,In_979);
or U363 (N_363,In_199,In_872);
nor U364 (N_364,In_671,In_496);
nand U365 (N_365,In_827,In_451);
nand U366 (N_366,In_936,In_431);
nand U367 (N_367,In_942,In_792);
and U368 (N_368,In_235,In_475);
or U369 (N_369,In_892,In_655);
nor U370 (N_370,In_616,In_388);
or U371 (N_371,In_40,In_848);
and U372 (N_372,In_56,In_42);
nand U373 (N_373,In_357,In_814);
and U374 (N_374,In_531,In_647);
nor U375 (N_375,In_859,In_811);
nor U376 (N_376,In_722,In_606);
nor U377 (N_377,In_598,In_731);
and U378 (N_378,In_992,In_397);
nor U379 (N_379,In_615,In_880);
nand U380 (N_380,In_44,In_192);
nor U381 (N_381,In_195,In_782);
and U382 (N_382,In_625,In_411);
nor U383 (N_383,In_470,In_742);
nand U384 (N_384,In_307,In_501);
nor U385 (N_385,In_265,In_304);
and U386 (N_386,In_679,In_999);
nor U387 (N_387,In_849,In_677);
nor U388 (N_388,In_385,In_86);
or U389 (N_389,In_766,In_573);
and U390 (N_390,In_182,In_479);
and U391 (N_391,In_752,In_389);
nor U392 (N_392,In_909,In_830);
and U393 (N_393,In_466,In_415);
and U394 (N_394,In_424,In_170);
and U395 (N_395,In_921,In_198);
and U396 (N_396,In_285,In_484);
nor U397 (N_397,In_624,In_754);
nor U398 (N_398,In_694,In_821);
nor U399 (N_399,In_637,In_591);
nand U400 (N_400,In_911,In_629);
nor U401 (N_401,In_791,In_480);
or U402 (N_402,In_73,In_879);
and U403 (N_403,In_947,In_181);
nand U404 (N_404,In_105,In_148);
nand U405 (N_405,In_554,In_520);
and U406 (N_406,In_614,In_290);
xnor U407 (N_407,In_773,In_611);
nor U408 (N_408,In_875,In_687);
nand U409 (N_409,In_828,In_219);
nor U410 (N_410,In_79,In_428);
and U411 (N_411,In_297,In_202);
and U412 (N_412,In_944,In_112);
or U413 (N_413,In_204,In_972);
nor U414 (N_414,In_884,In_196);
nor U415 (N_415,In_472,In_867);
nand U416 (N_416,In_543,In_836);
or U417 (N_417,In_322,In_12);
nand U418 (N_418,In_430,In_871);
xor U419 (N_419,In_187,In_721);
nor U420 (N_420,In_293,In_259);
nand U421 (N_421,In_648,In_985);
and U422 (N_422,In_303,In_29);
nor U423 (N_423,In_193,In_281);
and U424 (N_424,In_818,In_672);
and U425 (N_425,In_890,In_732);
xor U426 (N_426,In_838,In_906);
or U427 (N_427,In_320,In_603);
or U428 (N_428,In_630,In_166);
nor U429 (N_429,In_953,In_795);
and U430 (N_430,In_913,In_494);
or U431 (N_431,In_131,In_619);
or U432 (N_432,In_358,In_311);
or U433 (N_433,In_175,In_45);
xor U434 (N_434,In_935,In_770);
nor U435 (N_435,In_765,In_946);
and U436 (N_436,In_898,In_581);
nor U437 (N_437,In_934,In_332);
and U438 (N_438,In_594,In_423);
or U439 (N_439,In_416,In_617);
or U440 (N_440,In_261,In_750);
nor U441 (N_441,In_976,In_983);
nand U442 (N_442,In_22,In_477);
and U443 (N_443,In_975,In_63);
and U444 (N_444,In_139,In_700);
and U445 (N_445,In_252,In_481);
nor U446 (N_446,In_362,In_404);
nand U447 (N_447,In_866,In_954);
or U448 (N_448,In_157,In_833);
and U449 (N_449,In_144,In_536);
or U450 (N_450,In_949,In_429);
nor U451 (N_451,In_855,In_987);
and U452 (N_452,In_154,In_381);
or U453 (N_453,In_832,In_998);
and U454 (N_454,In_640,In_602);
nand U455 (N_455,In_653,In_858);
or U456 (N_456,In_72,In_822);
nand U457 (N_457,In_636,In_825);
and U458 (N_458,In_580,In_608);
or U459 (N_459,In_850,In_772);
nor U460 (N_460,In_706,In_755);
nand U461 (N_461,In_645,In_678);
nor U462 (N_462,In_262,In_902);
nor U463 (N_463,In_124,In_530);
nor U464 (N_464,In_100,In_32);
nor U465 (N_465,In_841,In_787);
nand U466 (N_466,In_161,In_25);
and U467 (N_467,In_160,In_74);
or U468 (N_468,In_68,In_370);
or U469 (N_469,In_869,In_324);
and U470 (N_470,In_980,In_75);
and U471 (N_471,In_305,In_465);
nand U472 (N_472,In_587,In_334);
nand U473 (N_473,In_886,In_69);
nor U474 (N_474,In_24,In_622);
nand U475 (N_475,In_831,In_860);
nand U476 (N_476,In_38,In_380);
and U477 (N_477,In_108,In_553);
nor U478 (N_478,In_375,In_537);
nand U479 (N_479,In_492,In_788);
xnor U480 (N_480,In_689,In_147);
nor U481 (N_481,In_835,In_300);
nand U482 (N_482,In_140,In_443);
nand U483 (N_483,In_256,In_586);
or U484 (N_484,In_971,In_674);
nand U485 (N_485,In_823,In_779);
nand U486 (N_486,In_233,In_454);
nor U487 (N_487,In_350,In_894);
nor U488 (N_488,In_813,In_406);
nor U489 (N_489,In_660,In_723);
nand U490 (N_490,In_132,In_519);
or U491 (N_491,In_215,In_434);
or U492 (N_492,In_93,In_579);
nand U493 (N_493,In_738,In_951);
xnor U494 (N_494,In_412,In_66);
nor U495 (N_495,In_122,In_294);
nor U496 (N_496,In_41,In_238);
and U497 (N_497,In_556,In_2);
nor U498 (N_498,In_156,In_681);
xnor U499 (N_499,In_709,In_263);
and U500 (N_500,In_531,In_268);
and U501 (N_501,In_644,In_45);
and U502 (N_502,In_394,In_626);
and U503 (N_503,In_356,In_304);
and U504 (N_504,In_997,In_577);
nand U505 (N_505,In_425,In_941);
nor U506 (N_506,In_167,In_490);
or U507 (N_507,In_280,In_223);
and U508 (N_508,In_434,In_363);
nand U509 (N_509,In_566,In_838);
nand U510 (N_510,In_427,In_812);
nor U511 (N_511,In_312,In_209);
nor U512 (N_512,In_236,In_955);
and U513 (N_513,In_199,In_921);
and U514 (N_514,In_608,In_395);
nand U515 (N_515,In_368,In_510);
nor U516 (N_516,In_401,In_470);
and U517 (N_517,In_47,In_403);
and U518 (N_518,In_889,In_418);
and U519 (N_519,In_173,In_838);
and U520 (N_520,In_180,In_679);
or U521 (N_521,In_428,In_349);
nand U522 (N_522,In_296,In_708);
nor U523 (N_523,In_66,In_506);
nand U524 (N_524,In_414,In_480);
nor U525 (N_525,In_179,In_277);
nor U526 (N_526,In_597,In_827);
or U527 (N_527,In_664,In_140);
and U528 (N_528,In_652,In_766);
nand U529 (N_529,In_515,In_447);
nand U530 (N_530,In_364,In_342);
and U531 (N_531,In_732,In_277);
nor U532 (N_532,In_860,In_791);
nor U533 (N_533,In_723,In_988);
nand U534 (N_534,In_929,In_651);
or U535 (N_535,In_906,In_430);
or U536 (N_536,In_676,In_243);
or U537 (N_537,In_920,In_102);
nor U538 (N_538,In_720,In_526);
or U539 (N_539,In_207,In_436);
and U540 (N_540,In_241,In_412);
or U541 (N_541,In_702,In_963);
nor U542 (N_542,In_680,In_639);
nor U543 (N_543,In_626,In_310);
and U544 (N_544,In_205,In_717);
nand U545 (N_545,In_471,In_996);
nand U546 (N_546,In_220,In_351);
and U547 (N_547,In_53,In_377);
or U548 (N_548,In_435,In_466);
and U549 (N_549,In_254,In_160);
and U550 (N_550,In_162,In_597);
or U551 (N_551,In_980,In_385);
or U552 (N_552,In_388,In_485);
nand U553 (N_553,In_650,In_614);
and U554 (N_554,In_431,In_817);
or U555 (N_555,In_429,In_315);
and U556 (N_556,In_776,In_242);
nand U557 (N_557,In_596,In_166);
and U558 (N_558,In_321,In_224);
or U559 (N_559,In_377,In_985);
nor U560 (N_560,In_1,In_166);
or U561 (N_561,In_765,In_80);
and U562 (N_562,In_577,In_717);
and U563 (N_563,In_979,In_343);
nor U564 (N_564,In_100,In_914);
nor U565 (N_565,In_315,In_40);
or U566 (N_566,In_218,In_539);
or U567 (N_567,In_270,In_542);
and U568 (N_568,In_334,In_246);
nor U569 (N_569,In_573,In_623);
or U570 (N_570,In_753,In_717);
or U571 (N_571,In_299,In_544);
nor U572 (N_572,In_156,In_562);
nor U573 (N_573,In_402,In_969);
or U574 (N_574,In_179,In_441);
nor U575 (N_575,In_280,In_439);
xnor U576 (N_576,In_47,In_204);
or U577 (N_577,In_915,In_674);
nor U578 (N_578,In_741,In_123);
nand U579 (N_579,In_476,In_572);
and U580 (N_580,In_760,In_202);
nand U581 (N_581,In_911,In_390);
nor U582 (N_582,In_444,In_328);
nor U583 (N_583,In_80,In_502);
nand U584 (N_584,In_785,In_921);
or U585 (N_585,In_95,In_236);
or U586 (N_586,In_791,In_264);
and U587 (N_587,In_157,In_741);
or U588 (N_588,In_979,In_753);
or U589 (N_589,In_62,In_942);
or U590 (N_590,In_364,In_389);
and U591 (N_591,In_415,In_126);
nand U592 (N_592,In_314,In_984);
nand U593 (N_593,In_965,In_149);
and U594 (N_594,In_698,In_430);
nor U595 (N_595,In_485,In_432);
nand U596 (N_596,In_291,In_589);
nand U597 (N_597,In_803,In_777);
nor U598 (N_598,In_717,In_72);
xor U599 (N_599,In_346,In_361);
or U600 (N_600,In_292,In_279);
nor U601 (N_601,In_720,In_99);
and U602 (N_602,In_343,In_47);
and U603 (N_603,In_381,In_734);
nor U604 (N_604,In_23,In_60);
and U605 (N_605,In_561,In_240);
or U606 (N_606,In_125,In_698);
and U607 (N_607,In_923,In_672);
and U608 (N_608,In_487,In_831);
nand U609 (N_609,In_347,In_607);
nor U610 (N_610,In_977,In_124);
or U611 (N_611,In_110,In_887);
nand U612 (N_612,In_823,In_485);
nand U613 (N_613,In_41,In_181);
or U614 (N_614,In_777,In_759);
and U615 (N_615,In_542,In_609);
nand U616 (N_616,In_744,In_92);
and U617 (N_617,In_295,In_484);
nand U618 (N_618,In_214,In_197);
nor U619 (N_619,In_248,In_535);
nand U620 (N_620,In_639,In_963);
nand U621 (N_621,In_742,In_988);
nor U622 (N_622,In_779,In_72);
or U623 (N_623,In_404,In_983);
and U624 (N_624,In_689,In_572);
nor U625 (N_625,In_547,In_702);
nor U626 (N_626,In_122,In_640);
nand U627 (N_627,In_560,In_792);
nor U628 (N_628,In_181,In_656);
and U629 (N_629,In_788,In_120);
nand U630 (N_630,In_445,In_103);
or U631 (N_631,In_298,In_67);
nand U632 (N_632,In_187,In_790);
nand U633 (N_633,In_235,In_773);
and U634 (N_634,In_298,In_401);
nor U635 (N_635,In_368,In_742);
and U636 (N_636,In_255,In_330);
nor U637 (N_637,In_940,In_917);
nand U638 (N_638,In_721,In_499);
and U639 (N_639,In_105,In_752);
nor U640 (N_640,In_907,In_140);
or U641 (N_641,In_994,In_951);
nand U642 (N_642,In_968,In_872);
and U643 (N_643,In_745,In_39);
nand U644 (N_644,In_591,In_23);
nor U645 (N_645,In_77,In_781);
xor U646 (N_646,In_365,In_26);
and U647 (N_647,In_172,In_617);
nand U648 (N_648,In_840,In_733);
and U649 (N_649,In_908,In_87);
or U650 (N_650,In_194,In_704);
and U651 (N_651,In_157,In_854);
and U652 (N_652,In_811,In_660);
nor U653 (N_653,In_446,In_672);
or U654 (N_654,In_732,In_930);
nand U655 (N_655,In_887,In_880);
nand U656 (N_656,In_736,In_12);
nor U657 (N_657,In_519,In_347);
nand U658 (N_658,In_706,In_588);
nand U659 (N_659,In_312,In_48);
and U660 (N_660,In_31,In_280);
xor U661 (N_661,In_464,In_80);
nor U662 (N_662,In_937,In_12);
and U663 (N_663,In_228,In_676);
nor U664 (N_664,In_853,In_35);
or U665 (N_665,In_584,In_157);
and U666 (N_666,In_150,In_854);
nor U667 (N_667,In_663,In_918);
nand U668 (N_668,In_972,In_565);
and U669 (N_669,In_984,In_445);
nor U670 (N_670,In_321,In_234);
nand U671 (N_671,In_45,In_219);
and U672 (N_672,In_598,In_457);
or U673 (N_673,In_705,In_213);
and U674 (N_674,In_398,In_583);
nand U675 (N_675,In_206,In_576);
and U676 (N_676,In_997,In_189);
nand U677 (N_677,In_74,In_93);
and U678 (N_678,In_344,In_217);
nor U679 (N_679,In_907,In_606);
nand U680 (N_680,In_361,In_695);
nand U681 (N_681,In_229,In_352);
nor U682 (N_682,In_988,In_423);
nor U683 (N_683,In_772,In_779);
and U684 (N_684,In_814,In_661);
nand U685 (N_685,In_286,In_926);
nand U686 (N_686,In_359,In_258);
and U687 (N_687,In_461,In_550);
or U688 (N_688,In_413,In_185);
and U689 (N_689,In_494,In_1);
and U690 (N_690,In_596,In_96);
or U691 (N_691,In_944,In_309);
nor U692 (N_692,In_379,In_50);
nand U693 (N_693,In_104,In_160);
or U694 (N_694,In_978,In_516);
nor U695 (N_695,In_454,In_228);
or U696 (N_696,In_696,In_624);
xor U697 (N_697,In_937,In_625);
nor U698 (N_698,In_158,In_770);
nor U699 (N_699,In_143,In_626);
and U700 (N_700,In_241,In_362);
nand U701 (N_701,In_474,In_123);
or U702 (N_702,In_27,In_581);
or U703 (N_703,In_815,In_820);
nand U704 (N_704,In_570,In_198);
and U705 (N_705,In_455,In_142);
xor U706 (N_706,In_899,In_814);
nand U707 (N_707,In_167,In_320);
nand U708 (N_708,In_77,In_780);
nor U709 (N_709,In_474,In_895);
and U710 (N_710,In_132,In_609);
nand U711 (N_711,In_418,In_659);
or U712 (N_712,In_224,In_278);
nand U713 (N_713,In_23,In_516);
nor U714 (N_714,In_117,In_39);
nor U715 (N_715,In_318,In_314);
nor U716 (N_716,In_835,In_698);
nand U717 (N_717,In_292,In_816);
nand U718 (N_718,In_871,In_980);
or U719 (N_719,In_305,In_85);
nor U720 (N_720,In_184,In_870);
and U721 (N_721,In_512,In_949);
nand U722 (N_722,In_135,In_869);
nor U723 (N_723,In_265,In_197);
or U724 (N_724,In_352,In_353);
and U725 (N_725,In_421,In_9);
or U726 (N_726,In_748,In_220);
or U727 (N_727,In_404,In_331);
and U728 (N_728,In_115,In_105);
nand U729 (N_729,In_4,In_204);
and U730 (N_730,In_186,In_926);
nor U731 (N_731,In_378,In_880);
or U732 (N_732,In_777,In_537);
nor U733 (N_733,In_854,In_101);
or U734 (N_734,In_434,In_37);
nand U735 (N_735,In_128,In_426);
nand U736 (N_736,In_377,In_64);
and U737 (N_737,In_481,In_408);
nor U738 (N_738,In_800,In_538);
and U739 (N_739,In_188,In_502);
or U740 (N_740,In_194,In_221);
and U741 (N_741,In_960,In_96);
nor U742 (N_742,In_38,In_464);
nand U743 (N_743,In_458,In_719);
and U744 (N_744,In_915,In_240);
nand U745 (N_745,In_545,In_164);
nor U746 (N_746,In_928,In_649);
nand U747 (N_747,In_252,In_672);
nor U748 (N_748,In_386,In_409);
and U749 (N_749,In_914,In_263);
nand U750 (N_750,In_723,In_564);
and U751 (N_751,In_842,In_972);
nor U752 (N_752,In_514,In_408);
or U753 (N_753,In_428,In_484);
and U754 (N_754,In_901,In_60);
nor U755 (N_755,In_204,In_771);
nor U756 (N_756,In_269,In_10);
and U757 (N_757,In_844,In_76);
nor U758 (N_758,In_415,In_815);
and U759 (N_759,In_996,In_530);
nand U760 (N_760,In_129,In_931);
nand U761 (N_761,In_538,In_518);
and U762 (N_762,In_633,In_60);
nand U763 (N_763,In_808,In_163);
xor U764 (N_764,In_500,In_290);
nor U765 (N_765,In_867,In_340);
nor U766 (N_766,In_634,In_672);
and U767 (N_767,In_494,In_7);
and U768 (N_768,In_287,In_337);
nand U769 (N_769,In_686,In_384);
nand U770 (N_770,In_447,In_553);
nand U771 (N_771,In_316,In_350);
nor U772 (N_772,In_607,In_454);
and U773 (N_773,In_349,In_310);
or U774 (N_774,In_631,In_505);
nor U775 (N_775,In_226,In_947);
or U776 (N_776,In_592,In_654);
nor U777 (N_777,In_661,In_17);
nand U778 (N_778,In_773,In_446);
nor U779 (N_779,In_174,In_195);
nor U780 (N_780,In_668,In_600);
nand U781 (N_781,In_670,In_333);
nand U782 (N_782,In_725,In_586);
or U783 (N_783,In_955,In_252);
nor U784 (N_784,In_538,In_708);
nand U785 (N_785,In_596,In_633);
and U786 (N_786,In_201,In_125);
and U787 (N_787,In_436,In_864);
nor U788 (N_788,In_100,In_947);
nand U789 (N_789,In_14,In_674);
and U790 (N_790,In_755,In_106);
or U791 (N_791,In_51,In_356);
nor U792 (N_792,In_646,In_706);
and U793 (N_793,In_207,In_777);
and U794 (N_794,In_995,In_677);
nand U795 (N_795,In_498,In_501);
nand U796 (N_796,In_640,In_128);
and U797 (N_797,In_340,In_433);
nor U798 (N_798,In_498,In_812);
xnor U799 (N_799,In_930,In_145);
nand U800 (N_800,In_7,In_725);
nand U801 (N_801,In_184,In_341);
nand U802 (N_802,In_845,In_958);
and U803 (N_803,In_999,In_392);
and U804 (N_804,In_355,In_295);
and U805 (N_805,In_177,In_696);
nor U806 (N_806,In_341,In_206);
nand U807 (N_807,In_945,In_794);
xor U808 (N_808,In_259,In_819);
nand U809 (N_809,In_380,In_841);
nand U810 (N_810,In_25,In_781);
nand U811 (N_811,In_141,In_401);
and U812 (N_812,In_453,In_318);
nand U813 (N_813,In_801,In_931);
nor U814 (N_814,In_570,In_728);
or U815 (N_815,In_25,In_477);
nand U816 (N_816,In_752,In_746);
and U817 (N_817,In_678,In_206);
or U818 (N_818,In_799,In_528);
nor U819 (N_819,In_994,In_262);
nor U820 (N_820,In_246,In_861);
nand U821 (N_821,In_133,In_840);
nor U822 (N_822,In_824,In_774);
or U823 (N_823,In_54,In_481);
nor U824 (N_824,In_311,In_574);
or U825 (N_825,In_289,In_214);
nor U826 (N_826,In_921,In_883);
nand U827 (N_827,In_516,In_879);
and U828 (N_828,In_140,In_494);
and U829 (N_829,In_159,In_609);
and U830 (N_830,In_784,In_552);
and U831 (N_831,In_426,In_335);
nand U832 (N_832,In_243,In_705);
nand U833 (N_833,In_711,In_852);
nor U834 (N_834,In_721,In_797);
nor U835 (N_835,In_74,In_417);
and U836 (N_836,In_6,In_964);
and U837 (N_837,In_103,In_765);
or U838 (N_838,In_80,In_955);
nor U839 (N_839,In_834,In_578);
nor U840 (N_840,In_818,In_445);
xnor U841 (N_841,In_239,In_880);
and U842 (N_842,In_43,In_671);
and U843 (N_843,In_663,In_208);
and U844 (N_844,In_509,In_890);
nor U845 (N_845,In_990,In_588);
and U846 (N_846,In_243,In_319);
or U847 (N_847,In_297,In_82);
and U848 (N_848,In_582,In_477);
nor U849 (N_849,In_651,In_943);
nor U850 (N_850,In_431,In_924);
and U851 (N_851,In_579,In_878);
nor U852 (N_852,In_470,In_943);
and U853 (N_853,In_273,In_479);
or U854 (N_854,In_810,In_155);
nor U855 (N_855,In_354,In_531);
and U856 (N_856,In_361,In_166);
nor U857 (N_857,In_238,In_84);
and U858 (N_858,In_926,In_797);
nor U859 (N_859,In_591,In_931);
or U860 (N_860,In_229,In_344);
nand U861 (N_861,In_265,In_735);
nand U862 (N_862,In_612,In_868);
nor U863 (N_863,In_793,In_803);
or U864 (N_864,In_0,In_337);
nor U865 (N_865,In_147,In_268);
nand U866 (N_866,In_231,In_905);
nor U867 (N_867,In_629,In_157);
or U868 (N_868,In_705,In_593);
or U869 (N_869,In_961,In_231);
nand U870 (N_870,In_713,In_409);
and U871 (N_871,In_39,In_52);
nor U872 (N_872,In_874,In_344);
and U873 (N_873,In_442,In_419);
nand U874 (N_874,In_405,In_895);
or U875 (N_875,In_429,In_406);
nor U876 (N_876,In_327,In_664);
and U877 (N_877,In_747,In_630);
nand U878 (N_878,In_523,In_195);
or U879 (N_879,In_9,In_199);
nand U880 (N_880,In_296,In_690);
or U881 (N_881,In_969,In_294);
nor U882 (N_882,In_864,In_442);
nor U883 (N_883,In_785,In_766);
and U884 (N_884,In_168,In_449);
or U885 (N_885,In_971,In_441);
nand U886 (N_886,In_623,In_809);
nand U887 (N_887,In_909,In_186);
nor U888 (N_888,In_857,In_509);
nor U889 (N_889,In_795,In_408);
or U890 (N_890,In_62,In_193);
or U891 (N_891,In_163,In_817);
or U892 (N_892,In_609,In_42);
nand U893 (N_893,In_928,In_793);
nand U894 (N_894,In_800,In_690);
nand U895 (N_895,In_812,In_544);
nand U896 (N_896,In_634,In_177);
nand U897 (N_897,In_63,In_998);
or U898 (N_898,In_536,In_474);
nand U899 (N_899,In_653,In_172);
and U900 (N_900,In_389,In_935);
or U901 (N_901,In_431,In_320);
nor U902 (N_902,In_794,In_311);
nor U903 (N_903,In_524,In_2);
nor U904 (N_904,In_735,In_14);
and U905 (N_905,In_273,In_165);
nand U906 (N_906,In_267,In_769);
or U907 (N_907,In_120,In_769);
and U908 (N_908,In_343,In_367);
and U909 (N_909,In_4,In_920);
and U910 (N_910,In_535,In_998);
or U911 (N_911,In_399,In_630);
nand U912 (N_912,In_730,In_234);
or U913 (N_913,In_313,In_223);
nand U914 (N_914,In_452,In_161);
nand U915 (N_915,In_817,In_545);
nor U916 (N_916,In_915,In_428);
nor U917 (N_917,In_516,In_188);
nand U918 (N_918,In_477,In_594);
and U919 (N_919,In_601,In_140);
and U920 (N_920,In_50,In_847);
and U921 (N_921,In_5,In_186);
or U922 (N_922,In_517,In_969);
or U923 (N_923,In_494,In_428);
nand U924 (N_924,In_371,In_168);
or U925 (N_925,In_428,In_68);
nor U926 (N_926,In_871,In_400);
or U927 (N_927,In_951,In_417);
and U928 (N_928,In_771,In_898);
nor U929 (N_929,In_227,In_860);
and U930 (N_930,In_211,In_667);
or U931 (N_931,In_448,In_943);
nor U932 (N_932,In_875,In_75);
nor U933 (N_933,In_490,In_660);
nand U934 (N_934,In_821,In_354);
or U935 (N_935,In_842,In_122);
or U936 (N_936,In_422,In_285);
or U937 (N_937,In_98,In_957);
and U938 (N_938,In_283,In_382);
or U939 (N_939,In_702,In_250);
nor U940 (N_940,In_450,In_587);
nor U941 (N_941,In_179,In_218);
and U942 (N_942,In_255,In_235);
nor U943 (N_943,In_97,In_386);
and U944 (N_944,In_437,In_408);
or U945 (N_945,In_481,In_285);
nand U946 (N_946,In_105,In_626);
nand U947 (N_947,In_292,In_460);
and U948 (N_948,In_144,In_540);
or U949 (N_949,In_724,In_749);
and U950 (N_950,In_105,In_202);
nand U951 (N_951,In_880,In_55);
and U952 (N_952,In_133,In_816);
or U953 (N_953,In_603,In_419);
nor U954 (N_954,In_856,In_879);
nand U955 (N_955,In_328,In_829);
and U956 (N_956,In_702,In_641);
nor U957 (N_957,In_387,In_959);
and U958 (N_958,In_510,In_316);
nand U959 (N_959,In_402,In_448);
and U960 (N_960,In_23,In_223);
nand U961 (N_961,In_605,In_957);
nor U962 (N_962,In_53,In_816);
and U963 (N_963,In_828,In_809);
nand U964 (N_964,In_537,In_720);
or U965 (N_965,In_40,In_350);
nand U966 (N_966,In_75,In_452);
nand U967 (N_967,In_803,In_938);
nor U968 (N_968,In_850,In_466);
or U969 (N_969,In_434,In_872);
nand U970 (N_970,In_236,In_688);
nand U971 (N_971,In_963,In_66);
nand U972 (N_972,In_276,In_320);
nor U973 (N_973,In_277,In_399);
nand U974 (N_974,In_997,In_915);
and U975 (N_975,In_97,In_59);
or U976 (N_976,In_832,In_982);
and U977 (N_977,In_815,In_37);
nor U978 (N_978,In_802,In_408);
nand U979 (N_979,In_423,In_427);
or U980 (N_980,In_163,In_330);
nand U981 (N_981,In_762,In_347);
xnor U982 (N_982,In_742,In_189);
nand U983 (N_983,In_990,In_614);
and U984 (N_984,In_417,In_634);
nand U985 (N_985,In_31,In_834);
nor U986 (N_986,In_246,In_825);
or U987 (N_987,In_100,In_653);
nand U988 (N_988,In_749,In_413);
nand U989 (N_989,In_581,In_174);
or U990 (N_990,In_772,In_361);
or U991 (N_991,In_448,In_546);
and U992 (N_992,In_727,In_235);
nand U993 (N_993,In_80,In_270);
and U994 (N_994,In_482,In_291);
nor U995 (N_995,In_156,In_865);
and U996 (N_996,In_329,In_336);
nor U997 (N_997,In_106,In_344);
and U998 (N_998,In_969,In_855);
and U999 (N_999,In_798,In_205);
nand U1000 (N_1000,In_706,In_686);
and U1001 (N_1001,In_950,In_205);
xor U1002 (N_1002,In_766,In_177);
nor U1003 (N_1003,In_510,In_849);
nor U1004 (N_1004,In_191,In_655);
nand U1005 (N_1005,In_899,In_958);
and U1006 (N_1006,In_807,In_461);
nand U1007 (N_1007,In_300,In_981);
or U1008 (N_1008,In_250,In_440);
nand U1009 (N_1009,In_984,In_896);
nand U1010 (N_1010,In_315,In_874);
or U1011 (N_1011,In_515,In_687);
and U1012 (N_1012,In_11,In_708);
nand U1013 (N_1013,In_545,In_782);
or U1014 (N_1014,In_185,In_331);
nor U1015 (N_1015,In_412,In_667);
nor U1016 (N_1016,In_425,In_825);
or U1017 (N_1017,In_254,In_452);
and U1018 (N_1018,In_185,In_938);
and U1019 (N_1019,In_890,In_860);
nand U1020 (N_1020,In_100,In_902);
xnor U1021 (N_1021,In_194,In_210);
nor U1022 (N_1022,In_874,In_592);
xnor U1023 (N_1023,In_155,In_510);
or U1024 (N_1024,In_546,In_537);
nand U1025 (N_1025,In_679,In_920);
nor U1026 (N_1026,In_857,In_542);
and U1027 (N_1027,In_496,In_193);
or U1028 (N_1028,In_637,In_531);
nand U1029 (N_1029,In_614,In_214);
nand U1030 (N_1030,In_653,In_763);
or U1031 (N_1031,In_425,In_96);
nor U1032 (N_1032,In_930,In_988);
and U1033 (N_1033,In_976,In_784);
nand U1034 (N_1034,In_246,In_504);
nand U1035 (N_1035,In_317,In_32);
and U1036 (N_1036,In_727,In_621);
and U1037 (N_1037,In_582,In_740);
nor U1038 (N_1038,In_209,In_630);
and U1039 (N_1039,In_120,In_457);
nand U1040 (N_1040,In_164,In_403);
and U1041 (N_1041,In_114,In_601);
nand U1042 (N_1042,In_661,In_624);
and U1043 (N_1043,In_615,In_25);
nand U1044 (N_1044,In_755,In_554);
nor U1045 (N_1045,In_341,In_494);
and U1046 (N_1046,In_315,In_232);
or U1047 (N_1047,In_259,In_311);
nor U1048 (N_1048,In_221,In_756);
or U1049 (N_1049,In_247,In_557);
nor U1050 (N_1050,In_140,In_8);
and U1051 (N_1051,In_980,In_391);
nand U1052 (N_1052,In_392,In_756);
nand U1053 (N_1053,In_622,In_734);
and U1054 (N_1054,In_683,In_687);
nor U1055 (N_1055,In_353,In_573);
nand U1056 (N_1056,In_554,In_614);
and U1057 (N_1057,In_956,In_271);
or U1058 (N_1058,In_626,In_780);
nand U1059 (N_1059,In_348,In_692);
or U1060 (N_1060,In_961,In_82);
or U1061 (N_1061,In_20,In_642);
nand U1062 (N_1062,In_778,In_878);
nand U1063 (N_1063,In_409,In_586);
and U1064 (N_1064,In_913,In_42);
nor U1065 (N_1065,In_614,In_792);
or U1066 (N_1066,In_125,In_520);
xor U1067 (N_1067,In_908,In_885);
or U1068 (N_1068,In_34,In_80);
xnor U1069 (N_1069,In_810,In_165);
nand U1070 (N_1070,In_237,In_129);
or U1071 (N_1071,In_57,In_529);
nand U1072 (N_1072,In_30,In_19);
nand U1073 (N_1073,In_806,In_558);
or U1074 (N_1074,In_190,In_315);
or U1075 (N_1075,In_925,In_120);
nand U1076 (N_1076,In_265,In_910);
or U1077 (N_1077,In_461,In_201);
and U1078 (N_1078,In_147,In_289);
and U1079 (N_1079,In_84,In_268);
nor U1080 (N_1080,In_785,In_148);
and U1081 (N_1081,In_456,In_848);
nand U1082 (N_1082,In_399,In_835);
and U1083 (N_1083,In_565,In_656);
nand U1084 (N_1084,In_11,In_148);
or U1085 (N_1085,In_912,In_67);
and U1086 (N_1086,In_893,In_503);
nor U1087 (N_1087,In_788,In_275);
nor U1088 (N_1088,In_387,In_840);
nor U1089 (N_1089,In_835,In_198);
nor U1090 (N_1090,In_606,In_39);
or U1091 (N_1091,In_857,In_913);
nor U1092 (N_1092,In_964,In_762);
nor U1093 (N_1093,In_191,In_353);
nor U1094 (N_1094,In_489,In_757);
and U1095 (N_1095,In_952,In_748);
and U1096 (N_1096,In_406,In_490);
nor U1097 (N_1097,In_832,In_483);
nor U1098 (N_1098,In_81,In_997);
nand U1099 (N_1099,In_891,In_968);
nor U1100 (N_1100,In_625,In_531);
nand U1101 (N_1101,In_69,In_421);
and U1102 (N_1102,In_688,In_260);
nand U1103 (N_1103,In_670,In_102);
or U1104 (N_1104,In_865,In_201);
and U1105 (N_1105,In_397,In_123);
and U1106 (N_1106,In_205,In_803);
nor U1107 (N_1107,In_446,In_113);
nor U1108 (N_1108,In_155,In_833);
nor U1109 (N_1109,In_632,In_941);
or U1110 (N_1110,In_993,In_609);
nor U1111 (N_1111,In_522,In_465);
and U1112 (N_1112,In_177,In_726);
or U1113 (N_1113,In_407,In_836);
and U1114 (N_1114,In_405,In_85);
nor U1115 (N_1115,In_91,In_857);
and U1116 (N_1116,In_976,In_449);
or U1117 (N_1117,In_341,In_263);
or U1118 (N_1118,In_256,In_410);
or U1119 (N_1119,In_648,In_461);
and U1120 (N_1120,In_342,In_888);
or U1121 (N_1121,In_543,In_143);
or U1122 (N_1122,In_442,In_813);
or U1123 (N_1123,In_702,In_817);
and U1124 (N_1124,In_725,In_204);
or U1125 (N_1125,In_926,In_207);
or U1126 (N_1126,In_361,In_448);
and U1127 (N_1127,In_468,In_372);
nand U1128 (N_1128,In_254,In_477);
and U1129 (N_1129,In_776,In_85);
nor U1130 (N_1130,In_616,In_376);
nor U1131 (N_1131,In_982,In_826);
nand U1132 (N_1132,In_684,In_283);
nor U1133 (N_1133,In_851,In_289);
and U1134 (N_1134,In_659,In_790);
or U1135 (N_1135,In_953,In_829);
or U1136 (N_1136,In_807,In_923);
nand U1137 (N_1137,In_155,In_408);
nand U1138 (N_1138,In_442,In_206);
or U1139 (N_1139,In_500,In_204);
nor U1140 (N_1140,In_687,In_812);
or U1141 (N_1141,In_629,In_858);
and U1142 (N_1142,In_138,In_595);
nand U1143 (N_1143,In_584,In_453);
or U1144 (N_1144,In_106,In_634);
nor U1145 (N_1145,In_626,In_360);
nor U1146 (N_1146,In_24,In_449);
nand U1147 (N_1147,In_311,In_678);
nand U1148 (N_1148,In_966,In_483);
and U1149 (N_1149,In_667,In_702);
and U1150 (N_1150,In_326,In_416);
nor U1151 (N_1151,In_27,In_116);
nor U1152 (N_1152,In_345,In_879);
and U1153 (N_1153,In_299,In_1);
or U1154 (N_1154,In_800,In_323);
nor U1155 (N_1155,In_777,In_769);
nand U1156 (N_1156,In_532,In_725);
nor U1157 (N_1157,In_157,In_625);
nand U1158 (N_1158,In_929,In_401);
nor U1159 (N_1159,In_284,In_31);
nand U1160 (N_1160,In_688,In_675);
or U1161 (N_1161,In_209,In_372);
and U1162 (N_1162,In_989,In_123);
nor U1163 (N_1163,In_582,In_152);
nor U1164 (N_1164,In_995,In_395);
and U1165 (N_1165,In_512,In_697);
nor U1166 (N_1166,In_156,In_211);
nor U1167 (N_1167,In_368,In_382);
nand U1168 (N_1168,In_280,In_414);
or U1169 (N_1169,In_719,In_970);
and U1170 (N_1170,In_918,In_17);
and U1171 (N_1171,In_639,In_591);
nor U1172 (N_1172,In_825,In_737);
nor U1173 (N_1173,In_474,In_917);
nand U1174 (N_1174,In_33,In_747);
nand U1175 (N_1175,In_580,In_129);
nor U1176 (N_1176,In_653,In_14);
nand U1177 (N_1177,In_441,In_491);
and U1178 (N_1178,In_609,In_468);
or U1179 (N_1179,In_138,In_710);
or U1180 (N_1180,In_177,In_489);
nand U1181 (N_1181,In_380,In_718);
or U1182 (N_1182,In_808,In_885);
or U1183 (N_1183,In_124,In_957);
and U1184 (N_1184,In_896,In_389);
nand U1185 (N_1185,In_921,In_456);
nand U1186 (N_1186,In_150,In_620);
nand U1187 (N_1187,In_878,In_0);
nor U1188 (N_1188,In_208,In_249);
nor U1189 (N_1189,In_448,In_409);
nor U1190 (N_1190,In_623,In_185);
nand U1191 (N_1191,In_731,In_931);
or U1192 (N_1192,In_491,In_550);
or U1193 (N_1193,In_491,In_783);
and U1194 (N_1194,In_644,In_933);
nand U1195 (N_1195,In_141,In_666);
or U1196 (N_1196,In_575,In_430);
nor U1197 (N_1197,In_858,In_956);
or U1198 (N_1198,In_727,In_901);
and U1199 (N_1199,In_81,In_532);
nand U1200 (N_1200,In_600,In_771);
nor U1201 (N_1201,In_536,In_69);
and U1202 (N_1202,In_83,In_810);
and U1203 (N_1203,In_505,In_629);
and U1204 (N_1204,In_104,In_811);
nor U1205 (N_1205,In_505,In_831);
and U1206 (N_1206,In_11,In_91);
and U1207 (N_1207,In_766,In_841);
or U1208 (N_1208,In_844,In_37);
nor U1209 (N_1209,In_314,In_462);
and U1210 (N_1210,In_964,In_999);
or U1211 (N_1211,In_838,In_81);
and U1212 (N_1212,In_949,In_742);
and U1213 (N_1213,In_480,In_706);
and U1214 (N_1214,In_609,In_14);
nor U1215 (N_1215,In_451,In_739);
and U1216 (N_1216,In_991,In_480);
and U1217 (N_1217,In_126,In_640);
nor U1218 (N_1218,In_77,In_446);
and U1219 (N_1219,In_786,In_964);
nand U1220 (N_1220,In_275,In_46);
nand U1221 (N_1221,In_294,In_568);
nor U1222 (N_1222,In_749,In_407);
or U1223 (N_1223,In_183,In_345);
nor U1224 (N_1224,In_834,In_819);
or U1225 (N_1225,In_693,In_708);
nor U1226 (N_1226,In_635,In_465);
or U1227 (N_1227,In_590,In_249);
and U1228 (N_1228,In_983,In_835);
and U1229 (N_1229,In_856,In_477);
and U1230 (N_1230,In_722,In_581);
nor U1231 (N_1231,In_961,In_43);
and U1232 (N_1232,In_595,In_505);
and U1233 (N_1233,In_351,In_745);
or U1234 (N_1234,In_577,In_298);
and U1235 (N_1235,In_554,In_344);
and U1236 (N_1236,In_464,In_96);
or U1237 (N_1237,In_847,In_958);
and U1238 (N_1238,In_415,In_458);
nand U1239 (N_1239,In_496,In_334);
and U1240 (N_1240,In_3,In_459);
or U1241 (N_1241,In_519,In_342);
or U1242 (N_1242,In_1,In_856);
or U1243 (N_1243,In_863,In_504);
nor U1244 (N_1244,In_491,In_228);
nor U1245 (N_1245,In_59,In_968);
nor U1246 (N_1246,In_168,In_715);
and U1247 (N_1247,In_1,In_488);
nor U1248 (N_1248,In_502,In_568);
nand U1249 (N_1249,In_449,In_815);
or U1250 (N_1250,In_912,In_738);
nor U1251 (N_1251,In_228,In_122);
or U1252 (N_1252,In_14,In_877);
nor U1253 (N_1253,In_379,In_600);
and U1254 (N_1254,In_750,In_273);
nor U1255 (N_1255,In_886,In_149);
or U1256 (N_1256,In_821,In_213);
or U1257 (N_1257,In_394,In_217);
nor U1258 (N_1258,In_284,In_292);
nand U1259 (N_1259,In_634,In_584);
or U1260 (N_1260,In_788,In_236);
or U1261 (N_1261,In_350,In_486);
or U1262 (N_1262,In_132,In_224);
nand U1263 (N_1263,In_467,In_752);
and U1264 (N_1264,In_935,In_821);
or U1265 (N_1265,In_727,In_614);
and U1266 (N_1266,In_565,In_44);
nand U1267 (N_1267,In_72,In_222);
nand U1268 (N_1268,In_581,In_16);
nand U1269 (N_1269,In_611,In_619);
and U1270 (N_1270,In_255,In_894);
nand U1271 (N_1271,In_813,In_349);
and U1272 (N_1272,In_91,In_219);
xor U1273 (N_1273,In_295,In_471);
and U1274 (N_1274,In_392,In_272);
nor U1275 (N_1275,In_512,In_848);
nand U1276 (N_1276,In_558,In_940);
nand U1277 (N_1277,In_838,In_153);
and U1278 (N_1278,In_929,In_45);
or U1279 (N_1279,In_554,In_320);
nand U1280 (N_1280,In_325,In_543);
and U1281 (N_1281,In_541,In_954);
nand U1282 (N_1282,In_61,In_607);
or U1283 (N_1283,In_684,In_200);
and U1284 (N_1284,In_56,In_155);
nand U1285 (N_1285,In_130,In_914);
and U1286 (N_1286,In_698,In_727);
or U1287 (N_1287,In_620,In_181);
and U1288 (N_1288,In_514,In_859);
nor U1289 (N_1289,In_662,In_645);
and U1290 (N_1290,In_708,In_824);
and U1291 (N_1291,In_482,In_522);
nor U1292 (N_1292,In_154,In_222);
nor U1293 (N_1293,In_100,In_336);
and U1294 (N_1294,In_30,In_858);
or U1295 (N_1295,In_120,In_874);
or U1296 (N_1296,In_987,In_72);
nand U1297 (N_1297,In_166,In_359);
nand U1298 (N_1298,In_240,In_488);
and U1299 (N_1299,In_218,In_264);
nor U1300 (N_1300,In_251,In_97);
and U1301 (N_1301,In_338,In_614);
nand U1302 (N_1302,In_654,In_87);
nand U1303 (N_1303,In_915,In_301);
and U1304 (N_1304,In_193,In_845);
nor U1305 (N_1305,In_166,In_90);
and U1306 (N_1306,In_794,In_359);
nor U1307 (N_1307,In_946,In_719);
or U1308 (N_1308,In_268,In_766);
and U1309 (N_1309,In_992,In_82);
nor U1310 (N_1310,In_760,In_468);
or U1311 (N_1311,In_766,In_326);
or U1312 (N_1312,In_805,In_353);
and U1313 (N_1313,In_738,In_335);
nor U1314 (N_1314,In_298,In_23);
nand U1315 (N_1315,In_871,In_129);
and U1316 (N_1316,In_868,In_872);
or U1317 (N_1317,In_739,In_407);
nor U1318 (N_1318,In_896,In_139);
nor U1319 (N_1319,In_689,In_769);
nor U1320 (N_1320,In_312,In_748);
or U1321 (N_1321,In_257,In_888);
nor U1322 (N_1322,In_352,In_5);
and U1323 (N_1323,In_442,In_678);
and U1324 (N_1324,In_645,In_53);
xor U1325 (N_1325,In_149,In_84);
or U1326 (N_1326,In_758,In_385);
nor U1327 (N_1327,In_86,In_440);
or U1328 (N_1328,In_384,In_925);
nor U1329 (N_1329,In_180,In_90);
and U1330 (N_1330,In_988,In_130);
and U1331 (N_1331,In_355,In_802);
nand U1332 (N_1332,In_351,In_774);
and U1333 (N_1333,In_581,In_741);
nor U1334 (N_1334,In_690,In_179);
and U1335 (N_1335,In_906,In_696);
and U1336 (N_1336,In_587,In_708);
nand U1337 (N_1337,In_573,In_105);
nand U1338 (N_1338,In_277,In_30);
and U1339 (N_1339,In_996,In_876);
or U1340 (N_1340,In_746,In_542);
nand U1341 (N_1341,In_853,In_165);
or U1342 (N_1342,In_575,In_599);
nand U1343 (N_1343,In_33,In_271);
and U1344 (N_1344,In_41,In_734);
or U1345 (N_1345,In_798,In_8);
nand U1346 (N_1346,In_847,In_325);
or U1347 (N_1347,In_181,In_351);
nor U1348 (N_1348,In_827,In_477);
nand U1349 (N_1349,In_32,In_596);
nand U1350 (N_1350,In_970,In_747);
or U1351 (N_1351,In_507,In_401);
nand U1352 (N_1352,In_730,In_47);
nor U1353 (N_1353,In_657,In_427);
or U1354 (N_1354,In_691,In_389);
nor U1355 (N_1355,In_507,In_392);
nor U1356 (N_1356,In_530,In_638);
nand U1357 (N_1357,In_348,In_609);
nor U1358 (N_1358,In_444,In_548);
xor U1359 (N_1359,In_299,In_975);
and U1360 (N_1360,In_404,In_952);
nand U1361 (N_1361,In_248,In_3);
or U1362 (N_1362,In_125,In_310);
and U1363 (N_1363,In_608,In_178);
and U1364 (N_1364,In_613,In_954);
xor U1365 (N_1365,In_974,In_407);
nor U1366 (N_1366,In_887,In_805);
nand U1367 (N_1367,In_857,In_510);
or U1368 (N_1368,In_729,In_9);
and U1369 (N_1369,In_730,In_718);
nor U1370 (N_1370,In_796,In_926);
or U1371 (N_1371,In_498,In_248);
xor U1372 (N_1372,In_308,In_919);
nand U1373 (N_1373,In_785,In_598);
nand U1374 (N_1374,In_537,In_662);
and U1375 (N_1375,In_56,In_608);
nor U1376 (N_1376,In_468,In_678);
nand U1377 (N_1377,In_120,In_261);
nor U1378 (N_1378,In_419,In_132);
or U1379 (N_1379,In_482,In_91);
nor U1380 (N_1380,In_136,In_729);
nor U1381 (N_1381,In_275,In_748);
or U1382 (N_1382,In_927,In_938);
or U1383 (N_1383,In_620,In_728);
and U1384 (N_1384,In_579,In_483);
nor U1385 (N_1385,In_841,In_644);
nand U1386 (N_1386,In_867,In_479);
and U1387 (N_1387,In_214,In_223);
or U1388 (N_1388,In_887,In_193);
or U1389 (N_1389,In_942,In_317);
or U1390 (N_1390,In_607,In_69);
and U1391 (N_1391,In_773,In_742);
or U1392 (N_1392,In_282,In_223);
nand U1393 (N_1393,In_836,In_60);
and U1394 (N_1394,In_851,In_867);
nand U1395 (N_1395,In_446,In_334);
or U1396 (N_1396,In_329,In_332);
xor U1397 (N_1397,In_384,In_559);
and U1398 (N_1398,In_268,In_134);
nor U1399 (N_1399,In_591,In_78);
nand U1400 (N_1400,In_803,In_316);
nor U1401 (N_1401,In_484,In_432);
and U1402 (N_1402,In_219,In_393);
nor U1403 (N_1403,In_154,In_93);
or U1404 (N_1404,In_292,In_141);
and U1405 (N_1405,In_947,In_977);
or U1406 (N_1406,In_589,In_637);
or U1407 (N_1407,In_229,In_833);
nand U1408 (N_1408,In_247,In_216);
nor U1409 (N_1409,In_786,In_507);
nand U1410 (N_1410,In_31,In_127);
nor U1411 (N_1411,In_852,In_906);
and U1412 (N_1412,In_102,In_966);
or U1413 (N_1413,In_852,In_933);
nor U1414 (N_1414,In_838,In_640);
and U1415 (N_1415,In_657,In_753);
and U1416 (N_1416,In_826,In_439);
or U1417 (N_1417,In_500,In_279);
or U1418 (N_1418,In_726,In_209);
or U1419 (N_1419,In_451,In_845);
nand U1420 (N_1420,In_513,In_835);
and U1421 (N_1421,In_849,In_821);
and U1422 (N_1422,In_395,In_341);
nand U1423 (N_1423,In_235,In_427);
nand U1424 (N_1424,In_73,In_293);
nand U1425 (N_1425,In_436,In_719);
or U1426 (N_1426,In_305,In_323);
nor U1427 (N_1427,In_152,In_79);
nand U1428 (N_1428,In_221,In_284);
and U1429 (N_1429,In_413,In_84);
or U1430 (N_1430,In_791,In_915);
and U1431 (N_1431,In_707,In_671);
nand U1432 (N_1432,In_181,In_234);
and U1433 (N_1433,In_568,In_74);
nor U1434 (N_1434,In_905,In_344);
nor U1435 (N_1435,In_680,In_675);
or U1436 (N_1436,In_719,In_452);
or U1437 (N_1437,In_548,In_426);
nor U1438 (N_1438,In_22,In_313);
and U1439 (N_1439,In_445,In_529);
nand U1440 (N_1440,In_987,In_15);
or U1441 (N_1441,In_198,In_473);
and U1442 (N_1442,In_687,In_563);
nand U1443 (N_1443,In_750,In_161);
nand U1444 (N_1444,In_457,In_621);
and U1445 (N_1445,In_419,In_440);
and U1446 (N_1446,In_898,In_606);
or U1447 (N_1447,In_467,In_966);
or U1448 (N_1448,In_252,In_362);
or U1449 (N_1449,In_578,In_36);
or U1450 (N_1450,In_310,In_200);
or U1451 (N_1451,In_109,In_839);
or U1452 (N_1452,In_378,In_873);
nand U1453 (N_1453,In_807,In_490);
or U1454 (N_1454,In_57,In_329);
nand U1455 (N_1455,In_179,In_450);
and U1456 (N_1456,In_476,In_386);
and U1457 (N_1457,In_768,In_744);
nand U1458 (N_1458,In_956,In_20);
nand U1459 (N_1459,In_213,In_728);
nand U1460 (N_1460,In_884,In_153);
nor U1461 (N_1461,In_97,In_150);
or U1462 (N_1462,In_664,In_284);
and U1463 (N_1463,In_59,In_335);
nand U1464 (N_1464,In_615,In_813);
nor U1465 (N_1465,In_104,In_837);
and U1466 (N_1466,In_64,In_809);
and U1467 (N_1467,In_173,In_877);
nand U1468 (N_1468,In_499,In_31);
nor U1469 (N_1469,In_923,In_244);
nor U1470 (N_1470,In_711,In_725);
nor U1471 (N_1471,In_123,In_939);
and U1472 (N_1472,In_586,In_748);
nand U1473 (N_1473,In_994,In_534);
nor U1474 (N_1474,In_558,In_829);
and U1475 (N_1475,In_801,In_643);
nand U1476 (N_1476,In_935,In_266);
or U1477 (N_1477,In_179,In_982);
or U1478 (N_1478,In_948,In_620);
nor U1479 (N_1479,In_17,In_816);
and U1480 (N_1480,In_131,In_177);
or U1481 (N_1481,In_230,In_562);
nor U1482 (N_1482,In_517,In_686);
nand U1483 (N_1483,In_532,In_259);
and U1484 (N_1484,In_271,In_632);
nor U1485 (N_1485,In_85,In_668);
or U1486 (N_1486,In_153,In_358);
nand U1487 (N_1487,In_984,In_356);
and U1488 (N_1488,In_433,In_989);
nor U1489 (N_1489,In_949,In_574);
xnor U1490 (N_1490,In_300,In_140);
nand U1491 (N_1491,In_668,In_369);
and U1492 (N_1492,In_872,In_826);
nand U1493 (N_1493,In_698,In_207);
nor U1494 (N_1494,In_147,In_953);
nand U1495 (N_1495,In_717,In_446);
or U1496 (N_1496,In_467,In_332);
or U1497 (N_1497,In_968,In_214);
or U1498 (N_1498,In_797,In_547);
nand U1499 (N_1499,In_259,In_609);
and U1500 (N_1500,In_776,In_667);
or U1501 (N_1501,In_666,In_354);
nand U1502 (N_1502,In_591,In_683);
or U1503 (N_1503,In_876,In_597);
and U1504 (N_1504,In_609,In_720);
nand U1505 (N_1505,In_710,In_28);
nand U1506 (N_1506,In_362,In_146);
and U1507 (N_1507,In_246,In_581);
nor U1508 (N_1508,In_386,In_990);
or U1509 (N_1509,In_977,In_122);
nand U1510 (N_1510,In_16,In_327);
nor U1511 (N_1511,In_325,In_134);
nor U1512 (N_1512,In_375,In_957);
and U1513 (N_1513,In_863,In_346);
nand U1514 (N_1514,In_106,In_105);
nor U1515 (N_1515,In_59,In_579);
nand U1516 (N_1516,In_248,In_41);
and U1517 (N_1517,In_677,In_238);
nor U1518 (N_1518,In_168,In_562);
nor U1519 (N_1519,In_850,In_120);
nand U1520 (N_1520,In_180,In_273);
nor U1521 (N_1521,In_451,In_375);
or U1522 (N_1522,In_554,In_111);
or U1523 (N_1523,In_594,In_623);
and U1524 (N_1524,In_165,In_399);
nor U1525 (N_1525,In_242,In_531);
or U1526 (N_1526,In_508,In_454);
nand U1527 (N_1527,In_656,In_757);
nand U1528 (N_1528,In_774,In_297);
or U1529 (N_1529,In_417,In_624);
nand U1530 (N_1530,In_417,In_117);
and U1531 (N_1531,In_25,In_222);
nor U1532 (N_1532,In_741,In_575);
or U1533 (N_1533,In_325,In_440);
nand U1534 (N_1534,In_391,In_988);
nand U1535 (N_1535,In_241,In_217);
or U1536 (N_1536,In_118,In_7);
or U1537 (N_1537,In_951,In_985);
or U1538 (N_1538,In_418,In_453);
and U1539 (N_1539,In_973,In_875);
nor U1540 (N_1540,In_744,In_131);
nor U1541 (N_1541,In_738,In_258);
or U1542 (N_1542,In_989,In_886);
nand U1543 (N_1543,In_227,In_369);
and U1544 (N_1544,In_489,In_851);
and U1545 (N_1545,In_202,In_98);
or U1546 (N_1546,In_853,In_558);
nand U1547 (N_1547,In_278,In_296);
nor U1548 (N_1548,In_211,In_698);
or U1549 (N_1549,In_294,In_306);
and U1550 (N_1550,In_622,In_362);
nand U1551 (N_1551,In_795,In_850);
nor U1552 (N_1552,In_386,In_621);
and U1553 (N_1553,In_631,In_497);
nor U1554 (N_1554,In_333,In_525);
nand U1555 (N_1555,In_185,In_214);
nor U1556 (N_1556,In_259,In_729);
nor U1557 (N_1557,In_217,In_786);
nand U1558 (N_1558,In_772,In_683);
or U1559 (N_1559,In_469,In_534);
nand U1560 (N_1560,In_38,In_188);
nor U1561 (N_1561,In_674,In_287);
and U1562 (N_1562,In_188,In_39);
xor U1563 (N_1563,In_645,In_66);
or U1564 (N_1564,In_812,In_78);
and U1565 (N_1565,In_611,In_846);
or U1566 (N_1566,In_482,In_924);
or U1567 (N_1567,In_755,In_150);
and U1568 (N_1568,In_1,In_564);
or U1569 (N_1569,In_11,In_281);
nor U1570 (N_1570,In_388,In_280);
or U1571 (N_1571,In_617,In_576);
and U1572 (N_1572,In_110,In_527);
nand U1573 (N_1573,In_514,In_277);
nand U1574 (N_1574,In_235,In_268);
and U1575 (N_1575,In_550,In_316);
nand U1576 (N_1576,In_431,In_329);
or U1577 (N_1577,In_677,In_518);
and U1578 (N_1578,In_175,In_461);
and U1579 (N_1579,In_441,In_542);
or U1580 (N_1580,In_452,In_191);
nor U1581 (N_1581,In_304,In_513);
or U1582 (N_1582,In_35,In_947);
and U1583 (N_1583,In_525,In_171);
nand U1584 (N_1584,In_327,In_642);
nand U1585 (N_1585,In_353,In_623);
or U1586 (N_1586,In_638,In_368);
nor U1587 (N_1587,In_507,In_813);
and U1588 (N_1588,In_877,In_790);
and U1589 (N_1589,In_767,In_516);
and U1590 (N_1590,In_968,In_645);
nor U1591 (N_1591,In_482,In_395);
nor U1592 (N_1592,In_868,In_489);
or U1593 (N_1593,In_940,In_995);
and U1594 (N_1594,In_960,In_460);
or U1595 (N_1595,In_853,In_968);
and U1596 (N_1596,In_364,In_161);
nor U1597 (N_1597,In_153,In_208);
nor U1598 (N_1598,In_507,In_795);
or U1599 (N_1599,In_675,In_564);
or U1600 (N_1600,In_974,In_591);
nand U1601 (N_1601,In_365,In_287);
nor U1602 (N_1602,In_358,In_567);
nand U1603 (N_1603,In_132,In_958);
or U1604 (N_1604,In_305,In_755);
nand U1605 (N_1605,In_80,In_311);
nand U1606 (N_1606,In_138,In_468);
nor U1607 (N_1607,In_559,In_754);
nor U1608 (N_1608,In_708,In_705);
nand U1609 (N_1609,In_433,In_184);
and U1610 (N_1610,In_109,In_48);
and U1611 (N_1611,In_361,In_557);
nor U1612 (N_1612,In_308,In_731);
and U1613 (N_1613,In_582,In_273);
and U1614 (N_1614,In_760,In_810);
nand U1615 (N_1615,In_821,In_685);
or U1616 (N_1616,In_356,In_147);
or U1617 (N_1617,In_337,In_669);
nor U1618 (N_1618,In_333,In_458);
or U1619 (N_1619,In_640,In_184);
or U1620 (N_1620,In_247,In_660);
or U1621 (N_1621,In_194,In_15);
nor U1622 (N_1622,In_7,In_835);
or U1623 (N_1623,In_13,In_456);
or U1624 (N_1624,In_632,In_200);
xnor U1625 (N_1625,In_442,In_625);
xnor U1626 (N_1626,In_560,In_736);
nand U1627 (N_1627,In_384,In_136);
or U1628 (N_1628,In_202,In_738);
nor U1629 (N_1629,In_183,In_726);
or U1630 (N_1630,In_208,In_928);
nor U1631 (N_1631,In_770,In_666);
nand U1632 (N_1632,In_335,In_264);
or U1633 (N_1633,In_982,In_142);
or U1634 (N_1634,In_169,In_352);
nand U1635 (N_1635,In_38,In_964);
nor U1636 (N_1636,In_851,In_114);
or U1637 (N_1637,In_703,In_89);
nor U1638 (N_1638,In_148,In_782);
nor U1639 (N_1639,In_813,In_520);
nor U1640 (N_1640,In_93,In_983);
or U1641 (N_1641,In_467,In_555);
or U1642 (N_1642,In_543,In_638);
or U1643 (N_1643,In_200,In_581);
nor U1644 (N_1644,In_507,In_498);
nand U1645 (N_1645,In_13,In_740);
nor U1646 (N_1646,In_368,In_5);
nor U1647 (N_1647,In_78,In_636);
nor U1648 (N_1648,In_193,In_648);
nand U1649 (N_1649,In_560,In_503);
nor U1650 (N_1650,In_755,In_34);
or U1651 (N_1651,In_701,In_578);
nor U1652 (N_1652,In_907,In_418);
or U1653 (N_1653,In_435,In_77);
and U1654 (N_1654,In_616,In_736);
and U1655 (N_1655,In_632,In_790);
and U1656 (N_1656,In_547,In_952);
nor U1657 (N_1657,In_467,In_255);
nor U1658 (N_1658,In_410,In_420);
and U1659 (N_1659,In_369,In_25);
nor U1660 (N_1660,In_575,In_821);
and U1661 (N_1661,In_461,In_736);
nor U1662 (N_1662,In_861,In_220);
and U1663 (N_1663,In_849,In_535);
and U1664 (N_1664,In_237,In_252);
and U1665 (N_1665,In_408,In_89);
nand U1666 (N_1666,In_752,In_298);
nand U1667 (N_1667,In_332,In_777);
or U1668 (N_1668,In_751,In_124);
nor U1669 (N_1669,In_739,In_361);
and U1670 (N_1670,In_732,In_566);
nand U1671 (N_1671,In_225,In_302);
or U1672 (N_1672,In_292,In_783);
and U1673 (N_1673,In_322,In_448);
and U1674 (N_1674,In_96,In_576);
nand U1675 (N_1675,In_206,In_350);
or U1676 (N_1676,In_365,In_718);
nand U1677 (N_1677,In_928,In_422);
and U1678 (N_1678,In_957,In_371);
nand U1679 (N_1679,In_831,In_916);
xnor U1680 (N_1680,In_510,In_163);
nor U1681 (N_1681,In_937,In_434);
or U1682 (N_1682,In_111,In_774);
nor U1683 (N_1683,In_115,In_460);
nand U1684 (N_1684,In_60,In_37);
and U1685 (N_1685,In_304,In_702);
nor U1686 (N_1686,In_415,In_950);
nor U1687 (N_1687,In_396,In_474);
or U1688 (N_1688,In_918,In_124);
and U1689 (N_1689,In_304,In_608);
nor U1690 (N_1690,In_282,In_641);
or U1691 (N_1691,In_162,In_104);
and U1692 (N_1692,In_755,In_105);
nand U1693 (N_1693,In_749,In_722);
or U1694 (N_1694,In_886,In_259);
nor U1695 (N_1695,In_458,In_459);
nand U1696 (N_1696,In_489,In_39);
or U1697 (N_1697,In_7,In_291);
and U1698 (N_1698,In_72,In_329);
nor U1699 (N_1699,In_477,In_780);
nor U1700 (N_1700,In_527,In_485);
nor U1701 (N_1701,In_408,In_731);
or U1702 (N_1702,In_119,In_631);
or U1703 (N_1703,In_594,In_251);
or U1704 (N_1704,In_623,In_416);
or U1705 (N_1705,In_526,In_569);
nand U1706 (N_1706,In_218,In_827);
nor U1707 (N_1707,In_522,In_737);
and U1708 (N_1708,In_312,In_715);
nor U1709 (N_1709,In_838,In_537);
nand U1710 (N_1710,In_632,In_510);
nand U1711 (N_1711,In_977,In_454);
nor U1712 (N_1712,In_816,In_813);
nor U1713 (N_1713,In_897,In_864);
nor U1714 (N_1714,In_913,In_590);
or U1715 (N_1715,In_204,In_28);
nor U1716 (N_1716,In_602,In_313);
or U1717 (N_1717,In_819,In_912);
nand U1718 (N_1718,In_196,In_582);
and U1719 (N_1719,In_900,In_325);
nor U1720 (N_1720,In_696,In_868);
or U1721 (N_1721,In_498,In_930);
or U1722 (N_1722,In_140,In_564);
or U1723 (N_1723,In_251,In_605);
and U1724 (N_1724,In_557,In_114);
or U1725 (N_1725,In_725,In_833);
or U1726 (N_1726,In_651,In_875);
nand U1727 (N_1727,In_738,In_67);
or U1728 (N_1728,In_958,In_314);
and U1729 (N_1729,In_519,In_988);
nor U1730 (N_1730,In_872,In_163);
or U1731 (N_1731,In_542,In_29);
or U1732 (N_1732,In_292,In_754);
or U1733 (N_1733,In_171,In_105);
and U1734 (N_1734,In_936,In_942);
nor U1735 (N_1735,In_864,In_22);
or U1736 (N_1736,In_429,In_519);
xor U1737 (N_1737,In_328,In_587);
and U1738 (N_1738,In_684,In_581);
or U1739 (N_1739,In_456,In_34);
nor U1740 (N_1740,In_99,In_815);
nor U1741 (N_1741,In_403,In_228);
nand U1742 (N_1742,In_44,In_961);
or U1743 (N_1743,In_434,In_502);
and U1744 (N_1744,In_322,In_108);
nand U1745 (N_1745,In_496,In_502);
or U1746 (N_1746,In_118,In_589);
and U1747 (N_1747,In_805,In_541);
nand U1748 (N_1748,In_510,In_354);
nand U1749 (N_1749,In_496,In_467);
nor U1750 (N_1750,In_360,In_674);
nand U1751 (N_1751,In_580,In_867);
nor U1752 (N_1752,In_318,In_955);
or U1753 (N_1753,In_924,In_867);
or U1754 (N_1754,In_386,In_951);
nand U1755 (N_1755,In_662,In_570);
nand U1756 (N_1756,In_180,In_219);
nand U1757 (N_1757,In_561,In_321);
nor U1758 (N_1758,In_93,In_882);
or U1759 (N_1759,In_617,In_653);
and U1760 (N_1760,In_898,In_585);
or U1761 (N_1761,In_573,In_707);
nor U1762 (N_1762,In_118,In_743);
nand U1763 (N_1763,In_580,In_804);
and U1764 (N_1764,In_164,In_686);
or U1765 (N_1765,In_367,In_161);
nand U1766 (N_1766,In_727,In_560);
or U1767 (N_1767,In_505,In_818);
or U1768 (N_1768,In_347,In_346);
and U1769 (N_1769,In_991,In_191);
or U1770 (N_1770,In_342,In_444);
nor U1771 (N_1771,In_454,In_845);
or U1772 (N_1772,In_272,In_742);
or U1773 (N_1773,In_651,In_530);
nand U1774 (N_1774,In_786,In_284);
xor U1775 (N_1775,In_781,In_648);
and U1776 (N_1776,In_652,In_77);
nand U1777 (N_1777,In_132,In_727);
and U1778 (N_1778,In_271,In_972);
or U1779 (N_1779,In_721,In_959);
nand U1780 (N_1780,In_498,In_712);
nor U1781 (N_1781,In_701,In_71);
nand U1782 (N_1782,In_820,In_210);
nand U1783 (N_1783,In_519,In_129);
nor U1784 (N_1784,In_393,In_869);
or U1785 (N_1785,In_118,In_328);
nor U1786 (N_1786,In_170,In_72);
nor U1787 (N_1787,In_944,In_430);
nor U1788 (N_1788,In_225,In_973);
or U1789 (N_1789,In_872,In_389);
nand U1790 (N_1790,In_980,In_378);
and U1791 (N_1791,In_979,In_362);
and U1792 (N_1792,In_816,In_444);
nor U1793 (N_1793,In_533,In_135);
and U1794 (N_1794,In_449,In_909);
nor U1795 (N_1795,In_910,In_455);
and U1796 (N_1796,In_494,In_329);
nor U1797 (N_1797,In_53,In_566);
or U1798 (N_1798,In_255,In_685);
or U1799 (N_1799,In_213,In_552);
nand U1800 (N_1800,In_722,In_627);
nor U1801 (N_1801,In_750,In_38);
nor U1802 (N_1802,In_352,In_172);
nand U1803 (N_1803,In_304,In_897);
or U1804 (N_1804,In_326,In_480);
nor U1805 (N_1805,In_844,In_820);
nand U1806 (N_1806,In_491,In_792);
nor U1807 (N_1807,In_521,In_144);
or U1808 (N_1808,In_97,In_856);
nand U1809 (N_1809,In_284,In_709);
nand U1810 (N_1810,In_849,In_284);
nor U1811 (N_1811,In_44,In_753);
nand U1812 (N_1812,In_90,In_649);
nor U1813 (N_1813,In_813,In_784);
nand U1814 (N_1814,In_174,In_717);
and U1815 (N_1815,In_634,In_985);
or U1816 (N_1816,In_223,In_982);
and U1817 (N_1817,In_466,In_842);
nand U1818 (N_1818,In_302,In_6);
nand U1819 (N_1819,In_171,In_925);
and U1820 (N_1820,In_159,In_309);
xor U1821 (N_1821,In_343,In_447);
nand U1822 (N_1822,In_603,In_871);
nand U1823 (N_1823,In_348,In_459);
or U1824 (N_1824,In_822,In_99);
or U1825 (N_1825,In_872,In_715);
or U1826 (N_1826,In_408,In_987);
nor U1827 (N_1827,In_342,In_184);
nand U1828 (N_1828,In_467,In_876);
nor U1829 (N_1829,In_469,In_658);
or U1830 (N_1830,In_53,In_448);
or U1831 (N_1831,In_603,In_105);
or U1832 (N_1832,In_954,In_293);
nand U1833 (N_1833,In_179,In_603);
nor U1834 (N_1834,In_204,In_664);
and U1835 (N_1835,In_71,In_405);
or U1836 (N_1836,In_29,In_943);
nor U1837 (N_1837,In_272,In_193);
and U1838 (N_1838,In_332,In_873);
nor U1839 (N_1839,In_451,In_231);
and U1840 (N_1840,In_442,In_305);
or U1841 (N_1841,In_197,In_52);
or U1842 (N_1842,In_533,In_626);
and U1843 (N_1843,In_398,In_649);
or U1844 (N_1844,In_116,In_961);
nand U1845 (N_1845,In_582,In_553);
nand U1846 (N_1846,In_924,In_622);
or U1847 (N_1847,In_227,In_133);
or U1848 (N_1848,In_662,In_700);
nor U1849 (N_1849,In_807,In_983);
or U1850 (N_1850,In_959,In_882);
or U1851 (N_1851,In_677,In_678);
or U1852 (N_1852,In_983,In_570);
nand U1853 (N_1853,In_4,In_33);
nand U1854 (N_1854,In_156,In_46);
or U1855 (N_1855,In_634,In_465);
nor U1856 (N_1856,In_477,In_115);
nor U1857 (N_1857,In_998,In_615);
and U1858 (N_1858,In_384,In_818);
and U1859 (N_1859,In_715,In_874);
or U1860 (N_1860,In_743,In_261);
and U1861 (N_1861,In_884,In_730);
and U1862 (N_1862,In_13,In_517);
and U1863 (N_1863,In_973,In_650);
and U1864 (N_1864,In_65,In_73);
nor U1865 (N_1865,In_112,In_599);
or U1866 (N_1866,In_123,In_943);
nor U1867 (N_1867,In_59,In_21);
nor U1868 (N_1868,In_579,In_81);
or U1869 (N_1869,In_454,In_185);
nand U1870 (N_1870,In_280,In_673);
nand U1871 (N_1871,In_108,In_173);
and U1872 (N_1872,In_356,In_404);
nor U1873 (N_1873,In_336,In_114);
and U1874 (N_1874,In_676,In_611);
nand U1875 (N_1875,In_321,In_505);
and U1876 (N_1876,In_524,In_558);
and U1877 (N_1877,In_358,In_840);
nand U1878 (N_1878,In_523,In_512);
and U1879 (N_1879,In_584,In_312);
or U1880 (N_1880,In_626,In_805);
nor U1881 (N_1881,In_662,In_692);
and U1882 (N_1882,In_205,In_598);
and U1883 (N_1883,In_318,In_393);
and U1884 (N_1884,In_234,In_737);
nor U1885 (N_1885,In_677,In_233);
and U1886 (N_1886,In_703,In_981);
or U1887 (N_1887,In_528,In_912);
nand U1888 (N_1888,In_36,In_794);
nand U1889 (N_1889,In_465,In_477);
and U1890 (N_1890,In_872,In_68);
and U1891 (N_1891,In_773,In_61);
nor U1892 (N_1892,In_446,In_563);
or U1893 (N_1893,In_554,In_275);
or U1894 (N_1894,In_721,In_373);
nor U1895 (N_1895,In_755,In_939);
nand U1896 (N_1896,In_706,In_283);
or U1897 (N_1897,In_565,In_910);
nand U1898 (N_1898,In_290,In_384);
or U1899 (N_1899,In_154,In_888);
nor U1900 (N_1900,In_80,In_302);
and U1901 (N_1901,In_65,In_710);
nor U1902 (N_1902,In_985,In_706);
or U1903 (N_1903,In_536,In_77);
nor U1904 (N_1904,In_64,In_356);
and U1905 (N_1905,In_731,In_875);
nor U1906 (N_1906,In_942,In_930);
nand U1907 (N_1907,In_938,In_322);
nor U1908 (N_1908,In_223,In_896);
and U1909 (N_1909,In_143,In_250);
and U1910 (N_1910,In_514,In_919);
and U1911 (N_1911,In_656,In_721);
and U1912 (N_1912,In_788,In_655);
and U1913 (N_1913,In_975,In_735);
or U1914 (N_1914,In_777,In_108);
or U1915 (N_1915,In_769,In_699);
and U1916 (N_1916,In_916,In_418);
nand U1917 (N_1917,In_729,In_535);
nand U1918 (N_1918,In_259,In_834);
and U1919 (N_1919,In_437,In_847);
nor U1920 (N_1920,In_770,In_998);
nor U1921 (N_1921,In_448,In_917);
nand U1922 (N_1922,In_168,In_438);
nand U1923 (N_1923,In_22,In_162);
and U1924 (N_1924,In_339,In_587);
or U1925 (N_1925,In_864,In_958);
and U1926 (N_1926,In_753,In_603);
and U1927 (N_1927,In_995,In_678);
or U1928 (N_1928,In_772,In_578);
and U1929 (N_1929,In_449,In_765);
or U1930 (N_1930,In_833,In_572);
xnor U1931 (N_1931,In_687,In_826);
or U1932 (N_1932,In_875,In_980);
and U1933 (N_1933,In_953,In_203);
and U1934 (N_1934,In_157,In_345);
and U1935 (N_1935,In_347,In_756);
and U1936 (N_1936,In_935,In_702);
and U1937 (N_1937,In_552,In_171);
or U1938 (N_1938,In_208,In_453);
nand U1939 (N_1939,In_563,In_606);
or U1940 (N_1940,In_481,In_665);
or U1941 (N_1941,In_747,In_69);
or U1942 (N_1942,In_993,In_877);
nor U1943 (N_1943,In_890,In_857);
nand U1944 (N_1944,In_496,In_726);
and U1945 (N_1945,In_631,In_303);
nand U1946 (N_1946,In_699,In_196);
or U1947 (N_1947,In_450,In_887);
nand U1948 (N_1948,In_389,In_631);
or U1949 (N_1949,In_92,In_94);
nand U1950 (N_1950,In_914,In_200);
or U1951 (N_1951,In_315,In_206);
and U1952 (N_1952,In_323,In_950);
and U1953 (N_1953,In_469,In_432);
nand U1954 (N_1954,In_18,In_799);
nor U1955 (N_1955,In_486,In_710);
nor U1956 (N_1956,In_719,In_853);
nand U1957 (N_1957,In_626,In_45);
or U1958 (N_1958,In_224,In_191);
xnor U1959 (N_1959,In_128,In_68);
or U1960 (N_1960,In_207,In_722);
nand U1961 (N_1961,In_54,In_830);
nor U1962 (N_1962,In_354,In_739);
nand U1963 (N_1963,In_53,In_280);
or U1964 (N_1964,In_426,In_767);
nor U1965 (N_1965,In_425,In_245);
nor U1966 (N_1966,In_423,In_431);
nand U1967 (N_1967,In_332,In_244);
and U1968 (N_1968,In_23,In_690);
and U1969 (N_1969,In_708,In_401);
nor U1970 (N_1970,In_398,In_348);
or U1971 (N_1971,In_798,In_245);
nand U1972 (N_1972,In_453,In_522);
or U1973 (N_1973,In_402,In_137);
nor U1974 (N_1974,In_899,In_800);
nor U1975 (N_1975,In_424,In_761);
nand U1976 (N_1976,In_120,In_255);
or U1977 (N_1977,In_102,In_300);
nand U1978 (N_1978,In_303,In_830);
or U1979 (N_1979,In_564,In_747);
and U1980 (N_1980,In_807,In_399);
nor U1981 (N_1981,In_983,In_761);
and U1982 (N_1982,In_154,In_91);
nand U1983 (N_1983,In_524,In_815);
and U1984 (N_1984,In_199,In_98);
nor U1985 (N_1985,In_199,In_337);
or U1986 (N_1986,In_193,In_464);
or U1987 (N_1987,In_307,In_634);
and U1988 (N_1988,In_293,In_25);
and U1989 (N_1989,In_554,In_607);
or U1990 (N_1990,In_559,In_727);
nor U1991 (N_1991,In_722,In_316);
nand U1992 (N_1992,In_703,In_843);
nand U1993 (N_1993,In_972,In_512);
or U1994 (N_1994,In_559,In_121);
nor U1995 (N_1995,In_234,In_547);
nor U1996 (N_1996,In_17,In_155);
nand U1997 (N_1997,In_380,In_204);
and U1998 (N_1998,In_63,In_843);
nand U1999 (N_1999,In_655,In_123);
and U2000 (N_2000,In_304,In_726);
or U2001 (N_2001,In_356,In_743);
nand U2002 (N_2002,In_966,In_728);
and U2003 (N_2003,In_372,In_88);
or U2004 (N_2004,In_332,In_136);
nand U2005 (N_2005,In_362,In_690);
or U2006 (N_2006,In_586,In_772);
and U2007 (N_2007,In_814,In_76);
or U2008 (N_2008,In_265,In_263);
nand U2009 (N_2009,In_778,In_648);
and U2010 (N_2010,In_26,In_160);
nand U2011 (N_2011,In_304,In_446);
and U2012 (N_2012,In_912,In_341);
or U2013 (N_2013,In_335,In_794);
and U2014 (N_2014,In_431,In_381);
nor U2015 (N_2015,In_867,In_77);
nor U2016 (N_2016,In_613,In_397);
nor U2017 (N_2017,In_521,In_26);
nand U2018 (N_2018,In_938,In_54);
and U2019 (N_2019,In_875,In_119);
and U2020 (N_2020,In_8,In_925);
nand U2021 (N_2021,In_525,In_20);
nor U2022 (N_2022,In_960,In_374);
or U2023 (N_2023,In_141,In_869);
or U2024 (N_2024,In_507,In_535);
nand U2025 (N_2025,In_946,In_883);
nor U2026 (N_2026,In_749,In_667);
and U2027 (N_2027,In_653,In_197);
or U2028 (N_2028,In_437,In_799);
nand U2029 (N_2029,In_224,In_513);
nand U2030 (N_2030,In_278,In_378);
nor U2031 (N_2031,In_6,In_60);
or U2032 (N_2032,In_999,In_650);
nor U2033 (N_2033,In_478,In_690);
or U2034 (N_2034,In_540,In_337);
or U2035 (N_2035,In_801,In_928);
nand U2036 (N_2036,In_271,In_871);
nand U2037 (N_2037,In_813,In_962);
and U2038 (N_2038,In_855,In_771);
or U2039 (N_2039,In_208,In_620);
and U2040 (N_2040,In_328,In_725);
or U2041 (N_2041,In_880,In_40);
nand U2042 (N_2042,In_995,In_77);
nor U2043 (N_2043,In_196,In_655);
nor U2044 (N_2044,In_620,In_729);
or U2045 (N_2045,In_330,In_630);
nor U2046 (N_2046,In_899,In_819);
xor U2047 (N_2047,In_918,In_20);
nand U2048 (N_2048,In_478,In_785);
nor U2049 (N_2049,In_20,In_776);
nand U2050 (N_2050,In_721,In_115);
and U2051 (N_2051,In_434,In_592);
nand U2052 (N_2052,In_462,In_860);
and U2053 (N_2053,In_428,In_585);
or U2054 (N_2054,In_682,In_524);
nor U2055 (N_2055,In_79,In_847);
nand U2056 (N_2056,In_242,In_624);
nand U2057 (N_2057,In_786,In_69);
and U2058 (N_2058,In_134,In_105);
nand U2059 (N_2059,In_908,In_877);
nand U2060 (N_2060,In_176,In_279);
nand U2061 (N_2061,In_847,In_210);
and U2062 (N_2062,In_426,In_839);
or U2063 (N_2063,In_173,In_463);
and U2064 (N_2064,In_323,In_571);
nor U2065 (N_2065,In_787,In_158);
nand U2066 (N_2066,In_172,In_631);
and U2067 (N_2067,In_192,In_726);
nand U2068 (N_2068,In_961,In_367);
nand U2069 (N_2069,In_183,In_881);
or U2070 (N_2070,In_444,In_763);
nand U2071 (N_2071,In_61,In_0);
or U2072 (N_2072,In_401,In_463);
nand U2073 (N_2073,In_704,In_737);
and U2074 (N_2074,In_66,In_108);
nand U2075 (N_2075,In_57,In_642);
nand U2076 (N_2076,In_279,In_73);
or U2077 (N_2077,In_362,In_225);
and U2078 (N_2078,In_42,In_988);
nor U2079 (N_2079,In_749,In_997);
nor U2080 (N_2080,In_731,In_325);
nor U2081 (N_2081,In_994,In_236);
xor U2082 (N_2082,In_226,In_671);
and U2083 (N_2083,In_589,In_455);
nor U2084 (N_2084,In_721,In_816);
nand U2085 (N_2085,In_659,In_603);
or U2086 (N_2086,In_79,In_127);
nor U2087 (N_2087,In_638,In_58);
nor U2088 (N_2088,In_925,In_795);
and U2089 (N_2089,In_478,In_188);
and U2090 (N_2090,In_113,In_54);
nand U2091 (N_2091,In_152,In_771);
or U2092 (N_2092,In_457,In_415);
and U2093 (N_2093,In_329,In_857);
and U2094 (N_2094,In_582,In_309);
and U2095 (N_2095,In_939,In_987);
xnor U2096 (N_2096,In_970,In_615);
nor U2097 (N_2097,In_203,In_360);
nand U2098 (N_2098,In_117,In_213);
or U2099 (N_2099,In_824,In_454);
nand U2100 (N_2100,In_890,In_309);
nor U2101 (N_2101,In_73,In_112);
nor U2102 (N_2102,In_780,In_716);
nor U2103 (N_2103,In_841,In_839);
or U2104 (N_2104,In_414,In_330);
or U2105 (N_2105,In_308,In_618);
or U2106 (N_2106,In_324,In_633);
nand U2107 (N_2107,In_270,In_740);
and U2108 (N_2108,In_454,In_100);
or U2109 (N_2109,In_870,In_345);
nand U2110 (N_2110,In_434,In_260);
nand U2111 (N_2111,In_14,In_515);
or U2112 (N_2112,In_147,In_135);
nand U2113 (N_2113,In_957,In_226);
nor U2114 (N_2114,In_706,In_779);
or U2115 (N_2115,In_340,In_762);
and U2116 (N_2116,In_318,In_620);
nand U2117 (N_2117,In_163,In_605);
and U2118 (N_2118,In_339,In_841);
and U2119 (N_2119,In_859,In_578);
and U2120 (N_2120,In_859,In_851);
nor U2121 (N_2121,In_478,In_944);
nor U2122 (N_2122,In_281,In_543);
and U2123 (N_2123,In_507,In_543);
nor U2124 (N_2124,In_71,In_643);
or U2125 (N_2125,In_583,In_684);
nor U2126 (N_2126,In_731,In_868);
nand U2127 (N_2127,In_361,In_639);
nand U2128 (N_2128,In_889,In_32);
nand U2129 (N_2129,In_151,In_734);
or U2130 (N_2130,In_958,In_960);
or U2131 (N_2131,In_262,In_856);
and U2132 (N_2132,In_528,In_371);
or U2133 (N_2133,In_437,In_165);
nand U2134 (N_2134,In_878,In_435);
and U2135 (N_2135,In_786,In_501);
and U2136 (N_2136,In_917,In_591);
nor U2137 (N_2137,In_576,In_288);
nor U2138 (N_2138,In_458,In_502);
nand U2139 (N_2139,In_167,In_977);
or U2140 (N_2140,In_538,In_299);
or U2141 (N_2141,In_342,In_363);
nor U2142 (N_2142,In_312,In_162);
and U2143 (N_2143,In_203,In_783);
nand U2144 (N_2144,In_535,In_59);
nor U2145 (N_2145,In_562,In_875);
nand U2146 (N_2146,In_508,In_662);
nor U2147 (N_2147,In_959,In_15);
nand U2148 (N_2148,In_61,In_561);
or U2149 (N_2149,In_160,In_963);
nor U2150 (N_2150,In_33,In_774);
or U2151 (N_2151,In_574,In_901);
or U2152 (N_2152,In_884,In_762);
or U2153 (N_2153,In_476,In_857);
and U2154 (N_2154,In_778,In_529);
and U2155 (N_2155,In_369,In_429);
nand U2156 (N_2156,In_555,In_684);
nand U2157 (N_2157,In_750,In_604);
and U2158 (N_2158,In_760,In_155);
nand U2159 (N_2159,In_736,In_34);
or U2160 (N_2160,In_979,In_885);
nor U2161 (N_2161,In_346,In_501);
or U2162 (N_2162,In_153,In_816);
or U2163 (N_2163,In_250,In_31);
nor U2164 (N_2164,In_559,In_235);
or U2165 (N_2165,In_426,In_813);
or U2166 (N_2166,In_518,In_630);
or U2167 (N_2167,In_279,In_122);
and U2168 (N_2168,In_632,In_562);
nand U2169 (N_2169,In_579,In_925);
or U2170 (N_2170,In_144,In_897);
nand U2171 (N_2171,In_637,In_585);
nand U2172 (N_2172,In_469,In_614);
nor U2173 (N_2173,In_202,In_522);
nor U2174 (N_2174,In_636,In_83);
or U2175 (N_2175,In_771,In_398);
and U2176 (N_2176,In_589,In_919);
or U2177 (N_2177,In_367,In_378);
and U2178 (N_2178,In_685,In_969);
nor U2179 (N_2179,In_833,In_129);
and U2180 (N_2180,In_659,In_806);
nor U2181 (N_2181,In_436,In_569);
nor U2182 (N_2182,In_485,In_394);
nand U2183 (N_2183,In_708,In_172);
nand U2184 (N_2184,In_789,In_630);
or U2185 (N_2185,In_370,In_362);
nand U2186 (N_2186,In_455,In_248);
or U2187 (N_2187,In_248,In_123);
or U2188 (N_2188,In_512,In_573);
or U2189 (N_2189,In_97,In_961);
or U2190 (N_2190,In_917,In_113);
and U2191 (N_2191,In_635,In_14);
nor U2192 (N_2192,In_741,In_975);
nand U2193 (N_2193,In_137,In_466);
nand U2194 (N_2194,In_231,In_853);
nand U2195 (N_2195,In_474,In_720);
nor U2196 (N_2196,In_414,In_629);
or U2197 (N_2197,In_714,In_313);
xnor U2198 (N_2198,In_408,In_905);
nor U2199 (N_2199,In_627,In_459);
or U2200 (N_2200,In_79,In_487);
or U2201 (N_2201,In_596,In_683);
and U2202 (N_2202,In_373,In_284);
and U2203 (N_2203,In_958,In_400);
nor U2204 (N_2204,In_75,In_36);
nand U2205 (N_2205,In_988,In_707);
and U2206 (N_2206,In_61,In_840);
nor U2207 (N_2207,In_987,In_24);
and U2208 (N_2208,In_831,In_350);
and U2209 (N_2209,In_897,In_161);
and U2210 (N_2210,In_602,In_584);
and U2211 (N_2211,In_206,In_310);
nand U2212 (N_2212,In_285,In_235);
and U2213 (N_2213,In_808,In_89);
or U2214 (N_2214,In_798,In_150);
nor U2215 (N_2215,In_38,In_227);
nand U2216 (N_2216,In_961,In_511);
or U2217 (N_2217,In_997,In_119);
and U2218 (N_2218,In_600,In_710);
or U2219 (N_2219,In_900,In_876);
nand U2220 (N_2220,In_172,In_534);
or U2221 (N_2221,In_178,In_619);
nor U2222 (N_2222,In_465,In_792);
nand U2223 (N_2223,In_233,In_657);
nand U2224 (N_2224,In_987,In_237);
or U2225 (N_2225,In_305,In_849);
or U2226 (N_2226,In_793,In_990);
or U2227 (N_2227,In_30,In_298);
nand U2228 (N_2228,In_443,In_803);
nand U2229 (N_2229,In_627,In_299);
or U2230 (N_2230,In_332,In_875);
or U2231 (N_2231,In_644,In_924);
or U2232 (N_2232,In_668,In_588);
nand U2233 (N_2233,In_553,In_171);
or U2234 (N_2234,In_668,In_18);
or U2235 (N_2235,In_743,In_361);
nor U2236 (N_2236,In_109,In_458);
nor U2237 (N_2237,In_889,In_746);
or U2238 (N_2238,In_625,In_270);
nor U2239 (N_2239,In_783,In_941);
or U2240 (N_2240,In_47,In_16);
nand U2241 (N_2241,In_886,In_518);
and U2242 (N_2242,In_839,In_672);
or U2243 (N_2243,In_287,In_208);
or U2244 (N_2244,In_135,In_317);
nor U2245 (N_2245,In_223,In_805);
nand U2246 (N_2246,In_974,In_122);
nand U2247 (N_2247,In_90,In_989);
or U2248 (N_2248,In_283,In_467);
nand U2249 (N_2249,In_246,In_665);
nor U2250 (N_2250,In_930,In_489);
nand U2251 (N_2251,In_596,In_334);
nor U2252 (N_2252,In_330,In_618);
or U2253 (N_2253,In_254,In_776);
and U2254 (N_2254,In_586,In_875);
nor U2255 (N_2255,In_957,In_565);
nand U2256 (N_2256,In_197,In_431);
nand U2257 (N_2257,In_727,In_889);
or U2258 (N_2258,In_504,In_851);
nor U2259 (N_2259,In_121,In_662);
nand U2260 (N_2260,In_147,In_868);
nand U2261 (N_2261,In_988,In_295);
nand U2262 (N_2262,In_316,In_296);
and U2263 (N_2263,In_772,In_192);
or U2264 (N_2264,In_100,In_398);
xnor U2265 (N_2265,In_602,In_327);
or U2266 (N_2266,In_11,In_808);
nand U2267 (N_2267,In_819,In_891);
nor U2268 (N_2268,In_31,In_916);
nand U2269 (N_2269,In_706,In_877);
nor U2270 (N_2270,In_496,In_121);
or U2271 (N_2271,In_613,In_593);
and U2272 (N_2272,In_351,In_641);
nand U2273 (N_2273,In_272,In_240);
and U2274 (N_2274,In_73,In_873);
nand U2275 (N_2275,In_533,In_359);
or U2276 (N_2276,In_58,In_302);
or U2277 (N_2277,In_326,In_829);
or U2278 (N_2278,In_25,In_11);
nor U2279 (N_2279,In_821,In_148);
nand U2280 (N_2280,In_135,In_694);
nand U2281 (N_2281,In_650,In_601);
or U2282 (N_2282,In_986,In_814);
and U2283 (N_2283,In_487,In_166);
nand U2284 (N_2284,In_701,In_255);
nand U2285 (N_2285,In_412,In_332);
or U2286 (N_2286,In_48,In_202);
or U2287 (N_2287,In_157,In_813);
nor U2288 (N_2288,In_229,In_72);
or U2289 (N_2289,In_602,In_120);
nand U2290 (N_2290,In_171,In_534);
nand U2291 (N_2291,In_216,In_385);
or U2292 (N_2292,In_191,In_478);
nor U2293 (N_2293,In_814,In_282);
and U2294 (N_2294,In_439,In_345);
nor U2295 (N_2295,In_120,In_189);
or U2296 (N_2296,In_558,In_545);
nor U2297 (N_2297,In_857,In_479);
nand U2298 (N_2298,In_95,In_173);
nand U2299 (N_2299,In_522,In_889);
nand U2300 (N_2300,In_432,In_236);
and U2301 (N_2301,In_425,In_540);
nor U2302 (N_2302,In_455,In_422);
or U2303 (N_2303,In_353,In_717);
or U2304 (N_2304,In_587,In_927);
nand U2305 (N_2305,In_437,In_511);
and U2306 (N_2306,In_449,In_869);
nor U2307 (N_2307,In_151,In_301);
nor U2308 (N_2308,In_676,In_4);
or U2309 (N_2309,In_234,In_957);
nor U2310 (N_2310,In_553,In_894);
nor U2311 (N_2311,In_410,In_844);
or U2312 (N_2312,In_898,In_896);
nor U2313 (N_2313,In_273,In_317);
nand U2314 (N_2314,In_416,In_286);
nand U2315 (N_2315,In_176,In_51);
nand U2316 (N_2316,In_592,In_974);
nand U2317 (N_2317,In_633,In_314);
or U2318 (N_2318,In_248,In_361);
and U2319 (N_2319,In_411,In_955);
or U2320 (N_2320,In_493,In_607);
nand U2321 (N_2321,In_580,In_575);
or U2322 (N_2322,In_843,In_666);
nor U2323 (N_2323,In_208,In_506);
or U2324 (N_2324,In_243,In_788);
and U2325 (N_2325,In_122,In_136);
or U2326 (N_2326,In_661,In_148);
nor U2327 (N_2327,In_455,In_131);
and U2328 (N_2328,In_994,In_784);
or U2329 (N_2329,In_972,In_843);
nand U2330 (N_2330,In_243,In_805);
nand U2331 (N_2331,In_625,In_860);
nor U2332 (N_2332,In_264,In_469);
nand U2333 (N_2333,In_545,In_764);
nor U2334 (N_2334,In_454,In_659);
nand U2335 (N_2335,In_274,In_254);
or U2336 (N_2336,In_670,In_572);
or U2337 (N_2337,In_386,In_450);
nand U2338 (N_2338,In_66,In_470);
and U2339 (N_2339,In_349,In_788);
or U2340 (N_2340,In_818,In_460);
xnor U2341 (N_2341,In_911,In_467);
nand U2342 (N_2342,In_876,In_856);
or U2343 (N_2343,In_263,In_160);
nor U2344 (N_2344,In_16,In_676);
and U2345 (N_2345,In_39,In_68);
nand U2346 (N_2346,In_583,In_709);
and U2347 (N_2347,In_270,In_157);
xor U2348 (N_2348,In_72,In_687);
nand U2349 (N_2349,In_578,In_472);
and U2350 (N_2350,In_598,In_303);
nor U2351 (N_2351,In_754,In_787);
or U2352 (N_2352,In_410,In_939);
nor U2353 (N_2353,In_424,In_181);
nand U2354 (N_2354,In_529,In_36);
nor U2355 (N_2355,In_965,In_543);
nand U2356 (N_2356,In_996,In_684);
nor U2357 (N_2357,In_75,In_712);
and U2358 (N_2358,In_900,In_932);
nand U2359 (N_2359,In_135,In_535);
nor U2360 (N_2360,In_41,In_513);
nand U2361 (N_2361,In_914,In_454);
nor U2362 (N_2362,In_557,In_183);
and U2363 (N_2363,In_657,In_476);
nand U2364 (N_2364,In_483,In_623);
nand U2365 (N_2365,In_7,In_973);
and U2366 (N_2366,In_114,In_672);
or U2367 (N_2367,In_808,In_10);
or U2368 (N_2368,In_309,In_105);
or U2369 (N_2369,In_574,In_488);
or U2370 (N_2370,In_929,In_101);
or U2371 (N_2371,In_985,In_312);
nor U2372 (N_2372,In_348,In_594);
nand U2373 (N_2373,In_363,In_264);
nand U2374 (N_2374,In_7,In_10);
nand U2375 (N_2375,In_150,In_264);
or U2376 (N_2376,In_892,In_971);
and U2377 (N_2377,In_357,In_300);
nor U2378 (N_2378,In_570,In_137);
or U2379 (N_2379,In_624,In_503);
or U2380 (N_2380,In_679,In_591);
nand U2381 (N_2381,In_173,In_733);
nand U2382 (N_2382,In_325,In_820);
nand U2383 (N_2383,In_379,In_87);
nor U2384 (N_2384,In_118,In_551);
xnor U2385 (N_2385,In_391,In_874);
and U2386 (N_2386,In_5,In_307);
or U2387 (N_2387,In_908,In_728);
nand U2388 (N_2388,In_804,In_164);
and U2389 (N_2389,In_608,In_625);
nand U2390 (N_2390,In_70,In_311);
or U2391 (N_2391,In_623,In_233);
or U2392 (N_2392,In_935,In_368);
xnor U2393 (N_2393,In_840,In_596);
nor U2394 (N_2394,In_761,In_902);
and U2395 (N_2395,In_395,In_381);
or U2396 (N_2396,In_964,In_810);
nand U2397 (N_2397,In_453,In_197);
nand U2398 (N_2398,In_814,In_328);
or U2399 (N_2399,In_442,In_321);
nand U2400 (N_2400,In_29,In_472);
or U2401 (N_2401,In_998,In_851);
or U2402 (N_2402,In_553,In_325);
nand U2403 (N_2403,In_635,In_621);
nor U2404 (N_2404,In_770,In_678);
nand U2405 (N_2405,In_471,In_515);
nor U2406 (N_2406,In_300,In_683);
and U2407 (N_2407,In_644,In_665);
and U2408 (N_2408,In_148,In_23);
or U2409 (N_2409,In_783,In_621);
and U2410 (N_2410,In_447,In_467);
or U2411 (N_2411,In_347,In_527);
and U2412 (N_2412,In_587,In_469);
nand U2413 (N_2413,In_159,In_539);
or U2414 (N_2414,In_430,In_762);
or U2415 (N_2415,In_170,In_695);
nor U2416 (N_2416,In_636,In_912);
or U2417 (N_2417,In_615,In_755);
nor U2418 (N_2418,In_464,In_979);
or U2419 (N_2419,In_964,In_175);
nor U2420 (N_2420,In_934,In_902);
nand U2421 (N_2421,In_366,In_673);
nor U2422 (N_2422,In_869,In_490);
nand U2423 (N_2423,In_141,In_227);
nor U2424 (N_2424,In_823,In_434);
nor U2425 (N_2425,In_932,In_947);
and U2426 (N_2426,In_448,In_221);
or U2427 (N_2427,In_847,In_20);
nor U2428 (N_2428,In_552,In_179);
nor U2429 (N_2429,In_701,In_846);
nor U2430 (N_2430,In_938,In_982);
nand U2431 (N_2431,In_685,In_193);
nand U2432 (N_2432,In_713,In_103);
nor U2433 (N_2433,In_630,In_656);
or U2434 (N_2434,In_334,In_23);
or U2435 (N_2435,In_470,In_85);
and U2436 (N_2436,In_427,In_489);
or U2437 (N_2437,In_195,In_320);
nand U2438 (N_2438,In_538,In_645);
or U2439 (N_2439,In_285,In_518);
or U2440 (N_2440,In_225,In_291);
nor U2441 (N_2441,In_803,In_18);
and U2442 (N_2442,In_938,In_365);
nand U2443 (N_2443,In_283,In_182);
nor U2444 (N_2444,In_714,In_131);
nor U2445 (N_2445,In_693,In_325);
or U2446 (N_2446,In_632,In_829);
or U2447 (N_2447,In_324,In_610);
nand U2448 (N_2448,In_696,In_368);
nor U2449 (N_2449,In_218,In_881);
nor U2450 (N_2450,In_325,In_217);
xor U2451 (N_2451,In_9,In_993);
nand U2452 (N_2452,In_74,In_11);
or U2453 (N_2453,In_59,In_576);
and U2454 (N_2454,In_382,In_712);
nor U2455 (N_2455,In_455,In_70);
nor U2456 (N_2456,In_709,In_769);
and U2457 (N_2457,In_534,In_663);
nand U2458 (N_2458,In_305,In_324);
nand U2459 (N_2459,In_806,In_398);
and U2460 (N_2460,In_391,In_627);
nor U2461 (N_2461,In_795,In_386);
and U2462 (N_2462,In_978,In_558);
nor U2463 (N_2463,In_169,In_661);
and U2464 (N_2464,In_26,In_906);
nor U2465 (N_2465,In_192,In_11);
and U2466 (N_2466,In_377,In_573);
nor U2467 (N_2467,In_108,In_656);
nor U2468 (N_2468,In_502,In_687);
nand U2469 (N_2469,In_405,In_519);
nor U2470 (N_2470,In_375,In_659);
or U2471 (N_2471,In_63,In_653);
or U2472 (N_2472,In_136,In_162);
nand U2473 (N_2473,In_824,In_108);
and U2474 (N_2474,In_197,In_102);
nor U2475 (N_2475,In_112,In_847);
or U2476 (N_2476,In_643,In_399);
and U2477 (N_2477,In_825,In_740);
or U2478 (N_2478,In_381,In_514);
nand U2479 (N_2479,In_382,In_295);
or U2480 (N_2480,In_744,In_385);
and U2481 (N_2481,In_218,In_260);
or U2482 (N_2482,In_335,In_749);
nand U2483 (N_2483,In_710,In_17);
nor U2484 (N_2484,In_220,In_329);
or U2485 (N_2485,In_828,In_174);
and U2486 (N_2486,In_7,In_250);
nand U2487 (N_2487,In_13,In_353);
nor U2488 (N_2488,In_202,In_241);
and U2489 (N_2489,In_433,In_145);
and U2490 (N_2490,In_120,In_724);
nor U2491 (N_2491,In_682,In_444);
nand U2492 (N_2492,In_787,In_182);
nor U2493 (N_2493,In_308,In_900);
or U2494 (N_2494,In_43,In_456);
nand U2495 (N_2495,In_545,In_827);
or U2496 (N_2496,In_4,In_278);
nand U2497 (N_2497,In_181,In_5);
nand U2498 (N_2498,In_187,In_480);
or U2499 (N_2499,In_480,In_595);
and U2500 (N_2500,In_302,In_764);
nor U2501 (N_2501,In_9,In_176);
nand U2502 (N_2502,In_76,In_119);
or U2503 (N_2503,In_228,In_989);
or U2504 (N_2504,In_330,In_889);
nand U2505 (N_2505,In_605,In_457);
nand U2506 (N_2506,In_812,In_870);
nand U2507 (N_2507,In_785,In_186);
and U2508 (N_2508,In_983,In_372);
nand U2509 (N_2509,In_260,In_913);
nand U2510 (N_2510,In_704,In_867);
or U2511 (N_2511,In_229,In_356);
and U2512 (N_2512,In_353,In_789);
or U2513 (N_2513,In_418,In_687);
and U2514 (N_2514,In_705,In_5);
or U2515 (N_2515,In_790,In_662);
xor U2516 (N_2516,In_794,In_568);
nor U2517 (N_2517,In_552,In_97);
and U2518 (N_2518,In_876,In_677);
and U2519 (N_2519,In_287,In_682);
nand U2520 (N_2520,In_431,In_768);
and U2521 (N_2521,In_594,In_980);
nor U2522 (N_2522,In_402,In_197);
and U2523 (N_2523,In_505,In_688);
nor U2524 (N_2524,In_238,In_799);
nor U2525 (N_2525,In_939,In_993);
and U2526 (N_2526,In_577,In_803);
and U2527 (N_2527,In_922,In_391);
nor U2528 (N_2528,In_351,In_816);
nor U2529 (N_2529,In_653,In_921);
or U2530 (N_2530,In_635,In_710);
nor U2531 (N_2531,In_817,In_318);
and U2532 (N_2532,In_673,In_737);
nor U2533 (N_2533,In_16,In_783);
nand U2534 (N_2534,In_156,In_772);
or U2535 (N_2535,In_145,In_115);
nand U2536 (N_2536,In_271,In_903);
and U2537 (N_2537,In_339,In_546);
or U2538 (N_2538,In_328,In_937);
nand U2539 (N_2539,In_577,In_683);
or U2540 (N_2540,In_538,In_8);
or U2541 (N_2541,In_225,In_807);
nor U2542 (N_2542,In_970,In_304);
nand U2543 (N_2543,In_774,In_858);
or U2544 (N_2544,In_320,In_846);
and U2545 (N_2545,In_181,In_545);
or U2546 (N_2546,In_998,In_758);
nand U2547 (N_2547,In_779,In_718);
nor U2548 (N_2548,In_284,In_693);
and U2549 (N_2549,In_237,In_736);
and U2550 (N_2550,In_681,In_222);
and U2551 (N_2551,In_640,In_926);
nand U2552 (N_2552,In_863,In_46);
and U2553 (N_2553,In_904,In_517);
nor U2554 (N_2554,In_131,In_484);
and U2555 (N_2555,In_880,In_83);
nor U2556 (N_2556,In_488,In_176);
nor U2557 (N_2557,In_405,In_246);
or U2558 (N_2558,In_103,In_987);
nand U2559 (N_2559,In_9,In_853);
and U2560 (N_2560,In_785,In_464);
nor U2561 (N_2561,In_182,In_331);
nor U2562 (N_2562,In_203,In_816);
nor U2563 (N_2563,In_212,In_805);
and U2564 (N_2564,In_173,In_14);
xor U2565 (N_2565,In_76,In_478);
or U2566 (N_2566,In_109,In_132);
and U2567 (N_2567,In_559,In_78);
and U2568 (N_2568,In_986,In_295);
and U2569 (N_2569,In_898,In_849);
or U2570 (N_2570,In_38,In_350);
nand U2571 (N_2571,In_670,In_349);
or U2572 (N_2572,In_496,In_638);
nor U2573 (N_2573,In_755,In_818);
nand U2574 (N_2574,In_77,In_627);
nand U2575 (N_2575,In_188,In_312);
nand U2576 (N_2576,In_660,In_66);
nand U2577 (N_2577,In_516,In_360);
or U2578 (N_2578,In_259,In_272);
and U2579 (N_2579,In_845,In_831);
nand U2580 (N_2580,In_563,In_448);
or U2581 (N_2581,In_440,In_463);
or U2582 (N_2582,In_808,In_107);
nand U2583 (N_2583,In_754,In_903);
and U2584 (N_2584,In_893,In_91);
nor U2585 (N_2585,In_212,In_184);
nor U2586 (N_2586,In_314,In_400);
nor U2587 (N_2587,In_308,In_527);
nand U2588 (N_2588,In_610,In_39);
nand U2589 (N_2589,In_885,In_176);
and U2590 (N_2590,In_4,In_942);
nand U2591 (N_2591,In_413,In_12);
nor U2592 (N_2592,In_820,In_742);
or U2593 (N_2593,In_983,In_489);
and U2594 (N_2594,In_488,In_651);
nor U2595 (N_2595,In_498,In_178);
nand U2596 (N_2596,In_361,In_792);
nand U2597 (N_2597,In_791,In_871);
or U2598 (N_2598,In_768,In_992);
nand U2599 (N_2599,In_202,In_334);
nand U2600 (N_2600,In_278,In_947);
or U2601 (N_2601,In_802,In_319);
nand U2602 (N_2602,In_179,In_548);
nor U2603 (N_2603,In_165,In_85);
nand U2604 (N_2604,In_228,In_427);
xor U2605 (N_2605,In_788,In_911);
nand U2606 (N_2606,In_142,In_861);
or U2607 (N_2607,In_305,In_951);
or U2608 (N_2608,In_955,In_184);
nand U2609 (N_2609,In_618,In_473);
and U2610 (N_2610,In_557,In_673);
or U2611 (N_2611,In_651,In_54);
nand U2612 (N_2612,In_767,In_597);
nor U2613 (N_2613,In_773,In_884);
and U2614 (N_2614,In_984,In_404);
and U2615 (N_2615,In_614,In_653);
nand U2616 (N_2616,In_767,In_379);
nor U2617 (N_2617,In_886,In_31);
or U2618 (N_2618,In_800,In_940);
or U2619 (N_2619,In_380,In_28);
and U2620 (N_2620,In_770,In_257);
and U2621 (N_2621,In_566,In_750);
nand U2622 (N_2622,In_916,In_206);
nand U2623 (N_2623,In_853,In_593);
nand U2624 (N_2624,In_118,In_775);
or U2625 (N_2625,In_723,In_729);
nor U2626 (N_2626,In_396,In_102);
nor U2627 (N_2627,In_556,In_464);
nand U2628 (N_2628,In_559,In_22);
nand U2629 (N_2629,In_347,In_332);
and U2630 (N_2630,In_530,In_50);
nor U2631 (N_2631,In_718,In_889);
or U2632 (N_2632,In_428,In_147);
nand U2633 (N_2633,In_448,In_626);
or U2634 (N_2634,In_269,In_292);
nand U2635 (N_2635,In_951,In_648);
nor U2636 (N_2636,In_808,In_61);
or U2637 (N_2637,In_709,In_762);
or U2638 (N_2638,In_243,In_324);
or U2639 (N_2639,In_987,In_62);
nor U2640 (N_2640,In_98,In_261);
or U2641 (N_2641,In_19,In_849);
nor U2642 (N_2642,In_816,In_741);
nor U2643 (N_2643,In_524,In_522);
nand U2644 (N_2644,In_263,In_345);
nand U2645 (N_2645,In_652,In_489);
nand U2646 (N_2646,In_771,In_527);
or U2647 (N_2647,In_451,In_336);
and U2648 (N_2648,In_40,In_493);
and U2649 (N_2649,In_181,In_894);
nand U2650 (N_2650,In_537,In_433);
and U2651 (N_2651,In_828,In_475);
nand U2652 (N_2652,In_124,In_264);
and U2653 (N_2653,In_861,In_380);
nor U2654 (N_2654,In_28,In_570);
and U2655 (N_2655,In_363,In_927);
or U2656 (N_2656,In_782,In_372);
nor U2657 (N_2657,In_13,In_858);
or U2658 (N_2658,In_680,In_882);
nand U2659 (N_2659,In_837,In_615);
nand U2660 (N_2660,In_391,In_224);
or U2661 (N_2661,In_209,In_747);
nor U2662 (N_2662,In_375,In_54);
and U2663 (N_2663,In_692,In_386);
or U2664 (N_2664,In_275,In_980);
and U2665 (N_2665,In_463,In_209);
nor U2666 (N_2666,In_147,In_343);
nor U2667 (N_2667,In_398,In_514);
nand U2668 (N_2668,In_137,In_533);
and U2669 (N_2669,In_549,In_237);
and U2670 (N_2670,In_772,In_518);
nand U2671 (N_2671,In_964,In_768);
or U2672 (N_2672,In_311,In_999);
or U2673 (N_2673,In_870,In_674);
nand U2674 (N_2674,In_545,In_315);
nand U2675 (N_2675,In_576,In_281);
or U2676 (N_2676,In_419,In_569);
and U2677 (N_2677,In_890,In_134);
or U2678 (N_2678,In_99,In_188);
nand U2679 (N_2679,In_213,In_777);
nand U2680 (N_2680,In_563,In_953);
nand U2681 (N_2681,In_518,In_993);
nor U2682 (N_2682,In_842,In_79);
nand U2683 (N_2683,In_683,In_333);
nor U2684 (N_2684,In_464,In_948);
and U2685 (N_2685,In_778,In_677);
or U2686 (N_2686,In_586,In_500);
nand U2687 (N_2687,In_446,In_71);
nand U2688 (N_2688,In_139,In_382);
or U2689 (N_2689,In_175,In_623);
nand U2690 (N_2690,In_574,In_704);
nor U2691 (N_2691,In_76,In_632);
nor U2692 (N_2692,In_402,In_498);
nor U2693 (N_2693,In_79,In_78);
and U2694 (N_2694,In_540,In_693);
and U2695 (N_2695,In_45,In_668);
nand U2696 (N_2696,In_18,In_669);
and U2697 (N_2697,In_119,In_306);
or U2698 (N_2698,In_491,In_283);
nor U2699 (N_2699,In_949,In_759);
and U2700 (N_2700,In_221,In_823);
and U2701 (N_2701,In_407,In_546);
nor U2702 (N_2702,In_826,In_437);
nor U2703 (N_2703,In_306,In_109);
nand U2704 (N_2704,In_108,In_398);
nand U2705 (N_2705,In_26,In_967);
and U2706 (N_2706,In_542,In_183);
or U2707 (N_2707,In_649,In_409);
or U2708 (N_2708,In_229,In_993);
nor U2709 (N_2709,In_262,In_147);
or U2710 (N_2710,In_874,In_903);
nand U2711 (N_2711,In_5,In_941);
nor U2712 (N_2712,In_80,In_837);
and U2713 (N_2713,In_337,In_409);
nor U2714 (N_2714,In_740,In_516);
nor U2715 (N_2715,In_235,In_240);
nand U2716 (N_2716,In_873,In_212);
or U2717 (N_2717,In_327,In_316);
and U2718 (N_2718,In_698,In_435);
nor U2719 (N_2719,In_801,In_29);
nor U2720 (N_2720,In_657,In_919);
or U2721 (N_2721,In_922,In_917);
and U2722 (N_2722,In_578,In_750);
nand U2723 (N_2723,In_188,In_424);
nor U2724 (N_2724,In_841,In_619);
nor U2725 (N_2725,In_458,In_918);
nor U2726 (N_2726,In_41,In_993);
or U2727 (N_2727,In_460,In_600);
nand U2728 (N_2728,In_204,In_979);
nor U2729 (N_2729,In_252,In_744);
nor U2730 (N_2730,In_111,In_155);
nor U2731 (N_2731,In_193,In_936);
nor U2732 (N_2732,In_96,In_10);
and U2733 (N_2733,In_719,In_237);
nor U2734 (N_2734,In_994,In_619);
or U2735 (N_2735,In_390,In_95);
nand U2736 (N_2736,In_798,In_587);
nand U2737 (N_2737,In_739,In_919);
nor U2738 (N_2738,In_480,In_786);
nor U2739 (N_2739,In_259,In_512);
nor U2740 (N_2740,In_306,In_597);
and U2741 (N_2741,In_106,In_913);
and U2742 (N_2742,In_535,In_811);
or U2743 (N_2743,In_86,In_276);
nor U2744 (N_2744,In_438,In_820);
nand U2745 (N_2745,In_444,In_909);
nand U2746 (N_2746,In_170,In_509);
nor U2747 (N_2747,In_93,In_572);
and U2748 (N_2748,In_356,In_763);
nand U2749 (N_2749,In_282,In_359);
nand U2750 (N_2750,In_311,In_360);
nor U2751 (N_2751,In_650,In_723);
and U2752 (N_2752,In_539,In_431);
nand U2753 (N_2753,In_553,In_640);
nor U2754 (N_2754,In_967,In_309);
nor U2755 (N_2755,In_600,In_711);
or U2756 (N_2756,In_470,In_896);
or U2757 (N_2757,In_428,In_256);
or U2758 (N_2758,In_943,In_972);
nor U2759 (N_2759,In_399,In_732);
nand U2760 (N_2760,In_388,In_949);
nor U2761 (N_2761,In_419,In_81);
or U2762 (N_2762,In_304,In_391);
and U2763 (N_2763,In_296,In_165);
and U2764 (N_2764,In_421,In_124);
and U2765 (N_2765,In_891,In_611);
nor U2766 (N_2766,In_998,In_544);
nand U2767 (N_2767,In_190,In_869);
nor U2768 (N_2768,In_308,In_224);
nand U2769 (N_2769,In_959,In_587);
nand U2770 (N_2770,In_611,In_576);
and U2771 (N_2771,In_863,In_901);
or U2772 (N_2772,In_634,In_827);
or U2773 (N_2773,In_106,In_751);
and U2774 (N_2774,In_853,In_283);
nand U2775 (N_2775,In_130,In_917);
nor U2776 (N_2776,In_925,In_163);
nor U2777 (N_2777,In_791,In_682);
nor U2778 (N_2778,In_650,In_436);
or U2779 (N_2779,In_622,In_467);
nand U2780 (N_2780,In_632,In_531);
or U2781 (N_2781,In_141,In_812);
nand U2782 (N_2782,In_116,In_414);
and U2783 (N_2783,In_699,In_679);
nand U2784 (N_2784,In_72,In_600);
nor U2785 (N_2785,In_170,In_414);
nor U2786 (N_2786,In_996,In_702);
or U2787 (N_2787,In_947,In_793);
nand U2788 (N_2788,In_543,In_692);
nand U2789 (N_2789,In_516,In_446);
nand U2790 (N_2790,In_769,In_597);
nor U2791 (N_2791,In_593,In_774);
nand U2792 (N_2792,In_95,In_910);
or U2793 (N_2793,In_544,In_91);
nor U2794 (N_2794,In_89,In_618);
or U2795 (N_2795,In_590,In_602);
and U2796 (N_2796,In_317,In_9);
and U2797 (N_2797,In_279,In_592);
nand U2798 (N_2798,In_63,In_331);
nand U2799 (N_2799,In_496,In_323);
or U2800 (N_2800,In_63,In_561);
and U2801 (N_2801,In_540,In_605);
nand U2802 (N_2802,In_514,In_275);
nand U2803 (N_2803,In_562,In_806);
or U2804 (N_2804,In_105,In_427);
nand U2805 (N_2805,In_326,In_609);
nor U2806 (N_2806,In_432,In_696);
nor U2807 (N_2807,In_584,In_619);
and U2808 (N_2808,In_248,In_567);
and U2809 (N_2809,In_285,In_893);
nand U2810 (N_2810,In_981,In_839);
nor U2811 (N_2811,In_618,In_472);
nor U2812 (N_2812,In_914,In_700);
or U2813 (N_2813,In_444,In_489);
nand U2814 (N_2814,In_325,In_942);
or U2815 (N_2815,In_750,In_110);
and U2816 (N_2816,In_604,In_119);
nor U2817 (N_2817,In_455,In_7);
nor U2818 (N_2818,In_199,In_523);
and U2819 (N_2819,In_184,In_704);
and U2820 (N_2820,In_709,In_728);
and U2821 (N_2821,In_502,In_268);
or U2822 (N_2822,In_206,In_252);
or U2823 (N_2823,In_654,In_885);
nor U2824 (N_2824,In_382,In_686);
nor U2825 (N_2825,In_534,In_170);
and U2826 (N_2826,In_314,In_521);
nand U2827 (N_2827,In_108,In_313);
nor U2828 (N_2828,In_405,In_122);
xnor U2829 (N_2829,In_120,In_127);
and U2830 (N_2830,In_828,In_608);
nor U2831 (N_2831,In_347,In_374);
nor U2832 (N_2832,In_400,In_730);
and U2833 (N_2833,In_896,In_975);
nor U2834 (N_2834,In_896,In_908);
nand U2835 (N_2835,In_522,In_774);
and U2836 (N_2836,In_745,In_920);
nand U2837 (N_2837,In_77,In_236);
nor U2838 (N_2838,In_149,In_156);
and U2839 (N_2839,In_744,In_547);
nand U2840 (N_2840,In_423,In_81);
or U2841 (N_2841,In_50,In_499);
and U2842 (N_2842,In_334,In_965);
nor U2843 (N_2843,In_250,In_421);
or U2844 (N_2844,In_950,In_886);
and U2845 (N_2845,In_159,In_231);
nor U2846 (N_2846,In_907,In_791);
nor U2847 (N_2847,In_683,In_464);
and U2848 (N_2848,In_255,In_487);
or U2849 (N_2849,In_380,In_616);
nor U2850 (N_2850,In_840,In_100);
and U2851 (N_2851,In_379,In_865);
and U2852 (N_2852,In_916,In_83);
nand U2853 (N_2853,In_959,In_311);
nand U2854 (N_2854,In_921,In_864);
or U2855 (N_2855,In_338,In_993);
and U2856 (N_2856,In_539,In_408);
nand U2857 (N_2857,In_846,In_816);
nor U2858 (N_2858,In_88,In_631);
or U2859 (N_2859,In_101,In_230);
or U2860 (N_2860,In_788,In_734);
nor U2861 (N_2861,In_137,In_284);
nand U2862 (N_2862,In_609,In_147);
or U2863 (N_2863,In_713,In_936);
nor U2864 (N_2864,In_42,In_355);
nand U2865 (N_2865,In_109,In_213);
or U2866 (N_2866,In_140,In_889);
or U2867 (N_2867,In_112,In_822);
and U2868 (N_2868,In_267,In_993);
or U2869 (N_2869,In_496,In_483);
nand U2870 (N_2870,In_260,In_305);
or U2871 (N_2871,In_957,In_285);
nand U2872 (N_2872,In_222,In_482);
nand U2873 (N_2873,In_703,In_262);
and U2874 (N_2874,In_424,In_991);
nor U2875 (N_2875,In_633,In_518);
or U2876 (N_2876,In_879,In_660);
and U2877 (N_2877,In_720,In_534);
and U2878 (N_2878,In_79,In_190);
nor U2879 (N_2879,In_559,In_946);
and U2880 (N_2880,In_974,In_756);
nand U2881 (N_2881,In_10,In_499);
or U2882 (N_2882,In_888,In_617);
and U2883 (N_2883,In_386,In_974);
nor U2884 (N_2884,In_276,In_239);
or U2885 (N_2885,In_938,In_547);
or U2886 (N_2886,In_457,In_188);
and U2887 (N_2887,In_436,In_150);
nand U2888 (N_2888,In_266,In_504);
nand U2889 (N_2889,In_668,In_466);
or U2890 (N_2890,In_885,In_456);
and U2891 (N_2891,In_711,In_531);
nor U2892 (N_2892,In_521,In_727);
and U2893 (N_2893,In_120,In_641);
or U2894 (N_2894,In_604,In_903);
nand U2895 (N_2895,In_803,In_463);
nand U2896 (N_2896,In_759,In_725);
and U2897 (N_2897,In_748,In_331);
nor U2898 (N_2898,In_635,In_612);
and U2899 (N_2899,In_670,In_339);
nand U2900 (N_2900,In_747,In_560);
and U2901 (N_2901,In_514,In_775);
and U2902 (N_2902,In_996,In_320);
xnor U2903 (N_2903,In_804,In_116);
nor U2904 (N_2904,In_542,In_581);
nand U2905 (N_2905,In_434,In_326);
nand U2906 (N_2906,In_547,In_625);
and U2907 (N_2907,In_677,In_74);
nor U2908 (N_2908,In_395,In_89);
nand U2909 (N_2909,In_148,In_768);
and U2910 (N_2910,In_884,In_745);
nor U2911 (N_2911,In_529,In_776);
and U2912 (N_2912,In_557,In_139);
nor U2913 (N_2913,In_62,In_813);
or U2914 (N_2914,In_406,In_274);
nor U2915 (N_2915,In_978,In_210);
xor U2916 (N_2916,In_401,In_2);
nor U2917 (N_2917,In_392,In_410);
or U2918 (N_2918,In_169,In_875);
or U2919 (N_2919,In_578,In_507);
and U2920 (N_2920,In_881,In_748);
and U2921 (N_2921,In_499,In_593);
nand U2922 (N_2922,In_380,In_802);
and U2923 (N_2923,In_203,In_653);
or U2924 (N_2924,In_864,In_893);
nor U2925 (N_2925,In_438,In_469);
nand U2926 (N_2926,In_525,In_963);
nor U2927 (N_2927,In_466,In_470);
and U2928 (N_2928,In_34,In_194);
and U2929 (N_2929,In_235,In_997);
nor U2930 (N_2930,In_314,In_448);
or U2931 (N_2931,In_835,In_132);
nor U2932 (N_2932,In_673,In_297);
nand U2933 (N_2933,In_124,In_509);
or U2934 (N_2934,In_997,In_23);
or U2935 (N_2935,In_805,In_514);
and U2936 (N_2936,In_131,In_412);
and U2937 (N_2937,In_780,In_427);
xnor U2938 (N_2938,In_533,In_407);
nor U2939 (N_2939,In_769,In_900);
or U2940 (N_2940,In_706,In_295);
nor U2941 (N_2941,In_291,In_975);
nand U2942 (N_2942,In_916,In_814);
nor U2943 (N_2943,In_86,In_265);
and U2944 (N_2944,In_265,In_790);
nand U2945 (N_2945,In_529,In_65);
or U2946 (N_2946,In_993,In_851);
nand U2947 (N_2947,In_778,In_929);
nor U2948 (N_2948,In_136,In_597);
nor U2949 (N_2949,In_141,In_272);
or U2950 (N_2950,In_350,In_865);
nand U2951 (N_2951,In_311,In_809);
and U2952 (N_2952,In_955,In_845);
nand U2953 (N_2953,In_985,In_48);
or U2954 (N_2954,In_191,In_852);
or U2955 (N_2955,In_508,In_530);
or U2956 (N_2956,In_81,In_151);
and U2957 (N_2957,In_958,In_815);
nand U2958 (N_2958,In_923,In_972);
or U2959 (N_2959,In_641,In_161);
nor U2960 (N_2960,In_141,In_547);
and U2961 (N_2961,In_273,In_94);
or U2962 (N_2962,In_133,In_61);
or U2963 (N_2963,In_235,In_695);
nand U2964 (N_2964,In_348,In_829);
and U2965 (N_2965,In_722,In_186);
or U2966 (N_2966,In_897,In_303);
or U2967 (N_2967,In_642,In_720);
nand U2968 (N_2968,In_987,In_596);
nor U2969 (N_2969,In_45,In_352);
or U2970 (N_2970,In_717,In_396);
or U2971 (N_2971,In_742,In_525);
and U2972 (N_2972,In_289,In_679);
and U2973 (N_2973,In_235,In_552);
nor U2974 (N_2974,In_48,In_521);
nor U2975 (N_2975,In_153,In_937);
nor U2976 (N_2976,In_920,In_565);
and U2977 (N_2977,In_213,In_548);
nor U2978 (N_2978,In_165,In_894);
nand U2979 (N_2979,In_407,In_541);
nand U2980 (N_2980,In_886,In_983);
nand U2981 (N_2981,In_523,In_366);
or U2982 (N_2982,In_0,In_408);
nor U2983 (N_2983,In_971,In_534);
or U2984 (N_2984,In_683,In_738);
or U2985 (N_2985,In_783,In_766);
or U2986 (N_2986,In_833,In_416);
nor U2987 (N_2987,In_25,In_719);
and U2988 (N_2988,In_673,In_12);
nand U2989 (N_2989,In_793,In_384);
nor U2990 (N_2990,In_183,In_698);
nor U2991 (N_2991,In_923,In_167);
or U2992 (N_2992,In_557,In_858);
nand U2993 (N_2993,In_985,In_367);
nand U2994 (N_2994,In_367,In_468);
or U2995 (N_2995,In_88,In_802);
nand U2996 (N_2996,In_908,In_301);
nand U2997 (N_2997,In_800,In_193);
nor U2998 (N_2998,In_562,In_280);
nand U2999 (N_2999,In_727,In_793);
or U3000 (N_3000,In_140,In_264);
and U3001 (N_3001,In_385,In_107);
nor U3002 (N_3002,In_270,In_662);
nand U3003 (N_3003,In_534,In_55);
nor U3004 (N_3004,In_562,In_691);
nor U3005 (N_3005,In_896,In_591);
or U3006 (N_3006,In_607,In_474);
and U3007 (N_3007,In_442,In_292);
and U3008 (N_3008,In_207,In_973);
nor U3009 (N_3009,In_220,In_183);
nor U3010 (N_3010,In_113,In_270);
or U3011 (N_3011,In_605,In_769);
or U3012 (N_3012,In_176,In_75);
nand U3013 (N_3013,In_985,In_672);
nand U3014 (N_3014,In_153,In_22);
and U3015 (N_3015,In_564,In_198);
nand U3016 (N_3016,In_77,In_737);
nor U3017 (N_3017,In_992,In_523);
nand U3018 (N_3018,In_109,In_990);
and U3019 (N_3019,In_194,In_588);
nor U3020 (N_3020,In_618,In_285);
nor U3021 (N_3021,In_88,In_153);
nand U3022 (N_3022,In_293,In_507);
and U3023 (N_3023,In_426,In_995);
nand U3024 (N_3024,In_642,In_509);
nor U3025 (N_3025,In_789,In_614);
nor U3026 (N_3026,In_136,In_580);
and U3027 (N_3027,In_325,In_705);
and U3028 (N_3028,In_106,In_322);
and U3029 (N_3029,In_78,In_616);
or U3030 (N_3030,In_24,In_129);
nor U3031 (N_3031,In_801,In_57);
or U3032 (N_3032,In_535,In_104);
and U3033 (N_3033,In_253,In_612);
nor U3034 (N_3034,In_486,In_982);
and U3035 (N_3035,In_650,In_198);
nor U3036 (N_3036,In_53,In_92);
and U3037 (N_3037,In_170,In_479);
and U3038 (N_3038,In_614,In_208);
nand U3039 (N_3039,In_288,In_15);
and U3040 (N_3040,In_348,In_180);
nand U3041 (N_3041,In_209,In_198);
nor U3042 (N_3042,In_192,In_941);
or U3043 (N_3043,In_504,In_24);
and U3044 (N_3044,In_931,In_423);
or U3045 (N_3045,In_593,In_472);
and U3046 (N_3046,In_435,In_5);
or U3047 (N_3047,In_252,In_407);
and U3048 (N_3048,In_659,In_419);
and U3049 (N_3049,In_249,In_429);
nor U3050 (N_3050,In_38,In_354);
or U3051 (N_3051,In_572,In_868);
nand U3052 (N_3052,In_593,In_486);
and U3053 (N_3053,In_376,In_955);
or U3054 (N_3054,In_30,In_430);
and U3055 (N_3055,In_504,In_10);
nor U3056 (N_3056,In_810,In_111);
or U3057 (N_3057,In_499,In_802);
and U3058 (N_3058,In_264,In_401);
or U3059 (N_3059,In_462,In_100);
or U3060 (N_3060,In_433,In_242);
or U3061 (N_3061,In_585,In_982);
and U3062 (N_3062,In_34,In_269);
and U3063 (N_3063,In_734,In_413);
and U3064 (N_3064,In_390,In_459);
nand U3065 (N_3065,In_943,In_804);
nor U3066 (N_3066,In_124,In_621);
nor U3067 (N_3067,In_34,In_79);
nand U3068 (N_3068,In_688,In_385);
or U3069 (N_3069,In_256,In_636);
nor U3070 (N_3070,In_428,In_414);
and U3071 (N_3071,In_151,In_331);
or U3072 (N_3072,In_339,In_66);
and U3073 (N_3073,In_246,In_725);
nand U3074 (N_3074,In_705,In_20);
or U3075 (N_3075,In_284,In_336);
nor U3076 (N_3076,In_813,In_547);
and U3077 (N_3077,In_186,In_740);
and U3078 (N_3078,In_214,In_705);
and U3079 (N_3079,In_245,In_166);
or U3080 (N_3080,In_640,In_506);
nor U3081 (N_3081,In_657,In_80);
and U3082 (N_3082,In_717,In_483);
nor U3083 (N_3083,In_686,In_625);
nand U3084 (N_3084,In_449,In_393);
or U3085 (N_3085,In_206,In_73);
nand U3086 (N_3086,In_136,In_699);
or U3087 (N_3087,In_716,In_361);
nand U3088 (N_3088,In_304,In_121);
nor U3089 (N_3089,In_495,In_658);
nand U3090 (N_3090,In_497,In_389);
or U3091 (N_3091,In_322,In_498);
xor U3092 (N_3092,In_101,In_443);
nor U3093 (N_3093,In_677,In_739);
and U3094 (N_3094,In_528,In_847);
nor U3095 (N_3095,In_714,In_490);
and U3096 (N_3096,In_927,In_996);
and U3097 (N_3097,In_721,In_866);
and U3098 (N_3098,In_415,In_649);
nor U3099 (N_3099,In_886,In_597);
nor U3100 (N_3100,In_589,In_629);
nor U3101 (N_3101,In_188,In_343);
nor U3102 (N_3102,In_630,In_296);
and U3103 (N_3103,In_306,In_893);
nor U3104 (N_3104,In_418,In_409);
or U3105 (N_3105,In_453,In_391);
nand U3106 (N_3106,In_666,In_218);
and U3107 (N_3107,In_895,In_527);
or U3108 (N_3108,In_743,In_26);
nor U3109 (N_3109,In_979,In_159);
nand U3110 (N_3110,In_654,In_198);
nor U3111 (N_3111,In_433,In_794);
nand U3112 (N_3112,In_531,In_257);
and U3113 (N_3113,In_331,In_666);
and U3114 (N_3114,In_947,In_286);
or U3115 (N_3115,In_847,In_561);
nand U3116 (N_3116,In_960,In_373);
or U3117 (N_3117,In_983,In_329);
and U3118 (N_3118,In_312,In_160);
or U3119 (N_3119,In_758,In_608);
nand U3120 (N_3120,In_355,In_644);
nand U3121 (N_3121,In_818,In_192);
and U3122 (N_3122,In_944,In_859);
and U3123 (N_3123,In_85,In_535);
nand U3124 (N_3124,In_137,In_738);
or U3125 (N_3125,In_719,In_662);
nand U3126 (N_3126,In_422,In_723);
or U3127 (N_3127,In_627,In_115);
xor U3128 (N_3128,In_563,In_617);
nand U3129 (N_3129,In_473,In_639);
or U3130 (N_3130,In_43,In_54);
or U3131 (N_3131,In_997,In_415);
nor U3132 (N_3132,In_964,In_236);
and U3133 (N_3133,In_603,In_536);
and U3134 (N_3134,In_156,In_99);
nor U3135 (N_3135,In_446,In_890);
nand U3136 (N_3136,In_47,In_503);
or U3137 (N_3137,In_688,In_50);
or U3138 (N_3138,In_760,In_204);
nor U3139 (N_3139,In_310,In_616);
nand U3140 (N_3140,In_850,In_617);
and U3141 (N_3141,In_746,In_789);
nor U3142 (N_3142,In_61,In_126);
or U3143 (N_3143,In_559,In_484);
nor U3144 (N_3144,In_953,In_689);
or U3145 (N_3145,In_941,In_666);
and U3146 (N_3146,In_86,In_12);
xor U3147 (N_3147,In_43,In_160);
or U3148 (N_3148,In_697,In_473);
or U3149 (N_3149,In_47,In_207);
nand U3150 (N_3150,In_577,In_104);
and U3151 (N_3151,In_963,In_245);
and U3152 (N_3152,In_29,In_433);
or U3153 (N_3153,In_518,In_109);
and U3154 (N_3154,In_491,In_610);
and U3155 (N_3155,In_906,In_262);
nor U3156 (N_3156,In_843,In_84);
and U3157 (N_3157,In_277,In_525);
nand U3158 (N_3158,In_562,In_801);
and U3159 (N_3159,In_955,In_141);
or U3160 (N_3160,In_841,In_883);
nor U3161 (N_3161,In_56,In_186);
nor U3162 (N_3162,In_90,In_437);
or U3163 (N_3163,In_817,In_321);
nand U3164 (N_3164,In_991,In_607);
nand U3165 (N_3165,In_964,In_461);
or U3166 (N_3166,In_212,In_324);
or U3167 (N_3167,In_521,In_8);
nand U3168 (N_3168,In_126,In_206);
nand U3169 (N_3169,In_70,In_742);
nor U3170 (N_3170,In_836,In_980);
or U3171 (N_3171,In_539,In_888);
or U3172 (N_3172,In_506,In_294);
xnor U3173 (N_3173,In_565,In_840);
nor U3174 (N_3174,In_113,In_198);
nand U3175 (N_3175,In_278,In_62);
and U3176 (N_3176,In_437,In_154);
and U3177 (N_3177,In_701,In_387);
nand U3178 (N_3178,In_875,In_342);
or U3179 (N_3179,In_862,In_978);
nor U3180 (N_3180,In_159,In_522);
and U3181 (N_3181,In_755,In_551);
nor U3182 (N_3182,In_665,In_459);
and U3183 (N_3183,In_613,In_359);
nand U3184 (N_3184,In_319,In_894);
and U3185 (N_3185,In_233,In_300);
xor U3186 (N_3186,In_196,In_787);
or U3187 (N_3187,In_975,In_882);
nor U3188 (N_3188,In_185,In_249);
nor U3189 (N_3189,In_422,In_470);
nand U3190 (N_3190,In_220,In_200);
nor U3191 (N_3191,In_507,In_329);
nand U3192 (N_3192,In_762,In_873);
nor U3193 (N_3193,In_37,In_739);
or U3194 (N_3194,In_762,In_20);
nand U3195 (N_3195,In_449,In_568);
and U3196 (N_3196,In_487,In_325);
nand U3197 (N_3197,In_984,In_254);
or U3198 (N_3198,In_125,In_925);
nor U3199 (N_3199,In_671,In_241);
nand U3200 (N_3200,In_62,In_389);
nor U3201 (N_3201,In_275,In_213);
nor U3202 (N_3202,In_635,In_104);
nand U3203 (N_3203,In_824,In_328);
or U3204 (N_3204,In_320,In_765);
nor U3205 (N_3205,In_106,In_950);
or U3206 (N_3206,In_555,In_386);
nand U3207 (N_3207,In_318,In_101);
nor U3208 (N_3208,In_62,In_505);
or U3209 (N_3209,In_449,In_384);
and U3210 (N_3210,In_430,In_423);
or U3211 (N_3211,In_261,In_181);
or U3212 (N_3212,In_9,In_722);
or U3213 (N_3213,In_184,In_646);
or U3214 (N_3214,In_364,In_52);
or U3215 (N_3215,In_176,In_538);
or U3216 (N_3216,In_285,In_871);
or U3217 (N_3217,In_783,In_230);
nor U3218 (N_3218,In_202,In_434);
nand U3219 (N_3219,In_775,In_266);
and U3220 (N_3220,In_562,In_439);
nor U3221 (N_3221,In_753,In_368);
nand U3222 (N_3222,In_22,In_971);
nor U3223 (N_3223,In_764,In_205);
and U3224 (N_3224,In_867,In_250);
or U3225 (N_3225,In_790,In_568);
and U3226 (N_3226,In_923,In_225);
nor U3227 (N_3227,In_956,In_381);
and U3228 (N_3228,In_624,In_570);
and U3229 (N_3229,In_615,In_726);
nand U3230 (N_3230,In_597,In_964);
nand U3231 (N_3231,In_656,In_366);
nor U3232 (N_3232,In_415,In_463);
nor U3233 (N_3233,In_258,In_433);
nor U3234 (N_3234,In_699,In_21);
xor U3235 (N_3235,In_864,In_169);
and U3236 (N_3236,In_372,In_361);
or U3237 (N_3237,In_330,In_314);
nor U3238 (N_3238,In_367,In_896);
nand U3239 (N_3239,In_0,In_383);
nand U3240 (N_3240,In_144,In_837);
nor U3241 (N_3241,In_16,In_786);
and U3242 (N_3242,In_222,In_461);
or U3243 (N_3243,In_862,In_485);
nor U3244 (N_3244,In_673,In_987);
and U3245 (N_3245,In_39,In_576);
nand U3246 (N_3246,In_954,In_491);
or U3247 (N_3247,In_836,In_117);
or U3248 (N_3248,In_330,In_773);
nor U3249 (N_3249,In_853,In_689);
nand U3250 (N_3250,In_431,In_691);
and U3251 (N_3251,In_706,In_240);
nand U3252 (N_3252,In_471,In_805);
nor U3253 (N_3253,In_631,In_722);
nand U3254 (N_3254,In_389,In_763);
and U3255 (N_3255,In_555,In_693);
or U3256 (N_3256,In_287,In_827);
nand U3257 (N_3257,In_422,In_861);
or U3258 (N_3258,In_7,In_306);
nand U3259 (N_3259,In_685,In_165);
or U3260 (N_3260,In_290,In_857);
and U3261 (N_3261,In_910,In_779);
or U3262 (N_3262,In_772,In_537);
nand U3263 (N_3263,In_963,In_589);
and U3264 (N_3264,In_738,In_695);
nor U3265 (N_3265,In_508,In_700);
or U3266 (N_3266,In_371,In_167);
or U3267 (N_3267,In_241,In_922);
nand U3268 (N_3268,In_92,In_398);
nand U3269 (N_3269,In_843,In_458);
nor U3270 (N_3270,In_219,In_441);
nand U3271 (N_3271,In_22,In_504);
and U3272 (N_3272,In_189,In_105);
nor U3273 (N_3273,In_377,In_193);
or U3274 (N_3274,In_898,In_49);
nand U3275 (N_3275,In_811,In_738);
and U3276 (N_3276,In_589,In_745);
or U3277 (N_3277,In_447,In_903);
or U3278 (N_3278,In_626,In_981);
and U3279 (N_3279,In_11,In_204);
or U3280 (N_3280,In_331,In_147);
nor U3281 (N_3281,In_646,In_808);
nand U3282 (N_3282,In_318,In_464);
or U3283 (N_3283,In_493,In_235);
and U3284 (N_3284,In_927,In_155);
and U3285 (N_3285,In_414,In_187);
or U3286 (N_3286,In_13,In_725);
nor U3287 (N_3287,In_88,In_552);
nor U3288 (N_3288,In_490,In_968);
or U3289 (N_3289,In_266,In_914);
and U3290 (N_3290,In_785,In_573);
and U3291 (N_3291,In_568,In_206);
and U3292 (N_3292,In_37,In_858);
nor U3293 (N_3293,In_705,In_237);
nor U3294 (N_3294,In_138,In_278);
and U3295 (N_3295,In_511,In_100);
nand U3296 (N_3296,In_212,In_507);
or U3297 (N_3297,In_188,In_454);
xor U3298 (N_3298,In_195,In_489);
nor U3299 (N_3299,In_52,In_761);
nor U3300 (N_3300,In_66,In_74);
nand U3301 (N_3301,In_739,In_107);
and U3302 (N_3302,In_150,In_41);
nand U3303 (N_3303,In_738,In_530);
nand U3304 (N_3304,In_751,In_695);
nand U3305 (N_3305,In_875,In_393);
and U3306 (N_3306,In_493,In_943);
nor U3307 (N_3307,In_117,In_715);
nand U3308 (N_3308,In_395,In_814);
or U3309 (N_3309,In_234,In_378);
or U3310 (N_3310,In_942,In_781);
nand U3311 (N_3311,In_247,In_955);
nor U3312 (N_3312,In_169,In_881);
nor U3313 (N_3313,In_780,In_638);
nand U3314 (N_3314,In_113,In_116);
nor U3315 (N_3315,In_424,In_344);
and U3316 (N_3316,In_861,In_804);
or U3317 (N_3317,In_946,In_625);
nand U3318 (N_3318,In_375,In_782);
nor U3319 (N_3319,In_135,In_720);
or U3320 (N_3320,In_31,In_305);
nand U3321 (N_3321,In_760,In_61);
and U3322 (N_3322,In_383,In_858);
or U3323 (N_3323,In_955,In_652);
or U3324 (N_3324,In_814,In_857);
nand U3325 (N_3325,In_453,In_150);
nor U3326 (N_3326,In_753,In_211);
nand U3327 (N_3327,In_160,In_354);
nand U3328 (N_3328,In_473,In_36);
or U3329 (N_3329,In_444,In_749);
nand U3330 (N_3330,In_301,In_832);
nor U3331 (N_3331,In_304,In_557);
and U3332 (N_3332,In_938,In_573);
nor U3333 (N_3333,In_739,In_517);
nand U3334 (N_3334,In_579,In_611);
and U3335 (N_3335,In_518,In_376);
and U3336 (N_3336,In_601,In_937);
and U3337 (N_3337,In_102,In_313);
or U3338 (N_3338,In_63,In_459);
nor U3339 (N_3339,In_100,In_864);
and U3340 (N_3340,In_495,In_373);
and U3341 (N_3341,In_563,In_112);
nor U3342 (N_3342,In_857,In_906);
nor U3343 (N_3343,In_570,In_587);
nand U3344 (N_3344,In_188,In_417);
or U3345 (N_3345,In_433,In_800);
or U3346 (N_3346,In_610,In_108);
and U3347 (N_3347,In_143,In_423);
or U3348 (N_3348,In_110,In_163);
nand U3349 (N_3349,In_104,In_339);
nand U3350 (N_3350,In_900,In_216);
or U3351 (N_3351,In_125,In_237);
or U3352 (N_3352,In_809,In_990);
and U3353 (N_3353,In_950,In_246);
and U3354 (N_3354,In_994,In_400);
or U3355 (N_3355,In_271,In_387);
or U3356 (N_3356,In_870,In_721);
nor U3357 (N_3357,In_690,In_92);
or U3358 (N_3358,In_114,In_236);
nor U3359 (N_3359,In_237,In_153);
and U3360 (N_3360,In_232,In_51);
nor U3361 (N_3361,In_197,In_718);
or U3362 (N_3362,In_697,In_635);
nand U3363 (N_3363,In_497,In_858);
nor U3364 (N_3364,In_134,In_856);
or U3365 (N_3365,In_893,In_99);
and U3366 (N_3366,In_306,In_469);
or U3367 (N_3367,In_164,In_644);
nor U3368 (N_3368,In_668,In_605);
or U3369 (N_3369,In_627,In_90);
or U3370 (N_3370,In_103,In_134);
or U3371 (N_3371,In_640,In_766);
and U3372 (N_3372,In_875,In_336);
or U3373 (N_3373,In_968,In_397);
nor U3374 (N_3374,In_766,In_172);
or U3375 (N_3375,In_575,In_545);
and U3376 (N_3376,In_62,In_927);
nor U3377 (N_3377,In_826,In_78);
nand U3378 (N_3378,In_648,In_428);
and U3379 (N_3379,In_164,In_289);
and U3380 (N_3380,In_148,In_796);
or U3381 (N_3381,In_765,In_157);
and U3382 (N_3382,In_719,In_769);
nand U3383 (N_3383,In_284,In_312);
nor U3384 (N_3384,In_735,In_20);
and U3385 (N_3385,In_218,In_59);
nand U3386 (N_3386,In_15,In_326);
or U3387 (N_3387,In_699,In_239);
nand U3388 (N_3388,In_827,In_384);
and U3389 (N_3389,In_889,In_247);
nand U3390 (N_3390,In_653,In_742);
nor U3391 (N_3391,In_193,In_802);
nor U3392 (N_3392,In_535,In_341);
nor U3393 (N_3393,In_86,In_71);
nand U3394 (N_3394,In_798,In_387);
and U3395 (N_3395,In_486,In_188);
or U3396 (N_3396,In_426,In_464);
or U3397 (N_3397,In_421,In_260);
or U3398 (N_3398,In_959,In_997);
or U3399 (N_3399,In_978,In_629);
nand U3400 (N_3400,In_959,In_129);
nor U3401 (N_3401,In_87,In_830);
and U3402 (N_3402,In_561,In_478);
or U3403 (N_3403,In_465,In_109);
nor U3404 (N_3404,In_572,In_464);
and U3405 (N_3405,In_173,In_512);
nor U3406 (N_3406,In_705,In_523);
nand U3407 (N_3407,In_430,In_507);
nor U3408 (N_3408,In_103,In_232);
or U3409 (N_3409,In_77,In_141);
nand U3410 (N_3410,In_618,In_873);
or U3411 (N_3411,In_116,In_745);
nand U3412 (N_3412,In_374,In_37);
and U3413 (N_3413,In_988,In_819);
nor U3414 (N_3414,In_788,In_774);
and U3415 (N_3415,In_452,In_833);
nand U3416 (N_3416,In_355,In_550);
nor U3417 (N_3417,In_171,In_905);
and U3418 (N_3418,In_616,In_317);
nand U3419 (N_3419,In_772,In_528);
or U3420 (N_3420,In_600,In_940);
xor U3421 (N_3421,In_417,In_541);
and U3422 (N_3422,In_523,In_155);
and U3423 (N_3423,In_413,In_336);
nand U3424 (N_3424,In_834,In_821);
nor U3425 (N_3425,In_370,In_960);
and U3426 (N_3426,In_663,In_756);
nand U3427 (N_3427,In_641,In_706);
or U3428 (N_3428,In_431,In_605);
nor U3429 (N_3429,In_100,In_518);
nor U3430 (N_3430,In_789,In_16);
nand U3431 (N_3431,In_856,In_691);
or U3432 (N_3432,In_923,In_729);
nor U3433 (N_3433,In_774,In_893);
or U3434 (N_3434,In_247,In_484);
nand U3435 (N_3435,In_168,In_425);
nand U3436 (N_3436,In_172,In_115);
nand U3437 (N_3437,In_872,In_7);
nand U3438 (N_3438,In_239,In_943);
or U3439 (N_3439,In_504,In_377);
and U3440 (N_3440,In_826,In_112);
or U3441 (N_3441,In_269,In_669);
nand U3442 (N_3442,In_662,In_11);
nand U3443 (N_3443,In_956,In_709);
or U3444 (N_3444,In_677,In_49);
nand U3445 (N_3445,In_502,In_178);
nor U3446 (N_3446,In_521,In_681);
nand U3447 (N_3447,In_675,In_994);
nand U3448 (N_3448,In_754,In_527);
nand U3449 (N_3449,In_446,In_876);
nand U3450 (N_3450,In_371,In_915);
nor U3451 (N_3451,In_867,In_273);
nor U3452 (N_3452,In_390,In_288);
and U3453 (N_3453,In_179,In_464);
or U3454 (N_3454,In_191,In_653);
nand U3455 (N_3455,In_628,In_774);
and U3456 (N_3456,In_917,In_439);
nand U3457 (N_3457,In_575,In_81);
nor U3458 (N_3458,In_151,In_494);
and U3459 (N_3459,In_880,In_802);
nor U3460 (N_3460,In_824,In_941);
and U3461 (N_3461,In_37,In_528);
or U3462 (N_3462,In_254,In_154);
and U3463 (N_3463,In_902,In_739);
nand U3464 (N_3464,In_559,In_33);
nor U3465 (N_3465,In_260,In_980);
and U3466 (N_3466,In_958,In_33);
nand U3467 (N_3467,In_917,In_683);
or U3468 (N_3468,In_784,In_536);
or U3469 (N_3469,In_150,In_724);
or U3470 (N_3470,In_491,In_382);
nand U3471 (N_3471,In_333,In_873);
and U3472 (N_3472,In_608,In_915);
nor U3473 (N_3473,In_923,In_545);
nor U3474 (N_3474,In_319,In_211);
nor U3475 (N_3475,In_671,In_956);
or U3476 (N_3476,In_509,In_480);
nor U3477 (N_3477,In_292,In_588);
nand U3478 (N_3478,In_748,In_737);
nor U3479 (N_3479,In_155,In_157);
nor U3480 (N_3480,In_955,In_537);
or U3481 (N_3481,In_879,In_902);
nor U3482 (N_3482,In_466,In_788);
nor U3483 (N_3483,In_376,In_424);
nor U3484 (N_3484,In_803,In_764);
nand U3485 (N_3485,In_397,In_693);
or U3486 (N_3486,In_840,In_242);
or U3487 (N_3487,In_451,In_588);
and U3488 (N_3488,In_160,In_878);
nor U3489 (N_3489,In_150,In_527);
nand U3490 (N_3490,In_374,In_59);
xnor U3491 (N_3491,In_961,In_37);
or U3492 (N_3492,In_205,In_722);
or U3493 (N_3493,In_230,In_983);
and U3494 (N_3494,In_757,In_639);
and U3495 (N_3495,In_805,In_803);
nor U3496 (N_3496,In_813,In_165);
nor U3497 (N_3497,In_821,In_621);
nor U3498 (N_3498,In_775,In_477);
or U3499 (N_3499,In_756,In_648);
or U3500 (N_3500,In_432,In_855);
and U3501 (N_3501,In_775,In_306);
or U3502 (N_3502,In_751,In_614);
or U3503 (N_3503,In_167,In_765);
nand U3504 (N_3504,In_406,In_720);
and U3505 (N_3505,In_769,In_165);
and U3506 (N_3506,In_111,In_595);
and U3507 (N_3507,In_323,In_622);
and U3508 (N_3508,In_709,In_686);
or U3509 (N_3509,In_299,In_385);
nand U3510 (N_3510,In_174,In_634);
nand U3511 (N_3511,In_13,In_887);
nand U3512 (N_3512,In_129,In_942);
or U3513 (N_3513,In_447,In_810);
nand U3514 (N_3514,In_527,In_814);
or U3515 (N_3515,In_40,In_274);
or U3516 (N_3516,In_614,In_58);
or U3517 (N_3517,In_79,In_513);
nor U3518 (N_3518,In_708,In_409);
or U3519 (N_3519,In_473,In_972);
and U3520 (N_3520,In_490,In_452);
or U3521 (N_3521,In_320,In_96);
nor U3522 (N_3522,In_775,In_45);
or U3523 (N_3523,In_315,In_441);
nor U3524 (N_3524,In_115,In_470);
nand U3525 (N_3525,In_416,In_921);
nor U3526 (N_3526,In_897,In_305);
and U3527 (N_3527,In_658,In_755);
nand U3528 (N_3528,In_97,In_308);
nor U3529 (N_3529,In_597,In_341);
nor U3530 (N_3530,In_913,In_316);
and U3531 (N_3531,In_320,In_216);
nor U3532 (N_3532,In_473,In_793);
nor U3533 (N_3533,In_295,In_235);
nor U3534 (N_3534,In_688,In_444);
nand U3535 (N_3535,In_722,In_719);
and U3536 (N_3536,In_763,In_100);
or U3537 (N_3537,In_385,In_886);
nor U3538 (N_3538,In_420,In_413);
nor U3539 (N_3539,In_566,In_136);
or U3540 (N_3540,In_299,In_731);
nand U3541 (N_3541,In_715,In_739);
nand U3542 (N_3542,In_246,In_839);
and U3543 (N_3543,In_411,In_122);
nand U3544 (N_3544,In_905,In_9);
nand U3545 (N_3545,In_177,In_324);
nand U3546 (N_3546,In_77,In_44);
nor U3547 (N_3547,In_941,In_870);
and U3548 (N_3548,In_758,In_309);
and U3549 (N_3549,In_736,In_716);
or U3550 (N_3550,In_416,In_870);
nor U3551 (N_3551,In_916,In_784);
nor U3552 (N_3552,In_134,In_291);
nor U3553 (N_3553,In_980,In_112);
nor U3554 (N_3554,In_181,In_777);
or U3555 (N_3555,In_715,In_589);
or U3556 (N_3556,In_266,In_172);
and U3557 (N_3557,In_673,In_605);
nand U3558 (N_3558,In_670,In_871);
and U3559 (N_3559,In_922,In_418);
xor U3560 (N_3560,In_28,In_480);
or U3561 (N_3561,In_34,In_3);
nor U3562 (N_3562,In_732,In_597);
and U3563 (N_3563,In_122,In_689);
or U3564 (N_3564,In_914,In_234);
or U3565 (N_3565,In_829,In_473);
nor U3566 (N_3566,In_213,In_680);
nand U3567 (N_3567,In_935,In_235);
nor U3568 (N_3568,In_644,In_4);
or U3569 (N_3569,In_744,In_265);
nor U3570 (N_3570,In_680,In_225);
nand U3571 (N_3571,In_629,In_55);
or U3572 (N_3572,In_89,In_680);
or U3573 (N_3573,In_608,In_329);
nor U3574 (N_3574,In_99,In_255);
and U3575 (N_3575,In_539,In_88);
and U3576 (N_3576,In_459,In_616);
nand U3577 (N_3577,In_984,In_731);
nor U3578 (N_3578,In_433,In_776);
nor U3579 (N_3579,In_422,In_760);
or U3580 (N_3580,In_410,In_753);
and U3581 (N_3581,In_721,In_883);
or U3582 (N_3582,In_632,In_436);
nor U3583 (N_3583,In_720,In_363);
and U3584 (N_3584,In_20,In_437);
and U3585 (N_3585,In_476,In_660);
or U3586 (N_3586,In_244,In_495);
nor U3587 (N_3587,In_319,In_529);
or U3588 (N_3588,In_780,In_994);
and U3589 (N_3589,In_579,In_71);
nor U3590 (N_3590,In_589,In_468);
or U3591 (N_3591,In_537,In_180);
nand U3592 (N_3592,In_981,In_450);
or U3593 (N_3593,In_194,In_237);
nand U3594 (N_3594,In_153,In_987);
or U3595 (N_3595,In_405,In_444);
or U3596 (N_3596,In_437,In_655);
nor U3597 (N_3597,In_799,In_554);
or U3598 (N_3598,In_119,In_290);
nor U3599 (N_3599,In_987,In_813);
nand U3600 (N_3600,In_184,In_773);
or U3601 (N_3601,In_465,In_217);
nor U3602 (N_3602,In_508,In_872);
and U3603 (N_3603,In_679,In_383);
or U3604 (N_3604,In_338,In_737);
nand U3605 (N_3605,In_10,In_642);
and U3606 (N_3606,In_81,In_923);
or U3607 (N_3607,In_359,In_125);
and U3608 (N_3608,In_471,In_166);
nor U3609 (N_3609,In_171,In_166);
nand U3610 (N_3610,In_603,In_170);
and U3611 (N_3611,In_617,In_847);
and U3612 (N_3612,In_441,In_866);
and U3613 (N_3613,In_147,In_762);
nor U3614 (N_3614,In_532,In_491);
nor U3615 (N_3615,In_525,In_314);
nand U3616 (N_3616,In_186,In_697);
or U3617 (N_3617,In_626,In_727);
and U3618 (N_3618,In_317,In_144);
nor U3619 (N_3619,In_909,In_942);
nand U3620 (N_3620,In_355,In_738);
nor U3621 (N_3621,In_470,In_254);
nand U3622 (N_3622,In_219,In_959);
or U3623 (N_3623,In_73,In_286);
or U3624 (N_3624,In_305,In_960);
xnor U3625 (N_3625,In_81,In_852);
nand U3626 (N_3626,In_876,In_502);
or U3627 (N_3627,In_557,In_679);
or U3628 (N_3628,In_610,In_318);
nand U3629 (N_3629,In_300,In_549);
nor U3630 (N_3630,In_119,In_712);
nand U3631 (N_3631,In_392,In_962);
and U3632 (N_3632,In_436,In_842);
or U3633 (N_3633,In_566,In_683);
nor U3634 (N_3634,In_213,In_570);
nor U3635 (N_3635,In_291,In_162);
and U3636 (N_3636,In_220,In_33);
nor U3637 (N_3637,In_573,In_505);
or U3638 (N_3638,In_701,In_770);
nor U3639 (N_3639,In_987,In_934);
or U3640 (N_3640,In_285,In_435);
or U3641 (N_3641,In_855,In_695);
and U3642 (N_3642,In_826,In_669);
and U3643 (N_3643,In_573,In_854);
and U3644 (N_3644,In_680,In_148);
and U3645 (N_3645,In_652,In_684);
nor U3646 (N_3646,In_3,In_16);
and U3647 (N_3647,In_86,In_621);
and U3648 (N_3648,In_190,In_280);
or U3649 (N_3649,In_84,In_177);
nand U3650 (N_3650,In_403,In_701);
and U3651 (N_3651,In_16,In_740);
and U3652 (N_3652,In_309,In_264);
xor U3653 (N_3653,In_48,In_685);
nor U3654 (N_3654,In_328,In_307);
nand U3655 (N_3655,In_565,In_14);
nor U3656 (N_3656,In_108,In_585);
nor U3657 (N_3657,In_587,In_365);
or U3658 (N_3658,In_214,In_507);
and U3659 (N_3659,In_96,In_432);
or U3660 (N_3660,In_484,In_987);
nand U3661 (N_3661,In_204,In_88);
xor U3662 (N_3662,In_483,In_949);
or U3663 (N_3663,In_388,In_931);
nor U3664 (N_3664,In_262,In_831);
nor U3665 (N_3665,In_161,In_943);
nor U3666 (N_3666,In_453,In_244);
nand U3667 (N_3667,In_769,In_819);
nand U3668 (N_3668,In_243,In_434);
nand U3669 (N_3669,In_5,In_348);
or U3670 (N_3670,In_550,In_7);
and U3671 (N_3671,In_311,In_469);
or U3672 (N_3672,In_28,In_92);
nor U3673 (N_3673,In_305,In_481);
nor U3674 (N_3674,In_909,In_727);
and U3675 (N_3675,In_248,In_617);
or U3676 (N_3676,In_95,In_476);
and U3677 (N_3677,In_883,In_497);
and U3678 (N_3678,In_548,In_734);
or U3679 (N_3679,In_86,In_899);
nand U3680 (N_3680,In_466,In_9);
and U3681 (N_3681,In_726,In_700);
nor U3682 (N_3682,In_747,In_445);
or U3683 (N_3683,In_875,In_752);
nor U3684 (N_3684,In_903,In_969);
nand U3685 (N_3685,In_472,In_348);
nand U3686 (N_3686,In_678,In_590);
or U3687 (N_3687,In_53,In_438);
nor U3688 (N_3688,In_596,In_108);
nand U3689 (N_3689,In_7,In_824);
nand U3690 (N_3690,In_666,In_290);
and U3691 (N_3691,In_108,In_821);
nor U3692 (N_3692,In_99,In_102);
nand U3693 (N_3693,In_165,In_986);
nor U3694 (N_3694,In_286,In_696);
nor U3695 (N_3695,In_799,In_7);
nor U3696 (N_3696,In_345,In_696);
nand U3697 (N_3697,In_380,In_526);
nand U3698 (N_3698,In_796,In_26);
and U3699 (N_3699,In_695,In_598);
and U3700 (N_3700,In_353,In_153);
nand U3701 (N_3701,In_832,In_124);
nand U3702 (N_3702,In_284,In_14);
or U3703 (N_3703,In_612,In_451);
or U3704 (N_3704,In_690,In_854);
and U3705 (N_3705,In_96,In_796);
and U3706 (N_3706,In_648,In_790);
nand U3707 (N_3707,In_890,In_583);
nor U3708 (N_3708,In_992,In_348);
nor U3709 (N_3709,In_907,In_485);
nand U3710 (N_3710,In_495,In_585);
nand U3711 (N_3711,In_283,In_580);
and U3712 (N_3712,In_241,In_646);
nand U3713 (N_3713,In_101,In_209);
nand U3714 (N_3714,In_626,In_587);
nor U3715 (N_3715,In_974,In_979);
and U3716 (N_3716,In_106,In_23);
nor U3717 (N_3717,In_611,In_834);
or U3718 (N_3718,In_835,In_498);
or U3719 (N_3719,In_410,In_148);
nor U3720 (N_3720,In_49,In_345);
or U3721 (N_3721,In_390,In_678);
and U3722 (N_3722,In_310,In_483);
nor U3723 (N_3723,In_99,In_472);
and U3724 (N_3724,In_365,In_327);
or U3725 (N_3725,In_101,In_279);
and U3726 (N_3726,In_325,In_265);
or U3727 (N_3727,In_264,In_789);
or U3728 (N_3728,In_576,In_113);
nand U3729 (N_3729,In_185,In_337);
nand U3730 (N_3730,In_982,In_809);
nor U3731 (N_3731,In_809,In_471);
and U3732 (N_3732,In_669,In_612);
or U3733 (N_3733,In_654,In_139);
and U3734 (N_3734,In_114,In_910);
or U3735 (N_3735,In_107,In_329);
or U3736 (N_3736,In_811,In_506);
nand U3737 (N_3737,In_983,In_204);
nand U3738 (N_3738,In_465,In_663);
and U3739 (N_3739,In_79,In_664);
or U3740 (N_3740,In_12,In_153);
and U3741 (N_3741,In_687,In_705);
nand U3742 (N_3742,In_720,In_970);
nand U3743 (N_3743,In_336,In_829);
or U3744 (N_3744,In_77,In_339);
nor U3745 (N_3745,In_536,In_903);
and U3746 (N_3746,In_448,In_734);
nor U3747 (N_3747,In_460,In_804);
or U3748 (N_3748,In_211,In_782);
or U3749 (N_3749,In_15,In_420);
and U3750 (N_3750,In_262,In_216);
or U3751 (N_3751,In_840,In_449);
and U3752 (N_3752,In_169,In_979);
or U3753 (N_3753,In_384,In_101);
nand U3754 (N_3754,In_566,In_547);
or U3755 (N_3755,In_660,In_417);
nor U3756 (N_3756,In_460,In_763);
nor U3757 (N_3757,In_959,In_838);
or U3758 (N_3758,In_978,In_119);
nor U3759 (N_3759,In_887,In_768);
and U3760 (N_3760,In_492,In_375);
nor U3761 (N_3761,In_891,In_203);
and U3762 (N_3762,In_581,In_78);
nor U3763 (N_3763,In_303,In_951);
nand U3764 (N_3764,In_169,In_822);
or U3765 (N_3765,In_219,In_696);
or U3766 (N_3766,In_403,In_725);
nor U3767 (N_3767,In_848,In_736);
and U3768 (N_3768,In_253,In_992);
or U3769 (N_3769,In_208,In_891);
and U3770 (N_3770,In_142,In_557);
nand U3771 (N_3771,In_896,In_512);
nand U3772 (N_3772,In_193,In_812);
nor U3773 (N_3773,In_465,In_317);
or U3774 (N_3774,In_734,In_15);
or U3775 (N_3775,In_57,In_884);
and U3776 (N_3776,In_787,In_808);
nand U3777 (N_3777,In_780,In_91);
and U3778 (N_3778,In_639,In_412);
or U3779 (N_3779,In_578,In_244);
and U3780 (N_3780,In_998,In_346);
nand U3781 (N_3781,In_923,In_599);
or U3782 (N_3782,In_773,In_402);
nand U3783 (N_3783,In_961,In_943);
and U3784 (N_3784,In_366,In_116);
and U3785 (N_3785,In_409,In_925);
nor U3786 (N_3786,In_627,In_861);
nor U3787 (N_3787,In_272,In_349);
or U3788 (N_3788,In_527,In_532);
nor U3789 (N_3789,In_202,In_660);
or U3790 (N_3790,In_813,In_401);
nand U3791 (N_3791,In_244,In_860);
nor U3792 (N_3792,In_564,In_287);
and U3793 (N_3793,In_647,In_93);
xor U3794 (N_3794,In_594,In_52);
and U3795 (N_3795,In_447,In_758);
nand U3796 (N_3796,In_893,In_901);
nand U3797 (N_3797,In_636,In_763);
nand U3798 (N_3798,In_943,In_176);
nand U3799 (N_3799,In_841,In_633);
nor U3800 (N_3800,In_94,In_297);
nor U3801 (N_3801,In_127,In_692);
or U3802 (N_3802,In_605,In_707);
or U3803 (N_3803,In_268,In_154);
and U3804 (N_3804,In_102,In_474);
nor U3805 (N_3805,In_36,In_490);
nand U3806 (N_3806,In_419,In_684);
nor U3807 (N_3807,In_797,In_317);
nand U3808 (N_3808,In_954,In_776);
and U3809 (N_3809,In_559,In_738);
nand U3810 (N_3810,In_677,In_762);
or U3811 (N_3811,In_820,In_869);
nand U3812 (N_3812,In_227,In_916);
nor U3813 (N_3813,In_935,In_4);
nor U3814 (N_3814,In_504,In_823);
and U3815 (N_3815,In_258,In_852);
and U3816 (N_3816,In_886,In_444);
nand U3817 (N_3817,In_298,In_877);
nor U3818 (N_3818,In_581,In_34);
or U3819 (N_3819,In_20,In_741);
nand U3820 (N_3820,In_23,In_936);
or U3821 (N_3821,In_984,In_457);
and U3822 (N_3822,In_641,In_545);
and U3823 (N_3823,In_515,In_85);
or U3824 (N_3824,In_644,In_256);
and U3825 (N_3825,In_150,In_777);
nor U3826 (N_3826,In_627,In_561);
nand U3827 (N_3827,In_904,In_934);
and U3828 (N_3828,In_150,In_893);
nor U3829 (N_3829,In_901,In_167);
nand U3830 (N_3830,In_594,In_714);
or U3831 (N_3831,In_238,In_101);
or U3832 (N_3832,In_886,In_102);
nand U3833 (N_3833,In_688,In_669);
nor U3834 (N_3834,In_138,In_328);
and U3835 (N_3835,In_112,In_414);
and U3836 (N_3836,In_734,In_731);
nand U3837 (N_3837,In_644,In_145);
nand U3838 (N_3838,In_735,In_738);
and U3839 (N_3839,In_760,In_189);
nand U3840 (N_3840,In_349,In_981);
or U3841 (N_3841,In_783,In_453);
and U3842 (N_3842,In_767,In_608);
nor U3843 (N_3843,In_650,In_853);
or U3844 (N_3844,In_754,In_831);
and U3845 (N_3845,In_925,In_998);
nand U3846 (N_3846,In_399,In_582);
and U3847 (N_3847,In_47,In_843);
and U3848 (N_3848,In_682,In_530);
and U3849 (N_3849,In_903,In_325);
and U3850 (N_3850,In_288,In_87);
nor U3851 (N_3851,In_421,In_487);
nor U3852 (N_3852,In_782,In_175);
nand U3853 (N_3853,In_83,In_528);
nor U3854 (N_3854,In_907,In_38);
nor U3855 (N_3855,In_172,In_637);
nor U3856 (N_3856,In_515,In_369);
nor U3857 (N_3857,In_578,In_548);
and U3858 (N_3858,In_886,In_795);
or U3859 (N_3859,In_924,In_620);
and U3860 (N_3860,In_22,In_571);
nand U3861 (N_3861,In_781,In_640);
and U3862 (N_3862,In_337,In_610);
and U3863 (N_3863,In_228,In_110);
nand U3864 (N_3864,In_746,In_859);
or U3865 (N_3865,In_747,In_942);
and U3866 (N_3866,In_491,In_798);
and U3867 (N_3867,In_859,In_101);
and U3868 (N_3868,In_828,In_75);
nand U3869 (N_3869,In_659,In_40);
nor U3870 (N_3870,In_361,In_527);
and U3871 (N_3871,In_940,In_91);
nor U3872 (N_3872,In_116,In_770);
nand U3873 (N_3873,In_238,In_706);
nor U3874 (N_3874,In_525,In_867);
nand U3875 (N_3875,In_356,In_770);
or U3876 (N_3876,In_895,In_994);
or U3877 (N_3877,In_582,In_304);
or U3878 (N_3878,In_974,In_470);
nor U3879 (N_3879,In_11,In_400);
or U3880 (N_3880,In_983,In_975);
or U3881 (N_3881,In_814,In_414);
nand U3882 (N_3882,In_204,In_588);
nor U3883 (N_3883,In_113,In_135);
and U3884 (N_3884,In_133,In_413);
or U3885 (N_3885,In_443,In_909);
nor U3886 (N_3886,In_234,In_992);
and U3887 (N_3887,In_463,In_431);
and U3888 (N_3888,In_719,In_948);
or U3889 (N_3889,In_495,In_470);
nand U3890 (N_3890,In_470,In_600);
and U3891 (N_3891,In_220,In_11);
and U3892 (N_3892,In_873,In_890);
nor U3893 (N_3893,In_306,In_474);
nand U3894 (N_3894,In_430,In_395);
nor U3895 (N_3895,In_13,In_605);
nor U3896 (N_3896,In_866,In_977);
and U3897 (N_3897,In_136,In_364);
and U3898 (N_3898,In_79,In_863);
nand U3899 (N_3899,In_186,In_625);
nand U3900 (N_3900,In_256,In_51);
nor U3901 (N_3901,In_686,In_809);
and U3902 (N_3902,In_77,In_504);
and U3903 (N_3903,In_783,In_7);
or U3904 (N_3904,In_793,In_927);
nor U3905 (N_3905,In_343,In_532);
nand U3906 (N_3906,In_119,In_564);
and U3907 (N_3907,In_158,In_531);
nand U3908 (N_3908,In_893,In_123);
or U3909 (N_3909,In_825,In_600);
nand U3910 (N_3910,In_422,In_335);
nor U3911 (N_3911,In_624,In_697);
and U3912 (N_3912,In_604,In_470);
and U3913 (N_3913,In_817,In_823);
nand U3914 (N_3914,In_863,In_270);
nand U3915 (N_3915,In_800,In_118);
nor U3916 (N_3916,In_113,In_881);
and U3917 (N_3917,In_545,In_859);
nand U3918 (N_3918,In_268,In_678);
and U3919 (N_3919,In_953,In_46);
nor U3920 (N_3920,In_68,In_791);
nand U3921 (N_3921,In_364,In_900);
or U3922 (N_3922,In_310,In_336);
nor U3923 (N_3923,In_692,In_697);
nand U3924 (N_3924,In_78,In_878);
and U3925 (N_3925,In_823,In_576);
nor U3926 (N_3926,In_973,In_918);
and U3927 (N_3927,In_768,In_258);
nor U3928 (N_3928,In_228,In_653);
or U3929 (N_3929,In_548,In_216);
nand U3930 (N_3930,In_480,In_974);
or U3931 (N_3931,In_770,In_497);
nor U3932 (N_3932,In_759,In_648);
nor U3933 (N_3933,In_73,In_604);
nand U3934 (N_3934,In_988,In_897);
nand U3935 (N_3935,In_239,In_278);
or U3936 (N_3936,In_532,In_370);
nor U3937 (N_3937,In_79,In_574);
and U3938 (N_3938,In_157,In_818);
and U3939 (N_3939,In_176,In_595);
or U3940 (N_3940,In_46,In_385);
nand U3941 (N_3941,In_449,In_52);
and U3942 (N_3942,In_222,In_617);
nand U3943 (N_3943,In_456,In_629);
and U3944 (N_3944,In_460,In_757);
or U3945 (N_3945,In_187,In_370);
and U3946 (N_3946,In_342,In_610);
nand U3947 (N_3947,In_988,In_474);
nor U3948 (N_3948,In_672,In_486);
or U3949 (N_3949,In_883,In_727);
or U3950 (N_3950,In_645,In_542);
or U3951 (N_3951,In_9,In_219);
nor U3952 (N_3952,In_648,In_93);
or U3953 (N_3953,In_827,In_524);
nor U3954 (N_3954,In_381,In_258);
and U3955 (N_3955,In_762,In_368);
and U3956 (N_3956,In_49,In_326);
nand U3957 (N_3957,In_321,In_168);
nor U3958 (N_3958,In_605,In_838);
nand U3959 (N_3959,In_754,In_904);
or U3960 (N_3960,In_839,In_828);
nand U3961 (N_3961,In_663,In_971);
and U3962 (N_3962,In_863,In_261);
and U3963 (N_3963,In_158,In_891);
nand U3964 (N_3964,In_184,In_359);
nand U3965 (N_3965,In_321,In_798);
nand U3966 (N_3966,In_398,In_346);
and U3967 (N_3967,In_95,In_966);
or U3968 (N_3968,In_633,In_872);
and U3969 (N_3969,In_473,In_169);
or U3970 (N_3970,In_917,In_743);
and U3971 (N_3971,In_348,In_366);
nor U3972 (N_3972,In_793,In_873);
nand U3973 (N_3973,In_832,In_869);
or U3974 (N_3974,In_751,In_236);
nor U3975 (N_3975,In_549,In_440);
nand U3976 (N_3976,In_475,In_601);
nand U3977 (N_3977,In_158,In_682);
or U3978 (N_3978,In_573,In_637);
or U3979 (N_3979,In_80,In_717);
and U3980 (N_3980,In_0,In_553);
or U3981 (N_3981,In_91,In_899);
and U3982 (N_3982,In_687,In_551);
xor U3983 (N_3983,In_386,In_525);
nand U3984 (N_3984,In_319,In_327);
nand U3985 (N_3985,In_664,In_173);
nand U3986 (N_3986,In_931,In_365);
or U3987 (N_3987,In_322,In_707);
or U3988 (N_3988,In_234,In_466);
and U3989 (N_3989,In_220,In_684);
nor U3990 (N_3990,In_244,In_954);
nand U3991 (N_3991,In_627,In_39);
or U3992 (N_3992,In_762,In_219);
or U3993 (N_3993,In_697,In_548);
nand U3994 (N_3994,In_715,In_632);
nand U3995 (N_3995,In_642,In_17);
or U3996 (N_3996,In_734,In_185);
nand U3997 (N_3997,In_533,In_715);
nor U3998 (N_3998,In_865,In_907);
nand U3999 (N_3999,In_195,In_811);
and U4000 (N_4000,In_226,In_755);
nor U4001 (N_4001,In_781,In_6);
or U4002 (N_4002,In_236,In_821);
nor U4003 (N_4003,In_68,In_217);
and U4004 (N_4004,In_622,In_45);
nor U4005 (N_4005,In_745,In_709);
nor U4006 (N_4006,In_262,In_493);
or U4007 (N_4007,In_345,In_635);
or U4008 (N_4008,In_703,In_607);
nand U4009 (N_4009,In_378,In_828);
and U4010 (N_4010,In_310,In_405);
nand U4011 (N_4011,In_476,In_794);
and U4012 (N_4012,In_210,In_254);
nand U4013 (N_4013,In_389,In_899);
and U4014 (N_4014,In_370,In_737);
and U4015 (N_4015,In_949,In_478);
nor U4016 (N_4016,In_167,In_505);
and U4017 (N_4017,In_144,In_49);
nand U4018 (N_4018,In_749,In_713);
nand U4019 (N_4019,In_639,In_529);
nand U4020 (N_4020,In_577,In_587);
nor U4021 (N_4021,In_31,In_3);
and U4022 (N_4022,In_537,In_744);
or U4023 (N_4023,In_692,In_975);
nor U4024 (N_4024,In_839,In_229);
xor U4025 (N_4025,In_477,In_464);
nor U4026 (N_4026,In_272,In_905);
or U4027 (N_4027,In_111,In_107);
nor U4028 (N_4028,In_507,In_733);
nand U4029 (N_4029,In_436,In_780);
or U4030 (N_4030,In_655,In_908);
or U4031 (N_4031,In_672,In_653);
or U4032 (N_4032,In_651,In_986);
or U4033 (N_4033,In_813,In_528);
or U4034 (N_4034,In_263,In_723);
or U4035 (N_4035,In_270,In_624);
and U4036 (N_4036,In_749,In_550);
or U4037 (N_4037,In_670,In_856);
nor U4038 (N_4038,In_11,In_644);
nor U4039 (N_4039,In_519,In_137);
or U4040 (N_4040,In_221,In_663);
nand U4041 (N_4041,In_8,In_457);
and U4042 (N_4042,In_807,In_94);
nand U4043 (N_4043,In_389,In_200);
and U4044 (N_4044,In_294,In_736);
nor U4045 (N_4045,In_411,In_692);
or U4046 (N_4046,In_822,In_511);
and U4047 (N_4047,In_5,In_198);
and U4048 (N_4048,In_398,In_212);
nor U4049 (N_4049,In_326,In_425);
or U4050 (N_4050,In_932,In_475);
nor U4051 (N_4051,In_802,In_462);
nor U4052 (N_4052,In_642,In_109);
nand U4053 (N_4053,In_776,In_664);
nor U4054 (N_4054,In_804,In_477);
or U4055 (N_4055,In_79,In_242);
and U4056 (N_4056,In_131,In_138);
or U4057 (N_4057,In_389,In_6);
nor U4058 (N_4058,In_87,In_646);
or U4059 (N_4059,In_887,In_646);
or U4060 (N_4060,In_33,In_50);
nor U4061 (N_4061,In_803,In_209);
and U4062 (N_4062,In_391,In_497);
or U4063 (N_4063,In_725,In_394);
or U4064 (N_4064,In_277,In_194);
and U4065 (N_4065,In_732,In_674);
nor U4066 (N_4066,In_7,In_977);
nor U4067 (N_4067,In_198,In_56);
and U4068 (N_4068,In_496,In_331);
nand U4069 (N_4069,In_847,In_358);
or U4070 (N_4070,In_559,In_426);
nor U4071 (N_4071,In_743,In_952);
or U4072 (N_4072,In_13,In_753);
nand U4073 (N_4073,In_313,In_656);
and U4074 (N_4074,In_925,In_264);
nand U4075 (N_4075,In_566,In_203);
nor U4076 (N_4076,In_277,In_878);
and U4077 (N_4077,In_26,In_475);
nor U4078 (N_4078,In_708,In_697);
nor U4079 (N_4079,In_748,In_429);
and U4080 (N_4080,In_234,In_802);
nor U4081 (N_4081,In_461,In_234);
or U4082 (N_4082,In_286,In_167);
or U4083 (N_4083,In_444,In_384);
nand U4084 (N_4084,In_981,In_789);
nor U4085 (N_4085,In_513,In_266);
and U4086 (N_4086,In_742,In_506);
nor U4087 (N_4087,In_490,In_516);
nand U4088 (N_4088,In_347,In_828);
and U4089 (N_4089,In_916,In_226);
and U4090 (N_4090,In_638,In_257);
nor U4091 (N_4091,In_278,In_622);
nor U4092 (N_4092,In_557,In_325);
or U4093 (N_4093,In_592,In_818);
nor U4094 (N_4094,In_129,In_893);
nor U4095 (N_4095,In_620,In_363);
nor U4096 (N_4096,In_921,In_62);
xor U4097 (N_4097,In_203,In_337);
nor U4098 (N_4098,In_563,In_31);
nand U4099 (N_4099,In_663,In_779);
and U4100 (N_4100,In_119,In_955);
xor U4101 (N_4101,In_963,In_196);
nor U4102 (N_4102,In_811,In_167);
nand U4103 (N_4103,In_905,In_696);
or U4104 (N_4104,In_161,In_543);
or U4105 (N_4105,In_939,In_559);
and U4106 (N_4106,In_157,In_819);
nor U4107 (N_4107,In_810,In_125);
nand U4108 (N_4108,In_544,In_963);
nor U4109 (N_4109,In_888,In_53);
nand U4110 (N_4110,In_756,In_189);
nand U4111 (N_4111,In_370,In_770);
nor U4112 (N_4112,In_611,In_142);
or U4113 (N_4113,In_336,In_703);
nor U4114 (N_4114,In_308,In_963);
and U4115 (N_4115,In_844,In_660);
nor U4116 (N_4116,In_275,In_668);
and U4117 (N_4117,In_962,In_484);
nor U4118 (N_4118,In_12,In_487);
or U4119 (N_4119,In_41,In_872);
or U4120 (N_4120,In_627,In_527);
nor U4121 (N_4121,In_108,In_982);
nand U4122 (N_4122,In_931,In_874);
xor U4123 (N_4123,In_810,In_590);
and U4124 (N_4124,In_348,In_245);
or U4125 (N_4125,In_922,In_950);
nor U4126 (N_4126,In_123,In_551);
or U4127 (N_4127,In_137,In_112);
and U4128 (N_4128,In_864,In_237);
and U4129 (N_4129,In_499,In_985);
and U4130 (N_4130,In_756,In_145);
and U4131 (N_4131,In_942,In_103);
nand U4132 (N_4132,In_285,In_476);
nor U4133 (N_4133,In_340,In_560);
nor U4134 (N_4134,In_243,In_297);
nor U4135 (N_4135,In_851,In_514);
nor U4136 (N_4136,In_460,In_74);
nand U4137 (N_4137,In_349,In_771);
and U4138 (N_4138,In_65,In_607);
and U4139 (N_4139,In_947,In_2);
or U4140 (N_4140,In_401,In_465);
xor U4141 (N_4141,In_421,In_495);
nor U4142 (N_4142,In_356,In_822);
nor U4143 (N_4143,In_896,In_66);
nand U4144 (N_4144,In_837,In_658);
nor U4145 (N_4145,In_192,In_246);
nor U4146 (N_4146,In_162,In_830);
nor U4147 (N_4147,In_845,In_126);
nor U4148 (N_4148,In_792,In_381);
or U4149 (N_4149,In_931,In_465);
and U4150 (N_4150,In_811,In_3);
and U4151 (N_4151,In_562,In_260);
or U4152 (N_4152,In_698,In_295);
nor U4153 (N_4153,In_381,In_793);
and U4154 (N_4154,In_173,In_906);
and U4155 (N_4155,In_347,In_856);
and U4156 (N_4156,In_243,In_14);
nand U4157 (N_4157,In_836,In_434);
nand U4158 (N_4158,In_818,In_86);
or U4159 (N_4159,In_973,In_997);
and U4160 (N_4160,In_599,In_400);
nor U4161 (N_4161,In_860,In_835);
or U4162 (N_4162,In_117,In_158);
xor U4163 (N_4163,In_499,In_23);
xor U4164 (N_4164,In_200,In_272);
or U4165 (N_4165,In_28,In_18);
and U4166 (N_4166,In_896,In_366);
nor U4167 (N_4167,In_76,In_391);
nor U4168 (N_4168,In_650,In_386);
nor U4169 (N_4169,In_52,In_472);
nor U4170 (N_4170,In_329,In_785);
nor U4171 (N_4171,In_394,In_407);
nor U4172 (N_4172,In_500,In_621);
or U4173 (N_4173,In_108,In_939);
and U4174 (N_4174,In_97,In_484);
and U4175 (N_4175,In_28,In_363);
nand U4176 (N_4176,In_925,In_707);
nand U4177 (N_4177,In_498,In_325);
nor U4178 (N_4178,In_104,In_720);
nor U4179 (N_4179,In_458,In_246);
or U4180 (N_4180,In_833,In_720);
and U4181 (N_4181,In_704,In_909);
or U4182 (N_4182,In_178,In_97);
and U4183 (N_4183,In_265,In_95);
nor U4184 (N_4184,In_12,In_536);
nor U4185 (N_4185,In_848,In_482);
nor U4186 (N_4186,In_86,In_731);
nand U4187 (N_4187,In_293,In_485);
nor U4188 (N_4188,In_92,In_925);
nor U4189 (N_4189,In_590,In_856);
or U4190 (N_4190,In_691,In_841);
nor U4191 (N_4191,In_239,In_578);
or U4192 (N_4192,In_895,In_454);
or U4193 (N_4193,In_561,In_438);
or U4194 (N_4194,In_715,In_921);
nor U4195 (N_4195,In_912,In_945);
nand U4196 (N_4196,In_953,In_480);
nor U4197 (N_4197,In_584,In_990);
or U4198 (N_4198,In_391,In_338);
nor U4199 (N_4199,In_21,In_580);
nor U4200 (N_4200,In_17,In_974);
nor U4201 (N_4201,In_958,In_401);
nor U4202 (N_4202,In_632,In_507);
nand U4203 (N_4203,In_37,In_516);
nand U4204 (N_4204,In_186,In_556);
nand U4205 (N_4205,In_860,In_726);
and U4206 (N_4206,In_191,In_274);
and U4207 (N_4207,In_127,In_13);
nor U4208 (N_4208,In_616,In_420);
nor U4209 (N_4209,In_794,In_557);
nand U4210 (N_4210,In_434,In_576);
and U4211 (N_4211,In_730,In_488);
and U4212 (N_4212,In_787,In_326);
nand U4213 (N_4213,In_552,In_33);
nor U4214 (N_4214,In_506,In_635);
nand U4215 (N_4215,In_436,In_520);
or U4216 (N_4216,In_192,In_857);
nand U4217 (N_4217,In_305,In_340);
nand U4218 (N_4218,In_832,In_339);
or U4219 (N_4219,In_779,In_889);
nand U4220 (N_4220,In_119,In_936);
nand U4221 (N_4221,In_218,In_993);
and U4222 (N_4222,In_521,In_554);
nor U4223 (N_4223,In_666,In_712);
nand U4224 (N_4224,In_610,In_13);
nand U4225 (N_4225,In_958,In_851);
nand U4226 (N_4226,In_324,In_618);
nor U4227 (N_4227,In_242,In_483);
nand U4228 (N_4228,In_794,In_484);
nor U4229 (N_4229,In_528,In_603);
nor U4230 (N_4230,In_244,In_262);
nand U4231 (N_4231,In_998,In_660);
nand U4232 (N_4232,In_117,In_667);
nor U4233 (N_4233,In_711,In_785);
nand U4234 (N_4234,In_53,In_868);
and U4235 (N_4235,In_317,In_811);
nor U4236 (N_4236,In_957,In_305);
nor U4237 (N_4237,In_447,In_809);
and U4238 (N_4238,In_746,In_218);
nor U4239 (N_4239,In_447,In_248);
or U4240 (N_4240,In_814,In_259);
and U4241 (N_4241,In_739,In_609);
or U4242 (N_4242,In_985,In_295);
or U4243 (N_4243,In_230,In_200);
nor U4244 (N_4244,In_837,In_741);
nand U4245 (N_4245,In_26,In_869);
and U4246 (N_4246,In_274,In_880);
or U4247 (N_4247,In_850,In_822);
nand U4248 (N_4248,In_785,In_561);
nor U4249 (N_4249,In_336,In_419);
or U4250 (N_4250,In_486,In_247);
and U4251 (N_4251,In_808,In_920);
and U4252 (N_4252,In_745,In_177);
nor U4253 (N_4253,In_225,In_377);
nor U4254 (N_4254,In_223,In_565);
nor U4255 (N_4255,In_629,In_773);
or U4256 (N_4256,In_876,In_420);
nor U4257 (N_4257,In_642,In_132);
or U4258 (N_4258,In_315,In_569);
and U4259 (N_4259,In_396,In_162);
or U4260 (N_4260,In_171,In_539);
nor U4261 (N_4261,In_372,In_464);
and U4262 (N_4262,In_578,In_725);
nor U4263 (N_4263,In_203,In_154);
nor U4264 (N_4264,In_968,In_685);
or U4265 (N_4265,In_17,In_24);
or U4266 (N_4266,In_547,In_701);
nor U4267 (N_4267,In_67,In_9);
nor U4268 (N_4268,In_108,In_959);
or U4269 (N_4269,In_932,In_468);
nand U4270 (N_4270,In_194,In_760);
nor U4271 (N_4271,In_635,In_347);
nand U4272 (N_4272,In_749,In_322);
and U4273 (N_4273,In_651,In_171);
and U4274 (N_4274,In_737,In_257);
nand U4275 (N_4275,In_994,In_693);
nor U4276 (N_4276,In_992,In_167);
nand U4277 (N_4277,In_670,In_56);
and U4278 (N_4278,In_904,In_87);
nor U4279 (N_4279,In_397,In_339);
or U4280 (N_4280,In_56,In_819);
nor U4281 (N_4281,In_96,In_751);
nand U4282 (N_4282,In_108,In_272);
nor U4283 (N_4283,In_629,In_467);
nand U4284 (N_4284,In_175,In_352);
and U4285 (N_4285,In_134,In_160);
and U4286 (N_4286,In_259,In_144);
nor U4287 (N_4287,In_702,In_415);
or U4288 (N_4288,In_364,In_308);
and U4289 (N_4289,In_989,In_302);
and U4290 (N_4290,In_854,In_272);
nor U4291 (N_4291,In_507,In_645);
and U4292 (N_4292,In_986,In_199);
or U4293 (N_4293,In_932,In_128);
and U4294 (N_4294,In_275,In_396);
and U4295 (N_4295,In_148,In_537);
nor U4296 (N_4296,In_339,In_75);
or U4297 (N_4297,In_634,In_158);
nor U4298 (N_4298,In_571,In_305);
and U4299 (N_4299,In_332,In_551);
or U4300 (N_4300,In_876,In_569);
or U4301 (N_4301,In_306,In_793);
nand U4302 (N_4302,In_533,In_678);
or U4303 (N_4303,In_827,In_7);
and U4304 (N_4304,In_505,In_701);
nand U4305 (N_4305,In_511,In_878);
nor U4306 (N_4306,In_18,In_876);
or U4307 (N_4307,In_67,In_811);
or U4308 (N_4308,In_861,In_460);
nor U4309 (N_4309,In_75,In_264);
nor U4310 (N_4310,In_595,In_559);
nand U4311 (N_4311,In_756,In_245);
nor U4312 (N_4312,In_825,In_170);
nand U4313 (N_4313,In_706,In_101);
or U4314 (N_4314,In_113,In_661);
nand U4315 (N_4315,In_913,In_287);
and U4316 (N_4316,In_63,In_425);
and U4317 (N_4317,In_892,In_905);
and U4318 (N_4318,In_205,In_708);
nand U4319 (N_4319,In_63,In_833);
nor U4320 (N_4320,In_93,In_833);
nand U4321 (N_4321,In_629,In_18);
and U4322 (N_4322,In_449,In_193);
nand U4323 (N_4323,In_49,In_354);
and U4324 (N_4324,In_143,In_98);
and U4325 (N_4325,In_199,In_387);
nand U4326 (N_4326,In_942,In_845);
or U4327 (N_4327,In_861,In_507);
nor U4328 (N_4328,In_478,In_378);
nand U4329 (N_4329,In_281,In_85);
and U4330 (N_4330,In_929,In_98);
or U4331 (N_4331,In_740,In_867);
nand U4332 (N_4332,In_147,In_203);
and U4333 (N_4333,In_934,In_25);
nand U4334 (N_4334,In_625,In_171);
or U4335 (N_4335,In_5,In_693);
and U4336 (N_4336,In_602,In_513);
xor U4337 (N_4337,In_355,In_637);
and U4338 (N_4338,In_307,In_286);
nor U4339 (N_4339,In_175,In_207);
and U4340 (N_4340,In_708,In_196);
and U4341 (N_4341,In_150,In_213);
nor U4342 (N_4342,In_789,In_142);
and U4343 (N_4343,In_9,In_359);
or U4344 (N_4344,In_782,In_557);
nor U4345 (N_4345,In_469,In_656);
or U4346 (N_4346,In_106,In_853);
nand U4347 (N_4347,In_126,In_478);
or U4348 (N_4348,In_832,In_949);
and U4349 (N_4349,In_482,In_996);
nand U4350 (N_4350,In_958,In_68);
nand U4351 (N_4351,In_622,In_967);
nor U4352 (N_4352,In_468,In_68);
or U4353 (N_4353,In_332,In_871);
or U4354 (N_4354,In_359,In_601);
nor U4355 (N_4355,In_111,In_164);
and U4356 (N_4356,In_901,In_44);
or U4357 (N_4357,In_632,In_912);
and U4358 (N_4358,In_414,In_878);
and U4359 (N_4359,In_737,In_200);
and U4360 (N_4360,In_665,In_549);
nand U4361 (N_4361,In_996,In_865);
or U4362 (N_4362,In_941,In_534);
nand U4363 (N_4363,In_831,In_297);
nand U4364 (N_4364,In_123,In_636);
nor U4365 (N_4365,In_497,In_805);
and U4366 (N_4366,In_724,In_21);
nor U4367 (N_4367,In_83,In_230);
and U4368 (N_4368,In_639,In_514);
and U4369 (N_4369,In_859,In_667);
and U4370 (N_4370,In_38,In_203);
nand U4371 (N_4371,In_810,In_897);
and U4372 (N_4372,In_859,In_669);
nor U4373 (N_4373,In_512,In_366);
nand U4374 (N_4374,In_999,In_883);
nand U4375 (N_4375,In_606,In_425);
nor U4376 (N_4376,In_726,In_456);
and U4377 (N_4377,In_227,In_533);
nor U4378 (N_4378,In_20,In_703);
or U4379 (N_4379,In_884,In_911);
and U4380 (N_4380,In_465,In_598);
or U4381 (N_4381,In_951,In_872);
and U4382 (N_4382,In_249,In_977);
or U4383 (N_4383,In_37,In_433);
nor U4384 (N_4384,In_325,In_427);
or U4385 (N_4385,In_776,In_253);
nand U4386 (N_4386,In_71,In_678);
nor U4387 (N_4387,In_965,In_384);
or U4388 (N_4388,In_772,In_373);
or U4389 (N_4389,In_266,In_208);
and U4390 (N_4390,In_487,In_377);
nor U4391 (N_4391,In_741,In_688);
nand U4392 (N_4392,In_64,In_539);
and U4393 (N_4393,In_570,In_258);
or U4394 (N_4394,In_873,In_285);
nor U4395 (N_4395,In_184,In_489);
nor U4396 (N_4396,In_447,In_239);
nor U4397 (N_4397,In_37,In_803);
nand U4398 (N_4398,In_21,In_375);
nand U4399 (N_4399,In_491,In_56);
nand U4400 (N_4400,In_699,In_890);
nand U4401 (N_4401,In_118,In_535);
or U4402 (N_4402,In_216,In_490);
nand U4403 (N_4403,In_125,In_212);
nand U4404 (N_4404,In_862,In_388);
or U4405 (N_4405,In_138,In_265);
or U4406 (N_4406,In_480,In_321);
and U4407 (N_4407,In_324,In_436);
nor U4408 (N_4408,In_535,In_333);
nand U4409 (N_4409,In_782,In_672);
nor U4410 (N_4410,In_166,In_776);
nand U4411 (N_4411,In_600,In_152);
nor U4412 (N_4412,In_379,In_890);
and U4413 (N_4413,In_396,In_442);
or U4414 (N_4414,In_142,In_712);
nor U4415 (N_4415,In_960,In_902);
nor U4416 (N_4416,In_637,In_461);
nand U4417 (N_4417,In_13,In_757);
and U4418 (N_4418,In_261,In_423);
and U4419 (N_4419,In_402,In_741);
or U4420 (N_4420,In_212,In_266);
or U4421 (N_4421,In_642,In_977);
or U4422 (N_4422,In_944,In_507);
nor U4423 (N_4423,In_843,In_983);
and U4424 (N_4424,In_98,In_737);
nand U4425 (N_4425,In_76,In_928);
and U4426 (N_4426,In_73,In_48);
and U4427 (N_4427,In_744,In_379);
and U4428 (N_4428,In_61,In_817);
and U4429 (N_4429,In_104,In_504);
nand U4430 (N_4430,In_297,In_463);
or U4431 (N_4431,In_591,In_435);
and U4432 (N_4432,In_301,In_611);
or U4433 (N_4433,In_20,In_104);
and U4434 (N_4434,In_131,In_51);
nand U4435 (N_4435,In_169,In_232);
and U4436 (N_4436,In_970,In_834);
nor U4437 (N_4437,In_512,In_753);
nand U4438 (N_4438,In_815,In_26);
or U4439 (N_4439,In_329,In_479);
nand U4440 (N_4440,In_2,In_415);
and U4441 (N_4441,In_955,In_741);
and U4442 (N_4442,In_506,In_636);
or U4443 (N_4443,In_231,In_392);
and U4444 (N_4444,In_176,In_239);
or U4445 (N_4445,In_95,In_136);
or U4446 (N_4446,In_502,In_671);
or U4447 (N_4447,In_544,In_467);
nor U4448 (N_4448,In_131,In_67);
nand U4449 (N_4449,In_995,In_180);
nand U4450 (N_4450,In_402,In_452);
and U4451 (N_4451,In_513,In_459);
nor U4452 (N_4452,In_890,In_503);
nand U4453 (N_4453,In_75,In_336);
nor U4454 (N_4454,In_145,In_773);
nand U4455 (N_4455,In_68,In_892);
nor U4456 (N_4456,In_558,In_337);
nand U4457 (N_4457,In_563,In_320);
nand U4458 (N_4458,In_366,In_995);
nor U4459 (N_4459,In_326,In_848);
nand U4460 (N_4460,In_101,In_406);
and U4461 (N_4461,In_475,In_667);
nand U4462 (N_4462,In_622,In_556);
nor U4463 (N_4463,In_116,In_103);
and U4464 (N_4464,In_845,In_112);
and U4465 (N_4465,In_805,In_446);
or U4466 (N_4466,In_223,In_19);
and U4467 (N_4467,In_625,In_950);
nor U4468 (N_4468,In_954,In_592);
nor U4469 (N_4469,In_269,In_521);
nand U4470 (N_4470,In_273,In_413);
and U4471 (N_4471,In_957,In_253);
and U4472 (N_4472,In_805,In_137);
or U4473 (N_4473,In_182,In_965);
or U4474 (N_4474,In_863,In_459);
nor U4475 (N_4475,In_224,In_226);
and U4476 (N_4476,In_201,In_392);
and U4477 (N_4477,In_260,In_9);
nand U4478 (N_4478,In_277,In_547);
and U4479 (N_4479,In_882,In_405);
nand U4480 (N_4480,In_376,In_213);
or U4481 (N_4481,In_689,In_286);
or U4482 (N_4482,In_139,In_203);
nand U4483 (N_4483,In_26,In_747);
nand U4484 (N_4484,In_886,In_210);
xnor U4485 (N_4485,In_854,In_85);
nor U4486 (N_4486,In_847,In_785);
and U4487 (N_4487,In_698,In_749);
and U4488 (N_4488,In_50,In_178);
or U4489 (N_4489,In_545,In_669);
nand U4490 (N_4490,In_860,In_971);
or U4491 (N_4491,In_234,In_985);
nand U4492 (N_4492,In_49,In_912);
nand U4493 (N_4493,In_176,In_774);
or U4494 (N_4494,In_933,In_811);
and U4495 (N_4495,In_637,In_143);
nand U4496 (N_4496,In_471,In_584);
and U4497 (N_4497,In_19,In_249);
or U4498 (N_4498,In_774,In_321);
and U4499 (N_4499,In_686,In_163);
nand U4500 (N_4500,In_824,In_147);
or U4501 (N_4501,In_679,In_636);
nor U4502 (N_4502,In_107,In_331);
and U4503 (N_4503,In_792,In_452);
nand U4504 (N_4504,In_942,In_449);
nor U4505 (N_4505,In_659,In_295);
nand U4506 (N_4506,In_331,In_400);
or U4507 (N_4507,In_827,In_228);
nor U4508 (N_4508,In_450,In_716);
nor U4509 (N_4509,In_68,In_113);
or U4510 (N_4510,In_992,In_367);
nand U4511 (N_4511,In_80,In_581);
or U4512 (N_4512,In_127,In_757);
and U4513 (N_4513,In_806,In_721);
nor U4514 (N_4514,In_729,In_34);
or U4515 (N_4515,In_873,In_922);
or U4516 (N_4516,In_344,In_912);
nor U4517 (N_4517,In_891,In_829);
or U4518 (N_4518,In_688,In_180);
nor U4519 (N_4519,In_945,In_49);
nand U4520 (N_4520,In_967,In_451);
and U4521 (N_4521,In_452,In_809);
nand U4522 (N_4522,In_658,In_76);
and U4523 (N_4523,In_683,In_413);
nand U4524 (N_4524,In_430,In_95);
and U4525 (N_4525,In_850,In_786);
and U4526 (N_4526,In_845,In_60);
and U4527 (N_4527,In_977,In_25);
or U4528 (N_4528,In_195,In_763);
nor U4529 (N_4529,In_301,In_742);
or U4530 (N_4530,In_757,In_412);
nor U4531 (N_4531,In_310,In_214);
nor U4532 (N_4532,In_467,In_145);
nand U4533 (N_4533,In_306,In_303);
or U4534 (N_4534,In_170,In_800);
nand U4535 (N_4535,In_307,In_136);
and U4536 (N_4536,In_630,In_158);
or U4537 (N_4537,In_667,In_964);
and U4538 (N_4538,In_887,In_51);
nand U4539 (N_4539,In_606,In_186);
and U4540 (N_4540,In_571,In_328);
or U4541 (N_4541,In_723,In_612);
and U4542 (N_4542,In_106,In_177);
nor U4543 (N_4543,In_948,In_828);
nand U4544 (N_4544,In_406,In_843);
or U4545 (N_4545,In_797,In_791);
and U4546 (N_4546,In_865,In_436);
nand U4547 (N_4547,In_793,In_543);
and U4548 (N_4548,In_735,In_168);
and U4549 (N_4549,In_428,In_88);
and U4550 (N_4550,In_607,In_258);
and U4551 (N_4551,In_794,In_120);
and U4552 (N_4552,In_782,In_661);
nor U4553 (N_4553,In_779,In_44);
nand U4554 (N_4554,In_877,In_309);
nand U4555 (N_4555,In_289,In_556);
and U4556 (N_4556,In_96,In_767);
and U4557 (N_4557,In_480,In_47);
nand U4558 (N_4558,In_285,In_62);
nor U4559 (N_4559,In_68,In_836);
or U4560 (N_4560,In_284,In_929);
or U4561 (N_4561,In_185,In_662);
nand U4562 (N_4562,In_363,In_785);
nor U4563 (N_4563,In_728,In_579);
and U4564 (N_4564,In_490,In_252);
or U4565 (N_4565,In_666,In_470);
nor U4566 (N_4566,In_856,In_686);
nand U4567 (N_4567,In_816,In_718);
and U4568 (N_4568,In_440,In_825);
nand U4569 (N_4569,In_105,In_772);
or U4570 (N_4570,In_625,In_339);
and U4571 (N_4571,In_679,In_470);
and U4572 (N_4572,In_824,In_930);
and U4573 (N_4573,In_278,In_289);
nor U4574 (N_4574,In_886,In_700);
or U4575 (N_4575,In_213,In_792);
nor U4576 (N_4576,In_544,In_392);
nand U4577 (N_4577,In_151,In_403);
or U4578 (N_4578,In_141,In_192);
or U4579 (N_4579,In_172,In_961);
nor U4580 (N_4580,In_844,In_584);
and U4581 (N_4581,In_352,In_553);
nand U4582 (N_4582,In_699,In_124);
nand U4583 (N_4583,In_216,In_199);
nor U4584 (N_4584,In_762,In_464);
and U4585 (N_4585,In_456,In_44);
or U4586 (N_4586,In_460,In_328);
nor U4587 (N_4587,In_273,In_89);
and U4588 (N_4588,In_925,In_173);
and U4589 (N_4589,In_365,In_463);
nand U4590 (N_4590,In_415,In_43);
or U4591 (N_4591,In_622,In_97);
and U4592 (N_4592,In_490,In_343);
or U4593 (N_4593,In_656,In_763);
nand U4594 (N_4594,In_655,In_68);
and U4595 (N_4595,In_333,In_47);
or U4596 (N_4596,In_308,In_903);
or U4597 (N_4597,In_850,In_892);
nor U4598 (N_4598,In_911,In_589);
nand U4599 (N_4599,In_329,In_344);
nor U4600 (N_4600,In_437,In_654);
nor U4601 (N_4601,In_778,In_26);
nor U4602 (N_4602,In_939,In_438);
nor U4603 (N_4603,In_467,In_714);
and U4604 (N_4604,In_620,In_257);
nor U4605 (N_4605,In_982,In_44);
or U4606 (N_4606,In_611,In_915);
nand U4607 (N_4607,In_533,In_114);
nand U4608 (N_4608,In_355,In_361);
nand U4609 (N_4609,In_849,In_851);
nand U4610 (N_4610,In_484,In_270);
and U4611 (N_4611,In_835,In_19);
nand U4612 (N_4612,In_948,In_43);
nor U4613 (N_4613,In_407,In_282);
nor U4614 (N_4614,In_73,In_769);
or U4615 (N_4615,In_899,In_224);
nand U4616 (N_4616,In_277,In_577);
nor U4617 (N_4617,In_652,In_809);
nand U4618 (N_4618,In_407,In_839);
or U4619 (N_4619,In_512,In_802);
and U4620 (N_4620,In_110,In_999);
and U4621 (N_4621,In_379,In_221);
nor U4622 (N_4622,In_686,In_376);
nand U4623 (N_4623,In_247,In_62);
nor U4624 (N_4624,In_801,In_923);
nand U4625 (N_4625,In_338,In_23);
or U4626 (N_4626,In_886,In_593);
nand U4627 (N_4627,In_37,In_188);
and U4628 (N_4628,In_711,In_729);
and U4629 (N_4629,In_221,In_977);
and U4630 (N_4630,In_330,In_702);
nand U4631 (N_4631,In_956,In_216);
nor U4632 (N_4632,In_361,In_998);
and U4633 (N_4633,In_18,In_339);
and U4634 (N_4634,In_477,In_710);
or U4635 (N_4635,In_870,In_431);
or U4636 (N_4636,In_964,In_176);
nand U4637 (N_4637,In_691,In_978);
or U4638 (N_4638,In_808,In_601);
and U4639 (N_4639,In_0,In_996);
nand U4640 (N_4640,In_465,In_660);
nor U4641 (N_4641,In_620,In_781);
or U4642 (N_4642,In_621,In_898);
nand U4643 (N_4643,In_624,In_129);
or U4644 (N_4644,In_699,In_107);
and U4645 (N_4645,In_543,In_673);
nor U4646 (N_4646,In_724,In_463);
or U4647 (N_4647,In_789,In_603);
and U4648 (N_4648,In_177,In_109);
and U4649 (N_4649,In_255,In_721);
or U4650 (N_4650,In_599,In_637);
nand U4651 (N_4651,In_610,In_879);
and U4652 (N_4652,In_955,In_173);
nor U4653 (N_4653,In_443,In_875);
nand U4654 (N_4654,In_380,In_976);
and U4655 (N_4655,In_674,In_255);
or U4656 (N_4656,In_767,In_835);
nor U4657 (N_4657,In_312,In_248);
nand U4658 (N_4658,In_39,In_917);
and U4659 (N_4659,In_36,In_127);
nor U4660 (N_4660,In_37,In_814);
nor U4661 (N_4661,In_927,In_700);
nor U4662 (N_4662,In_681,In_254);
nand U4663 (N_4663,In_304,In_683);
nand U4664 (N_4664,In_413,In_220);
or U4665 (N_4665,In_948,In_241);
and U4666 (N_4666,In_482,In_196);
and U4667 (N_4667,In_709,In_900);
or U4668 (N_4668,In_51,In_879);
nor U4669 (N_4669,In_799,In_551);
and U4670 (N_4670,In_744,In_806);
nand U4671 (N_4671,In_41,In_193);
nand U4672 (N_4672,In_191,In_829);
or U4673 (N_4673,In_389,In_50);
and U4674 (N_4674,In_146,In_255);
nor U4675 (N_4675,In_785,In_513);
nor U4676 (N_4676,In_696,In_283);
or U4677 (N_4677,In_648,In_950);
nor U4678 (N_4678,In_995,In_843);
and U4679 (N_4679,In_733,In_114);
and U4680 (N_4680,In_159,In_857);
nand U4681 (N_4681,In_81,In_125);
or U4682 (N_4682,In_586,In_306);
and U4683 (N_4683,In_564,In_645);
nand U4684 (N_4684,In_698,In_693);
or U4685 (N_4685,In_363,In_125);
and U4686 (N_4686,In_633,In_540);
or U4687 (N_4687,In_71,In_55);
nand U4688 (N_4688,In_390,In_550);
nand U4689 (N_4689,In_219,In_946);
nand U4690 (N_4690,In_879,In_344);
nor U4691 (N_4691,In_994,In_829);
xnor U4692 (N_4692,In_695,In_353);
nor U4693 (N_4693,In_918,In_991);
nor U4694 (N_4694,In_367,In_577);
nor U4695 (N_4695,In_481,In_205);
nor U4696 (N_4696,In_330,In_523);
nand U4697 (N_4697,In_763,In_316);
and U4698 (N_4698,In_437,In_127);
or U4699 (N_4699,In_503,In_280);
or U4700 (N_4700,In_503,In_882);
and U4701 (N_4701,In_798,In_853);
nor U4702 (N_4702,In_55,In_512);
and U4703 (N_4703,In_212,In_160);
nand U4704 (N_4704,In_702,In_783);
or U4705 (N_4705,In_910,In_816);
and U4706 (N_4706,In_675,In_207);
nand U4707 (N_4707,In_234,In_724);
nor U4708 (N_4708,In_393,In_804);
nand U4709 (N_4709,In_853,In_552);
and U4710 (N_4710,In_742,In_329);
or U4711 (N_4711,In_826,In_190);
nand U4712 (N_4712,In_77,In_479);
or U4713 (N_4713,In_712,In_665);
and U4714 (N_4714,In_506,In_869);
or U4715 (N_4715,In_705,In_776);
nand U4716 (N_4716,In_818,In_495);
and U4717 (N_4717,In_630,In_654);
or U4718 (N_4718,In_182,In_220);
nor U4719 (N_4719,In_379,In_430);
or U4720 (N_4720,In_609,In_530);
nor U4721 (N_4721,In_381,In_263);
nand U4722 (N_4722,In_524,In_632);
and U4723 (N_4723,In_833,In_64);
nor U4724 (N_4724,In_401,In_839);
nand U4725 (N_4725,In_452,In_11);
and U4726 (N_4726,In_98,In_529);
nor U4727 (N_4727,In_553,In_370);
nand U4728 (N_4728,In_815,In_995);
or U4729 (N_4729,In_818,In_488);
or U4730 (N_4730,In_886,In_357);
nor U4731 (N_4731,In_756,In_700);
and U4732 (N_4732,In_446,In_280);
or U4733 (N_4733,In_693,In_310);
nand U4734 (N_4734,In_855,In_399);
and U4735 (N_4735,In_877,In_935);
nor U4736 (N_4736,In_703,In_402);
and U4737 (N_4737,In_768,In_457);
or U4738 (N_4738,In_54,In_100);
nand U4739 (N_4739,In_624,In_164);
nand U4740 (N_4740,In_864,In_207);
and U4741 (N_4741,In_725,In_52);
nor U4742 (N_4742,In_143,In_891);
and U4743 (N_4743,In_377,In_457);
nor U4744 (N_4744,In_497,In_475);
nor U4745 (N_4745,In_552,In_753);
nor U4746 (N_4746,In_46,In_769);
nand U4747 (N_4747,In_225,In_606);
and U4748 (N_4748,In_770,In_933);
or U4749 (N_4749,In_695,In_241);
nand U4750 (N_4750,In_879,In_602);
nor U4751 (N_4751,In_639,In_813);
or U4752 (N_4752,In_303,In_627);
nor U4753 (N_4753,In_140,In_651);
nand U4754 (N_4754,In_905,In_76);
or U4755 (N_4755,In_980,In_25);
nor U4756 (N_4756,In_79,In_183);
and U4757 (N_4757,In_924,In_791);
and U4758 (N_4758,In_319,In_622);
or U4759 (N_4759,In_535,In_288);
xnor U4760 (N_4760,In_776,In_126);
and U4761 (N_4761,In_914,In_802);
or U4762 (N_4762,In_308,In_738);
nand U4763 (N_4763,In_354,In_68);
or U4764 (N_4764,In_943,In_772);
nor U4765 (N_4765,In_934,In_776);
or U4766 (N_4766,In_630,In_378);
or U4767 (N_4767,In_428,In_836);
or U4768 (N_4768,In_995,In_984);
nand U4769 (N_4769,In_397,In_720);
and U4770 (N_4770,In_197,In_822);
nand U4771 (N_4771,In_721,In_58);
and U4772 (N_4772,In_924,In_98);
nor U4773 (N_4773,In_28,In_597);
or U4774 (N_4774,In_549,In_733);
nand U4775 (N_4775,In_465,In_442);
nand U4776 (N_4776,In_273,In_546);
nor U4777 (N_4777,In_493,In_893);
nand U4778 (N_4778,In_112,In_583);
and U4779 (N_4779,In_490,In_107);
nand U4780 (N_4780,In_464,In_284);
nor U4781 (N_4781,In_716,In_444);
or U4782 (N_4782,In_238,In_686);
and U4783 (N_4783,In_560,In_884);
or U4784 (N_4784,In_391,In_275);
nor U4785 (N_4785,In_318,In_700);
nand U4786 (N_4786,In_173,In_467);
nor U4787 (N_4787,In_75,In_581);
nand U4788 (N_4788,In_393,In_870);
and U4789 (N_4789,In_207,In_817);
and U4790 (N_4790,In_467,In_791);
nor U4791 (N_4791,In_198,In_478);
or U4792 (N_4792,In_484,In_365);
nand U4793 (N_4793,In_283,In_666);
nand U4794 (N_4794,In_495,In_123);
or U4795 (N_4795,In_486,In_470);
and U4796 (N_4796,In_93,In_748);
and U4797 (N_4797,In_695,In_166);
nor U4798 (N_4798,In_571,In_186);
nand U4799 (N_4799,In_419,In_661);
or U4800 (N_4800,In_999,In_962);
nand U4801 (N_4801,In_497,In_459);
and U4802 (N_4802,In_978,In_635);
and U4803 (N_4803,In_515,In_374);
or U4804 (N_4804,In_484,In_747);
nand U4805 (N_4805,In_791,In_563);
nand U4806 (N_4806,In_780,In_805);
and U4807 (N_4807,In_23,In_335);
and U4808 (N_4808,In_634,In_476);
and U4809 (N_4809,In_623,In_532);
and U4810 (N_4810,In_589,In_674);
or U4811 (N_4811,In_64,In_465);
nand U4812 (N_4812,In_749,In_605);
nor U4813 (N_4813,In_205,In_276);
nand U4814 (N_4814,In_171,In_611);
nand U4815 (N_4815,In_82,In_968);
nor U4816 (N_4816,In_279,In_680);
nor U4817 (N_4817,In_519,In_299);
or U4818 (N_4818,In_951,In_693);
nor U4819 (N_4819,In_798,In_956);
or U4820 (N_4820,In_285,In_355);
and U4821 (N_4821,In_744,In_958);
or U4822 (N_4822,In_814,In_53);
nand U4823 (N_4823,In_554,In_247);
or U4824 (N_4824,In_977,In_213);
nor U4825 (N_4825,In_415,In_283);
and U4826 (N_4826,In_311,In_230);
nand U4827 (N_4827,In_27,In_51);
and U4828 (N_4828,In_297,In_354);
and U4829 (N_4829,In_951,In_599);
nor U4830 (N_4830,In_655,In_459);
or U4831 (N_4831,In_788,In_973);
nor U4832 (N_4832,In_724,In_835);
or U4833 (N_4833,In_553,In_998);
nand U4834 (N_4834,In_920,In_356);
nand U4835 (N_4835,In_299,In_101);
and U4836 (N_4836,In_371,In_674);
nand U4837 (N_4837,In_748,In_227);
or U4838 (N_4838,In_427,In_307);
nand U4839 (N_4839,In_215,In_663);
nor U4840 (N_4840,In_466,In_524);
nand U4841 (N_4841,In_282,In_245);
and U4842 (N_4842,In_303,In_384);
and U4843 (N_4843,In_688,In_885);
and U4844 (N_4844,In_79,In_193);
xor U4845 (N_4845,In_475,In_34);
nand U4846 (N_4846,In_781,In_287);
nand U4847 (N_4847,In_475,In_690);
and U4848 (N_4848,In_475,In_371);
nor U4849 (N_4849,In_197,In_130);
or U4850 (N_4850,In_708,In_487);
or U4851 (N_4851,In_555,In_41);
nor U4852 (N_4852,In_19,In_45);
nor U4853 (N_4853,In_813,In_46);
nor U4854 (N_4854,In_677,In_751);
and U4855 (N_4855,In_314,In_249);
nor U4856 (N_4856,In_487,In_535);
nor U4857 (N_4857,In_521,In_612);
and U4858 (N_4858,In_138,In_832);
or U4859 (N_4859,In_820,In_393);
nor U4860 (N_4860,In_277,In_161);
nor U4861 (N_4861,In_304,In_620);
and U4862 (N_4862,In_408,In_183);
nor U4863 (N_4863,In_88,In_669);
or U4864 (N_4864,In_309,In_2);
and U4865 (N_4865,In_643,In_114);
and U4866 (N_4866,In_512,In_107);
and U4867 (N_4867,In_834,In_57);
and U4868 (N_4868,In_33,In_23);
or U4869 (N_4869,In_771,In_447);
and U4870 (N_4870,In_35,In_225);
nor U4871 (N_4871,In_620,In_580);
and U4872 (N_4872,In_895,In_49);
or U4873 (N_4873,In_367,In_235);
and U4874 (N_4874,In_847,In_885);
nand U4875 (N_4875,In_390,In_47);
or U4876 (N_4876,In_317,In_75);
and U4877 (N_4877,In_227,In_398);
nor U4878 (N_4878,In_889,In_656);
and U4879 (N_4879,In_698,In_607);
or U4880 (N_4880,In_631,In_750);
nand U4881 (N_4881,In_864,In_611);
nor U4882 (N_4882,In_387,In_462);
or U4883 (N_4883,In_148,In_563);
or U4884 (N_4884,In_196,In_444);
nand U4885 (N_4885,In_576,In_259);
or U4886 (N_4886,In_145,In_879);
nand U4887 (N_4887,In_910,In_86);
and U4888 (N_4888,In_859,In_858);
or U4889 (N_4889,In_951,In_299);
nor U4890 (N_4890,In_362,In_229);
and U4891 (N_4891,In_403,In_451);
nor U4892 (N_4892,In_176,In_564);
or U4893 (N_4893,In_190,In_2);
or U4894 (N_4894,In_672,In_255);
and U4895 (N_4895,In_180,In_419);
nor U4896 (N_4896,In_186,In_460);
nor U4897 (N_4897,In_474,In_847);
and U4898 (N_4898,In_589,In_739);
nand U4899 (N_4899,In_89,In_413);
nor U4900 (N_4900,In_774,In_456);
or U4901 (N_4901,In_653,In_508);
nand U4902 (N_4902,In_482,In_274);
nand U4903 (N_4903,In_396,In_914);
nand U4904 (N_4904,In_298,In_983);
or U4905 (N_4905,In_948,In_448);
or U4906 (N_4906,In_500,In_933);
or U4907 (N_4907,In_52,In_284);
nor U4908 (N_4908,In_232,In_697);
and U4909 (N_4909,In_690,In_607);
nand U4910 (N_4910,In_715,In_584);
and U4911 (N_4911,In_473,In_808);
nand U4912 (N_4912,In_51,In_999);
and U4913 (N_4913,In_51,In_526);
xor U4914 (N_4914,In_954,In_702);
nor U4915 (N_4915,In_578,In_3);
and U4916 (N_4916,In_729,In_21);
nand U4917 (N_4917,In_92,In_687);
or U4918 (N_4918,In_47,In_732);
nor U4919 (N_4919,In_440,In_993);
and U4920 (N_4920,In_183,In_59);
nor U4921 (N_4921,In_548,In_382);
nor U4922 (N_4922,In_845,In_168);
nand U4923 (N_4923,In_642,In_592);
and U4924 (N_4924,In_138,In_178);
nand U4925 (N_4925,In_934,In_3);
nor U4926 (N_4926,In_366,In_979);
nor U4927 (N_4927,In_891,In_334);
or U4928 (N_4928,In_817,In_730);
or U4929 (N_4929,In_262,In_990);
nand U4930 (N_4930,In_123,In_777);
or U4931 (N_4931,In_821,In_252);
nor U4932 (N_4932,In_166,In_984);
or U4933 (N_4933,In_994,In_999);
and U4934 (N_4934,In_376,In_300);
and U4935 (N_4935,In_115,In_678);
or U4936 (N_4936,In_811,In_959);
nand U4937 (N_4937,In_835,In_218);
and U4938 (N_4938,In_117,In_396);
nor U4939 (N_4939,In_698,In_661);
nand U4940 (N_4940,In_826,In_585);
nand U4941 (N_4941,In_221,In_488);
nand U4942 (N_4942,In_858,In_205);
and U4943 (N_4943,In_600,In_787);
nand U4944 (N_4944,In_927,In_360);
nand U4945 (N_4945,In_663,In_371);
nand U4946 (N_4946,In_293,In_46);
or U4947 (N_4947,In_648,In_696);
and U4948 (N_4948,In_124,In_615);
or U4949 (N_4949,In_894,In_694);
and U4950 (N_4950,In_354,In_969);
or U4951 (N_4951,In_853,In_681);
or U4952 (N_4952,In_225,In_953);
nor U4953 (N_4953,In_22,In_866);
nand U4954 (N_4954,In_541,In_870);
or U4955 (N_4955,In_279,In_967);
and U4956 (N_4956,In_930,In_780);
and U4957 (N_4957,In_752,In_658);
nand U4958 (N_4958,In_506,In_314);
and U4959 (N_4959,In_584,In_137);
nor U4960 (N_4960,In_39,In_65);
and U4961 (N_4961,In_638,In_988);
nand U4962 (N_4962,In_243,In_797);
or U4963 (N_4963,In_734,In_65);
nor U4964 (N_4964,In_401,In_888);
nand U4965 (N_4965,In_463,In_243);
nand U4966 (N_4966,In_424,In_292);
or U4967 (N_4967,In_175,In_994);
or U4968 (N_4968,In_970,In_983);
nand U4969 (N_4969,In_868,In_372);
and U4970 (N_4970,In_865,In_717);
or U4971 (N_4971,In_494,In_938);
nand U4972 (N_4972,In_980,In_801);
or U4973 (N_4973,In_931,In_633);
nand U4974 (N_4974,In_268,In_156);
nor U4975 (N_4975,In_362,In_70);
or U4976 (N_4976,In_815,In_49);
nand U4977 (N_4977,In_883,In_750);
or U4978 (N_4978,In_756,In_158);
and U4979 (N_4979,In_593,In_38);
xor U4980 (N_4980,In_276,In_55);
nand U4981 (N_4981,In_33,In_37);
and U4982 (N_4982,In_153,In_270);
nand U4983 (N_4983,In_556,In_388);
nand U4984 (N_4984,In_579,In_359);
and U4985 (N_4985,In_669,In_626);
xor U4986 (N_4986,In_923,In_750);
nor U4987 (N_4987,In_602,In_364);
and U4988 (N_4988,In_366,In_380);
xnor U4989 (N_4989,In_443,In_104);
or U4990 (N_4990,In_911,In_863);
nand U4991 (N_4991,In_817,In_78);
nor U4992 (N_4992,In_664,In_296);
nand U4993 (N_4993,In_738,In_408);
nand U4994 (N_4994,In_590,In_786);
nand U4995 (N_4995,In_456,In_803);
nand U4996 (N_4996,In_441,In_50);
nor U4997 (N_4997,In_333,In_999);
xnor U4998 (N_4998,In_248,In_860);
or U4999 (N_4999,In_729,In_757);
nor U5000 (N_5000,N_2765,N_1843);
and U5001 (N_5001,N_3160,N_1116);
nand U5002 (N_5002,N_2347,N_2191);
or U5003 (N_5003,N_1575,N_3565);
and U5004 (N_5004,N_2965,N_1158);
nor U5005 (N_5005,N_4666,N_929);
and U5006 (N_5006,N_3383,N_2097);
and U5007 (N_5007,N_3562,N_2818);
and U5008 (N_5008,N_128,N_3749);
and U5009 (N_5009,N_748,N_353);
nand U5010 (N_5010,N_3816,N_3260);
or U5011 (N_5011,N_2015,N_3020);
or U5012 (N_5012,N_3857,N_3585);
and U5013 (N_5013,N_2859,N_4774);
and U5014 (N_5014,N_3985,N_1239);
and U5015 (N_5015,N_1052,N_3662);
nand U5016 (N_5016,N_1975,N_2138);
nand U5017 (N_5017,N_1324,N_4271);
nand U5018 (N_5018,N_1812,N_572);
and U5019 (N_5019,N_4218,N_513);
and U5020 (N_5020,N_472,N_4763);
nor U5021 (N_5021,N_673,N_4315);
nor U5022 (N_5022,N_1183,N_991);
nand U5023 (N_5023,N_385,N_4831);
nand U5024 (N_5024,N_4952,N_3616);
and U5025 (N_5025,N_3878,N_606);
nor U5026 (N_5026,N_1980,N_4237);
and U5027 (N_5027,N_2189,N_1279);
nand U5028 (N_5028,N_1300,N_517);
nand U5029 (N_5029,N_3079,N_3472);
nand U5030 (N_5030,N_2021,N_1780);
nand U5031 (N_5031,N_4712,N_2306);
or U5032 (N_5032,N_1261,N_3650);
or U5033 (N_5033,N_1177,N_4746);
nor U5034 (N_5034,N_3492,N_800);
or U5035 (N_5035,N_1049,N_1182);
or U5036 (N_5036,N_2889,N_30);
or U5037 (N_5037,N_2124,N_682);
and U5038 (N_5038,N_2041,N_1649);
nor U5039 (N_5039,N_817,N_2778);
nand U5040 (N_5040,N_2581,N_3009);
and U5041 (N_5041,N_1312,N_2327);
nor U5042 (N_5042,N_1664,N_837);
nor U5043 (N_5043,N_3950,N_2146);
or U5044 (N_5044,N_721,N_4032);
nand U5045 (N_5045,N_50,N_1817);
nor U5046 (N_5046,N_3428,N_4299);
or U5047 (N_5047,N_4996,N_3931);
and U5048 (N_5048,N_2266,N_2577);
and U5049 (N_5049,N_4071,N_1581);
nor U5050 (N_5050,N_3338,N_958);
and U5051 (N_5051,N_1631,N_3213);
nor U5052 (N_5052,N_822,N_4717);
nand U5053 (N_5053,N_4025,N_724);
nand U5054 (N_5054,N_4513,N_631);
and U5055 (N_5055,N_199,N_3192);
nand U5056 (N_5056,N_4878,N_781);
nor U5057 (N_5057,N_2722,N_4859);
nand U5058 (N_5058,N_446,N_1321);
or U5059 (N_5059,N_3015,N_409);
nor U5060 (N_5060,N_1090,N_2231);
nand U5061 (N_5061,N_4877,N_4749);
or U5062 (N_5062,N_2394,N_2708);
nor U5063 (N_5063,N_1006,N_1978);
nand U5064 (N_5064,N_200,N_1908);
or U5065 (N_5065,N_4053,N_2369);
and U5066 (N_5066,N_1128,N_1462);
or U5067 (N_5067,N_300,N_3342);
nand U5068 (N_5068,N_247,N_4214);
nand U5069 (N_5069,N_4034,N_19);
or U5070 (N_5070,N_1289,N_1651);
or U5071 (N_5071,N_3830,N_536);
or U5072 (N_5072,N_3324,N_2739);
nand U5073 (N_5073,N_4362,N_426);
and U5074 (N_5074,N_3803,N_4829);
or U5075 (N_5075,N_1373,N_2955);
nand U5076 (N_5076,N_2193,N_4103);
or U5077 (N_5077,N_2538,N_3457);
and U5078 (N_5078,N_2142,N_1751);
or U5079 (N_5079,N_4139,N_2961);
or U5080 (N_5080,N_1991,N_2058);
nor U5081 (N_5081,N_4597,N_4393);
nand U5082 (N_5082,N_4059,N_2157);
and U5083 (N_5083,N_4044,N_4659);
nor U5084 (N_5084,N_3559,N_2313);
or U5085 (N_5085,N_1240,N_547);
or U5086 (N_5086,N_4262,N_1486);
or U5087 (N_5087,N_3129,N_1816);
nand U5088 (N_5088,N_1837,N_576);
and U5089 (N_5089,N_862,N_311);
or U5090 (N_5090,N_998,N_3082);
or U5091 (N_5091,N_3867,N_3994);
and U5092 (N_5092,N_4502,N_1074);
nor U5093 (N_5093,N_1915,N_440);
or U5094 (N_5094,N_753,N_3843);
and U5095 (N_5095,N_1446,N_610);
nand U5096 (N_5096,N_1684,N_3016);
nor U5097 (N_5097,N_3511,N_491);
or U5098 (N_5098,N_3879,N_3360);
and U5099 (N_5099,N_4165,N_236);
and U5100 (N_5100,N_769,N_183);
nand U5101 (N_5101,N_1126,N_4799);
and U5102 (N_5102,N_1635,N_55);
nor U5103 (N_5103,N_1277,N_1734);
or U5104 (N_5104,N_1459,N_2563);
or U5105 (N_5105,N_672,N_968);
and U5106 (N_5106,N_256,N_4110);
and U5107 (N_5107,N_2329,N_4111);
or U5108 (N_5108,N_4445,N_3050);
nor U5109 (N_5109,N_4000,N_1850);
or U5110 (N_5110,N_3651,N_4121);
nor U5111 (N_5111,N_1112,N_4084);
nand U5112 (N_5112,N_2701,N_3914);
and U5113 (N_5113,N_4402,N_3486);
nor U5114 (N_5114,N_3707,N_2683);
or U5115 (N_5115,N_592,N_2805);
and U5116 (N_5116,N_3032,N_2448);
and U5117 (N_5117,N_511,N_4089);
or U5118 (N_5118,N_8,N_4838);
and U5119 (N_5119,N_2880,N_2596);
or U5120 (N_5120,N_4474,N_3370);
and U5121 (N_5121,N_3400,N_4215);
nand U5122 (N_5122,N_2413,N_96);
or U5123 (N_5123,N_4368,N_2526);
nor U5124 (N_5124,N_3422,N_3150);
nand U5125 (N_5125,N_1223,N_402);
nand U5126 (N_5126,N_3633,N_2046);
or U5127 (N_5127,N_1318,N_4327);
and U5128 (N_5128,N_1609,N_4684);
and U5129 (N_5129,N_4897,N_3885);
nor U5130 (N_5130,N_2429,N_4702);
nor U5131 (N_5131,N_3097,N_1093);
nor U5132 (N_5132,N_4989,N_3109);
nor U5133 (N_5133,N_2482,N_3584);
and U5134 (N_5134,N_1395,N_2901);
or U5135 (N_5135,N_562,N_2235);
or U5136 (N_5136,N_427,N_2451);
nor U5137 (N_5137,N_1208,N_1473);
and U5138 (N_5138,N_1701,N_3941);
nor U5139 (N_5139,N_3283,N_3410);
nand U5140 (N_5140,N_4510,N_543);
or U5141 (N_5141,N_3574,N_2198);
and U5142 (N_5142,N_3561,N_146);
xor U5143 (N_5143,N_4933,N_4867);
nor U5144 (N_5144,N_1372,N_1622);
or U5145 (N_5145,N_2381,N_3452);
nor U5146 (N_5146,N_3946,N_3627);
nand U5147 (N_5147,N_3365,N_4696);
nand U5148 (N_5148,N_1759,N_4258);
nand U5149 (N_5149,N_3233,N_3987);
or U5150 (N_5150,N_1970,N_2207);
nor U5151 (N_5151,N_2111,N_3144);
nand U5152 (N_5152,N_3025,N_3421);
nor U5153 (N_5153,N_1385,N_3376);
nor U5154 (N_5154,N_2492,N_3450);
or U5155 (N_5155,N_2152,N_886);
or U5156 (N_5156,N_1347,N_3958);
and U5157 (N_5157,N_4586,N_2192);
nand U5158 (N_5158,N_2917,N_2171);
or U5159 (N_5159,N_372,N_4546);
nor U5160 (N_5160,N_4055,N_398);
or U5161 (N_5161,N_1207,N_2332);
nand U5162 (N_5162,N_4431,N_1465);
and U5163 (N_5163,N_4890,N_4718);
nor U5164 (N_5164,N_561,N_2209);
or U5165 (N_5165,N_681,N_838);
or U5166 (N_5166,N_1016,N_4954);
nor U5167 (N_5167,N_2996,N_453);
nor U5168 (N_5168,N_3766,N_3928);
or U5169 (N_5169,N_1353,N_4574);
or U5170 (N_5170,N_1165,N_4429);
or U5171 (N_5171,N_4051,N_4275);
or U5172 (N_5172,N_4419,N_1345);
nor U5173 (N_5173,N_2617,N_3459);
nor U5174 (N_5174,N_2629,N_3877);
and U5175 (N_5175,N_888,N_4359);
xnor U5176 (N_5176,N_2618,N_2280);
nor U5177 (N_5177,N_2582,N_3845);
nor U5178 (N_5178,N_4043,N_2364);
or U5179 (N_5179,N_451,N_2325);
or U5180 (N_5180,N_819,N_1466);
nand U5181 (N_5181,N_4832,N_2031);
or U5182 (N_5182,N_2864,N_4353);
and U5183 (N_5183,N_1351,N_2789);
or U5184 (N_5184,N_4150,N_734);
nand U5185 (N_5185,N_2499,N_1648);
and U5186 (N_5186,N_4776,N_979);
nand U5187 (N_5187,N_4968,N_4576);
nor U5188 (N_5188,N_4547,N_4222);
and U5189 (N_5189,N_1808,N_4013);
and U5190 (N_5190,N_3060,N_3299);
nand U5191 (N_5191,N_3959,N_2087);
and U5192 (N_5192,N_4822,N_4664);
nor U5193 (N_5193,N_645,N_3688);
nand U5194 (N_5194,N_1705,N_4489);
nor U5195 (N_5195,N_2262,N_2139);
nor U5196 (N_5196,N_3146,N_2084);
nand U5197 (N_5197,N_1425,N_4078);
nand U5198 (N_5198,N_990,N_1911);
and U5199 (N_5199,N_826,N_2348);
nand U5200 (N_5200,N_1814,N_4906);
or U5201 (N_5201,N_1845,N_456);
nand U5202 (N_5202,N_1500,N_3273);
or U5203 (N_5203,N_266,N_2853);
nor U5204 (N_5204,N_3489,N_500);
nor U5205 (N_5205,N_2587,N_1679);
nor U5206 (N_5206,N_1480,N_2745);
and U5207 (N_5207,N_4918,N_1402);
nand U5208 (N_5208,N_1452,N_2892);
and U5209 (N_5209,N_2841,N_404);
or U5210 (N_5210,N_4754,N_4980);
or U5211 (N_5211,N_4660,N_4300);
and U5212 (N_5212,N_3770,N_330);
nor U5213 (N_5213,N_3251,N_4852);
nand U5214 (N_5214,N_772,N_930);
xor U5215 (N_5215,N_714,N_770);
and U5216 (N_5216,N_1543,N_3403);
nor U5217 (N_5217,N_3840,N_367);
or U5218 (N_5218,N_3323,N_1572);
and U5219 (N_5219,N_2958,N_2439);
or U5220 (N_5220,N_4066,N_4261);
or U5221 (N_5221,N_133,N_4594);
nand U5222 (N_5222,N_4475,N_1520);
nor U5223 (N_5223,N_4973,N_1134);
or U5224 (N_5224,N_157,N_4565);
and U5225 (N_5225,N_322,N_2500);
and U5226 (N_5226,N_1797,N_594);
nand U5227 (N_5227,N_2574,N_2260);
nand U5228 (N_5228,N_413,N_1589);
nand U5229 (N_5229,N_2383,N_3141);
or U5230 (N_5230,N_2102,N_1085);
or U5231 (N_5231,N_4142,N_4658);
nor U5232 (N_5232,N_864,N_4179);
nor U5233 (N_5233,N_1528,N_2375);
or U5234 (N_5234,N_2456,N_2076);
nand U5235 (N_5235,N_3173,N_3963);
nand U5236 (N_5236,N_3970,N_739);
or U5237 (N_5237,N_3152,N_358);
or U5238 (N_5238,N_1636,N_2599);
nor U5239 (N_5239,N_1083,N_2743);
or U5240 (N_5240,N_1327,N_3405);
or U5241 (N_5241,N_1731,N_1795);
nor U5242 (N_5242,N_845,N_1031);
nand U5243 (N_5243,N_4620,N_3257);
and U5244 (N_5244,N_712,N_246);
nor U5245 (N_5245,N_602,N_4416);
nand U5246 (N_5246,N_1450,N_4585);
or U5247 (N_5247,N_2363,N_2893);
or U5248 (N_5248,N_3143,N_4579);
xnor U5249 (N_5249,N_4983,N_393);
and U5250 (N_5250,N_2975,N_2672);
and U5251 (N_5251,N_337,N_963);
or U5252 (N_5252,N_3256,N_988);
or U5253 (N_5253,N_4881,N_1941);
nor U5254 (N_5254,N_3654,N_595);
or U5255 (N_5255,N_112,N_1089);
nor U5256 (N_5256,N_468,N_969);
and U5257 (N_5257,N_3200,N_4770);
nor U5258 (N_5258,N_972,N_2398);
nand U5259 (N_5259,N_3350,N_601);
and U5260 (N_5260,N_3480,N_3859);
or U5261 (N_5261,N_3021,N_4926);
nor U5262 (N_5262,N_477,N_3435);
nand U5263 (N_5263,N_3617,N_4638);
and U5264 (N_5264,N_2547,N_531);
nor U5265 (N_5265,N_1955,N_3634);
and U5266 (N_5266,N_1346,N_4540);
or U5267 (N_5267,N_3898,N_4714);
nor U5268 (N_5268,N_2253,N_2529);
nand U5269 (N_5269,N_2099,N_4534);
nand U5270 (N_5270,N_4313,N_3753);
nor U5271 (N_5271,N_2643,N_3449);
and U5272 (N_5272,N_801,N_3530);
nand U5273 (N_5273,N_4760,N_1214);
or U5274 (N_5274,N_2150,N_3301);
or U5275 (N_5275,N_1639,N_4241);
and U5276 (N_5276,N_1906,N_2452);
or U5277 (N_5277,N_213,N_3085);
and U5278 (N_5278,N_2872,N_3099);
nand U5279 (N_5279,N_3953,N_774);
and U5280 (N_5280,N_3521,N_3929);
and U5281 (N_5281,N_2852,N_2963);
nor U5282 (N_5282,N_867,N_4971);
nand U5283 (N_5283,N_1786,N_4285);
and U5284 (N_5284,N_3075,N_1519);
or U5285 (N_5285,N_613,N_853);
nor U5286 (N_5286,N_3269,N_2552);
nor U5287 (N_5287,N_2704,N_4135);
nand U5288 (N_5288,N_827,N_4951);
nor U5289 (N_5289,N_399,N_235);
nor U5290 (N_5290,N_2758,N_3613);
or U5291 (N_5291,N_1272,N_3871);
nor U5292 (N_5292,N_1606,N_1907);
nand U5293 (N_5293,N_4719,N_4999);
nand U5294 (N_5294,N_657,N_2432);
nor U5295 (N_5295,N_3829,N_1073);
nand U5296 (N_5296,N_539,N_1996);
nor U5297 (N_5297,N_943,N_2871);
nand U5298 (N_5298,N_2940,N_2803);
nand U5299 (N_5299,N_2395,N_4598);
or U5300 (N_5300,N_1719,N_4766);
and U5301 (N_5301,N_3033,N_3258);
and U5302 (N_5302,N_1698,N_956);
or U5303 (N_5303,N_4872,N_1139);
nor U5304 (N_5304,N_691,N_2894);
and U5305 (N_5305,N_737,N_3884);
nor U5306 (N_5306,N_1971,N_1894);
and U5307 (N_5307,N_3102,N_1896);
and U5308 (N_5308,N_2811,N_3208);
and U5309 (N_5309,N_354,N_3820);
nor U5310 (N_5310,N_578,N_570);
and U5311 (N_5311,N_622,N_614);
nand U5312 (N_5312,N_1594,N_263);
nor U5313 (N_5313,N_1718,N_4372);
nand U5314 (N_5314,N_3755,N_4942);
or U5315 (N_5315,N_1824,N_2341);
or U5316 (N_5316,N_1789,N_3682);
xnor U5317 (N_5317,N_34,N_381);
or U5318 (N_5318,N_3469,N_1947);
nand U5319 (N_5319,N_4703,N_3606);
or U5320 (N_5320,N_885,N_2378);
nand U5321 (N_5321,N_3372,N_1204);
or U5322 (N_5322,N_4946,N_1762);
or U5323 (N_5323,N_277,N_3197);
and U5324 (N_5324,N_2952,N_1454);
nor U5325 (N_5325,N_2312,N_2457);
or U5326 (N_5326,N_2184,N_1133);
nor U5327 (N_5327,N_4675,N_2173);
and U5328 (N_5328,N_102,N_2918);
nand U5329 (N_5329,N_4512,N_1009);
nor U5330 (N_5330,N_1711,N_4750);
nor U5331 (N_5331,N_2750,N_455);
nand U5332 (N_5332,N_4736,N_1494);
nand U5333 (N_5333,N_2026,N_3503);
nand U5334 (N_5334,N_1417,N_3702);
nor U5335 (N_5335,N_75,N_492);
nand U5336 (N_5336,N_662,N_2767);
and U5337 (N_5337,N_3703,N_2588);
nor U5338 (N_5338,N_4289,N_3069);
nand U5339 (N_5339,N_2977,N_3215);
nand U5340 (N_5340,N_1325,N_4167);
nand U5341 (N_5341,N_1923,N_1655);
or U5342 (N_5342,N_3206,N_145);
nand U5343 (N_5343,N_4081,N_2621);
nor U5344 (N_5344,N_3356,N_2830);
nor U5345 (N_5345,N_4470,N_4833);
nor U5346 (N_5346,N_2120,N_828);
and U5347 (N_5347,N_176,N_43);
or U5348 (N_5348,N_416,N_3842);
and U5349 (N_5349,N_1316,N_1378);
nor U5350 (N_5350,N_883,N_3664);
and U5351 (N_5351,N_3599,N_11);
nor U5352 (N_5352,N_4338,N_2244);
or U5353 (N_5353,N_1953,N_3722);
or U5354 (N_5354,N_2211,N_2783);
and U5355 (N_5355,N_4813,N_4154);
nor U5356 (N_5356,N_3321,N_1984);
and U5357 (N_5357,N_2453,N_3673);
nand U5358 (N_5358,N_1764,N_1926);
or U5359 (N_5359,N_4132,N_2277);
nor U5360 (N_5360,N_4782,N_3618);
or U5361 (N_5361,N_1497,N_1369);
or U5362 (N_5362,N_3547,N_4217);
and U5363 (N_5363,N_482,N_2247);
xor U5364 (N_5364,N_4708,N_1043);
nor U5365 (N_5365,N_1666,N_3346);
or U5366 (N_5366,N_3474,N_1833);
nand U5367 (N_5367,N_3727,N_1106);
nor U5368 (N_5368,N_3937,N_764);
nor U5369 (N_5369,N_1173,N_3769);
and U5370 (N_5370,N_2914,N_4681);
or U5371 (N_5371,N_4633,N_2685);
or U5372 (N_5372,N_2490,N_3539);
and U5373 (N_5373,N_4373,N_4907);
nand U5374 (N_5374,N_3303,N_121);
xor U5375 (N_5375,N_670,N_4757);
and U5376 (N_5376,N_3757,N_3322);
nor U5377 (N_5377,N_3636,N_2678);
or U5378 (N_5378,N_412,N_1196);
and U5379 (N_5379,N_88,N_3359);
and U5380 (N_5380,N_3,N_3989);
or U5381 (N_5381,N_2697,N_2705);
nor U5382 (N_5382,N_2151,N_4922);
and U5383 (N_5383,N_255,N_3858);
or U5384 (N_5384,N_1107,N_4269);
and U5385 (N_5385,N_4152,N_2328);
and U5386 (N_5386,N_2402,N_421);
or U5387 (N_5387,N_2731,N_741);
nor U5388 (N_5388,N_3437,N_2649);
nand U5389 (N_5389,N_1060,N_2707);
nand U5390 (N_5390,N_4558,N_2507);
and U5391 (N_5391,N_2674,N_3741);
nand U5392 (N_5392,N_3164,N_73);
or U5393 (N_5393,N_1026,N_1782);
and U5394 (N_5394,N_1460,N_140);
nand U5395 (N_5395,N_6,N_107);
nor U5396 (N_5396,N_4380,N_1171);
nor U5397 (N_5397,N_467,N_4496);
and U5398 (N_5398,N_4065,N_857);
xnor U5399 (N_5399,N_3477,N_4888);
and U5400 (N_5400,N_2520,N_2278);
or U5401 (N_5401,N_4188,N_4521);
and U5402 (N_5402,N_4169,N_3398);
nor U5403 (N_5403,N_4136,N_3005);
and U5404 (N_5404,N_175,N_2806);
and U5405 (N_5405,N_1769,N_3187);
or U5406 (N_5406,N_967,N_2733);
nand U5407 (N_5407,N_4420,N_1766);
and U5408 (N_5408,N_4628,N_3710);
or U5409 (N_5409,N_4934,N_4570);
or U5410 (N_5410,N_2223,N_1358);
nand U5411 (N_5411,N_1265,N_3775);
nor U5412 (N_5412,N_3748,N_299);
or U5413 (N_5413,N_1146,N_2968);
nor U5414 (N_5414,N_2256,N_1331);
nor U5415 (N_5415,N_2090,N_2673);
or U5416 (N_5416,N_2790,N_1835);
and U5417 (N_5417,N_3776,N_2236);
nand U5418 (N_5418,N_3542,N_1281);
or U5419 (N_5419,N_2530,N_167);
or U5420 (N_5420,N_4069,N_2167);
nand U5421 (N_5421,N_2155,N_1340);
or U5422 (N_5422,N_1244,N_3681);
and U5423 (N_5423,N_620,N_51);
nor U5424 (N_5424,N_2075,N_3479);
or U5425 (N_5425,N_2195,N_2634);
nand U5426 (N_5426,N_4566,N_4722);
and U5427 (N_5427,N_4015,N_108);
and U5428 (N_5428,N_2792,N_3527);
or U5429 (N_5429,N_1976,N_4254);
and U5430 (N_5430,N_4387,N_2445);
nor U5431 (N_5431,N_4438,N_2980);
nand U5432 (N_5432,N_2768,N_3546);
nand U5433 (N_5433,N_3620,N_900);
and U5434 (N_5434,N_2506,N_312);
nor U5435 (N_5435,N_1754,N_3579);
or U5436 (N_5436,N_4350,N_54);
nand U5437 (N_5437,N_884,N_3524);
nor U5438 (N_5438,N_4147,N_47);
or U5439 (N_5439,N_1067,N_3185);
nand U5440 (N_5440,N_4469,N_805);
nand U5441 (N_5441,N_2459,N_1199);
nand U5442 (N_5442,N_4201,N_2289);
nor U5443 (N_5443,N_3481,N_4609);
and U5444 (N_5444,N_4472,N_4936);
nand U5445 (N_5445,N_1038,N_515);
xnor U5446 (N_5446,N_3059,N_1053);
or U5447 (N_5447,N_814,N_2062);
and U5448 (N_5448,N_3487,N_4392);
nor U5449 (N_5449,N_3210,N_787);
nand U5450 (N_5450,N_4182,N_4711);
nor U5451 (N_5451,N_4086,N_3343);
or U5452 (N_5452,N_441,N_600);
and U5453 (N_5453,N_2091,N_1348);
nand U5454 (N_5454,N_3309,N_1582);
or U5455 (N_5455,N_1296,N_3715);
nand U5456 (N_5456,N_2870,N_201);
and U5457 (N_5457,N_2094,N_4274);
or U5458 (N_5458,N_1379,N_2639);
or U5459 (N_5459,N_4482,N_2929);
nand U5460 (N_5460,N_1806,N_1891);
or U5461 (N_5461,N_4742,N_2764);
and U5462 (N_5462,N_3084,N_866);
or U5463 (N_5463,N_326,N_3183);
and U5464 (N_5464,N_4840,N_1504);
or U5465 (N_5465,N_3984,N_4582);
and U5466 (N_5466,N_4564,N_4191);
nor U5467 (N_5467,N_665,N_3207);
and U5468 (N_5468,N_3096,N_4276);
and U5469 (N_5469,N_2950,N_98);
or U5470 (N_5470,N_591,N_1662);
nand U5471 (N_5471,N_2680,N_3483);
or U5472 (N_5472,N_2989,N_4531);
nor U5473 (N_5473,N_2884,N_3010);
nor U5474 (N_5474,N_2291,N_1401);
nand U5475 (N_5475,N_2935,N_3880);
xor U5476 (N_5476,N_4197,N_3534);
nand U5477 (N_5477,N_2351,N_3981);
or U5478 (N_5478,N_1015,N_1405);
nand U5479 (N_5479,N_2447,N_3625);
and U5480 (N_5480,N_483,N_4287);
nor U5481 (N_5481,N_2744,N_4264);
and U5482 (N_5482,N_1418,N_3860);
nand U5483 (N_5483,N_2073,N_4138);
nor U5484 (N_5484,N_4771,N_935);
nor U5485 (N_5485,N_2791,N_4932);
or U5486 (N_5486,N_3999,N_1374);
and U5487 (N_5487,N_1579,N_668);
nor U5488 (N_5488,N_3232,N_3712);
and U5489 (N_5489,N_2480,N_3191);
and U5490 (N_5490,N_1632,N_1691);
nand U5491 (N_5491,N_3866,N_4875);
nand U5492 (N_5492,N_549,N_3965);
and U5493 (N_5493,N_792,N_1935);
nor U5494 (N_5494,N_1467,N_4621);
or U5495 (N_5495,N_4707,N_4375);
nor U5496 (N_5496,N_4383,N_3238);
or U5497 (N_5497,N_2470,N_4593);
or U5498 (N_5498,N_340,N_2959);
or U5499 (N_5499,N_4505,N_420);
and U5500 (N_5500,N_788,N_3761);
nor U5501 (N_5501,N_4654,N_2125);
nand U5502 (N_5502,N_1097,N_3116);
and U5503 (N_5503,N_3091,N_1298);
or U5504 (N_5504,N_2298,N_2772);
nor U5505 (N_5505,N_4140,N_2367);
nand U5506 (N_5506,N_3348,N_2515);
nand U5507 (N_5507,N_2164,N_2716);
or U5508 (N_5508,N_3882,N_177);
and U5509 (N_5509,N_2122,N_3944);
nor U5510 (N_5510,N_1209,N_4526);
or U5511 (N_5511,N_25,N_2873);
or U5512 (N_5512,N_4239,N_1578);
nand U5513 (N_5513,N_447,N_669);
nor U5514 (N_5514,N_2798,N_2337);
and U5515 (N_5515,N_1903,N_2135);
nor U5516 (N_5516,N_29,N_675);
and U5517 (N_5517,N_623,N_2408);
nor U5518 (N_5518,N_2237,N_1860);
nand U5519 (N_5519,N_3224,N_400);
and U5520 (N_5520,N_3508,N_3123);
nor U5521 (N_5521,N_2134,N_3949);
nand U5522 (N_5522,N_2905,N_795);
nor U5523 (N_5523,N_3319,N_2147);
nand U5524 (N_5524,N_452,N_3926);
nand U5525 (N_5525,N_1939,N_221);
or U5526 (N_5526,N_1542,N_23);
or U5527 (N_5527,N_727,N_2902);
xor U5528 (N_5528,N_4243,N_987);
nand U5529 (N_5529,N_3042,N_1895);
nand U5530 (N_5530,N_3281,N_1304);
nand U5531 (N_5531,N_3093,N_1027);
or U5532 (N_5532,N_1933,N_4483);
and U5533 (N_5533,N_2801,N_345);
nand U5534 (N_5534,N_3728,N_3001);
nand U5535 (N_5535,N_2360,N_3725);
and U5536 (N_5536,N_2808,N_3386);
nand U5537 (N_5537,N_2655,N_4480);
xnor U5538 (N_5538,N_4204,N_2850);
or U5539 (N_5539,N_746,N_1142);
or U5540 (N_5540,N_4137,N_245);
nor U5541 (N_5541,N_1757,N_4561);
and U5542 (N_5542,N_4058,N_1853);
nor U5543 (N_5543,N_2276,N_696);
or U5544 (N_5544,N_4231,N_2458);
and U5545 (N_5545,N_4964,N_2454);
nand U5546 (N_5546,N_4186,N_1952);
nand U5547 (N_5547,N_2982,N_3935);
nand U5548 (N_5548,N_3700,N_4166);
nand U5549 (N_5549,N_1387,N_3073);
nand U5550 (N_5550,N_571,N_4583);
nor U5551 (N_5551,N_2344,N_4097);
and U5552 (N_5552,N_135,N_1120);
nor U5553 (N_5553,N_3894,N_3611);
nor U5554 (N_5554,N_4894,N_4109);
nand U5555 (N_5555,N_486,N_3968);
or U5556 (N_5556,N_3029,N_4676);
nand U5557 (N_5557,N_4921,N_3196);
nand U5558 (N_5558,N_2477,N_2340);
or U5559 (N_5559,N_2194,N_3156);
nor U5560 (N_5560,N_368,N_2051);
nand U5561 (N_5561,N_3120,N_4298);
nor U5562 (N_5562,N_2392,N_1036);
nor U5563 (N_5563,N_940,N_1934);
nand U5564 (N_5564,N_2407,N_142);
nand U5565 (N_5565,N_2342,N_4796);
or U5566 (N_5566,N_2695,N_3220);
or U5567 (N_5567,N_4690,N_4733);
nor U5568 (N_5568,N_2187,N_2305);
nor U5569 (N_5569,N_2810,N_4661);
nor U5570 (N_5570,N_4709,N_2724);
or U5571 (N_5571,N_425,N_626);
nand U5572 (N_5572,N_2620,N_3754);
or U5573 (N_5573,N_2269,N_1741);
and U5574 (N_5574,N_435,N_2030);
or U5575 (N_5575,N_4550,N_4543);
or U5576 (N_5576,N_2624,N_4716);
or U5577 (N_5577,N_58,N_2263);
or U5578 (N_5578,N_1195,N_2773);
and U5579 (N_5579,N_3638,N_3558);
or U5580 (N_5580,N_2938,N_210);
nor U5581 (N_5581,N_3337,N_2865);
and U5582 (N_5582,N_545,N_2436);
nand U5583 (N_5583,N_1966,N_2887);
nor U5584 (N_5584,N_1874,N_3750);
or U5585 (N_5585,N_298,N_193);
or U5586 (N_5586,N_803,N_627);
or U5587 (N_5587,N_3013,N_3475);
and U5588 (N_5588,N_4575,N_3827);
nor U5589 (N_5589,N_4417,N_2144);
and U5590 (N_5590,N_2539,N_2330);
or U5591 (N_5591,N_1438,N_2911);
nand U5592 (N_5592,N_1930,N_1212);
nand U5593 (N_5593,N_3752,N_244);
nor U5594 (N_5594,N_1222,N_473);
nor U5595 (N_5595,N_4478,N_4520);
nand U5596 (N_5596,N_2060,N_3805);
or U5597 (N_5597,N_2322,N_2230);
nor U5598 (N_5598,N_2561,N_3122);
nor U5599 (N_5599,N_4747,N_703);
nor U5600 (N_5600,N_1389,N_76);
nand U5601 (N_5601,N_1796,N_3333);
nand U5602 (N_5602,N_3395,N_4366);
nand U5603 (N_5603,N_2424,N_1830);
nor U5604 (N_5604,N_1130,N_3431);
and U5605 (N_5605,N_1001,N_1630);
nor U5606 (N_5606,N_4670,N_3130);
nand U5607 (N_5607,N_679,N_1255);
nand U5608 (N_5608,N_4283,N_1862);
and U5609 (N_5609,N_3876,N_3913);
or U5610 (N_5610,N_4281,N_470);
and U5611 (N_5611,N_3756,N_2537);
or U5612 (N_5612,N_4073,N_824);
nand U5613 (N_5613,N_1230,N_3942);
or U5614 (N_5614,N_2573,N_1070);
nand U5615 (N_5615,N_3510,N_3666);
nor U5616 (N_5616,N_361,N_126);
nand U5617 (N_5617,N_815,N_1129);
or U5618 (N_5618,N_3171,N_351);
and U5619 (N_5619,N_3687,N_1435);
nand U5620 (N_5620,N_1197,N_291);
nand U5621 (N_5621,N_2059,N_360);
nand U5622 (N_5622,N_3920,N_2054);
nand U5623 (N_5623,N_3112,N_2688);
or U5624 (N_5624,N_843,N_1437);
nand U5625 (N_5625,N_2354,N_3195);
and U5626 (N_5626,N_1537,N_1712);
or U5627 (N_5627,N_397,N_2558);
or U5628 (N_5628,N_2721,N_4726);
and U5629 (N_5629,N_1527,N_1088);
nor U5630 (N_5630,N_2576,N_3789);
or U5631 (N_5631,N_914,N_1050);
nand U5632 (N_5632,N_1175,N_282);
nand U5633 (N_5633,N_522,N_702);
or U5634 (N_5634,N_2564,N_676);
nor U5635 (N_5635,N_1997,N_3297);
nand U5636 (N_5636,N_3992,N_1468);
nor U5637 (N_5637,N_3062,N_1022);
nor U5638 (N_5638,N_4815,N_1778);
nor U5639 (N_5639,N_4720,N_4618);
nor U5640 (N_5640,N_569,N_4500);
and U5641 (N_5641,N_1695,N_4022);
nor U5642 (N_5642,N_2825,N_3983);
nor U5643 (N_5643,N_1621,N_2028);
nand U5644 (N_5644,N_2519,N_3847);
nand U5645 (N_5645,N_1118,N_1066);
nand U5646 (N_5646,N_4223,N_4790);
and U5647 (N_5647,N_3433,N_1964);
and U5648 (N_5648,N_3478,N_633);
nand U5649 (N_5649,N_264,N_2593);
or U5650 (N_5650,N_3685,N_1828);
nor U5651 (N_5651,N_1266,N_3869);
or U5652 (N_5652,N_4866,N_3990);
nor U5653 (N_5653,N_3392,N_3267);
nand U5654 (N_5654,N_4553,N_1748);
and U5655 (N_5655,N_418,N_2511);
nand U5656 (N_5656,N_957,N_4629);
nand U5657 (N_5657,N_1071,N_3908);
and U5658 (N_5658,N_1634,N_2279);
and U5659 (N_5659,N_4108,N_2874);
or U5660 (N_5660,N_3051,N_3619);
or U5661 (N_5661,N_2832,N_664);
or U5662 (N_5662,N_1856,N_493);
and U5663 (N_5663,N_1062,N_1852);
and U5664 (N_5664,N_2315,N_3250);
and U5665 (N_5665,N_1918,N_1627);
and U5666 (N_5666,N_4900,N_2579);
nand U5667 (N_5667,N_2181,N_1412);
xor U5668 (N_5668,N_653,N_1203);
nor U5669 (N_5669,N_2441,N_1863);
and U5670 (N_5670,N_4088,N_3295);
nor U5671 (N_5671,N_2216,N_2414);
nand U5672 (N_5672,N_4573,N_4612);
or U5673 (N_5673,N_261,N_1160);
nand U5674 (N_5674,N_1246,N_2834);
nor U5675 (N_5675,N_1322,N_3054);
and U5676 (N_5676,N_3212,N_2132);
and U5677 (N_5677,N_2771,N_1616);
or U5678 (N_5678,N_1888,N_392);
or U5679 (N_5679,N_1993,N_4199);
nand U5680 (N_5680,N_944,N_3991);
nand U5681 (N_5681,N_4895,N_1556);
and U5682 (N_5682,N_2085,N_3278);
or U5683 (N_5683,N_4943,N_4164);
nor U5684 (N_5684,N_2412,N_4114);
or U5685 (N_5685,N_4581,N_2657);
nand U5686 (N_5686,N_3107,N_3603);
and U5687 (N_5687,N_812,N_619);
nand U5688 (N_5688,N_2405,N_1362);
nand U5689 (N_5689,N_3604,N_1729);
nor U5690 (N_5690,N_4950,N_62);
or U5691 (N_5691,N_268,N_2603);
or U5692 (N_5692,N_2096,N_757);
nand U5693 (N_5693,N_2056,N_4792);
nand U5694 (N_5694,N_3810,N_97);
or U5695 (N_5695,N_2960,N_869);
or U5696 (N_5696,N_1242,N_2990);
nor U5697 (N_5697,N_1535,N_3500);
nand U5698 (N_5698,N_2845,N_4422);
nor U5699 (N_5699,N_1638,N_527);
nor U5700 (N_5700,N_3602,N_1601);
and U5701 (N_5701,N_1391,N_2240);
and U5702 (N_5702,N_4325,N_4772);
nand U5703 (N_5703,N_4649,N_2326);
nor U5704 (N_5704,N_542,N_2205);
and U5705 (N_5705,N_1124,N_1761);
and U5706 (N_5706,N_4101,N_87);
and U5707 (N_5707,N_3034,N_364);
or U5708 (N_5708,N_2027,N_4456);
nor U5709 (N_5709,N_1882,N_3589);
nor U5710 (N_5710,N_585,N_3982);
nand U5711 (N_5711,N_3939,N_1722);
nor U5712 (N_5712,N_2815,N_4440);
nor U5713 (N_5713,N_3855,N_2355);
or U5714 (N_5714,N_4653,N_3781);
or U5715 (N_5715,N_374,N_732);
and U5716 (N_5716,N_3158,N_3763);
and U5717 (N_5717,N_39,N_3417);
or U5718 (N_5718,N_3596,N_4865);
nand U5719 (N_5719,N_4322,N_747);
or U5720 (N_5720,N_17,N_730);
and U5721 (N_5721,N_3739,N_1667);
nor U5722 (N_5722,N_2040,N_4640);
nor U5723 (N_5723,N_1206,N_2921);
xnor U5724 (N_5724,N_83,N_1530);
and U5725 (N_5725,N_3671,N_2255);
or U5726 (N_5726,N_3131,N_1111);
and U5727 (N_5727,N_3653,N_3090);
and U5728 (N_5728,N_3986,N_4645);
nor U5729 (N_5729,N_1857,N_851);
nand U5730 (N_5730,N_2523,N_4871);
or U5731 (N_5731,N_1424,N_1104);
nor U5732 (N_5732,N_2709,N_1274);
nand U5733 (N_5733,N_677,N_4826);
nor U5734 (N_5734,N_2010,N_4780);
nor U5735 (N_5735,N_726,N_3169);
nor U5736 (N_5736,N_4057,N_2361);
nor U5737 (N_5737,N_4630,N_3661);
and U5738 (N_5738,N_1685,N_2036);
nand U5739 (N_5739,N_2895,N_2297);
nand U5740 (N_5740,N_2524,N_2345);
nor U5741 (N_5741,N_2023,N_1720);
nand U5742 (N_5742,N_3704,N_265);
and U5743 (N_5743,N_736,N_2148);
nor U5744 (N_5744,N_3699,N_1670);
nand U5745 (N_5745,N_3056,N_1758);
or U5746 (N_5746,N_4447,N_2421);
nor U5747 (N_5747,N_2560,N_2541);
or U5748 (N_5748,N_442,N_2224);
nand U5749 (N_5749,N_92,N_3041);
nand U5750 (N_5750,N_1886,N_3067);
and U5751 (N_5751,N_4376,N_3783);
nand U5752 (N_5752,N_4981,N_3667);
nand U5753 (N_5753,N_2969,N_1827);
and U5754 (N_5754,N_4768,N_1375);
nand U5755 (N_5755,N_3745,N_1045);
nand U5756 (N_5756,N_1471,N_3853);
nor U5757 (N_5757,N_564,N_3167);
nand U5758 (N_5758,N_332,N_4842);
nor U5759 (N_5759,N_2177,N_2159);
or U5760 (N_5760,N_3854,N_2785);
nor U5761 (N_5761,N_323,N_4985);
or U5762 (N_5762,N_3764,N_2004);
and U5763 (N_5763,N_3822,N_683);
and U5764 (N_5764,N_2000,N_2916);
or U5765 (N_5765,N_1644,N_164);
nand U5766 (N_5766,N_1278,N_667);
and U5767 (N_5767,N_2605,N_433);
nor U5768 (N_5768,N_1270,N_1057);
nand U5769 (N_5769,N_804,N_2613);
and U5770 (N_5770,N_1310,N_2664);
or U5771 (N_5771,N_2493,N_3583);
or U5772 (N_5772,N_754,N_4082);
or U5773 (N_5773,N_4614,N_414);
nor U5774 (N_5774,N_42,N_1364);
xor U5775 (N_5775,N_1735,N_1008);
and U5776 (N_5776,N_2714,N_205);
nor U5777 (N_5777,N_4023,N_2284);
nand U5778 (N_5778,N_4787,N_939);
and U5779 (N_5779,N_4104,N_2754);
and U5780 (N_5780,N_2357,N_4310);
nand U5781 (N_5781,N_2933,N_2909);
or U5782 (N_5782,N_3155,N_308);
xnor U5783 (N_5783,N_390,N_2653);
nand U5784 (N_5784,N_4296,N_3162);
or U5785 (N_5785,N_913,N_959);
and U5786 (N_5786,N_310,N_996);
or U5787 (N_5787,N_2641,N_3921);
or U5788 (N_5788,N_912,N_1295);
nand U5789 (N_5789,N_4795,N_4759);
or U5790 (N_5790,N_3838,N_733);
or U5791 (N_5791,N_4155,N_671);
nand U5792 (N_5792,N_1713,N_4737);
and U5793 (N_5793,N_3399,N_538);
or U5794 (N_5794,N_328,N_343);
nand U5795 (N_5795,N_465,N_4008);
and U5796 (N_5796,N_3135,N_3737);
or U5797 (N_5797,N_1818,N_3513);
or U5798 (N_5798,N_1432,N_3649);
and U5799 (N_5799,N_4247,N_336);
nor U5800 (N_5800,N_3545,N_3689);
or U5801 (N_5801,N_3509,N_2131);
and U5802 (N_5802,N_2654,N_384);
or U5803 (N_5803,N_4814,N_4537);
or U5804 (N_5804,N_3732,N_3241);
and U5805 (N_5805,N_4396,N_2130);
or U5806 (N_5806,N_284,N_4591);
or U5807 (N_5807,N_464,N_1338);
nor U5808 (N_5808,N_4291,N_4250);
nand U5809 (N_5809,N_1968,N_2353);
nand U5810 (N_5810,N_4346,N_4691);
nand U5811 (N_5811,N_4020,N_4748);
nand U5812 (N_5812,N_4411,N_1961);
and U5813 (N_5813,N_4451,N_2774);
and U5814 (N_5814,N_3774,N_3153);
and U5815 (N_5815,N_2440,N_1597);
nor U5816 (N_5816,N_4190,N_4492);
nor U5817 (N_5817,N_1885,N_2948);
nor U5818 (N_5818,N_831,N_181);
nand U5819 (N_5819,N_3147,N_4624);
and U5820 (N_5820,N_816,N_2717);
nand U5821 (N_5821,N_4672,N_4473);
nand U5822 (N_5822,N_2912,N_1339);
nor U5823 (N_5823,N_449,N_3176);
nor U5824 (N_5824,N_2625,N_4364);
or U5825 (N_5825,N_53,N_559);
and U5826 (N_5826,N_1765,N_3856);
or U5827 (N_5827,N_4481,N_2141);
nor U5828 (N_5828,N_514,N_1189);
nand U5829 (N_5829,N_3188,N_137);
and U5830 (N_5830,N_1110,N_1048);
nand U5831 (N_5831,N_3658,N_3074);
and U5832 (N_5832,N_4584,N_2689);
nor U5833 (N_5833,N_3824,N_4751);
nor U5834 (N_5834,N_3263,N_541);
or U5835 (N_5835,N_4332,N_537);
or U5836 (N_5836,N_2611,N_1730);
and U5837 (N_5837,N_127,N_1314);
nand U5838 (N_5838,N_2787,N_4277);
nand U5839 (N_5839,N_955,N_2072);
or U5840 (N_5840,N_3385,N_325);
and U5841 (N_5841,N_2939,N_3229);
nand U5842 (N_5842,N_4893,N_3436);
or U5843 (N_5843,N_2221,N_1608);
nand U5844 (N_5844,N_1626,N_369);
or U5845 (N_5845,N_4007,N_348);
and U5846 (N_5846,N_147,N_784);
and U5847 (N_5847,N_4458,N_3765);
and U5848 (N_5848,N_2032,N_1485);
nor U5849 (N_5849,N_1125,N_4568);
or U5850 (N_5850,N_650,N_1951);
or U5851 (N_5851,N_3111,N_4835);
nand U5852 (N_5852,N_1790,N_154);
nand U5853 (N_5853,N_3831,N_275);
or U5854 (N_5854,N_700,N_4441);
and U5855 (N_5855,N_2487,N_4145);
nand U5856 (N_5856,N_2170,N_2779);
or U5857 (N_5857,N_2932,N_2206);
nor U5858 (N_5858,N_1488,N_1505);
and U5859 (N_5859,N_565,N_3691);
or U5860 (N_5860,N_2129,N_4449);
nand U5861 (N_5861,N_2831,N_2308);
nor U5862 (N_5862,N_1870,N_18);
nor U5863 (N_5863,N_2186,N_3731);
nor U5864 (N_5864,N_1335,N_4118);
nor U5865 (N_5865,N_1755,N_2048);
and U5866 (N_5866,N_1484,N_1370);
or U5867 (N_5867,N_2016,N_1075);
or U5868 (N_5868,N_973,N_2257);
or U5869 (N_5869,N_2734,N_4236);
or U5870 (N_5870,N_3228,N_3642);
and U5871 (N_5871,N_2973,N_3092);
xnor U5872 (N_5872,N_3057,N_2478);
nand U5873 (N_5873,N_3438,N_4979);
or U5874 (N_5874,N_4896,N_186);
and U5875 (N_5875,N_868,N_2503);
or U5876 (N_5876,N_966,N_782);
nor U5877 (N_5877,N_1875,N_3243);
or U5878 (N_5878,N_3900,N_4595);
nor U5879 (N_5879,N_503,N_4255);
nor U5880 (N_5880,N_2450,N_2468);
nand U5881 (N_5881,N_2627,N_2105);
or U5882 (N_5882,N_4788,N_3996);
nand U5883 (N_5883,N_3471,N_743);
and U5884 (N_5884,N_2847,N_4767);
nor U5885 (N_5885,N_4099,N_78);
xor U5886 (N_5886,N_1082,N_713);
and U5887 (N_5887,N_3844,N_2333);
or U5888 (N_5888,N_309,N_1320);
and U5889 (N_5889,N_3065,N_4305);
and U5890 (N_5890,N_4453,N_2521);
or U5891 (N_5891,N_396,N_2080);
nand U5892 (N_5892,N_2915,N_4235);
and U5893 (N_5893,N_1152,N_933);
nor U5894 (N_5894,N_2078,N_2012);
nand U5895 (N_5895,N_2715,N_4116);
nor U5896 (N_5896,N_3312,N_1577);
and U5897 (N_5897,N_4245,N_1478);
nand U5898 (N_5898,N_1704,N_1065);
nand U5899 (N_5899,N_1215,N_4304);
nand U5900 (N_5900,N_2385,N_178);
nor U5901 (N_5901,N_3108,N_2349);
nor U5902 (N_5902,N_4798,N_2676);
and U5903 (N_5903,N_4229,N_2020);
or U5904 (N_5904,N_3656,N_852);
or U5905 (N_5905,N_941,N_4484);
nand U5906 (N_5906,N_3277,N_4024);
nand U5907 (N_5907,N_3439,N_975);
or U5908 (N_5908,N_2551,N_839);
nor U5909 (N_5909,N_904,N_2533);
nor U5910 (N_5910,N_1307,N_2828);
nor U5911 (N_5911,N_1613,N_262);
or U5912 (N_5912,N_1986,N_223);
nand U5913 (N_5913,N_4060,N_4183);
nand U5914 (N_5914,N_222,N_3516);
or U5915 (N_5915,N_1584,N_692);
nor U5916 (N_5916,N_2504,N_948);
and U5917 (N_5917,N_1673,N_4956);
nand U5918 (N_5918,N_1585,N_318);
or U5919 (N_5919,N_1443,N_3310);
and U5920 (N_5920,N_3531,N_1078);
or U5921 (N_5921,N_1700,N_2633);
nor U5922 (N_5922,N_2302,N_4384);
or U5923 (N_5923,N_4054,N_3826);
or U5924 (N_5924,N_341,N_3259);
and U5925 (N_5925,N_148,N_4406);
and U5926 (N_5926,N_4830,N_1297);
nor U5927 (N_5927,N_307,N_3340);
or U5928 (N_5928,N_2174,N_90);
and U5929 (N_5929,N_4207,N_2411);
or U5930 (N_5930,N_1960,N_1973);
nor U5931 (N_5931,N_1162,N_4391);
or U5932 (N_5932,N_2008,N_873);
nor U5933 (N_5933,N_4884,N_1573);
nand U5934 (N_5934,N_2420,N_1035);
nand U5935 (N_5935,N_2419,N_1849);
nor U5936 (N_5936,N_2796,N_3594);
and U5937 (N_5937,N_2876,N_4577);
nor U5938 (N_5938,N_2376,N_1919);
nand U5939 (N_5939,N_3448,N_226);
or U5940 (N_5940,N_214,N_820);
or U5941 (N_5941,N_4610,N_2516);
or U5942 (N_5942,N_4536,N_4580);
nor U5943 (N_5943,N_2690,N_1103);
nor U5944 (N_5944,N_1123,N_2532);
or U5945 (N_5945,N_3494,N_4828);
and U5946 (N_5946,N_190,N_2239);
or U5947 (N_5947,N_3628,N_2476);
nand U5948 (N_5948,N_1461,N_1436);
nand U5949 (N_5949,N_1169,N_3572);
nor U5950 (N_5950,N_2047,N_810);
or U5951 (N_5951,N_3784,N_1736);
nand U5952 (N_5952,N_1992,N_3182);
or U5953 (N_5953,N_3706,N_2518);
nor U5954 (N_5954,N_1464,N_321);
nor U5955 (N_5955,N_1910,N_1801);
and U5956 (N_5956,N_1598,N_4914);
or U5957 (N_5957,N_3888,N_898);
nand U5958 (N_5958,N_909,N_4435);
and U5959 (N_5959,N_4331,N_2610);
nand U5960 (N_5960,N_2571,N_1260);
nor U5961 (N_5961,N_227,N_3938);
xnor U5962 (N_5962,N_4769,N_194);
nor U5963 (N_5963,N_3514,N_301);
and U5964 (N_5964,N_3569,N_2208);
or U5965 (N_5965,N_4234,N_583);
or U5966 (N_5966,N_2931,N_350);
or U5967 (N_5967,N_3268,N_391);
and U5968 (N_5968,N_4005,N_3204);
nand U5969 (N_5969,N_3381,N_932);
or U5970 (N_5970,N_1367,N_3526);
nand U5971 (N_5971,N_3482,N_3720);
nor U5972 (N_5972,N_1745,N_4076);
or U5973 (N_5973,N_2891,N_217);
and U5974 (N_5974,N_4923,N_3136);
nor U5975 (N_5975,N_4124,N_3291);
nor U5976 (N_5976,N_2275,N_2572);
nor U5977 (N_5977,N_2956,N_4590);
nand U5978 (N_5978,N_877,N_1516);
nor U5979 (N_5979,N_2809,N_1551);
and U5980 (N_5980,N_2998,N_523);
nand U5981 (N_5981,N_2443,N_4280);
or U5982 (N_5982,N_429,N_3875);
nor U5983 (N_5983,N_4462,N_4539);
nor U5984 (N_5984,N_3529,N_4698);
nand U5985 (N_5985,N_2365,N_1258);
nor U5986 (N_5986,N_579,N_648);
and U5987 (N_5987,N_3506,N_4745);
nand U5988 (N_5988,N_283,N_475);
nor U5989 (N_5989,N_1095,N_2024);
nor U5990 (N_5990,N_4329,N_3461);
and U5991 (N_5991,N_4486,N_1840);
nor U5992 (N_5992,N_2166,N_3089);
nand U5993 (N_5993,N_172,N_742);
nor U5994 (N_5994,N_66,N_2117);
or U5995 (N_5995,N_1946,N_1721);
or U5996 (N_5996,N_1117,N_1293);
nor U5997 (N_5997,N_3641,N_2339);
nand U5998 (N_5998,N_1099,N_3817);
nand U5999 (N_5999,N_2455,N_3862);
and U6000 (N_6000,N_2165,N_806);
and U6001 (N_6001,N_2234,N_3006);
nor U6002 (N_6002,N_553,N_4011);
or U6003 (N_6003,N_2544,N_2505);
nand U6004 (N_6004,N_2775,N_759);
and U6005 (N_6005,N_68,N_1023);
nand U6006 (N_6006,N_1273,N_196);
nand U6007 (N_6007,N_1936,N_1328);
and U6008 (N_6008,N_646,N_4929);
and U6009 (N_6009,N_1867,N_2622);
or U6010 (N_6010,N_1017,N_701);
nor U6011 (N_6011,N_4284,N_2366);
or U6012 (N_6012,N_2602,N_1587);
nand U6013 (N_6013,N_4825,N_3614);
and U6014 (N_6014,N_1388,N_2877);
and U6015 (N_6015,N_3528,N_1681);
nand U6016 (N_6016,N_74,N_612);
or U6017 (N_6017,N_3157,N_2776);
and U6018 (N_6018,N_760,N_1319);
nand U6019 (N_6019,N_3286,N_3714);
nand U6020 (N_6020,N_2934,N_1423);
or U6021 (N_6021,N_2900,N_1166);
or U6022 (N_6022,N_2338,N_1440);
and U6023 (N_6023,N_4027,N_3038);
and U6024 (N_6024,N_3716,N_2483);
or U6025 (N_6025,N_118,N_3893);
or U6026 (N_6026,N_4049,N_218);
or U6027 (N_6027,N_1562,N_3446);
and U6028 (N_6028,N_3815,N_2416);
nand U6029 (N_6029,N_4407,N_2158);
and U6030 (N_6030,N_4834,N_1547);
or U6031 (N_6031,N_2465,N_961);
and U6032 (N_6032,N_4381,N_4715);
nand U6033 (N_6033,N_3549,N_1114);
nand U6034 (N_6034,N_3137,N_4656);
nand U6035 (N_6035,N_3255,N_4604);
nand U6036 (N_6036,N_4874,N_9);
and U6037 (N_6037,N_684,N_635);
nand U6038 (N_6038,N_4430,N_872);
and U6039 (N_6039,N_160,N_1416);
and U6040 (N_6040,N_1750,N_2549);
and U6041 (N_6041,N_2609,N_2512);
nor U6042 (N_6042,N_3507,N_2995);
nor U6043 (N_6043,N_4120,N_287);
nor U6044 (N_6044,N_4960,N_3945);
or U6045 (N_6045,N_2522,N_2848);
or U6046 (N_6046,N_3022,N_1942);
nor U6047 (N_6047,N_4818,N_3254);
and U6048 (N_6048,N_1637,N_1714);
nand U6049 (N_6049,N_3285,N_1275);
nand U6050 (N_6050,N_2022,N_2890);
or U6051 (N_6051,N_1285,N_1920);
and U6052 (N_6052,N_2112,N_4454);
nand U6053 (N_6053,N_4613,N_976);
nor U6054 (N_6054,N_461,N_2813);
and U6055 (N_6055,N_2590,N_3523);
nand U6056 (N_6056,N_4042,N_169);
or U6057 (N_6057,N_15,N_3786);
and U6058 (N_6058,N_132,N_2726);
and U6059 (N_6059,N_2228,N_1900);
nand U6060 (N_6060,N_3790,N_4211);
and U6061 (N_6061,N_3868,N_2628);
and U6062 (N_6062,N_91,N_2757);
or U6063 (N_6063,N_699,N_4797);
or U6064 (N_6064,N_2396,N_1426);
nand U6065 (N_6065,N_3375,N_2992);
or U6066 (N_6066,N_587,N_1878);
or U6067 (N_6067,N_2126,N_3665);
nand U6068 (N_6068,N_4817,N_1540);
and U6069 (N_6069,N_4002,N_1024);
or U6070 (N_6070,N_2352,N_1371);
nand U6071 (N_6071,N_1890,N_3379);
and U6072 (N_6072,N_1558,N_2296);
or U6073 (N_6073,N_2088,N_4003);
or U6074 (N_6074,N_4778,N_4982);
nor U6075 (N_6075,N_2433,N_4809);
or U6076 (N_6076,N_1682,N_2025);
or U6077 (N_6077,N_755,N_4948);
and U6078 (N_6078,N_3289,N_3735);
nand U6079 (N_6079,N_1866,N_2670);
nand U6080 (N_6080,N_878,N_4955);
nor U6081 (N_6081,N_1487,N_1536);
nand U6082 (N_6082,N_765,N_3601);
nor U6083 (N_6083,N_3905,N_1586);
or U6084 (N_6084,N_1654,N_155);
nand U6085 (N_6085,N_3979,N_1513);
or U6086 (N_6086,N_1442,N_1985);
or U6087 (N_6087,N_4530,N_4303);
nor U6088 (N_6088,N_3567,N_1733);
xor U6089 (N_6089,N_3416,N_366);
nor U6090 (N_6090,N_3804,N_731);
nor U6091 (N_6091,N_2922,N_71);
or U6092 (N_6092,N_63,N_1434);
nand U6093 (N_6093,N_3239,N_2751);
or U6094 (N_6094,N_1724,N_4976);
nand U6095 (N_6095,N_1846,N_2140);
nand U6096 (N_6096,N_2466,N_4498);
or U6097 (N_6097,N_3717,N_952);
and U6098 (N_6098,N_4442,N_1041);
nor U6099 (N_6099,N_1428,N_2271);
and U6100 (N_6100,N_1928,N_3290);
and U6101 (N_6101,N_2927,N_1063);
nor U6102 (N_6102,N_4695,N_2687);
nand U6103 (N_6103,N_3849,N_2883);
or U6104 (N_6104,N_3744,N_3552);
or U6105 (N_6105,N_3023,N_4163);
nand U6106 (N_6106,N_297,N_3639);
xnor U6107 (N_6107,N_4106,N_3978);
nand U6108 (N_6108,N_1619,N_1398);
and U6109 (N_6109,N_1349,N_1776);
and U6110 (N_6110,N_4967,N_2781);
or U6111 (N_6111,N_3327,N_3730);
or U6112 (N_6112,N_2782,N_3525);
or U6113 (N_6113,N_2942,N_2838);
and U6114 (N_6114,N_3095,N_4673);
nand U6115 (N_6115,N_3668,N_2119);
and U6116 (N_6116,N_4947,N_3318);
nand U6117 (N_6117,N_3170,N_3363);
nand U6118 (N_6118,N_3694,N_4704);
nand U6119 (N_6119,N_4333,N_4636);
nand U6120 (N_6120,N_450,N_99);
nand U6121 (N_6121,N_516,N_950);
nor U6122 (N_6122,N_2491,N_2861);
nand U6123 (N_6123,N_2168,N_861);
nand U6124 (N_6124,N_4783,N_4801);
or U6125 (N_6125,N_4360,N_3052);
and U6126 (N_6126,N_855,N_3284);
nor U6127 (N_6127,N_4348,N_3836);
nand U6128 (N_6128,N_0,N_4342);
nand U6129 (N_6129,N_3568,N_238);
nand U6130 (N_6130,N_4619,N_2050);
or U6131 (N_6131,N_577,N_4093);
or U6132 (N_6132,N_4085,N_1179);
nand U6133 (N_6133,N_3907,N_65);
nor U6134 (N_6134,N_3622,N_947);
nor U6135 (N_6135,N_278,N_4523);
nor U6136 (N_6136,N_1496,N_2508);
nand U6137 (N_6137,N_4764,N_1591);
nand U6138 (N_6138,N_763,N_4036);
or U6139 (N_6139,N_1380,N_4732);
nor U6140 (N_6140,N_776,N_1645);
nand U6141 (N_6141,N_2370,N_4641);
and U6142 (N_6142,N_4176,N_3078);
nand U6143 (N_6143,N_1408,N_403);
and U6144 (N_6144,N_1956,N_3821);
and U6145 (N_6145,N_3663,N_3357);
nor U6146 (N_6146,N_4507,N_80);
nand U6147 (N_6147,N_4048,N_2684);
nand U6148 (N_6148,N_1264,N_3314);
or U6149 (N_6149,N_1905,N_3501);
nand U6150 (N_6150,N_695,N_1663);
nand U6151 (N_6151,N_2380,N_4141);
and U6152 (N_6152,N_1383,N_3828);
or U6153 (N_6153,N_2246,N_4753);
nand U6154 (N_6154,N_881,N_3088);
nand U6155 (N_6155,N_2100,N_3292);
and U6156 (N_6156,N_655,N_3127);
or U6157 (N_6157,N_428,N_2747);
nand U6158 (N_6158,N_1749,N_4294);
and U6159 (N_6159,N_130,N_2299);
or U6160 (N_6160,N_1697,N_3899);
nand U6161 (N_6161,N_243,N_1916);
and U6162 (N_6162,N_2258,N_1805);
nand U6163 (N_6163,N_4545,N_3344);
nor U6164 (N_6164,N_992,N_191);
nor U6165 (N_6165,N_4162,N_2136);
nand U6166 (N_6166,N_4655,N_3874);
nand U6167 (N_6167,N_2675,N_3222);
nand U6168 (N_6168,N_2607,N_203);
and U6169 (N_6169,N_4461,N_2691);
and U6170 (N_6170,N_2542,N_2837);
or U6171 (N_6171,N_422,N_4035);
and U6172 (N_6172,N_2285,N_2659);
nand U6173 (N_6173,N_2301,N_1101);
nor U6174 (N_6174,N_3948,N_16);
or U6175 (N_6175,N_151,N_4637);
nor U6176 (N_6176,N_2382,N_829);
nor U6177 (N_6177,N_1988,N_892);
nand U6178 (N_6178,N_430,N_106);
or U6179 (N_6179,N_4227,N_1441);
and U6180 (N_6180,N_3846,N_251);
or U6181 (N_6181,N_4647,N_3336);
nand U6182 (N_6182,N_2372,N_3719);
and U6183 (N_6183,N_3178,N_1549);
nand U6184 (N_6184,N_1489,N_4200);
or U6185 (N_6185,N_3734,N_4389);
nor U6186 (N_6186,N_1400,N_1393);
nor U6187 (N_6187,N_4562,N_4557);
nor U6188 (N_6188,N_2212,N_4529);
and U6189 (N_6189,N_498,N_1225);
and U6190 (N_6190,N_4105,N_3861);
and U6191 (N_6191,N_3311,N_95);
or U6192 (N_6192,N_2092,N_3657);
nor U6193 (N_6193,N_3593,N_3799);
nor U6194 (N_6194,N_4052,N_3903);
nand U6195 (N_6195,N_2003,N_680);
nand U6196 (N_6196,N_1732,N_2736);
nand U6197 (N_6197,N_2069,N_1292);
or U6198 (N_6198,N_3237,N_2748);
nor U6199 (N_6199,N_995,N_1948);
or U6200 (N_6200,N_3225,N_1661);
and U6201 (N_6201,N_4090,N_3887);
nor U6202 (N_6202,N_2438,N_2679);
or U6203 (N_6203,N_156,N_4171);
nand U6204 (N_6204,N_3353,N_1002);
and U6205 (N_6205,N_4127,N_1798);
nand U6206 (N_6206,N_77,N_1854);
or U6207 (N_6207,N_1122,N_1576);
and U6208 (N_6208,N_1834,N_2295);
and U6209 (N_6209,N_259,N_4077);
or U6210 (N_6210,N_3217,N_3624);
and U6211 (N_6211,N_3771,N_2535);
or U6212 (N_6212,N_1550,N_2600);
and U6213 (N_6213,N_4944,N_1475);
nand U6214 (N_6214,N_3934,N_2983);
nor U6215 (N_6215,N_260,N_2446);
nand U6216 (N_6216,N_2178,N_2043);
nand U6217 (N_6217,N_563,N_927);
and U6218 (N_6218,N_3637,N_1411);
and U6219 (N_6219,N_3597,N_4839);
and U6220 (N_6220,N_2110,N_1829);
and U6221 (N_6221,N_1357,N_2052);
nand U6222 (N_6222,N_2226,N_2331);
or U6223 (N_6223,N_4394,N_2310);
nor U6224 (N_6224,N_104,N_1785);
and U6225 (N_6225,N_1257,N_285);
nor U6226 (N_6226,N_2971,N_1625);
nor U6227 (N_6227,N_660,N_1623);
nor U6228 (N_6228,N_2666,N_3367);
and U6229 (N_6229,N_2115,N_2336);
nor U6230 (N_6230,N_3351,N_494);
nor U6231 (N_6231,N_1361,N_2086);
and U6232 (N_6232,N_1181,N_2578);
nor U6233 (N_6233,N_2233,N_4662);
nor U6234 (N_6234,N_2986,N_4410);
and U6235 (N_6235,N_2509,N_2098);
nand U6236 (N_6236,N_4316,N_1511);
nor U6237 (N_6237,N_2926,N_3669);
nor U6238 (N_6238,N_525,N_2274);
nor U6239 (N_6239,N_3672,N_2978);
nand U6240 (N_6240,N_3588,N_2706);
nand U6241 (N_6241,N_647,N_1233);
nand U6242 (N_6242,N_3573,N_4295);
nor U6243 (N_6243,N_4399,N_2127);
nand U6244 (N_6244,N_3444,N_1280);
nor U6245 (N_6245,N_4862,N_4468);
nor U6246 (N_6246,N_3362,N_1844);
or U6247 (N_6247,N_1541,N_2694);
nand U6248 (N_6248,N_2108,N_2474);
nor U6249 (N_6249,N_72,N_1354);
nand U6250 (N_6250,N_1013,N_3242);
nand U6251 (N_6251,N_3647,N_4569);
and U6252 (N_6252,N_4040,N_1301);
nor U6253 (N_6253,N_59,N_4282);
and U6254 (N_6254,N_4134,N_2288);
and U6255 (N_6255,N_3740,N_2527);
nor U6256 (N_6256,N_4752,N_1228);
nand U6257 (N_6257,N_2488,N_4068);
and U6258 (N_6258,N_1342,N_3969);
nor U6259 (N_6259,N_3747,N_749);
nand U6260 (N_6260,N_2699,N_981);
nand U6261 (N_6261,N_250,N_2017);
nor U6262 (N_6262,N_3100,N_1810);
nand U6263 (N_6263,N_3380,N_2153);
nand U6264 (N_6264,N_1080,N_2002);
nor U6265 (N_6265,N_654,N_2225);
or U6266 (N_6266,N_4339,N_1529);
nand U6267 (N_6267,N_1716,N_1241);
nand U6268 (N_6268,N_2868,N_376);
nand U6269 (N_6269,N_4724,N_4532);
or U6270 (N_6270,N_1967,N_49);
or U6271 (N_6271,N_2732,N_1250);
nand U6272 (N_6272,N_2462,N_1901);
or U6273 (N_6273,N_379,N_1742);
nand U6274 (N_6274,N_4917,N_729);
nand U6275 (N_6275,N_1235,N_2437);
or U6276 (N_6276,N_2700,N_3424);
or U6277 (N_6277,N_3434,N_663);
and U6278 (N_6278,N_1145,N_1479);
nor U6279 (N_6279,N_1821,N_4117);
and U6280 (N_6280,N_1566,N_2562);
nand U6281 (N_6281,N_2,N_841);
nand U6282 (N_6282,N_3553,N_1472);
and U6283 (N_6283,N_1588,N_4761);
nand U6284 (N_6284,N_2444,N_597);
and U6285 (N_6285,N_3316,N_2742);
and U6286 (N_6286,N_4997,N_1675);
nor U6287 (N_6287,N_4535,N_2763);
and U6288 (N_6288,N_4671,N_3071);
or U6289 (N_6289,N_3556,N_4632);
or U6290 (N_6290,N_835,N_3402);
nor U6291 (N_6291,N_4816,N_1140);
nor U6292 (N_6292,N_4056,N_3179);
or U6293 (N_6293,N_117,N_2570);
nor U6294 (N_6294,N_2283,N_2616);
and U6295 (N_6295,N_529,N_3227);
or U6296 (N_6296,N_4209,N_2358);
xor U6297 (N_6297,N_879,N_4266);
or U6298 (N_6298,N_2403,N_2642);
nand U6299 (N_6299,N_2517,N_439);
nand U6300 (N_6300,N_2565,N_2878);
nand U6301 (N_6301,N_1688,N_1552);
nand U6302 (N_6302,N_833,N_1481);
nor U6303 (N_6303,N_2661,N_2200);
nand U6304 (N_6304,N_208,N_2070);
nor U6305 (N_6305,N_2250,N_1355);
or U6306 (N_6306,N_469,N_1788);
nor U6307 (N_6307,N_4021,N_2559);
or U6308 (N_6308,N_4602,N_2919);
or U6309 (N_6309,N_4623,N_1176);
or U6310 (N_6310,N_4444,N_4596);
nand U6311 (N_6311,N_2662,N_224);
nor U6312 (N_6312,N_4992,N_1781);
or U6313 (N_6313,N_32,N_3902);
nor U6314 (N_6314,N_1046,N_3443);
nand U6315 (N_6315,N_327,N_3081);
or U6316 (N_6316,N_1262,N_4963);
and U6317 (N_6317,N_1876,N_4683);
or U6318 (N_6318,N_3693,N_1221);
and U6319 (N_6319,N_566,N_4898);
nor U6320 (N_6320,N_4070,N_4793);
nand U6321 (N_6321,N_4345,N_723);
and U6322 (N_6322,N_1410,N_611);
nand U6323 (N_6323,N_694,N_2113);
nor U6324 (N_6324,N_2356,N_2749);
nor U6325 (N_6325,N_3368,N_1477);
and U6326 (N_6326,N_4693,N_4126);
nor U6327 (N_6327,N_2282,N_3244);
nor U6328 (N_6328,N_1226,N_273);
nor U6329 (N_6329,N_666,N_173);
and U6330 (N_6330,N_4903,N_3711);
nand U6331 (N_6331,N_4563,N_4739);
and U6332 (N_6332,N_499,N_230);
or U6333 (N_6333,N_2583,N_3388);
or U6334 (N_6334,N_4466,N_1051);
and U6335 (N_6335,N_637,N_4870);
nand U6336 (N_6336,N_4511,N_206);
nor U6337 (N_6337,N_3377,N_4423);
nor U6338 (N_6338,N_4485,N_2849);
or U6339 (N_6339,N_4242,N_1407);
or U6340 (N_6340,N_1517,N_3964);
and U6341 (N_6341,N_1807,N_4891);
and U6342 (N_6342,N_4925,N_2945);
nor U6343 (N_6343,N_3139,N_603);
and U6344 (N_6344,N_4743,N_3046);
or U6345 (N_6345,N_777,N_2494);
and U6346 (N_6346,N_1132,N_1515);
nand U6347 (N_6347,N_1802,N_1121);
nand U6348 (N_6348,N_4491,N_4412);
nand U6349 (N_6349,N_4990,N_4961);
nand U6350 (N_6350,N_3980,N_4571);
and U6351 (N_6351,N_1056,N_3018);
or U6352 (N_6352,N_974,N_589);
nand U6353 (N_6353,N_3201,N_1800);
nor U6354 (N_6354,N_4827,N_719);
and U6355 (N_6355,N_2730,N_4639);
xnor U6356 (N_6356,N_3317,N_3364);
or U6357 (N_6357,N_4206,N_4213);
nor U6358 (N_6358,N_2320,N_2300);
or U6359 (N_6359,N_2489,N_899);
nor U6360 (N_6360,N_3035,N_2966);
or U6361 (N_6361,N_306,N_2217);
nor U6362 (N_6362,N_3049,N_4528);
nor U6363 (N_6363,N_4625,N_3214);
nor U6364 (N_6364,N_3485,N_3648);
or U6365 (N_6365,N_462,N_1689);
and U6366 (N_6366,N_1826,N_2988);
nor U6367 (N_6367,N_1727,N_4551);
and U6368 (N_6368,N_2987,N_4476);
and U6369 (N_6369,N_64,N_1770);
or U6370 (N_6370,N_3358,N_1972);
nand U6371 (N_6371,N_4212,N_524);
and U6372 (N_6372,N_485,N_978);
or U6373 (N_6373,N_2681,N_149);
nor U6374 (N_6374,N_4810,N_2822);
nand U6375 (N_6375,N_4916,N_3294);
or U6376 (N_6376,N_3709,N_2415);
nand U6377 (N_6377,N_4347,N_3518);
nand U6378 (N_6378,N_2595,N_2180);
and U6379 (N_6379,N_4846,N_4824);
nor U6380 (N_6380,N_1420,N_4721);
and U6381 (N_6381,N_2795,N_4988);
nand U6382 (N_6382,N_3802,N_2272);
nor U6383 (N_6383,N_445,N_3288);
nand U6384 (N_6384,N_3930,N_3551);
nand U6385 (N_6385,N_31,N_2199);
nor U6386 (N_6386,N_3609,N_4413);
or U6387 (N_6387,N_1620,N_847);
nand U6388 (N_6388,N_4644,N_4680);
and U6389 (N_6389,N_4919,N_2536);
or U6390 (N_6390,N_139,N_304);
or U6391 (N_6391,N_1259,N_4738);
nand U6392 (N_6392,N_807,N_2401);
nand U6393 (N_6393,N_540,N_1076);
nor U6394 (N_6394,N_3174,N_4083);
nor U6395 (N_6395,N_532,N_4634);
nand U6396 (N_6396,N_4288,N_4701);
and U6397 (N_6397,N_4268,N_931);
nor U6398 (N_6398,N_1091,N_4397);
or U6399 (N_6399,N_1752,N_4257);
nor U6400 (N_6400,N_1607,N_4019);
nor U6401 (N_6401,N_908,N_3909);
nand U6402 (N_6402,N_2485,N_4030);
nand U6403 (N_6403,N_1220,N_2196);
nand U6404 (N_6404,N_3072,N_2435);
nand U6405 (N_6405,N_270,N_1294);
and U6406 (N_6406,N_3401,N_1559);
nand U6407 (N_6407,N_1105,N_4252);
nand U6408 (N_6408,N_355,N_3906);
nor U6409 (N_6409,N_3425,N_3743);
nand U6410 (N_6410,N_3334,N_593);
nor U6411 (N_6411,N_1131,N_2741);
and U6412 (N_6412,N_2251,N_2179);
nand U6413 (N_6413,N_2817,N_3270);
or U6414 (N_6414,N_1811,N_279);
nor U6415 (N_6415,N_3918,N_3841);
nand U6416 (N_6416,N_3115,N_359);
or U6417 (N_6417,N_598,N_4729);
or U6418 (N_6418,N_573,N_4123);
or U6419 (N_6419,N_4432,N_3456);
nor U6420 (N_6420,N_3451,N_314);
nand U6421 (N_6421,N_86,N_4606);
or U6422 (N_6422,N_1010,N_2759);
nor U6423 (N_6423,N_1746,N_4615);
nor U6424 (N_6424,N_1033,N_4219);
or U6425 (N_6425,N_3635,N_689);
or U6426 (N_6426,N_3499,N_1922);
and U6427 (N_6427,N_4669,N_3848);
and U6428 (N_6428,N_4426,N_1696);
or U6429 (N_6429,N_4244,N_3012);
nand U6430 (N_6430,N_3252,N_4080);
or U6431 (N_6431,N_109,N_3341);
or U6432 (N_6432,N_240,N_2882);
or U6433 (N_6433,N_143,N_3922);
nand U6434 (N_6434,N_1618,N_1832);
nand U6435 (N_6435,N_4369,N_4026);
nand U6436 (N_6436,N_4418,N_3118);
or U6437 (N_6437,N_629,N_3502);
or U6438 (N_6438,N_2467,N_2648);
nand U6439 (N_6439,N_4986,N_2554);
nand U6440 (N_6440,N_1617,N_3374);
nand U6441 (N_6441,N_3045,N_4688);
nand U6442 (N_6442,N_2316,N_1493);
and U6443 (N_6443,N_1202,N_1526);
and U6444 (N_6444,N_3028,N_4503);
nand U6445 (N_6445,N_344,N_1568);
or U6446 (N_6446,N_3615,N_166);
nand U6447 (N_6447,N_4175,N_2067);
and U6448 (N_6448,N_3814,N_1977);
nor U6449 (N_6449,N_3612,N_1610);
or U6450 (N_6450,N_4549,N_1794);
and U6451 (N_6451,N_338,N_3031);
nor U6452 (N_6452,N_257,N_2101);
and U6453 (N_6453,N_986,N_1784);
nor U6454 (N_6454,N_3808,N_2898);
nand U6455 (N_6455,N_4405,N_2925);
or U6456 (N_6456,N_556,N_1188);
or U6457 (N_6457,N_4318,N_4012);
nand U6458 (N_6458,N_1447,N_4860);
and U6459 (N_6459,N_3247,N_2156);
nor U6460 (N_6460,N_4572,N_4953);
and U6461 (N_6461,N_3493,N_405);
nor U6462 (N_6462,N_1282,N_4504);
nand U6463 (N_6463,N_4821,N_1238);
nor U6464 (N_6464,N_2343,N_2116);
nand U6465 (N_6465,N_1269,N_2123);
nor U6466 (N_6466,N_1683,N_690);
nand U6467 (N_6467,N_4975,N_1290);
nor U6468 (N_6468,N_3923,N_1605);
and U6469 (N_6469,N_502,N_2121);
and U6470 (N_6470,N_856,N_3791);
and U6471 (N_6471,N_1474,N_1344);
and U6472 (N_6472,N_3190,N_1574);
and U6473 (N_6473,N_1161,N_168);
nand U6474 (N_6474,N_4819,N_1096);
or U6475 (N_6475,N_4962,N_2812);
and U6476 (N_6476,N_2089,N_2924);
and U6477 (N_6477,N_4723,N_1768);
nand U6478 (N_6478,N_1763,N_480);
and U6479 (N_6479,N_2068,N_4443);
or U6480 (N_6480,N_2907,N_4259);
and U6481 (N_6481,N_4386,N_2703);
nor U6482 (N_6482,N_785,N_1822);
and U6483 (N_6483,N_136,N_630);
nor U6484 (N_6484,N_120,N_4542);
nand U6485 (N_6485,N_1924,N_4765);
or U6486 (N_6486,N_4686,N_4460);
and U6487 (N_6487,N_1884,N_751);
or U6488 (N_6488,N_4184,N_103);
nor U6489 (N_6489,N_1299,N_1414);
nor U6490 (N_6490,N_2106,N_3515);
nor U6491 (N_6491,N_1168,N_382);
or U6492 (N_6492,N_4328,N_3165);
and U6493 (N_6493,N_834,N_983);
nor U6494 (N_6494,N_4246,N_4820);
nand U6495 (N_6495,N_1842,N_1671);
and U6496 (N_6496,N_639,N_1687);
or U6497 (N_6497,N_3411,N_2636);
nor U6498 (N_6498,N_234,N_3464);
and U6499 (N_6499,N_3652,N_4273);
nand U6500 (N_6500,N_3972,N_4004);
or U6501 (N_6501,N_3773,N_387);
or U6502 (N_6502,N_3779,N_4446);
or U6503 (N_6503,N_2154,N_2586);
and U6504 (N_6504,N_3912,N_2281);
nor U6505 (N_6505,N_632,N_560);
nor U6506 (N_6506,N_2202,N_4713);
or U6507 (N_6507,N_1545,N_2379);
or U6508 (N_6508,N_3491,N_1308);
nand U6509 (N_6509,N_4527,N_4202);
nor U6510 (N_6510,N_303,N_2725);
xnor U6511 (N_6511,N_1287,N_4940);
nand U6512 (N_6512,N_1333,N_3993);
nor U6513 (N_6513,N_4958,N_1284);
nor U6514 (N_6514,N_1302,N_1352);
and U6515 (N_6515,N_3205,N_3863);
nand U6516 (N_6516,N_3504,N_4977);
nand U6517 (N_6517,N_1823,N_636);
nand U6518 (N_6518,N_924,N_3253);
or U6519 (N_6519,N_3924,N_3797);
and U6520 (N_6520,N_3587,N_3837);
and U6521 (N_6521,N_4622,N_371);
or U6522 (N_6522,N_989,N_3851);
and U6523 (N_6523,N_4853,N_3819);
nand U6524 (N_6524,N_1005,N_2081);
and U6525 (N_6525,N_1981,N_3325);
or U6526 (N_6526,N_3973,N_3138);
and U6527 (N_6527,N_380,N_768);
nand U6528 (N_6528,N_1525,N_3792);
and U6529 (N_6529,N_1707,N_3236);
nor U6530 (N_6530,N_116,N_4657);
nor U6531 (N_6531,N_2710,N_1227);
and U6532 (N_6532,N_249,N_4371);
nor U6533 (N_6533,N_2238,N_2566);
nand U6534 (N_6534,N_3396,N_1141);
nand U6535 (N_6535,N_1710,N_555);
nand U6536 (N_6536,N_3110,N_4319);
nand U6537 (N_6537,N_1157,N_2720);
or U6538 (N_6538,N_3563,N_546);
and U6539 (N_6539,N_3429,N_3595);
or U6540 (N_6540,N_1386,N_1170);
nand U6541 (N_6541,N_3063,N_2469);
nand U6542 (N_6542,N_1453,N_4700);
xor U6543 (N_6543,N_3000,N_4263);
nor U6544 (N_6544,N_2769,N_4355);
nand U6545 (N_6545,N_3124,N_3427);
nand U6546 (N_6546,N_188,N_3674);
or U6547 (N_6547,N_2270,N_4028);
or U6548 (N_6548,N_296,N_417);
nor U6549 (N_6549,N_1245,N_1880);
nor U6550 (N_6550,N_1288,N_2430);
and U6551 (N_6551,N_2820,N_3163);
nor U6552 (N_6552,N_1921,N_3505);
nand U6553 (N_6553,N_4525,N_1653);
and U6554 (N_6554,N_1723,N_2311);
nand U6555 (N_6555,N_4158,N_3670);
nor U6556 (N_6556,N_4994,N_3106);
nand U6557 (N_6557,N_1457,N_3767);
nand U6558 (N_6558,N_3441,N_4667);
nor U6559 (N_6559,N_1237,N_1509);
nand U6560 (N_6560,N_3462,N_3695);
nand U6561 (N_6561,N_3864,N_4367);
nor U6562 (N_6562,N_258,N_3564);
or U6563 (N_6563,N_3194,N_2844);
nor U6564 (N_6564,N_4920,N_1979);
or U6565 (N_6565,N_3701,N_4959);
and U6566 (N_6566,N_1864,N_3014);
nor U6567 (N_6567,N_4351,N_1583);
nand U6568 (N_6568,N_825,N_4031);
nand U6569 (N_6569,N_1938,N_4522);
or U6570 (N_6570,N_3915,N_4016);
or U6571 (N_6571,N_1841,N_4401);
nand U6572 (N_6572,N_4072,N_383);
nand U6573 (N_6573,N_1753,N_1490);
nor U6574 (N_6574,N_4439,N_3834);
and U6575 (N_6575,N_1677,N_4314);
nand U6576 (N_6576,N_1055,N_2640);
nor U6577 (N_6577,N_3630,N_3646);
or U6578 (N_6578,N_615,N_2713);
or U6579 (N_6579,N_2899,N_2334);
and U6580 (N_6580,N_4517,N_661);
or U6581 (N_6581,N_1138,N_3976);
and U6582 (N_6582,N_3952,N_707);
or U6583 (N_6583,N_2946,N_2007);
and U6584 (N_6584,N_434,N_1198);
and U6585 (N_6585,N_1087,N_3408);
nor U6586 (N_6586,N_4189,N_3586);
nor U6587 (N_6587,N_1193,N_2786);
and U6588 (N_6588,N_3543,N_459);
and U6589 (N_6589,N_4910,N_3331);
nor U6590 (N_6590,N_3180,N_27);
and U6591 (N_6591,N_4588,N_2486);
nor U6592 (N_6592,N_4129,N_4195);
nor U6593 (N_6593,N_3415,N_1538);
or U6594 (N_6594,N_3956,N_476);
and U6595 (N_6595,N_215,N_3540);
nand U6596 (N_6596,N_401,N_2064);
and U6597 (N_6597,N_3387,N_2083);
nor U6598 (N_6598,N_3768,N_3053);
or U6599 (N_6599,N_10,N_3751);
nand U6600 (N_6600,N_1092,N_3231);
or U6601 (N_6601,N_1044,N_1433);
nor U6602 (N_6602,N_4238,N_897);
nor U6603 (N_6603,N_3409,N_2346);
or U6604 (N_6604,N_2897,N_317);
or U6605 (N_6605,N_1000,N_2543);
or U6606 (N_6606,N_4336,N_1444);
nand U6607 (N_6607,N_1247,N_2728);
nor U6608 (N_6608,N_187,N_3145);
nor U6609 (N_6609,N_320,N_1771);
and U6610 (N_6610,N_4941,N_4648);
and U6611 (N_6611,N_3760,N_1058);
or U6612 (N_6612,N_693,N_651);
or U6613 (N_6613,N_4931,N_3114);
nand U6614 (N_6614,N_3300,N_2548);
and U6615 (N_6615,N_4554,N_289);
nand U6616 (N_6616,N_3121,N_3026);
nand U6617 (N_6617,N_710,N_1306);
nor U6618 (N_6618,N_1686,N_4174);
nor U6619 (N_6619,N_4224,N_1803);
xnor U6620 (N_6620,N_946,N_706);
and U6621 (N_6621,N_4087,N_1859);
and U6622 (N_6622,N_4879,N_4560);
nand U6623 (N_6623,N_4781,N_4868);
nand U6624 (N_6624,N_377,N_110);
nand U6625 (N_6625,N_2719,N_4341);
nor U6626 (N_6626,N_1216,N_1313);
or U6627 (N_6627,N_463,N_122);
nor U6628 (N_6628,N_3954,N_791);
or U6629 (N_6629,N_1668,N_1570);
nor U6630 (N_6630,N_158,N_280);
nor U6631 (N_6631,N_4094,N_2598);
or U6632 (N_6632,N_1518,N_1061);
and U6633 (N_6633,N_3458,N_84);
and U6634 (N_6634,N_373,N_1819);
nor U6635 (N_6635,N_936,N_4194);
and U6636 (N_6636,N_2644,N_1084);
and U6637 (N_6637,N_1463,N_1185);
nor U6638 (N_6638,N_1449,N_2484);
nand U6639 (N_6639,N_85,N_4928);
and U6640 (N_6640,N_4603,N_2981);
and U6641 (N_6641,N_1912,N_3947);
or U6642 (N_6642,N_24,N_3891);
and U6643 (N_6643,N_1439,N_832);
or U6644 (N_6644,N_3098,N_3660);
or U6645 (N_6645,N_3313,N_607);
or U6646 (N_6646,N_1229,N_4168);
nor U6647 (N_6647,N_4974,N_1470);
and U6648 (N_6648,N_1210,N_4286);
or U6649 (N_6649,N_2976,N_3498);
or U6650 (N_6650,N_894,N_2109);
nand U6651 (N_6651,N_1838,N_3962);
or U6652 (N_6652,N_3030,N_1167);
nand U6653 (N_6653,N_67,N_3226);
and U6654 (N_6654,N_4196,N_1381);
nand U6655 (N_6655,N_2970,N_2114);
or U6656 (N_6656,N_1147,N_554);
nor U6657 (N_6657,N_3680,N_1883);
or U6658 (N_6658,N_1495,N_2391);
nand U6659 (N_6659,N_2908,N_2254);
nand U6660 (N_6660,N_2268,N_4178);
and U6661 (N_6661,N_2729,N_3576);
nand U6662 (N_6662,N_644,N_4499);
or U6663 (N_6663,N_4845,N_1669);
and U6664 (N_6664,N_3631,N_114);
or U6665 (N_6665,N_2727,N_119);
nor U6666 (N_6666,N_2481,N_3036);
or U6667 (N_6667,N_3304,N_4488);
and U6668 (N_6668,N_3335,N_638);
and U6669 (N_6669,N_3305,N_558);
nand U6670 (N_6670,N_859,N_2065);
and U6671 (N_6671,N_4323,N_1877);
or U6672 (N_6672,N_3733,N_945);
and U6673 (N_6673,N_2243,N_4133);
or U6674 (N_6674,N_3697,N_4857);
nand U6675 (N_6675,N_232,N_1336);
nand U6676 (N_6676,N_2426,N_4519);
nand U6677 (N_6677,N_4382,N_2936);
nor U6678 (N_6678,N_1064,N_4886);
and U6679 (N_6679,N_4149,N_474);
and U6680 (N_6680,N_490,N_3640);
and U6681 (N_6681,N_735,N_4248);
nand U6682 (N_6682,N_1917,N_3742);
xor U6683 (N_6683,N_2608,N_1999);
or U6684 (N_6684,N_1007,N_977);
nand U6685 (N_6685,N_994,N_2149);
and U6686 (N_6686,N_1957,N_3967);
and U6687 (N_6687,N_2829,N_48);
and U6688 (N_6688,N_3094,N_903);
nor U6689 (N_6689,N_4882,N_535);
nand U6690 (N_6690,N_3008,N_4146);
nor U6691 (N_6691,N_4600,N_4037);
nor U6692 (N_6692,N_386,N_370);
nor U6693 (N_6693,N_2953,N_3517);
or U6694 (N_6694,N_4904,N_3809);
or U6695 (N_6695,N_3736,N_481);
nor U6696 (N_6696,N_4290,N_2425);
nor U6697 (N_6697,N_3019,N_2846);
and U6698 (N_6698,N_4966,N_4293);
or U6699 (N_6699,N_4403,N_2557);
and U6700 (N_6700,N_3027,N_1624);
nand U6701 (N_6701,N_2175,N_161);
nor U6702 (N_6702,N_423,N_3621);
nand U6703 (N_6703,N_2362,N_288);
nand U6704 (N_6704,N_2107,N_3975);
or U6705 (N_6705,N_3873,N_3219);
nor U6706 (N_6706,N_460,N_1094);
nor U6707 (N_6707,N_2954,N_3339);
or U6708 (N_6708,N_1656,N_305);
nor U6709 (N_6709,N_4509,N_1740);
and U6710 (N_6710,N_1040,N_2460);
xnor U6711 (N_6711,N_254,N_2145);
or U6712 (N_6712,N_315,N_3577);
nand U6713 (N_6713,N_1028,N_1564);
nor U6714 (N_6714,N_4939,N_618);
nor U6715 (N_6715,N_3892,N_159);
or U6716 (N_6716,N_395,N_4876);
nand U6717 (N_6717,N_848,N_4552);
nand U6718 (N_6718,N_625,N_1599);
and U6719 (N_6719,N_3800,N_2479);
nand U6720 (N_6720,N_3308,N_1641);
nand U6721 (N_6721,N_3151,N_1869);
nand U6722 (N_6722,N_267,N_1427);
and U6723 (N_6723,N_2906,N_4192);
nor U6724 (N_6724,N_1376,N_2663);
nand U6725 (N_6725,N_3248,N_704);
and U6726 (N_6726,N_3870,N_649);
nand U6727 (N_6727,N_783,N_3355);
and U6728 (N_6728,N_4755,N_1419);
and U6729 (N_6729,N_1522,N_2384);
or U6730 (N_6730,N_4153,N_443);
and U6731 (N_6731,N_489,N_171);
or U6732 (N_6732,N_3904,N_2816);
and U6733 (N_6733,N_4969,N_3571);
nand U6734 (N_6734,N_407,N_1868);
and U6735 (N_6735,N_2555,N_4674);
and U6736 (N_6736,N_4177,N_2760);
or U6737 (N_6737,N_4902,N_4357);
and U6738 (N_6738,N_4685,N_830);
and U6739 (N_6739,N_4075,N_2991);
nor U6740 (N_6740,N_198,N_4773);
nor U6741 (N_6741,N_1706,N_3883);
or U6742 (N_6742,N_1201,N_4682);
or U6743 (N_6743,N_4330,N_3940);
nand U6744 (N_6744,N_3895,N_656);
and U6745 (N_6745,N_1431,N_4803);
nor U6746 (N_6746,N_4450,N_4911);
or U6747 (N_6747,N_3708,N_4524);
nor U6748 (N_6748,N_1404,N_3382);
nor U6749 (N_6749,N_4185,N_2756);
nor U6750 (N_6750,N_1665,N_4156);
and U6751 (N_6751,N_4515,N_3117);
and U6752 (N_6752,N_4452,N_3218);
nor U6753 (N_6753,N_4232,N_4358);
nor U6754 (N_6754,N_2855,N_3420);
nor U6755 (N_6755,N_3007,N_1503);
xnor U6756 (N_6756,N_1989,N_153);
nand U6757 (N_6757,N_1809,N_4471);
or U6758 (N_6758,N_4317,N_138);
and U6759 (N_6759,N_4278,N_4459);
nand U6760 (N_6760,N_1560,N_895);
nor U6761 (N_6761,N_242,N_874);
and U6762 (N_6762,N_1151,N_2265);
or U6763 (N_6763,N_1332,N_1456);
nor U6764 (N_6764,N_3230,N_1902);
nand U6765 (N_6765,N_2035,N_2597);
or U6766 (N_6766,N_4758,N_2857);
nand U6767 (N_6767,N_4157,N_1693);
and U6768 (N_6768,N_1115,N_687);
xor U6769 (N_6769,N_1865,N_4301);
xor U6770 (N_6770,N_2546,N_2417);
or U6771 (N_6771,N_2388,N_3537);
nand U6772 (N_6772,N_4326,N_4006);
or U6773 (N_6773,N_2039,N_4354);
nor U6774 (N_6774,N_4477,N_2303);
nand U6775 (N_6775,N_35,N_3245);
or U6776 (N_6776,N_1368,N_4170);
nand U6777 (N_6777,N_4385,N_2972);
nor U6778 (N_6778,N_2647,N_3581);
and U6779 (N_6779,N_1243,N_2930);
nor U6780 (N_6780,N_2556,N_1692);
and U6781 (N_6781,N_2545,N_1263);
or U6782 (N_6782,N_3723,N_70);
nor U6783 (N_6783,N_604,N_3076);
nand U6784 (N_6784,N_3890,N_4297);
and U6785 (N_6785,N_3476,N_605);
and U6786 (N_6786,N_2169,N_4379);
and U6787 (N_6787,N_3582,N_2309);
nand U6788 (N_6788,N_209,N_818);
or U6789 (N_6789,N_4356,N_3520);
nand U6790 (N_6790,N_1717,N_170);
or U6791 (N_6791,N_4508,N_1512);
nor U6792 (N_6792,N_1422,N_1476);
or U6793 (N_6793,N_4334,N_2665);
or U6794 (N_6794,N_896,N_4873);
nor U6795 (N_6795,N_1192,N_4697);
and U6796 (N_6796,N_2650,N_621);
and U6797 (N_6797,N_2821,N_302);
or U6798 (N_6798,N_3272,N_1642);
or U6799 (N_6799,N_2531,N_2197);
or U6800 (N_6800,N_4009,N_798);
nand U6801 (N_6801,N_1982,N_960);
nor U6802 (N_6802,N_3296,N_2738);
or U6803 (N_6803,N_3718,N_4400);
xor U6804 (N_6804,N_4786,N_3017);
or U6805 (N_6805,N_2962,N_3393);
nand U6806 (N_6806,N_794,N_46);
or U6807 (N_6807,N_1403,N_1532);
or U6808 (N_6808,N_4017,N_2249);
nand U6809 (N_6809,N_1708,N_567);
nor U6810 (N_6810,N_4388,N_4650);
or U6811 (N_6811,N_971,N_105);
or U6812 (N_6812,N_4131,N_3778);
nor U6813 (N_6813,N_901,N_890);
or U6814 (N_6814,N_590,N_3713);
nor U6815 (N_6815,N_294,N_272);
or U6816 (N_6816,N_1596,N_2584);
nor U6817 (N_6817,N_2227,N_750);
or U6818 (N_6818,N_1557,N_2635);
or U6819 (N_6819,N_3354,N_1271);
or U6820 (N_6820,N_3997,N_3445);
and U6821 (N_6821,N_165,N_3788);
nor U6822 (N_6822,N_938,N_36);
and U6823 (N_6823,N_1643,N_4160);
or U6824 (N_6824,N_4437,N_60);
and U6825 (N_6825,N_1553,N_580);
nand U6826 (N_6826,N_2752,N_3184);
nand U6827 (N_6827,N_20,N_4148);
nand U6828 (N_6828,N_1998,N_3468);
and U6829 (N_6829,N_1113,N_2229);
and U6830 (N_6830,N_4970,N_802);
nand U6831 (N_6831,N_2951,N_907);
nand U6832 (N_6832,N_1514,N_448);
or U6833 (N_6833,N_2161,N_3373);
nor U6834 (N_6834,N_2377,N_3698);
and U6835 (N_6835,N_2788,N_1363);
nand U6836 (N_6836,N_942,N_1153);
and U6837 (N_6837,N_1219,N_3676);
nand U6838 (N_6838,N_3044,N_2693);
nand U6839 (N_6839,N_738,N_1659);
and U6840 (N_6840,N_1020,N_4233);
nand U6841 (N_6841,N_3798,N_3724);
and U6842 (N_6842,N_3463,N_3086);
or U6843 (N_6843,N_388,N_1102);
or U6844 (N_6844,N_2863,N_365);
nand U6845 (N_6845,N_709,N_1614);
nand U6846 (N_6846,N_3643,N_4844);
and U6847 (N_6847,N_241,N_346);
and U6848 (N_6848,N_530,N_61);
nor U6849 (N_6849,N_1079,N_550);
or U6850 (N_6850,N_3221,N_2780);
nor U6851 (N_6851,N_4775,N_4694);
and U6852 (N_6852,N_3832,N_3287);
nand U6853 (N_6853,N_4807,N_3696);
nor U6854 (N_6854,N_3453,N_3175);
nor U6855 (N_6855,N_3328,N_2833);
and U6856 (N_6856,N_4436,N_1783);
nand U6857 (N_6857,N_2879,N_94);
nor U6858 (N_6858,N_1945,N_1676);
and U6859 (N_6859,N_4309,N_1291);
and U6860 (N_6860,N_3246,N_2241);
and U6861 (N_6861,N_557,N_698);
nand U6862 (N_6862,N_1248,N_2623);
nand U6863 (N_6863,N_937,N_349);
nor U6864 (N_6864,N_4187,N_906);
or U6865 (N_6865,N_2686,N_2799);
nor U6866 (N_6866,N_1037,N_2449);
xor U6867 (N_6867,N_708,N_1072);
nand U6868 (N_6868,N_3039,N_4567);
and U6869 (N_6869,N_2128,N_3488);
or U6870 (N_6870,N_526,N_789);
and U6871 (N_6871,N_922,N_4115);
nor U6872 (N_6872,N_1899,N_3394);
and U6873 (N_6873,N_2513,N_2682);
and U6874 (N_6874,N_2222,N_2463);
or U6875 (N_6875,N_4805,N_705);
or U6876 (N_6876,N_889,N_951);
nor U6877 (N_6877,N_1326,N_2220);
and U6878 (N_6878,N_4841,N_2232);
nand U6879 (N_6879,N_3384,N_1555);
and U6880 (N_6880,N_1217,N_1646);
or U6881 (N_6881,N_3598,N_4740);
and U6882 (N_6882,N_2082,N_3234);
nor U6883 (N_6883,N_293,N_2248);
nand U6884 (N_6884,N_1699,N_89);
nor U6885 (N_6885,N_211,N_1658);
nand U6886 (N_6886,N_4320,N_3782);
nor U6887 (N_6887,N_4608,N_3125);
or U6888 (N_6888,N_389,N_1309);
nand U6889 (N_6889,N_4806,N_4804);
nor U6890 (N_6890,N_2869,N_2074);
or U6891 (N_6891,N_295,N_4267);
nor U6892 (N_6892,N_762,N_269);
or U6893 (N_6893,N_1554,N_3349);
nor U6894 (N_6894,N_1974,N_586);
or U6895 (N_6895,N_1858,N_910);
and U6896 (N_6896,N_4506,N_1744);
and U6897 (N_6897,N_152,N_3910);
nand U6898 (N_6898,N_3140,N_3128);
and U6899 (N_6899,N_4395,N_3413);
nor U6900 (N_6900,N_4378,N_12);
and U6901 (N_6901,N_231,N_1777);
or U6902 (N_6902,N_4699,N_4487);
and U6903 (N_6903,N_324,N_4497);
and U6904 (N_6904,N_3149,N_2290);
nor U6905 (N_6905,N_2534,N_1458);
nor U6906 (N_6906,N_3397,N_1672);
nand U6907 (N_6907,N_2292,N_3352);
nor U6908 (N_6908,N_1774,N_4899);
or U6909 (N_6909,N_2259,N_4642);
nand U6910 (N_6910,N_1690,N_4494);
or U6911 (N_6911,N_4913,N_2498);
nor U6912 (N_6912,N_3345,N_1678);
or U6913 (N_6913,N_640,N_1004);
nand U6914 (N_6914,N_4279,N_1839);
nor U6915 (N_6915,N_394,N_2133);
nand U6916 (N_6916,N_2273,N_528);
and U6917 (N_6917,N_2019,N_3548);
or U6918 (N_6918,N_408,N_3040);
nand U6919 (N_6919,N_1019,N_1680);
nor U6920 (N_6920,N_4631,N_1507);
and U6921 (N_6921,N_4039,N_466);
nand U6922 (N_6922,N_2011,N_4668);
or U6923 (N_6923,N_3684,N_3623);
nor U6924 (N_6924,N_1086,N_1032);
and U6925 (N_6925,N_718,N_758);
or U6926 (N_6926,N_2723,N_2143);
and U6927 (N_6927,N_4404,N_628);
and U6928 (N_6928,N_4228,N_4652);
or U6929 (N_6929,N_3223,N_179);
nand U6930 (N_6930,N_180,N_2335);
or U6931 (N_6931,N_2210,N_1156);
xnor U6932 (N_6932,N_3003,N_1737);
and U6933 (N_6933,N_1940,N_1994);
nor U6934 (N_6934,N_4847,N_4029);
nand U6935 (N_6935,N_2063,N_3677);
or U6936 (N_6936,N_1409,N_2804);
nand U6937 (N_6937,N_1205,N_4001);
and U6938 (N_6938,N_2172,N_4725);
or U6939 (N_6939,N_2242,N_3414);
nand U6940 (N_6940,N_3302,N_4119);
nand U6941 (N_6941,N_1343,N_2711);
nor U6942 (N_6942,N_4425,N_4514);
nand U6943 (N_6943,N_4390,N_799);
and U6944 (N_6944,N_3280,N_717);
and U6945 (N_6945,N_4010,N_3557);
nor U6946 (N_6946,N_3419,N_1501);
or U6947 (N_6947,N_1390,N_2245);
nor U6948 (N_6948,N_424,N_1861);
or U6949 (N_6949,N_3544,N_1042);
nor U6950 (N_6950,N_1276,N_686);
and U6951 (N_6951,N_2903,N_1604);
nand U6952 (N_6952,N_2692,N_3971);
nor U6953 (N_6953,N_2472,N_3282);
or U6954 (N_6954,N_357,N_821);
and U6955 (N_6955,N_1820,N_1914);
or U6956 (N_6956,N_406,N_1137);
nand U6957 (N_6957,N_3721,N_4883);
and U6958 (N_6958,N_3839,N_3645);
and U6959 (N_6959,N_4311,N_2252);
nand U6960 (N_6960,N_3465,N_444);
and U6961 (N_6961,N_4210,N_1021);
or U6962 (N_6962,N_4260,N_4045);
nand U6963 (N_6963,N_4064,N_4935);
nor U6964 (N_6964,N_1174,N_212);
and U6965 (N_6965,N_1178,N_1469);
and U6966 (N_6966,N_3787,N_4555);
or U6967 (N_6967,N_1871,N_2638);
nand U6968 (N_6968,N_1931,N_4972);
or U6969 (N_6969,N_3726,N_2350);
nand U6970 (N_6970,N_3591,N_4802);
or U6971 (N_6971,N_3610,N_1963);
nor U6972 (N_6972,N_3522,N_2314);
nand U6973 (N_6973,N_4518,N_438);
nand U6974 (N_6974,N_204,N_4455);
and U6975 (N_6975,N_3087,N_4122);
nand U6976 (N_6976,N_3495,N_2501);
nand U6977 (N_6977,N_4744,N_2800);
nand U6978 (N_6978,N_1567,N_780);
nor U6979 (N_6979,N_3181,N_1047);
nand U6980 (N_6980,N_4074,N_2442);
nor U6981 (N_6981,N_26,N_3813);
nand U6982 (N_6982,N_808,N_4837);
or U6983 (N_6983,N_4363,N_495);
and U6984 (N_6984,N_1633,N_4256);
nor U6985 (N_6985,N_4937,N_3447);
nor U6986 (N_6986,N_57,N_1159);
nor U6987 (N_6987,N_2013,N_4361);
and U6988 (N_6988,N_3209,N_997);
or U6989 (N_6989,N_4601,N_3455);
nor U6990 (N_6990,N_4556,N_2014);
nand U6991 (N_6991,N_4046,N_4414);
nand U6992 (N_6992,N_2287,N_3193);
nand U6993 (N_6993,N_2321,N_2896);
nor U6994 (N_6994,N_2913,N_3850);
nand U6995 (N_6995,N_1969,N_1726);
nor U6996 (N_6996,N_902,N_4589);
and U6997 (N_6997,N_1329,N_4221);
or U6998 (N_6998,N_1738,N_3690);
nor U6999 (N_6999,N_4302,N_3004);
nor U7000 (N_7000,N_1356,N_1909);
nand U7001 (N_7001,N_3533,N_4984);
or U7002 (N_7002,N_2735,N_871);
nor U7003 (N_7003,N_2317,N_4599);
and U7004 (N_7004,N_4651,N_1330);
nand U7005 (N_7005,N_4374,N_4611);
xor U7006 (N_7006,N_1792,N_893);
or U7007 (N_7007,N_2400,N_4678);
or U7008 (N_7008,N_773,N_2319);
nor U7009 (N_7009,N_697,N_1360);
or U7010 (N_7010,N_985,N_582);
nor U7011 (N_7011,N_1039,N_2261);
nand U7012 (N_7012,N_923,N_634);
nor U7013 (N_7013,N_471,N_505);
and U7014 (N_7014,N_2964,N_2368);
or U7015 (N_7015,N_4193,N_1950);
nand U7016 (N_7016,N_3925,N_347);
and U7017 (N_7017,N_3159,N_1029);
and U7018 (N_7018,N_3279,N_4370);
nand U7019 (N_7019,N_1366,N_2528);
nand U7020 (N_7020,N_4092,N_1881);
nand U7021 (N_7021,N_4777,N_1068);
nand U7022 (N_7022,N_3833,N_1889);
and U7023 (N_7023,N_3271,N_3048);
or U7024 (N_7024,N_2525,N_1394);
and U7025 (N_7025,N_4041,N_411);
and U7026 (N_7026,N_2696,N_3332);
nand U7027 (N_7027,N_2854,N_129);
nand U7028 (N_7028,N_616,N_4501);
nand U7029 (N_7029,N_4098,N_2510);
and U7030 (N_7030,N_4306,N_2646);
or U7031 (N_7031,N_228,N_2592);
nand U7032 (N_7032,N_617,N_1365);
nor U7033 (N_7033,N_2881,N_3168);
or U7034 (N_7034,N_100,N_239);
nor U7035 (N_7035,N_3070,N_229);
and U7036 (N_7036,N_3240,N_4559);
and U7037 (N_7037,N_3678,N_916);
and U7038 (N_7038,N_1793,N_4731);
and U7039 (N_7039,N_1937,N_271);
xnor U7040 (N_7040,N_124,N_1406);
and U7041 (N_7041,N_2888,N_1492);
nand U7042 (N_7042,N_506,N_4800);
nand U7043 (N_7043,N_1602,N_69);
nand U7044 (N_7044,N_496,N_4789);
or U7045 (N_7045,N_3966,N_609);
nand U7046 (N_7046,N_1799,N_2324);
nor U7047 (N_7047,N_184,N_2044);
and U7048 (N_7048,N_574,N_1600);
or U7049 (N_7049,N_3919,N_3759);
and U7050 (N_7050,N_2856,N_1506);
and U7051 (N_7051,N_316,N_2671);
nor U7052 (N_7052,N_3936,N_608);
nand U7053 (N_7053,N_2267,N_431);
nand U7054 (N_7054,N_3679,N_4307);
and U7055 (N_7055,N_4159,N_3683);
nand U7056 (N_7056,N_3852,N_1932);
or U7057 (N_7057,N_3911,N_14);
and U7058 (N_7058,N_1323,N_4880);
and U7059 (N_7059,N_1848,N_876);
nor U7060 (N_7060,N_575,N_965);
nand U7061 (N_7061,N_2604,N_3738);
or U7062 (N_7062,N_2835,N_1224);
and U7063 (N_7063,N_3644,N_775);
and U7064 (N_7064,N_1629,N_3407);
nand U7065 (N_7065,N_2389,N_3607);
and U7066 (N_7066,N_331,N_4957);
nor U7067 (N_7067,N_4463,N_1194);
and U7068 (N_7068,N_3202,N_3872);
nand U7069 (N_7069,N_2475,N_4365);
nor U7070 (N_7070,N_984,N_1739);
nor U7071 (N_7071,N_3484,N_4756);
nor U7072 (N_7072,N_3801,N_1650);
and U7073 (N_7073,N_1660,N_2923);
and U7074 (N_7074,N_3566,N_3418);
or U7075 (N_7075,N_4945,N_2840);
nor U7076 (N_7076,N_4646,N_652);
nand U7077 (N_7077,N_1534,N_233);
and U7078 (N_7078,N_1502,N_1430);
and U7079 (N_7079,N_4181,N_4220);
and U7080 (N_7080,N_4063,N_4161);
nor U7081 (N_7081,N_4843,N_1954);
nor U7082 (N_7082,N_182,N_286);
or U7083 (N_7083,N_3943,N_1350);
nor U7084 (N_7084,N_1234,N_4858);
nor U7085 (N_7085,N_3927,N_4434);
nand U7086 (N_7086,N_3896,N_2984);
and U7087 (N_7087,N_1897,N_2631);
xnor U7088 (N_7088,N_1628,N_4061);
or U7089 (N_7089,N_1069,N_4292);
and U7090 (N_7090,N_533,N_4692);
and U7091 (N_7091,N_3066,N_1892);
nand U7092 (N_7092,N_2867,N_220);
and U7093 (N_7093,N_3519,N_1184);
nand U7094 (N_7094,N_1011,N_225);
nand U7095 (N_7095,N_3320,N_4851);
or U7096 (N_7096,N_352,N_33);
and U7097 (N_7097,N_4626,N_752);
nor U7098 (N_7098,N_4924,N_4479);
nor U7099 (N_7099,N_2393,N_2427);
and U7100 (N_7100,N_1359,N_512);
nor U7101 (N_7101,N_2591,N_2858);
nand U7102 (N_7102,N_454,N_3901);
or U7103 (N_7103,N_761,N_519);
and U7104 (N_7104,N_2862,N_4993);
xnor U7105 (N_7105,N_2307,N_4592);
nand U7106 (N_7106,N_786,N_3369);
and U7107 (N_7107,N_2553,N_3580);
nand U7108 (N_7108,N_4578,N_3675);
and U7109 (N_7109,N_375,N_1791);
nor U7110 (N_7110,N_362,N_3105);
nand U7111 (N_7111,N_1109,N_2066);
nor U7112 (N_7112,N_115,N_2163);
and U7113 (N_7113,N_1943,N_2928);
and U7114 (N_7114,N_4823,N_520);
and U7115 (N_7115,N_1164,N_237);
or U7116 (N_7116,N_4208,N_487);
nor U7117 (N_7117,N_2612,N_4421);
or U7118 (N_7118,N_2740,N_4791);
and U7119 (N_7119,N_1531,N_1252);
nand U7120 (N_7120,N_3793,N_3886);
nand U7121 (N_7121,N_2866,N_3758);
or U7122 (N_7122,N_1421,N_1546);
xor U7123 (N_7123,N_2746,N_3199);
nand U7124 (N_7124,N_4762,N_1804);
nand U7125 (N_7125,N_1025,N_1592);
nor U7126 (N_7126,N_3807,N_1267);
nand U7127 (N_7127,N_4495,N_274);
nor U7128 (N_7128,N_4836,N_858);
or U7129 (N_7129,N_497,N_4377);
nor U7130 (N_7130,N_1334,N_144);
nand U7131 (N_7131,N_925,N_4908);
or U7132 (N_7132,N_1929,N_111);
and U7133 (N_7133,N_4095,N_113);
xor U7134 (N_7134,N_2077,N_1615);
nand U7135 (N_7135,N_4727,N_4352);
nand U7136 (N_7136,N_921,N_432);
nand U7137 (N_7137,N_1154,N_1136);
nor U7138 (N_7138,N_2619,N_1251);
nand U7139 (N_7139,N_1018,N_2201);
and U7140 (N_7140,N_1054,N_2993);
or U7141 (N_7141,N_1831,N_3211);
or U7142 (N_7142,N_3390,N_3466);
and U7143 (N_7143,N_52,N_1813);
and U7144 (N_7144,N_1144,N_4643);
and U7145 (N_7145,N_1148,N_507);
nor U7146 (N_7146,N_3361,N_2018);
nand U7147 (N_7147,N_510,N_3796);
and U7148 (N_7148,N_581,N_3186);
and U7149 (N_7149,N_4216,N_2944);
and U7150 (N_7150,N_2318,N_2999);
nor U7151 (N_7151,N_685,N_3932);
and U7152 (N_7152,N_3423,N_3865);
nor U7153 (N_7153,N_4079,N_2057);
nand U7154 (N_7154,N_1455,N_3692);
or U7155 (N_7155,N_4930,N_4864);
nor U7156 (N_7156,N_875,N_3988);
nand U7157 (N_7157,N_3889,N_797);
or U7158 (N_7158,N_1510,N_3077);
and U7159 (N_7159,N_584,N_2323);
nand U7160 (N_7160,N_1014,N_4909);
and U7161 (N_7161,N_3467,N_3460);
nand U7162 (N_7162,N_1100,N_1077);
nand U7163 (N_7163,N_2589,N_4128);
and U7164 (N_7164,N_3275,N_419);
nor U7165 (N_7165,N_1595,N_3917);
nand U7166 (N_7166,N_722,N_3497);
or U7167 (N_7167,N_2374,N_4995);
nand U7168 (N_7168,N_4905,N_3177);
nor U7169 (N_7169,N_2568,N_3142);
and U7170 (N_7170,N_458,N_1949);
or U7171 (N_7171,N_410,N_891);
nor U7172 (N_7172,N_1081,N_4130);
nor U7173 (N_7173,N_3818,N_2947);
nor U7174 (N_7174,N_1429,N_4091);
and U7175 (N_7175,N_3686,N_4779);
or U7176 (N_7176,N_1218,N_1959);
or U7177 (N_7177,N_2885,N_1098);
or U7178 (N_7178,N_2203,N_56);
nand U7179 (N_7179,N_4861,N_4734);
nand U7180 (N_7180,N_2294,N_4225);
and U7181 (N_7181,N_1728,N_3103);
nand U7182 (N_7182,N_756,N_4047);
nor U7183 (N_7183,N_2937,N_2218);
nor U7184 (N_7184,N_3406,N_4230);
or U7185 (N_7185,N_3605,N_1603);
or U7186 (N_7186,N_1702,N_216);
and U7187 (N_7187,N_1775,N_290);
or U7188 (N_7188,N_4607,N_720);
or U7189 (N_7189,N_4408,N_1213);
nor U7190 (N_7190,N_3203,N_1397);
nor U7191 (N_7191,N_3371,N_4205);
or U7192 (N_7192,N_4100,N_2702);
and U7193 (N_7193,N_1451,N_1003);
and U7194 (N_7194,N_2104,N_2162);
and U7195 (N_7195,N_905,N_1415);
and U7196 (N_7196,N_1311,N_1815);
nor U7197 (N_7197,N_1172,N_982);
nand U7198 (N_7198,N_809,N_2304);
or U7199 (N_7199,N_596,N_2652);
nand U7200 (N_7200,N_2293,N_2766);
nor U7201 (N_7201,N_2656,N_642);
or U7202 (N_7202,N_4548,N_1384);
nor U7203 (N_7203,N_342,N_1303);
nand U7204 (N_7204,N_3132,N_3113);
or U7205 (N_7205,N_919,N_1253);
or U7206 (N_7206,N_4892,N_4850);
and U7207 (N_7207,N_2957,N_4848);
nand U7208 (N_7208,N_1898,N_767);
xor U7209 (N_7209,N_2399,N_2941);
or U7210 (N_7210,N_641,N_2204);
and U7211 (N_7211,N_189,N_3216);
and U7212 (N_7212,N_1652,N_4889);
nor U7213 (N_7213,N_3133,N_3043);
and U7214 (N_7214,N_252,N_658);
or U7215 (N_7215,N_3161,N_484);
or U7216 (N_7216,N_2397,N_711);
and U7217 (N_7217,N_3960,N_3266);
nor U7218 (N_7218,N_4854,N_4794);
nor U7219 (N_7219,N_1760,N_101);
or U7220 (N_7220,N_329,N_674);
nand U7221 (N_7221,N_3608,N_1544);
and U7222 (N_7222,N_3659,N_2431);
nand U7223 (N_7223,N_2802,N_3762);
nand U7224 (N_7224,N_4312,N_2793);
and U7225 (N_7225,N_4728,N_2406);
nand U7226 (N_7226,N_2807,N_3134);
nand U7227 (N_7227,N_504,N_2645);
nor U7228 (N_7228,N_836,N_3541);
xor U7229 (N_7229,N_2985,N_3101);
and U7230 (N_7230,N_844,N_3002);
and U7231 (N_7231,N_4014,N_1836);
and U7232 (N_7232,N_3823,N_4706);
and U7233 (N_7233,N_2886,N_4448);
nor U7234 (N_7234,N_4855,N_3825);
nor U7235 (N_7235,N_202,N_4415);
nor U7236 (N_7236,N_2797,N_2038);
nor U7237 (N_7237,N_4869,N_4927);
nand U7238 (N_7238,N_2071,N_2182);
or U7239 (N_7239,N_4457,N_2387);
nand U7240 (N_7240,N_123,N_3600);
or U7241 (N_7241,N_3172,N_2176);
nand U7242 (N_7242,N_771,N_3951);
xnor U7243 (N_7243,N_1571,N_3037);
nand U7244 (N_7244,N_4427,N_887);
nand U7245 (N_7245,N_4272,N_4785);
nor U7246 (N_7246,N_1232,N_3933);
or U7247 (N_7247,N_2814,N_4949);
or U7248 (N_7248,N_1524,N_457);
nand U7249 (N_7249,N_1612,N_4180);
nor U7250 (N_7250,N_3262,N_3974);
nand U7251 (N_7251,N_1413,N_4428);
and U7252 (N_7252,N_3795,N_2404);
nand U7253 (N_7253,N_335,N_870);
or U7254 (N_7254,N_3550,N_688);
nand U7255 (N_7255,N_953,N_2997);
and U7256 (N_7256,N_2055,N_1747);
or U7257 (N_7257,N_363,N_544);
and U7258 (N_7258,N_599,N_2668);
or U7259 (N_7259,N_4198,N_1337);
and U7260 (N_7260,N_3432,N_4863);
nand U7261 (N_7261,N_3592,N_854);
nor U7262 (N_7262,N_3366,N_1150);
nor U7263 (N_7263,N_823,N_2045);
and U7264 (N_7264,N_2540,N_1127);
nor U7265 (N_7265,N_3264,N_3538);
nor U7266 (N_7266,N_4493,N_4687);
nor U7267 (N_7267,N_2839,N_880);
nor U7268 (N_7268,N_4811,N_3555);
nor U7269 (N_7269,N_863,N_1887);
and U7270 (N_7270,N_3148,N_1523);
or U7271 (N_7271,N_4173,N_2390);
and U7272 (N_7272,N_3955,N_917);
nand U7273 (N_7273,N_2794,N_4885);
and U7274 (N_7274,N_4849,N_4113);
nand U7275 (N_7275,N_1548,N_1382);
or U7276 (N_7276,N_1539,N_150);
or U7277 (N_7277,N_3391,N_3442);
or U7278 (N_7278,N_4465,N_44);
and U7279 (N_7279,N_3083,N_2667);
and U7280 (N_7280,N_4784,N_568);
nor U7281 (N_7281,N_2160,N_1508);
nand U7282 (N_7282,N_292,N_1286);
and U7283 (N_7283,N_3806,N_1944);
or U7284 (N_7284,N_4635,N_2214);
nor U7285 (N_7285,N_2979,N_3470);
and U7286 (N_7286,N_1772,N_333);
xnor U7287 (N_7287,N_4965,N_2042);
nand U7288 (N_7288,N_934,N_4730);
or U7289 (N_7289,N_3785,N_192);
and U7290 (N_7290,N_479,N_2286);
nor U7291 (N_7291,N_4424,N_2827);
or U7292 (N_7292,N_842,N_3535);
nor U7293 (N_7293,N_93,N_4587);
nor U7294 (N_7294,N_2718,N_4321);
and U7295 (N_7295,N_3655,N_2761);
and U7296 (N_7296,N_518,N_4067);
nand U7297 (N_7297,N_1855,N_4912);
nand U7298 (N_7298,N_3329,N_3426);
and U7299 (N_7299,N_4062,N_276);
nor U7300 (N_7300,N_962,N_131);
nand U7301 (N_7301,N_81,N_2213);
nor U7302 (N_7302,N_1445,N_4226);
nand U7303 (N_7303,N_2669,N_2755);
and U7304 (N_7304,N_3729,N_4663);
nor U7305 (N_7305,N_1787,N_2219);
and U7306 (N_7306,N_488,N_659);
and U7307 (N_7307,N_3080,N_2053);
or U7308 (N_7308,N_2614,N_2770);
or U7309 (N_7309,N_5,N_4344);
or U7310 (N_7310,N_1694,N_920);
nor U7311 (N_7311,N_980,N_1657);
or U7312 (N_7312,N_4689,N_2949);
nor U7313 (N_7313,N_45,N_3166);
and U7314 (N_7314,N_2823,N_4705);
nor U7315 (N_7315,N_1191,N_2630);
nand U7316 (N_7316,N_745,N_4050);
or U7317 (N_7317,N_1983,N_3777);
or U7318 (N_7318,N_4627,N_2698);
and U7319 (N_7319,N_2006,N_2514);
or U7320 (N_7320,N_3961,N_4741);
nand U7321 (N_7321,N_21,N_3705);
or U7322 (N_7322,N_3154,N_3307);
nand U7323 (N_7323,N_813,N_2632);
and U7324 (N_7324,N_3293,N_849);
and U7325 (N_7325,N_4398,N_865);
xnor U7326 (N_7326,N_3276,N_3590);
nand U7327 (N_7327,N_3055,N_2095);
and U7328 (N_7328,N_716,N_1872);
or U7329 (N_7329,N_1913,N_1483);
nor U7330 (N_7330,N_2418,N_3189);
nor U7331 (N_7331,N_1640,N_3378);
and U7332 (N_7332,N_1211,N_195);
nor U7333 (N_7333,N_3794,N_2502);
and U7334 (N_7334,N_1958,N_4324);
nor U7335 (N_7335,N_1851,N_4125);
nand U7336 (N_7336,N_37,N_1561);
and U7337 (N_7337,N_2753,N_2033);
nor U7338 (N_7338,N_125,N_4533);
nor U7339 (N_7339,N_2567,N_2606);
nor U7340 (N_7340,N_1674,N_2575);
and U7341 (N_7341,N_2034,N_1491);
and U7342 (N_7342,N_3570,N_2497);
nand U7343 (N_7343,N_4,N_4679);
and U7344 (N_7344,N_2215,N_1569);
and U7345 (N_7345,N_1756,N_4308);
and U7346 (N_7346,N_2836,N_4538);
nor U7347 (N_7347,N_4033,N_3068);
and U7348 (N_7348,N_850,N_4340);
and U7349 (N_7349,N_2660,N_4617);
nand U7350 (N_7350,N_3347,N_2037);
and U7351 (N_7351,N_2061,N_3626);
nand U7352 (N_7352,N_1925,N_1563);
and U7353 (N_7353,N_1725,N_4251);
nor U7354 (N_7354,N_2473,N_521);
nor U7355 (N_7355,N_1498,N_2009);
and U7356 (N_7356,N_1377,N_7);
nand U7357 (N_7357,N_2386,N_3772);
or U7358 (N_7358,N_2409,N_3835);
nor U7359 (N_7359,N_3061,N_1703);
and U7360 (N_7360,N_1593,N_22);
nand U7361 (N_7361,N_1565,N_1268);
and U7362 (N_7362,N_2784,N_185);
and U7363 (N_7363,N_3265,N_339);
nand U7364 (N_7364,N_860,N_811);
or U7365 (N_7365,N_3473,N_4172);
xor U7366 (N_7366,N_281,N_588);
nand U7367 (N_7367,N_4409,N_4335);
and U7368 (N_7368,N_1305,N_3011);
nor U7369 (N_7369,N_2651,N_313);
nand U7370 (N_7370,N_2434,N_3298);
nor U7371 (N_7371,N_2001,N_1743);
and U7372 (N_7372,N_2615,N_2005);
nand U7373 (N_7373,N_2049,N_1927);
or U7374 (N_7374,N_1315,N_219);
or U7375 (N_7375,N_4467,N_911);
and U7376 (N_7376,N_3454,N_954);
or U7377 (N_7377,N_4938,N_2967);
nor U7378 (N_7378,N_4490,N_1962);
nor U7379 (N_7379,N_4915,N_4433);
or U7380 (N_7380,N_534,N_174);
nand U7381 (N_7381,N_2904,N_1186);
or U7382 (N_7382,N_3532,N_846);
and U7383 (N_7383,N_2029,N_2824);
nor U7384 (N_7384,N_3916,N_2103);
nor U7385 (N_7385,N_1392,N_436);
nor U7386 (N_7386,N_4887,N_2601);
nor U7387 (N_7387,N_4901,N_4102);
and U7388 (N_7388,N_4349,N_1149);
and U7389 (N_7389,N_2875,N_548);
and U7390 (N_7390,N_41,N_248);
nor U7391 (N_7391,N_964,N_4978);
nand U7392 (N_7392,N_552,N_1990);
or U7393 (N_7393,N_1873,N_2920);
and U7394 (N_7394,N_38,N_4710);
or U7395 (N_7395,N_3119,N_3064);
or U7396 (N_7396,N_4240,N_4038);
nor U7397 (N_7397,N_4735,N_1904);
nand U7398 (N_7398,N_3881,N_1030);
or U7399 (N_7399,N_1893,N_2422);
nor U7400 (N_7400,N_4265,N_1767);
nor U7401 (N_7401,N_3632,N_197);
and U7402 (N_7402,N_253,N_4143);
and U7403 (N_7403,N_2183,N_2190);
nor U7404 (N_7404,N_1256,N_3554);
nor U7405 (N_7405,N_915,N_4544);
and U7406 (N_7406,N_2550,N_1987);
nor U7407 (N_7407,N_2079,N_766);
nor U7408 (N_7408,N_415,N_1715);
nand U7409 (N_7409,N_3058,N_725);
and U7410 (N_7410,N_993,N_2359);
or U7411 (N_7411,N_378,N_840);
and U7412 (N_7412,N_1155,N_2093);
or U7413 (N_7413,N_3578,N_715);
nor U7414 (N_7414,N_2826,N_4018);
or U7415 (N_7415,N_926,N_1399);
nor U7416 (N_7416,N_1580,N_3496);
and U7417 (N_7417,N_4541,N_3047);
nand U7418 (N_7418,N_82,N_13);
or U7419 (N_7419,N_2626,N_1533);
and U7420 (N_7420,N_1059,N_1254);
nor U7421 (N_7421,N_2423,N_3104);
or U7422 (N_7422,N_3811,N_1611);
nand U7423 (N_7423,N_207,N_4856);
nor U7424 (N_7424,N_2264,N_2594);
or U7425 (N_7425,N_508,N_1249);
or U7426 (N_7426,N_4516,N_1847);
and U7427 (N_7427,N_1647,N_1825);
nand U7428 (N_7428,N_2496,N_3024);
or U7429 (N_7429,N_1779,N_4270);
or U7430 (N_7430,N_3404,N_918);
nor U7431 (N_7431,N_793,N_4998);
nor U7432 (N_7432,N_2819,N_643);
nor U7433 (N_7433,N_1521,N_2842);
or U7434 (N_7434,N_728,N_4464);
nor U7435 (N_7435,N_4991,N_1879);
nor U7436 (N_7436,N_2428,N_1034);
nor U7437 (N_7437,N_134,N_2737);
or U7438 (N_7438,N_3249,N_1231);
and U7439 (N_7439,N_1190,N_3977);
and U7440 (N_7440,N_778,N_1317);
nor U7441 (N_7441,N_3274,N_3126);
nand U7442 (N_7442,N_1143,N_1200);
or U7443 (N_7443,N_2373,N_3957);
and U7444 (N_7444,N_79,N_163);
and U7445 (N_7445,N_3746,N_4605);
nor U7446 (N_7446,N_1396,N_4677);
and U7447 (N_7447,N_2910,N_1995);
or U7448 (N_7448,N_1108,N_3389);
nor U7449 (N_7449,N_141,N_3261);
or U7450 (N_7450,N_162,N_3897);
nand U7451 (N_7451,N_2762,N_1163);
and U7452 (N_7452,N_3235,N_796);
and U7453 (N_7453,N_2471,N_2118);
nor U7454 (N_7454,N_1012,N_1482);
or U7455 (N_7455,N_4987,N_4343);
or U7456 (N_7456,N_4812,N_1773);
and U7457 (N_7457,N_3629,N_509);
nor U7458 (N_7458,N_2371,N_3995);
or U7459 (N_7459,N_2994,N_2677);
or U7460 (N_7460,N_2585,N_2860);
nor U7461 (N_7461,N_882,N_3330);
nand U7462 (N_7462,N_790,N_1187);
and U7463 (N_7463,N_3812,N_4249);
and U7464 (N_7464,N_1341,N_28);
and U7465 (N_7465,N_2712,N_3315);
nand U7466 (N_7466,N_3575,N_437);
and U7467 (N_7467,N_999,N_2137);
and U7468 (N_7468,N_2569,N_2637);
and U7469 (N_7469,N_1965,N_1709);
or U7470 (N_7470,N_2851,N_2658);
and U7471 (N_7471,N_2843,N_4665);
or U7472 (N_7472,N_3490,N_2943);
and U7473 (N_7473,N_2777,N_2464);
and U7474 (N_7474,N_4253,N_3998);
nor U7475 (N_7475,N_1499,N_740);
and U7476 (N_7476,N_3430,N_3306);
nand U7477 (N_7477,N_356,N_334);
nand U7478 (N_7478,N_1119,N_3560);
or U7479 (N_7479,N_2188,N_1590);
nand U7480 (N_7480,N_3198,N_624);
or U7481 (N_7481,N_2410,N_4616);
nand U7482 (N_7482,N_501,N_3326);
nand U7483 (N_7483,N_1,N_4151);
or U7484 (N_7484,N_4144,N_3412);
nand U7485 (N_7485,N_744,N_3536);
nand U7486 (N_7486,N_551,N_2580);
and U7487 (N_7487,N_40,N_2974);
nand U7488 (N_7488,N_2495,N_319);
nand U7489 (N_7489,N_1135,N_1180);
xor U7490 (N_7490,N_4112,N_2185);
nor U7491 (N_7491,N_1283,N_779);
and U7492 (N_7492,N_928,N_3440);
and U7493 (N_7493,N_4107,N_1236);
or U7494 (N_7494,N_949,N_4337);
and U7495 (N_7495,N_678,N_4096);
nand U7496 (N_7496,N_970,N_478);
nor U7497 (N_7497,N_4808,N_2461);
or U7498 (N_7498,N_3512,N_3780);
nand U7499 (N_7499,N_4203,N_1448);
or U7500 (N_7500,N_273,N_81);
and U7501 (N_7501,N_492,N_2460);
and U7502 (N_7502,N_1279,N_3617);
xor U7503 (N_7503,N_4436,N_127);
nand U7504 (N_7504,N_494,N_4451);
or U7505 (N_7505,N_102,N_2364);
and U7506 (N_7506,N_3666,N_4615);
nand U7507 (N_7507,N_1255,N_2124);
nor U7508 (N_7508,N_3597,N_2842);
and U7509 (N_7509,N_4186,N_2161);
nor U7510 (N_7510,N_4177,N_2937);
and U7511 (N_7511,N_1107,N_3533);
nor U7512 (N_7512,N_4866,N_1562);
and U7513 (N_7513,N_298,N_2753);
and U7514 (N_7514,N_1920,N_877);
or U7515 (N_7515,N_2091,N_3319);
or U7516 (N_7516,N_4373,N_1077);
nand U7517 (N_7517,N_8,N_3867);
and U7518 (N_7518,N_4820,N_3341);
nor U7519 (N_7519,N_1796,N_4320);
or U7520 (N_7520,N_3934,N_1951);
and U7521 (N_7521,N_1406,N_1525);
nor U7522 (N_7522,N_3981,N_3887);
or U7523 (N_7523,N_3108,N_541);
or U7524 (N_7524,N_3642,N_4606);
and U7525 (N_7525,N_193,N_4901);
or U7526 (N_7526,N_3074,N_2432);
nor U7527 (N_7527,N_3616,N_1131);
nand U7528 (N_7528,N_4103,N_2865);
and U7529 (N_7529,N_1276,N_3507);
nor U7530 (N_7530,N_1986,N_2145);
nand U7531 (N_7531,N_3440,N_3651);
nor U7532 (N_7532,N_3907,N_4028);
nor U7533 (N_7533,N_1837,N_4762);
and U7534 (N_7534,N_1405,N_855);
and U7535 (N_7535,N_1754,N_1352);
nor U7536 (N_7536,N_1157,N_726);
nor U7537 (N_7537,N_1279,N_1856);
or U7538 (N_7538,N_4044,N_303);
or U7539 (N_7539,N_513,N_3914);
nor U7540 (N_7540,N_1424,N_3829);
and U7541 (N_7541,N_3210,N_537);
nand U7542 (N_7542,N_626,N_3364);
or U7543 (N_7543,N_1230,N_1203);
or U7544 (N_7544,N_640,N_3888);
nor U7545 (N_7545,N_3904,N_3847);
nor U7546 (N_7546,N_276,N_4132);
or U7547 (N_7547,N_1765,N_1161);
or U7548 (N_7548,N_3129,N_3728);
or U7549 (N_7549,N_1707,N_2976);
nand U7550 (N_7550,N_226,N_631);
nand U7551 (N_7551,N_4174,N_4137);
nor U7552 (N_7552,N_1759,N_706);
and U7553 (N_7553,N_244,N_112);
nor U7554 (N_7554,N_592,N_4425);
or U7555 (N_7555,N_4891,N_4890);
and U7556 (N_7556,N_4980,N_1556);
nand U7557 (N_7557,N_1169,N_1709);
or U7558 (N_7558,N_1248,N_131);
nor U7559 (N_7559,N_3663,N_545);
nor U7560 (N_7560,N_332,N_3994);
nand U7561 (N_7561,N_4181,N_2739);
and U7562 (N_7562,N_1174,N_2952);
nand U7563 (N_7563,N_1745,N_2081);
nor U7564 (N_7564,N_1701,N_2937);
nor U7565 (N_7565,N_4574,N_1567);
nor U7566 (N_7566,N_4727,N_813);
and U7567 (N_7567,N_1292,N_684);
nand U7568 (N_7568,N_781,N_2622);
nor U7569 (N_7569,N_3860,N_3065);
nand U7570 (N_7570,N_3246,N_1640);
nand U7571 (N_7571,N_3036,N_794);
and U7572 (N_7572,N_1154,N_317);
or U7573 (N_7573,N_4814,N_2232);
and U7574 (N_7574,N_2759,N_1926);
nand U7575 (N_7575,N_2603,N_608);
nand U7576 (N_7576,N_3727,N_2460);
and U7577 (N_7577,N_498,N_404);
or U7578 (N_7578,N_263,N_1954);
nor U7579 (N_7579,N_147,N_3370);
and U7580 (N_7580,N_4781,N_456);
and U7581 (N_7581,N_2706,N_4094);
nor U7582 (N_7582,N_4137,N_2008);
nand U7583 (N_7583,N_2558,N_814);
nand U7584 (N_7584,N_4474,N_2597);
and U7585 (N_7585,N_4617,N_2775);
and U7586 (N_7586,N_3770,N_2053);
and U7587 (N_7587,N_940,N_4867);
nor U7588 (N_7588,N_4118,N_4530);
nor U7589 (N_7589,N_4895,N_4352);
and U7590 (N_7590,N_3836,N_1589);
or U7591 (N_7591,N_1781,N_4163);
and U7592 (N_7592,N_4171,N_12);
nor U7593 (N_7593,N_1213,N_1676);
and U7594 (N_7594,N_2402,N_423);
nand U7595 (N_7595,N_257,N_4820);
nor U7596 (N_7596,N_3554,N_2315);
and U7597 (N_7597,N_2335,N_4857);
nor U7598 (N_7598,N_1995,N_4660);
nor U7599 (N_7599,N_4416,N_308);
nor U7600 (N_7600,N_1146,N_4668);
nand U7601 (N_7601,N_3337,N_971);
nor U7602 (N_7602,N_2596,N_4313);
nand U7603 (N_7603,N_4016,N_4615);
nor U7604 (N_7604,N_4459,N_158);
nor U7605 (N_7605,N_4935,N_4890);
or U7606 (N_7606,N_2693,N_292);
nand U7607 (N_7607,N_2292,N_590);
or U7608 (N_7608,N_1493,N_7);
and U7609 (N_7609,N_4301,N_4583);
and U7610 (N_7610,N_4593,N_4368);
and U7611 (N_7611,N_2149,N_634);
or U7612 (N_7612,N_272,N_4039);
and U7613 (N_7613,N_860,N_1673);
nand U7614 (N_7614,N_914,N_188);
or U7615 (N_7615,N_1915,N_4993);
and U7616 (N_7616,N_3466,N_4187);
and U7617 (N_7617,N_4120,N_4662);
and U7618 (N_7618,N_2878,N_2317);
nand U7619 (N_7619,N_3871,N_294);
nand U7620 (N_7620,N_1335,N_3991);
and U7621 (N_7621,N_1306,N_3844);
and U7622 (N_7622,N_3586,N_2527);
nand U7623 (N_7623,N_2,N_3015);
or U7624 (N_7624,N_2668,N_833);
or U7625 (N_7625,N_4138,N_3771);
nand U7626 (N_7626,N_181,N_4544);
or U7627 (N_7627,N_509,N_1637);
nand U7628 (N_7628,N_1966,N_518);
nor U7629 (N_7629,N_89,N_4371);
nor U7630 (N_7630,N_4939,N_4481);
or U7631 (N_7631,N_51,N_2810);
and U7632 (N_7632,N_326,N_3858);
nand U7633 (N_7633,N_3572,N_3071);
nand U7634 (N_7634,N_370,N_1761);
nand U7635 (N_7635,N_984,N_612);
and U7636 (N_7636,N_344,N_390);
or U7637 (N_7637,N_3397,N_2940);
nor U7638 (N_7638,N_2076,N_587);
nor U7639 (N_7639,N_36,N_1399);
xor U7640 (N_7640,N_209,N_1702);
nand U7641 (N_7641,N_781,N_1349);
and U7642 (N_7642,N_4322,N_2797);
nor U7643 (N_7643,N_10,N_1546);
nand U7644 (N_7644,N_2015,N_2312);
or U7645 (N_7645,N_1198,N_2785);
and U7646 (N_7646,N_4178,N_4926);
nor U7647 (N_7647,N_4772,N_2290);
and U7648 (N_7648,N_2520,N_650);
nor U7649 (N_7649,N_3054,N_1293);
nand U7650 (N_7650,N_1495,N_4909);
nor U7651 (N_7651,N_4868,N_6);
nand U7652 (N_7652,N_2905,N_3275);
and U7653 (N_7653,N_96,N_3175);
nand U7654 (N_7654,N_662,N_2223);
nor U7655 (N_7655,N_3102,N_4534);
and U7656 (N_7656,N_1183,N_2898);
nand U7657 (N_7657,N_863,N_4113);
or U7658 (N_7658,N_668,N_2220);
or U7659 (N_7659,N_858,N_547);
and U7660 (N_7660,N_3938,N_2552);
nor U7661 (N_7661,N_4295,N_232);
nor U7662 (N_7662,N_4749,N_4256);
or U7663 (N_7663,N_3933,N_3605);
or U7664 (N_7664,N_2574,N_4849);
or U7665 (N_7665,N_3244,N_4035);
and U7666 (N_7666,N_4878,N_876);
and U7667 (N_7667,N_4885,N_2957);
or U7668 (N_7668,N_128,N_870);
nor U7669 (N_7669,N_3138,N_2936);
nand U7670 (N_7670,N_2780,N_2157);
or U7671 (N_7671,N_4360,N_2445);
nand U7672 (N_7672,N_466,N_769);
or U7673 (N_7673,N_1842,N_4387);
and U7674 (N_7674,N_1753,N_3831);
or U7675 (N_7675,N_3061,N_3229);
or U7676 (N_7676,N_4409,N_4063);
or U7677 (N_7677,N_1338,N_1605);
and U7678 (N_7678,N_4558,N_1113);
xor U7679 (N_7679,N_3900,N_3730);
nand U7680 (N_7680,N_204,N_4204);
or U7681 (N_7681,N_1511,N_1420);
or U7682 (N_7682,N_246,N_2701);
nor U7683 (N_7683,N_1350,N_4327);
or U7684 (N_7684,N_3151,N_4697);
or U7685 (N_7685,N_652,N_3684);
or U7686 (N_7686,N_355,N_4784);
nand U7687 (N_7687,N_3683,N_1983);
or U7688 (N_7688,N_3035,N_3287);
nand U7689 (N_7689,N_2824,N_1424);
or U7690 (N_7690,N_4463,N_4313);
nand U7691 (N_7691,N_3303,N_2101);
and U7692 (N_7692,N_3194,N_4384);
nor U7693 (N_7693,N_3383,N_1317);
nand U7694 (N_7694,N_3264,N_3016);
or U7695 (N_7695,N_1322,N_1422);
or U7696 (N_7696,N_2665,N_3683);
nor U7697 (N_7697,N_2435,N_3126);
nor U7698 (N_7698,N_551,N_2533);
and U7699 (N_7699,N_1658,N_2913);
nand U7700 (N_7700,N_534,N_2799);
or U7701 (N_7701,N_4962,N_4092);
nand U7702 (N_7702,N_1152,N_2241);
xnor U7703 (N_7703,N_289,N_4017);
nand U7704 (N_7704,N_4364,N_1639);
or U7705 (N_7705,N_35,N_3631);
or U7706 (N_7706,N_3244,N_3476);
nor U7707 (N_7707,N_4788,N_72);
nand U7708 (N_7708,N_880,N_719);
nand U7709 (N_7709,N_4733,N_3216);
or U7710 (N_7710,N_2951,N_1993);
nand U7711 (N_7711,N_4428,N_3810);
or U7712 (N_7712,N_1978,N_1582);
and U7713 (N_7713,N_4131,N_3197);
nor U7714 (N_7714,N_2676,N_2414);
and U7715 (N_7715,N_2529,N_4745);
or U7716 (N_7716,N_1154,N_1137);
nand U7717 (N_7717,N_1038,N_2260);
nor U7718 (N_7718,N_211,N_587);
nor U7719 (N_7719,N_1014,N_868);
and U7720 (N_7720,N_3392,N_1315);
nand U7721 (N_7721,N_1270,N_4703);
nand U7722 (N_7722,N_2593,N_591);
nor U7723 (N_7723,N_4306,N_3945);
or U7724 (N_7724,N_825,N_4150);
nor U7725 (N_7725,N_4649,N_2558);
nand U7726 (N_7726,N_289,N_4694);
or U7727 (N_7727,N_2160,N_2704);
or U7728 (N_7728,N_4538,N_1353);
nor U7729 (N_7729,N_2609,N_3270);
or U7730 (N_7730,N_2035,N_3564);
nand U7731 (N_7731,N_2814,N_4991);
and U7732 (N_7732,N_2022,N_1938);
or U7733 (N_7733,N_4706,N_3782);
nand U7734 (N_7734,N_1631,N_3894);
xnor U7735 (N_7735,N_2024,N_3400);
or U7736 (N_7736,N_3435,N_3089);
and U7737 (N_7737,N_2240,N_4792);
and U7738 (N_7738,N_0,N_3241);
and U7739 (N_7739,N_2594,N_226);
nor U7740 (N_7740,N_3495,N_2670);
nand U7741 (N_7741,N_4397,N_4077);
nand U7742 (N_7742,N_4787,N_3057);
nor U7743 (N_7743,N_3210,N_2902);
or U7744 (N_7744,N_3633,N_1663);
and U7745 (N_7745,N_2596,N_1919);
nor U7746 (N_7746,N_788,N_336);
nand U7747 (N_7747,N_748,N_572);
nor U7748 (N_7748,N_3567,N_1955);
or U7749 (N_7749,N_2994,N_1900);
nand U7750 (N_7750,N_4209,N_1296);
nand U7751 (N_7751,N_1719,N_3499);
or U7752 (N_7752,N_3732,N_4550);
xnor U7753 (N_7753,N_3563,N_714);
nand U7754 (N_7754,N_1306,N_2599);
nor U7755 (N_7755,N_435,N_60);
nand U7756 (N_7756,N_3988,N_3577);
or U7757 (N_7757,N_4190,N_1215);
nand U7758 (N_7758,N_2631,N_4954);
nand U7759 (N_7759,N_1118,N_1244);
nor U7760 (N_7760,N_284,N_4717);
and U7761 (N_7761,N_1705,N_3236);
and U7762 (N_7762,N_897,N_1928);
or U7763 (N_7763,N_1162,N_4046);
nor U7764 (N_7764,N_4222,N_1565);
nor U7765 (N_7765,N_4270,N_1053);
nor U7766 (N_7766,N_398,N_2873);
and U7767 (N_7767,N_2614,N_936);
or U7768 (N_7768,N_1572,N_386);
nand U7769 (N_7769,N_2957,N_1696);
xnor U7770 (N_7770,N_114,N_4446);
nor U7771 (N_7771,N_4566,N_989);
or U7772 (N_7772,N_2103,N_2256);
nand U7773 (N_7773,N_2277,N_3973);
and U7774 (N_7774,N_675,N_3646);
nor U7775 (N_7775,N_2466,N_2324);
nand U7776 (N_7776,N_4078,N_2836);
nand U7777 (N_7777,N_2578,N_3187);
nand U7778 (N_7778,N_741,N_4029);
or U7779 (N_7779,N_4446,N_3075);
and U7780 (N_7780,N_2891,N_3762);
nor U7781 (N_7781,N_4142,N_2483);
or U7782 (N_7782,N_1619,N_2390);
or U7783 (N_7783,N_1405,N_1600);
nand U7784 (N_7784,N_628,N_2130);
nand U7785 (N_7785,N_4406,N_4277);
nand U7786 (N_7786,N_4953,N_1826);
or U7787 (N_7787,N_2011,N_3938);
nor U7788 (N_7788,N_4769,N_1105);
and U7789 (N_7789,N_613,N_685);
or U7790 (N_7790,N_1000,N_4327);
and U7791 (N_7791,N_4317,N_181);
nor U7792 (N_7792,N_1693,N_2816);
and U7793 (N_7793,N_3989,N_3760);
and U7794 (N_7794,N_4146,N_3527);
and U7795 (N_7795,N_268,N_2693);
nand U7796 (N_7796,N_2861,N_2850);
xnor U7797 (N_7797,N_2895,N_2463);
xnor U7798 (N_7798,N_4199,N_4506);
or U7799 (N_7799,N_1745,N_1603);
or U7800 (N_7800,N_542,N_4511);
or U7801 (N_7801,N_2513,N_4530);
nor U7802 (N_7802,N_2115,N_321);
and U7803 (N_7803,N_178,N_102);
nand U7804 (N_7804,N_4579,N_873);
nor U7805 (N_7805,N_3803,N_4318);
and U7806 (N_7806,N_2667,N_4604);
and U7807 (N_7807,N_3539,N_2527);
nand U7808 (N_7808,N_590,N_2716);
nor U7809 (N_7809,N_3089,N_2199);
nand U7810 (N_7810,N_1801,N_873);
nor U7811 (N_7811,N_4653,N_3398);
nor U7812 (N_7812,N_3195,N_386);
nand U7813 (N_7813,N_3765,N_1217);
and U7814 (N_7814,N_1303,N_394);
and U7815 (N_7815,N_4356,N_2838);
nor U7816 (N_7816,N_2594,N_166);
nand U7817 (N_7817,N_3275,N_293);
nor U7818 (N_7818,N_1008,N_362);
or U7819 (N_7819,N_3935,N_4133);
and U7820 (N_7820,N_327,N_425);
nand U7821 (N_7821,N_2675,N_1527);
and U7822 (N_7822,N_4053,N_2199);
nor U7823 (N_7823,N_4768,N_1666);
or U7824 (N_7824,N_3852,N_179);
or U7825 (N_7825,N_2349,N_4229);
or U7826 (N_7826,N_2949,N_1104);
and U7827 (N_7827,N_1441,N_3184);
or U7828 (N_7828,N_910,N_435);
and U7829 (N_7829,N_4905,N_2616);
and U7830 (N_7830,N_1003,N_2287);
and U7831 (N_7831,N_1825,N_1146);
nor U7832 (N_7832,N_351,N_2021);
nand U7833 (N_7833,N_2799,N_819);
and U7834 (N_7834,N_1191,N_2835);
nand U7835 (N_7835,N_4444,N_2880);
or U7836 (N_7836,N_770,N_4586);
nand U7837 (N_7837,N_4709,N_2575);
nor U7838 (N_7838,N_1545,N_1496);
nand U7839 (N_7839,N_2862,N_1007);
and U7840 (N_7840,N_3296,N_2038);
nor U7841 (N_7841,N_1326,N_2073);
or U7842 (N_7842,N_4851,N_4640);
nand U7843 (N_7843,N_634,N_2415);
and U7844 (N_7844,N_4111,N_3916);
or U7845 (N_7845,N_907,N_3685);
nand U7846 (N_7846,N_198,N_888);
nand U7847 (N_7847,N_4691,N_1802);
or U7848 (N_7848,N_4617,N_4707);
nor U7849 (N_7849,N_2091,N_4353);
nand U7850 (N_7850,N_2598,N_3677);
nor U7851 (N_7851,N_1354,N_322);
and U7852 (N_7852,N_4454,N_1988);
nor U7853 (N_7853,N_4974,N_2000);
and U7854 (N_7854,N_1235,N_2599);
nand U7855 (N_7855,N_2833,N_697);
nor U7856 (N_7856,N_390,N_3799);
xnor U7857 (N_7857,N_472,N_4430);
and U7858 (N_7858,N_2499,N_780);
nand U7859 (N_7859,N_411,N_30);
nand U7860 (N_7860,N_2103,N_1903);
or U7861 (N_7861,N_3464,N_2792);
or U7862 (N_7862,N_4325,N_3487);
and U7863 (N_7863,N_2498,N_1590);
nand U7864 (N_7864,N_2690,N_2129);
and U7865 (N_7865,N_4071,N_4331);
and U7866 (N_7866,N_23,N_614);
and U7867 (N_7867,N_543,N_593);
nand U7868 (N_7868,N_2403,N_4072);
nand U7869 (N_7869,N_2301,N_4548);
nand U7870 (N_7870,N_3971,N_613);
nand U7871 (N_7871,N_2934,N_948);
and U7872 (N_7872,N_2424,N_1330);
nor U7873 (N_7873,N_2691,N_564);
nand U7874 (N_7874,N_998,N_2030);
and U7875 (N_7875,N_1835,N_3484);
and U7876 (N_7876,N_675,N_2362);
and U7877 (N_7877,N_386,N_1915);
nand U7878 (N_7878,N_4575,N_1708);
nand U7879 (N_7879,N_2912,N_4389);
nand U7880 (N_7880,N_774,N_1699);
nor U7881 (N_7881,N_2945,N_116);
nor U7882 (N_7882,N_766,N_1911);
or U7883 (N_7883,N_710,N_457);
and U7884 (N_7884,N_2169,N_3018);
or U7885 (N_7885,N_2161,N_3705);
or U7886 (N_7886,N_4760,N_846);
nor U7887 (N_7887,N_2937,N_616);
and U7888 (N_7888,N_3291,N_4959);
nor U7889 (N_7889,N_2121,N_2444);
nand U7890 (N_7890,N_2508,N_2115);
nor U7891 (N_7891,N_4223,N_1670);
and U7892 (N_7892,N_3362,N_4449);
or U7893 (N_7893,N_4463,N_4660);
or U7894 (N_7894,N_3064,N_375);
and U7895 (N_7895,N_2705,N_2875);
and U7896 (N_7896,N_2671,N_260);
and U7897 (N_7897,N_1684,N_637);
and U7898 (N_7898,N_4627,N_1300);
nand U7899 (N_7899,N_1005,N_1173);
and U7900 (N_7900,N_3786,N_979);
and U7901 (N_7901,N_3824,N_2909);
and U7902 (N_7902,N_3208,N_4637);
nand U7903 (N_7903,N_4418,N_1395);
or U7904 (N_7904,N_2255,N_943);
nand U7905 (N_7905,N_3815,N_2522);
nor U7906 (N_7906,N_336,N_1854);
nand U7907 (N_7907,N_1758,N_4128);
nor U7908 (N_7908,N_4621,N_2453);
or U7909 (N_7909,N_1430,N_2563);
and U7910 (N_7910,N_829,N_1440);
nand U7911 (N_7911,N_3475,N_4518);
or U7912 (N_7912,N_4510,N_4993);
and U7913 (N_7913,N_4506,N_1455);
and U7914 (N_7914,N_2688,N_1466);
and U7915 (N_7915,N_4108,N_2667);
or U7916 (N_7916,N_3141,N_676);
nand U7917 (N_7917,N_228,N_2984);
nor U7918 (N_7918,N_1304,N_2840);
and U7919 (N_7919,N_3958,N_972);
and U7920 (N_7920,N_3646,N_3650);
nor U7921 (N_7921,N_3487,N_3788);
or U7922 (N_7922,N_3483,N_4461);
nand U7923 (N_7923,N_10,N_2626);
or U7924 (N_7924,N_2602,N_2304);
and U7925 (N_7925,N_2584,N_3144);
and U7926 (N_7926,N_4889,N_1386);
nand U7927 (N_7927,N_4846,N_866);
nand U7928 (N_7928,N_4103,N_4991);
and U7929 (N_7929,N_4703,N_2659);
nand U7930 (N_7930,N_1606,N_801);
nand U7931 (N_7931,N_3357,N_2351);
or U7932 (N_7932,N_1236,N_4971);
and U7933 (N_7933,N_3455,N_4682);
or U7934 (N_7934,N_1570,N_391);
nor U7935 (N_7935,N_2647,N_2449);
nor U7936 (N_7936,N_3539,N_2267);
or U7937 (N_7937,N_3788,N_1017);
or U7938 (N_7938,N_750,N_4328);
nor U7939 (N_7939,N_3951,N_2152);
or U7940 (N_7940,N_726,N_672);
or U7941 (N_7941,N_2097,N_622);
and U7942 (N_7942,N_375,N_1991);
nor U7943 (N_7943,N_4452,N_4828);
or U7944 (N_7944,N_2680,N_180);
and U7945 (N_7945,N_4645,N_2771);
or U7946 (N_7946,N_2626,N_2250);
and U7947 (N_7947,N_747,N_1754);
nor U7948 (N_7948,N_4109,N_3437);
and U7949 (N_7949,N_997,N_886);
nand U7950 (N_7950,N_3001,N_1769);
or U7951 (N_7951,N_1406,N_4539);
and U7952 (N_7952,N_2493,N_4579);
and U7953 (N_7953,N_2237,N_172);
nor U7954 (N_7954,N_4468,N_1494);
or U7955 (N_7955,N_2417,N_3097);
nor U7956 (N_7956,N_65,N_3724);
nand U7957 (N_7957,N_3266,N_137);
nand U7958 (N_7958,N_4507,N_1662);
or U7959 (N_7959,N_3892,N_806);
and U7960 (N_7960,N_967,N_3681);
or U7961 (N_7961,N_1701,N_746);
and U7962 (N_7962,N_566,N_1025);
nor U7963 (N_7963,N_2631,N_3892);
nand U7964 (N_7964,N_1432,N_409);
nor U7965 (N_7965,N_883,N_622);
nand U7966 (N_7966,N_961,N_3147);
and U7967 (N_7967,N_3296,N_4744);
nand U7968 (N_7968,N_3355,N_2111);
or U7969 (N_7969,N_2148,N_1984);
nand U7970 (N_7970,N_4278,N_4937);
or U7971 (N_7971,N_2185,N_1738);
xor U7972 (N_7972,N_1886,N_763);
nand U7973 (N_7973,N_4560,N_695);
and U7974 (N_7974,N_3861,N_3641);
nor U7975 (N_7975,N_703,N_1859);
nor U7976 (N_7976,N_2206,N_2948);
or U7977 (N_7977,N_371,N_1476);
nor U7978 (N_7978,N_1382,N_4677);
nor U7979 (N_7979,N_182,N_2680);
nor U7980 (N_7980,N_1214,N_2805);
nor U7981 (N_7981,N_4186,N_179);
nor U7982 (N_7982,N_2729,N_406);
and U7983 (N_7983,N_4288,N_3373);
or U7984 (N_7984,N_754,N_4869);
xor U7985 (N_7985,N_4361,N_1075);
nand U7986 (N_7986,N_4113,N_3310);
nor U7987 (N_7987,N_2614,N_2710);
and U7988 (N_7988,N_1792,N_4831);
or U7989 (N_7989,N_2244,N_3346);
and U7990 (N_7990,N_3955,N_2593);
nand U7991 (N_7991,N_917,N_1521);
or U7992 (N_7992,N_1794,N_4832);
or U7993 (N_7993,N_3328,N_900);
and U7994 (N_7994,N_3807,N_3540);
nor U7995 (N_7995,N_930,N_2011);
or U7996 (N_7996,N_2370,N_1281);
nor U7997 (N_7997,N_1868,N_344);
or U7998 (N_7998,N_2196,N_4719);
and U7999 (N_7999,N_711,N_3194);
nand U8000 (N_8000,N_524,N_1008);
or U8001 (N_8001,N_1230,N_640);
and U8002 (N_8002,N_3027,N_2701);
or U8003 (N_8003,N_2225,N_4890);
or U8004 (N_8004,N_2816,N_4066);
nor U8005 (N_8005,N_4151,N_4964);
and U8006 (N_8006,N_1795,N_2673);
xor U8007 (N_8007,N_4576,N_2543);
or U8008 (N_8008,N_691,N_1337);
nand U8009 (N_8009,N_2271,N_4113);
or U8010 (N_8010,N_592,N_1550);
or U8011 (N_8011,N_971,N_3138);
nand U8012 (N_8012,N_251,N_3820);
and U8013 (N_8013,N_49,N_45);
or U8014 (N_8014,N_4292,N_341);
or U8015 (N_8015,N_2429,N_27);
nor U8016 (N_8016,N_305,N_1034);
nand U8017 (N_8017,N_4180,N_761);
or U8018 (N_8018,N_2342,N_2489);
nor U8019 (N_8019,N_1817,N_454);
nand U8020 (N_8020,N_2036,N_3665);
and U8021 (N_8021,N_1294,N_698);
and U8022 (N_8022,N_443,N_3310);
or U8023 (N_8023,N_2843,N_463);
xnor U8024 (N_8024,N_614,N_2170);
nand U8025 (N_8025,N_4545,N_4189);
and U8026 (N_8026,N_4746,N_1317);
nand U8027 (N_8027,N_71,N_2312);
and U8028 (N_8028,N_2471,N_1443);
and U8029 (N_8029,N_3384,N_210);
or U8030 (N_8030,N_3580,N_3702);
or U8031 (N_8031,N_2013,N_266);
and U8032 (N_8032,N_1405,N_3072);
nor U8033 (N_8033,N_3512,N_4502);
nor U8034 (N_8034,N_870,N_3790);
and U8035 (N_8035,N_4287,N_3771);
or U8036 (N_8036,N_2230,N_4033);
nor U8037 (N_8037,N_1124,N_4030);
nor U8038 (N_8038,N_2178,N_1388);
or U8039 (N_8039,N_4834,N_2255);
nand U8040 (N_8040,N_2058,N_1276);
and U8041 (N_8041,N_1814,N_1301);
and U8042 (N_8042,N_4939,N_4729);
and U8043 (N_8043,N_2038,N_803);
nand U8044 (N_8044,N_1530,N_3725);
nor U8045 (N_8045,N_2258,N_4453);
nand U8046 (N_8046,N_3523,N_510);
nand U8047 (N_8047,N_392,N_1492);
and U8048 (N_8048,N_4662,N_2429);
and U8049 (N_8049,N_688,N_1152);
nor U8050 (N_8050,N_413,N_2369);
and U8051 (N_8051,N_840,N_3121);
nor U8052 (N_8052,N_1409,N_4345);
and U8053 (N_8053,N_4451,N_98);
or U8054 (N_8054,N_66,N_2384);
nand U8055 (N_8055,N_4706,N_2363);
or U8056 (N_8056,N_2630,N_3934);
nand U8057 (N_8057,N_3082,N_4015);
or U8058 (N_8058,N_1533,N_2311);
and U8059 (N_8059,N_643,N_1719);
nor U8060 (N_8060,N_245,N_2224);
nor U8061 (N_8061,N_1024,N_910);
nand U8062 (N_8062,N_2920,N_3650);
and U8063 (N_8063,N_1120,N_1034);
or U8064 (N_8064,N_574,N_2079);
nand U8065 (N_8065,N_165,N_2452);
or U8066 (N_8066,N_3924,N_1507);
or U8067 (N_8067,N_4088,N_4111);
and U8068 (N_8068,N_2547,N_3640);
and U8069 (N_8069,N_538,N_2383);
and U8070 (N_8070,N_3248,N_4183);
or U8071 (N_8071,N_2894,N_3295);
nor U8072 (N_8072,N_4229,N_1753);
xnor U8073 (N_8073,N_2136,N_3074);
nand U8074 (N_8074,N_3532,N_300);
nor U8075 (N_8075,N_3364,N_3487);
nand U8076 (N_8076,N_2956,N_1258);
and U8077 (N_8077,N_1046,N_2287);
and U8078 (N_8078,N_1956,N_273);
xnor U8079 (N_8079,N_3291,N_1806);
nor U8080 (N_8080,N_1649,N_156);
and U8081 (N_8081,N_3804,N_4217);
nand U8082 (N_8082,N_894,N_759);
and U8083 (N_8083,N_3078,N_2353);
nand U8084 (N_8084,N_2413,N_3996);
and U8085 (N_8085,N_526,N_4276);
or U8086 (N_8086,N_4584,N_3304);
or U8087 (N_8087,N_1057,N_3895);
nand U8088 (N_8088,N_1098,N_4006);
nor U8089 (N_8089,N_751,N_37);
nand U8090 (N_8090,N_1853,N_3731);
xnor U8091 (N_8091,N_3860,N_1047);
nor U8092 (N_8092,N_999,N_1098);
nand U8093 (N_8093,N_839,N_2976);
and U8094 (N_8094,N_4040,N_2087);
nor U8095 (N_8095,N_1524,N_874);
or U8096 (N_8096,N_1087,N_2635);
and U8097 (N_8097,N_630,N_1315);
nor U8098 (N_8098,N_4458,N_2755);
nand U8099 (N_8099,N_1726,N_2300);
or U8100 (N_8100,N_2124,N_774);
nand U8101 (N_8101,N_3328,N_3016);
nand U8102 (N_8102,N_2406,N_49);
nor U8103 (N_8103,N_4094,N_2139);
and U8104 (N_8104,N_4405,N_2155);
nand U8105 (N_8105,N_217,N_3209);
nor U8106 (N_8106,N_4420,N_3231);
nand U8107 (N_8107,N_4807,N_1535);
or U8108 (N_8108,N_1158,N_4360);
and U8109 (N_8109,N_3252,N_4832);
nor U8110 (N_8110,N_1624,N_3421);
nand U8111 (N_8111,N_4495,N_1269);
and U8112 (N_8112,N_2277,N_3175);
and U8113 (N_8113,N_4030,N_4478);
nand U8114 (N_8114,N_3846,N_2822);
or U8115 (N_8115,N_4519,N_3196);
nand U8116 (N_8116,N_3511,N_3017);
and U8117 (N_8117,N_2516,N_1838);
and U8118 (N_8118,N_665,N_446);
and U8119 (N_8119,N_4756,N_3390);
and U8120 (N_8120,N_20,N_1345);
and U8121 (N_8121,N_3898,N_2733);
and U8122 (N_8122,N_2748,N_2867);
or U8123 (N_8123,N_976,N_2488);
nand U8124 (N_8124,N_2363,N_3208);
and U8125 (N_8125,N_2620,N_2109);
nand U8126 (N_8126,N_3392,N_376);
and U8127 (N_8127,N_2793,N_159);
or U8128 (N_8128,N_3793,N_2724);
or U8129 (N_8129,N_647,N_180);
nand U8130 (N_8130,N_3903,N_3356);
and U8131 (N_8131,N_975,N_3867);
and U8132 (N_8132,N_4802,N_1236);
nand U8133 (N_8133,N_4410,N_4556);
and U8134 (N_8134,N_720,N_3136);
nand U8135 (N_8135,N_1117,N_4648);
nand U8136 (N_8136,N_2650,N_1532);
and U8137 (N_8137,N_1027,N_2135);
nand U8138 (N_8138,N_2395,N_1105);
nor U8139 (N_8139,N_4624,N_1193);
nand U8140 (N_8140,N_1958,N_4527);
nor U8141 (N_8141,N_1459,N_3985);
nor U8142 (N_8142,N_1373,N_4278);
and U8143 (N_8143,N_371,N_4044);
and U8144 (N_8144,N_4848,N_2552);
or U8145 (N_8145,N_1021,N_1158);
or U8146 (N_8146,N_1166,N_3121);
or U8147 (N_8147,N_642,N_2784);
nand U8148 (N_8148,N_3651,N_2762);
or U8149 (N_8149,N_2451,N_3208);
and U8150 (N_8150,N_1573,N_3665);
nor U8151 (N_8151,N_4033,N_447);
nand U8152 (N_8152,N_187,N_3045);
and U8153 (N_8153,N_1767,N_59);
nor U8154 (N_8154,N_507,N_817);
or U8155 (N_8155,N_1686,N_1405);
nor U8156 (N_8156,N_1747,N_4323);
nor U8157 (N_8157,N_4062,N_4867);
and U8158 (N_8158,N_2021,N_1454);
nand U8159 (N_8159,N_4555,N_3357);
nand U8160 (N_8160,N_3603,N_1137);
or U8161 (N_8161,N_2194,N_2470);
nand U8162 (N_8162,N_2052,N_2137);
and U8163 (N_8163,N_955,N_1285);
nand U8164 (N_8164,N_2738,N_2128);
nor U8165 (N_8165,N_2109,N_1215);
nor U8166 (N_8166,N_1308,N_1553);
and U8167 (N_8167,N_2604,N_3579);
or U8168 (N_8168,N_2937,N_1760);
and U8169 (N_8169,N_2129,N_4453);
and U8170 (N_8170,N_2807,N_3135);
nor U8171 (N_8171,N_3387,N_105);
nor U8172 (N_8172,N_1762,N_4361);
nand U8173 (N_8173,N_4287,N_4970);
nor U8174 (N_8174,N_3822,N_593);
nand U8175 (N_8175,N_2763,N_657);
or U8176 (N_8176,N_4517,N_1496);
nand U8177 (N_8177,N_3120,N_3042);
nor U8178 (N_8178,N_3983,N_982);
and U8179 (N_8179,N_1619,N_2655);
nor U8180 (N_8180,N_1681,N_2987);
nand U8181 (N_8181,N_3709,N_1079);
and U8182 (N_8182,N_4949,N_43);
and U8183 (N_8183,N_2507,N_4766);
or U8184 (N_8184,N_2656,N_4447);
and U8185 (N_8185,N_1933,N_2884);
nand U8186 (N_8186,N_2723,N_2768);
nand U8187 (N_8187,N_2097,N_1757);
and U8188 (N_8188,N_3466,N_2429);
nor U8189 (N_8189,N_122,N_8);
and U8190 (N_8190,N_2882,N_3631);
and U8191 (N_8191,N_1816,N_752);
or U8192 (N_8192,N_4309,N_4346);
nand U8193 (N_8193,N_571,N_1553);
nor U8194 (N_8194,N_2622,N_971);
and U8195 (N_8195,N_3228,N_4788);
nor U8196 (N_8196,N_122,N_1873);
nand U8197 (N_8197,N_749,N_491);
and U8198 (N_8198,N_1669,N_1985);
and U8199 (N_8199,N_4554,N_874);
nand U8200 (N_8200,N_648,N_4819);
or U8201 (N_8201,N_1618,N_1105);
nand U8202 (N_8202,N_750,N_1068);
and U8203 (N_8203,N_4242,N_4591);
or U8204 (N_8204,N_1711,N_3496);
and U8205 (N_8205,N_4066,N_3890);
nand U8206 (N_8206,N_2246,N_3519);
or U8207 (N_8207,N_1063,N_996);
nor U8208 (N_8208,N_3859,N_741);
or U8209 (N_8209,N_558,N_2643);
nor U8210 (N_8210,N_58,N_1945);
nand U8211 (N_8211,N_1714,N_2087);
or U8212 (N_8212,N_1037,N_4361);
and U8213 (N_8213,N_737,N_3142);
nand U8214 (N_8214,N_2282,N_4971);
nor U8215 (N_8215,N_4013,N_3694);
and U8216 (N_8216,N_400,N_3260);
and U8217 (N_8217,N_3419,N_4509);
and U8218 (N_8218,N_2275,N_935);
or U8219 (N_8219,N_4646,N_747);
or U8220 (N_8220,N_4726,N_2484);
and U8221 (N_8221,N_3716,N_479);
nor U8222 (N_8222,N_990,N_3728);
and U8223 (N_8223,N_2322,N_2414);
nand U8224 (N_8224,N_964,N_3217);
and U8225 (N_8225,N_2693,N_161);
nor U8226 (N_8226,N_3928,N_962);
and U8227 (N_8227,N_2610,N_776);
nor U8228 (N_8228,N_2853,N_3368);
nand U8229 (N_8229,N_1260,N_4155);
or U8230 (N_8230,N_1222,N_3253);
and U8231 (N_8231,N_2215,N_3366);
or U8232 (N_8232,N_3302,N_963);
nand U8233 (N_8233,N_4837,N_4174);
or U8234 (N_8234,N_3805,N_447);
nor U8235 (N_8235,N_3966,N_4377);
nand U8236 (N_8236,N_4027,N_3988);
or U8237 (N_8237,N_1628,N_3209);
nand U8238 (N_8238,N_593,N_4895);
or U8239 (N_8239,N_3729,N_2187);
nor U8240 (N_8240,N_4068,N_755);
nand U8241 (N_8241,N_326,N_1248);
nand U8242 (N_8242,N_3268,N_847);
nor U8243 (N_8243,N_3803,N_2397);
and U8244 (N_8244,N_2629,N_1968);
nor U8245 (N_8245,N_4345,N_3128);
nor U8246 (N_8246,N_945,N_4195);
nand U8247 (N_8247,N_514,N_3359);
nor U8248 (N_8248,N_2202,N_243);
and U8249 (N_8249,N_2898,N_2226);
nand U8250 (N_8250,N_3169,N_2483);
nand U8251 (N_8251,N_143,N_3758);
and U8252 (N_8252,N_939,N_640);
or U8253 (N_8253,N_3624,N_4837);
or U8254 (N_8254,N_2859,N_2912);
nand U8255 (N_8255,N_2609,N_2489);
or U8256 (N_8256,N_1744,N_208);
and U8257 (N_8257,N_78,N_2644);
xnor U8258 (N_8258,N_602,N_3411);
nor U8259 (N_8259,N_2520,N_2065);
or U8260 (N_8260,N_2977,N_3918);
or U8261 (N_8261,N_1300,N_640);
nor U8262 (N_8262,N_3874,N_862);
or U8263 (N_8263,N_3893,N_413);
and U8264 (N_8264,N_3283,N_2104);
nor U8265 (N_8265,N_4933,N_3180);
and U8266 (N_8266,N_3907,N_3615);
and U8267 (N_8267,N_151,N_2384);
or U8268 (N_8268,N_623,N_3557);
and U8269 (N_8269,N_1393,N_1090);
or U8270 (N_8270,N_247,N_30);
nand U8271 (N_8271,N_4673,N_4817);
and U8272 (N_8272,N_1381,N_393);
and U8273 (N_8273,N_311,N_2811);
nand U8274 (N_8274,N_1548,N_1743);
nand U8275 (N_8275,N_2103,N_1280);
nor U8276 (N_8276,N_3392,N_4199);
nor U8277 (N_8277,N_3442,N_4663);
and U8278 (N_8278,N_2557,N_1560);
nand U8279 (N_8279,N_3171,N_335);
or U8280 (N_8280,N_520,N_2050);
or U8281 (N_8281,N_404,N_1869);
nand U8282 (N_8282,N_2380,N_4166);
and U8283 (N_8283,N_4121,N_2248);
nor U8284 (N_8284,N_4132,N_4530);
nand U8285 (N_8285,N_193,N_2428);
nand U8286 (N_8286,N_3268,N_598);
and U8287 (N_8287,N_1964,N_4952);
and U8288 (N_8288,N_3189,N_1537);
and U8289 (N_8289,N_1171,N_4892);
or U8290 (N_8290,N_4963,N_1558);
or U8291 (N_8291,N_2584,N_608);
or U8292 (N_8292,N_4982,N_3370);
and U8293 (N_8293,N_4022,N_4767);
nand U8294 (N_8294,N_4266,N_1729);
or U8295 (N_8295,N_2905,N_4018);
and U8296 (N_8296,N_3757,N_2645);
nand U8297 (N_8297,N_133,N_1693);
nor U8298 (N_8298,N_3399,N_2627);
nand U8299 (N_8299,N_603,N_4557);
or U8300 (N_8300,N_305,N_3854);
or U8301 (N_8301,N_780,N_4089);
or U8302 (N_8302,N_2909,N_1806);
or U8303 (N_8303,N_3078,N_404);
nor U8304 (N_8304,N_3702,N_2334);
and U8305 (N_8305,N_3895,N_3414);
or U8306 (N_8306,N_4345,N_4461);
nor U8307 (N_8307,N_4596,N_1750);
or U8308 (N_8308,N_3697,N_1153);
nand U8309 (N_8309,N_3257,N_4176);
and U8310 (N_8310,N_1214,N_1789);
nor U8311 (N_8311,N_1729,N_2656);
or U8312 (N_8312,N_2784,N_234);
or U8313 (N_8313,N_597,N_893);
or U8314 (N_8314,N_3810,N_3016);
or U8315 (N_8315,N_1632,N_2595);
nand U8316 (N_8316,N_2913,N_4259);
or U8317 (N_8317,N_4508,N_3535);
or U8318 (N_8318,N_3616,N_2313);
nand U8319 (N_8319,N_2054,N_1281);
or U8320 (N_8320,N_3985,N_1892);
or U8321 (N_8321,N_2027,N_2655);
nand U8322 (N_8322,N_1187,N_3246);
nand U8323 (N_8323,N_4015,N_146);
or U8324 (N_8324,N_672,N_1902);
nand U8325 (N_8325,N_3099,N_1812);
or U8326 (N_8326,N_456,N_4211);
and U8327 (N_8327,N_3543,N_3448);
or U8328 (N_8328,N_4647,N_3680);
and U8329 (N_8329,N_899,N_2171);
nand U8330 (N_8330,N_3067,N_3588);
nor U8331 (N_8331,N_1592,N_2374);
or U8332 (N_8332,N_97,N_80);
nand U8333 (N_8333,N_327,N_3713);
nor U8334 (N_8334,N_82,N_1734);
or U8335 (N_8335,N_3110,N_1256);
or U8336 (N_8336,N_1436,N_3878);
nand U8337 (N_8337,N_1748,N_2543);
nor U8338 (N_8338,N_1686,N_1514);
or U8339 (N_8339,N_2672,N_3698);
nor U8340 (N_8340,N_662,N_2388);
nor U8341 (N_8341,N_726,N_3993);
or U8342 (N_8342,N_458,N_844);
nand U8343 (N_8343,N_1737,N_3235);
or U8344 (N_8344,N_2090,N_2616);
or U8345 (N_8345,N_95,N_3549);
and U8346 (N_8346,N_670,N_1694);
nand U8347 (N_8347,N_2408,N_4485);
or U8348 (N_8348,N_2714,N_4425);
nand U8349 (N_8349,N_325,N_958);
and U8350 (N_8350,N_934,N_1470);
nand U8351 (N_8351,N_4209,N_3428);
or U8352 (N_8352,N_441,N_4306);
nor U8353 (N_8353,N_2236,N_2653);
nand U8354 (N_8354,N_4711,N_3024);
nor U8355 (N_8355,N_1193,N_3938);
and U8356 (N_8356,N_435,N_3260);
or U8357 (N_8357,N_1540,N_4907);
and U8358 (N_8358,N_3896,N_377);
or U8359 (N_8359,N_3821,N_3883);
and U8360 (N_8360,N_284,N_3647);
nor U8361 (N_8361,N_4498,N_4255);
nor U8362 (N_8362,N_3571,N_3229);
nand U8363 (N_8363,N_3211,N_1329);
nand U8364 (N_8364,N_1715,N_981);
and U8365 (N_8365,N_3804,N_434);
and U8366 (N_8366,N_4184,N_2557);
nand U8367 (N_8367,N_2739,N_1639);
and U8368 (N_8368,N_1638,N_4305);
or U8369 (N_8369,N_1410,N_954);
nand U8370 (N_8370,N_4057,N_2559);
nand U8371 (N_8371,N_3700,N_1818);
nand U8372 (N_8372,N_4940,N_279);
and U8373 (N_8373,N_946,N_1186);
and U8374 (N_8374,N_2458,N_1035);
xnor U8375 (N_8375,N_1218,N_466);
or U8376 (N_8376,N_39,N_267);
or U8377 (N_8377,N_4481,N_3414);
or U8378 (N_8378,N_2639,N_2225);
and U8379 (N_8379,N_3216,N_590);
or U8380 (N_8380,N_4397,N_130);
and U8381 (N_8381,N_3638,N_4337);
nor U8382 (N_8382,N_3262,N_4649);
and U8383 (N_8383,N_2332,N_4772);
and U8384 (N_8384,N_2670,N_717);
nor U8385 (N_8385,N_576,N_1222);
nand U8386 (N_8386,N_4350,N_2008);
nor U8387 (N_8387,N_4673,N_3774);
and U8388 (N_8388,N_2277,N_3222);
or U8389 (N_8389,N_13,N_3961);
or U8390 (N_8390,N_3386,N_447);
and U8391 (N_8391,N_2621,N_2235);
and U8392 (N_8392,N_3300,N_377);
nor U8393 (N_8393,N_1369,N_895);
or U8394 (N_8394,N_1499,N_2490);
nand U8395 (N_8395,N_2575,N_365);
or U8396 (N_8396,N_3408,N_1444);
nor U8397 (N_8397,N_1349,N_4813);
or U8398 (N_8398,N_1485,N_2067);
nand U8399 (N_8399,N_3046,N_757);
xor U8400 (N_8400,N_637,N_508);
nor U8401 (N_8401,N_3686,N_4087);
or U8402 (N_8402,N_1068,N_4476);
nand U8403 (N_8403,N_4828,N_3150);
nand U8404 (N_8404,N_1590,N_2440);
nor U8405 (N_8405,N_3463,N_1449);
nor U8406 (N_8406,N_2688,N_1889);
or U8407 (N_8407,N_2445,N_1323);
nor U8408 (N_8408,N_3593,N_589);
nor U8409 (N_8409,N_1788,N_1824);
and U8410 (N_8410,N_1250,N_1755);
nor U8411 (N_8411,N_2019,N_3930);
nor U8412 (N_8412,N_1317,N_2784);
or U8413 (N_8413,N_1353,N_265);
nand U8414 (N_8414,N_2100,N_4956);
nor U8415 (N_8415,N_4815,N_3862);
and U8416 (N_8416,N_3789,N_1181);
and U8417 (N_8417,N_4347,N_1713);
nor U8418 (N_8418,N_2427,N_4763);
nand U8419 (N_8419,N_3243,N_3159);
nor U8420 (N_8420,N_2256,N_1811);
and U8421 (N_8421,N_1899,N_944);
and U8422 (N_8422,N_3283,N_3997);
nor U8423 (N_8423,N_240,N_923);
and U8424 (N_8424,N_1719,N_2649);
and U8425 (N_8425,N_2544,N_3071);
nand U8426 (N_8426,N_2587,N_4006);
and U8427 (N_8427,N_54,N_4652);
or U8428 (N_8428,N_1974,N_3231);
or U8429 (N_8429,N_4497,N_2615);
nor U8430 (N_8430,N_747,N_4759);
and U8431 (N_8431,N_886,N_1613);
nand U8432 (N_8432,N_4465,N_3705);
or U8433 (N_8433,N_1012,N_794);
or U8434 (N_8434,N_2205,N_773);
nand U8435 (N_8435,N_708,N_2492);
nor U8436 (N_8436,N_3627,N_1464);
and U8437 (N_8437,N_5,N_3124);
nor U8438 (N_8438,N_4729,N_2672);
or U8439 (N_8439,N_4754,N_3662);
and U8440 (N_8440,N_1671,N_4634);
or U8441 (N_8441,N_1632,N_4508);
nand U8442 (N_8442,N_3223,N_4420);
and U8443 (N_8443,N_3203,N_1417);
or U8444 (N_8444,N_842,N_4838);
nand U8445 (N_8445,N_4089,N_3986);
nor U8446 (N_8446,N_3499,N_1628);
or U8447 (N_8447,N_1780,N_448);
and U8448 (N_8448,N_1334,N_3707);
nand U8449 (N_8449,N_4143,N_118);
and U8450 (N_8450,N_4395,N_58);
nand U8451 (N_8451,N_1319,N_3295);
nand U8452 (N_8452,N_1987,N_765);
nand U8453 (N_8453,N_273,N_255);
and U8454 (N_8454,N_1731,N_3093);
and U8455 (N_8455,N_3210,N_3189);
nand U8456 (N_8456,N_3689,N_4688);
nor U8457 (N_8457,N_4169,N_790);
nand U8458 (N_8458,N_4196,N_2570);
or U8459 (N_8459,N_1455,N_2660);
or U8460 (N_8460,N_1437,N_4040);
nor U8461 (N_8461,N_1918,N_4395);
nor U8462 (N_8462,N_3450,N_3171);
and U8463 (N_8463,N_1674,N_798);
nand U8464 (N_8464,N_4331,N_3092);
nand U8465 (N_8465,N_1230,N_3396);
nand U8466 (N_8466,N_3316,N_2473);
or U8467 (N_8467,N_3935,N_3194);
nand U8468 (N_8468,N_3386,N_2952);
nor U8469 (N_8469,N_1082,N_119);
nand U8470 (N_8470,N_2795,N_1387);
nand U8471 (N_8471,N_4283,N_3520);
nand U8472 (N_8472,N_2280,N_1564);
nand U8473 (N_8473,N_2704,N_3242);
nor U8474 (N_8474,N_759,N_3191);
or U8475 (N_8475,N_2847,N_3945);
and U8476 (N_8476,N_579,N_3428);
and U8477 (N_8477,N_53,N_4902);
nor U8478 (N_8478,N_3732,N_4788);
nand U8479 (N_8479,N_4746,N_4781);
xor U8480 (N_8480,N_2832,N_553);
nor U8481 (N_8481,N_1457,N_1855);
nand U8482 (N_8482,N_3442,N_1531);
and U8483 (N_8483,N_1116,N_4237);
and U8484 (N_8484,N_3335,N_3947);
or U8485 (N_8485,N_3239,N_447);
and U8486 (N_8486,N_2828,N_4212);
nand U8487 (N_8487,N_1924,N_2412);
nand U8488 (N_8488,N_2977,N_4379);
or U8489 (N_8489,N_3877,N_290);
or U8490 (N_8490,N_2680,N_4026);
nor U8491 (N_8491,N_2210,N_1311);
and U8492 (N_8492,N_4611,N_919);
nor U8493 (N_8493,N_2776,N_523);
nor U8494 (N_8494,N_3253,N_726);
nor U8495 (N_8495,N_4755,N_4376);
or U8496 (N_8496,N_1812,N_293);
nand U8497 (N_8497,N_4583,N_3759);
and U8498 (N_8498,N_1835,N_3003);
nand U8499 (N_8499,N_1399,N_365);
nand U8500 (N_8500,N_1391,N_552);
or U8501 (N_8501,N_4937,N_926);
nor U8502 (N_8502,N_1171,N_4699);
nor U8503 (N_8503,N_516,N_1469);
nor U8504 (N_8504,N_1098,N_3957);
nor U8505 (N_8505,N_4779,N_421);
nor U8506 (N_8506,N_2544,N_3347);
nor U8507 (N_8507,N_2720,N_636);
and U8508 (N_8508,N_3456,N_3860);
and U8509 (N_8509,N_419,N_669);
nor U8510 (N_8510,N_4048,N_3705);
and U8511 (N_8511,N_3237,N_1504);
nor U8512 (N_8512,N_2346,N_1825);
and U8513 (N_8513,N_2466,N_608);
nand U8514 (N_8514,N_4233,N_578);
nand U8515 (N_8515,N_773,N_3487);
nor U8516 (N_8516,N_901,N_2446);
and U8517 (N_8517,N_3133,N_1431);
and U8518 (N_8518,N_3869,N_2527);
nand U8519 (N_8519,N_2231,N_389);
nand U8520 (N_8520,N_1171,N_902);
nand U8521 (N_8521,N_2976,N_1061);
nand U8522 (N_8522,N_942,N_2789);
and U8523 (N_8523,N_3441,N_3987);
nand U8524 (N_8524,N_2253,N_4477);
nor U8525 (N_8525,N_3036,N_1060);
nand U8526 (N_8526,N_1436,N_1030);
or U8527 (N_8527,N_4963,N_2181);
nor U8528 (N_8528,N_1562,N_2995);
and U8529 (N_8529,N_644,N_4919);
nand U8530 (N_8530,N_328,N_4277);
and U8531 (N_8531,N_317,N_1471);
and U8532 (N_8532,N_4462,N_2586);
or U8533 (N_8533,N_1258,N_4026);
nor U8534 (N_8534,N_2922,N_1101);
and U8535 (N_8535,N_4375,N_1903);
and U8536 (N_8536,N_3001,N_1511);
and U8537 (N_8537,N_2471,N_1401);
nor U8538 (N_8538,N_4893,N_4412);
nor U8539 (N_8539,N_1867,N_4123);
nor U8540 (N_8540,N_3782,N_2445);
nor U8541 (N_8541,N_1265,N_1369);
nor U8542 (N_8542,N_785,N_3025);
and U8543 (N_8543,N_3819,N_3469);
or U8544 (N_8544,N_1184,N_3065);
nor U8545 (N_8545,N_3217,N_1742);
or U8546 (N_8546,N_3346,N_3401);
or U8547 (N_8547,N_751,N_2177);
or U8548 (N_8548,N_4619,N_1121);
or U8549 (N_8549,N_2414,N_3554);
or U8550 (N_8550,N_4772,N_4846);
and U8551 (N_8551,N_918,N_4577);
nand U8552 (N_8552,N_4033,N_433);
or U8553 (N_8553,N_2282,N_2263);
or U8554 (N_8554,N_2172,N_1088);
nand U8555 (N_8555,N_358,N_889);
or U8556 (N_8556,N_1202,N_2271);
nor U8557 (N_8557,N_1511,N_2387);
or U8558 (N_8558,N_4120,N_2430);
and U8559 (N_8559,N_3894,N_4837);
nor U8560 (N_8560,N_2888,N_494);
nand U8561 (N_8561,N_1985,N_482);
or U8562 (N_8562,N_1933,N_2896);
or U8563 (N_8563,N_648,N_1841);
and U8564 (N_8564,N_3805,N_346);
nand U8565 (N_8565,N_291,N_4712);
nand U8566 (N_8566,N_1648,N_1183);
nand U8567 (N_8567,N_2695,N_2703);
nand U8568 (N_8568,N_2156,N_3747);
and U8569 (N_8569,N_3922,N_3810);
nor U8570 (N_8570,N_2486,N_316);
or U8571 (N_8571,N_3808,N_4963);
or U8572 (N_8572,N_4164,N_3086);
nand U8573 (N_8573,N_4348,N_920);
or U8574 (N_8574,N_111,N_889);
nor U8575 (N_8575,N_3184,N_3864);
and U8576 (N_8576,N_1172,N_329);
and U8577 (N_8577,N_1502,N_2557);
nand U8578 (N_8578,N_2206,N_1330);
or U8579 (N_8579,N_1929,N_2771);
nand U8580 (N_8580,N_3766,N_1084);
nand U8581 (N_8581,N_2830,N_3656);
or U8582 (N_8582,N_2949,N_3105);
nand U8583 (N_8583,N_1244,N_1579);
or U8584 (N_8584,N_2307,N_3185);
and U8585 (N_8585,N_3133,N_163);
or U8586 (N_8586,N_4255,N_407);
nor U8587 (N_8587,N_3574,N_2116);
or U8588 (N_8588,N_3262,N_3886);
nand U8589 (N_8589,N_2098,N_386);
nand U8590 (N_8590,N_1192,N_2554);
and U8591 (N_8591,N_1708,N_1267);
nor U8592 (N_8592,N_510,N_4524);
or U8593 (N_8593,N_521,N_3548);
nor U8594 (N_8594,N_3508,N_1213);
and U8595 (N_8595,N_3159,N_3501);
nor U8596 (N_8596,N_4470,N_1925);
or U8597 (N_8597,N_4373,N_4807);
or U8598 (N_8598,N_3969,N_1702);
or U8599 (N_8599,N_36,N_2027);
nand U8600 (N_8600,N_1738,N_2039);
or U8601 (N_8601,N_231,N_4053);
and U8602 (N_8602,N_3212,N_609);
and U8603 (N_8603,N_2074,N_1571);
xnor U8604 (N_8604,N_2219,N_3587);
or U8605 (N_8605,N_1886,N_795);
or U8606 (N_8606,N_4227,N_892);
or U8607 (N_8607,N_2596,N_3192);
and U8608 (N_8608,N_3256,N_703);
nor U8609 (N_8609,N_1653,N_23);
or U8610 (N_8610,N_4752,N_3770);
nand U8611 (N_8611,N_453,N_4372);
or U8612 (N_8612,N_1691,N_1939);
nand U8613 (N_8613,N_1388,N_3917);
nand U8614 (N_8614,N_4825,N_4816);
or U8615 (N_8615,N_3859,N_4548);
or U8616 (N_8616,N_51,N_2212);
and U8617 (N_8617,N_1320,N_2012);
and U8618 (N_8618,N_4084,N_3930);
nand U8619 (N_8619,N_2979,N_2466);
and U8620 (N_8620,N_653,N_2433);
or U8621 (N_8621,N_3008,N_342);
or U8622 (N_8622,N_1006,N_2352);
nor U8623 (N_8623,N_4507,N_2870);
and U8624 (N_8624,N_807,N_1192);
and U8625 (N_8625,N_1916,N_4466);
nand U8626 (N_8626,N_4424,N_2349);
and U8627 (N_8627,N_2562,N_3874);
nor U8628 (N_8628,N_4232,N_3695);
nor U8629 (N_8629,N_3928,N_3749);
and U8630 (N_8630,N_4281,N_138);
and U8631 (N_8631,N_2098,N_3328);
or U8632 (N_8632,N_4757,N_1805);
nor U8633 (N_8633,N_1349,N_1652);
nor U8634 (N_8634,N_3881,N_284);
nor U8635 (N_8635,N_1935,N_3872);
or U8636 (N_8636,N_653,N_3939);
nor U8637 (N_8637,N_3689,N_4051);
or U8638 (N_8638,N_2533,N_1898);
nor U8639 (N_8639,N_4245,N_314);
and U8640 (N_8640,N_1116,N_3666);
or U8641 (N_8641,N_4975,N_1658);
nor U8642 (N_8642,N_2121,N_3322);
nor U8643 (N_8643,N_689,N_1863);
and U8644 (N_8644,N_4696,N_3415);
nor U8645 (N_8645,N_460,N_3897);
nand U8646 (N_8646,N_389,N_3347);
and U8647 (N_8647,N_2526,N_655);
and U8648 (N_8648,N_600,N_4592);
xnor U8649 (N_8649,N_4843,N_555);
or U8650 (N_8650,N_677,N_402);
nor U8651 (N_8651,N_4044,N_3855);
nand U8652 (N_8652,N_3575,N_3847);
or U8653 (N_8653,N_1133,N_2065);
or U8654 (N_8654,N_2144,N_4271);
or U8655 (N_8655,N_3721,N_230);
or U8656 (N_8656,N_3635,N_2511);
xor U8657 (N_8657,N_2647,N_1132);
nor U8658 (N_8658,N_2060,N_2539);
xor U8659 (N_8659,N_1676,N_2728);
and U8660 (N_8660,N_1011,N_4624);
and U8661 (N_8661,N_65,N_3550);
nand U8662 (N_8662,N_2847,N_4309);
and U8663 (N_8663,N_35,N_4198);
and U8664 (N_8664,N_2270,N_4945);
xor U8665 (N_8665,N_1796,N_3415);
or U8666 (N_8666,N_2066,N_1041);
and U8667 (N_8667,N_2962,N_964);
and U8668 (N_8668,N_4190,N_857);
and U8669 (N_8669,N_3739,N_3450);
nor U8670 (N_8670,N_3516,N_4888);
nand U8671 (N_8671,N_1703,N_4518);
or U8672 (N_8672,N_1056,N_402);
nor U8673 (N_8673,N_2831,N_901);
nor U8674 (N_8674,N_4143,N_4169);
nand U8675 (N_8675,N_17,N_1125);
and U8676 (N_8676,N_1548,N_722);
nand U8677 (N_8677,N_501,N_3955);
nand U8678 (N_8678,N_2444,N_3448);
and U8679 (N_8679,N_2094,N_4894);
nand U8680 (N_8680,N_4429,N_560);
or U8681 (N_8681,N_3222,N_2333);
and U8682 (N_8682,N_4418,N_4864);
nand U8683 (N_8683,N_2141,N_3352);
nand U8684 (N_8684,N_4406,N_2840);
xnor U8685 (N_8685,N_4834,N_2728);
or U8686 (N_8686,N_4637,N_1476);
and U8687 (N_8687,N_841,N_4229);
and U8688 (N_8688,N_2968,N_1834);
nor U8689 (N_8689,N_2237,N_4670);
nor U8690 (N_8690,N_4798,N_4177);
or U8691 (N_8691,N_167,N_4633);
nand U8692 (N_8692,N_3527,N_1790);
or U8693 (N_8693,N_1851,N_1535);
and U8694 (N_8694,N_2585,N_820);
nand U8695 (N_8695,N_3098,N_732);
and U8696 (N_8696,N_4797,N_1646);
or U8697 (N_8697,N_682,N_2753);
or U8698 (N_8698,N_2619,N_4783);
nand U8699 (N_8699,N_960,N_1697);
nor U8700 (N_8700,N_3501,N_2733);
and U8701 (N_8701,N_3253,N_1211);
and U8702 (N_8702,N_4105,N_3087);
and U8703 (N_8703,N_2567,N_1397);
nand U8704 (N_8704,N_4928,N_648);
nand U8705 (N_8705,N_3805,N_298);
and U8706 (N_8706,N_656,N_562);
nand U8707 (N_8707,N_828,N_4169);
and U8708 (N_8708,N_2468,N_3279);
and U8709 (N_8709,N_3921,N_1175);
or U8710 (N_8710,N_890,N_1887);
nor U8711 (N_8711,N_606,N_2358);
nand U8712 (N_8712,N_4252,N_1606);
nor U8713 (N_8713,N_1900,N_4114);
nor U8714 (N_8714,N_1806,N_913);
and U8715 (N_8715,N_3635,N_1233);
nand U8716 (N_8716,N_3444,N_1093);
xor U8717 (N_8717,N_1849,N_3654);
and U8718 (N_8718,N_4854,N_4902);
nor U8719 (N_8719,N_3537,N_3798);
nor U8720 (N_8720,N_441,N_1000);
and U8721 (N_8721,N_1037,N_4319);
nand U8722 (N_8722,N_2685,N_2061);
nand U8723 (N_8723,N_2237,N_1051);
nor U8724 (N_8724,N_4663,N_1891);
nand U8725 (N_8725,N_1303,N_1522);
or U8726 (N_8726,N_2721,N_3821);
nand U8727 (N_8727,N_2137,N_3381);
or U8728 (N_8728,N_1714,N_2749);
and U8729 (N_8729,N_4706,N_1539);
nor U8730 (N_8730,N_2125,N_2641);
or U8731 (N_8731,N_2518,N_787);
nand U8732 (N_8732,N_1808,N_1338);
or U8733 (N_8733,N_2632,N_3523);
or U8734 (N_8734,N_2210,N_3035);
and U8735 (N_8735,N_1059,N_3457);
and U8736 (N_8736,N_2453,N_4153);
nor U8737 (N_8737,N_655,N_76);
nand U8738 (N_8738,N_4064,N_4308);
or U8739 (N_8739,N_4702,N_3267);
or U8740 (N_8740,N_4269,N_1488);
and U8741 (N_8741,N_4761,N_2191);
or U8742 (N_8742,N_3413,N_1669);
and U8743 (N_8743,N_2876,N_4373);
and U8744 (N_8744,N_2943,N_3462);
nor U8745 (N_8745,N_3259,N_3639);
nor U8746 (N_8746,N_2201,N_2179);
or U8747 (N_8747,N_3821,N_480);
and U8748 (N_8748,N_3903,N_1475);
or U8749 (N_8749,N_3109,N_3265);
nand U8750 (N_8750,N_2487,N_2751);
nand U8751 (N_8751,N_3784,N_2185);
nor U8752 (N_8752,N_865,N_4245);
nand U8753 (N_8753,N_1957,N_752);
and U8754 (N_8754,N_1576,N_3534);
or U8755 (N_8755,N_101,N_3773);
nor U8756 (N_8756,N_4780,N_527);
or U8757 (N_8757,N_1564,N_3162);
nand U8758 (N_8758,N_4058,N_4019);
nor U8759 (N_8759,N_546,N_4991);
or U8760 (N_8760,N_280,N_3156);
or U8761 (N_8761,N_3267,N_3589);
or U8762 (N_8762,N_539,N_4636);
nand U8763 (N_8763,N_389,N_4549);
nand U8764 (N_8764,N_3502,N_3932);
nor U8765 (N_8765,N_4584,N_303);
nand U8766 (N_8766,N_4152,N_733);
nand U8767 (N_8767,N_951,N_2990);
nand U8768 (N_8768,N_2548,N_1179);
nand U8769 (N_8769,N_1387,N_2073);
nor U8770 (N_8770,N_4413,N_2350);
nor U8771 (N_8771,N_2433,N_2964);
nor U8772 (N_8772,N_693,N_3887);
or U8773 (N_8773,N_1426,N_513);
nor U8774 (N_8774,N_1682,N_333);
or U8775 (N_8775,N_1359,N_578);
and U8776 (N_8776,N_3958,N_3477);
or U8777 (N_8777,N_3271,N_4977);
and U8778 (N_8778,N_2557,N_4254);
nor U8779 (N_8779,N_1721,N_1803);
nor U8780 (N_8780,N_1085,N_1649);
nor U8781 (N_8781,N_1040,N_4650);
nor U8782 (N_8782,N_518,N_61);
or U8783 (N_8783,N_1291,N_786);
or U8784 (N_8784,N_1506,N_918);
nand U8785 (N_8785,N_969,N_1053);
and U8786 (N_8786,N_2842,N_2790);
or U8787 (N_8787,N_4888,N_2575);
nand U8788 (N_8788,N_2236,N_4498);
nor U8789 (N_8789,N_2220,N_3181);
or U8790 (N_8790,N_4579,N_4059);
nor U8791 (N_8791,N_991,N_4372);
and U8792 (N_8792,N_3611,N_1887);
nand U8793 (N_8793,N_1122,N_1044);
and U8794 (N_8794,N_533,N_2836);
or U8795 (N_8795,N_3291,N_2378);
nor U8796 (N_8796,N_3643,N_4126);
and U8797 (N_8797,N_2330,N_820);
nand U8798 (N_8798,N_3634,N_259);
or U8799 (N_8799,N_1629,N_3114);
or U8800 (N_8800,N_3315,N_4075);
nor U8801 (N_8801,N_2003,N_1930);
and U8802 (N_8802,N_1705,N_4217);
nand U8803 (N_8803,N_123,N_3785);
nor U8804 (N_8804,N_3546,N_3935);
and U8805 (N_8805,N_3580,N_4907);
nand U8806 (N_8806,N_4772,N_2457);
nor U8807 (N_8807,N_2103,N_1262);
nor U8808 (N_8808,N_465,N_580);
or U8809 (N_8809,N_4398,N_2500);
nand U8810 (N_8810,N_2636,N_4631);
nand U8811 (N_8811,N_861,N_2569);
or U8812 (N_8812,N_2627,N_123);
or U8813 (N_8813,N_3631,N_3022);
or U8814 (N_8814,N_1610,N_2865);
and U8815 (N_8815,N_4137,N_1049);
or U8816 (N_8816,N_4707,N_945);
or U8817 (N_8817,N_3857,N_1326);
or U8818 (N_8818,N_317,N_4248);
nand U8819 (N_8819,N_4853,N_4550);
nor U8820 (N_8820,N_314,N_4073);
and U8821 (N_8821,N_4977,N_4043);
nor U8822 (N_8822,N_3303,N_4254);
or U8823 (N_8823,N_2367,N_1070);
nor U8824 (N_8824,N_1086,N_2193);
xnor U8825 (N_8825,N_1635,N_4361);
or U8826 (N_8826,N_2912,N_1133);
nand U8827 (N_8827,N_1414,N_4034);
and U8828 (N_8828,N_4868,N_2466);
nor U8829 (N_8829,N_99,N_906);
nand U8830 (N_8830,N_4554,N_4960);
nor U8831 (N_8831,N_760,N_3925);
or U8832 (N_8832,N_1774,N_2978);
nand U8833 (N_8833,N_2667,N_2229);
and U8834 (N_8834,N_1996,N_4796);
or U8835 (N_8835,N_859,N_2583);
or U8836 (N_8836,N_2128,N_196);
and U8837 (N_8837,N_4087,N_3568);
nand U8838 (N_8838,N_5,N_4816);
nor U8839 (N_8839,N_534,N_17);
or U8840 (N_8840,N_2820,N_208);
xor U8841 (N_8841,N_2718,N_1263);
or U8842 (N_8842,N_1118,N_3062);
nand U8843 (N_8843,N_4611,N_1505);
or U8844 (N_8844,N_429,N_2981);
nor U8845 (N_8845,N_1393,N_2380);
nor U8846 (N_8846,N_2585,N_489);
and U8847 (N_8847,N_3362,N_4698);
or U8848 (N_8848,N_4997,N_2627);
nand U8849 (N_8849,N_2164,N_2029);
or U8850 (N_8850,N_1928,N_4775);
and U8851 (N_8851,N_538,N_1833);
nand U8852 (N_8852,N_4289,N_698);
nor U8853 (N_8853,N_3736,N_1930);
nand U8854 (N_8854,N_1684,N_3402);
nor U8855 (N_8855,N_1384,N_309);
nand U8856 (N_8856,N_72,N_4045);
or U8857 (N_8857,N_1302,N_1063);
nand U8858 (N_8858,N_355,N_3911);
nor U8859 (N_8859,N_2506,N_3567);
nand U8860 (N_8860,N_1758,N_3226);
nand U8861 (N_8861,N_1983,N_936);
nor U8862 (N_8862,N_3247,N_4309);
nand U8863 (N_8863,N_2621,N_4996);
nand U8864 (N_8864,N_1842,N_4959);
or U8865 (N_8865,N_4698,N_963);
and U8866 (N_8866,N_359,N_4372);
nand U8867 (N_8867,N_3817,N_3203);
or U8868 (N_8868,N_14,N_3326);
and U8869 (N_8869,N_4475,N_245);
and U8870 (N_8870,N_3775,N_4825);
and U8871 (N_8871,N_2299,N_2874);
nand U8872 (N_8872,N_1976,N_2174);
nand U8873 (N_8873,N_367,N_2102);
and U8874 (N_8874,N_660,N_3517);
nand U8875 (N_8875,N_4015,N_1265);
nand U8876 (N_8876,N_1246,N_2675);
nand U8877 (N_8877,N_3149,N_738);
nor U8878 (N_8878,N_4447,N_2697);
nor U8879 (N_8879,N_321,N_3762);
nor U8880 (N_8880,N_1605,N_1317);
nand U8881 (N_8881,N_2780,N_2628);
nor U8882 (N_8882,N_4099,N_797);
or U8883 (N_8883,N_4259,N_445);
and U8884 (N_8884,N_3221,N_1102);
and U8885 (N_8885,N_3946,N_4490);
and U8886 (N_8886,N_1349,N_3385);
or U8887 (N_8887,N_3556,N_1900);
or U8888 (N_8888,N_3415,N_944);
nand U8889 (N_8889,N_716,N_4397);
and U8890 (N_8890,N_4044,N_1083);
and U8891 (N_8891,N_3058,N_2887);
or U8892 (N_8892,N_3123,N_377);
nand U8893 (N_8893,N_1618,N_4155);
nor U8894 (N_8894,N_4314,N_356);
or U8895 (N_8895,N_589,N_1224);
nor U8896 (N_8896,N_1049,N_2874);
and U8897 (N_8897,N_714,N_2476);
or U8898 (N_8898,N_3461,N_629);
nor U8899 (N_8899,N_881,N_2386);
nand U8900 (N_8900,N_2042,N_904);
or U8901 (N_8901,N_2407,N_451);
nand U8902 (N_8902,N_3515,N_3983);
nor U8903 (N_8903,N_2144,N_2801);
or U8904 (N_8904,N_3795,N_2384);
and U8905 (N_8905,N_1589,N_1386);
nor U8906 (N_8906,N_1460,N_2210);
nand U8907 (N_8907,N_1449,N_650);
nand U8908 (N_8908,N_1685,N_3884);
nand U8909 (N_8909,N_718,N_2318);
and U8910 (N_8910,N_3237,N_3061);
or U8911 (N_8911,N_3501,N_4729);
nor U8912 (N_8912,N_1798,N_2405);
or U8913 (N_8913,N_420,N_674);
nand U8914 (N_8914,N_2893,N_1461);
or U8915 (N_8915,N_2401,N_1578);
nor U8916 (N_8916,N_1060,N_605);
nand U8917 (N_8917,N_274,N_3406);
and U8918 (N_8918,N_3220,N_3260);
nand U8919 (N_8919,N_1009,N_739);
and U8920 (N_8920,N_227,N_1622);
and U8921 (N_8921,N_2128,N_2898);
or U8922 (N_8922,N_4099,N_1869);
nand U8923 (N_8923,N_1704,N_3422);
nor U8924 (N_8924,N_1958,N_1134);
nand U8925 (N_8925,N_3288,N_3470);
nand U8926 (N_8926,N_2520,N_4041);
and U8927 (N_8927,N_1210,N_2358);
nand U8928 (N_8928,N_3191,N_3905);
nor U8929 (N_8929,N_3699,N_3);
nor U8930 (N_8930,N_3675,N_4288);
nand U8931 (N_8931,N_3280,N_644);
nor U8932 (N_8932,N_4422,N_965);
and U8933 (N_8933,N_2360,N_3967);
nor U8934 (N_8934,N_2787,N_4808);
nor U8935 (N_8935,N_2771,N_304);
or U8936 (N_8936,N_1644,N_2543);
nand U8937 (N_8937,N_2832,N_1786);
nor U8938 (N_8938,N_3258,N_1336);
and U8939 (N_8939,N_4468,N_1732);
and U8940 (N_8940,N_4160,N_145);
and U8941 (N_8941,N_3589,N_1052);
nor U8942 (N_8942,N_1989,N_1687);
nor U8943 (N_8943,N_1638,N_3373);
and U8944 (N_8944,N_3433,N_797);
nor U8945 (N_8945,N_4192,N_1860);
or U8946 (N_8946,N_4652,N_2553);
nor U8947 (N_8947,N_2918,N_4753);
nand U8948 (N_8948,N_2647,N_3311);
nand U8949 (N_8949,N_2317,N_4657);
nor U8950 (N_8950,N_1570,N_2980);
nor U8951 (N_8951,N_4178,N_1917);
nand U8952 (N_8952,N_2559,N_716);
or U8953 (N_8953,N_2278,N_124);
or U8954 (N_8954,N_3777,N_3399);
nand U8955 (N_8955,N_986,N_142);
nand U8956 (N_8956,N_110,N_1253);
or U8957 (N_8957,N_3484,N_3884);
or U8958 (N_8958,N_3892,N_3116);
or U8959 (N_8959,N_2907,N_424);
and U8960 (N_8960,N_4244,N_2975);
or U8961 (N_8961,N_3302,N_4538);
and U8962 (N_8962,N_3174,N_2556);
and U8963 (N_8963,N_2158,N_710);
nor U8964 (N_8964,N_3689,N_1693);
and U8965 (N_8965,N_4569,N_900);
or U8966 (N_8966,N_4150,N_583);
or U8967 (N_8967,N_3458,N_1297);
nand U8968 (N_8968,N_1430,N_1299);
or U8969 (N_8969,N_3822,N_3753);
or U8970 (N_8970,N_1380,N_3421);
nand U8971 (N_8971,N_583,N_3538);
or U8972 (N_8972,N_1084,N_4944);
nor U8973 (N_8973,N_3878,N_2929);
nand U8974 (N_8974,N_2684,N_3280);
nand U8975 (N_8975,N_1141,N_3118);
and U8976 (N_8976,N_2746,N_4410);
nand U8977 (N_8977,N_4194,N_1296);
and U8978 (N_8978,N_2455,N_444);
and U8979 (N_8979,N_268,N_2148);
nand U8980 (N_8980,N_2188,N_3877);
and U8981 (N_8981,N_3891,N_997);
nand U8982 (N_8982,N_3594,N_4204);
nand U8983 (N_8983,N_985,N_2944);
nor U8984 (N_8984,N_3751,N_4437);
nand U8985 (N_8985,N_629,N_4996);
nand U8986 (N_8986,N_3371,N_3400);
and U8987 (N_8987,N_2546,N_560);
or U8988 (N_8988,N_2199,N_2557);
and U8989 (N_8989,N_2644,N_4521);
or U8990 (N_8990,N_1432,N_1696);
nor U8991 (N_8991,N_2835,N_2689);
nor U8992 (N_8992,N_3801,N_4463);
nor U8993 (N_8993,N_4403,N_4524);
and U8994 (N_8994,N_3717,N_931);
nor U8995 (N_8995,N_4706,N_1401);
nor U8996 (N_8996,N_4371,N_4715);
nor U8997 (N_8997,N_1199,N_1681);
nor U8998 (N_8998,N_912,N_3024);
nor U8999 (N_8999,N_3223,N_4013);
nor U9000 (N_9000,N_509,N_2281);
or U9001 (N_9001,N_509,N_4652);
and U9002 (N_9002,N_1821,N_3450);
and U9003 (N_9003,N_4720,N_1293);
nand U9004 (N_9004,N_3856,N_3806);
nand U9005 (N_9005,N_4897,N_3399);
or U9006 (N_9006,N_4049,N_1903);
or U9007 (N_9007,N_2420,N_278);
nand U9008 (N_9008,N_4450,N_1583);
nand U9009 (N_9009,N_2534,N_1664);
or U9010 (N_9010,N_215,N_2883);
and U9011 (N_9011,N_4218,N_1529);
nor U9012 (N_9012,N_1065,N_4039);
nand U9013 (N_9013,N_81,N_3551);
nor U9014 (N_9014,N_2037,N_3307);
and U9015 (N_9015,N_116,N_1218);
and U9016 (N_9016,N_1937,N_3273);
nor U9017 (N_9017,N_1365,N_466);
and U9018 (N_9018,N_1555,N_1315);
and U9019 (N_9019,N_1343,N_2694);
xor U9020 (N_9020,N_3046,N_4684);
nor U9021 (N_9021,N_4820,N_1521);
and U9022 (N_9022,N_948,N_582);
and U9023 (N_9023,N_2517,N_4584);
nor U9024 (N_9024,N_1324,N_4668);
nand U9025 (N_9025,N_505,N_62);
or U9026 (N_9026,N_4592,N_137);
and U9027 (N_9027,N_3711,N_4708);
nor U9028 (N_9028,N_4541,N_1836);
and U9029 (N_9029,N_3096,N_2146);
nor U9030 (N_9030,N_3974,N_1355);
and U9031 (N_9031,N_2899,N_4999);
nand U9032 (N_9032,N_3815,N_4403);
nor U9033 (N_9033,N_1610,N_77);
nand U9034 (N_9034,N_1392,N_3279);
nand U9035 (N_9035,N_4106,N_2848);
and U9036 (N_9036,N_1810,N_617);
nand U9037 (N_9037,N_29,N_1757);
or U9038 (N_9038,N_34,N_3044);
or U9039 (N_9039,N_2084,N_1462);
nand U9040 (N_9040,N_893,N_2321);
or U9041 (N_9041,N_2969,N_1851);
nand U9042 (N_9042,N_1423,N_2579);
or U9043 (N_9043,N_2742,N_1619);
and U9044 (N_9044,N_612,N_3676);
nand U9045 (N_9045,N_4877,N_2388);
and U9046 (N_9046,N_3312,N_3859);
nand U9047 (N_9047,N_326,N_1245);
nor U9048 (N_9048,N_2816,N_2283);
nor U9049 (N_9049,N_3445,N_3636);
and U9050 (N_9050,N_3111,N_2107);
nor U9051 (N_9051,N_387,N_1610);
nand U9052 (N_9052,N_4680,N_2535);
nand U9053 (N_9053,N_4103,N_1181);
nor U9054 (N_9054,N_345,N_4875);
or U9055 (N_9055,N_1875,N_2265);
and U9056 (N_9056,N_3098,N_1605);
and U9057 (N_9057,N_1566,N_1903);
nand U9058 (N_9058,N_4721,N_615);
and U9059 (N_9059,N_3539,N_3447);
nor U9060 (N_9060,N_2560,N_2002);
nor U9061 (N_9061,N_1401,N_1843);
nor U9062 (N_9062,N_2714,N_1185);
nand U9063 (N_9063,N_1468,N_2107);
nor U9064 (N_9064,N_800,N_774);
and U9065 (N_9065,N_1476,N_3024);
and U9066 (N_9066,N_4714,N_4792);
nand U9067 (N_9067,N_3696,N_537);
nor U9068 (N_9068,N_2645,N_3565);
or U9069 (N_9069,N_2798,N_1217);
nor U9070 (N_9070,N_3803,N_994);
or U9071 (N_9071,N_2897,N_2143);
nor U9072 (N_9072,N_1617,N_1131);
and U9073 (N_9073,N_3538,N_2105);
and U9074 (N_9074,N_4612,N_2121);
nor U9075 (N_9075,N_4555,N_1108);
nor U9076 (N_9076,N_132,N_1642);
or U9077 (N_9077,N_3262,N_4373);
and U9078 (N_9078,N_2431,N_4484);
nand U9079 (N_9079,N_4588,N_1727);
or U9080 (N_9080,N_2030,N_3134);
or U9081 (N_9081,N_803,N_728);
or U9082 (N_9082,N_1334,N_4249);
and U9083 (N_9083,N_4383,N_483);
nor U9084 (N_9084,N_3793,N_4144);
or U9085 (N_9085,N_1922,N_2312);
nand U9086 (N_9086,N_4268,N_1426);
nor U9087 (N_9087,N_3682,N_4297);
nand U9088 (N_9088,N_2166,N_559);
nor U9089 (N_9089,N_1372,N_3688);
nor U9090 (N_9090,N_4804,N_2313);
or U9091 (N_9091,N_300,N_183);
nor U9092 (N_9092,N_1454,N_1940);
and U9093 (N_9093,N_1738,N_4254);
nor U9094 (N_9094,N_1338,N_4958);
nand U9095 (N_9095,N_1759,N_3018);
or U9096 (N_9096,N_1431,N_4773);
or U9097 (N_9097,N_4518,N_491);
or U9098 (N_9098,N_1051,N_3622);
nor U9099 (N_9099,N_1967,N_1327);
nand U9100 (N_9100,N_1145,N_288);
or U9101 (N_9101,N_4397,N_4459);
nand U9102 (N_9102,N_1006,N_816);
nand U9103 (N_9103,N_3095,N_2909);
nand U9104 (N_9104,N_4128,N_289);
or U9105 (N_9105,N_2759,N_2735);
and U9106 (N_9106,N_2728,N_108);
nor U9107 (N_9107,N_4770,N_4011);
and U9108 (N_9108,N_753,N_2774);
nor U9109 (N_9109,N_3253,N_4993);
nand U9110 (N_9110,N_2331,N_2737);
or U9111 (N_9111,N_4555,N_4605);
nand U9112 (N_9112,N_2486,N_4304);
and U9113 (N_9113,N_633,N_384);
nor U9114 (N_9114,N_2782,N_4199);
or U9115 (N_9115,N_1001,N_4066);
and U9116 (N_9116,N_3533,N_3746);
or U9117 (N_9117,N_2898,N_1122);
and U9118 (N_9118,N_2319,N_926);
nand U9119 (N_9119,N_1843,N_1275);
nor U9120 (N_9120,N_1393,N_3547);
or U9121 (N_9121,N_2221,N_86);
or U9122 (N_9122,N_1291,N_496);
nor U9123 (N_9123,N_1152,N_2843);
or U9124 (N_9124,N_2091,N_1767);
nor U9125 (N_9125,N_4990,N_455);
nor U9126 (N_9126,N_2219,N_595);
or U9127 (N_9127,N_3687,N_4794);
or U9128 (N_9128,N_4246,N_4602);
and U9129 (N_9129,N_1686,N_1693);
nand U9130 (N_9130,N_4532,N_324);
or U9131 (N_9131,N_4110,N_820);
and U9132 (N_9132,N_2242,N_4510);
or U9133 (N_9133,N_2854,N_363);
nand U9134 (N_9134,N_945,N_4749);
or U9135 (N_9135,N_2293,N_3824);
or U9136 (N_9136,N_2441,N_4884);
nand U9137 (N_9137,N_839,N_1201);
nand U9138 (N_9138,N_2937,N_194);
and U9139 (N_9139,N_3953,N_2855);
and U9140 (N_9140,N_127,N_4043);
and U9141 (N_9141,N_3087,N_1437);
or U9142 (N_9142,N_1304,N_383);
or U9143 (N_9143,N_3439,N_837);
nand U9144 (N_9144,N_561,N_4418);
nor U9145 (N_9145,N_2189,N_3717);
nor U9146 (N_9146,N_3948,N_2566);
and U9147 (N_9147,N_2306,N_293);
and U9148 (N_9148,N_2341,N_1482);
nor U9149 (N_9149,N_1702,N_4484);
nor U9150 (N_9150,N_1482,N_1249);
or U9151 (N_9151,N_4303,N_1191);
or U9152 (N_9152,N_1703,N_676);
nand U9153 (N_9153,N_3846,N_3223);
nor U9154 (N_9154,N_1521,N_4061);
nor U9155 (N_9155,N_3822,N_1984);
and U9156 (N_9156,N_2344,N_744);
nor U9157 (N_9157,N_1512,N_710);
and U9158 (N_9158,N_468,N_3738);
and U9159 (N_9159,N_696,N_1362);
nor U9160 (N_9160,N_2055,N_3851);
nor U9161 (N_9161,N_640,N_4684);
and U9162 (N_9162,N_2683,N_2096);
nor U9163 (N_9163,N_3827,N_1465);
or U9164 (N_9164,N_2847,N_4967);
or U9165 (N_9165,N_4091,N_361);
or U9166 (N_9166,N_1031,N_3886);
nor U9167 (N_9167,N_2515,N_1393);
or U9168 (N_9168,N_4845,N_1904);
nor U9169 (N_9169,N_1114,N_3926);
nand U9170 (N_9170,N_1243,N_352);
and U9171 (N_9171,N_553,N_433);
or U9172 (N_9172,N_463,N_2372);
and U9173 (N_9173,N_84,N_2276);
and U9174 (N_9174,N_211,N_1558);
and U9175 (N_9175,N_3047,N_2069);
and U9176 (N_9176,N_864,N_2054);
or U9177 (N_9177,N_3892,N_974);
and U9178 (N_9178,N_381,N_4470);
or U9179 (N_9179,N_3151,N_4975);
nand U9180 (N_9180,N_1710,N_4581);
nand U9181 (N_9181,N_432,N_3493);
and U9182 (N_9182,N_2951,N_2709);
nor U9183 (N_9183,N_3262,N_63);
xnor U9184 (N_9184,N_961,N_1910);
nor U9185 (N_9185,N_2968,N_2114);
nand U9186 (N_9186,N_3535,N_4894);
or U9187 (N_9187,N_3889,N_2600);
nand U9188 (N_9188,N_2832,N_2823);
and U9189 (N_9189,N_627,N_2136);
nand U9190 (N_9190,N_631,N_1999);
or U9191 (N_9191,N_443,N_638);
nor U9192 (N_9192,N_2155,N_3554);
or U9193 (N_9193,N_2629,N_3178);
or U9194 (N_9194,N_2898,N_1161);
nor U9195 (N_9195,N_4132,N_2029);
nor U9196 (N_9196,N_666,N_4746);
nand U9197 (N_9197,N_2424,N_3694);
nand U9198 (N_9198,N_4296,N_1490);
or U9199 (N_9199,N_3166,N_541);
nand U9200 (N_9200,N_3838,N_4913);
nand U9201 (N_9201,N_4950,N_2893);
nor U9202 (N_9202,N_647,N_4596);
and U9203 (N_9203,N_4480,N_3643);
nand U9204 (N_9204,N_1691,N_4016);
nor U9205 (N_9205,N_1544,N_2236);
and U9206 (N_9206,N_2448,N_1523);
nor U9207 (N_9207,N_1838,N_314);
nor U9208 (N_9208,N_2672,N_3928);
nor U9209 (N_9209,N_1020,N_4593);
nand U9210 (N_9210,N_4311,N_4220);
nand U9211 (N_9211,N_1714,N_4715);
and U9212 (N_9212,N_3621,N_1542);
or U9213 (N_9213,N_4685,N_2093);
nor U9214 (N_9214,N_4450,N_1007);
nand U9215 (N_9215,N_1464,N_4712);
nor U9216 (N_9216,N_1695,N_3149);
and U9217 (N_9217,N_1002,N_3946);
nand U9218 (N_9218,N_2258,N_3490);
nand U9219 (N_9219,N_3379,N_802);
nand U9220 (N_9220,N_3133,N_1117);
or U9221 (N_9221,N_3971,N_4225);
nor U9222 (N_9222,N_4056,N_379);
nor U9223 (N_9223,N_3314,N_2215);
nand U9224 (N_9224,N_4446,N_3626);
nand U9225 (N_9225,N_1041,N_3094);
nand U9226 (N_9226,N_1937,N_4730);
nor U9227 (N_9227,N_2542,N_3991);
and U9228 (N_9228,N_2874,N_3937);
and U9229 (N_9229,N_3687,N_4270);
nor U9230 (N_9230,N_3903,N_1877);
nor U9231 (N_9231,N_3224,N_2325);
nand U9232 (N_9232,N_2520,N_1963);
nor U9233 (N_9233,N_1147,N_323);
nor U9234 (N_9234,N_2432,N_2554);
and U9235 (N_9235,N_2924,N_4722);
or U9236 (N_9236,N_2707,N_4972);
nand U9237 (N_9237,N_877,N_2261);
or U9238 (N_9238,N_3056,N_3280);
or U9239 (N_9239,N_4625,N_4563);
or U9240 (N_9240,N_3668,N_3106);
and U9241 (N_9241,N_1508,N_4698);
or U9242 (N_9242,N_79,N_3343);
nor U9243 (N_9243,N_403,N_3505);
and U9244 (N_9244,N_3882,N_2949);
nand U9245 (N_9245,N_3470,N_1411);
nand U9246 (N_9246,N_2784,N_1709);
nand U9247 (N_9247,N_4127,N_4935);
and U9248 (N_9248,N_4638,N_2040);
or U9249 (N_9249,N_4838,N_4913);
nor U9250 (N_9250,N_1781,N_2299);
nand U9251 (N_9251,N_55,N_3174);
and U9252 (N_9252,N_3516,N_1351);
nand U9253 (N_9253,N_760,N_3817);
and U9254 (N_9254,N_4551,N_4604);
nand U9255 (N_9255,N_3800,N_4083);
nand U9256 (N_9256,N_2430,N_63);
or U9257 (N_9257,N_4053,N_4725);
and U9258 (N_9258,N_4661,N_117);
and U9259 (N_9259,N_4658,N_40);
and U9260 (N_9260,N_2552,N_4677);
and U9261 (N_9261,N_3932,N_4834);
or U9262 (N_9262,N_2948,N_4512);
and U9263 (N_9263,N_422,N_3015);
and U9264 (N_9264,N_1861,N_3256);
nand U9265 (N_9265,N_944,N_1354);
and U9266 (N_9266,N_2434,N_4971);
or U9267 (N_9267,N_3147,N_261);
nand U9268 (N_9268,N_1348,N_3902);
and U9269 (N_9269,N_3020,N_2761);
nor U9270 (N_9270,N_2452,N_956);
and U9271 (N_9271,N_3946,N_881);
nand U9272 (N_9272,N_481,N_2548);
nand U9273 (N_9273,N_4603,N_4439);
or U9274 (N_9274,N_4138,N_305);
xor U9275 (N_9275,N_2476,N_1360);
or U9276 (N_9276,N_4817,N_2123);
xnor U9277 (N_9277,N_734,N_4979);
or U9278 (N_9278,N_13,N_3282);
or U9279 (N_9279,N_1885,N_4921);
and U9280 (N_9280,N_3032,N_4551);
nand U9281 (N_9281,N_3773,N_4342);
nand U9282 (N_9282,N_3611,N_4979);
and U9283 (N_9283,N_2188,N_4434);
or U9284 (N_9284,N_4997,N_2386);
nand U9285 (N_9285,N_528,N_3108);
or U9286 (N_9286,N_4224,N_2435);
and U9287 (N_9287,N_4385,N_2);
nand U9288 (N_9288,N_2990,N_6);
or U9289 (N_9289,N_2406,N_4279);
or U9290 (N_9290,N_575,N_3450);
and U9291 (N_9291,N_2041,N_2316);
nand U9292 (N_9292,N_1635,N_284);
nor U9293 (N_9293,N_4972,N_4262);
and U9294 (N_9294,N_132,N_301);
and U9295 (N_9295,N_3045,N_3278);
and U9296 (N_9296,N_4408,N_3224);
nor U9297 (N_9297,N_837,N_2370);
or U9298 (N_9298,N_664,N_4478);
nand U9299 (N_9299,N_306,N_3589);
nand U9300 (N_9300,N_3167,N_1694);
nand U9301 (N_9301,N_3139,N_4055);
or U9302 (N_9302,N_3449,N_1016);
nand U9303 (N_9303,N_4232,N_1668);
or U9304 (N_9304,N_3187,N_1408);
and U9305 (N_9305,N_2830,N_733);
or U9306 (N_9306,N_1991,N_4259);
or U9307 (N_9307,N_639,N_1528);
nand U9308 (N_9308,N_951,N_4325);
xnor U9309 (N_9309,N_585,N_3375);
nor U9310 (N_9310,N_3797,N_3710);
and U9311 (N_9311,N_2183,N_1023);
or U9312 (N_9312,N_2418,N_4716);
nor U9313 (N_9313,N_3357,N_4969);
nor U9314 (N_9314,N_4624,N_2695);
nand U9315 (N_9315,N_1028,N_4007);
or U9316 (N_9316,N_2123,N_3862);
nand U9317 (N_9317,N_779,N_1180);
nor U9318 (N_9318,N_1575,N_4611);
or U9319 (N_9319,N_871,N_3729);
or U9320 (N_9320,N_254,N_67);
nand U9321 (N_9321,N_3000,N_4287);
or U9322 (N_9322,N_4842,N_3366);
and U9323 (N_9323,N_2480,N_1163);
nor U9324 (N_9324,N_3223,N_3181);
nand U9325 (N_9325,N_997,N_2188);
or U9326 (N_9326,N_3902,N_2601);
or U9327 (N_9327,N_2570,N_442);
nand U9328 (N_9328,N_1936,N_1268);
nand U9329 (N_9329,N_800,N_614);
nor U9330 (N_9330,N_3651,N_1883);
or U9331 (N_9331,N_2943,N_1763);
nor U9332 (N_9332,N_500,N_765);
and U9333 (N_9333,N_1139,N_1763);
nor U9334 (N_9334,N_4642,N_1020);
or U9335 (N_9335,N_959,N_514);
or U9336 (N_9336,N_4139,N_1921);
nand U9337 (N_9337,N_3028,N_4583);
or U9338 (N_9338,N_1349,N_1671);
nor U9339 (N_9339,N_4544,N_4879);
or U9340 (N_9340,N_798,N_1783);
nand U9341 (N_9341,N_2867,N_2182);
or U9342 (N_9342,N_3932,N_1440);
or U9343 (N_9343,N_3452,N_2504);
or U9344 (N_9344,N_3930,N_2781);
and U9345 (N_9345,N_2030,N_1401);
and U9346 (N_9346,N_179,N_633);
and U9347 (N_9347,N_1157,N_4726);
and U9348 (N_9348,N_3742,N_251);
and U9349 (N_9349,N_503,N_1958);
or U9350 (N_9350,N_994,N_2271);
or U9351 (N_9351,N_2708,N_1417);
and U9352 (N_9352,N_565,N_1860);
nor U9353 (N_9353,N_11,N_4245);
nand U9354 (N_9354,N_641,N_458);
or U9355 (N_9355,N_3693,N_4081);
xnor U9356 (N_9356,N_894,N_4699);
or U9357 (N_9357,N_3371,N_4487);
or U9358 (N_9358,N_4061,N_2817);
and U9359 (N_9359,N_1623,N_3779);
nand U9360 (N_9360,N_2831,N_1132);
and U9361 (N_9361,N_3193,N_1938);
nor U9362 (N_9362,N_3354,N_2304);
or U9363 (N_9363,N_4617,N_1853);
and U9364 (N_9364,N_2058,N_395);
nor U9365 (N_9365,N_2134,N_3111);
or U9366 (N_9366,N_4809,N_1866);
or U9367 (N_9367,N_3186,N_1204);
or U9368 (N_9368,N_2012,N_1165);
or U9369 (N_9369,N_1759,N_4436);
nand U9370 (N_9370,N_1576,N_2237);
nor U9371 (N_9371,N_3930,N_2180);
or U9372 (N_9372,N_4812,N_4511);
nand U9373 (N_9373,N_2214,N_111);
and U9374 (N_9374,N_2371,N_4091);
nand U9375 (N_9375,N_4093,N_2649);
or U9376 (N_9376,N_3069,N_2608);
and U9377 (N_9377,N_4765,N_526);
and U9378 (N_9378,N_2357,N_4024);
nand U9379 (N_9379,N_554,N_3149);
xor U9380 (N_9380,N_4648,N_1308);
nand U9381 (N_9381,N_3161,N_4697);
or U9382 (N_9382,N_3357,N_1910);
nor U9383 (N_9383,N_1687,N_2725);
or U9384 (N_9384,N_3993,N_3018);
and U9385 (N_9385,N_1772,N_4874);
and U9386 (N_9386,N_2649,N_3163);
nand U9387 (N_9387,N_3779,N_3846);
and U9388 (N_9388,N_4823,N_2263);
or U9389 (N_9389,N_294,N_2468);
and U9390 (N_9390,N_906,N_886);
nor U9391 (N_9391,N_4318,N_4267);
nand U9392 (N_9392,N_300,N_3734);
and U9393 (N_9393,N_1111,N_2836);
nand U9394 (N_9394,N_2185,N_3979);
nor U9395 (N_9395,N_1961,N_4805);
nor U9396 (N_9396,N_2997,N_2926);
nand U9397 (N_9397,N_3340,N_4269);
nor U9398 (N_9398,N_3952,N_3004);
nor U9399 (N_9399,N_1705,N_2160);
or U9400 (N_9400,N_1130,N_2355);
and U9401 (N_9401,N_2805,N_4418);
or U9402 (N_9402,N_4805,N_3162);
nor U9403 (N_9403,N_3509,N_2569);
and U9404 (N_9404,N_3958,N_3003);
nand U9405 (N_9405,N_3578,N_4383);
xor U9406 (N_9406,N_4178,N_752);
or U9407 (N_9407,N_1255,N_24);
and U9408 (N_9408,N_1956,N_142);
xor U9409 (N_9409,N_2395,N_1290);
or U9410 (N_9410,N_2603,N_2546);
nor U9411 (N_9411,N_2544,N_252);
nor U9412 (N_9412,N_1081,N_117);
nand U9413 (N_9413,N_3248,N_94);
nand U9414 (N_9414,N_198,N_2803);
and U9415 (N_9415,N_108,N_1183);
or U9416 (N_9416,N_4747,N_3236);
and U9417 (N_9417,N_1172,N_3261);
and U9418 (N_9418,N_1827,N_2076);
nand U9419 (N_9419,N_410,N_3240);
and U9420 (N_9420,N_2313,N_5);
nor U9421 (N_9421,N_707,N_2697);
or U9422 (N_9422,N_3542,N_941);
nor U9423 (N_9423,N_1506,N_4922);
and U9424 (N_9424,N_1864,N_3077);
nand U9425 (N_9425,N_652,N_740);
nand U9426 (N_9426,N_3017,N_847);
and U9427 (N_9427,N_1956,N_4717);
xor U9428 (N_9428,N_4601,N_3415);
nand U9429 (N_9429,N_1347,N_4716);
and U9430 (N_9430,N_3637,N_3245);
nand U9431 (N_9431,N_526,N_690);
or U9432 (N_9432,N_629,N_3890);
and U9433 (N_9433,N_3896,N_933);
or U9434 (N_9434,N_990,N_165);
nand U9435 (N_9435,N_732,N_3600);
and U9436 (N_9436,N_1739,N_263);
nand U9437 (N_9437,N_120,N_3353);
nor U9438 (N_9438,N_1711,N_4759);
nor U9439 (N_9439,N_1322,N_2236);
nand U9440 (N_9440,N_4320,N_4464);
or U9441 (N_9441,N_4626,N_1841);
nor U9442 (N_9442,N_2855,N_115);
nor U9443 (N_9443,N_2399,N_1213);
and U9444 (N_9444,N_4748,N_2666);
or U9445 (N_9445,N_2064,N_3266);
nor U9446 (N_9446,N_4474,N_1474);
and U9447 (N_9447,N_3957,N_4966);
nor U9448 (N_9448,N_3202,N_0);
nand U9449 (N_9449,N_2688,N_4614);
and U9450 (N_9450,N_349,N_4720);
and U9451 (N_9451,N_3384,N_65);
or U9452 (N_9452,N_2791,N_1063);
nand U9453 (N_9453,N_1331,N_4085);
nand U9454 (N_9454,N_748,N_2635);
nor U9455 (N_9455,N_1426,N_337);
or U9456 (N_9456,N_1498,N_508);
or U9457 (N_9457,N_3375,N_1127);
nor U9458 (N_9458,N_2185,N_3708);
and U9459 (N_9459,N_1720,N_4950);
nand U9460 (N_9460,N_3809,N_1870);
and U9461 (N_9461,N_132,N_2414);
nor U9462 (N_9462,N_4484,N_3301);
nand U9463 (N_9463,N_998,N_3166);
or U9464 (N_9464,N_1683,N_4665);
nand U9465 (N_9465,N_2251,N_2381);
nor U9466 (N_9466,N_1628,N_4309);
or U9467 (N_9467,N_581,N_4875);
and U9468 (N_9468,N_1387,N_647);
or U9469 (N_9469,N_1454,N_1083);
nor U9470 (N_9470,N_1477,N_4198);
nand U9471 (N_9471,N_289,N_4553);
and U9472 (N_9472,N_4921,N_574);
and U9473 (N_9473,N_2346,N_644);
nand U9474 (N_9474,N_3950,N_843);
nor U9475 (N_9475,N_1084,N_4472);
and U9476 (N_9476,N_32,N_514);
or U9477 (N_9477,N_4157,N_810);
nor U9478 (N_9478,N_4735,N_1546);
and U9479 (N_9479,N_2852,N_2636);
nor U9480 (N_9480,N_17,N_242);
nor U9481 (N_9481,N_4241,N_1228);
nor U9482 (N_9482,N_2495,N_3755);
or U9483 (N_9483,N_3002,N_1872);
nor U9484 (N_9484,N_3156,N_2731);
nor U9485 (N_9485,N_1178,N_3007);
and U9486 (N_9486,N_2171,N_3500);
nor U9487 (N_9487,N_1379,N_1107);
or U9488 (N_9488,N_1607,N_2877);
nand U9489 (N_9489,N_817,N_1628);
or U9490 (N_9490,N_4280,N_1246);
and U9491 (N_9491,N_210,N_2559);
nand U9492 (N_9492,N_2947,N_2330);
or U9493 (N_9493,N_3031,N_771);
and U9494 (N_9494,N_612,N_1080);
and U9495 (N_9495,N_479,N_965);
nand U9496 (N_9496,N_52,N_4002);
nor U9497 (N_9497,N_4731,N_4249);
nand U9498 (N_9498,N_981,N_4753);
and U9499 (N_9499,N_509,N_4669);
and U9500 (N_9500,N_3190,N_705);
nand U9501 (N_9501,N_720,N_3220);
or U9502 (N_9502,N_141,N_4204);
nand U9503 (N_9503,N_2143,N_284);
xnor U9504 (N_9504,N_4194,N_4480);
nand U9505 (N_9505,N_3045,N_1855);
nand U9506 (N_9506,N_2676,N_2914);
nor U9507 (N_9507,N_3634,N_4926);
nor U9508 (N_9508,N_3754,N_2604);
or U9509 (N_9509,N_4760,N_538);
or U9510 (N_9510,N_704,N_1459);
nor U9511 (N_9511,N_3148,N_2985);
or U9512 (N_9512,N_3049,N_4466);
or U9513 (N_9513,N_4325,N_1984);
and U9514 (N_9514,N_2877,N_2264);
or U9515 (N_9515,N_2541,N_4724);
or U9516 (N_9516,N_1749,N_2743);
or U9517 (N_9517,N_2414,N_2622);
or U9518 (N_9518,N_3735,N_4149);
xnor U9519 (N_9519,N_4443,N_3191);
nand U9520 (N_9520,N_1442,N_2189);
or U9521 (N_9521,N_1780,N_3008);
or U9522 (N_9522,N_4538,N_3091);
or U9523 (N_9523,N_4890,N_4830);
nand U9524 (N_9524,N_4344,N_811);
nor U9525 (N_9525,N_1907,N_905);
or U9526 (N_9526,N_2301,N_2794);
nand U9527 (N_9527,N_1577,N_38);
nor U9528 (N_9528,N_1646,N_2525);
nor U9529 (N_9529,N_2227,N_4474);
nor U9530 (N_9530,N_4409,N_3770);
nand U9531 (N_9531,N_2091,N_1699);
and U9532 (N_9532,N_3829,N_1590);
or U9533 (N_9533,N_4743,N_1266);
or U9534 (N_9534,N_4192,N_4899);
nor U9535 (N_9535,N_338,N_975);
or U9536 (N_9536,N_1948,N_2384);
or U9537 (N_9537,N_4622,N_1556);
nand U9538 (N_9538,N_2233,N_4493);
and U9539 (N_9539,N_4970,N_2659);
nand U9540 (N_9540,N_2007,N_416);
nor U9541 (N_9541,N_1589,N_4037);
or U9542 (N_9542,N_3917,N_2809);
and U9543 (N_9543,N_3021,N_1803);
nor U9544 (N_9544,N_3549,N_2317);
nand U9545 (N_9545,N_2397,N_454);
and U9546 (N_9546,N_1403,N_1244);
nor U9547 (N_9547,N_3813,N_2034);
or U9548 (N_9548,N_626,N_180);
nand U9549 (N_9549,N_2493,N_1784);
nor U9550 (N_9550,N_3193,N_1913);
and U9551 (N_9551,N_3116,N_2999);
xnor U9552 (N_9552,N_1488,N_392);
or U9553 (N_9553,N_2214,N_1130);
and U9554 (N_9554,N_979,N_614);
nand U9555 (N_9555,N_410,N_4701);
or U9556 (N_9556,N_718,N_2196);
or U9557 (N_9557,N_2584,N_1235);
or U9558 (N_9558,N_3931,N_3563);
or U9559 (N_9559,N_4975,N_2330);
nor U9560 (N_9560,N_445,N_4775);
or U9561 (N_9561,N_485,N_65);
nor U9562 (N_9562,N_2631,N_362);
or U9563 (N_9563,N_3452,N_685);
nand U9564 (N_9564,N_193,N_1723);
nand U9565 (N_9565,N_23,N_2202);
nor U9566 (N_9566,N_3855,N_3149);
or U9567 (N_9567,N_3224,N_4520);
or U9568 (N_9568,N_1738,N_2049);
and U9569 (N_9569,N_1571,N_4014);
or U9570 (N_9570,N_2153,N_4257);
nand U9571 (N_9571,N_2303,N_4292);
or U9572 (N_9572,N_2227,N_2866);
or U9573 (N_9573,N_530,N_1394);
xor U9574 (N_9574,N_2229,N_2581);
nor U9575 (N_9575,N_1401,N_1937);
and U9576 (N_9576,N_1663,N_3617);
or U9577 (N_9577,N_762,N_3076);
nand U9578 (N_9578,N_3069,N_3800);
and U9579 (N_9579,N_64,N_650);
nand U9580 (N_9580,N_1787,N_3888);
nand U9581 (N_9581,N_2040,N_4183);
and U9582 (N_9582,N_2702,N_1500);
and U9583 (N_9583,N_250,N_3586);
nand U9584 (N_9584,N_3281,N_2692);
nand U9585 (N_9585,N_2399,N_1036);
or U9586 (N_9586,N_3246,N_1894);
or U9587 (N_9587,N_3502,N_342);
and U9588 (N_9588,N_3586,N_4792);
nand U9589 (N_9589,N_2097,N_1299);
nor U9590 (N_9590,N_1177,N_1202);
or U9591 (N_9591,N_3470,N_99);
or U9592 (N_9592,N_2207,N_2225);
and U9593 (N_9593,N_4838,N_3636);
nand U9594 (N_9594,N_3484,N_4262);
and U9595 (N_9595,N_480,N_3075);
or U9596 (N_9596,N_1436,N_2573);
xnor U9597 (N_9597,N_2856,N_1485);
and U9598 (N_9598,N_4084,N_1918);
nand U9599 (N_9599,N_3809,N_1261);
nand U9600 (N_9600,N_472,N_2031);
nor U9601 (N_9601,N_2839,N_4949);
or U9602 (N_9602,N_4025,N_275);
or U9603 (N_9603,N_1646,N_1236);
nand U9604 (N_9604,N_619,N_3285);
or U9605 (N_9605,N_1644,N_1646);
nand U9606 (N_9606,N_2353,N_515);
or U9607 (N_9607,N_3129,N_3684);
nand U9608 (N_9608,N_3133,N_2943);
or U9609 (N_9609,N_1846,N_4381);
and U9610 (N_9610,N_4216,N_2256);
nor U9611 (N_9611,N_1422,N_3165);
nor U9612 (N_9612,N_302,N_2058);
nand U9613 (N_9613,N_2536,N_1776);
or U9614 (N_9614,N_1950,N_4122);
nand U9615 (N_9615,N_740,N_4193);
nand U9616 (N_9616,N_2805,N_3413);
nor U9617 (N_9617,N_148,N_3709);
nand U9618 (N_9618,N_822,N_3093);
and U9619 (N_9619,N_4446,N_2738);
or U9620 (N_9620,N_1086,N_850);
or U9621 (N_9621,N_4570,N_3754);
nor U9622 (N_9622,N_1011,N_2793);
and U9623 (N_9623,N_3625,N_2150);
nor U9624 (N_9624,N_1446,N_4747);
and U9625 (N_9625,N_3067,N_1042);
and U9626 (N_9626,N_2907,N_67);
or U9627 (N_9627,N_1090,N_1072);
or U9628 (N_9628,N_4406,N_2441);
or U9629 (N_9629,N_2981,N_4990);
nor U9630 (N_9630,N_3731,N_4557);
and U9631 (N_9631,N_3017,N_3474);
and U9632 (N_9632,N_1519,N_1077);
or U9633 (N_9633,N_4302,N_2141);
nand U9634 (N_9634,N_3077,N_3528);
nand U9635 (N_9635,N_4747,N_3470);
nand U9636 (N_9636,N_1805,N_2015);
nand U9637 (N_9637,N_4693,N_58);
nand U9638 (N_9638,N_1398,N_3620);
and U9639 (N_9639,N_2147,N_3366);
or U9640 (N_9640,N_152,N_4384);
nand U9641 (N_9641,N_3413,N_3353);
or U9642 (N_9642,N_4676,N_1363);
or U9643 (N_9643,N_1600,N_429);
or U9644 (N_9644,N_4469,N_3151);
nand U9645 (N_9645,N_1635,N_275);
nor U9646 (N_9646,N_1201,N_2119);
xnor U9647 (N_9647,N_195,N_4415);
nor U9648 (N_9648,N_1251,N_124);
nand U9649 (N_9649,N_3907,N_3371);
nor U9650 (N_9650,N_2615,N_2282);
or U9651 (N_9651,N_2293,N_2362);
and U9652 (N_9652,N_3932,N_144);
or U9653 (N_9653,N_4672,N_2665);
nor U9654 (N_9654,N_3854,N_3000);
and U9655 (N_9655,N_1466,N_3344);
nand U9656 (N_9656,N_4400,N_1233);
or U9657 (N_9657,N_1486,N_3846);
nand U9658 (N_9658,N_3543,N_3999);
nor U9659 (N_9659,N_1784,N_2961);
or U9660 (N_9660,N_3676,N_3498);
and U9661 (N_9661,N_1038,N_4462);
and U9662 (N_9662,N_4508,N_2998);
and U9663 (N_9663,N_3341,N_4967);
nor U9664 (N_9664,N_3578,N_742);
nand U9665 (N_9665,N_316,N_3103);
nor U9666 (N_9666,N_4232,N_3978);
or U9667 (N_9667,N_307,N_1916);
nand U9668 (N_9668,N_3938,N_278);
nor U9669 (N_9669,N_3221,N_507);
or U9670 (N_9670,N_3029,N_1868);
and U9671 (N_9671,N_1830,N_2020);
nand U9672 (N_9672,N_1855,N_4149);
nand U9673 (N_9673,N_2335,N_2640);
nand U9674 (N_9674,N_2454,N_2204);
nand U9675 (N_9675,N_1642,N_2930);
nor U9676 (N_9676,N_2056,N_1666);
and U9677 (N_9677,N_1125,N_4596);
and U9678 (N_9678,N_2596,N_4187);
nand U9679 (N_9679,N_1419,N_4573);
and U9680 (N_9680,N_2265,N_4265);
nand U9681 (N_9681,N_3700,N_1952);
nand U9682 (N_9682,N_2098,N_731);
nand U9683 (N_9683,N_764,N_1016);
nor U9684 (N_9684,N_3164,N_136);
or U9685 (N_9685,N_3569,N_1392);
nor U9686 (N_9686,N_4010,N_3653);
nor U9687 (N_9687,N_897,N_3829);
nand U9688 (N_9688,N_945,N_3037);
nand U9689 (N_9689,N_268,N_4731);
nor U9690 (N_9690,N_4601,N_2345);
nand U9691 (N_9691,N_2371,N_521);
and U9692 (N_9692,N_3837,N_1543);
xor U9693 (N_9693,N_4255,N_1909);
nor U9694 (N_9694,N_1903,N_1117);
and U9695 (N_9695,N_842,N_2417);
and U9696 (N_9696,N_3639,N_580);
or U9697 (N_9697,N_1807,N_1617);
or U9698 (N_9698,N_4794,N_1193);
nor U9699 (N_9699,N_4569,N_379);
or U9700 (N_9700,N_2138,N_453);
or U9701 (N_9701,N_409,N_2713);
or U9702 (N_9702,N_1481,N_4266);
and U9703 (N_9703,N_2088,N_4997);
and U9704 (N_9704,N_4488,N_1794);
nor U9705 (N_9705,N_2460,N_1700);
or U9706 (N_9706,N_4318,N_4439);
nor U9707 (N_9707,N_2966,N_657);
or U9708 (N_9708,N_4204,N_3776);
nand U9709 (N_9709,N_1994,N_4607);
nor U9710 (N_9710,N_701,N_2142);
and U9711 (N_9711,N_2758,N_3831);
nand U9712 (N_9712,N_683,N_3635);
or U9713 (N_9713,N_4015,N_553);
nand U9714 (N_9714,N_644,N_769);
nor U9715 (N_9715,N_1567,N_3961);
nand U9716 (N_9716,N_1117,N_803);
nor U9717 (N_9717,N_49,N_3819);
or U9718 (N_9718,N_466,N_3971);
nor U9719 (N_9719,N_2578,N_2886);
or U9720 (N_9720,N_1518,N_2465);
and U9721 (N_9721,N_4929,N_3747);
or U9722 (N_9722,N_2223,N_2844);
nor U9723 (N_9723,N_3035,N_2653);
or U9724 (N_9724,N_3873,N_97);
or U9725 (N_9725,N_3321,N_3225);
and U9726 (N_9726,N_1765,N_1399);
nand U9727 (N_9727,N_2761,N_1105);
nor U9728 (N_9728,N_1833,N_392);
and U9729 (N_9729,N_4659,N_585);
and U9730 (N_9730,N_2516,N_3594);
nor U9731 (N_9731,N_4161,N_373);
nor U9732 (N_9732,N_2788,N_205);
and U9733 (N_9733,N_991,N_2268);
nor U9734 (N_9734,N_2342,N_4226);
and U9735 (N_9735,N_1711,N_1013);
nor U9736 (N_9736,N_4469,N_2801);
or U9737 (N_9737,N_1475,N_913);
nor U9738 (N_9738,N_3026,N_328);
nor U9739 (N_9739,N_947,N_1405);
nor U9740 (N_9740,N_3951,N_4598);
nand U9741 (N_9741,N_835,N_2705);
nand U9742 (N_9742,N_1338,N_1509);
and U9743 (N_9743,N_3401,N_1695);
or U9744 (N_9744,N_1614,N_85);
nand U9745 (N_9745,N_4557,N_2777);
nor U9746 (N_9746,N_838,N_4113);
or U9747 (N_9747,N_4557,N_2367);
nand U9748 (N_9748,N_4911,N_1370);
and U9749 (N_9749,N_3554,N_4824);
and U9750 (N_9750,N_2501,N_1345);
nor U9751 (N_9751,N_1908,N_3273);
and U9752 (N_9752,N_3459,N_1943);
nor U9753 (N_9753,N_3768,N_2503);
nor U9754 (N_9754,N_753,N_4456);
nor U9755 (N_9755,N_2952,N_2798);
and U9756 (N_9756,N_829,N_57);
and U9757 (N_9757,N_4255,N_4802);
nor U9758 (N_9758,N_2257,N_3596);
nand U9759 (N_9759,N_2249,N_469);
xnor U9760 (N_9760,N_1402,N_2604);
nand U9761 (N_9761,N_530,N_176);
nand U9762 (N_9762,N_3245,N_276);
and U9763 (N_9763,N_2293,N_3412);
or U9764 (N_9764,N_4958,N_2721);
or U9765 (N_9765,N_1618,N_1194);
and U9766 (N_9766,N_3177,N_2397);
and U9767 (N_9767,N_557,N_1810);
nor U9768 (N_9768,N_1015,N_2816);
nor U9769 (N_9769,N_1859,N_823);
xnor U9770 (N_9770,N_1471,N_1518);
or U9771 (N_9771,N_4318,N_3819);
nor U9772 (N_9772,N_1003,N_4978);
nand U9773 (N_9773,N_2715,N_3382);
and U9774 (N_9774,N_2385,N_1308);
nand U9775 (N_9775,N_1733,N_9);
and U9776 (N_9776,N_3174,N_1356);
and U9777 (N_9777,N_606,N_273);
nor U9778 (N_9778,N_1794,N_2146);
or U9779 (N_9779,N_1735,N_28);
nand U9780 (N_9780,N_3939,N_4557);
or U9781 (N_9781,N_337,N_2237);
nand U9782 (N_9782,N_1483,N_4998);
nor U9783 (N_9783,N_3502,N_1179);
and U9784 (N_9784,N_854,N_2768);
nor U9785 (N_9785,N_4908,N_986);
or U9786 (N_9786,N_837,N_1740);
nand U9787 (N_9787,N_1919,N_3613);
or U9788 (N_9788,N_781,N_4799);
nand U9789 (N_9789,N_4427,N_1660);
and U9790 (N_9790,N_259,N_3588);
or U9791 (N_9791,N_1195,N_3072);
and U9792 (N_9792,N_2114,N_4454);
nor U9793 (N_9793,N_4516,N_1333);
or U9794 (N_9794,N_2552,N_1323);
nand U9795 (N_9795,N_2191,N_4888);
and U9796 (N_9796,N_2749,N_3453);
nand U9797 (N_9797,N_1103,N_1219);
nand U9798 (N_9798,N_3266,N_192);
or U9799 (N_9799,N_4912,N_4695);
and U9800 (N_9800,N_4011,N_262);
or U9801 (N_9801,N_890,N_2990);
and U9802 (N_9802,N_1072,N_2696);
xor U9803 (N_9803,N_3699,N_2823);
nand U9804 (N_9804,N_857,N_904);
or U9805 (N_9805,N_739,N_3642);
nor U9806 (N_9806,N_676,N_32);
nand U9807 (N_9807,N_2313,N_4510);
nand U9808 (N_9808,N_3283,N_1180);
nor U9809 (N_9809,N_3079,N_1625);
nor U9810 (N_9810,N_633,N_4326);
or U9811 (N_9811,N_408,N_1968);
nand U9812 (N_9812,N_4417,N_2490);
and U9813 (N_9813,N_2461,N_1773);
nand U9814 (N_9814,N_247,N_1217);
nor U9815 (N_9815,N_1765,N_1648);
nand U9816 (N_9816,N_4185,N_290);
and U9817 (N_9817,N_3967,N_2929);
or U9818 (N_9818,N_4722,N_1449);
nor U9819 (N_9819,N_3530,N_3646);
nand U9820 (N_9820,N_1550,N_4176);
nor U9821 (N_9821,N_1037,N_4410);
nand U9822 (N_9822,N_1443,N_2963);
and U9823 (N_9823,N_3581,N_3279);
nor U9824 (N_9824,N_477,N_1270);
nor U9825 (N_9825,N_3807,N_4666);
nor U9826 (N_9826,N_3911,N_4584);
nor U9827 (N_9827,N_2805,N_4317);
nand U9828 (N_9828,N_31,N_4891);
or U9829 (N_9829,N_843,N_2954);
and U9830 (N_9830,N_2146,N_3972);
or U9831 (N_9831,N_959,N_4634);
nor U9832 (N_9832,N_818,N_2561);
nor U9833 (N_9833,N_384,N_1336);
nor U9834 (N_9834,N_2824,N_1343);
or U9835 (N_9835,N_224,N_1056);
nor U9836 (N_9836,N_3375,N_1909);
nand U9837 (N_9837,N_4790,N_2506);
nand U9838 (N_9838,N_2509,N_2030);
nand U9839 (N_9839,N_1462,N_2497);
xnor U9840 (N_9840,N_2093,N_304);
or U9841 (N_9841,N_2095,N_385);
or U9842 (N_9842,N_2496,N_4056);
or U9843 (N_9843,N_4364,N_3990);
or U9844 (N_9844,N_3308,N_1259);
nor U9845 (N_9845,N_3296,N_2659);
and U9846 (N_9846,N_2057,N_916);
nor U9847 (N_9847,N_1066,N_2096);
nor U9848 (N_9848,N_3555,N_1977);
nor U9849 (N_9849,N_3429,N_4729);
nand U9850 (N_9850,N_954,N_4237);
and U9851 (N_9851,N_1996,N_1081);
and U9852 (N_9852,N_1246,N_2078);
nand U9853 (N_9853,N_2220,N_4160);
nand U9854 (N_9854,N_3180,N_4833);
and U9855 (N_9855,N_493,N_1058);
or U9856 (N_9856,N_3254,N_1830);
nor U9857 (N_9857,N_3744,N_2479);
or U9858 (N_9858,N_2980,N_4938);
and U9859 (N_9859,N_1932,N_138);
or U9860 (N_9860,N_3925,N_688);
or U9861 (N_9861,N_3140,N_3170);
nand U9862 (N_9862,N_4931,N_4782);
and U9863 (N_9863,N_725,N_2289);
and U9864 (N_9864,N_105,N_3295);
or U9865 (N_9865,N_785,N_1202);
and U9866 (N_9866,N_4917,N_3176);
xnor U9867 (N_9867,N_2588,N_4136);
or U9868 (N_9868,N_658,N_4202);
or U9869 (N_9869,N_2215,N_462);
or U9870 (N_9870,N_3098,N_887);
nand U9871 (N_9871,N_3517,N_867);
or U9872 (N_9872,N_1993,N_4440);
nor U9873 (N_9873,N_2552,N_2208);
and U9874 (N_9874,N_1317,N_418);
nand U9875 (N_9875,N_3169,N_1060);
or U9876 (N_9876,N_540,N_2795);
nor U9877 (N_9877,N_3500,N_678);
and U9878 (N_9878,N_4808,N_4194);
and U9879 (N_9879,N_3860,N_2639);
nor U9880 (N_9880,N_1118,N_2481);
or U9881 (N_9881,N_4789,N_3041);
or U9882 (N_9882,N_4651,N_3588);
or U9883 (N_9883,N_3570,N_2432);
or U9884 (N_9884,N_2497,N_2025);
nand U9885 (N_9885,N_4908,N_934);
or U9886 (N_9886,N_2759,N_4449);
and U9887 (N_9887,N_1508,N_1625);
and U9888 (N_9888,N_2748,N_3874);
nand U9889 (N_9889,N_181,N_2452);
nor U9890 (N_9890,N_2491,N_2208);
and U9891 (N_9891,N_4056,N_4980);
nand U9892 (N_9892,N_3428,N_1644);
nor U9893 (N_9893,N_2260,N_2457);
and U9894 (N_9894,N_4023,N_1124);
and U9895 (N_9895,N_2365,N_4502);
nor U9896 (N_9896,N_3744,N_1382);
and U9897 (N_9897,N_1852,N_533);
or U9898 (N_9898,N_4581,N_3017);
or U9899 (N_9899,N_4748,N_446);
or U9900 (N_9900,N_4345,N_981);
nand U9901 (N_9901,N_349,N_492);
or U9902 (N_9902,N_534,N_4642);
nand U9903 (N_9903,N_3825,N_3912);
or U9904 (N_9904,N_488,N_1654);
or U9905 (N_9905,N_424,N_975);
nand U9906 (N_9906,N_1738,N_2420);
and U9907 (N_9907,N_598,N_2937);
or U9908 (N_9908,N_337,N_1940);
nor U9909 (N_9909,N_4821,N_316);
nor U9910 (N_9910,N_4072,N_3252);
and U9911 (N_9911,N_1889,N_22);
nor U9912 (N_9912,N_2329,N_4680);
xor U9913 (N_9913,N_1802,N_4045);
and U9914 (N_9914,N_4108,N_2827);
or U9915 (N_9915,N_3541,N_3289);
or U9916 (N_9916,N_1897,N_1785);
nand U9917 (N_9917,N_3279,N_1253);
or U9918 (N_9918,N_2010,N_740);
nand U9919 (N_9919,N_296,N_1977);
or U9920 (N_9920,N_756,N_1066);
nor U9921 (N_9921,N_1881,N_3767);
or U9922 (N_9922,N_584,N_1065);
nand U9923 (N_9923,N_3407,N_1671);
nand U9924 (N_9924,N_2557,N_2049);
xor U9925 (N_9925,N_4864,N_141);
and U9926 (N_9926,N_161,N_4788);
or U9927 (N_9927,N_4031,N_1450);
or U9928 (N_9928,N_928,N_1989);
or U9929 (N_9929,N_2292,N_3124);
and U9930 (N_9930,N_3609,N_4332);
nor U9931 (N_9931,N_2245,N_3086);
nor U9932 (N_9932,N_1708,N_126);
nand U9933 (N_9933,N_4850,N_4133);
or U9934 (N_9934,N_4534,N_3800);
nand U9935 (N_9935,N_2280,N_3713);
nor U9936 (N_9936,N_2675,N_3902);
nand U9937 (N_9937,N_1289,N_2615);
and U9938 (N_9938,N_1515,N_3152);
or U9939 (N_9939,N_1340,N_1707);
and U9940 (N_9940,N_153,N_1216);
or U9941 (N_9941,N_3146,N_2115);
nor U9942 (N_9942,N_2509,N_2278);
nor U9943 (N_9943,N_1045,N_1066);
nor U9944 (N_9944,N_4870,N_1068);
nand U9945 (N_9945,N_1668,N_32);
nor U9946 (N_9946,N_4730,N_4647);
nand U9947 (N_9947,N_4709,N_1156);
and U9948 (N_9948,N_629,N_693);
nor U9949 (N_9949,N_2473,N_3364);
nor U9950 (N_9950,N_2540,N_870);
nand U9951 (N_9951,N_2979,N_3854);
or U9952 (N_9952,N_4483,N_14);
nand U9953 (N_9953,N_1544,N_2901);
xnor U9954 (N_9954,N_3922,N_3101);
and U9955 (N_9955,N_3832,N_139);
or U9956 (N_9956,N_1678,N_568);
and U9957 (N_9957,N_214,N_2428);
nor U9958 (N_9958,N_4296,N_3151);
nand U9959 (N_9959,N_4808,N_1009);
nor U9960 (N_9960,N_212,N_1998);
and U9961 (N_9961,N_2501,N_1636);
nor U9962 (N_9962,N_4664,N_4612);
and U9963 (N_9963,N_682,N_1148);
and U9964 (N_9964,N_3887,N_4603);
nor U9965 (N_9965,N_3957,N_3083);
or U9966 (N_9966,N_205,N_1352);
and U9967 (N_9967,N_909,N_1215);
nor U9968 (N_9968,N_2210,N_4486);
or U9969 (N_9969,N_3736,N_758);
or U9970 (N_9970,N_358,N_4085);
nor U9971 (N_9971,N_54,N_3088);
nand U9972 (N_9972,N_2936,N_2812);
or U9973 (N_9973,N_2845,N_2327);
or U9974 (N_9974,N_552,N_569);
nor U9975 (N_9975,N_3560,N_3595);
or U9976 (N_9976,N_278,N_4707);
and U9977 (N_9977,N_1044,N_1582);
and U9978 (N_9978,N_3160,N_2108);
or U9979 (N_9979,N_77,N_302);
nand U9980 (N_9980,N_3247,N_1531);
nand U9981 (N_9981,N_856,N_2115);
and U9982 (N_9982,N_335,N_3863);
or U9983 (N_9983,N_3376,N_3893);
and U9984 (N_9984,N_3595,N_1195);
nand U9985 (N_9985,N_2449,N_3536);
xor U9986 (N_9986,N_549,N_2096);
and U9987 (N_9987,N_189,N_4532);
nand U9988 (N_9988,N_2874,N_116);
nand U9989 (N_9989,N_1706,N_3129);
and U9990 (N_9990,N_2603,N_4477);
nor U9991 (N_9991,N_1434,N_4647);
or U9992 (N_9992,N_518,N_2238);
and U9993 (N_9993,N_2461,N_1495);
or U9994 (N_9994,N_2749,N_3543);
and U9995 (N_9995,N_1618,N_398);
and U9996 (N_9996,N_259,N_3051);
nand U9997 (N_9997,N_1087,N_3447);
or U9998 (N_9998,N_3435,N_996);
nor U9999 (N_9999,N_4154,N_2450);
nand UO_0 (O_0,N_5987,N_5507);
and UO_1 (O_1,N_7576,N_5758);
nor UO_2 (O_2,N_9977,N_9612);
nor UO_3 (O_3,N_7474,N_6077);
or UO_4 (O_4,N_7328,N_8169);
xnor UO_5 (O_5,N_8862,N_6027);
nand UO_6 (O_6,N_5044,N_7982);
nor UO_7 (O_7,N_8780,N_7744);
and UO_8 (O_8,N_7007,N_9691);
and UO_9 (O_9,N_8111,N_9581);
and UO_10 (O_10,N_7588,N_8317);
nand UO_11 (O_11,N_7693,N_9006);
nand UO_12 (O_12,N_8255,N_9451);
or UO_13 (O_13,N_9959,N_5585);
nor UO_14 (O_14,N_9415,N_6231);
xnor UO_15 (O_15,N_7061,N_7227);
nand UO_16 (O_16,N_8783,N_5519);
or UO_17 (O_17,N_6790,N_5254);
nand UO_18 (O_18,N_9738,N_6358);
nor UO_19 (O_19,N_9992,N_7129);
nor UO_20 (O_20,N_5551,N_9608);
and UO_21 (O_21,N_9060,N_8728);
nand UO_22 (O_22,N_5942,N_9828);
or UO_23 (O_23,N_9754,N_5993);
or UO_24 (O_24,N_6101,N_6068);
nor UO_25 (O_25,N_9286,N_9855);
or UO_26 (O_26,N_6079,N_8598);
or UO_27 (O_27,N_9439,N_5946);
nor UO_28 (O_28,N_5653,N_9586);
or UO_29 (O_29,N_7411,N_5672);
and UO_30 (O_30,N_8729,N_9623);
nor UO_31 (O_31,N_6642,N_7049);
nand UO_32 (O_32,N_7393,N_8386);
or UO_33 (O_33,N_8716,N_8515);
nand UO_34 (O_34,N_7368,N_8307);
nand UO_35 (O_35,N_5623,N_9821);
nand UO_36 (O_36,N_6701,N_7500);
and UO_37 (O_37,N_7151,N_6181);
nand UO_38 (O_38,N_7220,N_8252);
or UO_39 (O_39,N_9253,N_5954);
nand UO_40 (O_40,N_6932,N_7910);
nand UO_41 (O_41,N_7923,N_8550);
or UO_42 (O_42,N_8376,N_5194);
nand UO_43 (O_43,N_8482,N_7684);
nor UO_44 (O_44,N_7115,N_9962);
or UO_45 (O_45,N_5515,N_7914);
nor UO_46 (O_46,N_5393,N_8087);
nor UO_47 (O_47,N_7716,N_7184);
nand UO_48 (O_48,N_7330,N_8795);
nor UO_49 (O_49,N_8181,N_8960);
or UO_50 (O_50,N_7252,N_5786);
or UO_51 (O_51,N_6646,N_6756);
nor UO_52 (O_52,N_6906,N_5315);
and UO_53 (O_53,N_9081,N_7435);
or UO_54 (O_54,N_8410,N_9130);
nor UO_55 (O_55,N_8671,N_5659);
and UO_56 (O_56,N_7333,N_7996);
and UO_57 (O_57,N_5249,N_6964);
and UO_58 (O_58,N_6596,N_9592);
and UO_59 (O_59,N_7859,N_8428);
and UO_60 (O_60,N_5674,N_8366);
or UO_61 (O_61,N_6023,N_8691);
or UO_62 (O_62,N_5982,N_8528);
nor UO_63 (O_63,N_9607,N_5330);
nand UO_64 (O_64,N_9310,N_7027);
nor UO_65 (O_65,N_5056,N_6622);
xnor UO_66 (O_66,N_9011,N_5354);
xor UO_67 (O_67,N_8526,N_5616);
nand UO_68 (O_68,N_6322,N_6422);
nor UO_69 (O_69,N_5245,N_6008);
nor UO_70 (O_70,N_8015,N_8083);
and UO_71 (O_71,N_6103,N_7460);
or UO_72 (O_72,N_8072,N_6564);
or UO_73 (O_73,N_5295,N_5521);
nor UO_74 (O_74,N_9405,N_7089);
nor UO_75 (O_75,N_7556,N_9414);
or UO_76 (O_76,N_6892,N_7503);
and UO_77 (O_77,N_6286,N_7337);
nand UO_78 (O_78,N_5848,N_8435);
or UO_79 (O_79,N_7839,N_9770);
and UO_80 (O_80,N_9054,N_9655);
nor UO_81 (O_81,N_9242,N_6227);
or UO_82 (O_82,N_9596,N_6198);
and UO_83 (O_83,N_9049,N_5378);
nand UO_84 (O_84,N_8997,N_7413);
or UO_85 (O_85,N_6581,N_8305);
or UO_86 (O_86,N_9733,N_9705);
and UO_87 (O_87,N_5911,N_7936);
nor UO_88 (O_88,N_8361,N_7791);
nor UO_89 (O_89,N_5910,N_7825);
and UO_90 (O_90,N_5029,N_8928);
nor UO_91 (O_91,N_6202,N_5779);
or UO_92 (O_92,N_9635,N_8814);
or UO_93 (O_93,N_7107,N_7776);
and UO_94 (O_94,N_7070,N_5630);
nor UO_95 (O_95,N_6902,N_5132);
nand UO_96 (O_96,N_6125,N_8383);
or UO_97 (O_97,N_9270,N_9555);
nor UO_98 (O_98,N_5572,N_6330);
nor UO_99 (O_99,N_6277,N_9219);
or UO_100 (O_100,N_8670,N_8961);
or UO_101 (O_101,N_5545,N_5005);
and UO_102 (O_102,N_5069,N_5685);
nor UO_103 (O_103,N_5880,N_8657);
nor UO_104 (O_104,N_8885,N_5951);
and UO_105 (O_105,N_5924,N_8552);
nor UO_106 (O_106,N_5328,N_6108);
or UO_107 (O_107,N_6343,N_8119);
nor UO_108 (O_108,N_5472,N_8655);
nand UO_109 (O_109,N_6005,N_7283);
nand UO_110 (O_110,N_8952,N_7865);
nand UO_111 (O_111,N_6132,N_8241);
nand UO_112 (O_112,N_9099,N_8029);
nand UO_113 (O_113,N_8067,N_8093);
and UO_114 (O_114,N_7924,N_7090);
xnor UO_115 (O_115,N_8702,N_6130);
or UO_116 (O_116,N_5373,N_7675);
nor UO_117 (O_117,N_6752,N_5799);
nor UO_118 (O_118,N_7781,N_9845);
nor UO_119 (O_119,N_7495,N_7629);
nor UO_120 (O_120,N_5857,N_8881);
nor UO_121 (O_121,N_8866,N_9047);
nand UO_122 (O_122,N_6354,N_6266);
and UO_123 (O_123,N_6712,N_5497);
nor UO_124 (O_124,N_9268,N_6200);
and UO_125 (O_125,N_7285,N_9290);
or UO_126 (O_126,N_8463,N_8726);
nand UO_127 (O_127,N_5412,N_9352);
or UO_128 (O_128,N_9443,N_8249);
nand UO_129 (O_129,N_8799,N_7445);
or UO_130 (O_130,N_8583,N_5844);
and UO_131 (O_131,N_6190,N_6318);
and UO_132 (O_132,N_8009,N_8576);
or UO_133 (O_133,N_6185,N_8356);
and UO_134 (O_134,N_6876,N_8445);
and UO_135 (O_135,N_6805,N_8967);
nand UO_136 (O_136,N_7112,N_9810);
and UO_137 (O_137,N_7075,N_9762);
or UO_138 (O_138,N_8461,N_7235);
nor UO_139 (O_139,N_8240,N_5004);
or UO_140 (O_140,N_8642,N_5753);
nand UO_141 (O_141,N_6569,N_8634);
or UO_142 (O_142,N_9940,N_9170);
or UO_143 (O_143,N_7980,N_9914);
nand UO_144 (O_144,N_5589,N_6235);
and UO_145 (O_145,N_7827,N_5777);
nand UO_146 (O_146,N_5578,N_8519);
nand UO_147 (O_147,N_7973,N_5022);
and UO_148 (O_148,N_9122,N_8633);
or UO_149 (O_149,N_6612,N_5617);
nor UO_150 (O_150,N_7671,N_7212);
or UO_151 (O_151,N_5549,N_7456);
nor UO_152 (O_152,N_9866,N_7573);
and UO_153 (O_153,N_5528,N_9839);
and UO_154 (O_154,N_8216,N_9617);
nand UO_155 (O_155,N_7078,N_6798);
nor UO_156 (O_156,N_8123,N_7356);
nor UO_157 (O_157,N_6696,N_6697);
nand UO_158 (O_158,N_5757,N_7259);
nor UO_159 (O_159,N_5428,N_7086);
nor UO_160 (O_160,N_5426,N_6104);
nor UO_161 (O_161,N_7785,N_7172);
nor UO_162 (O_162,N_7940,N_8338);
or UO_163 (O_163,N_5172,N_6315);
and UO_164 (O_164,N_8516,N_8924);
or UO_165 (O_165,N_8759,N_6020);
and UO_166 (O_166,N_6944,N_5730);
nor UO_167 (O_167,N_6471,N_9747);
nand UO_168 (O_168,N_7249,N_6774);
and UO_169 (O_169,N_6758,N_9388);
and UO_170 (O_170,N_6081,N_5156);
and UO_171 (O_171,N_9547,N_8213);
nand UO_172 (O_172,N_8946,N_6159);
nand UO_173 (O_173,N_9653,N_9492);
nor UO_174 (O_174,N_7690,N_5838);
or UO_175 (O_175,N_9028,N_7853);
nand UO_176 (O_176,N_8048,N_6968);
and UO_177 (O_177,N_7346,N_7901);
nand UO_178 (O_178,N_8030,N_8116);
or UO_179 (O_179,N_5227,N_5881);
nand UO_180 (O_180,N_8693,N_5579);
nand UO_181 (O_181,N_6351,N_6895);
and UO_182 (O_182,N_5647,N_5350);
or UO_183 (O_183,N_9213,N_5023);
nand UO_184 (O_184,N_6561,N_9735);
or UO_185 (O_185,N_6938,N_9141);
nand UO_186 (O_186,N_9965,N_5812);
nor UO_187 (O_187,N_5986,N_6538);
nand UO_188 (O_188,N_5506,N_7260);
or UO_189 (O_189,N_9792,N_6967);
or UO_190 (O_190,N_6905,N_9363);
nand UO_191 (O_191,N_8848,N_5675);
xnor UO_192 (O_192,N_6110,N_7429);
nand UO_193 (O_193,N_9306,N_7846);
nor UO_194 (O_194,N_9699,N_9228);
nand UO_195 (O_195,N_9157,N_5532);
nand UO_196 (O_196,N_6060,N_7786);
or UO_197 (O_197,N_6601,N_6526);
or UO_198 (O_198,N_5268,N_9591);
and UO_199 (O_199,N_6808,N_7746);
nor UO_200 (O_200,N_8341,N_8419);
or UO_201 (O_201,N_8151,N_7861);
nor UO_202 (O_202,N_8209,N_6848);
or UO_203 (O_203,N_9647,N_9666);
nor UO_204 (O_204,N_8948,N_9947);
nor UO_205 (O_205,N_8073,N_5325);
nand UO_206 (O_206,N_5503,N_5781);
nor UO_207 (O_207,N_8556,N_7388);
or UO_208 (O_208,N_9276,N_9800);
or UO_209 (O_209,N_7611,N_7211);
and UO_210 (O_210,N_9065,N_5389);
or UO_211 (O_211,N_5700,N_9421);
nor UO_212 (O_212,N_8478,N_8856);
and UO_213 (O_213,N_7189,N_9086);
and UO_214 (O_214,N_8704,N_8411);
nand UO_215 (O_215,N_9868,N_6673);
nor UO_216 (O_216,N_5547,N_9614);
or UO_217 (O_217,N_5207,N_5006);
xor UO_218 (O_218,N_6312,N_8715);
nor UO_219 (O_219,N_8719,N_6737);
or UO_220 (O_220,N_9568,N_5376);
or UO_221 (O_221,N_9546,N_6771);
and UO_222 (O_222,N_9437,N_5273);
nand UO_223 (O_223,N_7567,N_6233);
nor UO_224 (O_224,N_5368,N_9178);
and UO_225 (O_225,N_7165,N_5992);
nand UO_226 (O_226,N_8497,N_6925);
and UO_227 (O_227,N_9527,N_9008);
nor UO_228 (O_228,N_7308,N_6177);
nor UO_229 (O_229,N_7595,N_7479);
nand UO_230 (O_230,N_6241,N_9600);
nor UO_231 (O_231,N_5037,N_8248);
or UO_232 (O_232,N_9365,N_5255);
and UO_233 (O_233,N_8607,N_6559);
or UO_234 (O_234,N_7226,N_8271);
nor UO_235 (O_235,N_7054,N_7634);
or UO_236 (O_236,N_6082,N_9037);
or UO_237 (O_237,N_7480,N_8756);
or UO_238 (O_238,N_6704,N_8569);
nand UO_239 (O_239,N_9474,N_8650);
nor UO_240 (O_240,N_8760,N_6634);
and UO_241 (O_241,N_6827,N_9820);
and UO_242 (O_242,N_6188,N_9171);
and UO_243 (O_243,N_9860,N_7101);
and UO_244 (O_244,N_6206,N_7096);
or UO_245 (O_245,N_6062,N_7416);
nor UO_246 (O_246,N_6083,N_6787);
nand UO_247 (O_247,N_7674,N_8420);
nor UO_248 (O_248,N_7907,N_9826);
and UO_249 (O_249,N_7902,N_9695);
nor UO_250 (O_250,N_5116,N_6603);
or UO_251 (O_251,N_7857,N_6232);
nand UO_252 (O_252,N_5726,N_8930);
or UO_253 (O_253,N_6380,N_7888);
and UO_254 (O_254,N_6723,N_7397);
xnor UO_255 (O_255,N_5884,N_5573);
nand UO_256 (O_256,N_8754,N_6153);
and UO_257 (O_257,N_6209,N_6393);
nor UO_258 (O_258,N_9261,N_6810);
nand UO_259 (O_259,N_7365,N_5727);
or UO_260 (O_260,N_7467,N_8549);
nor UO_261 (O_261,N_8602,N_9500);
xor UO_262 (O_262,N_7403,N_5692);
and UO_263 (O_263,N_5562,N_7522);
and UO_264 (O_264,N_6698,N_7446);
or UO_265 (O_265,N_7989,N_8816);
nor UO_266 (O_266,N_9687,N_5160);
nand UO_267 (O_267,N_9216,N_6017);
nand UO_268 (O_268,N_8235,N_5062);
and UO_269 (O_269,N_8162,N_5224);
or UO_270 (O_270,N_6523,N_9796);
and UO_271 (O_271,N_7349,N_9034);
nor UO_272 (O_272,N_6293,N_7679);
or UO_273 (O_273,N_8730,N_7970);
and UO_274 (O_274,N_7312,N_5770);
nand UO_275 (O_275,N_9952,N_9284);
nor UO_276 (O_276,N_6796,N_6617);
nand UO_277 (O_277,N_7275,N_7072);
or UO_278 (O_278,N_9324,N_9605);
or UO_279 (O_279,N_6971,N_9911);
nor UO_280 (O_280,N_5110,N_7138);
nand UO_281 (O_281,N_8582,N_9549);
xnor UO_282 (O_282,N_5842,N_8931);
nand UO_283 (O_283,N_9958,N_5855);
nor UO_284 (O_284,N_5424,N_9470);
nor UO_285 (O_285,N_9282,N_9700);
nand UO_286 (O_286,N_5403,N_6901);
nor UO_287 (O_287,N_6089,N_5015);
nor UO_288 (O_288,N_8585,N_9133);
nand UO_289 (O_289,N_5731,N_5349);
xor UO_290 (O_290,N_6297,N_5491);
nor UO_291 (O_291,N_5712,N_8061);
nand UO_292 (O_292,N_6327,N_6969);
nor UO_293 (O_293,N_9435,N_6091);
and UO_294 (O_294,N_6678,N_5720);
nand UO_295 (O_295,N_7624,N_6792);
or UO_296 (O_296,N_7191,N_6150);
or UO_297 (O_297,N_8299,N_9515);
and UO_298 (O_298,N_5441,N_8328);
and UO_299 (O_299,N_8078,N_6437);
nor UO_300 (O_300,N_6695,N_7152);
nor UO_301 (O_301,N_7176,N_8918);
nor UO_302 (O_302,N_5152,N_9996);
nand UO_303 (O_303,N_9158,N_6438);
and UO_304 (O_304,N_8471,N_5401);
and UO_305 (O_305,N_9145,N_5063);
nand UO_306 (O_306,N_5643,N_5978);
and UO_307 (O_307,N_8781,N_8220);
and UO_308 (O_308,N_5668,N_8016);
or UO_309 (O_309,N_6677,N_5974);
nand UO_310 (O_310,N_7771,N_6854);
or UO_311 (O_311,N_9672,N_8770);
and UO_312 (O_312,N_7733,N_5442);
nand UO_313 (O_313,N_8899,N_8019);
or UO_314 (O_314,N_9062,N_8813);
nand UO_315 (O_315,N_8329,N_9633);
nor UO_316 (O_316,N_9750,N_6835);
nor UO_317 (O_317,N_5768,N_8685);
xnor UO_318 (O_318,N_8055,N_5701);
or UO_319 (O_319,N_5086,N_5101);
nand UO_320 (O_320,N_9651,N_6379);
and UO_321 (O_321,N_6862,N_8441);
and UO_322 (O_322,N_6240,N_5833);
nor UO_323 (O_323,N_5377,N_7058);
and UO_324 (O_324,N_5673,N_5597);
nand UO_325 (O_325,N_8052,N_8263);
nand UO_326 (O_326,N_6176,N_9342);
nand UO_327 (O_327,N_6489,N_6705);
and UO_328 (O_328,N_7642,N_7498);
nor UO_329 (O_329,N_9638,N_6171);
or UO_330 (O_330,N_9066,N_7631);
nor UO_331 (O_331,N_6527,N_6050);
or UO_332 (O_332,N_6914,N_5546);
nand UO_333 (O_333,N_5238,N_7046);
nand UO_334 (O_334,N_8457,N_6418);
or UO_335 (O_335,N_6229,N_9425);
nor UO_336 (O_336,N_6165,N_8611);
nor UO_337 (O_337,N_9938,N_5899);
nand UO_338 (O_338,N_5743,N_6246);
and UO_339 (O_339,N_6700,N_8125);
nand UO_340 (O_340,N_6382,N_9485);
or UO_341 (O_341,N_5133,N_8283);
or UO_342 (O_342,N_5906,N_8787);
nor UO_343 (O_343,N_6311,N_6288);
nor UO_344 (O_344,N_9937,N_7657);
nand UO_345 (O_345,N_8266,N_9375);
nand UO_346 (O_346,N_5134,N_8292);
or UO_347 (O_347,N_9483,N_8158);
nand UO_348 (O_348,N_8674,N_9245);
and UO_349 (O_349,N_7955,N_9366);
nor UO_350 (O_350,N_6543,N_6813);
nor UO_351 (O_351,N_9794,N_7324);
and UO_352 (O_352,N_9051,N_8094);
and UO_353 (O_353,N_6133,N_9552);
nand UO_354 (O_354,N_5118,N_5289);
nor UO_355 (O_355,N_7323,N_7062);
and UO_356 (O_356,N_6264,N_7311);
and UO_357 (O_357,N_9950,N_8751);
nand UO_358 (O_358,N_5433,N_9226);
nand UO_359 (O_359,N_8335,N_7793);
or UO_360 (O_360,N_7120,N_7706);
nand UO_361 (O_361,N_6279,N_6802);
and UO_362 (O_362,N_7713,N_9340);
nor UO_363 (O_363,N_7625,N_8004);
and UO_364 (O_364,N_7991,N_5905);
and UO_365 (O_365,N_6113,N_8182);
nor UO_366 (O_366,N_8802,N_6878);
or UO_367 (O_367,N_7080,N_8316);
xnor UO_368 (O_368,N_9807,N_8057);
and UO_369 (O_369,N_7903,N_6006);
nand UO_370 (O_370,N_8652,N_8393);
nand UO_371 (O_371,N_7571,N_9682);
nor UO_372 (O_372,N_7250,N_7041);
nand UO_373 (O_373,N_6979,N_6531);
nor UO_374 (O_374,N_6292,N_5922);
nand UO_375 (O_375,N_8827,N_9248);
and UO_376 (O_376,N_6528,N_6497);
xnor UO_377 (O_377,N_6204,N_5830);
nor UO_378 (O_378,N_8036,N_9015);
nand UO_379 (O_379,N_7929,N_5934);
and UO_380 (O_380,N_5494,N_9928);
and UO_381 (O_381,N_6466,N_8599);
or UO_382 (O_382,N_5026,N_7011);
nand UO_383 (O_383,N_6116,N_7650);
nand UO_384 (O_384,N_9854,N_5123);
nor UO_385 (O_385,N_6276,N_5252);
or UO_386 (O_386,N_5140,N_9347);
or UO_387 (O_387,N_6219,N_6481);
and UO_388 (O_388,N_9476,N_9696);
nor UO_389 (O_389,N_8649,N_7803);
nor UO_390 (O_390,N_8981,N_8350);
nor UO_391 (O_391,N_5710,N_9882);
or UO_392 (O_392,N_7060,N_9579);
and UO_393 (O_393,N_8929,N_6419);
nand UO_394 (O_394,N_7339,N_8184);
or UO_395 (O_395,N_6178,N_9539);
nor UO_396 (O_396,N_5979,N_7019);
nand UO_397 (O_397,N_7423,N_5556);
nand UO_398 (O_398,N_7038,N_9232);
nand UO_399 (O_399,N_6769,N_9734);
nor UO_400 (O_400,N_5078,N_9382);
and UO_401 (O_401,N_9444,N_9999);
nand UO_402 (O_402,N_6284,N_6166);
or UO_403 (O_403,N_6811,N_6960);
and UO_404 (O_404,N_8834,N_8402);
and UO_405 (O_405,N_8088,N_7052);
or UO_406 (O_406,N_5068,N_5930);
nand UO_407 (O_407,N_5300,N_9254);
or UO_408 (O_408,N_7351,N_5530);
or UO_409 (O_409,N_5177,N_7597);
nor UO_410 (O_410,N_7554,N_7593);
nand UO_411 (O_411,N_6838,N_9314);
nand UO_412 (O_412,N_5124,N_5776);
nand UO_413 (O_413,N_8855,N_7641);
nand UO_414 (O_414,N_7754,N_7313);
or UO_415 (O_415,N_8215,N_8577);
xnor UO_416 (O_416,N_6766,N_6585);
and UO_417 (O_417,N_5559,N_9869);
nand UO_418 (O_418,N_6408,N_8175);
nand UO_419 (O_419,N_8551,N_9477);
or UO_420 (O_420,N_8204,N_5011);
nand UO_421 (O_421,N_8502,N_5914);
nand UO_422 (O_422,N_9106,N_5170);
and UO_423 (O_423,N_6447,N_7960);
and UO_424 (O_424,N_8499,N_8342);
or UO_425 (O_425,N_5155,N_6186);
or UO_426 (O_426,N_6891,N_8978);
or UO_427 (O_427,N_6899,N_8149);
or UO_428 (O_428,N_9718,N_5183);
or UO_429 (O_429,N_7219,N_6921);
nor UO_430 (O_430,N_9986,N_6726);
nor UO_431 (O_431,N_5281,N_9832);
and UO_432 (O_432,N_9075,N_9423);
nor UO_433 (O_433,N_7581,N_9720);
nand UO_434 (O_434,N_5102,N_7229);
and UO_435 (O_435,N_7967,N_7251);
or UO_436 (O_436,N_7681,N_8849);
nor UO_437 (O_437,N_7767,N_9809);
and UO_438 (O_438,N_8110,N_9128);
or UO_439 (O_439,N_9799,N_5317);
nand UO_440 (O_440,N_6461,N_8498);
or UO_441 (O_441,N_6943,N_6674);
and UO_442 (O_442,N_7427,N_6075);
and UO_443 (O_443,N_9438,N_5678);
and UO_444 (O_444,N_7407,N_8446);
nor UO_445 (O_445,N_5752,N_9512);
nor UO_446 (O_446,N_6255,N_6203);
nor UO_447 (O_447,N_5473,N_5602);
or UO_448 (O_448,N_7253,N_6245);
or UO_449 (O_449,N_8700,N_9208);
and UO_450 (O_450,N_5091,N_6360);
or UO_451 (O_451,N_9513,N_7852);
nor UO_452 (O_452,N_6953,N_6778);
or UO_453 (O_453,N_9772,N_8301);
nor UO_454 (O_454,N_8629,N_6716);
nand UO_455 (O_455,N_8090,N_7057);
or UO_456 (O_456,N_9831,N_9639);
and UO_457 (O_457,N_8980,N_7552);
or UO_458 (O_458,N_5485,N_5603);
or UO_459 (O_459,N_5984,N_7979);
or UO_460 (O_460,N_9409,N_8534);
and UO_461 (O_461,N_6722,N_5136);
and UO_462 (O_462,N_5972,N_5875);
or UO_463 (O_463,N_5417,N_9067);
nor UO_464 (O_464,N_9356,N_8690);
nor UO_465 (O_465,N_8973,N_7748);
and UO_466 (O_466,N_9077,N_8062);
and UO_467 (O_467,N_9844,N_5805);
or UO_468 (O_468,N_9864,N_7257);
or UO_469 (O_469,N_8803,N_9896);
and UO_470 (O_470,N_5894,N_7032);
nand UO_471 (O_471,N_5593,N_8321);
nand UO_472 (O_472,N_6031,N_7589);
and UO_473 (O_473,N_7303,N_5478);
nor UO_474 (O_474,N_6500,N_7157);
or UO_475 (O_475,N_5619,N_6409);
nor UO_476 (O_476,N_8805,N_5971);
or UO_477 (O_477,N_6034,N_7999);
nor UO_478 (O_478,N_9825,N_9956);
nand UO_479 (O_479,N_8415,N_7097);
nor UO_480 (O_480,N_6645,N_9294);
or UO_481 (O_481,N_8348,N_8174);
nand UO_482 (O_482,N_5737,N_7099);
nor UO_483 (O_483,N_8012,N_5274);
nor UO_484 (O_484,N_5297,N_5671);
and UO_485 (O_485,N_9706,N_5775);
and UO_486 (O_486,N_9308,N_9878);
or UO_487 (O_487,N_5806,N_9348);
nor UO_488 (O_488,N_6900,N_9954);
xnor UO_489 (O_489,N_8605,N_8259);
nor UO_490 (O_490,N_5126,N_5210);
or UO_491 (O_491,N_8965,N_6767);
and UO_492 (O_492,N_9450,N_5874);
nor UO_493 (O_493,N_9867,N_6659);
or UO_494 (O_494,N_7020,N_8481);
and UO_495 (O_495,N_9578,N_8343);
nand UO_496 (O_496,N_9353,N_6348);
or UO_497 (O_497,N_5553,N_5411);
or UO_498 (O_498,N_7093,N_9737);
nand UO_499 (O_499,N_8508,N_5965);
or UO_500 (O_500,N_6029,N_8339);
and UO_501 (O_501,N_6764,N_5476);
nor UO_502 (O_502,N_8990,N_6149);
or UO_503 (O_503,N_6468,N_8086);
or UO_504 (O_504,N_9288,N_9004);
or UO_505 (O_505,N_8819,N_9472);
and UO_506 (O_506,N_7173,N_8291);
nand UO_507 (O_507,N_6924,N_9741);
and UO_508 (O_508,N_8560,N_5218);
nand UO_509 (O_509,N_8008,N_8733);
nor UO_510 (O_510,N_5284,N_6517);
nor UO_511 (O_511,N_7702,N_9805);
and UO_512 (O_512,N_7835,N_9943);
and UO_513 (O_513,N_8112,N_8836);
and UO_514 (O_514,N_8392,N_9123);
nand UO_515 (O_515,N_9302,N_8991);
nand UO_516 (O_516,N_5014,N_8477);
or UO_517 (O_517,N_7217,N_5642);
nor UO_518 (O_518,N_6158,N_7068);
or UO_519 (O_519,N_7764,N_9389);
nor UO_520 (O_520,N_5822,N_7922);
nor UO_521 (O_521,N_9753,N_6864);
nand UO_522 (O_522,N_8340,N_5039);
nand UO_523 (O_523,N_5247,N_5361);
and UO_524 (O_524,N_7433,N_7558);
or UO_525 (O_525,N_5266,N_7883);
nand UO_526 (O_526,N_7347,N_6604);
nor UO_527 (O_527,N_8432,N_9312);
nor UO_528 (O_528,N_9757,N_9266);
nor UO_529 (O_529,N_7410,N_6649);
and UO_530 (O_530,N_5636,N_7774);
or UO_531 (O_531,N_6037,N_5159);
or UO_532 (O_532,N_7336,N_9112);
or UO_533 (O_533,N_8367,N_5076);
nor UO_534 (O_534,N_9328,N_5660);
nand UO_535 (O_535,N_5677,N_8613);
nand UO_536 (O_536,N_7307,N_9606);
and UO_537 (O_537,N_6151,N_6222);
and UO_538 (O_538,N_7400,N_9544);
nand UO_539 (O_539,N_5862,N_5687);
and UO_540 (O_540,N_8101,N_8039);
or UO_541 (O_541,N_8370,N_7067);
and UO_542 (O_542,N_8872,N_6234);
nor UO_543 (O_543,N_8955,N_9749);
or UO_544 (O_544,N_5169,N_9766);
or UO_545 (O_545,N_6717,N_5606);
nor UO_546 (O_546,N_7290,N_8947);
or UO_547 (O_547,N_5734,N_5018);
or UO_548 (O_548,N_6533,N_9267);
nor UO_549 (O_549,N_5052,N_5338);
and UO_550 (O_550,N_5908,N_6120);
nor UO_551 (O_551,N_7672,N_7660);
and UO_552 (O_552,N_6799,N_6859);
or UO_553 (O_553,N_8912,N_9722);
nor UO_554 (O_554,N_7937,N_7224);
nor UO_555 (O_555,N_7442,N_6650);
nor UO_556 (O_556,N_6667,N_7205);
or UO_557 (O_557,N_6839,N_7222);
nand UO_558 (O_558,N_6627,N_6144);
nor UO_559 (O_559,N_9742,N_5229);
and UO_560 (O_560,N_9033,N_9084);
nor UO_561 (O_561,N_8187,N_7348);
and UO_562 (O_562,N_5484,N_9945);
or UO_563 (O_563,N_8571,N_8395);
and UO_564 (O_564,N_5913,N_9159);
or UO_565 (O_565,N_8987,N_6857);
or UO_566 (O_566,N_9494,N_7738);
nor UO_567 (O_567,N_7830,N_7758);
or UO_568 (O_568,N_8986,N_7539);
and UO_569 (O_569,N_9519,N_8500);
and UO_570 (O_570,N_5464,N_7586);
or UO_571 (O_571,N_6356,N_5117);
or UO_572 (O_572,N_6458,N_9571);
nand UO_573 (O_573,N_5879,N_5919);
xor UO_574 (O_574,N_9721,N_9360);
or UO_575 (O_575,N_6412,N_5027);
or UO_576 (O_576,N_7542,N_5932);
and UO_577 (O_577,N_9387,N_6598);
or UO_578 (O_578,N_9625,N_9833);
and UO_579 (O_579,N_6636,N_9379);
or UO_580 (O_580,N_7073,N_6337);
nor UO_581 (O_581,N_7241,N_6195);
nand UO_582 (O_582,N_5293,N_9506);
and UO_583 (O_583,N_7376,N_8745);
and UO_584 (O_584,N_6164,N_7459);
or UO_585 (O_585,N_6793,N_6454);
or UO_586 (O_586,N_9147,N_7787);
nand UO_587 (O_587,N_8466,N_9109);
nor UO_588 (O_588,N_7387,N_8847);
nand UO_589 (O_589,N_5352,N_7661);
nand UO_590 (O_590,N_7899,N_7505);
or UO_591 (O_591,N_9587,N_5337);
or UO_592 (O_592,N_7133,N_9953);
or UO_593 (O_593,N_9393,N_6557);
nand UO_594 (O_594,N_5051,N_7472);
nor UO_595 (O_595,N_5686,N_5109);
and UO_596 (O_596,N_5467,N_6094);
nand UO_597 (O_597,N_9643,N_7318);
nor UO_598 (O_598,N_6244,N_8251);
or UO_599 (O_599,N_5406,N_6154);
nand UO_600 (O_600,N_7598,N_9331);
nand UO_601 (O_601,N_8403,N_9196);
nand UO_602 (O_602,N_6080,N_8812);
nand UO_603 (O_603,N_7678,N_5702);
or UO_604 (O_604,N_7008,N_6747);
and UO_605 (O_605,N_6242,N_7238);
nor UO_606 (O_606,N_8573,N_9204);
nand UO_607 (O_607,N_7540,N_9783);
nor UO_608 (O_608,N_7134,N_7181);
and UO_609 (O_609,N_9055,N_5832);
and UO_610 (O_610,N_6929,N_6995);
nor UO_611 (O_611,N_8372,N_5385);
or UO_612 (O_612,N_8128,N_9061);
nand UO_613 (O_613,N_9396,N_7644);
nor UO_614 (O_614,N_6401,N_8423);
and UO_615 (O_615,N_7806,N_5423);
and UO_616 (O_616,N_6057,N_8319);
or UO_617 (O_617,N_9487,N_6699);
or UO_618 (O_618,N_9481,N_9305);
nor UO_619 (O_619,N_6916,N_8437);
and UO_620 (O_620,N_8013,N_7039);
nand UO_621 (O_621,N_6840,N_7698);
and UO_622 (O_622,N_9272,N_7688);
nand UO_623 (O_623,N_7037,N_7836);
nand UO_624 (O_624,N_9823,N_8096);
and UO_625 (O_625,N_5469,N_7248);
or UO_626 (O_626,N_6630,N_5278);
nand UO_627 (O_627,N_8851,N_8114);
or UO_628 (O_628,N_6044,N_8897);
or UO_629 (O_629,N_9939,N_5128);
or UO_630 (O_630,N_6141,N_6658);
and UO_631 (O_631,N_9143,N_6096);
nand UO_632 (O_632,N_9627,N_9767);
nor UO_633 (O_633,N_8068,N_7869);
or UO_634 (O_634,N_5945,N_9644);
and UO_635 (O_635,N_6294,N_6357);
or UO_636 (O_636,N_9017,N_5847);
nand UO_637 (O_637,N_6404,N_8260);
and UO_638 (O_638,N_5501,N_7452);
and UO_639 (O_639,N_9104,N_8064);
and UO_640 (O_640,N_7945,N_7831);
and UO_641 (O_641,N_8409,N_5310);
and UO_642 (O_642,N_8926,N_8589);
nor UO_643 (O_643,N_8021,N_5233);
nand UO_644 (O_644,N_6220,N_9319);
or UO_645 (O_645,N_7696,N_6230);
and UO_646 (O_646,N_8491,N_6988);
nor UO_647 (O_647,N_9948,N_6370);
and UO_648 (O_648,N_9223,N_9138);
and UO_649 (O_649,N_9070,N_5463);
nand UO_650 (O_650,N_5835,N_6870);
nand UO_651 (O_651,N_7736,N_5962);
nor UO_652 (O_652,N_6801,N_5513);
and UO_653 (O_653,N_6323,N_9449);
or UO_654 (O_654,N_9001,N_6262);
nor UO_655 (O_655,N_7557,N_7860);
nand UO_656 (O_656,N_5739,N_9043);
or UO_657 (O_657,N_6963,N_5093);
and UO_658 (O_658,N_8053,N_8077);
nor UO_659 (O_659,N_6385,N_7053);
and UO_660 (O_660,N_7800,N_6654);
nor UO_661 (O_661,N_8663,N_7496);
nand UO_662 (O_662,N_5396,N_9155);
and UO_663 (O_663,N_7103,N_6494);
and UO_664 (O_664,N_9230,N_5237);
or UO_665 (O_665,N_8721,N_5313);
nand UO_666 (O_666,N_9227,N_5845);
and UO_667 (O_667,N_6826,N_9836);
or UO_668 (O_668,N_7431,N_7166);
and UO_669 (O_669,N_6274,N_5564);
and UO_670 (O_670,N_6844,N_5158);
nor UO_671 (O_671,N_5622,N_6541);
nor UO_672 (O_672,N_9468,N_9486);
or UO_673 (O_673,N_8797,N_7833);
nor UO_674 (O_674,N_6930,N_9697);
or UO_675 (O_675,N_7514,N_7659);
or UO_676 (O_676,N_7325,N_8586);
and UO_677 (O_677,N_6539,N_9787);
nand UO_678 (O_678,N_8694,N_9289);
and UO_679 (O_679,N_8479,N_5656);
nand UO_680 (O_680,N_7051,N_9212);
or UO_681 (O_681,N_5119,N_6545);
nand UO_682 (O_682,N_6926,N_7926);
and UO_683 (O_683,N_6407,N_8050);
nand UO_684 (O_684,N_7995,N_9374);
nand UO_685 (O_685,N_5903,N_8537);
nand UO_686 (O_686,N_8345,N_6550);
nand UO_687 (O_687,N_7055,N_7095);
or UO_688 (O_688,N_9525,N_7626);
or UO_689 (O_689,N_6515,N_5742);
or UO_690 (O_690,N_9646,N_6417);
and UO_691 (O_691,N_8977,N_6320);
and UO_692 (O_692,N_5460,N_6945);
nor UO_693 (O_693,N_9537,N_8103);
and UO_694 (O_694,N_8763,N_8937);
or UO_695 (O_695,N_6573,N_8774);
nor UO_696 (O_696,N_5891,N_5316);
nand UO_697 (O_697,N_9073,N_6207);
nand UO_698 (O_698,N_5137,N_7372);
nor UO_699 (O_699,N_9041,N_5998);
nand UO_700 (O_700,N_9025,N_9269);
nand UO_701 (O_701,N_6095,N_9050);
nor UO_702 (O_702,N_7566,N_5046);
nor UO_703 (O_703,N_6549,N_5228);
and UO_704 (O_704,N_7383,N_7016);
nand UO_705 (O_705,N_9880,N_7292);
and UO_706 (O_706,N_6614,N_7695);
and UO_707 (O_707,N_8172,N_7933);
nor UO_708 (O_708,N_5688,N_7939);
and UO_709 (O_709,N_7137,N_8738);
xnor UO_710 (O_710,N_6632,N_6886);
nand UO_711 (O_711,N_7950,N_9784);
nand UO_712 (O_712,N_5364,N_5950);
nor UO_713 (O_713,N_6624,N_9299);
xor UO_714 (O_714,N_5362,N_8495);
or UO_715 (O_715,N_7056,N_7515);
nand UO_716 (O_716,N_9376,N_6451);
nor UO_717 (O_717,N_5658,N_7004);
nand UO_718 (O_718,N_5926,N_7630);
nor UO_719 (O_719,N_8089,N_6252);
and UO_720 (O_720,N_8992,N_9575);
nor UO_721 (O_721,N_8902,N_7583);
nor UO_722 (O_722,N_7662,N_5605);
or UO_723 (O_723,N_7981,N_6552);
nor UO_724 (O_724,N_8632,N_6592);
nor UO_725 (O_725,N_7218,N_8771);
and UO_726 (O_726,N_8486,N_7875);
and UO_727 (O_727,N_6179,N_8740);
and UO_728 (O_728,N_8857,N_6729);
or UO_729 (O_729,N_5088,N_7141);
nor UO_730 (O_730,N_6849,N_6137);
or UO_731 (O_731,N_6097,N_8277);
or UO_732 (O_732,N_5163,N_9765);
or UO_733 (O_733,N_9400,N_6342);
nor UO_734 (O_734,N_5360,N_9645);
nor UO_735 (O_735,N_5358,N_9658);
or UO_736 (O_736,N_7782,N_5802);
nor UO_737 (O_737,N_5277,N_8609);
nand UO_738 (O_738,N_7048,N_6711);
and UO_739 (O_739,N_8817,N_9790);
or UO_740 (O_740,N_9390,N_8910);
nand UO_741 (O_741,N_9475,N_9085);
or UO_742 (O_742,N_9611,N_8426);
and UO_743 (O_743,N_6441,N_7108);
and UO_744 (O_744,N_9829,N_6600);
nand UO_745 (O_745,N_7579,N_8853);
or UO_746 (O_746,N_6555,N_5104);
or UO_747 (O_747,N_7225,N_6009);
nor UO_748 (O_748,N_7990,N_5299);
nand UO_749 (O_749,N_5608,N_9949);
nand UO_750 (O_750,N_5877,N_5963);
and UO_751 (O_751,N_5620,N_7976);
and UO_752 (O_752,N_8939,N_7352);
and UO_753 (O_753,N_6492,N_8612);
nand UO_754 (O_754,N_7610,N_7194);
and UO_755 (O_755,N_5261,N_7334);
nor UO_756 (O_756,N_9910,N_8966);
and UO_757 (O_757,N_7392,N_8243);
and UO_758 (O_758,N_8788,N_9599);
nor UO_759 (O_759,N_7826,N_8996);
and UO_760 (O_760,N_6226,N_6763);
nand UO_761 (O_761,N_5820,N_7709);
and UO_762 (O_762,N_6162,N_9793);
nand UO_763 (O_763,N_6978,N_5756);
or UO_764 (O_764,N_5090,N_7563);
nor UO_765 (O_765,N_9121,N_6135);
and UO_766 (O_766,N_8171,N_8320);
nor UO_767 (O_767,N_8137,N_9295);
or UO_768 (O_768,N_5861,N_9031);
and UO_769 (O_769,N_8503,N_6977);
or UO_770 (O_770,N_5017,N_6467);
nand UO_771 (O_771,N_7341,N_6155);
or UO_772 (O_772,N_6329,N_8462);
nor UO_773 (O_773,N_6828,N_7297);
nor UO_774 (O_774,N_9944,N_6710);
and UO_775 (O_775,N_5355,N_7304);
and UO_776 (O_776,N_7206,N_7934);
and UO_777 (O_777,N_8882,N_8035);
or UO_778 (O_778,N_8669,N_7003);
and UO_779 (O_779,N_5173,N_6919);
or UO_780 (O_780,N_6328,N_5801);
nor UO_781 (O_781,N_9467,N_6275);
nor UO_782 (O_782,N_6444,N_5304);
and UO_783 (O_783,N_9162,N_9271);
nand UO_784 (O_784,N_7559,N_7705);
nand UO_785 (O_785,N_8911,N_5475);
nor UO_786 (O_786,N_5980,N_7799);
nand UO_787 (O_787,N_5929,N_9092);
nand UO_788 (O_788,N_9064,N_6221);
nand UO_789 (O_789,N_5253,N_5841);
nor UO_790 (O_790,N_9479,N_9030);
and UO_791 (O_791,N_9367,N_8401);
nand UO_792 (O_792,N_7548,N_9553);
nor UO_793 (O_793,N_7605,N_7242);
and UO_794 (O_794,N_8579,N_7794);
and UO_795 (O_795,N_5780,N_8268);
and UO_796 (O_796,N_6685,N_6540);
and UO_797 (O_797,N_9683,N_7187);
nand UO_798 (O_798,N_9330,N_8570);
or UO_799 (O_799,N_5085,N_8359);
or UO_800 (O_800,N_6631,N_8594);
nand UO_801 (O_801,N_6054,N_7501);
nor UO_802 (O_802,N_6446,N_9981);
nand UO_803 (O_803,N_6371,N_8720);
nor UO_804 (O_804,N_9429,N_8917);
nand UO_805 (O_805,N_8592,N_8159);
or UO_806 (O_806,N_6666,N_7160);
or UO_807 (O_807,N_8353,N_6885);
or UO_808 (O_808,N_8154,N_5311);
and UO_809 (O_809,N_7208,N_9251);
nand UO_810 (O_810,N_9873,N_6670);
nand UO_811 (O_811,N_6021,N_6435);
nand UO_812 (O_812,N_5933,N_6124);
or UO_813 (O_813,N_8547,N_8118);
or UO_814 (O_814,N_5080,N_5670);
and UO_815 (O_815,N_9134,N_5662);
nand UO_816 (O_816,N_9256,N_7155);
nand UO_817 (O_817,N_6856,N_7994);
and UO_818 (O_818,N_9951,N_8564);
nand UO_819 (O_819,N_9110,N_5817);
nor UO_820 (O_820,N_5189,N_9101);
and UO_821 (O_821,N_9895,N_7601);
or UO_822 (O_822,N_6271,N_5318);
nor UO_823 (O_823,N_8117,N_6736);
nand UO_824 (O_824,N_9321,N_5909);
xor UO_825 (O_825,N_9887,N_5949);
nand UO_826 (O_826,N_7953,N_5259);
nor UO_827 (O_827,N_7608,N_5202);
and UO_828 (O_828,N_8107,N_5754);
nor UO_829 (O_829,N_7064,N_9620);
nand UO_830 (O_830,N_5153,N_7959);
nand UO_831 (O_831,N_8279,N_5746);
and UO_832 (O_832,N_8538,N_8993);
nor UO_833 (O_833,N_7692,N_5953);
or UO_834 (O_834,N_5787,N_7844);
or UO_835 (O_835,N_9318,N_6739);
or UO_836 (O_836,N_5380,N_7353);
and UO_837 (O_837,N_7110,N_8010);
or UO_838 (O_838,N_6966,N_6090);
or UO_839 (O_839,N_5520,N_8318);
or UO_840 (O_840,N_6653,N_6707);
nand UO_841 (O_841,N_5956,N_8368);
nand UO_842 (O_842,N_5791,N_8887);
nand UO_843 (O_843,N_9827,N_8876);
and UO_844 (O_844,N_6355,N_5860);
nor UO_845 (O_845,N_7188,N_7638);
or UO_846 (O_846,N_8976,N_6822);
and UO_847 (O_847,N_9381,N_8076);
xnor UO_848 (O_848,N_5723,N_6139);
and UO_849 (O_849,N_6824,N_6635);
and UO_850 (O_850,N_7364,N_7288);
nand UO_851 (O_851,N_5815,N_7240);
nor UO_852 (O_852,N_7651,N_8620);
nor UO_853 (O_853,N_7401,N_7088);
nor UO_854 (O_854,N_8003,N_7541);
and UO_855 (O_855,N_7834,N_7721);
nor UO_856 (O_856,N_8298,N_7012);
and UO_857 (O_857,N_8786,N_9224);
or UO_858 (O_858,N_9142,N_7808);
nor UO_859 (O_859,N_6479,N_9530);
or UO_860 (O_860,N_8267,N_5327);
and UO_861 (O_861,N_9830,N_7546);
nand UO_862 (O_862,N_8226,N_6109);
nor UO_863 (O_863,N_5738,N_5000);
nand UO_864 (O_864,N_6998,N_5867);
nor UO_865 (O_865,N_7543,N_6450);
nand UO_866 (O_866,N_7578,N_7200);
nor UO_867 (O_867,N_5699,N_6087);
nor UO_868 (O_868,N_6831,N_5456);
or UO_869 (O_869,N_9452,N_5935);
or UO_870 (O_870,N_7109,N_7028);
nand UO_871 (O_871,N_7710,N_7358);
and UO_872 (O_872,N_5540,N_5492);
or UO_873 (O_873,N_6004,N_6621);
nand UO_874 (O_874,N_6459,N_9846);
nand UO_875 (O_875,N_6520,N_5367);
and UO_876 (O_876,N_7121,N_6683);
nor UO_877 (O_877,N_8718,N_9659);
nor UO_878 (O_878,N_8925,N_5735);
or UO_879 (O_879,N_6502,N_9283);
nor UO_880 (O_880,N_8555,N_9816);
or UO_881 (O_881,N_7451,N_6299);
nand UO_882 (O_882,N_9899,N_9969);
or UO_883 (O_883,N_5522,N_5645);
or UO_884 (O_884,N_5523,N_7816);
nor UO_885 (O_885,N_8032,N_6400);
and UO_886 (O_886,N_9416,N_8229);
or UO_887 (O_887,N_5682,N_8278);
or UO_888 (O_888,N_5138,N_6287);
nand UO_889 (O_889,N_6332,N_6353);
and UO_890 (O_890,N_6690,N_9988);
and UO_891 (O_891,N_5142,N_5374);
nand UO_892 (O_892,N_7284,N_8678);
and UO_893 (O_893,N_8818,N_5190);
or UO_894 (O_894,N_7750,N_5443);
and UO_895 (O_895,N_7171,N_8310);
nand UO_896 (O_896,N_7391,N_5648);
nand UO_897 (O_897,N_7453,N_9013);
or UO_898 (O_898,N_7477,N_8464);
nor UO_899 (O_899,N_5161,N_7464);
nand UO_900 (O_900,N_8063,N_9535);
nor UO_901 (O_901,N_8042,N_6465);
nor UO_902 (O_902,N_8595,N_6487);
nor UO_903 (O_903,N_6917,N_9129);
and UO_904 (O_904,N_9574,N_8675);
and UO_905 (O_905,N_9018,N_7529);
nor UO_906 (O_906,N_8152,N_8195);
and UO_907 (O_907,N_5661,N_5477);
or UO_908 (O_908,N_6725,N_5448);
or UO_909 (O_909,N_5219,N_9489);
and UO_910 (O_910,N_5591,N_5058);
and UO_911 (O_911,N_8864,N_8779);
xnor UO_912 (O_912,N_7291,N_5511);
or UO_913 (O_913,N_9603,N_8870);
nand UO_914 (O_914,N_8443,N_9859);
or UO_915 (O_915,N_9679,N_6114);
nor UO_916 (O_916,N_7894,N_5359);
or UO_917 (O_917,N_5437,N_8606);
nor UO_918 (O_918,N_7511,N_7509);
or UO_919 (O_919,N_8189,N_8531);
nor UO_920 (O_920,N_9090,N_8011);
or UO_921 (O_921,N_8603,N_5452);
nor UO_922 (O_922,N_8871,N_7555);
nor UO_923 (O_923,N_5638,N_8192);
and UO_924 (O_924,N_5814,N_5976);
or UO_925 (O_925,N_6267,N_8972);
or UO_926 (O_926,N_6633,N_8791);
or UO_927 (O_927,N_7278,N_6381);
nor UO_928 (O_928,N_8542,N_5145);
and UO_929 (O_929,N_8850,N_5379);
and UO_930 (O_930,N_6001,N_5803);
nand UO_931 (O_931,N_8351,N_8102);
nand UO_932 (O_932,N_5298,N_7178);
and UO_933 (O_933,N_8711,N_5543);
or UO_934 (O_934,N_6580,N_6842);
and UO_935 (O_935,N_7895,N_5283);
nand UO_936 (O_936,N_5235,N_5271);
and UO_937 (O_937,N_5127,N_8180);
nand UO_938 (O_938,N_7321,N_5788);
nor UO_939 (O_939,N_6032,N_7462);
nor UO_940 (O_940,N_8134,N_7169);
and UO_941 (O_941,N_7045,N_7031);
nand UO_942 (O_942,N_8163,N_6041);
and UO_943 (O_943,N_7143,N_6761);
and UO_944 (O_944,N_8146,N_6795);
nor UO_945 (O_945,N_6482,N_8286);
or UO_946 (O_946,N_8934,N_5563);
nand UO_947 (O_947,N_7422,N_7213);
and UO_948 (O_948,N_8069,N_6668);
nand UO_949 (O_949,N_5897,N_6610);
nand UO_950 (O_950,N_6036,N_8294);
or UO_951 (O_951,N_5689,N_7504);
nand UO_952 (O_952,N_7919,N_5329);
and UO_953 (O_953,N_7066,N_5055);
or UO_954 (O_954,N_6702,N_8127);
nor UO_955 (O_955,N_6238,N_6836);
nand UO_956 (O_956,N_9168,N_7562);
nand UO_957 (O_957,N_9597,N_5151);
nor UO_958 (O_958,N_6506,N_6554);
nor UO_959 (O_959,N_9876,N_7951);
nor UO_960 (O_960,N_6588,N_7867);
nor UO_961 (O_961,N_8135,N_7792);
nand UO_962 (O_962,N_6268,N_6803);
nor UO_963 (O_963,N_9566,N_9795);
nor UO_964 (O_964,N_8665,N_6475);
and UO_965 (O_965,N_8394,N_6476);
nand UO_966 (O_966,N_9976,N_6338);
and UO_967 (O_967,N_6367,N_9325);
nor UO_968 (O_968,N_6837,N_7743);
and UO_969 (O_969,N_9538,N_8894);
and UO_970 (O_970,N_5209,N_7271);
or UO_971 (O_971,N_8148,N_9343);
nor UO_972 (O_972,N_5952,N_8563);
nor UO_973 (O_973,N_6974,N_9717);
nor UO_974 (O_974,N_5272,N_5471);
or UO_975 (O_975,N_9464,N_9813);
or UO_976 (O_976,N_5499,N_5200);
nand UO_977 (O_977,N_8909,N_5191);
nand UO_978 (O_978,N_6365,N_6590);
nand UO_979 (O_979,N_5607,N_9788);
and UO_980 (O_980,N_9704,N_6243);
nor UO_981 (O_981,N_7691,N_7476);
or UO_982 (O_982,N_9480,N_5527);
or UO_983 (O_983,N_9404,N_6460);
or UO_984 (O_984,N_8873,N_5565);
nand UO_985 (O_985,N_8023,N_8098);
or UO_986 (O_986,N_8637,N_9746);
and UO_987 (O_987,N_8696,N_9263);
and UO_988 (O_988,N_7475,N_8230);
nor UO_989 (O_989,N_7215,N_7486);
nor UO_990 (O_990,N_7261,N_8536);
and UO_991 (O_991,N_6443,N_8200);
and UO_992 (O_992,N_5422,N_5996);
nor UO_993 (O_993,N_8801,N_8422);
nand UO_994 (O_994,N_5241,N_7938);
nand UO_995 (O_995,N_5174,N_8767);
and UO_996 (O_996,N_8510,N_7345);
nand UO_997 (O_997,N_7828,N_5262);
nand UO_998 (O_998,N_7294,N_5625);
and UO_999 (O_999,N_5599,N_7300);
nand UO_1000 (O_1000,N_9149,N_5312);
and UO_1001 (O_1001,N_8447,N_8959);
nand UO_1002 (O_1002,N_6434,N_6843);
and UO_1003 (O_1003,N_6026,N_8810);
nor UO_1004 (O_1004,N_5525,N_5094);
nor UO_1005 (O_1005,N_9681,N_8662);
nand UO_1006 (O_1006,N_6986,N_5474);
nor UO_1007 (O_1007,N_9108,N_5749);
nor UO_1008 (O_1008,N_5936,N_6949);
nand UO_1009 (O_1009,N_8458,N_8161);
nand UO_1010 (O_1010,N_7359,N_7687);
nand UO_1011 (O_1011,N_9445,N_7470);
or UO_1012 (O_1012,N_7670,N_6215);
nor UO_1013 (O_1013,N_7730,N_8300);
nand UO_1014 (O_1014,N_9036,N_6768);
nor UO_1015 (O_1015,N_8164,N_7635);
nand UO_1016 (O_1016,N_9893,N_6345);
and UO_1017 (O_1017,N_6033,N_8687);
nor UO_1018 (O_1018,N_5049,N_8639);
nor UO_1019 (O_1019,N_5690,N_7159);
or UO_1020 (O_1020,N_5977,N_8242);
nand UO_1021 (O_1021,N_7701,N_7405);
or UO_1022 (O_1022,N_7845,N_7130);
nor UO_1023 (O_1023,N_5536,N_6582);
nor UO_1024 (O_1024,N_7320,N_6989);
or UO_1025 (O_1025,N_9401,N_6871);
and UO_1026 (O_1026,N_7954,N_7406);
xnor UO_1027 (O_1027,N_9497,N_8122);
and UO_1028 (O_1028,N_8058,N_7309);
and UO_1029 (O_1029,N_6740,N_7373);
and UO_1030 (O_1030,N_8104,N_5921);
or UO_1031 (O_1031,N_8725,N_8698);
nor UO_1032 (O_1032,N_8989,N_7111);
nand UO_1033 (O_1033,N_6283,N_7720);
and UO_1034 (O_1034,N_8806,N_5236);
or UO_1035 (O_1035,N_6484,N_9146);
nand UO_1036 (O_1036,N_8109,N_5548);
nand UO_1037 (O_1037,N_9275,N_9630);
nor UO_1038 (O_1038,N_9301,N_6868);
or UO_1039 (O_1039,N_7668,N_7199);
nand UO_1040 (O_1040,N_6877,N_7105);
nor UO_1041 (O_1041,N_5755,N_9058);
and UO_1042 (O_1042,N_5741,N_8968);
and UO_1043 (O_1043,N_5369,N_8166);
and UO_1044 (O_1044,N_6821,N_9908);
and UO_1045 (O_1045,N_5041,N_7729);
or UO_1046 (O_1046,N_8472,N_6040);
or UO_1047 (O_1047,N_8379,N_8347);
and UO_1048 (O_1048,N_6259,N_7653);
nand UO_1049 (O_1049,N_9955,N_5326);
and UO_1050 (O_1050,N_5785,N_9337);
and UO_1051 (O_1051,N_8170,N_7927);
nand UO_1052 (O_1052,N_7085,N_9856);
and UO_1053 (O_1053,N_8202,N_9842);
and UO_1054 (O_1054,N_7769,N_5676);
nand UO_1055 (O_1055,N_8442,N_9448);
nand UO_1056 (O_1056,N_6341,N_5920);
nand UO_1057 (O_1057,N_5115,N_9545);
nand UO_1058 (O_1058,N_6874,N_7992);
or UO_1059 (O_1059,N_5489,N_8276);
and UO_1060 (O_1060,N_7814,N_5728);
nand UO_1061 (O_1061,N_9843,N_6783);
or UO_1062 (O_1062,N_6143,N_8998);
or UO_1063 (O_1063,N_8176,N_9322);
and UO_1064 (O_1064,N_6583,N_6019);
nor UO_1065 (O_1065,N_7408,N_6693);
and UO_1066 (O_1066,N_8284,N_7126);
or UO_1067 (O_1067,N_5680,N_6002);
or UO_1068 (O_1068,N_7609,N_6093);
or UO_1069 (O_1069,N_7473,N_8900);
nor UO_1070 (O_1070,N_9048,N_7602);
or UO_1071 (O_1071,N_9755,N_8695);
or UO_1072 (O_1072,N_6904,N_5772);
nor UO_1073 (O_1073,N_5275,N_5135);
or UO_1074 (O_1074,N_5032,N_5413);
nand UO_1075 (O_1075,N_6391,N_9803);
or UO_1076 (O_1076,N_7851,N_7697);
nand UO_1077 (O_1077,N_7911,N_6644);
or UO_1078 (O_1078,N_6270,N_8153);
nand UO_1079 (O_1079,N_6335,N_6565);
and UO_1080 (O_1080,N_6786,N_7872);
nor UO_1081 (O_1081,N_5871,N_7018);
nand UO_1082 (O_1082,N_6934,N_7870);
nor UO_1083 (O_1083,N_9384,N_6923);
and UO_1084 (O_1084,N_7006,N_6657);
nor UO_1085 (O_1085,N_5400,N_7232);
or UO_1086 (O_1086,N_7614,N_6280);
nand UO_1087 (O_1087,N_6626,N_8130);
and UO_1088 (O_1088,N_7448,N_5973);
and UO_1089 (O_1089,N_5267,N_8397);
nand UO_1090 (O_1090,N_6278,N_5420);
or UO_1091 (O_1091,N_7686,N_7772);
nor UO_1092 (O_1092,N_8840,N_6961);
and UO_1093 (O_1093,N_6349,N_5529);
nor UO_1094 (O_1094,N_9761,N_8842);
nor UO_1095 (O_1095,N_9584,N_8688);
and UO_1096 (O_1096,N_7489,N_5695);
and UO_1097 (O_1097,N_5542,N_8636);
and UO_1098 (O_1098,N_5650,N_9719);
and UO_1099 (O_1099,N_7447,N_9618);
nor UO_1100 (O_1100,N_6797,N_7239);
and UO_1101 (O_1101,N_8375,N_9751);
or UO_1102 (O_1102,N_8380,N_8558);
and UO_1103 (O_1103,N_5121,N_9411);
nand UO_1104 (O_1104,N_9521,N_7900);
or UO_1105 (O_1105,N_9621,N_5939);
or UO_1106 (O_1106,N_7454,N_8138);
and UO_1107 (O_1107,N_5399,N_8661);
nand UO_1108 (O_1108,N_7986,N_6281);
nand UO_1109 (O_1109,N_6940,N_9964);
nand UO_1110 (O_1110,N_6537,N_9677);
or UO_1111 (O_1111,N_5092,N_5059);
nor UO_1112 (O_1112,N_9534,N_8210);
nand UO_1113 (O_1113,N_7807,N_9277);
or UO_1114 (O_1114,N_5990,N_5722);
and UO_1115 (O_1115,N_7014,N_8095);
nor UO_1116 (O_1116,N_7010,N_6374);
nand UO_1117 (O_1117,N_6505,N_7893);
xor UO_1118 (O_1118,N_7817,N_6719);
or UO_1119 (O_1119,N_8302,N_8377);
or UO_1120 (O_1120,N_5571,N_6893);
and UO_1121 (O_1121,N_8815,N_9585);
or UO_1122 (O_1122,N_5302,N_5099);
nor UO_1123 (O_1123,N_7230,N_7158);
nor UO_1124 (O_1124,N_5796,N_7943);
or UO_1125 (O_1125,N_8034,N_9362);
nand UO_1126 (O_1126,N_8369,N_6269);
and UO_1127 (O_1127,N_7527,N_6727);
and UO_1128 (O_1128,N_5733,N_5408);
and UO_1129 (O_1129,N_9071,N_6260);
nor UO_1130 (O_1130,N_6629,N_8686);
and UO_1131 (O_1131,N_6307,N_7098);
or UO_1132 (O_1132,N_8156,N_7884);
or UO_1133 (O_1133,N_7680,N_6228);
and UO_1134 (O_1134,N_6638,N_5715);
or UO_1135 (O_1135,N_9237,N_7506);
or UO_1136 (O_1136,N_6572,N_6172);
or UO_1137 (O_1137,N_9024,N_6703);
or UO_1138 (O_1138,N_8580,N_6820);
nor UO_1139 (O_1139,N_9516,N_7930);
nand UO_1140 (O_1140,N_6168,N_7377);
and UO_1141 (O_1141,N_6908,N_6834);
nor UO_1142 (O_1142,N_6387,N_5410);
nor UO_1143 (O_1143,N_6536,N_9089);
and UO_1144 (O_1144,N_6265,N_8206);
and UO_1145 (O_1145,N_5705,N_9541);
nor UO_1146 (O_1146,N_9551,N_5435);
and UO_1147 (O_1147,N_9297,N_7463);
nor UO_1148 (O_1148,N_7656,N_5366);
nor UO_1149 (O_1149,N_6950,N_5344);
or UO_1150 (O_1150,N_9680,N_5640);
nand UO_1151 (O_1151,N_7544,N_6071);
or UO_1152 (O_1152,N_9412,N_7521);
nor UO_1153 (O_1153,N_7258,N_7394);
nor UO_1154 (O_1154,N_6016,N_7761);
or UO_1155 (O_1155,N_9461,N_8027);
nor UO_1156 (O_1156,N_6595,N_7362);
nand UO_1157 (O_1157,N_7389,N_8940);
or UO_1158 (O_1158,N_9582,N_5846);
nand UO_1159 (O_1159,N_5657,N_6972);
and UO_1160 (O_1160,N_7874,N_8190);
and UO_1161 (O_1161,N_7813,N_5666);
nor UO_1162 (O_1162,N_7128,N_7756);
nor UO_1163 (O_1163,N_9380,N_8371);
and UO_1164 (O_1164,N_8548,N_7603);
nor UO_1165 (O_1165,N_9309,N_5843);
nand UO_1166 (O_1166,N_5714,N_7590);
or UO_1167 (O_1167,N_7370,N_8750);
or UO_1168 (O_1168,N_8459,N_9894);
or UO_1169 (O_1169,N_7267,N_7673);
and UO_1170 (O_1170,N_8982,N_6915);
or UO_1171 (O_1171,N_7385,N_7587);
nand UO_1172 (O_1172,N_9554,N_8167);
nand UO_1173 (O_1173,N_8666,N_5537);
nand UO_1174 (O_1174,N_6939,N_6684);
and UO_1175 (O_1175,N_8236,N_7745);
or UO_1176 (O_1176,N_5108,N_5696);
or UO_1177 (O_1177,N_6931,N_9744);
nor UO_1178 (O_1178,N_6339,N_7281);
nand UO_1179 (O_1179,N_9265,N_8826);
nor UO_1180 (O_1180,N_8186,N_9637);
and UO_1181 (O_1181,N_5033,N_5095);
or UO_1182 (O_1182,N_6122,N_6817);
nand UO_1183 (O_1183,N_5402,N_8060);
nand UO_1184 (O_1184,N_9729,N_5613);
and UO_1185 (O_1185,N_6749,N_9957);
nor UO_1186 (O_1186,N_5149,N_9778);
nor UO_1187 (O_1187,N_8692,N_7233);
nor UO_1188 (O_1188,N_9493,N_9150);
nand UO_1189 (O_1189,N_8953,N_9303);
and UO_1190 (O_1190,N_5348,N_8140);
nand UO_1191 (O_1191,N_7009,N_5637);
or UO_1192 (O_1192,N_5991,N_8610);
nand UO_1193 (O_1193,N_6503,N_7461);
and UO_1194 (O_1194,N_8707,N_8221);
nand UO_1195 (O_1195,N_9934,N_6714);
nand UO_1196 (O_1196,N_7114,N_6123);
nor UO_1197 (O_1197,N_5012,N_6160);
and UO_1198 (O_1198,N_9984,N_5947);
or UO_1199 (O_1199,N_5320,N_6347);
nor UO_1200 (O_1200,N_8597,N_8892);
or UO_1201 (O_1201,N_5125,N_5089);
nor UO_1202 (O_1202,N_8285,N_8084);
or UO_1203 (O_1203,N_8450,N_8108);
nand UO_1204 (O_1204,N_6628,N_5626);
xor UO_1205 (O_1205,N_9886,N_9459);
or UO_1206 (O_1206,N_5234,N_5508);
and UO_1207 (O_1207,N_9418,N_5999);
nor UO_1208 (O_1208,N_5634,N_9078);
or UO_1209 (O_1209,N_6129,N_9771);
nand UO_1210 (O_1210,N_5175,N_8349);
or UO_1211 (O_1211,N_7809,N_6326);
and UO_1212 (O_1212,N_5569,N_8017);
and UO_1213 (O_1213,N_7417,N_9059);
nand UO_1214 (O_1214,N_6105,N_9197);
and UO_1215 (O_1215,N_8789,N_9016);
nor UO_1216 (O_1216,N_9610,N_8336);
or UO_1217 (O_1217,N_8051,N_9673);
or UO_1218 (O_1218,N_5103,N_7947);
nor UO_1219 (O_1219,N_6688,N_9496);
nand UO_1220 (O_1220,N_7640,N_9315);
xnor UO_1221 (O_1221,N_9763,N_6983);
or UO_1222 (O_1222,N_5765,N_7768);
or UO_1223 (O_1223,N_5074,N_6256);
or UO_1224 (O_1224,N_8360,N_8520);
xor UO_1225 (O_1225,N_5614,N_7360);
or UO_1226 (O_1226,N_5586,N_5113);
nand UO_1227 (O_1227,N_8059,N_7997);
or UO_1228 (O_1228,N_9774,N_7879);
and UO_1229 (O_1229,N_7837,N_9010);
nand UO_1230 (O_1230,N_7850,N_6411);
nand UO_1231 (O_1231,N_7810,N_7998);
or UO_1232 (O_1232,N_5064,N_5195);
nand UO_1233 (O_1233,N_5558,N_7882);
or UO_1234 (O_1234,N_9920,N_6053);
or UO_1235 (O_1235,N_6022,N_8054);
nor UO_1236 (O_1236,N_5859,N_6180);
nor UO_1237 (O_1237,N_9661,N_9626);
or UO_1238 (O_1238,N_7122,N_7854);
nand UO_1239 (O_1239,N_8823,N_5831);
nand UO_1240 (O_1240,N_8567,N_6920);
nor UO_1241 (O_1241,N_6361,N_9074);
and UO_1242 (O_1242,N_6602,N_8326);
nor UO_1243 (O_1243,N_5013,N_6530);
and UO_1244 (O_1244,N_9009,N_6043);
and UO_1245 (O_1245,N_7762,N_6194);
and UO_1246 (O_1246,N_7780,N_8581);
and UO_1247 (O_1247,N_9105,N_8334);
nand UO_1248 (O_1248,N_7528,N_7957);
and UO_1249 (O_1249,N_6909,N_5243);
nor UO_1250 (O_1250,N_5165,N_8785);
nor UO_1251 (O_1251,N_5182,N_7282);
and UO_1252 (O_1252,N_5073,N_6586);
nand UO_1253 (O_1253,N_7819,N_8701);
and UO_1254 (O_1254,N_5003,N_5795);
or UO_1255 (O_1255,N_6303,N_6991);
or UO_1256 (O_1256,N_7113,N_7618);
nor UO_1257 (O_1257,N_5834,N_6579);
and UO_1258 (O_1258,N_7584,N_8483);
nand UO_1259 (O_1259,N_9368,N_7190);
and UO_1260 (O_1260,N_6049,N_8007);
nor UO_1261 (O_1261,N_6735,N_8985);
nand UO_1262 (O_1262,N_6992,N_5916);
nor UO_1263 (O_1263,N_6396,N_9936);
and UO_1264 (O_1264,N_5627,N_7862);
or UO_1265 (O_1265,N_8049,N_6420);
and UO_1266 (O_1266,N_9558,N_9285);
or UO_1267 (O_1267,N_7150,N_6833);
nand UO_1268 (O_1268,N_6421,N_8293);
nor UO_1269 (O_1269,N_5531,N_8274);
or UO_1270 (O_1270,N_7538,N_8179);
or UO_1271 (O_1271,N_6248,N_9879);
or UO_1272 (O_1272,N_9460,N_6197);
nand UO_1273 (O_1273,N_7829,N_5716);
nand UO_1274 (O_1274,N_9814,N_6183);
and UO_1275 (O_1275,N_5610,N_6359);
nand UO_1276 (O_1276,N_6092,N_5863);
or UO_1277 (O_1277,N_6675,N_8389);
nor UO_1278 (O_1278,N_6161,N_9711);
nand UO_1279 (O_1279,N_7842,N_9311);
and UO_1280 (O_1280,N_9407,N_9884);
nor UO_1281 (O_1281,N_8830,N_6664);
or UO_1282 (O_1282,N_9564,N_8313);
nand UO_1283 (O_1283,N_6804,N_9350);
nor UO_1284 (O_1284,N_7355,N_5387);
nand UO_1285 (O_1285,N_9132,N_9218);
and UO_1286 (O_1286,N_6477,N_5759);
or UO_1287 (O_1287,N_9902,N_6605);
nor UO_1288 (O_1288,N_7777,N_9189);
nor UO_1289 (O_1289,N_6510,N_9019);
or UO_1290 (O_1290,N_6464,N_6640);
or UO_1291 (O_1291,N_8288,N_9979);
and UO_1292 (O_1292,N_8014,N_9247);
and UO_1293 (O_1293,N_7000,N_6591);
or UO_1294 (O_1294,N_5888,N_9027);
nor UO_1295 (O_1295,N_9116,N_5751);
and UO_1296 (O_1296,N_5453,N_6544);
and UO_1297 (O_1297,N_7896,N_6491);
and UO_1298 (O_1298,N_5849,N_8157);
and UO_1299 (O_1299,N_8507,N_7648);
and UO_1300 (O_1300,N_9002,N_7523);
or UO_1301 (O_1301,N_7332,N_9215);
and UO_1302 (O_1302,N_9087,N_9752);
or UO_1303 (O_1303,N_5713,N_6184);
nand UO_1304 (O_1304,N_7728,N_7574);
nand UO_1305 (O_1305,N_9773,N_8297);
nand UO_1306 (O_1306,N_7647,N_9241);
or UO_1307 (O_1307,N_6619,N_6718);
and UO_1308 (O_1308,N_7526,N_8469);
and UO_1309 (O_1309,N_7492,N_9978);
or UO_1310 (O_1310,N_7627,N_8304);
and UO_1311 (O_1311,N_9079,N_8627);
nand UO_1312 (O_1312,N_5621,N_7898);
and UO_1313 (O_1313,N_9930,N_5449);
or UO_1314 (O_1314,N_5324,N_5321);
nor UO_1315 (O_1315,N_6955,N_8233);
and UO_1316 (O_1316,N_8761,N_7179);
nor UO_1317 (O_1317,N_6880,N_7876);
and UO_1318 (O_1318,N_5322,N_9183);
or UO_1319 (O_1319,N_7375,N_8811);
nor UO_1320 (O_1320,N_8211,N_8575);
and UO_1321 (O_1321,N_5171,N_9456);
nor UO_1322 (O_1322,N_6615,N_5030);
nor UO_1323 (O_1323,N_5301,N_9789);
and UO_1324 (O_1324,N_6368,N_9528);
nor UO_1325 (O_1325,N_5539,N_5035);
or UO_1326 (O_1326,N_6013,N_7905);
nand UO_1327 (O_1327,N_9186,N_6734);
nand UO_1328 (O_1328,N_5186,N_8640);
nand UO_1329 (O_1329,N_5724,N_7805);
nand UO_1330 (O_1330,N_8792,N_9671);
nand UO_1331 (O_1331,N_8081,N_6333);
nor UO_1332 (O_1332,N_7712,N_5823);
or UO_1333 (O_1333,N_7832,N_5211);
nor UO_1334 (O_1334,N_6486,N_9703);
and UO_1335 (O_1335,N_8800,N_5323);
and UO_1336 (O_1336,N_6867,N_9238);
nand UO_1337 (O_1337,N_8496,N_7015);
and UO_1338 (O_1338,N_5588,N_9634);
or UO_1339 (O_1339,N_9427,N_7234);
or UO_1340 (O_1340,N_6007,N_8858);
nor UO_1341 (O_1341,N_6754,N_9740);
and UO_1342 (O_1342,N_9417,N_9225);
nand UO_1343 (O_1343,N_9670,N_7784);
and UO_1344 (O_1344,N_8136,N_5319);
or UO_1345 (O_1345,N_7033,N_6148);
nor UO_1346 (O_1346,N_8845,N_5969);
or UO_1347 (O_1347,N_5560,N_8468);
nor UO_1348 (O_1348,N_5691,N_9298);
and UO_1349 (O_1349,N_5872,N_8038);
or UO_1350 (O_1350,N_8867,N_7279);
and UO_1351 (O_1351,N_7319,N_8915);
and UO_1352 (O_1352,N_6208,N_9117);
nor UO_1353 (O_1353,N_8261,N_7482);
or UO_1354 (O_1354,N_6913,N_7374);
nand UO_1355 (O_1355,N_5612,N_8532);
and UO_1356 (O_1356,N_8244,N_7568);
nand UO_1357 (O_1357,N_5356,N_6078);
and UO_1358 (O_1358,N_8492,N_9657);
nand UO_1359 (O_1359,N_9148,N_8904);
and UO_1360 (O_1360,N_8672,N_8626);
and UO_1361 (O_1361,N_7022,N_9968);
and UO_1362 (O_1362,N_6138,N_6933);
and UO_1363 (O_1363,N_5036,N_5139);
nand UO_1364 (O_1364,N_7001,N_8596);
nor UO_1365 (O_1365,N_5918,N_9403);
or UO_1366 (O_1366,N_9370,N_6720);
nand UO_1367 (O_1367,N_6055,N_8439);
or UO_1368 (O_1368,N_5615,N_5968);
and UO_1369 (O_1369,N_6395,N_8956);
or UO_1370 (O_1370,N_8868,N_5707);
nand UO_1371 (O_1371,N_5488,N_9056);
nor UO_1372 (O_1372,N_5576,N_9307);
or UO_1373 (O_1373,N_8456,N_8561);
nand UO_1374 (O_1374,N_9858,N_9131);
nand UO_1375 (O_1375,N_5276,N_8546);
and UO_1376 (O_1376,N_7726,N_9961);
nand UO_1377 (O_1377,N_7125,N_6192);
and UO_1378 (O_1378,N_9174,N_9152);
nand UO_1379 (O_1379,N_6694,N_9454);
nand UO_1380 (O_1380,N_7265,N_6340);
nor UO_1381 (O_1381,N_5384,N_5308);
and UO_1382 (O_1382,N_9003,N_8455);
nor UO_1383 (O_1383,N_9220,N_6000);
and UO_1384 (O_1384,N_9759,N_6445);
and UO_1385 (O_1385,N_6882,N_9708);
nor UO_1386 (O_1386,N_6730,N_9125);
nor UO_1387 (O_1387,N_7428,N_7550);
and UO_1388 (O_1388,N_9536,N_9713);
nand UO_1389 (O_1389,N_7342,N_8844);
nand UO_1390 (O_1390,N_5447,N_8623);
nor UO_1391 (O_1391,N_9190,N_6562);
nand UO_1392 (O_1392,N_9354,N_9649);
xnor UO_1393 (O_1393,N_7131,N_6781);
and UO_1394 (O_1394,N_5193,N_8765);
nand UO_1395 (O_1395,N_8168,N_8196);
nand UO_1396 (O_1396,N_8454,N_9870);
and UO_1397 (O_1397,N_9865,N_9777);
nor UO_1398 (O_1398,N_6028,N_7760);
and UO_1399 (O_1399,N_6620,N_9507);
nor UO_1400 (O_1400,N_8488,N_9818);
or UO_1401 (O_1401,N_6509,N_6606);
nand UO_1402 (O_1402,N_5504,N_9710);
nand UO_1403 (O_1403,N_5462,N_6981);
or UO_1404 (O_1404,N_5669,N_8254);
and UO_1405 (O_1405,N_7682,N_7891);
or UO_1406 (O_1406,N_5810,N_8494);
nand UO_1407 (O_1407,N_8604,N_7145);
and UO_1408 (O_1408,N_9636,N_7719);
nor UO_1409 (O_1409,N_9903,N_9193);
and UO_1410 (O_1410,N_5667,N_7079);
nand UO_1411 (O_1411,N_8859,N_6765);
and UO_1412 (O_1412,N_5580,N_8747);
nand UO_1413 (O_1413,N_7600,N_6317);
nand UO_1414 (O_1414,N_9715,N_9093);
and UO_1415 (O_1415,N_5516,N_7530);
xor UO_1416 (O_1416,N_8421,N_8227);
nor UO_1417 (O_1417,N_7301,N_5386);
and UO_1418 (O_1418,N_7983,N_5505);
nand UO_1419 (O_1419,N_7974,N_7161);
or UO_1420 (O_1420,N_6818,N_9690);
and UO_1421 (O_1421,N_9338,N_8374);
nand UO_1422 (O_1422,N_5904,N_9915);
or UO_1423 (O_1423,N_8082,N_8681);
or UO_1424 (O_1424,N_5450,N_5604);
or UO_1425 (O_1425,N_8676,N_8436);
nand UO_1426 (O_1426,N_6147,N_7025);
nand UO_1427 (O_1427,N_9217,N_8914);
nor UO_1428 (O_1428,N_6570,N_5568);
or UO_1429 (O_1429,N_6490,N_5807);
nor UO_1430 (O_1430,N_5225,N_8566);
or UO_1431 (O_1431,N_5600,N_9748);
or UO_1432 (O_1432,N_5825,N_8289);
and UO_1433 (O_1433,N_8493,N_7424);
or UO_1434 (O_1434,N_5697,N_7993);
nand UO_1435 (O_1435,N_8325,N_7941);
nor UO_1436 (O_1436,N_9632,N_7823);
nor UO_1437 (O_1437,N_7912,N_8097);
xor UO_1438 (O_1438,N_8438,N_6851);
and UO_1439 (O_1439,N_8018,N_5583);
nor UO_1440 (O_1440,N_9641,N_5072);
nor UO_1441 (O_1441,N_7270,N_5824);
xor UO_1442 (O_1442,N_5544,N_8731);
and UO_1443 (O_1443,N_9590,N_6142);
nand UO_1444 (O_1444,N_9441,N_5500);
nor UO_1445 (O_1445,N_7186,N_9406);
nor UO_1446 (O_1446,N_9169,N_8041);
and UO_1447 (O_1447,N_6175,N_5514);
and UO_1448 (O_1448,N_6661,N_7763);
nor UO_1449 (O_1449,N_5286,N_6962);
xnor UO_1450 (O_1450,N_8173,N_7142);
and UO_1451 (O_1451,N_7717,N_7432);
nand UO_1452 (O_1452,N_7519,N_8258);
or UO_1453 (O_1453,N_7029,N_8388);
nor UO_1454 (O_1454,N_9336,N_8272);
nor UO_1455 (O_1455,N_7402,N_9642);
nor UO_1456 (O_1456,N_5010,N_5957);
or UO_1457 (O_1457,N_6850,N_5282);
nor UO_1458 (O_1458,N_9214,N_8396);
and UO_1459 (O_1459,N_9583,N_8778);
and UO_1460 (O_1460,N_5729,N_6456);
nand UO_1461 (O_1461,N_7737,N_9327);
and UO_1462 (O_1462,N_8024,N_8835);
nand UO_1463 (O_1463,N_7920,N_7246);
and UO_1464 (O_1464,N_5470,N_9900);
or UO_1465 (O_1465,N_9118,N_9745);
and UO_1466 (O_1466,N_9669,N_6575);
or UO_1467 (O_1467,N_7487,N_8000);
or UO_1468 (O_1468,N_5646,N_6254);
nand UO_1469 (O_1469,N_5248,N_9739);
nor UO_1470 (O_1470,N_9279,N_9723);
nor UO_1471 (O_1471,N_9918,N_6907);
or UO_1472 (O_1472,N_8194,N_6189);
nand UO_1473 (O_1473,N_7398,N_5427);
nand UO_1474 (O_1474,N_7361,N_5665);
or UO_1475 (O_1475,N_7343,N_9038);
nand UO_1476 (O_1476,N_8056,N_8906);
nor UO_1477 (O_1477,N_6218,N_9960);
nor UO_1478 (O_1478,N_8514,N_8105);
nor UO_1479 (O_1479,N_9686,N_6364);
nand UO_1480 (O_1480,N_7140,N_9293);
nor UO_1481 (O_1481,N_9917,N_8355);
and UO_1482 (O_1482,N_5706,N_8773);
nor UO_1483 (O_1483,N_6383,N_5938);
or UO_1484 (O_1484,N_8207,N_9447);
or UO_1485 (O_1485,N_8878,N_8474);
or UO_1486 (O_1486,N_6671,N_6212);
nand UO_1487 (O_1487,N_5975,N_7906);
nand UO_1488 (O_1488,N_5285,N_7666);
nor UO_1489 (O_1489,N_6884,N_8682);
nor UO_1490 (O_1490,N_9613,N_6800);
nor UO_1491 (O_1491,N_6513,N_5821);
nand UO_1492 (O_1492,N_9648,N_6213);
nand UO_1493 (O_1493,N_8743,N_5445);
nand UO_1494 (O_1494,N_8656,N_9053);
or UO_1495 (O_1495,N_8653,N_8085);
or UO_1496 (O_1496,N_9736,N_8957);
or UO_1497 (O_1497,N_9022,N_5683);
or UO_1498 (O_1498,N_6889,N_6334);
xor UO_1499 (O_1499,N_7942,N_7437);
endmodule