module basic_2000_20000_2500_4_levels_5xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
nor U0 (N_0,In_796,In_731);
nand U1 (N_1,In_172,In_1343);
and U2 (N_2,In_390,In_946);
and U3 (N_3,In_1144,In_65);
and U4 (N_4,In_721,In_950);
and U5 (N_5,In_867,In_1029);
nand U6 (N_6,In_815,In_1862);
or U7 (N_7,In_1026,In_1466);
nand U8 (N_8,In_26,In_962);
and U9 (N_9,In_52,In_1666);
or U10 (N_10,In_368,In_677);
nor U11 (N_11,In_1967,In_580);
and U12 (N_12,In_215,In_318);
and U13 (N_13,In_596,In_736);
nor U14 (N_14,In_489,In_901);
and U15 (N_15,In_1519,In_1965);
nor U16 (N_16,In_177,In_937);
or U17 (N_17,In_16,In_196);
and U18 (N_18,In_1152,In_192);
nand U19 (N_19,In_926,In_919);
and U20 (N_20,In_1512,In_1728);
nor U21 (N_21,In_133,In_1312);
or U22 (N_22,In_1940,In_233);
nor U23 (N_23,In_1602,In_746);
nor U24 (N_24,In_1897,In_1799);
and U25 (N_25,In_1402,In_1219);
and U26 (N_26,In_406,In_13);
nor U27 (N_27,In_1808,In_420);
nor U28 (N_28,In_612,In_1982);
or U29 (N_29,In_1290,In_1615);
or U30 (N_30,In_1114,In_1420);
xnor U31 (N_31,In_491,In_747);
nor U32 (N_32,In_1522,In_1950);
nor U33 (N_33,In_1568,In_1687);
xor U34 (N_34,In_751,In_112);
and U35 (N_35,In_487,In_31);
xnor U36 (N_36,In_1451,In_391);
and U37 (N_37,In_73,In_1651);
nand U38 (N_38,In_1720,In_713);
or U39 (N_39,In_1056,In_1741);
or U40 (N_40,In_269,In_1831);
nor U41 (N_41,In_1887,In_1159);
nand U42 (N_42,In_1815,In_602);
nor U43 (N_43,In_735,In_1949);
nand U44 (N_44,In_1059,In_241);
xnor U45 (N_45,In_495,In_1279);
and U46 (N_46,In_1623,In_170);
and U47 (N_47,In_1205,In_705);
nor U48 (N_48,In_1300,In_323);
or U49 (N_49,In_1679,In_1721);
or U50 (N_50,In_1012,In_1776);
nand U51 (N_51,In_1994,In_182);
and U52 (N_52,In_753,In_1302);
and U53 (N_53,In_1662,In_733);
xnor U54 (N_54,In_128,In_1491);
and U55 (N_55,In_862,In_1080);
or U56 (N_56,In_1200,In_1525);
nand U57 (N_57,In_299,In_1754);
nor U58 (N_58,In_165,In_1415);
nand U59 (N_59,In_1696,In_800);
nor U60 (N_60,In_82,In_873);
nand U61 (N_61,In_517,In_1806);
nand U62 (N_62,In_151,In_187);
nand U63 (N_63,In_22,In_1939);
nand U64 (N_64,In_895,In_571);
nor U65 (N_65,In_1468,In_1683);
xnor U66 (N_66,In_864,In_1021);
and U67 (N_67,In_1820,In_1546);
nor U68 (N_68,In_174,In_1524);
and U69 (N_69,In_3,In_680);
nand U70 (N_70,In_147,In_1295);
nand U71 (N_71,In_849,In_667);
nand U72 (N_72,In_1090,In_441);
nor U73 (N_73,In_989,In_971);
xor U74 (N_74,In_1296,In_767);
nor U75 (N_75,In_450,In_1108);
xor U76 (N_76,In_141,In_395);
nand U77 (N_77,In_486,In_1654);
and U78 (N_78,In_1660,In_587);
nor U79 (N_79,In_1231,In_1819);
and U80 (N_80,In_481,In_1401);
or U81 (N_81,In_1510,In_1341);
nand U82 (N_82,In_1122,In_286);
nor U83 (N_83,In_1562,In_214);
or U84 (N_84,In_1680,In_1585);
or U85 (N_85,In_329,In_1945);
or U86 (N_86,In_913,In_925);
or U87 (N_87,In_1607,In_1639);
or U88 (N_88,In_1237,In_1304);
nor U89 (N_89,In_1533,In_1576);
and U90 (N_90,In_1476,In_980);
nor U91 (N_91,In_319,In_514);
and U92 (N_92,In_1907,In_790);
and U93 (N_93,In_993,In_1277);
nor U94 (N_94,In_1655,In_1880);
or U95 (N_95,In_912,In_1398);
nand U96 (N_96,In_774,In_1065);
nand U97 (N_97,In_723,In_1204);
and U98 (N_98,In_1482,In_1860);
nand U99 (N_99,In_42,In_1619);
or U100 (N_100,In_288,In_1271);
nand U101 (N_101,In_1315,In_186);
nand U102 (N_102,In_876,In_675);
nand U103 (N_103,In_1857,In_786);
nor U104 (N_104,In_1280,In_34);
or U105 (N_105,In_1483,In_1192);
nor U106 (N_106,In_1578,In_1264);
nand U107 (N_107,In_1076,In_358);
nor U108 (N_108,In_827,In_2);
nand U109 (N_109,In_1354,In_274);
or U110 (N_110,In_1650,In_683);
or U111 (N_111,In_615,In_503);
and U112 (N_112,In_1394,In_1143);
and U113 (N_113,In_1210,In_454);
and U114 (N_114,In_1325,In_1281);
or U115 (N_115,In_700,In_1778);
nor U116 (N_116,In_1698,In_1125);
nor U117 (N_117,In_1837,In_1485);
nor U118 (N_118,In_651,In_673);
and U119 (N_119,In_1384,In_1591);
and U120 (N_120,In_1901,In_1196);
and U121 (N_121,In_1046,In_1409);
and U122 (N_122,In_1891,In_1183);
and U123 (N_123,In_243,In_403);
xnor U124 (N_124,In_351,In_33);
and U125 (N_125,In_892,In_1288);
and U126 (N_126,In_750,In_419);
xnor U127 (N_127,In_88,In_664);
nor U128 (N_128,In_55,In_917);
nand U129 (N_129,In_1479,In_510);
and U130 (N_130,In_1003,In_1750);
or U131 (N_131,In_1189,In_1207);
and U132 (N_132,In_1034,In_1771);
or U133 (N_133,In_1243,In_600);
or U134 (N_134,In_992,In_1570);
or U135 (N_135,In_860,In_113);
and U136 (N_136,In_1433,In_375);
and U137 (N_137,In_1043,In_1274);
or U138 (N_138,In_1774,In_327);
nor U139 (N_139,In_986,In_1717);
xnor U140 (N_140,In_622,In_671);
or U141 (N_141,In_1282,In_1853);
or U142 (N_142,In_979,In_1472);
nand U143 (N_143,In_300,In_1141);
or U144 (N_144,In_843,In_447);
nand U145 (N_145,In_807,In_1814);
and U146 (N_146,In_437,In_140);
nor U147 (N_147,In_702,In_1805);
and U148 (N_148,In_1250,In_1782);
and U149 (N_149,In_674,In_1058);
nand U150 (N_150,In_291,In_1993);
or U151 (N_151,In_1648,In_1121);
and U152 (N_152,In_131,In_1405);
xor U153 (N_153,In_949,In_1574);
or U154 (N_154,In_1344,In_759);
and U155 (N_155,In_648,In_1583);
and U156 (N_156,In_234,In_367);
nor U157 (N_157,In_1381,In_888);
and U158 (N_158,In_1987,In_332);
and U159 (N_159,In_1064,In_1766);
xnor U160 (N_160,In_1133,In_1010);
xor U161 (N_161,In_1202,In_1240);
and U162 (N_162,In_1278,In_479);
nor U163 (N_163,In_194,In_1035);
xnor U164 (N_164,In_1084,In_104);
nand U165 (N_165,In_1167,In_222);
or U166 (N_166,In_1112,In_1763);
nand U167 (N_167,In_1361,In_883);
nand U168 (N_168,In_259,In_1719);
nand U169 (N_169,In_1475,In_1177);
nor U170 (N_170,In_1935,In_1115);
or U171 (N_171,In_282,In_1262);
xnor U172 (N_172,In_740,In_427);
or U173 (N_173,In_1735,In_1587);
and U174 (N_174,In_1917,In_833);
nor U175 (N_175,In_292,In_1375);
nand U176 (N_176,In_1732,In_1872);
or U177 (N_177,In_1626,In_1486);
xnor U178 (N_178,In_810,In_1577);
nor U179 (N_179,In_1608,In_579);
xor U180 (N_180,In_1740,In_1111);
and U181 (N_181,In_822,In_1136);
nand U182 (N_182,In_445,In_1028);
or U183 (N_183,In_1975,In_439);
and U184 (N_184,In_1895,In_1388);
nor U185 (N_185,In_953,In_1647);
or U186 (N_186,In_1633,In_1553);
or U187 (N_187,In_127,In_59);
nand U188 (N_188,In_1446,In_1671);
or U189 (N_189,In_689,In_556);
or U190 (N_190,In_1147,In_1865);
and U191 (N_191,In_394,In_1850);
and U192 (N_192,In_118,In_1423);
nor U193 (N_193,In_739,In_676);
nor U194 (N_194,In_1670,In_1470);
nand U195 (N_195,In_698,In_1211);
or U196 (N_196,In_175,In_696);
and U197 (N_197,In_30,In_1727);
or U198 (N_198,In_95,In_1223);
nor U199 (N_199,In_477,In_1554);
nand U200 (N_200,In_1033,In_820);
nand U201 (N_201,In_263,In_1802);
and U202 (N_202,In_1984,In_398);
and U203 (N_203,In_1270,In_1188);
and U204 (N_204,In_326,In_1724);
and U205 (N_205,In_1532,In_1438);
nor U206 (N_206,In_832,In_1225);
and U207 (N_207,In_123,In_737);
and U208 (N_208,In_195,In_10);
and U209 (N_209,In_471,In_1611);
and U210 (N_210,In_435,In_158);
nand U211 (N_211,In_1057,In_628);
nor U212 (N_212,In_541,In_1378);
nand U213 (N_213,In_262,In_1503);
nand U214 (N_214,In_200,In_1508);
nor U215 (N_215,In_500,In_1879);
or U216 (N_216,In_1756,In_38);
nand U217 (N_217,In_1582,In_1991);
and U218 (N_218,In_738,In_1916);
nand U219 (N_219,In_1008,In_799);
or U220 (N_220,In_1962,In_900);
nor U221 (N_221,In_1822,In_887);
and U222 (N_222,In_1934,In_159);
nor U223 (N_223,In_732,In_442);
nor U224 (N_224,In_1170,In_492);
and U225 (N_225,In_1074,In_1933);
nor U226 (N_226,In_654,In_1215);
nand U227 (N_227,In_775,In_787);
nor U228 (N_228,In_101,In_388);
and U229 (N_229,In_1429,In_585);
and U230 (N_230,In_794,In_1002);
xor U231 (N_231,In_826,In_1359);
or U232 (N_232,In_252,In_754);
nand U233 (N_233,In_577,In_1197);
or U234 (N_234,In_1997,In_1142);
or U235 (N_235,In_1807,In_1382);
nor U236 (N_236,In_1408,In_1017);
and U237 (N_237,In_611,In_1908);
and U238 (N_238,In_1921,In_1406);
and U239 (N_239,In_1529,In_1703);
xor U240 (N_240,In_1365,In_119);
and U241 (N_241,In_429,In_934);
nor U242 (N_242,In_861,In_1314);
nor U243 (N_243,In_1567,In_1713);
nand U244 (N_244,In_1928,In_51);
xor U245 (N_245,In_1927,In_426);
and U246 (N_246,In_988,In_385);
or U247 (N_247,In_1640,In_217);
and U248 (N_248,In_1337,In_576);
and U249 (N_249,In_434,In_226);
or U250 (N_250,In_261,In_1878);
nor U251 (N_251,In_1168,In_761);
or U252 (N_252,In_1863,In_562);
or U253 (N_253,In_637,In_1464);
nand U254 (N_254,In_1998,In_812);
nor U255 (N_255,In_1909,In_566);
nand U256 (N_256,In_478,In_672);
nand U257 (N_257,In_1851,In_1494);
nor U258 (N_258,In_582,In_1481);
nor U259 (N_259,In_14,In_1877);
or U260 (N_260,In_610,In_1442);
nor U261 (N_261,In_595,In_60);
and U262 (N_262,In_574,In_890);
nor U263 (N_263,In_185,In_1787);
and U264 (N_264,In_1081,In_678);
nand U265 (N_265,In_1768,In_268);
nand U266 (N_266,In_1521,In_1595);
nor U267 (N_267,In_115,In_1417);
and U268 (N_268,In_1009,In_885);
and U269 (N_269,In_1004,In_1929);
nor U270 (N_270,In_45,In_758);
nor U271 (N_271,In_161,In_1022);
nor U272 (N_272,In_197,In_1617);
nor U273 (N_273,In_117,In_805);
or U274 (N_274,In_1552,In_1005);
nor U275 (N_275,In_1664,In_449);
and U276 (N_276,In_1313,In_1463);
nor U277 (N_277,In_945,In_1007);
nor U278 (N_278,In_1234,In_1955);
nor U279 (N_279,In_1943,In_982);
nor U280 (N_280,In_1449,In_1160);
and U281 (N_281,In_1723,In_1212);
nand U282 (N_282,In_920,In_711);
nand U283 (N_283,In_125,In_103);
or U284 (N_284,In_1625,In_802);
xnor U285 (N_285,In_225,In_1888);
nor U286 (N_286,In_636,In_1931);
nor U287 (N_287,In_981,In_246);
or U288 (N_288,In_1627,In_164);
nor U289 (N_289,In_1705,In_136);
nor U290 (N_290,In_1099,In_1985);
or U291 (N_291,In_474,In_18);
and U292 (N_292,In_278,In_1707);
and U293 (N_293,In_1657,In_266);
or U294 (N_294,In_1674,In_1572);
and U295 (N_295,In_922,In_967);
and U296 (N_296,In_1153,In_545);
nand U297 (N_297,In_586,In_961);
or U298 (N_298,In_938,In_1801);
nand U299 (N_299,In_1593,In_1624);
and U300 (N_300,In_995,In_1612);
and U301 (N_301,In_1628,In_310);
or U302 (N_302,In_814,In_276);
nor U303 (N_303,In_287,In_592);
and U304 (N_304,In_1961,In_1914);
nand U305 (N_305,In_190,In_384);
or U306 (N_306,In_516,In_293);
nand U307 (N_307,In_819,In_1493);
or U308 (N_308,In_1247,In_604);
nor U309 (N_309,In_1156,In_53);
nor U310 (N_310,In_712,In_728);
nor U311 (N_311,In_1286,In_789);
nand U312 (N_312,In_563,In_1362);
nand U313 (N_313,In_1104,In_144);
or U314 (N_314,In_1739,In_1765);
and U315 (N_315,In_455,In_157);
and U316 (N_316,In_339,In_605);
or U317 (N_317,In_526,In_1445);
xnor U318 (N_318,In_1643,In_829);
nand U319 (N_319,In_212,In_1387);
or U320 (N_320,In_373,In_1905);
and U321 (N_321,In_1902,In_1659);
xor U322 (N_322,In_251,In_1255);
nor U323 (N_323,In_1500,In_844);
or U324 (N_324,In_353,In_518);
and U325 (N_325,In_330,In_681);
and U326 (N_326,In_1380,In_496);
or U327 (N_327,In_974,In_188);
nand U328 (N_328,In_1890,In_86);
nor U329 (N_329,In_1435,In_1180);
or U330 (N_330,In_1839,In_943);
and U331 (N_331,In_824,In_1060);
or U332 (N_332,In_1328,In_1944);
or U333 (N_333,In_1709,In_208);
nor U334 (N_334,In_1474,In_1373);
or U335 (N_335,In_464,In_813);
nand U336 (N_336,In_1040,In_1963);
or U337 (N_337,In_71,In_865);
xnor U338 (N_338,In_572,In_1812);
or U339 (N_339,In_1516,In_1867);
xnor U340 (N_340,In_1498,In_244);
or U341 (N_341,In_325,In_1742);
nand U342 (N_342,In_532,In_1427);
or U343 (N_343,In_975,In_825);
and U344 (N_344,In_19,In_1922);
nor U345 (N_345,In_418,In_583);
and U346 (N_346,In_1652,In_1020);
nor U347 (N_347,In_1886,In_265);
nand U348 (N_348,In_996,In_1140);
or U349 (N_349,In_1261,In_1560);
and U350 (N_350,In_923,In_46);
xnor U351 (N_351,In_1118,In_506);
or U352 (N_352,In_590,In_1575);
and U353 (N_353,In_156,In_472);
or U354 (N_354,In_773,In_1258);
nand U355 (N_355,In_1199,In_780);
and U356 (N_356,In_238,In_1273);
and U357 (N_357,In_1360,In_284);
xnor U358 (N_358,In_1798,In_97);
or U359 (N_359,In_1722,In_1695);
nor U360 (N_360,In_224,In_954);
nor U361 (N_361,In_1335,In_1214);
xnor U362 (N_362,In_765,In_443);
nand U363 (N_363,In_303,In_1644);
nor U364 (N_364,In_1638,In_535);
xor U365 (N_365,In_617,In_357);
nand U366 (N_366,In_361,In_1884);
or U367 (N_367,In_584,In_539);
xnor U368 (N_368,In_1072,In_1747);
xnor U369 (N_369,In_1980,In_473);
nand U370 (N_370,In_924,In_1792);
and U371 (N_371,In_89,In_321);
and U372 (N_372,In_1299,In_875);
and U373 (N_373,In_66,In_1269);
nor U374 (N_374,In_853,In_1697);
or U375 (N_375,In_1996,In_1598);
nand U376 (N_376,In_591,In_550);
nor U377 (N_377,In_1368,In_757);
nor U378 (N_378,In_1811,In_27);
or U379 (N_379,In_1127,In_1777);
or U380 (N_380,In_1293,In_614);
nand U381 (N_381,In_1356,In_257);
xnor U382 (N_382,In_227,In_868);
nand U383 (N_383,In_1253,In_1176);
nand U384 (N_384,In_1032,In_1403);
nand U385 (N_385,In_1773,In_24);
nor U386 (N_386,In_482,In_564);
nand U387 (N_387,In_178,In_855);
nand U388 (N_388,In_1690,In_1559);
xor U389 (N_389,In_84,In_697);
and U390 (N_390,In_1013,In_1761);
and U391 (N_391,In_1653,In_1414);
and U392 (N_392,In_626,In_1845);
xor U393 (N_393,In_494,In_499);
or U394 (N_394,In_1049,In_768);
or U395 (N_395,In_100,In_551);
and U396 (N_396,In_240,In_4);
and U397 (N_397,In_189,In_1370);
nand U398 (N_398,In_124,In_163);
nor U399 (N_399,In_856,In_841);
xor U400 (N_400,In_1637,In_1283);
and U401 (N_401,In_1338,In_1689);
nand U402 (N_402,In_703,In_891);
nand U403 (N_403,In_1999,In_1241);
nor U404 (N_404,In_997,In_126);
or U405 (N_405,In_1131,In_415);
nor U406 (N_406,In_304,In_315);
nand U407 (N_407,In_169,In_905);
or U408 (N_408,In_1110,In_307);
nor U409 (N_409,In_1209,In_1119);
or U410 (N_410,In_817,In_1327);
nand U411 (N_411,In_1301,In_154);
nand U412 (N_412,In_1106,In_1342);
and U413 (N_413,In_594,In_70);
or U414 (N_414,In_1622,In_1107);
nor U415 (N_415,In_1620,In_521);
or U416 (N_416,In_1454,In_397);
and U417 (N_417,In_1097,In_1855);
nand U418 (N_418,In_1006,In_29);
or U419 (N_419,In_609,In_655);
nand U420 (N_420,In_897,In_1050);
nor U421 (N_421,In_1227,In_834);
and U422 (N_422,In_1775,In_15);
xnor U423 (N_423,In_249,In_1609);
nand U424 (N_424,In_1473,In_277);
and U425 (N_425,In_1055,In_1336);
nor U426 (N_426,In_1549,In_1413);
and U427 (N_427,In_272,In_523);
nor U428 (N_428,In_206,In_598);
and U429 (N_429,In_722,In_618);
nand U430 (N_430,In_546,In_1564);
xnor U431 (N_431,In_1919,In_138);
nor U432 (N_432,In_665,In_509);
nor U433 (N_433,In_312,In_1903);
xnor U434 (N_434,In_1488,In_1610);
nand U435 (N_435,In_1162,In_1715);
nor U436 (N_436,In_1244,In_1489);
or U437 (N_437,In_1018,In_520);
nand U438 (N_438,In_1100,In_578);
nor U439 (N_439,In_633,In_1936);
xor U440 (N_440,In_1986,In_769);
nand U441 (N_441,In_1230,In_424);
and U442 (N_442,In_1706,In_425);
and U443 (N_443,In_297,In_806);
nor U444 (N_444,In_305,In_719);
nand U445 (N_445,In_1171,In_1673);
or U446 (N_446,In_1421,In_531);
nor U447 (N_447,In_1000,In_1419);
or U448 (N_448,In_910,In_407);
nand U449 (N_449,In_67,In_1263);
or U450 (N_450,In_1471,In_1910);
nor U451 (N_451,In_1490,In_940);
nand U452 (N_452,In_184,In_1334);
and U453 (N_453,In_1428,In_1091);
nand U454 (N_454,In_606,In_342);
nor U455 (N_455,In_830,In_781);
and U456 (N_456,In_36,In_695);
and U457 (N_457,In_528,In_1392);
or U458 (N_458,In_383,In_374);
nor U459 (N_459,In_554,In_216);
and U460 (N_460,In_1736,In_1254);
or U461 (N_461,In_1881,In_752);
xnor U462 (N_462,In_1731,In_1605);
nor U463 (N_463,In_1462,In_1232);
nor U464 (N_464,In_1804,In_296);
or U465 (N_465,In_203,In_1946);
and U466 (N_466,In_1139,In_1584);
xor U467 (N_467,In_1267,In_1957);
and U468 (N_468,In_1749,In_627);
or U469 (N_469,In_1113,In_795);
and U470 (N_470,In_1710,In_1746);
nand U471 (N_471,In_47,In_525);
nor U472 (N_472,In_50,In_498);
xor U473 (N_473,In_1440,In_1541);
nand U474 (N_474,In_1458,In_1686);
or U475 (N_475,In_1540,In_1970);
nor U476 (N_476,In_1501,In_1459);
or U477 (N_477,In_210,In_7);
xnor U478 (N_478,In_1841,In_273);
or U479 (N_479,In_1067,In_488);
and U480 (N_480,In_1093,In_1737);
nor U481 (N_481,In_428,In_1876);
nand U482 (N_482,In_734,In_1954);
xor U483 (N_483,In_1088,In_1852);
and U484 (N_484,In_1318,In_1588);
xor U485 (N_485,In_1308,In_1291);
xnor U486 (N_486,In_456,In_459);
xor U487 (N_487,In_1569,In_152);
nor U488 (N_488,In_1181,In_717);
and U489 (N_489,In_909,In_1738);
xnor U490 (N_490,In_1228,In_1346);
nor U491 (N_491,In_1636,In_656);
nand U492 (N_492,In_972,In_872);
or U493 (N_493,In_242,In_1047);
nor U494 (N_494,In_1586,In_1520);
nor U495 (N_495,In_295,In_977);
or U496 (N_496,In_1614,In_749);
nor U497 (N_497,In_1355,In_1596);
nand U498 (N_498,In_1550,In_1460);
nor U499 (N_499,In_1249,In_285);
or U500 (N_500,In_1484,In_1869);
and U501 (N_501,In_1527,In_1718);
nor U502 (N_502,In_294,In_1322);
nand U503 (N_503,In_1818,In_1496);
nor U504 (N_504,In_1439,In_1926);
and U505 (N_505,In_1779,In_438);
or U506 (N_506,In_1827,In_1348);
and U507 (N_507,In_63,In_1701);
or U508 (N_508,In_870,In_589);
xnor U509 (N_509,In_850,In_639);
xnor U510 (N_510,In_846,In_402);
nand U511 (N_511,In_1145,In_1832);
nor U512 (N_512,In_1526,In_1681);
or U513 (N_513,In_1041,In_641);
and U514 (N_514,In_1078,In_1186);
and U515 (N_515,In_918,In_380);
nand U516 (N_516,In_301,In_1734);
or U517 (N_517,In_1894,In_801);
and U518 (N_518,In_389,In_245);
nor U519 (N_519,In_1329,In_1573);
nor U520 (N_520,In_932,In_1758);
nor U521 (N_521,In_621,In_898);
nand U522 (N_522,In_968,In_1889);
nor U523 (N_523,In_258,In_1478);
and U524 (N_524,In_1942,In_1492);
nand U525 (N_525,In_366,In_1102);
and U526 (N_526,In_20,In_1173);
or U527 (N_527,In_762,In_324);
nor U528 (N_528,In_1538,In_349);
xnor U529 (N_529,In_707,In_619);
or U530 (N_530,In_139,In_1216);
and U531 (N_531,In_785,In_1642);
nand U532 (N_532,In_1594,In_1893);
nand U533 (N_533,In_608,In_1284);
or U534 (N_534,In_1981,In_485);
xor U535 (N_535,In_90,In_1748);
and U536 (N_536,In_569,In_1656);
nand U537 (N_537,In_1789,In_466);
nand U538 (N_538,In_58,In_1959);
nor U539 (N_539,In_797,In_642);
and U540 (N_540,In_72,In_1515);
nor U541 (N_541,In_1320,In_191);
nor U542 (N_542,In_1206,In_155);
or U543 (N_543,In_204,In_1836);
or U544 (N_544,In_1883,In_1871);
nand U545 (N_545,In_760,In_171);
xor U546 (N_546,In_818,In_399);
nor U547 (N_547,In_1073,In_1345);
xnor U548 (N_548,In_1457,In_1450);
or U549 (N_549,In_647,In_94);
nand U550 (N_550,In_201,In_1132);
nand U551 (N_551,In_1135,In_1752);
nand U552 (N_552,In_640,In_44);
xnor U553 (N_553,In_1220,In_772);
and U554 (N_554,In_558,In_1116);
or U555 (N_555,In_1151,In_1618);
or U556 (N_556,In_555,In_1658);
nand U557 (N_557,In_1682,In_469);
or U558 (N_558,In_565,In_239);
xnor U559 (N_559,In_62,In_878);
and U560 (N_560,In_632,In_1803);
or U561 (N_561,In_1580,In_1733);
xor U562 (N_562,In_928,In_137);
nor U563 (N_563,In_1646,In_56);
or U564 (N_564,In_1123,In_958);
and U565 (N_565,In_25,In_714);
nor U566 (N_566,In_567,In_256);
or U567 (N_567,In_43,In_1678);
xnor U568 (N_568,In_379,In_620);
nand U569 (N_569,In_1469,In_98);
nand U570 (N_570,In_1561,In_798);
nor U571 (N_571,In_1395,In_1309);
nand U572 (N_572,In_1918,In_1989);
nand U573 (N_573,In_959,In_37);
or U574 (N_574,In_1544,In_142);
nand U575 (N_575,In_247,In_1146);
nor U576 (N_576,In_1311,In_250);
nand U577 (N_577,In_336,In_1545);
nor U578 (N_578,In_1054,In_1014);
or U579 (N_579,In_362,In_1691);
and U580 (N_580,In_889,In_505);
nand U581 (N_581,In_804,In_877);
and U582 (N_582,In_235,In_1397);
and U583 (N_583,In_306,In_1729);
and U584 (N_584,In_857,In_28);
or U585 (N_585,In_1,In_470);
nor U586 (N_586,In_1426,In_1307);
or U587 (N_587,In_624,In_809);
or U588 (N_588,In_1391,In_1829);
or U589 (N_589,In_1367,In_369);
nor U590 (N_590,In_275,In_930);
nand U591 (N_591,In_1556,In_309);
or U592 (N_592,In_1530,In_1120);
nor U593 (N_593,In_976,In_1369);
and U594 (N_594,In_776,In_1268);
or U595 (N_595,In_1885,In_68);
nor U596 (N_596,In_560,In_317);
or U597 (N_597,In_726,In_1630);
nand U598 (N_598,In_1523,In_1386);
and U599 (N_599,In_941,In_547);
and U600 (N_600,In_916,In_1105);
nor U601 (N_601,In_1071,In_507);
nor U602 (N_602,In_1383,In_348);
and U603 (N_603,In_1566,In_1495);
xor U604 (N_604,In_1195,In_230);
nor U605 (N_605,In_755,In_460);
or U606 (N_606,In_475,In_542);
nor U607 (N_607,In_512,In_221);
nor U608 (N_608,In_724,In_858);
and U609 (N_609,In_1848,In_316);
and U610 (N_610,In_166,In_1794);
nand U611 (N_611,In_662,In_1744);
or U612 (N_612,In_5,In_1906);
nand U613 (N_613,In_433,In_129);
nor U614 (N_614,In_1685,In_1536);
nor U615 (N_615,In_1854,In_1129);
or U616 (N_616,In_729,In_480);
or U617 (N_617,In_39,In_688);
and U618 (N_618,In_106,In_1379);
and U619 (N_619,In_392,In_1094);
nand U620 (N_620,In_1184,In_716);
or U621 (N_621,In_1861,In_6);
or U622 (N_622,In_1410,In_1235);
and U623 (N_623,In_1645,In_422);
nand U624 (N_624,In_1432,In_936);
or U625 (N_625,In_859,In_1785);
nand U626 (N_626,In_354,In_231);
nor U627 (N_627,In_1937,In_1062);
or U628 (N_628,In_987,In_1726);
nand U629 (N_629,In_915,In_409);
or U630 (N_630,In_1866,In_1874);
and U631 (N_631,In_969,In_1781);
nand U632 (N_632,In_1310,In_630);
nand U633 (N_633,In_1565,In_1051);
or U634 (N_634,In_281,In_851);
nor U635 (N_635,In_1896,In_1038);
xor U636 (N_636,In_828,In_652);
nand U637 (N_637,In_725,In_1079);
and U638 (N_638,In_223,In_87);
and U639 (N_639,In_1868,In_645);
and U640 (N_640,In_405,In_1161);
and U641 (N_641,In_1092,In_83);
or U642 (N_642,In_1938,In_411);
or U643 (N_643,In_1303,In_1015);
xor U644 (N_644,In_1960,In_1870);
nor U645 (N_645,In_708,In_1714);
and U646 (N_646,In_1289,In_382);
nand U647 (N_647,In_658,In_1407);
nand U648 (N_648,In_1251,In_1751);
nand U649 (N_649,In_1830,In_1995);
or U650 (N_650,In_1175,In_1075);
or U651 (N_651,In_793,In_302);
nor U652 (N_652,In_1517,In_978);
and U653 (N_653,In_337,In_1404);
and U654 (N_654,In_1326,In_575);
or U655 (N_655,In_381,In_289);
and U656 (N_656,In_838,In_350);
or U657 (N_657,In_529,In_1331);
nor U658 (N_658,In_1817,In_1514);
xnor U659 (N_659,In_502,In_866);
and U660 (N_660,In_657,In_1983);
and U661 (N_661,In_80,In_770);
or U662 (N_662,In_440,In_8);
nand U663 (N_663,In_763,In_553);
and U664 (N_664,In_232,In_1956);
nand U665 (N_665,In_1846,In_682);
nor U666 (N_666,In_1317,In_1613);
nand U667 (N_667,In_1684,In_1672);
nand U668 (N_668,In_668,In_1589);
and U669 (N_669,In_1665,In_1436);
or U670 (N_670,In_1461,In_548);
and U671 (N_671,In_1925,In_283);
or U672 (N_672,In_690,In_1797);
and U673 (N_673,In_121,In_727);
nand U674 (N_674,In_661,In_290);
nand U675 (N_675,In_947,In_646);
and U676 (N_676,In_1828,In_1528);
nor U677 (N_677,In_1358,In_1823);
nand U678 (N_678,In_1422,In_338);
nor U679 (N_679,In_791,In_370);
or U680 (N_680,In_1198,In_538);
or U681 (N_681,In_1083,In_530);
or U682 (N_682,In_1555,In_1150);
nor U683 (N_683,In_1858,In_1725);
nand U684 (N_684,In_519,In_1036);
nand U685 (N_685,In_906,In_854);
and U686 (N_686,In_110,In_320);
or U687 (N_687,In_1699,In_199);
or U688 (N_688,In_1229,In_218);
or U689 (N_689,In_335,In_1024);
nand U690 (N_690,In_644,In_414);
nor U691 (N_691,In_96,In_816);
or U692 (N_692,In_1424,In_1743);
and U693 (N_693,In_1031,In_1238);
or U694 (N_694,In_1371,In_1201);
nand U695 (N_695,In_882,In_209);
and U696 (N_696,In_12,In_1109);
and U697 (N_697,In_465,In_205);
or U698 (N_698,In_468,In_490);
nor U699 (N_699,In_1130,In_638);
or U700 (N_700,In_396,In_1042);
and U701 (N_701,In_984,In_1912);
nand U702 (N_702,In_1692,In_132);
xor U703 (N_703,In_694,In_1821);
and U704 (N_704,In_1287,In_359);
xor U705 (N_705,In_311,In_1913);
or U706 (N_706,In_911,In_1172);
and U707 (N_707,In_183,In_1770);
or U708 (N_708,In_1242,In_1399);
nand U709 (N_709,In_1892,In_1708);
nor U710 (N_710,In_1069,In_593);
nor U711 (N_711,In_1780,In_1103);
and U712 (N_712,In_1411,In_1224);
or U713 (N_713,In_1844,In_1953);
nand U714 (N_714,In_340,In_1248);
or U715 (N_715,In_180,In_334);
and U716 (N_716,In_322,In_1385);
or U717 (N_717,In_417,In_1363);
nor U718 (N_718,In_1070,In_1788);
and U719 (N_719,In_202,In_1364);
nand U720 (N_720,In_0,In_811);
nor U721 (N_721,In_150,In_886);
nor U722 (N_722,In_421,In_1082);
or U723 (N_723,In_896,In_1272);
nor U724 (N_724,In_808,In_23);
and U725 (N_725,In_1537,In_308);
nand U726 (N_726,In_1641,In_730);
and U727 (N_727,In_985,In_1236);
nand U728 (N_728,In_453,In_994);
nand U729 (N_729,In_1068,In_939);
or U730 (N_730,In_1063,In_782);
and U731 (N_731,In_1923,In_1694);
and U732 (N_732,In_1226,In_213);
or U733 (N_733,In_1208,In_581);
nor U734 (N_734,In_1191,In_64);
nor U735 (N_735,In_1480,In_704);
nand U736 (N_736,In_79,In_145);
nand U737 (N_737,In_880,In_1155);
nor U738 (N_738,In_1547,In_179);
or U739 (N_739,In_1904,In_1712);
nand U740 (N_740,In_1511,In_1477);
nand U741 (N_741,In_784,In_1669);
nand U742 (N_742,In_193,In_207);
and U743 (N_743,In_314,In_1372);
and U744 (N_744,In_534,In_869);
or U745 (N_745,In_840,In_1126);
xnor U746 (N_746,In_603,In_1366);
xnor U747 (N_747,In_1376,In_1632);
and U748 (N_748,In_540,In_764);
or U749 (N_749,In_1661,In_1951);
xor U750 (N_750,In_1539,In_544);
nand U751 (N_751,In_837,In_1257);
or U752 (N_752,In_742,In_884);
nand U753 (N_753,In_105,In_552);
nand U754 (N_754,In_1353,In_706);
xnor U755 (N_755,In_623,In_423);
and U756 (N_756,In_999,In_1305);
and U757 (N_757,In_462,In_1285);
nor U758 (N_758,In_1400,In_1676);
or U759 (N_759,In_248,In_684);
xor U760 (N_760,In_9,In_356);
nor U761 (N_761,In_1389,In_914);
nand U762 (N_762,In_279,In_1873);
or U763 (N_763,In_54,In_176);
and U764 (N_764,In_74,In_879);
nor U765 (N_765,In_1087,In_1349);
or U766 (N_766,In_76,In_21);
nor U767 (N_767,In_1333,In_741);
nand U768 (N_768,In_1194,In_1030);
nor U769 (N_769,In_1824,In_1138);
xnor U770 (N_770,In_1930,In_561);
nand U771 (N_771,In_1688,In_255);
and U772 (N_772,In_1911,In_783);
xor U773 (N_773,In_484,In_1431);
nor U774 (N_774,In_1920,In_1875);
and U775 (N_775,In_1599,In_444);
and U776 (N_776,In_1154,In_1430);
nand U777 (N_777,In_823,In_1441);
nor U778 (N_778,In_1456,In_1958);
or U779 (N_779,In_1169,In_313);
or U780 (N_780,In_219,In_343);
nand U781 (N_781,In_1164,In_1505);
nor U782 (N_782,In_852,In_1027);
nand U783 (N_783,In_1952,In_1581);
nand U784 (N_784,In_328,In_1543);
nand U785 (N_785,In_1969,In_1117);
nand U786 (N_786,In_271,In_1924);
xor U787 (N_787,In_1019,In_957);
nand U788 (N_788,In_1535,In_1833);
or U789 (N_789,In_1518,In_111);
nor U790 (N_790,In_613,In_756);
or U791 (N_791,In_134,In_1557);
nand U792 (N_792,In_686,In_894);
and U793 (N_793,In_333,In_748);
xnor U794 (N_794,In_254,In_881);
or U795 (N_795,In_1077,In_1859);
nand U796 (N_796,In_1499,In_360);
and U797 (N_797,In_839,In_377);
nor U798 (N_798,In_476,In_355);
or U799 (N_799,In_1590,In_49);
nor U800 (N_800,In_691,In_352);
and U801 (N_801,In_1813,In_1061);
nand U802 (N_802,In_1629,In_601);
and U803 (N_803,In_270,In_1233);
and U804 (N_804,In_378,In_1443);
and U805 (N_805,In_663,In_1276);
nand U806 (N_806,In_363,In_1899);
or U807 (N_807,In_1606,In_452);
nor U808 (N_808,In_650,In_625);
and U809 (N_809,In_904,In_35);
nor U810 (N_810,In_344,In_1393);
nand U811 (N_811,In_120,In_836);
and U812 (N_812,In_1667,In_75);
nor U813 (N_813,In_1783,In_1039);
nand U814 (N_814,In_1603,In_1265);
nand U815 (N_815,In_1352,In_1898);
and U816 (N_816,In_960,In_515);
nand U817 (N_817,In_93,In_1174);
and U818 (N_818,In_766,In_146);
and U819 (N_819,In_1816,In_1444);
xor U820 (N_820,In_1534,In_1086);
nand U821 (N_821,In_458,In_1790);
nor U822 (N_822,In_116,In_1497);
xnor U823 (N_823,In_597,In_387);
nand U824 (N_824,In_57,In_1124);
nand U825 (N_825,In_1096,In_835);
and U826 (N_826,In_1730,In_1592);
xor U827 (N_827,In_874,In_1239);
nand U828 (N_828,In_1504,In_1052);
nand U829 (N_829,In_1351,In_149);
and U830 (N_830,In_40,In_1764);
or U831 (N_831,In_122,In_670);
or U832 (N_832,In_1023,In_693);
nor U833 (N_833,In_929,In_845);
or U834 (N_834,In_17,In_1324);
or U835 (N_835,In_1745,In_1571);
or U836 (N_836,In_1971,In_931);
nor U837 (N_837,In_1668,In_863);
xor U838 (N_838,In_493,In_260);
nand U839 (N_839,In_1621,In_1843);
nand U840 (N_840,In_944,In_1835);
and U841 (N_841,In_1711,In_114);
and U842 (N_842,In_1165,In_1842);
nand U843 (N_843,In_1298,In_1693);
xnor U844 (N_844,In_666,In_92);
nand U845 (N_845,In_1259,In_966);
nor U846 (N_846,In_448,In_568);
or U847 (N_847,In_160,In_1203);
or U848 (N_848,In_1834,In_513);
nand U849 (N_849,In_1252,In_32);
and U850 (N_850,In_1579,In_1784);
or U851 (N_851,In_168,In_1166);
xor U852 (N_852,In_1631,In_1825);
or U853 (N_853,In_779,In_1635);
or U854 (N_854,In_952,In_1964);
or U855 (N_855,In_1616,In_893);
xnor U856 (N_856,In_660,In_1978);
and U857 (N_857,In_998,In_1048);
and U858 (N_858,In_410,In_948);
and U859 (N_859,In_927,In_902);
or U860 (N_860,In_692,In_1245);
and U861 (N_861,In_1416,In_1634);
or U862 (N_862,In_1542,In_1412);
or U863 (N_863,In_659,In_1182);
and U864 (N_864,In_720,In_341);
nor U865 (N_865,In_549,In_400);
and U866 (N_866,In_1390,In_1753);
nor U867 (N_867,In_1977,In_1306);
nor U868 (N_868,In_431,In_85);
xnor U869 (N_869,In_1597,In_143);
or U870 (N_870,In_1437,In_1297);
or U871 (N_871,In_718,In_497);
or U872 (N_872,In_1178,In_990);
nand U873 (N_873,In_557,In_404);
and U874 (N_874,In_501,In_461);
and U875 (N_875,In_745,In_135);
nor U876 (N_876,In_1649,In_607);
or U877 (N_877,In_41,In_649);
nor U878 (N_878,In_107,In_1294);
nand U879 (N_879,In_331,In_701);
xnor U880 (N_880,In_1163,In_1966);
nor U881 (N_881,In_236,In_1001);
or U882 (N_882,In_1702,In_237);
nand U883 (N_883,In_401,In_1990);
or U884 (N_884,In_536,In_821);
nor U885 (N_885,In_1506,In_1847);
nand U886 (N_886,In_1793,In_504);
xor U887 (N_887,In_109,In_298);
nand U888 (N_888,In_78,In_1767);
nor U889 (N_889,In_1179,In_1292);
and U890 (N_890,In_1011,In_1357);
xor U891 (N_891,In_457,In_983);
xnor U892 (N_892,In_899,In_942);
nor U893 (N_893,In_1213,In_921);
and U894 (N_894,In_1085,In_1221);
xor U895 (N_895,In_771,In_543);
and U896 (N_896,In_1675,In_1600);
nor U897 (N_897,In_1418,In_907);
nor U898 (N_898,In_1374,In_963);
and U899 (N_899,In_537,In_1772);
nor U900 (N_900,In_1757,In_955);
or U901 (N_901,In_347,In_1968);
nor U902 (N_902,In_413,In_1453);
nor U903 (N_903,In_1760,In_743);
or U904 (N_904,In_1089,In_69);
nor U905 (N_905,In_1447,In_1551);
nor U906 (N_906,In_1190,In_1974);
and U907 (N_907,In_685,In_211);
xor U908 (N_908,In_229,In_1316);
or U909 (N_909,In_991,In_376);
and U910 (N_910,In_653,In_1137);
xnor U911 (N_911,In_1786,In_970);
or U912 (N_912,In_1604,In_559);
or U913 (N_913,In_1864,In_1321);
and U914 (N_914,In_1101,In_744);
or U915 (N_915,In_935,In_570);
nand U916 (N_916,In_710,In_1149);
or U917 (N_917,In_1700,In_933);
nand U918 (N_918,In_1319,In_1187);
or U919 (N_919,In_631,In_687);
or U920 (N_920,In_1045,In_264);
nor U921 (N_921,In_346,In_81);
nand U922 (N_922,In_430,In_1275);
and U923 (N_923,In_588,In_162);
nand U924 (N_924,In_77,In_48);
nand U925 (N_925,In_267,In_1548);
nor U926 (N_926,In_715,In_1976);
nor U927 (N_927,In_1487,In_778);
nor U928 (N_928,In_1973,In_951);
nand U929 (N_929,In_1988,In_1396);
or U930 (N_930,In_1509,In_228);
and U931 (N_931,In_1347,In_1016);
or U932 (N_932,In_364,In_1972);
xor U933 (N_933,In_788,In_1323);
or U934 (N_934,In_1663,In_153);
nand U935 (N_935,In_1222,In_102);
and U936 (N_936,In_842,In_1425);
xnor U937 (N_937,In_1840,In_1218);
xor U938 (N_938,In_108,In_508);
and U939 (N_939,In_1948,In_1759);
xnor U940 (N_940,In_99,In_1563);
or U941 (N_941,In_1809,In_432);
and U942 (N_942,In_956,In_253);
or U943 (N_943,In_1826,In_408);
or U944 (N_944,In_1791,In_573);
or U945 (N_945,In_1941,In_483);
nor U946 (N_946,In_1025,In_848);
nor U947 (N_947,In_616,In_1762);
or U948 (N_948,In_709,In_1193);
and U949 (N_949,In_1053,In_1037);
nand U950 (N_950,In_386,In_1448);
and U951 (N_951,In_1455,In_1979);
nor U952 (N_952,In_1158,In_1531);
nand U953 (N_953,In_1502,In_1350);
or U954 (N_954,In_371,In_365);
nor U955 (N_955,In_1332,In_1157);
xor U956 (N_956,In_148,In_831);
nand U957 (N_957,In_1677,In_1256);
or U958 (N_958,In_1915,In_964);
and U959 (N_959,In_511,In_1377);
or U960 (N_960,In_1266,In_167);
and U961 (N_961,In_803,In_1134);
nand U962 (N_962,In_1095,In_393);
nand U963 (N_963,In_345,In_1148);
or U964 (N_964,In_446,In_699);
and U965 (N_965,In_130,In_1882);
nor U966 (N_966,In_1507,In_1465);
nand U967 (N_967,In_1810,In_1434);
or U968 (N_968,In_1185,In_1340);
nand U969 (N_969,In_451,In_1558);
nand U970 (N_970,In_1716,In_792);
nor U971 (N_971,In_524,In_1330);
and U972 (N_972,In_412,In_1900);
and U973 (N_973,In_1066,In_1849);
nor U974 (N_974,In_220,In_1838);
nand U975 (N_975,In_1601,In_871);
xor U976 (N_976,In_1260,In_416);
or U977 (N_977,In_908,In_1128);
nor U978 (N_978,In_467,In_903);
and U979 (N_979,In_973,In_1795);
nand U980 (N_980,In_634,In_1800);
or U981 (N_981,In_1992,In_1467);
and U982 (N_982,In_1932,In_372);
and U983 (N_983,In_1856,In_847);
or U984 (N_984,In_280,In_91);
and U985 (N_985,In_1339,In_1796);
or U986 (N_986,In_1217,In_1452);
nor U987 (N_987,In_181,In_1769);
nand U988 (N_988,In_61,In_643);
and U989 (N_989,In_198,In_1704);
and U990 (N_990,In_522,In_1513);
or U991 (N_991,In_11,In_777);
or U992 (N_992,In_965,In_1947);
nor U993 (N_993,In_173,In_463);
or U994 (N_994,In_635,In_436);
and U995 (N_995,In_1246,In_1755);
or U996 (N_996,In_599,In_669);
or U997 (N_997,In_629,In_1098);
nand U998 (N_998,In_1044,In_679);
or U999 (N_999,In_533,In_527);
nand U1000 (N_1000,In_1017,In_1506);
and U1001 (N_1001,In_85,In_1569);
or U1002 (N_1002,In_1326,In_913);
nand U1003 (N_1003,In_183,In_1194);
or U1004 (N_1004,In_1108,In_586);
nand U1005 (N_1005,In_400,In_362);
nor U1006 (N_1006,In_579,In_1790);
and U1007 (N_1007,In_1250,In_688);
xor U1008 (N_1008,In_1730,In_44);
and U1009 (N_1009,In_1824,In_1066);
and U1010 (N_1010,In_590,In_1888);
and U1011 (N_1011,In_346,In_902);
nand U1012 (N_1012,In_1486,In_190);
and U1013 (N_1013,In_1891,In_1728);
nand U1014 (N_1014,In_1202,In_1442);
or U1015 (N_1015,In_867,In_163);
nand U1016 (N_1016,In_1258,In_1276);
nand U1017 (N_1017,In_384,In_1817);
nand U1018 (N_1018,In_1807,In_1325);
and U1019 (N_1019,In_929,In_1708);
and U1020 (N_1020,In_1386,In_1444);
xnor U1021 (N_1021,In_1507,In_1142);
nand U1022 (N_1022,In_54,In_517);
and U1023 (N_1023,In_856,In_1283);
or U1024 (N_1024,In_1260,In_524);
or U1025 (N_1025,In_1132,In_113);
nand U1026 (N_1026,In_55,In_1522);
or U1027 (N_1027,In_658,In_589);
and U1028 (N_1028,In_685,In_1023);
or U1029 (N_1029,In_1482,In_580);
and U1030 (N_1030,In_563,In_189);
nor U1031 (N_1031,In_995,In_740);
or U1032 (N_1032,In_430,In_1046);
and U1033 (N_1033,In_844,In_7);
xnor U1034 (N_1034,In_1978,In_511);
or U1035 (N_1035,In_1088,In_1185);
and U1036 (N_1036,In_241,In_554);
xor U1037 (N_1037,In_175,In_822);
xor U1038 (N_1038,In_138,In_105);
xor U1039 (N_1039,In_1014,In_14);
nor U1040 (N_1040,In_123,In_1402);
nand U1041 (N_1041,In_1208,In_598);
and U1042 (N_1042,In_40,In_52);
or U1043 (N_1043,In_1704,In_1985);
nand U1044 (N_1044,In_1018,In_1085);
nand U1045 (N_1045,In_734,In_1670);
nand U1046 (N_1046,In_1901,In_1666);
or U1047 (N_1047,In_166,In_1266);
xor U1048 (N_1048,In_1915,In_806);
nor U1049 (N_1049,In_1108,In_114);
xor U1050 (N_1050,In_1985,In_1628);
nor U1051 (N_1051,In_642,In_959);
and U1052 (N_1052,In_1131,In_1885);
nor U1053 (N_1053,In_691,In_1381);
nor U1054 (N_1054,In_429,In_1758);
nand U1055 (N_1055,In_228,In_487);
nand U1056 (N_1056,In_291,In_420);
and U1057 (N_1057,In_1841,In_1952);
nor U1058 (N_1058,In_1088,In_573);
or U1059 (N_1059,In_15,In_1141);
or U1060 (N_1060,In_1956,In_85);
and U1061 (N_1061,In_1229,In_691);
or U1062 (N_1062,In_258,In_1674);
nand U1063 (N_1063,In_875,In_927);
xnor U1064 (N_1064,In_297,In_1041);
nor U1065 (N_1065,In_1578,In_1043);
or U1066 (N_1066,In_854,In_1591);
and U1067 (N_1067,In_1539,In_328);
or U1068 (N_1068,In_758,In_1238);
or U1069 (N_1069,In_1755,In_882);
or U1070 (N_1070,In_423,In_325);
or U1071 (N_1071,In_841,In_1458);
nor U1072 (N_1072,In_644,In_1650);
and U1073 (N_1073,In_443,In_672);
xor U1074 (N_1074,In_555,In_753);
and U1075 (N_1075,In_409,In_1020);
nor U1076 (N_1076,In_652,In_1879);
and U1077 (N_1077,In_1112,In_599);
nand U1078 (N_1078,In_252,In_1);
nor U1079 (N_1079,In_1938,In_104);
nand U1080 (N_1080,In_1573,In_1271);
or U1081 (N_1081,In_29,In_297);
nor U1082 (N_1082,In_924,In_1212);
xnor U1083 (N_1083,In_1152,In_493);
xnor U1084 (N_1084,In_822,In_1947);
or U1085 (N_1085,In_1115,In_770);
or U1086 (N_1086,In_78,In_1717);
and U1087 (N_1087,In_842,In_999);
nor U1088 (N_1088,In_1718,In_1536);
and U1089 (N_1089,In_1598,In_1473);
or U1090 (N_1090,In_1565,In_1001);
xor U1091 (N_1091,In_522,In_52);
or U1092 (N_1092,In_1064,In_1419);
or U1093 (N_1093,In_1298,In_1595);
nor U1094 (N_1094,In_1801,In_233);
xnor U1095 (N_1095,In_488,In_1965);
nand U1096 (N_1096,In_1196,In_1446);
and U1097 (N_1097,In_1180,In_1669);
nor U1098 (N_1098,In_581,In_540);
or U1099 (N_1099,In_1640,In_408);
and U1100 (N_1100,In_371,In_276);
xor U1101 (N_1101,In_300,In_1345);
or U1102 (N_1102,In_298,In_1309);
or U1103 (N_1103,In_63,In_331);
nor U1104 (N_1104,In_1635,In_142);
and U1105 (N_1105,In_570,In_1921);
and U1106 (N_1106,In_945,In_1416);
or U1107 (N_1107,In_108,In_649);
nor U1108 (N_1108,In_1404,In_1944);
nand U1109 (N_1109,In_895,In_1387);
xnor U1110 (N_1110,In_367,In_1961);
or U1111 (N_1111,In_167,In_1828);
nand U1112 (N_1112,In_87,In_982);
and U1113 (N_1113,In_1295,In_122);
and U1114 (N_1114,In_1533,In_1440);
xnor U1115 (N_1115,In_914,In_1343);
xor U1116 (N_1116,In_746,In_287);
and U1117 (N_1117,In_1485,In_1601);
xor U1118 (N_1118,In_955,In_461);
xor U1119 (N_1119,In_1320,In_1983);
nor U1120 (N_1120,In_1185,In_1958);
nor U1121 (N_1121,In_1678,In_1787);
or U1122 (N_1122,In_1740,In_684);
nor U1123 (N_1123,In_1732,In_650);
nand U1124 (N_1124,In_779,In_505);
xnor U1125 (N_1125,In_677,In_627);
and U1126 (N_1126,In_125,In_560);
nand U1127 (N_1127,In_541,In_1979);
and U1128 (N_1128,In_1283,In_1445);
and U1129 (N_1129,In_1773,In_496);
and U1130 (N_1130,In_662,In_1141);
and U1131 (N_1131,In_501,In_1820);
and U1132 (N_1132,In_1894,In_1790);
or U1133 (N_1133,In_1930,In_188);
nand U1134 (N_1134,In_1451,In_70);
nor U1135 (N_1135,In_384,In_1210);
xnor U1136 (N_1136,In_1103,In_121);
nor U1137 (N_1137,In_461,In_1957);
xor U1138 (N_1138,In_131,In_1308);
nor U1139 (N_1139,In_1224,In_131);
nor U1140 (N_1140,In_351,In_1755);
nor U1141 (N_1141,In_114,In_1253);
or U1142 (N_1142,In_374,In_877);
and U1143 (N_1143,In_326,In_1472);
or U1144 (N_1144,In_1576,In_901);
nor U1145 (N_1145,In_973,In_453);
nand U1146 (N_1146,In_216,In_1225);
or U1147 (N_1147,In_1685,In_97);
nand U1148 (N_1148,In_693,In_129);
nand U1149 (N_1149,In_1820,In_752);
nand U1150 (N_1150,In_1465,In_344);
xnor U1151 (N_1151,In_329,In_209);
or U1152 (N_1152,In_1637,In_650);
nor U1153 (N_1153,In_1021,In_222);
nand U1154 (N_1154,In_511,In_444);
nand U1155 (N_1155,In_939,In_1837);
and U1156 (N_1156,In_276,In_1496);
nor U1157 (N_1157,In_1945,In_1057);
xor U1158 (N_1158,In_1559,In_1022);
or U1159 (N_1159,In_439,In_485);
xnor U1160 (N_1160,In_343,In_750);
nor U1161 (N_1161,In_99,In_937);
or U1162 (N_1162,In_1491,In_1269);
nand U1163 (N_1163,In_1035,In_796);
nor U1164 (N_1164,In_394,In_777);
nand U1165 (N_1165,In_1334,In_1396);
nand U1166 (N_1166,In_997,In_1114);
or U1167 (N_1167,In_770,In_902);
and U1168 (N_1168,In_1321,In_125);
or U1169 (N_1169,In_293,In_169);
or U1170 (N_1170,In_1330,In_1221);
nand U1171 (N_1171,In_1903,In_404);
and U1172 (N_1172,In_1635,In_227);
nor U1173 (N_1173,In_464,In_1);
nor U1174 (N_1174,In_200,In_1282);
nand U1175 (N_1175,In_1058,In_1173);
xor U1176 (N_1176,In_1484,In_1468);
and U1177 (N_1177,In_1590,In_1699);
and U1178 (N_1178,In_1277,In_1249);
or U1179 (N_1179,In_1474,In_1546);
nor U1180 (N_1180,In_1283,In_380);
nand U1181 (N_1181,In_1970,In_488);
and U1182 (N_1182,In_1920,In_1915);
nand U1183 (N_1183,In_133,In_1035);
and U1184 (N_1184,In_1658,In_1018);
nand U1185 (N_1185,In_642,In_1921);
xor U1186 (N_1186,In_1885,In_1111);
nor U1187 (N_1187,In_1609,In_1210);
or U1188 (N_1188,In_1967,In_1028);
or U1189 (N_1189,In_726,In_855);
and U1190 (N_1190,In_1259,In_778);
nor U1191 (N_1191,In_1202,In_844);
xor U1192 (N_1192,In_1814,In_1966);
xor U1193 (N_1193,In_1117,In_1036);
and U1194 (N_1194,In_1975,In_274);
and U1195 (N_1195,In_1822,In_1876);
or U1196 (N_1196,In_347,In_1815);
or U1197 (N_1197,In_124,In_951);
and U1198 (N_1198,In_1919,In_1556);
nand U1199 (N_1199,In_1200,In_1239);
nand U1200 (N_1200,In_1552,In_984);
nor U1201 (N_1201,In_150,In_508);
xnor U1202 (N_1202,In_770,In_1908);
nor U1203 (N_1203,In_343,In_855);
and U1204 (N_1204,In_1081,In_321);
nor U1205 (N_1205,In_1672,In_1188);
or U1206 (N_1206,In_1004,In_1759);
nor U1207 (N_1207,In_1747,In_1613);
nand U1208 (N_1208,In_177,In_765);
nor U1209 (N_1209,In_513,In_141);
nand U1210 (N_1210,In_1309,In_1377);
or U1211 (N_1211,In_121,In_1815);
nor U1212 (N_1212,In_1170,In_1569);
xnor U1213 (N_1213,In_219,In_687);
nand U1214 (N_1214,In_1303,In_247);
nand U1215 (N_1215,In_1856,In_1023);
or U1216 (N_1216,In_1707,In_76);
xor U1217 (N_1217,In_160,In_791);
nor U1218 (N_1218,In_1823,In_156);
or U1219 (N_1219,In_524,In_1623);
and U1220 (N_1220,In_1997,In_1715);
and U1221 (N_1221,In_171,In_27);
and U1222 (N_1222,In_887,In_1735);
nor U1223 (N_1223,In_1823,In_1718);
nand U1224 (N_1224,In_119,In_1389);
or U1225 (N_1225,In_1119,In_1800);
or U1226 (N_1226,In_1986,In_541);
and U1227 (N_1227,In_506,In_1781);
nand U1228 (N_1228,In_1559,In_593);
or U1229 (N_1229,In_328,In_144);
and U1230 (N_1230,In_364,In_1407);
nand U1231 (N_1231,In_1169,In_105);
and U1232 (N_1232,In_225,In_1734);
nor U1233 (N_1233,In_1627,In_598);
nand U1234 (N_1234,In_440,In_1330);
xor U1235 (N_1235,In_196,In_86);
nor U1236 (N_1236,In_1556,In_650);
nor U1237 (N_1237,In_1105,In_1929);
or U1238 (N_1238,In_226,In_196);
or U1239 (N_1239,In_1773,In_1050);
or U1240 (N_1240,In_114,In_236);
xnor U1241 (N_1241,In_526,In_1060);
nand U1242 (N_1242,In_1528,In_922);
or U1243 (N_1243,In_857,In_216);
nor U1244 (N_1244,In_1013,In_45);
and U1245 (N_1245,In_1618,In_705);
nor U1246 (N_1246,In_1826,In_1189);
and U1247 (N_1247,In_781,In_1867);
nor U1248 (N_1248,In_1192,In_1564);
xor U1249 (N_1249,In_542,In_1046);
and U1250 (N_1250,In_1991,In_1333);
or U1251 (N_1251,In_1750,In_982);
or U1252 (N_1252,In_1102,In_253);
nor U1253 (N_1253,In_1339,In_1941);
nand U1254 (N_1254,In_105,In_728);
or U1255 (N_1255,In_1178,In_1287);
nor U1256 (N_1256,In_1072,In_172);
nor U1257 (N_1257,In_161,In_1152);
nand U1258 (N_1258,In_1084,In_333);
and U1259 (N_1259,In_1246,In_1287);
nand U1260 (N_1260,In_115,In_904);
or U1261 (N_1261,In_768,In_1642);
or U1262 (N_1262,In_1598,In_694);
and U1263 (N_1263,In_383,In_674);
nand U1264 (N_1264,In_1552,In_770);
or U1265 (N_1265,In_54,In_1584);
nor U1266 (N_1266,In_1911,In_1695);
nor U1267 (N_1267,In_1127,In_390);
nand U1268 (N_1268,In_979,In_1958);
or U1269 (N_1269,In_1786,In_307);
or U1270 (N_1270,In_229,In_864);
or U1271 (N_1271,In_1491,In_1006);
nor U1272 (N_1272,In_1199,In_1584);
and U1273 (N_1273,In_1310,In_1728);
nor U1274 (N_1274,In_471,In_664);
nand U1275 (N_1275,In_1832,In_1304);
and U1276 (N_1276,In_255,In_1065);
nor U1277 (N_1277,In_560,In_574);
nand U1278 (N_1278,In_577,In_311);
nor U1279 (N_1279,In_835,In_1406);
or U1280 (N_1280,In_893,In_968);
and U1281 (N_1281,In_1862,In_100);
or U1282 (N_1282,In_8,In_69);
nand U1283 (N_1283,In_14,In_742);
or U1284 (N_1284,In_1766,In_1269);
nor U1285 (N_1285,In_687,In_1525);
and U1286 (N_1286,In_170,In_343);
or U1287 (N_1287,In_1756,In_76);
and U1288 (N_1288,In_1960,In_776);
nand U1289 (N_1289,In_1008,In_1928);
nor U1290 (N_1290,In_1278,In_764);
and U1291 (N_1291,In_739,In_1139);
and U1292 (N_1292,In_1083,In_1192);
or U1293 (N_1293,In_1336,In_1128);
nand U1294 (N_1294,In_795,In_891);
nand U1295 (N_1295,In_546,In_209);
nand U1296 (N_1296,In_654,In_1893);
nand U1297 (N_1297,In_477,In_1475);
nand U1298 (N_1298,In_1067,In_536);
nand U1299 (N_1299,In_1186,In_1419);
and U1300 (N_1300,In_933,In_1630);
and U1301 (N_1301,In_1043,In_4);
and U1302 (N_1302,In_22,In_1870);
nor U1303 (N_1303,In_366,In_442);
nor U1304 (N_1304,In_1393,In_1789);
and U1305 (N_1305,In_1423,In_415);
nor U1306 (N_1306,In_463,In_1024);
and U1307 (N_1307,In_1977,In_663);
nor U1308 (N_1308,In_1989,In_1367);
and U1309 (N_1309,In_1508,In_399);
or U1310 (N_1310,In_195,In_1977);
and U1311 (N_1311,In_1504,In_1299);
nor U1312 (N_1312,In_1592,In_1450);
and U1313 (N_1313,In_1948,In_1896);
nor U1314 (N_1314,In_280,In_1417);
and U1315 (N_1315,In_1357,In_351);
nand U1316 (N_1316,In_924,In_829);
nor U1317 (N_1317,In_1678,In_1395);
and U1318 (N_1318,In_749,In_1751);
nand U1319 (N_1319,In_1296,In_406);
nand U1320 (N_1320,In_1610,In_841);
nand U1321 (N_1321,In_1989,In_1654);
nor U1322 (N_1322,In_388,In_51);
nor U1323 (N_1323,In_260,In_515);
nor U1324 (N_1324,In_984,In_366);
xor U1325 (N_1325,In_1334,In_1249);
nor U1326 (N_1326,In_490,In_785);
nor U1327 (N_1327,In_1877,In_1654);
nand U1328 (N_1328,In_1833,In_507);
nand U1329 (N_1329,In_1894,In_223);
or U1330 (N_1330,In_14,In_168);
nor U1331 (N_1331,In_835,In_380);
nor U1332 (N_1332,In_981,In_1668);
nor U1333 (N_1333,In_1211,In_915);
or U1334 (N_1334,In_252,In_883);
xor U1335 (N_1335,In_378,In_958);
or U1336 (N_1336,In_290,In_946);
nand U1337 (N_1337,In_1186,In_1659);
or U1338 (N_1338,In_1386,In_775);
and U1339 (N_1339,In_363,In_1351);
or U1340 (N_1340,In_698,In_1062);
and U1341 (N_1341,In_1961,In_1955);
xor U1342 (N_1342,In_1003,In_794);
nor U1343 (N_1343,In_1011,In_1087);
xnor U1344 (N_1344,In_1055,In_995);
nor U1345 (N_1345,In_1249,In_1394);
nand U1346 (N_1346,In_1633,In_1092);
and U1347 (N_1347,In_1940,In_1839);
or U1348 (N_1348,In_1770,In_235);
and U1349 (N_1349,In_1672,In_724);
nor U1350 (N_1350,In_844,In_378);
and U1351 (N_1351,In_1673,In_120);
nor U1352 (N_1352,In_50,In_421);
nor U1353 (N_1353,In_1563,In_516);
nand U1354 (N_1354,In_752,In_597);
or U1355 (N_1355,In_576,In_153);
nand U1356 (N_1356,In_962,In_1478);
nand U1357 (N_1357,In_244,In_619);
nand U1358 (N_1358,In_1768,In_957);
xor U1359 (N_1359,In_1746,In_932);
xnor U1360 (N_1360,In_1988,In_764);
xnor U1361 (N_1361,In_527,In_431);
and U1362 (N_1362,In_1030,In_521);
nor U1363 (N_1363,In_635,In_1684);
nand U1364 (N_1364,In_1135,In_833);
nand U1365 (N_1365,In_544,In_603);
nand U1366 (N_1366,In_1005,In_1711);
nand U1367 (N_1367,In_1819,In_1569);
and U1368 (N_1368,In_1875,In_1733);
or U1369 (N_1369,In_1767,In_976);
nor U1370 (N_1370,In_882,In_462);
and U1371 (N_1371,In_1264,In_1353);
nor U1372 (N_1372,In_17,In_717);
or U1373 (N_1373,In_1502,In_58);
and U1374 (N_1374,In_282,In_88);
nand U1375 (N_1375,In_538,In_1086);
and U1376 (N_1376,In_1940,In_1393);
and U1377 (N_1377,In_467,In_630);
nand U1378 (N_1378,In_1131,In_1374);
or U1379 (N_1379,In_1628,In_998);
xnor U1380 (N_1380,In_16,In_1301);
or U1381 (N_1381,In_505,In_1510);
and U1382 (N_1382,In_1965,In_902);
and U1383 (N_1383,In_398,In_873);
nand U1384 (N_1384,In_1616,In_1414);
and U1385 (N_1385,In_405,In_345);
nand U1386 (N_1386,In_1421,In_1117);
and U1387 (N_1387,In_1112,In_718);
nand U1388 (N_1388,In_1969,In_843);
nand U1389 (N_1389,In_782,In_892);
or U1390 (N_1390,In_1750,In_756);
or U1391 (N_1391,In_1284,In_1037);
or U1392 (N_1392,In_1767,In_1861);
nor U1393 (N_1393,In_1019,In_724);
nand U1394 (N_1394,In_1392,In_1592);
nand U1395 (N_1395,In_946,In_1225);
or U1396 (N_1396,In_690,In_1620);
or U1397 (N_1397,In_1493,In_974);
nand U1398 (N_1398,In_446,In_1918);
or U1399 (N_1399,In_146,In_1295);
nand U1400 (N_1400,In_128,In_550);
nor U1401 (N_1401,In_322,In_785);
or U1402 (N_1402,In_1370,In_426);
nor U1403 (N_1403,In_506,In_405);
nand U1404 (N_1404,In_1024,In_1786);
xnor U1405 (N_1405,In_1775,In_1270);
and U1406 (N_1406,In_693,In_1887);
and U1407 (N_1407,In_403,In_509);
nand U1408 (N_1408,In_32,In_1610);
or U1409 (N_1409,In_640,In_544);
or U1410 (N_1410,In_906,In_1440);
and U1411 (N_1411,In_1622,In_647);
xnor U1412 (N_1412,In_707,In_686);
or U1413 (N_1413,In_1239,In_1064);
nand U1414 (N_1414,In_1934,In_1546);
nor U1415 (N_1415,In_190,In_1122);
or U1416 (N_1416,In_1235,In_222);
or U1417 (N_1417,In_225,In_843);
or U1418 (N_1418,In_1755,In_1237);
nand U1419 (N_1419,In_656,In_561);
nor U1420 (N_1420,In_1289,In_1408);
nor U1421 (N_1421,In_1811,In_396);
and U1422 (N_1422,In_1265,In_1437);
nand U1423 (N_1423,In_1056,In_980);
or U1424 (N_1424,In_1698,In_239);
and U1425 (N_1425,In_310,In_528);
or U1426 (N_1426,In_465,In_717);
nand U1427 (N_1427,In_986,In_339);
or U1428 (N_1428,In_654,In_1431);
nand U1429 (N_1429,In_787,In_1297);
and U1430 (N_1430,In_929,In_1852);
nand U1431 (N_1431,In_1459,In_134);
or U1432 (N_1432,In_1011,In_1660);
and U1433 (N_1433,In_1041,In_1135);
nand U1434 (N_1434,In_316,In_379);
nand U1435 (N_1435,In_898,In_1060);
and U1436 (N_1436,In_1529,In_1753);
and U1437 (N_1437,In_226,In_1890);
nand U1438 (N_1438,In_1016,In_1564);
nand U1439 (N_1439,In_1292,In_651);
or U1440 (N_1440,In_1107,In_352);
or U1441 (N_1441,In_49,In_623);
nor U1442 (N_1442,In_1833,In_342);
nand U1443 (N_1443,In_1163,In_1694);
or U1444 (N_1444,In_1898,In_109);
xnor U1445 (N_1445,In_1654,In_680);
and U1446 (N_1446,In_931,In_193);
or U1447 (N_1447,In_1481,In_33);
nand U1448 (N_1448,In_296,In_1139);
nand U1449 (N_1449,In_617,In_1540);
nand U1450 (N_1450,In_1820,In_1457);
and U1451 (N_1451,In_450,In_600);
and U1452 (N_1452,In_520,In_1247);
nand U1453 (N_1453,In_1213,In_706);
nand U1454 (N_1454,In_1076,In_1503);
nand U1455 (N_1455,In_1493,In_309);
nand U1456 (N_1456,In_979,In_422);
or U1457 (N_1457,In_1664,In_415);
or U1458 (N_1458,In_1952,In_1586);
or U1459 (N_1459,In_254,In_1322);
xor U1460 (N_1460,In_1645,In_716);
nor U1461 (N_1461,In_1464,In_820);
nor U1462 (N_1462,In_1998,In_1638);
nor U1463 (N_1463,In_1776,In_884);
or U1464 (N_1464,In_960,In_25);
and U1465 (N_1465,In_1336,In_770);
xnor U1466 (N_1466,In_1698,In_1216);
nand U1467 (N_1467,In_804,In_151);
nor U1468 (N_1468,In_535,In_866);
nor U1469 (N_1469,In_981,In_365);
and U1470 (N_1470,In_944,In_531);
nand U1471 (N_1471,In_704,In_1615);
nor U1472 (N_1472,In_477,In_545);
or U1473 (N_1473,In_618,In_765);
nand U1474 (N_1474,In_1339,In_458);
xnor U1475 (N_1475,In_398,In_1199);
or U1476 (N_1476,In_1286,In_919);
xnor U1477 (N_1477,In_85,In_877);
and U1478 (N_1478,In_98,In_420);
nand U1479 (N_1479,In_1974,In_792);
or U1480 (N_1480,In_1147,In_1322);
xnor U1481 (N_1481,In_958,In_367);
and U1482 (N_1482,In_1296,In_84);
xor U1483 (N_1483,In_1155,In_152);
nor U1484 (N_1484,In_513,In_21);
and U1485 (N_1485,In_1559,In_1152);
nand U1486 (N_1486,In_1400,In_1688);
and U1487 (N_1487,In_1926,In_299);
and U1488 (N_1488,In_1796,In_1730);
or U1489 (N_1489,In_1695,In_975);
nor U1490 (N_1490,In_1754,In_406);
nor U1491 (N_1491,In_818,In_550);
or U1492 (N_1492,In_599,In_1972);
and U1493 (N_1493,In_557,In_670);
nand U1494 (N_1494,In_60,In_1584);
and U1495 (N_1495,In_1461,In_902);
or U1496 (N_1496,In_27,In_681);
or U1497 (N_1497,In_1225,In_1319);
nand U1498 (N_1498,In_615,In_202);
nor U1499 (N_1499,In_820,In_91);
or U1500 (N_1500,In_1859,In_1436);
nor U1501 (N_1501,In_381,In_26);
nor U1502 (N_1502,In_1204,In_437);
xnor U1503 (N_1503,In_456,In_1736);
nor U1504 (N_1504,In_1811,In_579);
or U1505 (N_1505,In_501,In_59);
and U1506 (N_1506,In_186,In_1448);
xor U1507 (N_1507,In_869,In_422);
or U1508 (N_1508,In_955,In_559);
or U1509 (N_1509,In_1288,In_1046);
or U1510 (N_1510,In_1686,In_214);
and U1511 (N_1511,In_104,In_27);
or U1512 (N_1512,In_197,In_1905);
nor U1513 (N_1513,In_1109,In_130);
or U1514 (N_1514,In_1278,In_1951);
and U1515 (N_1515,In_212,In_1347);
nand U1516 (N_1516,In_105,In_78);
or U1517 (N_1517,In_1138,In_204);
and U1518 (N_1518,In_1293,In_647);
or U1519 (N_1519,In_1959,In_1853);
xnor U1520 (N_1520,In_606,In_1188);
nand U1521 (N_1521,In_1147,In_1932);
nand U1522 (N_1522,In_1679,In_439);
or U1523 (N_1523,In_1374,In_55);
or U1524 (N_1524,In_1089,In_1621);
nor U1525 (N_1525,In_484,In_1750);
and U1526 (N_1526,In_1619,In_1804);
nand U1527 (N_1527,In_1758,In_536);
and U1528 (N_1528,In_638,In_1237);
and U1529 (N_1529,In_219,In_1839);
nor U1530 (N_1530,In_1154,In_326);
or U1531 (N_1531,In_750,In_844);
or U1532 (N_1532,In_1861,In_1392);
and U1533 (N_1533,In_283,In_1376);
nor U1534 (N_1534,In_108,In_726);
nor U1535 (N_1535,In_1172,In_629);
or U1536 (N_1536,In_1293,In_1258);
and U1537 (N_1537,In_1511,In_1644);
nor U1538 (N_1538,In_1216,In_174);
or U1539 (N_1539,In_1324,In_1254);
or U1540 (N_1540,In_1440,In_667);
nor U1541 (N_1541,In_514,In_1133);
or U1542 (N_1542,In_761,In_457);
and U1543 (N_1543,In_835,In_1594);
xor U1544 (N_1544,In_1752,In_240);
nand U1545 (N_1545,In_1406,In_1201);
and U1546 (N_1546,In_1081,In_918);
nor U1547 (N_1547,In_372,In_1439);
xnor U1548 (N_1548,In_920,In_1893);
nand U1549 (N_1549,In_622,In_212);
or U1550 (N_1550,In_620,In_1184);
nand U1551 (N_1551,In_664,In_957);
or U1552 (N_1552,In_1157,In_180);
nand U1553 (N_1553,In_945,In_781);
nor U1554 (N_1554,In_1467,In_1596);
xnor U1555 (N_1555,In_363,In_1860);
nand U1556 (N_1556,In_1753,In_764);
or U1557 (N_1557,In_1908,In_1378);
nor U1558 (N_1558,In_1201,In_185);
nand U1559 (N_1559,In_269,In_1565);
and U1560 (N_1560,In_873,In_1795);
nor U1561 (N_1561,In_704,In_562);
and U1562 (N_1562,In_864,In_1986);
and U1563 (N_1563,In_914,In_1733);
and U1564 (N_1564,In_1449,In_423);
and U1565 (N_1565,In_815,In_168);
or U1566 (N_1566,In_191,In_290);
xnor U1567 (N_1567,In_210,In_128);
xnor U1568 (N_1568,In_697,In_1616);
xor U1569 (N_1569,In_1877,In_1268);
xnor U1570 (N_1570,In_656,In_1408);
and U1571 (N_1571,In_1746,In_434);
nand U1572 (N_1572,In_533,In_868);
and U1573 (N_1573,In_1002,In_346);
or U1574 (N_1574,In_728,In_1455);
and U1575 (N_1575,In_1802,In_1552);
nand U1576 (N_1576,In_616,In_689);
nand U1577 (N_1577,In_356,In_1171);
nor U1578 (N_1578,In_529,In_756);
and U1579 (N_1579,In_1827,In_403);
nand U1580 (N_1580,In_909,In_499);
and U1581 (N_1581,In_761,In_919);
and U1582 (N_1582,In_1327,In_1554);
nand U1583 (N_1583,In_1875,In_1551);
nand U1584 (N_1584,In_398,In_326);
and U1585 (N_1585,In_1321,In_548);
nor U1586 (N_1586,In_544,In_1518);
nand U1587 (N_1587,In_1775,In_534);
or U1588 (N_1588,In_8,In_449);
and U1589 (N_1589,In_724,In_698);
and U1590 (N_1590,In_1508,In_272);
nand U1591 (N_1591,In_154,In_1477);
nor U1592 (N_1592,In_1723,In_445);
nor U1593 (N_1593,In_873,In_711);
xnor U1594 (N_1594,In_842,In_741);
nand U1595 (N_1595,In_704,In_927);
and U1596 (N_1596,In_785,In_1746);
nand U1597 (N_1597,In_993,In_987);
nand U1598 (N_1598,In_27,In_879);
xor U1599 (N_1599,In_744,In_1599);
and U1600 (N_1600,In_1063,In_58);
nor U1601 (N_1601,In_1042,In_1135);
nand U1602 (N_1602,In_621,In_1414);
or U1603 (N_1603,In_3,In_1237);
nand U1604 (N_1604,In_1200,In_584);
nor U1605 (N_1605,In_1505,In_949);
nand U1606 (N_1606,In_1963,In_331);
and U1607 (N_1607,In_1704,In_288);
nor U1608 (N_1608,In_469,In_101);
and U1609 (N_1609,In_484,In_546);
or U1610 (N_1610,In_691,In_1353);
nand U1611 (N_1611,In_160,In_1143);
nor U1612 (N_1612,In_794,In_186);
or U1613 (N_1613,In_1095,In_570);
or U1614 (N_1614,In_94,In_848);
and U1615 (N_1615,In_1026,In_319);
xor U1616 (N_1616,In_1985,In_183);
and U1617 (N_1617,In_1334,In_1913);
and U1618 (N_1618,In_1826,In_1716);
nand U1619 (N_1619,In_278,In_1583);
nor U1620 (N_1620,In_71,In_1264);
nor U1621 (N_1621,In_818,In_1834);
or U1622 (N_1622,In_405,In_1060);
nor U1623 (N_1623,In_1182,In_1375);
nand U1624 (N_1624,In_1352,In_887);
and U1625 (N_1625,In_1143,In_505);
and U1626 (N_1626,In_956,In_513);
or U1627 (N_1627,In_491,In_1184);
and U1628 (N_1628,In_582,In_1506);
and U1629 (N_1629,In_1642,In_961);
nor U1630 (N_1630,In_718,In_208);
and U1631 (N_1631,In_939,In_964);
and U1632 (N_1632,In_591,In_214);
or U1633 (N_1633,In_1812,In_1912);
xor U1634 (N_1634,In_976,In_513);
xor U1635 (N_1635,In_1536,In_431);
xnor U1636 (N_1636,In_439,In_1598);
and U1637 (N_1637,In_287,In_210);
or U1638 (N_1638,In_1887,In_775);
nand U1639 (N_1639,In_1837,In_95);
and U1640 (N_1640,In_1754,In_1693);
nand U1641 (N_1641,In_1606,In_580);
or U1642 (N_1642,In_1331,In_1964);
nor U1643 (N_1643,In_701,In_794);
and U1644 (N_1644,In_951,In_1313);
and U1645 (N_1645,In_236,In_308);
and U1646 (N_1646,In_1321,In_86);
or U1647 (N_1647,In_698,In_1791);
nor U1648 (N_1648,In_1760,In_994);
nor U1649 (N_1649,In_386,In_1248);
and U1650 (N_1650,In_607,In_1463);
nor U1651 (N_1651,In_1427,In_1780);
nand U1652 (N_1652,In_1972,In_1466);
or U1653 (N_1653,In_1635,In_821);
and U1654 (N_1654,In_821,In_1452);
nand U1655 (N_1655,In_1559,In_789);
nand U1656 (N_1656,In_680,In_1379);
nor U1657 (N_1657,In_595,In_1745);
or U1658 (N_1658,In_1631,In_1711);
and U1659 (N_1659,In_1051,In_1892);
nand U1660 (N_1660,In_1681,In_704);
and U1661 (N_1661,In_1722,In_108);
or U1662 (N_1662,In_416,In_881);
nor U1663 (N_1663,In_954,In_1926);
and U1664 (N_1664,In_1859,In_951);
and U1665 (N_1665,In_1828,In_769);
nor U1666 (N_1666,In_1238,In_515);
and U1667 (N_1667,In_915,In_1122);
or U1668 (N_1668,In_842,In_878);
nand U1669 (N_1669,In_892,In_299);
or U1670 (N_1670,In_1180,In_765);
nor U1671 (N_1671,In_1019,In_417);
nor U1672 (N_1672,In_1871,In_1038);
nand U1673 (N_1673,In_1832,In_1201);
nand U1674 (N_1674,In_854,In_1664);
or U1675 (N_1675,In_1322,In_824);
nor U1676 (N_1676,In_590,In_907);
and U1677 (N_1677,In_547,In_1426);
or U1678 (N_1678,In_431,In_385);
or U1679 (N_1679,In_664,In_124);
nor U1680 (N_1680,In_1599,In_615);
nand U1681 (N_1681,In_1780,In_1309);
xnor U1682 (N_1682,In_1771,In_606);
nor U1683 (N_1683,In_1021,In_900);
and U1684 (N_1684,In_824,In_907);
nand U1685 (N_1685,In_1606,In_1030);
or U1686 (N_1686,In_29,In_800);
and U1687 (N_1687,In_1811,In_204);
or U1688 (N_1688,In_969,In_460);
and U1689 (N_1689,In_912,In_1300);
nand U1690 (N_1690,In_958,In_1645);
and U1691 (N_1691,In_900,In_1056);
xnor U1692 (N_1692,In_1293,In_505);
nor U1693 (N_1693,In_1023,In_386);
and U1694 (N_1694,In_369,In_1732);
and U1695 (N_1695,In_1469,In_1066);
nor U1696 (N_1696,In_1515,In_380);
nand U1697 (N_1697,In_748,In_1695);
and U1698 (N_1698,In_964,In_1555);
xor U1699 (N_1699,In_793,In_1559);
nand U1700 (N_1700,In_118,In_1146);
and U1701 (N_1701,In_1606,In_392);
and U1702 (N_1702,In_1544,In_1559);
nor U1703 (N_1703,In_1185,In_716);
xor U1704 (N_1704,In_1130,In_1110);
or U1705 (N_1705,In_698,In_6);
and U1706 (N_1706,In_704,In_576);
nand U1707 (N_1707,In_1844,In_344);
or U1708 (N_1708,In_487,In_458);
and U1709 (N_1709,In_1915,In_460);
or U1710 (N_1710,In_688,In_1139);
and U1711 (N_1711,In_463,In_863);
or U1712 (N_1712,In_1785,In_1112);
and U1713 (N_1713,In_1256,In_1021);
xor U1714 (N_1714,In_1728,In_598);
or U1715 (N_1715,In_1075,In_1419);
xor U1716 (N_1716,In_1386,In_1968);
and U1717 (N_1717,In_662,In_434);
xor U1718 (N_1718,In_1723,In_43);
or U1719 (N_1719,In_1313,In_453);
nand U1720 (N_1720,In_371,In_641);
or U1721 (N_1721,In_1540,In_97);
and U1722 (N_1722,In_1236,In_473);
xnor U1723 (N_1723,In_886,In_1305);
nand U1724 (N_1724,In_690,In_948);
or U1725 (N_1725,In_1808,In_170);
nand U1726 (N_1726,In_1845,In_1489);
nor U1727 (N_1727,In_217,In_1098);
nor U1728 (N_1728,In_1375,In_1790);
xor U1729 (N_1729,In_1089,In_15);
nor U1730 (N_1730,In_843,In_1128);
and U1731 (N_1731,In_1083,In_261);
or U1732 (N_1732,In_636,In_1246);
and U1733 (N_1733,In_193,In_1445);
or U1734 (N_1734,In_1366,In_761);
and U1735 (N_1735,In_1900,In_1997);
xnor U1736 (N_1736,In_958,In_1894);
nand U1737 (N_1737,In_293,In_1071);
nand U1738 (N_1738,In_472,In_552);
and U1739 (N_1739,In_565,In_285);
xnor U1740 (N_1740,In_1581,In_1132);
or U1741 (N_1741,In_670,In_1471);
and U1742 (N_1742,In_572,In_1396);
nor U1743 (N_1743,In_734,In_652);
or U1744 (N_1744,In_1055,In_1194);
nor U1745 (N_1745,In_1656,In_544);
xnor U1746 (N_1746,In_1059,In_282);
and U1747 (N_1747,In_764,In_1534);
and U1748 (N_1748,In_494,In_1993);
nand U1749 (N_1749,In_297,In_221);
nor U1750 (N_1750,In_1840,In_1988);
nor U1751 (N_1751,In_1007,In_830);
and U1752 (N_1752,In_145,In_616);
or U1753 (N_1753,In_1712,In_1342);
or U1754 (N_1754,In_247,In_1230);
nor U1755 (N_1755,In_392,In_1691);
or U1756 (N_1756,In_534,In_280);
or U1757 (N_1757,In_1392,In_1666);
or U1758 (N_1758,In_1662,In_1925);
and U1759 (N_1759,In_1083,In_281);
nand U1760 (N_1760,In_1932,In_1995);
or U1761 (N_1761,In_468,In_1952);
nand U1762 (N_1762,In_1420,In_305);
nand U1763 (N_1763,In_1723,In_1122);
nor U1764 (N_1764,In_294,In_1068);
nand U1765 (N_1765,In_1638,In_1673);
or U1766 (N_1766,In_256,In_1622);
and U1767 (N_1767,In_538,In_749);
or U1768 (N_1768,In_1204,In_660);
xnor U1769 (N_1769,In_1206,In_15);
or U1770 (N_1770,In_1458,In_1777);
nand U1771 (N_1771,In_1622,In_395);
nor U1772 (N_1772,In_267,In_1396);
and U1773 (N_1773,In_993,In_753);
nor U1774 (N_1774,In_1173,In_955);
nand U1775 (N_1775,In_491,In_1579);
and U1776 (N_1776,In_1938,In_1979);
and U1777 (N_1777,In_1005,In_1302);
xor U1778 (N_1778,In_1943,In_498);
and U1779 (N_1779,In_914,In_1703);
nand U1780 (N_1780,In_920,In_981);
and U1781 (N_1781,In_654,In_1996);
nand U1782 (N_1782,In_1085,In_1940);
or U1783 (N_1783,In_506,In_574);
or U1784 (N_1784,In_62,In_1711);
nor U1785 (N_1785,In_1610,In_608);
nor U1786 (N_1786,In_95,In_841);
nor U1787 (N_1787,In_114,In_42);
and U1788 (N_1788,In_1162,In_234);
nand U1789 (N_1789,In_677,In_689);
and U1790 (N_1790,In_1748,In_1843);
and U1791 (N_1791,In_1164,In_1120);
and U1792 (N_1792,In_226,In_97);
nand U1793 (N_1793,In_575,In_1472);
and U1794 (N_1794,In_632,In_638);
nand U1795 (N_1795,In_1072,In_636);
nor U1796 (N_1796,In_1962,In_1062);
nor U1797 (N_1797,In_374,In_695);
nand U1798 (N_1798,In_1176,In_1365);
and U1799 (N_1799,In_651,In_152);
xor U1800 (N_1800,In_1445,In_1157);
nor U1801 (N_1801,In_101,In_1123);
nand U1802 (N_1802,In_1642,In_1874);
nor U1803 (N_1803,In_1749,In_1440);
or U1804 (N_1804,In_1688,In_1054);
and U1805 (N_1805,In_495,In_1584);
nor U1806 (N_1806,In_546,In_140);
or U1807 (N_1807,In_1098,In_490);
or U1808 (N_1808,In_1909,In_1549);
or U1809 (N_1809,In_1603,In_1785);
and U1810 (N_1810,In_977,In_877);
or U1811 (N_1811,In_156,In_1968);
or U1812 (N_1812,In_66,In_747);
xnor U1813 (N_1813,In_777,In_1400);
or U1814 (N_1814,In_737,In_1598);
nor U1815 (N_1815,In_1128,In_357);
nand U1816 (N_1816,In_79,In_944);
or U1817 (N_1817,In_1172,In_1014);
nor U1818 (N_1818,In_485,In_1313);
xor U1819 (N_1819,In_1104,In_1089);
or U1820 (N_1820,In_231,In_1539);
nand U1821 (N_1821,In_283,In_1675);
nand U1822 (N_1822,In_1200,In_730);
or U1823 (N_1823,In_1680,In_527);
or U1824 (N_1824,In_354,In_1509);
or U1825 (N_1825,In_1499,In_24);
or U1826 (N_1826,In_1710,In_334);
or U1827 (N_1827,In_1730,In_941);
and U1828 (N_1828,In_923,In_742);
nand U1829 (N_1829,In_1618,In_978);
nor U1830 (N_1830,In_960,In_303);
and U1831 (N_1831,In_605,In_415);
or U1832 (N_1832,In_75,In_1207);
nand U1833 (N_1833,In_1529,In_1121);
and U1834 (N_1834,In_1110,In_365);
nand U1835 (N_1835,In_1400,In_729);
nor U1836 (N_1836,In_892,In_435);
nand U1837 (N_1837,In_1483,In_1057);
or U1838 (N_1838,In_1444,In_657);
nand U1839 (N_1839,In_870,In_1554);
and U1840 (N_1840,In_568,In_1389);
or U1841 (N_1841,In_173,In_413);
xnor U1842 (N_1842,In_857,In_14);
or U1843 (N_1843,In_940,In_364);
or U1844 (N_1844,In_317,In_1758);
nand U1845 (N_1845,In_750,In_646);
xor U1846 (N_1846,In_1456,In_1817);
nor U1847 (N_1847,In_1269,In_743);
xor U1848 (N_1848,In_1424,In_1003);
or U1849 (N_1849,In_357,In_1837);
or U1850 (N_1850,In_1962,In_1820);
nand U1851 (N_1851,In_1839,In_902);
and U1852 (N_1852,In_878,In_1769);
and U1853 (N_1853,In_897,In_1386);
nor U1854 (N_1854,In_1255,In_649);
nor U1855 (N_1855,In_140,In_511);
and U1856 (N_1856,In_745,In_792);
nand U1857 (N_1857,In_461,In_544);
and U1858 (N_1858,In_510,In_617);
nor U1859 (N_1859,In_138,In_1333);
nand U1860 (N_1860,In_1071,In_1654);
and U1861 (N_1861,In_916,In_880);
or U1862 (N_1862,In_1408,In_1630);
or U1863 (N_1863,In_1393,In_514);
nor U1864 (N_1864,In_1838,In_585);
xnor U1865 (N_1865,In_1972,In_774);
or U1866 (N_1866,In_1242,In_1134);
nand U1867 (N_1867,In_1214,In_1164);
or U1868 (N_1868,In_1904,In_726);
or U1869 (N_1869,In_1720,In_1144);
nor U1870 (N_1870,In_516,In_1078);
nor U1871 (N_1871,In_177,In_711);
nand U1872 (N_1872,In_1546,In_1655);
nor U1873 (N_1873,In_67,In_883);
nand U1874 (N_1874,In_655,In_1943);
nor U1875 (N_1875,In_450,In_1774);
and U1876 (N_1876,In_1432,In_21);
nor U1877 (N_1877,In_1462,In_1129);
and U1878 (N_1878,In_1724,In_1152);
and U1879 (N_1879,In_498,In_999);
and U1880 (N_1880,In_281,In_1712);
nand U1881 (N_1881,In_622,In_1160);
xnor U1882 (N_1882,In_1396,In_1157);
nor U1883 (N_1883,In_427,In_982);
nand U1884 (N_1884,In_1807,In_422);
xor U1885 (N_1885,In_744,In_1076);
nand U1886 (N_1886,In_824,In_773);
or U1887 (N_1887,In_900,In_1652);
or U1888 (N_1888,In_1141,In_1402);
nor U1889 (N_1889,In_1072,In_1117);
or U1890 (N_1890,In_137,In_1395);
nor U1891 (N_1891,In_1298,In_1726);
nand U1892 (N_1892,In_891,In_1816);
nor U1893 (N_1893,In_1949,In_768);
nor U1894 (N_1894,In_1914,In_1456);
nand U1895 (N_1895,In_1464,In_519);
nand U1896 (N_1896,In_219,In_1650);
or U1897 (N_1897,In_327,In_1666);
nand U1898 (N_1898,In_1315,In_736);
xor U1899 (N_1899,In_329,In_393);
nand U1900 (N_1900,In_713,In_1602);
xor U1901 (N_1901,In_1051,In_1700);
or U1902 (N_1902,In_1588,In_1520);
and U1903 (N_1903,In_240,In_579);
and U1904 (N_1904,In_873,In_85);
and U1905 (N_1905,In_1060,In_1471);
nor U1906 (N_1906,In_890,In_1816);
nand U1907 (N_1907,In_502,In_1082);
nand U1908 (N_1908,In_791,In_206);
or U1909 (N_1909,In_1735,In_1823);
and U1910 (N_1910,In_109,In_225);
nand U1911 (N_1911,In_1488,In_1678);
nor U1912 (N_1912,In_1854,In_125);
and U1913 (N_1913,In_1308,In_737);
nand U1914 (N_1914,In_1201,In_167);
and U1915 (N_1915,In_1194,In_1126);
and U1916 (N_1916,In_1156,In_403);
nor U1917 (N_1917,In_695,In_1562);
or U1918 (N_1918,In_521,In_675);
or U1919 (N_1919,In_680,In_597);
nor U1920 (N_1920,In_1053,In_651);
nand U1921 (N_1921,In_1577,In_1367);
nor U1922 (N_1922,In_1563,In_513);
and U1923 (N_1923,In_1802,In_1941);
and U1924 (N_1924,In_414,In_1293);
and U1925 (N_1925,In_1042,In_61);
xor U1926 (N_1926,In_845,In_791);
or U1927 (N_1927,In_1728,In_1480);
nand U1928 (N_1928,In_860,In_1412);
nand U1929 (N_1929,In_1758,In_199);
nor U1930 (N_1930,In_1962,In_1173);
and U1931 (N_1931,In_1614,In_1980);
and U1932 (N_1932,In_190,In_1993);
nor U1933 (N_1933,In_987,In_1182);
xor U1934 (N_1934,In_954,In_1486);
nor U1935 (N_1935,In_928,In_976);
and U1936 (N_1936,In_121,In_1117);
and U1937 (N_1937,In_1154,In_536);
xor U1938 (N_1938,In_584,In_1833);
nor U1939 (N_1939,In_1053,In_1995);
nand U1940 (N_1940,In_930,In_287);
nor U1941 (N_1941,In_705,In_363);
and U1942 (N_1942,In_699,In_1997);
or U1943 (N_1943,In_820,In_1585);
and U1944 (N_1944,In_1071,In_1978);
and U1945 (N_1945,In_1566,In_1688);
nand U1946 (N_1946,In_1774,In_1541);
or U1947 (N_1947,In_1349,In_1572);
nor U1948 (N_1948,In_7,In_1695);
or U1949 (N_1949,In_846,In_1762);
nor U1950 (N_1950,In_1228,In_1976);
nand U1951 (N_1951,In_737,In_403);
and U1952 (N_1952,In_506,In_1235);
nand U1953 (N_1953,In_1060,In_970);
or U1954 (N_1954,In_1022,In_1566);
and U1955 (N_1955,In_1891,In_1133);
xnor U1956 (N_1956,In_360,In_1653);
nand U1957 (N_1957,In_1130,In_166);
xor U1958 (N_1958,In_1900,In_1848);
nor U1959 (N_1959,In_544,In_163);
and U1960 (N_1960,In_1374,In_816);
nor U1961 (N_1961,In_324,In_1282);
or U1962 (N_1962,In_172,In_1389);
nand U1963 (N_1963,In_1070,In_813);
xor U1964 (N_1964,In_1025,In_718);
nor U1965 (N_1965,In_638,In_1589);
and U1966 (N_1966,In_803,In_1350);
nor U1967 (N_1967,In_1064,In_1355);
xor U1968 (N_1968,In_1563,In_1433);
xnor U1969 (N_1969,In_347,In_651);
nor U1970 (N_1970,In_1999,In_706);
nand U1971 (N_1971,In_1344,In_1888);
nor U1972 (N_1972,In_959,In_267);
xnor U1973 (N_1973,In_1009,In_641);
nor U1974 (N_1974,In_1609,In_852);
and U1975 (N_1975,In_1525,In_1262);
and U1976 (N_1976,In_273,In_395);
and U1977 (N_1977,In_224,In_918);
nand U1978 (N_1978,In_1325,In_591);
nor U1979 (N_1979,In_912,In_1724);
and U1980 (N_1980,In_1115,In_1972);
or U1981 (N_1981,In_16,In_513);
or U1982 (N_1982,In_331,In_1127);
and U1983 (N_1983,In_206,In_392);
or U1984 (N_1984,In_1894,In_1823);
xnor U1985 (N_1985,In_97,In_227);
nand U1986 (N_1986,In_59,In_1474);
or U1987 (N_1987,In_1181,In_136);
or U1988 (N_1988,In_1092,In_1720);
xor U1989 (N_1989,In_861,In_71);
nand U1990 (N_1990,In_1481,In_227);
and U1991 (N_1991,In_280,In_630);
xnor U1992 (N_1992,In_1044,In_529);
nor U1993 (N_1993,In_1845,In_204);
or U1994 (N_1994,In_1405,In_1966);
xnor U1995 (N_1995,In_247,In_1274);
or U1996 (N_1996,In_1566,In_84);
nand U1997 (N_1997,In_1915,In_1919);
xor U1998 (N_1998,In_811,In_1601);
and U1999 (N_1999,In_251,In_206);
and U2000 (N_2000,In_1154,In_1171);
nor U2001 (N_2001,In_680,In_1082);
nor U2002 (N_2002,In_1886,In_1385);
and U2003 (N_2003,In_274,In_1414);
or U2004 (N_2004,In_382,In_783);
or U2005 (N_2005,In_389,In_339);
or U2006 (N_2006,In_589,In_179);
or U2007 (N_2007,In_1726,In_1463);
and U2008 (N_2008,In_1821,In_895);
or U2009 (N_2009,In_317,In_1162);
or U2010 (N_2010,In_1329,In_66);
and U2011 (N_2011,In_1215,In_1190);
and U2012 (N_2012,In_1520,In_1944);
nand U2013 (N_2013,In_233,In_690);
nor U2014 (N_2014,In_734,In_1807);
and U2015 (N_2015,In_305,In_368);
or U2016 (N_2016,In_715,In_846);
and U2017 (N_2017,In_1933,In_615);
nand U2018 (N_2018,In_1459,In_140);
nor U2019 (N_2019,In_286,In_1726);
or U2020 (N_2020,In_388,In_297);
nor U2021 (N_2021,In_501,In_570);
nand U2022 (N_2022,In_1421,In_1204);
or U2023 (N_2023,In_1785,In_433);
nand U2024 (N_2024,In_945,In_1880);
nand U2025 (N_2025,In_368,In_542);
nor U2026 (N_2026,In_320,In_796);
or U2027 (N_2027,In_741,In_352);
or U2028 (N_2028,In_337,In_1631);
nand U2029 (N_2029,In_1367,In_846);
or U2030 (N_2030,In_838,In_693);
and U2031 (N_2031,In_1379,In_350);
xor U2032 (N_2032,In_476,In_397);
and U2033 (N_2033,In_601,In_1637);
nand U2034 (N_2034,In_1785,In_114);
and U2035 (N_2035,In_664,In_1690);
xor U2036 (N_2036,In_37,In_1090);
or U2037 (N_2037,In_117,In_1928);
nand U2038 (N_2038,In_1991,In_4);
and U2039 (N_2039,In_1123,In_1375);
nor U2040 (N_2040,In_1576,In_1949);
nand U2041 (N_2041,In_1334,In_258);
nor U2042 (N_2042,In_421,In_1310);
xnor U2043 (N_2043,In_529,In_1351);
nor U2044 (N_2044,In_257,In_455);
nor U2045 (N_2045,In_539,In_1402);
nor U2046 (N_2046,In_201,In_921);
or U2047 (N_2047,In_702,In_875);
or U2048 (N_2048,In_1462,In_129);
or U2049 (N_2049,In_1928,In_327);
and U2050 (N_2050,In_472,In_1912);
xor U2051 (N_2051,In_795,In_749);
nor U2052 (N_2052,In_713,In_255);
and U2053 (N_2053,In_136,In_1920);
and U2054 (N_2054,In_1067,In_335);
or U2055 (N_2055,In_74,In_110);
nand U2056 (N_2056,In_200,In_126);
xnor U2057 (N_2057,In_513,In_159);
nor U2058 (N_2058,In_975,In_1895);
nor U2059 (N_2059,In_1048,In_869);
and U2060 (N_2060,In_1324,In_1644);
nand U2061 (N_2061,In_87,In_69);
or U2062 (N_2062,In_415,In_807);
nor U2063 (N_2063,In_54,In_13);
nand U2064 (N_2064,In_1082,In_1186);
or U2065 (N_2065,In_353,In_1687);
or U2066 (N_2066,In_1877,In_1211);
nand U2067 (N_2067,In_638,In_1504);
or U2068 (N_2068,In_899,In_927);
or U2069 (N_2069,In_429,In_635);
nand U2070 (N_2070,In_1703,In_21);
nor U2071 (N_2071,In_1433,In_1581);
or U2072 (N_2072,In_205,In_1503);
nor U2073 (N_2073,In_437,In_1307);
xnor U2074 (N_2074,In_1731,In_1056);
nor U2075 (N_2075,In_402,In_361);
and U2076 (N_2076,In_1783,In_1044);
or U2077 (N_2077,In_962,In_20);
nor U2078 (N_2078,In_855,In_268);
and U2079 (N_2079,In_312,In_1835);
and U2080 (N_2080,In_1663,In_1166);
or U2081 (N_2081,In_501,In_1943);
nor U2082 (N_2082,In_645,In_276);
nand U2083 (N_2083,In_767,In_923);
xor U2084 (N_2084,In_1092,In_608);
nand U2085 (N_2085,In_1481,In_1880);
xnor U2086 (N_2086,In_538,In_90);
xnor U2087 (N_2087,In_1335,In_207);
nand U2088 (N_2088,In_1552,In_86);
and U2089 (N_2089,In_374,In_1636);
nor U2090 (N_2090,In_1945,In_1617);
nor U2091 (N_2091,In_1743,In_1758);
or U2092 (N_2092,In_1751,In_538);
nor U2093 (N_2093,In_175,In_1618);
and U2094 (N_2094,In_409,In_612);
and U2095 (N_2095,In_421,In_765);
and U2096 (N_2096,In_1194,In_1705);
and U2097 (N_2097,In_191,In_1234);
nor U2098 (N_2098,In_999,In_1270);
and U2099 (N_2099,In_507,In_723);
nand U2100 (N_2100,In_1415,In_791);
nand U2101 (N_2101,In_594,In_562);
and U2102 (N_2102,In_160,In_1218);
or U2103 (N_2103,In_1120,In_705);
nor U2104 (N_2104,In_1922,In_1907);
or U2105 (N_2105,In_1646,In_451);
nor U2106 (N_2106,In_1292,In_1525);
nand U2107 (N_2107,In_931,In_1780);
nor U2108 (N_2108,In_832,In_245);
or U2109 (N_2109,In_1910,In_786);
and U2110 (N_2110,In_1071,In_1833);
nand U2111 (N_2111,In_1011,In_943);
nand U2112 (N_2112,In_725,In_1979);
or U2113 (N_2113,In_1755,In_76);
nand U2114 (N_2114,In_402,In_397);
or U2115 (N_2115,In_1400,In_1773);
nor U2116 (N_2116,In_1438,In_86);
or U2117 (N_2117,In_1585,In_1549);
nor U2118 (N_2118,In_381,In_373);
nor U2119 (N_2119,In_330,In_1160);
or U2120 (N_2120,In_1272,In_697);
and U2121 (N_2121,In_496,In_346);
and U2122 (N_2122,In_1201,In_1653);
or U2123 (N_2123,In_172,In_1266);
or U2124 (N_2124,In_156,In_1168);
or U2125 (N_2125,In_1516,In_536);
nor U2126 (N_2126,In_1050,In_123);
or U2127 (N_2127,In_640,In_265);
nor U2128 (N_2128,In_483,In_974);
nand U2129 (N_2129,In_431,In_776);
nand U2130 (N_2130,In_1876,In_33);
xor U2131 (N_2131,In_331,In_131);
and U2132 (N_2132,In_1974,In_1050);
and U2133 (N_2133,In_1996,In_1961);
and U2134 (N_2134,In_1075,In_1103);
nor U2135 (N_2135,In_387,In_505);
nor U2136 (N_2136,In_1094,In_362);
nor U2137 (N_2137,In_304,In_636);
or U2138 (N_2138,In_1792,In_793);
nand U2139 (N_2139,In_1935,In_0);
or U2140 (N_2140,In_221,In_1891);
nor U2141 (N_2141,In_1173,In_1801);
or U2142 (N_2142,In_1306,In_276);
or U2143 (N_2143,In_1227,In_176);
nor U2144 (N_2144,In_1213,In_1770);
nor U2145 (N_2145,In_1121,In_852);
nor U2146 (N_2146,In_833,In_501);
nand U2147 (N_2147,In_1086,In_1545);
nand U2148 (N_2148,In_1126,In_1048);
and U2149 (N_2149,In_1269,In_296);
nand U2150 (N_2150,In_141,In_1971);
nor U2151 (N_2151,In_1808,In_1543);
xor U2152 (N_2152,In_17,In_1636);
and U2153 (N_2153,In_1711,In_735);
and U2154 (N_2154,In_207,In_1645);
nor U2155 (N_2155,In_1198,In_1723);
and U2156 (N_2156,In_1022,In_777);
xnor U2157 (N_2157,In_1343,In_1954);
nor U2158 (N_2158,In_390,In_403);
or U2159 (N_2159,In_955,In_1762);
nand U2160 (N_2160,In_1129,In_826);
and U2161 (N_2161,In_1554,In_1595);
nor U2162 (N_2162,In_977,In_1005);
nor U2163 (N_2163,In_1896,In_949);
or U2164 (N_2164,In_1785,In_291);
nor U2165 (N_2165,In_472,In_1145);
nor U2166 (N_2166,In_147,In_856);
or U2167 (N_2167,In_1662,In_1989);
nor U2168 (N_2168,In_1945,In_1202);
and U2169 (N_2169,In_1071,In_1441);
and U2170 (N_2170,In_144,In_1770);
nor U2171 (N_2171,In_359,In_1830);
and U2172 (N_2172,In_313,In_741);
or U2173 (N_2173,In_1563,In_1625);
and U2174 (N_2174,In_1672,In_199);
and U2175 (N_2175,In_700,In_306);
and U2176 (N_2176,In_827,In_1410);
or U2177 (N_2177,In_684,In_1997);
nor U2178 (N_2178,In_532,In_1074);
and U2179 (N_2179,In_607,In_6);
or U2180 (N_2180,In_993,In_808);
xnor U2181 (N_2181,In_448,In_4);
and U2182 (N_2182,In_1185,In_268);
nand U2183 (N_2183,In_290,In_1682);
nand U2184 (N_2184,In_245,In_840);
and U2185 (N_2185,In_1168,In_1278);
and U2186 (N_2186,In_1705,In_1451);
nand U2187 (N_2187,In_663,In_1242);
nand U2188 (N_2188,In_141,In_1623);
and U2189 (N_2189,In_926,In_1767);
xor U2190 (N_2190,In_1004,In_1162);
or U2191 (N_2191,In_951,In_1833);
nand U2192 (N_2192,In_1635,In_447);
nand U2193 (N_2193,In_1981,In_1347);
nor U2194 (N_2194,In_1475,In_1151);
or U2195 (N_2195,In_1885,In_1269);
nor U2196 (N_2196,In_1290,In_486);
and U2197 (N_2197,In_1565,In_1258);
nor U2198 (N_2198,In_1346,In_1124);
xor U2199 (N_2199,In_1901,In_624);
xor U2200 (N_2200,In_31,In_1364);
nor U2201 (N_2201,In_1227,In_1402);
nor U2202 (N_2202,In_397,In_419);
xor U2203 (N_2203,In_169,In_193);
xnor U2204 (N_2204,In_799,In_1291);
and U2205 (N_2205,In_1529,In_16);
nor U2206 (N_2206,In_572,In_386);
or U2207 (N_2207,In_1396,In_1266);
nor U2208 (N_2208,In_1780,In_1246);
or U2209 (N_2209,In_1006,In_558);
nor U2210 (N_2210,In_129,In_125);
and U2211 (N_2211,In_659,In_1422);
nand U2212 (N_2212,In_1004,In_56);
and U2213 (N_2213,In_380,In_1050);
nand U2214 (N_2214,In_414,In_304);
or U2215 (N_2215,In_34,In_1573);
and U2216 (N_2216,In_1613,In_1137);
nand U2217 (N_2217,In_1440,In_443);
nor U2218 (N_2218,In_953,In_199);
nor U2219 (N_2219,In_1518,In_1043);
nor U2220 (N_2220,In_1324,In_1911);
nor U2221 (N_2221,In_521,In_1564);
and U2222 (N_2222,In_66,In_1265);
nand U2223 (N_2223,In_1368,In_1956);
and U2224 (N_2224,In_956,In_741);
and U2225 (N_2225,In_746,In_1111);
and U2226 (N_2226,In_158,In_108);
xnor U2227 (N_2227,In_1913,In_1642);
nor U2228 (N_2228,In_959,In_662);
nor U2229 (N_2229,In_410,In_638);
or U2230 (N_2230,In_1479,In_1186);
or U2231 (N_2231,In_707,In_1150);
or U2232 (N_2232,In_591,In_134);
nor U2233 (N_2233,In_508,In_64);
nor U2234 (N_2234,In_740,In_1732);
or U2235 (N_2235,In_1051,In_404);
and U2236 (N_2236,In_1627,In_1940);
xnor U2237 (N_2237,In_467,In_815);
and U2238 (N_2238,In_90,In_207);
or U2239 (N_2239,In_917,In_1021);
or U2240 (N_2240,In_289,In_302);
xor U2241 (N_2241,In_680,In_1810);
nand U2242 (N_2242,In_1850,In_1);
or U2243 (N_2243,In_493,In_1861);
nand U2244 (N_2244,In_1972,In_286);
and U2245 (N_2245,In_1028,In_1216);
nor U2246 (N_2246,In_324,In_617);
nand U2247 (N_2247,In_1243,In_807);
and U2248 (N_2248,In_1428,In_935);
and U2249 (N_2249,In_756,In_1440);
nand U2250 (N_2250,In_1815,In_326);
nor U2251 (N_2251,In_788,In_421);
and U2252 (N_2252,In_1522,In_1318);
nor U2253 (N_2253,In_446,In_1143);
and U2254 (N_2254,In_1619,In_1091);
and U2255 (N_2255,In_1868,In_49);
nand U2256 (N_2256,In_1898,In_1421);
nand U2257 (N_2257,In_1064,In_422);
nor U2258 (N_2258,In_1526,In_966);
nor U2259 (N_2259,In_495,In_309);
and U2260 (N_2260,In_1173,In_142);
and U2261 (N_2261,In_1168,In_766);
xnor U2262 (N_2262,In_637,In_1246);
and U2263 (N_2263,In_946,In_1193);
and U2264 (N_2264,In_1500,In_1238);
or U2265 (N_2265,In_592,In_575);
nor U2266 (N_2266,In_1404,In_1567);
and U2267 (N_2267,In_974,In_560);
nor U2268 (N_2268,In_1205,In_1858);
or U2269 (N_2269,In_1784,In_0);
xnor U2270 (N_2270,In_703,In_30);
nor U2271 (N_2271,In_913,In_700);
or U2272 (N_2272,In_265,In_1551);
nor U2273 (N_2273,In_331,In_1659);
nand U2274 (N_2274,In_1927,In_862);
and U2275 (N_2275,In_1000,In_1585);
nand U2276 (N_2276,In_271,In_1158);
nor U2277 (N_2277,In_1342,In_936);
or U2278 (N_2278,In_703,In_1665);
or U2279 (N_2279,In_577,In_804);
and U2280 (N_2280,In_573,In_752);
or U2281 (N_2281,In_781,In_1502);
nor U2282 (N_2282,In_546,In_1535);
nor U2283 (N_2283,In_1808,In_1885);
nor U2284 (N_2284,In_1750,In_826);
or U2285 (N_2285,In_610,In_667);
xor U2286 (N_2286,In_551,In_1190);
or U2287 (N_2287,In_670,In_1711);
and U2288 (N_2288,In_1850,In_568);
or U2289 (N_2289,In_282,In_255);
and U2290 (N_2290,In_604,In_1111);
nand U2291 (N_2291,In_1123,In_6);
or U2292 (N_2292,In_407,In_153);
nor U2293 (N_2293,In_374,In_1654);
and U2294 (N_2294,In_1108,In_471);
nor U2295 (N_2295,In_1112,In_213);
nand U2296 (N_2296,In_1067,In_26);
or U2297 (N_2297,In_883,In_1568);
nor U2298 (N_2298,In_1282,In_334);
nor U2299 (N_2299,In_1208,In_1709);
and U2300 (N_2300,In_725,In_1492);
and U2301 (N_2301,In_739,In_1046);
xor U2302 (N_2302,In_1219,In_652);
nor U2303 (N_2303,In_83,In_178);
nor U2304 (N_2304,In_556,In_224);
and U2305 (N_2305,In_1081,In_943);
or U2306 (N_2306,In_1270,In_1346);
nor U2307 (N_2307,In_1398,In_1472);
and U2308 (N_2308,In_1459,In_1242);
nand U2309 (N_2309,In_301,In_1202);
or U2310 (N_2310,In_298,In_1304);
nand U2311 (N_2311,In_583,In_1045);
or U2312 (N_2312,In_937,In_712);
nand U2313 (N_2313,In_1160,In_1910);
and U2314 (N_2314,In_1901,In_1700);
nor U2315 (N_2315,In_490,In_684);
and U2316 (N_2316,In_1094,In_209);
nand U2317 (N_2317,In_1899,In_1841);
nand U2318 (N_2318,In_252,In_1436);
nor U2319 (N_2319,In_294,In_184);
nor U2320 (N_2320,In_183,In_1364);
and U2321 (N_2321,In_1656,In_1503);
and U2322 (N_2322,In_1482,In_1666);
or U2323 (N_2323,In_1842,In_1975);
or U2324 (N_2324,In_821,In_1541);
nand U2325 (N_2325,In_1495,In_827);
nor U2326 (N_2326,In_1842,In_906);
or U2327 (N_2327,In_908,In_1024);
nor U2328 (N_2328,In_685,In_722);
xor U2329 (N_2329,In_1516,In_1632);
and U2330 (N_2330,In_1320,In_1114);
and U2331 (N_2331,In_360,In_641);
nand U2332 (N_2332,In_1283,In_852);
nor U2333 (N_2333,In_1825,In_594);
or U2334 (N_2334,In_441,In_1674);
and U2335 (N_2335,In_271,In_1980);
nand U2336 (N_2336,In_466,In_563);
or U2337 (N_2337,In_902,In_324);
nand U2338 (N_2338,In_738,In_1679);
nor U2339 (N_2339,In_313,In_1942);
and U2340 (N_2340,In_1632,In_687);
or U2341 (N_2341,In_1711,In_726);
nand U2342 (N_2342,In_347,In_1473);
xor U2343 (N_2343,In_1837,In_1051);
nor U2344 (N_2344,In_1337,In_1857);
or U2345 (N_2345,In_1777,In_447);
and U2346 (N_2346,In_858,In_913);
and U2347 (N_2347,In_92,In_705);
nand U2348 (N_2348,In_884,In_241);
nand U2349 (N_2349,In_894,In_303);
and U2350 (N_2350,In_14,In_1272);
and U2351 (N_2351,In_1249,In_717);
nor U2352 (N_2352,In_1728,In_1934);
or U2353 (N_2353,In_1702,In_1022);
and U2354 (N_2354,In_1017,In_554);
nor U2355 (N_2355,In_599,In_146);
nand U2356 (N_2356,In_1828,In_1249);
nor U2357 (N_2357,In_951,In_264);
nor U2358 (N_2358,In_1762,In_51);
xnor U2359 (N_2359,In_541,In_662);
or U2360 (N_2360,In_1158,In_1663);
and U2361 (N_2361,In_1985,In_1939);
or U2362 (N_2362,In_521,In_589);
or U2363 (N_2363,In_1866,In_885);
or U2364 (N_2364,In_1112,In_457);
or U2365 (N_2365,In_252,In_1248);
or U2366 (N_2366,In_1305,In_751);
xnor U2367 (N_2367,In_787,In_1299);
nor U2368 (N_2368,In_1970,In_1090);
or U2369 (N_2369,In_1650,In_1626);
and U2370 (N_2370,In_895,In_909);
nor U2371 (N_2371,In_1814,In_1844);
or U2372 (N_2372,In_3,In_1315);
and U2373 (N_2373,In_1391,In_1549);
nand U2374 (N_2374,In_883,In_1131);
or U2375 (N_2375,In_928,In_1485);
nand U2376 (N_2376,In_564,In_1946);
nor U2377 (N_2377,In_1203,In_306);
nand U2378 (N_2378,In_670,In_461);
nand U2379 (N_2379,In_548,In_1120);
nand U2380 (N_2380,In_415,In_1584);
xor U2381 (N_2381,In_664,In_421);
or U2382 (N_2382,In_1913,In_1967);
nand U2383 (N_2383,In_812,In_1664);
nor U2384 (N_2384,In_1037,In_1337);
and U2385 (N_2385,In_1897,In_1763);
xnor U2386 (N_2386,In_1962,In_1220);
nand U2387 (N_2387,In_360,In_883);
nor U2388 (N_2388,In_667,In_1672);
or U2389 (N_2389,In_846,In_434);
nand U2390 (N_2390,In_1022,In_1796);
or U2391 (N_2391,In_44,In_875);
nor U2392 (N_2392,In_185,In_1746);
and U2393 (N_2393,In_968,In_1253);
or U2394 (N_2394,In_385,In_987);
and U2395 (N_2395,In_246,In_554);
or U2396 (N_2396,In_1578,In_1282);
and U2397 (N_2397,In_598,In_299);
and U2398 (N_2398,In_1464,In_472);
xnor U2399 (N_2399,In_1875,In_324);
nor U2400 (N_2400,In_1857,In_382);
nor U2401 (N_2401,In_1144,In_175);
nor U2402 (N_2402,In_469,In_565);
or U2403 (N_2403,In_118,In_273);
nand U2404 (N_2404,In_1665,In_1779);
and U2405 (N_2405,In_1659,In_1649);
nand U2406 (N_2406,In_561,In_1849);
nand U2407 (N_2407,In_110,In_1165);
and U2408 (N_2408,In_417,In_1767);
or U2409 (N_2409,In_1031,In_335);
xor U2410 (N_2410,In_12,In_1721);
or U2411 (N_2411,In_1796,In_1103);
xor U2412 (N_2412,In_1987,In_1413);
and U2413 (N_2413,In_1904,In_1591);
or U2414 (N_2414,In_5,In_1624);
nand U2415 (N_2415,In_1141,In_470);
nand U2416 (N_2416,In_1881,In_1103);
or U2417 (N_2417,In_706,In_1714);
nand U2418 (N_2418,In_1142,In_427);
nor U2419 (N_2419,In_1747,In_113);
xor U2420 (N_2420,In_1825,In_1700);
or U2421 (N_2421,In_753,In_1251);
or U2422 (N_2422,In_905,In_1488);
or U2423 (N_2423,In_1438,In_1481);
and U2424 (N_2424,In_1616,In_264);
xor U2425 (N_2425,In_679,In_1906);
nor U2426 (N_2426,In_307,In_1139);
and U2427 (N_2427,In_1388,In_1493);
or U2428 (N_2428,In_913,In_1866);
and U2429 (N_2429,In_1823,In_692);
and U2430 (N_2430,In_997,In_1322);
or U2431 (N_2431,In_1735,In_825);
or U2432 (N_2432,In_356,In_84);
and U2433 (N_2433,In_1544,In_1550);
nor U2434 (N_2434,In_1653,In_1533);
and U2435 (N_2435,In_1577,In_927);
or U2436 (N_2436,In_1772,In_110);
and U2437 (N_2437,In_775,In_1620);
nand U2438 (N_2438,In_1189,In_615);
or U2439 (N_2439,In_883,In_1886);
and U2440 (N_2440,In_227,In_1952);
or U2441 (N_2441,In_477,In_1942);
nand U2442 (N_2442,In_127,In_1099);
and U2443 (N_2443,In_193,In_837);
nand U2444 (N_2444,In_1069,In_1064);
or U2445 (N_2445,In_865,In_1247);
xnor U2446 (N_2446,In_606,In_516);
nand U2447 (N_2447,In_1834,In_1193);
or U2448 (N_2448,In_1376,In_1385);
nand U2449 (N_2449,In_1559,In_212);
nor U2450 (N_2450,In_883,In_1342);
nor U2451 (N_2451,In_832,In_248);
and U2452 (N_2452,In_772,In_1047);
and U2453 (N_2453,In_1946,In_838);
and U2454 (N_2454,In_624,In_1313);
xor U2455 (N_2455,In_1757,In_383);
or U2456 (N_2456,In_1851,In_45);
xnor U2457 (N_2457,In_1417,In_1491);
nor U2458 (N_2458,In_1020,In_1533);
xnor U2459 (N_2459,In_1898,In_974);
nand U2460 (N_2460,In_1156,In_689);
and U2461 (N_2461,In_419,In_14);
and U2462 (N_2462,In_1191,In_1464);
nand U2463 (N_2463,In_1872,In_995);
or U2464 (N_2464,In_298,In_1405);
xnor U2465 (N_2465,In_673,In_650);
nor U2466 (N_2466,In_1712,In_1213);
nand U2467 (N_2467,In_46,In_482);
nor U2468 (N_2468,In_1650,In_563);
or U2469 (N_2469,In_1607,In_55);
or U2470 (N_2470,In_400,In_1024);
or U2471 (N_2471,In_1704,In_1559);
nand U2472 (N_2472,In_1507,In_1584);
nand U2473 (N_2473,In_1678,In_1525);
or U2474 (N_2474,In_1563,In_1345);
or U2475 (N_2475,In_1140,In_772);
or U2476 (N_2476,In_1659,In_284);
nor U2477 (N_2477,In_758,In_231);
or U2478 (N_2478,In_590,In_457);
nand U2479 (N_2479,In_1654,In_1166);
nand U2480 (N_2480,In_593,In_116);
nand U2481 (N_2481,In_70,In_772);
nand U2482 (N_2482,In_19,In_890);
nor U2483 (N_2483,In_1817,In_191);
or U2484 (N_2484,In_1163,In_1569);
nand U2485 (N_2485,In_295,In_133);
or U2486 (N_2486,In_1270,In_1513);
and U2487 (N_2487,In_320,In_945);
and U2488 (N_2488,In_623,In_1988);
xnor U2489 (N_2489,In_671,In_756);
or U2490 (N_2490,In_1645,In_540);
or U2491 (N_2491,In_934,In_1710);
and U2492 (N_2492,In_1264,In_773);
nor U2493 (N_2493,In_1351,In_94);
or U2494 (N_2494,In_1152,In_1620);
and U2495 (N_2495,In_1896,In_528);
and U2496 (N_2496,In_1901,In_988);
or U2497 (N_2497,In_1465,In_1675);
and U2498 (N_2498,In_1374,In_1370);
nor U2499 (N_2499,In_1781,In_1946);
nand U2500 (N_2500,In_1613,In_996);
nor U2501 (N_2501,In_277,In_1081);
or U2502 (N_2502,In_351,In_34);
and U2503 (N_2503,In_138,In_1703);
or U2504 (N_2504,In_504,In_121);
and U2505 (N_2505,In_1316,In_1910);
xor U2506 (N_2506,In_1363,In_1382);
or U2507 (N_2507,In_1019,In_282);
or U2508 (N_2508,In_1010,In_247);
nand U2509 (N_2509,In_98,In_674);
and U2510 (N_2510,In_1271,In_409);
nand U2511 (N_2511,In_941,In_1992);
or U2512 (N_2512,In_1756,In_1967);
nor U2513 (N_2513,In_422,In_725);
and U2514 (N_2514,In_1332,In_1779);
nor U2515 (N_2515,In_587,In_1729);
and U2516 (N_2516,In_853,In_386);
and U2517 (N_2517,In_150,In_1153);
or U2518 (N_2518,In_1247,In_993);
nor U2519 (N_2519,In_1466,In_1359);
or U2520 (N_2520,In_1701,In_674);
and U2521 (N_2521,In_1270,In_677);
nand U2522 (N_2522,In_741,In_928);
nor U2523 (N_2523,In_1624,In_1238);
or U2524 (N_2524,In_1237,In_237);
nand U2525 (N_2525,In_1120,In_1497);
and U2526 (N_2526,In_1854,In_238);
or U2527 (N_2527,In_638,In_800);
and U2528 (N_2528,In_1771,In_479);
nor U2529 (N_2529,In_414,In_1089);
nor U2530 (N_2530,In_337,In_1023);
nor U2531 (N_2531,In_1504,In_70);
nor U2532 (N_2532,In_489,In_713);
nor U2533 (N_2533,In_1124,In_1161);
nor U2534 (N_2534,In_389,In_1607);
xor U2535 (N_2535,In_1329,In_1513);
and U2536 (N_2536,In_1783,In_334);
nand U2537 (N_2537,In_983,In_1561);
nor U2538 (N_2538,In_1009,In_1752);
or U2539 (N_2539,In_59,In_1289);
nor U2540 (N_2540,In_660,In_1914);
nand U2541 (N_2541,In_1544,In_1598);
and U2542 (N_2542,In_1683,In_141);
and U2543 (N_2543,In_324,In_1202);
and U2544 (N_2544,In_1462,In_257);
nand U2545 (N_2545,In_229,In_1705);
or U2546 (N_2546,In_265,In_992);
nand U2547 (N_2547,In_1463,In_913);
xor U2548 (N_2548,In_753,In_1571);
nor U2549 (N_2549,In_1696,In_430);
nor U2550 (N_2550,In_1731,In_977);
xnor U2551 (N_2551,In_1554,In_663);
nor U2552 (N_2552,In_1033,In_1221);
nand U2553 (N_2553,In_175,In_983);
nand U2554 (N_2554,In_64,In_1888);
and U2555 (N_2555,In_1815,In_272);
nand U2556 (N_2556,In_225,In_339);
nor U2557 (N_2557,In_205,In_257);
nor U2558 (N_2558,In_1645,In_1653);
or U2559 (N_2559,In_120,In_1299);
or U2560 (N_2560,In_1594,In_1729);
nand U2561 (N_2561,In_311,In_447);
nand U2562 (N_2562,In_1173,In_296);
nand U2563 (N_2563,In_1417,In_313);
or U2564 (N_2564,In_419,In_1156);
nand U2565 (N_2565,In_1678,In_421);
nor U2566 (N_2566,In_1584,In_447);
nand U2567 (N_2567,In_1541,In_1484);
and U2568 (N_2568,In_1160,In_64);
nand U2569 (N_2569,In_1280,In_288);
xnor U2570 (N_2570,In_761,In_713);
and U2571 (N_2571,In_1452,In_1276);
xnor U2572 (N_2572,In_658,In_342);
nor U2573 (N_2573,In_1709,In_112);
and U2574 (N_2574,In_763,In_251);
xnor U2575 (N_2575,In_983,In_1386);
and U2576 (N_2576,In_968,In_17);
nor U2577 (N_2577,In_240,In_686);
nand U2578 (N_2578,In_1871,In_1245);
nor U2579 (N_2579,In_1109,In_1912);
and U2580 (N_2580,In_620,In_1614);
nand U2581 (N_2581,In_827,In_1849);
nor U2582 (N_2582,In_258,In_1896);
nor U2583 (N_2583,In_1857,In_1240);
or U2584 (N_2584,In_834,In_121);
or U2585 (N_2585,In_210,In_213);
nor U2586 (N_2586,In_142,In_618);
xnor U2587 (N_2587,In_915,In_425);
and U2588 (N_2588,In_679,In_365);
and U2589 (N_2589,In_902,In_1797);
nor U2590 (N_2590,In_1527,In_711);
xor U2591 (N_2591,In_1110,In_1860);
xnor U2592 (N_2592,In_1721,In_1684);
nand U2593 (N_2593,In_1075,In_1142);
nor U2594 (N_2594,In_1547,In_1666);
and U2595 (N_2595,In_1875,In_1755);
or U2596 (N_2596,In_503,In_267);
and U2597 (N_2597,In_1210,In_1045);
nand U2598 (N_2598,In_460,In_1198);
or U2599 (N_2599,In_999,In_117);
xor U2600 (N_2600,In_1779,In_1115);
nor U2601 (N_2601,In_1293,In_1161);
and U2602 (N_2602,In_1534,In_1111);
and U2603 (N_2603,In_112,In_556);
and U2604 (N_2604,In_1038,In_1076);
and U2605 (N_2605,In_253,In_797);
nor U2606 (N_2606,In_610,In_978);
or U2607 (N_2607,In_1257,In_1912);
and U2608 (N_2608,In_525,In_1140);
or U2609 (N_2609,In_1232,In_516);
or U2610 (N_2610,In_389,In_660);
nor U2611 (N_2611,In_296,In_458);
xor U2612 (N_2612,In_665,In_996);
or U2613 (N_2613,In_1365,In_1704);
and U2614 (N_2614,In_126,In_346);
nand U2615 (N_2615,In_624,In_1186);
nor U2616 (N_2616,In_12,In_1790);
or U2617 (N_2617,In_1228,In_1463);
or U2618 (N_2618,In_1853,In_1227);
and U2619 (N_2619,In_1993,In_637);
nand U2620 (N_2620,In_664,In_1122);
xnor U2621 (N_2621,In_580,In_928);
xor U2622 (N_2622,In_1829,In_1449);
and U2623 (N_2623,In_897,In_1127);
and U2624 (N_2624,In_458,In_1039);
and U2625 (N_2625,In_1053,In_750);
nand U2626 (N_2626,In_275,In_1581);
nor U2627 (N_2627,In_563,In_426);
and U2628 (N_2628,In_1080,In_179);
and U2629 (N_2629,In_941,In_1624);
nand U2630 (N_2630,In_1888,In_275);
or U2631 (N_2631,In_1683,In_1798);
or U2632 (N_2632,In_1469,In_424);
nor U2633 (N_2633,In_1667,In_1412);
or U2634 (N_2634,In_1801,In_297);
nand U2635 (N_2635,In_913,In_186);
and U2636 (N_2636,In_1724,In_1624);
and U2637 (N_2637,In_123,In_1367);
nor U2638 (N_2638,In_974,In_1891);
nand U2639 (N_2639,In_1577,In_801);
nor U2640 (N_2640,In_107,In_155);
xor U2641 (N_2641,In_1001,In_35);
or U2642 (N_2642,In_1599,In_668);
or U2643 (N_2643,In_458,In_741);
nand U2644 (N_2644,In_332,In_57);
nand U2645 (N_2645,In_1388,In_43);
xnor U2646 (N_2646,In_690,In_469);
nand U2647 (N_2647,In_648,In_1349);
nand U2648 (N_2648,In_752,In_1897);
and U2649 (N_2649,In_431,In_1370);
nand U2650 (N_2650,In_1766,In_1146);
or U2651 (N_2651,In_1204,In_1849);
xor U2652 (N_2652,In_284,In_120);
or U2653 (N_2653,In_1713,In_1948);
and U2654 (N_2654,In_1469,In_1910);
or U2655 (N_2655,In_1887,In_362);
or U2656 (N_2656,In_1461,In_1447);
or U2657 (N_2657,In_617,In_1917);
nor U2658 (N_2658,In_780,In_491);
nand U2659 (N_2659,In_606,In_1054);
xor U2660 (N_2660,In_565,In_1538);
xor U2661 (N_2661,In_1013,In_1342);
and U2662 (N_2662,In_1268,In_974);
nor U2663 (N_2663,In_1515,In_80);
nand U2664 (N_2664,In_1877,In_231);
nor U2665 (N_2665,In_805,In_737);
and U2666 (N_2666,In_1740,In_1703);
and U2667 (N_2667,In_1775,In_1961);
nand U2668 (N_2668,In_893,In_1117);
nor U2669 (N_2669,In_1070,In_569);
and U2670 (N_2670,In_1438,In_615);
xnor U2671 (N_2671,In_771,In_1772);
or U2672 (N_2672,In_681,In_1788);
and U2673 (N_2673,In_216,In_171);
or U2674 (N_2674,In_166,In_808);
nand U2675 (N_2675,In_1335,In_219);
xor U2676 (N_2676,In_417,In_1875);
xor U2677 (N_2677,In_1251,In_1138);
nor U2678 (N_2678,In_1530,In_1185);
or U2679 (N_2679,In_598,In_397);
and U2680 (N_2680,In_1845,In_892);
nand U2681 (N_2681,In_486,In_1712);
xor U2682 (N_2682,In_1217,In_1768);
nand U2683 (N_2683,In_1804,In_594);
and U2684 (N_2684,In_202,In_1769);
nor U2685 (N_2685,In_1216,In_1123);
nand U2686 (N_2686,In_1745,In_364);
or U2687 (N_2687,In_192,In_659);
nor U2688 (N_2688,In_1159,In_82);
nand U2689 (N_2689,In_1915,In_668);
or U2690 (N_2690,In_281,In_1871);
and U2691 (N_2691,In_1629,In_1766);
xor U2692 (N_2692,In_1546,In_387);
nand U2693 (N_2693,In_1924,In_8);
nand U2694 (N_2694,In_557,In_357);
nor U2695 (N_2695,In_1019,In_238);
or U2696 (N_2696,In_34,In_371);
and U2697 (N_2697,In_699,In_1477);
and U2698 (N_2698,In_1592,In_1127);
or U2699 (N_2699,In_1030,In_630);
or U2700 (N_2700,In_1382,In_895);
or U2701 (N_2701,In_516,In_484);
or U2702 (N_2702,In_847,In_1343);
nand U2703 (N_2703,In_1554,In_1636);
and U2704 (N_2704,In_1967,In_1138);
and U2705 (N_2705,In_555,In_1215);
nand U2706 (N_2706,In_1255,In_904);
nand U2707 (N_2707,In_1805,In_1991);
nor U2708 (N_2708,In_1747,In_1649);
xnor U2709 (N_2709,In_1380,In_261);
nand U2710 (N_2710,In_291,In_1759);
and U2711 (N_2711,In_1846,In_122);
or U2712 (N_2712,In_1242,In_378);
nor U2713 (N_2713,In_1962,In_1933);
nor U2714 (N_2714,In_655,In_710);
nor U2715 (N_2715,In_1468,In_1273);
nor U2716 (N_2716,In_302,In_1857);
nor U2717 (N_2717,In_622,In_932);
and U2718 (N_2718,In_420,In_1623);
or U2719 (N_2719,In_1486,In_714);
or U2720 (N_2720,In_1222,In_871);
nor U2721 (N_2721,In_890,In_1269);
or U2722 (N_2722,In_896,In_103);
or U2723 (N_2723,In_1499,In_1435);
or U2724 (N_2724,In_380,In_229);
nor U2725 (N_2725,In_865,In_1272);
nor U2726 (N_2726,In_1311,In_373);
nor U2727 (N_2727,In_145,In_239);
nor U2728 (N_2728,In_1977,In_1071);
or U2729 (N_2729,In_1322,In_1238);
nand U2730 (N_2730,In_581,In_201);
nand U2731 (N_2731,In_1462,In_1244);
nand U2732 (N_2732,In_1469,In_1727);
nand U2733 (N_2733,In_1829,In_1730);
nor U2734 (N_2734,In_1723,In_972);
and U2735 (N_2735,In_506,In_1164);
and U2736 (N_2736,In_375,In_668);
and U2737 (N_2737,In_1974,In_424);
nor U2738 (N_2738,In_1527,In_1295);
and U2739 (N_2739,In_1550,In_767);
nor U2740 (N_2740,In_1956,In_1530);
and U2741 (N_2741,In_209,In_1406);
xnor U2742 (N_2742,In_1090,In_1665);
or U2743 (N_2743,In_1395,In_692);
and U2744 (N_2744,In_677,In_112);
nor U2745 (N_2745,In_16,In_259);
nand U2746 (N_2746,In_1856,In_703);
or U2747 (N_2747,In_668,In_1118);
nor U2748 (N_2748,In_1114,In_25);
or U2749 (N_2749,In_1444,In_736);
nand U2750 (N_2750,In_970,In_932);
nor U2751 (N_2751,In_37,In_1814);
nand U2752 (N_2752,In_534,In_555);
xor U2753 (N_2753,In_1944,In_1164);
and U2754 (N_2754,In_487,In_1169);
xnor U2755 (N_2755,In_670,In_289);
or U2756 (N_2756,In_1614,In_1316);
or U2757 (N_2757,In_457,In_329);
xnor U2758 (N_2758,In_1899,In_1940);
and U2759 (N_2759,In_1699,In_924);
and U2760 (N_2760,In_1312,In_38);
or U2761 (N_2761,In_1070,In_1843);
nor U2762 (N_2762,In_447,In_1558);
nor U2763 (N_2763,In_510,In_463);
and U2764 (N_2764,In_1236,In_52);
nor U2765 (N_2765,In_933,In_1645);
nor U2766 (N_2766,In_0,In_345);
or U2767 (N_2767,In_1228,In_522);
nand U2768 (N_2768,In_1543,In_1625);
or U2769 (N_2769,In_1442,In_495);
nand U2770 (N_2770,In_1129,In_253);
and U2771 (N_2771,In_121,In_1286);
and U2772 (N_2772,In_1299,In_1209);
or U2773 (N_2773,In_28,In_1382);
xor U2774 (N_2774,In_270,In_161);
nand U2775 (N_2775,In_783,In_520);
nand U2776 (N_2776,In_1502,In_842);
and U2777 (N_2777,In_15,In_975);
nand U2778 (N_2778,In_972,In_1159);
nor U2779 (N_2779,In_705,In_1486);
nand U2780 (N_2780,In_957,In_176);
nor U2781 (N_2781,In_839,In_896);
and U2782 (N_2782,In_580,In_339);
nand U2783 (N_2783,In_1922,In_928);
nor U2784 (N_2784,In_759,In_819);
or U2785 (N_2785,In_1706,In_2);
nor U2786 (N_2786,In_1986,In_188);
and U2787 (N_2787,In_602,In_112);
nor U2788 (N_2788,In_953,In_1195);
and U2789 (N_2789,In_235,In_322);
nand U2790 (N_2790,In_1727,In_1475);
and U2791 (N_2791,In_489,In_1659);
nand U2792 (N_2792,In_125,In_914);
and U2793 (N_2793,In_1264,In_1618);
nand U2794 (N_2794,In_1324,In_1509);
nand U2795 (N_2795,In_209,In_1153);
or U2796 (N_2796,In_1915,In_1476);
or U2797 (N_2797,In_744,In_1693);
or U2798 (N_2798,In_96,In_1761);
and U2799 (N_2799,In_574,In_962);
or U2800 (N_2800,In_1510,In_637);
nor U2801 (N_2801,In_1384,In_1374);
nor U2802 (N_2802,In_1009,In_37);
nand U2803 (N_2803,In_907,In_1086);
and U2804 (N_2804,In_248,In_79);
and U2805 (N_2805,In_948,In_1421);
nand U2806 (N_2806,In_1256,In_1028);
or U2807 (N_2807,In_499,In_498);
nand U2808 (N_2808,In_442,In_1042);
and U2809 (N_2809,In_1344,In_590);
or U2810 (N_2810,In_1735,In_1740);
nor U2811 (N_2811,In_1507,In_949);
nor U2812 (N_2812,In_825,In_748);
nor U2813 (N_2813,In_1971,In_22);
and U2814 (N_2814,In_1821,In_1619);
and U2815 (N_2815,In_1683,In_1799);
nor U2816 (N_2816,In_198,In_1784);
xnor U2817 (N_2817,In_1647,In_374);
and U2818 (N_2818,In_816,In_433);
and U2819 (N_2819,In_84,In_1579);
or U2820 (N_2820,In_649,In_1094);
nor U2821 (N_2821,In_833,In_1120);
nor U2822 (N_2822,In_1928,In_1410);
nor U2823 (N_2823,In_1198,In_1752);
nand U2824 (N_2824,In_1479,In_1688);
and U2825 (N_2825,In_1678,In_852);
nand U2826 (N_2826,In_213,In_1326);
nor U2827 (N_2827,In_1651,In_133);
nor U2828 (N_2828,In_794,In_1152);
xnor U2829 (N_2829,In_733,In_1062);
nand U2830 (N_2830,In_1341,In_52);
nor U2831 (N_2831,In_1935,In_29);
xor U2832 (N_2832,In_1764,In_470);
nor U2833 (N_2833,In_340,In_1676);
nor U2834 (N_2834,In_1467,In_581);
nand U2835 (N_2835,In_1829,In_1949);
xnor U2836 (N_2836,In_1446,In_37);
xnor U2837 (N_2837,In_444,In_781);
or U2838 (N_2838,In_1235,In_118);
and U2839 (N_2839,In_1679,In_1369);
nor U2840 (N_2840,In_565,In_1478);
nor U2841 (N_2841,In_1314,In_125);
or U2842 (N_2842,In_558,In_1593);
and U2843 (N_2843,In_1657,In_845);
xor U2844 (N_2844,In_1412,In_1678);
nand U2845 (N_2845,In_935,In_1326);
and U2846 (N_2846,In_775,In_386);
nor U2847 (N_2847,In_418,In_770);
xor U2848 (N_2848,In_1405,In_1775);
or U2849 (N_2849,In_1748,In_419);
or U2850 (N_2850,In_36,In_8);
xnor U2851 (N_2851,In_1280,In_1028);
xnor U2852 (N_2852,In_1156,In_163);
and U2853 (N_2853,In_837,In_1612);
or U2854 (N_2854,In_824,In_1896);
nand U2855 (N_2855,In_386,In_1432);
nand U2856 (N_2856,In_29,In_1433);
nor U2857 (N_2857,In_1137,In_1419);
nor U2858 (N_2858,In_521,In_733);
nor U2859 (N_2859,In_319,In_767);
nand U2860 (N_2860,In_1240,In_1933);
and U2861 (N_2861,In_1225,In_5);
nor U2862 (N_2862,In_673,In_200);
and U2863 (N_2863,In_1,In_835);
nor U2864 (N_2864,In_1155,In_623);
xor U2865 (N_2865,In_157,In_604);
nand U2866 (N_2866,In_997,In_1501);
and U2867 (N_2867,In_1511,In_877);
and U2868 (N_2868,In_638,In_470);
nand U2869 (N_2869,In_1358,In_1450);
nand U2870 (N_2870,In_266,In_1408);
or U2871 (N_2871,In_280,In_1947);
nor U2872 (N_2872,In_1414,In_1043);
and U2873 (N_2873,In_302,In_1265);
xor U2874 (N_2874,In_1864,In_1332);
nor U2875 (N_2875,In_172,In_617);
and U2876 (N_2876,In_1075,In_81);
or U2877 (N_2877,In_5,In_1616);
and U2878 (N_2878,In_265,In_214);
or U2879 (N_2879,In_1531,In_1478);
nand U2880 (N_2880,In_1293,In_1642);
or U2881 (N_2881,In_352,In_597);
nor U2882 (N_2882,In_617,In_1810);
and U2883 (N_2883,In_1540,In_1811);
or U2884 (N_2884,In_1479,In_125);
xnor U2885 (N_2885,In_740,In_1854);
or U2886 (N_2886,In_956,In_1075);
nand U2887 (N_2887,In_1748,In_1232);
nor U2888 (N_2888,In_1314,In_50);
and U2889 (N_2889,In_1284,In_283);
or U2890 (N_2890,In_1006,In_1311);
or U2891 (N_2891,In_1106,In_1132);
nor U2892 (N_2892,In_1387,In_1666);
xor U2893 (N_2893,In_1328,In_98);
and U2894 (N_2894,In_1055,In_1781);
or U2895 (N_2895,In_131,In_1605);
nand U2896 (N_2896,In_1311,In_238);
nand U2897 (N_2897,In_1797,In_1641);
and U2898 (N_2898,In_491,In_962);
nand U2899 (N_2899,In_1405,In_1196);
or U2900 (N_2900,In_895,In_404);
nand U2901 (N_2901,In_1118,In_1195);
nand U2902 (N_2902,In_675,In_1104);
or U2903 (N_2903,In_514,In_1604);
or U2904 (N_2904,In_1557,In_1138);
nor U2905 (N_2905,In_1162,In_1822);
or U2906 (N_2906,In_1912,In_1158);
nand U2907 (N_2907,In_439,In_1301);
nand U2908 (N_2908,In_732,In_1983);
nand U2909 (N_2909,In_380,In_1971);
or U2910 (N_2910,In_277,In_489);
xnor U2911 (N_2911,In_123,In_831);
and U2912 (N_2912,In_15,In_1407);
or U2913 (N_2913,In_1847,In_1641);
nand U2914 (N_2914,In_1780,In_808);
nand U2915 (N_2915,In_251,In_932);
xor U2916 (N_2916,In_1586,In_1470);
or U2917 (N_2917,In_1648,In_1924);
nand U2918 (N_2918,In_963,In_45);
nand U2919 (N_2919,In_1576,In_1097);
and U2920 (N_2920,In_1127,In_752);
nor U2921 (N_2921,In_672,In_339);
and U2922 (N_2922,In_626,In_67);
or U2923 (N_2923,In_640,In_278);
nand U2924 (N_2924,In_1524,In_1931);
and U2925 (N_2925,In_1010,In_819);
or U2926 (N_2926,In_1904,In_1447);
nand U2927 (N_2927,In_53,In_306);
nor U2928 (N_2928,In_536,In_49);
or U2929 (N_2929,In_1163,In_1708);
nand U2930 (N_2930,In_1652,In_736);
nand U2931 (N_2931,In_1918,In_785);
nor U2932 (N_2932,In_143,In_1073);
nor U2933 (N_2933,In_1680,In_1375);
xor U2934 (N_2934,In_1048,In_1907);
nand U2935 (N_2935,In_528,In_1038);
or U2936 (N_2936,In_1566,In_343);
and U2937 (N_2937,In_35,In_1621);
or U2938 (N_2938,In_1607,In_1043);
xor U2939 (N_2939,In_402,In_1517);
or U2940 (N_2940,In_1194,In_670);
nand U2941 (N_2941,In_1767,In_442);
nand U2942 (N_2942,In_1630,In_15);
nand U2943 (N_2943,In_55,In_599);
nor U2944 (N_2944,In_234,In_953);
and U2945 (N_2945,In_666,In_567);
xor U2946 (N_2946,In_1388,In_500);
nor U2947 (N_2947,In_628,In_1280);
xor U2948 (N_2948,In_1672,In_1640);
nor U2949 (N_2949,In_1195,In_20);
nand U2950 (N_2950,In_407,In_1916);
nor U2951 (N_2951,In_695,In_820);
nand U2952 (N_2952,In_1540,In_536);
or U2953 (N_2953,In_164,In_72);
nor U2954 (N_2954,In_895,In_893);
nor U2955 (N_2955,In_961,In_881);
nand U2956 (N_2956,In_1586,In_1175);
or U2957 (N_2957,In_778,In_525);
nand U2958 (N_2958,In_828,In_1509);
and U2959 (N_2959,In_1823,In_1578);
nor U2960 (N_2960,In_930,In_929);
or U2961 (N_2961,In_1870,In_437);
nand U2962 (N_2962,In_1103,In_1404);
nand U2963 (N_2963,In_877,In_1014);
and U2964 (N_2964,In_836,In_285);
or U2965 (N_2965,In_1205,In_1662);
and U2966 (N_2966,In_1517,In_1125);
nand U2967 (N_2967,In_650,In_1956);
nor U2968 (N_2968,In_1434,In_1697);
nand U2969 (N_2969,In_196,In_979);
and U2970 (N_2970,In_1167,In_1499);
or U2971 (N_2971,In_1819,In_1858);
or U2972 (N_2972,In_1599,In_1492);
and U2973 (N_2973,In_873,In_1111);
and U2974 (N_2974,In_869,In_838);
nand U2975 (N_2975,In_901,In_1147);
and U2976 (N_2976,In_1377,In_1681);
or U2977 (N_2977,In_56,In_12);
nor U2978 (N_2978,In_191,In_786);
xor U2979 (N_2979,In_1200,In_112);
xnor U2980 (N_2980,In_702,In_86);
or U2981 (N_2981,In_982,In_469);
or U2982 (N_2982,In_680,In_442);
nor U2983 (N_2983,In_792,In_1079);
nor U2984 (N_2984,In_1061,In_1070);
and U2985 (N_2985,In_1311,In_641);
nand U2986 (N_2986,In_942,In_1176);
and U2987 (N_2987,In_109,In_792);
xnor U2988 (N_2988,In_653,In_1157);
nor U2989 (N_2989,In_400,In_1259);
xnor U2990 (N_2990,In_245,In_1965);
nor U2991 (N_2991,In_455,In_462);
or U2992 (N_2992,In_567,In_42);
nor U2993 (N_2993,In_111,In_1830);
nand U2994 (N_2994,In_252,In_1344);
or U2995 (N_2995,In_1715,In_915);
nand U2996 (N_2996,In_1151,In_503);
and U2997 (N_2997,In_1456,In_375);
nand U2998 (N_2998,In_24,In_896);
or U2999 (N_2999,In_858,In_1011);
nand U3000 (N_3000,In_813,In_884);
nor U3001 (N_3001,In_77,In_336);
nand U3002 (N_3002,In_850,In_1059);
xnor U3003 (N_3003,In_1479,In_201);
nor U3004 (N_3004,In_962,In_1821);
or U3005 (N_3005,In_1709,In_952);
or U3006 (N_3006,In_428,In_471);
xor U3007 (N_3007,In_1338,In_361);
or U3008 (N_3008,In_928,In_14);
and U3009 (N_3009,In_1181,In_1847);
and U3010 (N_3010,In_433,In_560);
and U3011 (N_3011,In_583,In_1658);
xor U3012 (N_3012,In_20,In_603);
or U3013 (N_3013,In_205,In_901);
and U3014 (N_3014,In_145,In_866);
or U3015 (N_3015,In_306,In_1880);
and U3016 (N_3016,In_1023,In_418);
nand U3017 (N_3017,In_427,In_1930);
or U3018 (N_3018,In_736,In_1511);
or U3019 (N_3019,In_514,In_376);
nor U3020 (N_3020,In_980,In_581);
nand U3021 (N_3021,In_355,In_852);
nand U3022 (N_3022,In_564,In_1556);
xnor U3023 (N_3023,In_1819,In_1795);
or U3024 (N_3024,In_1536,In_261);
nor U3025 (N_3025,In_1844,In_1134);
nor U3026 (N_3026,In_965,In_1336);
and U3027 (N_3027,In_578,In_302);
or U3028 (N_3028,In_1670,In_937);
or U3029 (N_3029,In_1532,In_1168);
or U3030 (N_3030,In_114,In_1592);
nand U3031 (N_3031,In_1273,In_805);
or U3032 (N_3032,In_403,In_300);
and U3033 (N_3033,In_843,In_1098);
and U3034 (N_3034,In_1004,In_1968);
nand U3035 (N_3035,In_381,In_1192);
nand U3036 (N_3036,In_230,In_1899);
nor U3037 (N_3037,In_31,In_758);
or U3038 (N_3038,In_1407,In_1002);
or U3039 (N_3039,In_1869,In_1903);
or U3040 (N_3040,In_958,In_568);
nor U3041 (N_3041,In_57,In_1676);
and U3042 (N_3042,In_1139,In_892);
or U3043 (N_3043,In_1530,In_327);
and U3044 (N_3044,In_1842,In_1390);
and U3045 (N_3045,In_782,In_1717);
nor U3046 (N_3046,In_1341,In_1533);
nor U3047 (N_3047,In_291,In_783);
or U3048 (N_3048,In_623,In_770);
and U3049 (N_3049,In_719,In_148);
or U3050 (N_3050,In_698,In_1644);
nand U3051 (N_3051,In_181,In_1666);
xor U3052 (N_3052,In_1241,In_844);
nand U3053 (N_3053,In_1156,In_1568);
nor U3054 (N_3054,In_930,In_134);
or U3055 (N_3055,In_471,In_936);
or U3056 (N_3056,In_184,In_169);
and U3057 (N_3057,In_1589,In_1543);
nand U3058 (N_3058,In_355,In_1984);
or U3059 (N_3059,In_490,In_1242);
nor U3060 (N_3060,In_1616,In_850);
or U3061 (N_3061,In_795,In_1031);
nand U3062 (N_3062,In_688,In_1984);
and U3063 (N_3063,In_175,In_767);
nor U3064 (N_3064,In_810,In_1933);
and U3065 (N_3065,In_1091,In_1615);
nor U3066 (N_3066,In_1480,In_1551);
nor U3067 (N_3067,In_1449,In_27);
or U3068 (N_3068,In_964,In_934);
and U3069 (N_3069,In_1441,In_177);
or U3070 (N_3070,In_1360,In_500);
nor U3071 (N_3071,In_1895,In_222);
or U3072 (N_3072,In_1539,In_777);
nor U3073 (N_3073,In_154,In_1273);
nor U3074 (N_3074,In_1697,In_836);
and U3075 (N_3075,In_1408,In_1142);
xnor U3076 (N_3076,In_160,In_1036);
and U3077 (N_3077,In_1062,In_1576);
nand U3078 (N_3078,In_1195,In_384);
xnor U3079 (N_3079,In_1685,In_1566);
or U3080 (N_3080,In_158,In_1413);
and U3081 (N_3081,In_1583,In_1984);
nand U3082 (N_3082,In_484,In_1983);
or U3083 (N_3083,In_456,In_746);
xnor U3084 (N_3084,In_406,In_120);
or U3085 (N_3085,In_826,In_1802);
or U3086 (N_3086,In_828,In_841);
nand U3087 (N_3087,In_1966,In_163);
or U3088 (N_3088,In_1376,In_703);
xor U3089 (N_3089,In_319,In_1042);
nand U3090 (N_3090,In_336,In_1884);
xor U3091 (N_3091,In_1149,In_432);
nor U3092 (N_3092,In_1032,In_1091);
or U3093 (N_3093,In_1179,In_591);
or U3094 (N_3094,In_1920,In_1795);
or U3095 (N_3095,In_462,In_1944);
nand U3096 (N_3096,In_1785,In_342);
xnor U3097 (N_3097,In_1739,In_265);
or U3098 (N_3098,In_385,In_724);
or U3099 (N_3099,In_1691,In_206);
nor U3100 (N_3100,In_1855,In_1432);
or U3101 (N_3101,In_1856,In_430);
xnor U3102 (N_3102,In_1856,In_1283);
xnor U3103 (N_3103,In_893,In_892);
and U3104 (N_3104,In_36,In_1486);
nand U3105 (N_3105,In_892,In_1066);
and U3106 (N_3106,In_330,In_1606);
nor U3107 (N_3107,In_131,In_552);
and U3108 (N_3108,In_1075,In_1481);
xnor U3109 (N_3109,In_467,In_521);
or U3110 (N_3110,In_1430,In_785);
nor U3111 (N_3111,In_1639,In_1593);
or U3112 (N_3112,In_803,In_842);
xor U3113 (N_3113,In_1611,In_424);
xnor U3114 (N_3114,In_1021,In_167);
nor U3115 (N_3115,In_477,In_1802);
nor U3116 (N_3116,In_895,In_43);
nand U3117 (N_3117,In_80,In_1724);
and U3118 (N_3118,In_466,In_355);
and U3119 (N_3119,In_1719,In_1242);
or U3120 (N_3120,In_1545,In_1046);
nand U3121 (N_3121,In_1171,In_1392);
or U3122 (N_3122,In_477,In_693);
nor U3123 (N_3123,In_1214,In_628);
nand U3124 (N_3124,In_509,In_316);
nand U3125 (N_3125,In_930,In_1469);
or U3126 (N_3126,In_1320,In_914);
and U3127 (N_3127,In_584,In_243);
and U3128 (N_3128,In_436,In_1477);
and U3129 (N_3129,In_326,In_1475);
xnor U3130 (N_3130,In_478,In_1372);
nand U3131 (N_3131,In_372,In_1736);
xnor U3132 (N_3132,In_561,In_489);
or U3133 (N_3133,In_314,In_1256);
or U3134 (N_3134,In_1800,In_127);
nor U3135 (N_3135,In_210,In_869);
and U3136 (N_3136,In_1795,In_1520);
or U3137 (N_3137,In_135,In_1031);
and U3138 (N_3138,In_1133,In_1549);
and U3139 (N_3139,In_337,In_1129);
nor U3140 (N_3140,In_1342,In_1167);
nand U3141 (N_3141,In_1071,In_1258);
nor U3142 (N_3142,In_1830,In_689);
nor U3143 (N_3143,In_370,In_1686);
xnor U3144 (N_3144,In_1393,In_1092);
nand U3145 (N_3145,In_202,In_1606);
nand U3146 (N_3146,In_610,In_484);
nand U3147 (N_3147,In_48,In_1977);
nor U3148 (N_3148,In_643,In_1535);
xor U3149 (N_3149,In_931,In_1348);
nor U3150 (N_3150,In_329,In_1713);
or U3151 (N_3151,In_1968,In_1862);
or U3152 (N_3152,In_1380,In_570);
nor U3153 (N_3153,In_1868,In_363);
or U3154 (N_3154,In_845,In_1413);
xnor U3155 (N_3155,In_733,In_1277);
nand U3156 (N_3156,In_1978,In_678);
xnor U3157 (N_3157,In_1678,In_285);
or U3158 (N_3158,In_1963,In_456);
nor U3159 (N_3159,In_534,In_407);
nand U3160 (N_3160,In_1043,In_722);
or U3161 (N_3161,In_757,In_334);
nand U3162 (N_3162,In_730,In_1252);
and U3163 (N_3163,In_683,In_71);
and U3164 (N_3164,In_1662,In_1809);
or U3165 (N_3165,In_974,In_1295);
nor U3166 (N_3166,In_1296,In_1197);
or U3167 (N_3167,In_534,In_926);
or U3168 (N_3168,In_155,In_1506);
or U3169 (N_3169,In_662,In_1446);
or U3170 (N_3170,In_469,In_188);
or U3171 (N_3171,In_1392,In_1055);
nor U3172 (N_3172,In_1738,In_1457);
nand U3173 (N_3173,In_1968,In_1291);
and U3174 (N_3174,In_1252,In_591);
or U3175 (N_3175,In_538,In_1584);
or U3176 (N_3176,In_608,In_1278);
or U3177 (N_3177,In_881,In_1598);
and U3178 (N_3178,In_1598,In_1086);
xor U3179 (N_3179,In_23,In_1150);
and U3180 (N_3180,In_613,In_1186);
xor U3181 (N_3181,In_415,In_1160);
or U3182 (N_3182,In_984,In_1121);
nor U3183 (N_3183,In_90,In_1219);
nor U3184 (N_3184,In_922,In_1306);
and U3185 (N_3185,In_76,In_1740);
xor U3186 (N_3186,In_76,In_142);
or U3187 (N_3187,In_894,In_1998);
and U3188 (N_3188,In_980,In_996);
nor U3189 (N_3189,In_499,In_1647);
nor U3190 (N_3190,In_1705,In_740);
nor U3191 (N_3191,In_1685,In_604);
nand U3192 (N_3192,In_1511,In_995);
nand U3193 (N_3193,In_1172,In_1343);
xnor U3194 (N_3194,In_400,In_1280);
and U3195 (N_3195,In_1737,In_346);
nand U3196 (N_3196,In_703,In_1964);
nand U3197 (N_3197,In_302,In_922);
and U3198 (N_3198,In_38,In_1182);
nand U3199 (N_3199,In_833,In_606);
or U3200 (N_3200,In_1993,In_1882);
or U3201 (N_3201,In_1133,In_1177);
nand U3202 (N_3202,In_538,In_579);
nand U3203 (N_3203,In_1865,In_121);
xor U3204 (N_3204,In_1350,In_410);
nand U3205 (N_3205,In_1452,In_329);
and U3206 (N_3206,In_346,In_551);
nor U3207 (N_3207,In_1193,In_986);
and U3208 (N_3208,In_1503,In_1567);
and U3209 (N_3209,In_257,In_1758);
nor U3210 (N_3210,In_357,In_149);
and U3211 (N_3211,In_1040,In_1740);
or U3212 (N_3212,In_1119,In_1456);
or U3213 (N_3213,In_828,In_152);
or U3214 (N_3214,In_1807,In_1561);
xor U3215 (N_3215,In_510,In_421);
nor U3216 (N_3216,In_208,In_1210);
and U3217 (N_3217,In_1033,In_1266);
and U3218 (N_3218,In_1044,In_1467);
nand U3219 (N_3219,In_1285,In_190);
nand U3220 (N_3220,In_1173,In_654);
nor U3221 (N_3221,In_1034,In_1032);
nor U3222 (N_3222,In_127,In_1703);
or U3223 (N_3223,In_175,In_40);
nand U3224 (N_3224,In_1145,In_663);
nand U3225 (N_3225,In_1706,In_199);
xnor U3226 (N_3226,In_253,In_1813);
nor U3227 (N_3227,In_1504,In_204);
nor U3228 (N_3228,In_366,In_1778);
nand U3229 (N_3229,In_1201,In_1700);
nand U3230 (N_3230,In_1827,In_1419);
nor U3231 (N_3231,In_1474,In_210);
and U3232 (N_3232,In_1408,In_1385);
or U3233 (N_3233,In_1038,In_1783);
and U3234 (N_3234,In_851,In_1837);
nor U3235 (N_3235,In_955,In_1907);
and U3236 (N_3236,In_1655,In_1721);
and U3237 (N_3237,In_1084,In_1115);
nand U3238 (N_3238,In_1840,In_1183);
or U3239 (N_3239,In_1598,In_590);
and U3240 (N_3240,In_1069,In_1976);
or U3241 (N_3241,In_855,In_1025);
nand U3242 (N_3242,In_1326,In_1467);
nor U3243 (N_3243,In_1126,In_316);
nor U3244 (N_3244,In_190,In_820);
nand U3245 (N_3245,In_1679,In_1117);
nand U3246 (N_3246,In_751,In_662);
or U3247 (N_3247,In_273,In_932);
nand U3248 (N_3248,In_1980,In_511);
nor U3249 (N_3249,In_1264,In_449);
nand U3250 (N_3250,In_1981,In_282);
and U3251 (N_3251,In_1754,In_982);
nor U3252 (N_3252,In_1136,In_456);
nor U3253 (N_3253,In_1294,In_939);
nor U3254 (N_3254,In_1165,In_1076);
nor U3255 (N_3255,In_520,In_1973);
or U3256 (N_3256,In_197,In_1991);
nor U3257 (N_3257,In_1732,In_1833);
or U3258 (N_3258,In_296,In_1857);
and U3259 (N_3259,In_1570,In_1783);
or U3260 (N_3260,In_864,In_945);
and U3261 (N_3261,In_1152,In_452);
and U3262 (N_3262,In_349,In_747);
or U3263 (N_3263,In_1774,In_1771);
and U3264 (N_3264,In_236,In_230);
nand U3265 (N_3265,In_579,In_937);
or U3266 (N_3266,In_953,In_543);
and U3267 (N_3267,In_1496,In_302);
or U3268 (N_3268,In_1655,In_882);
nand U3269 (N_3269,In_623,In_1437);
nand U3270 (N_3270,In_1916,In_660);
nand U3271 (N_3271,In_1928,In_44);
nor U3272 (N_3272,In_997,In_527);
nand U3273 (N_3273,In_1390,In_175);
and U3274 (N_3274,In_861,In_1421);
nor U3275 (N_3275,In_204,In_637);
or U3276 (N_3276,In_340,In_1877);
or U3277 (N_3277,In_392,In_1213);
nand U3278 (N_3278,In_991,In_634);
nand U3279 (N_3279,In_1402,In_1514);
or U3280 (N_3280,In_1439,In_356);
nor U3281 (N_3281,In_1748,In_1861);
or U3282 (N_3282,In_1135,In_1846);
nand U3283 (N_3283,In_124,In_1479);
or U3284 (N_3284,In_808,In_1650);
nand U3285 (N_3285,In_1928,In_1338);
nand U3286 (N_3286,In_934,In_57);
or U3287 (N_3287,In_863,In_1672);
nor U3288 (N_3288,In_424,In_1299);
xor U3289 (N_3289,In_795,In_324);
nor U3290 (N_3290,In_889,In_1918);
nand U3291 (N_3291,In_34,In_1961);
nor U3292 (N_3292,In_1530,In_977);
nor U3293 (N_3293,In_33,In_514);
or U3294 (N_3294,In_1873,In_1542);
nor U3295 (N_3295,In_1175,In_420);
nand U3296 (N_3296,In_263,In_222);
and U3297 (N_3297,In_1282,In_1008);
and U3298 (N_3298,In_1262,In_1996);
nor U3299 (N_3299,In_1394,In_1077);
nand U3300 (N_3300,In_1837,In_1873);
nand U3301 (N_3301,In_879,In_673);
or U3302 (N_3302,In_106,In_788);
and U3303 (N_3303,In_1830,In_3);
nor U3304 (N_3304,In_141,In_1187);
nor U3305 (N_3305,In_1710,In_1512);
nand U3306 (N_3306,In_654,In_113);
nor U3307 (N_3307,In_1107,In_1223);
nand U3308 (N_3308,In_133,In_3);
nand U3309 (N_3309,In_662,In_1388);
nor U3310 (N_3310,In_1327,In_646);
nor U3311 (N_3311,In_48,In_1559);
or U3312 (N_3312,In_1906,In_889);
nor U3313 (N_3313,In_1331,In_1210);
and U3314 (N_3314,In_1420,In_143);
nor U3315 (N_3315,In_85,In_415);
or U3316 (N_3316,In_1824,In_1903);
nand U3317 (N_3317,In_1193,In_1584);
and U3318 (N_3318,In_1359,In_1577);
nand U3319 (N_3319,In_295,In_292);
or U3320 (N_3320,In_602,In_1237);
or U3321 (N_3321,In_1307,In_216);
xnor U3322 (N_3322,In_130,In_798);
nor U3323 (N_3323,In_575,In_1270);
or U3324 (N_3324,In_1103,In_153);
and U3325 (N_3325,In_1729,In_339);
xnor U3326 (N_3326,In_1658,In_993);
or U3327 (N_3327,In_315,In_1764);
and U3328 (N_3328,In_276,In_1778);
and U3329 (N_3329,In_1981,In_1113);
nor U3330 (N_3330,In_951,In_1151);
nand U3331 (N_3331,In_1262,In_468);
nor U3332 (N_3332,In_956,In_776);
and U3333 (N_3333,In_494,In_138);
and U3334 (N_3334,In_1998,In_1589);
or U3335 (N_3335,In_1762,In_176);
and U3336 (N_3336,In_305,In_1660);
or U3337 (N_3337,In_369,In_402);
nand U3338 (N_3338,In_1019,In_1666);
nor U3339 (N_3339,In_70,In_1003);
nand U3340 (N_3340,In_1183,In_718);
and U3341 (N_3341,In_282,In_115);
or U3342 (N_3342,In_1740,In_1872);
nand U3343 (N_3343,In_183,In_979);
nor U3344 (N_3344,In_558,In_1481);
xor U3345 (N_3345,In_1053,In_1902);
and U3346 (N_3346,In_93,In_786);
nand U3347 (N_3347,In_923,In_300);
nand U3348 (N_3348,In_421,In_998);
nand U3349 (N_3349,In_292,In_520);
or U3350 (N_3350,In_784,In_340);
and U3351 (N_3351,In_332,In_427);
nor U3352 (N_3352,In_1843,In_799);
and U3353 (N_3353,In_1212,In_853);
and U3354 (N_3354,In_1128,In_608);
nor U3355 (N_3355,In_13,In_1530);
or U3356 (N_3356,In_597,In_562);
nor U3357 (N_3357,In_1477,In_1478);
nor U3358 (N_3358,In_778,In_368);
nor U3359 (N_3359,In_593,In_1940);
nor U3360 (N_3360,In_704,In_384);
or U3361 (N_3361,In_1291,In_1672);
nand U3362 (N_3362,In_969,In_1659);
or U3363 (N_3363,In_371,In_1248);
nand U3364 (N_3364,In_1614,In_1817);
or U3365 (N_3365,In_382,In_1009);
nor U3366 (N_3366,In_1780,In_1379);
xor U3367 (N_3367,In_431,In_1019);
and U3368 (N_3368,In_263,In_6);
nor U3369 (N_3369,In_333,In_224);
nor U3370 (N_3370,In_706,In_1950);
nand U3371 (N_3371,In_559,In_1558);
or U3372 (N_3372,In_1462,In_374);
nand U3373 (N_3373,In_933,In_1383);
and U3374 (N_3374,In_457,In_524);
nand U3375 (N_3375,In_995,In_1994);
and U3376 (N_3376,In_626,In_908);
and U3377 (N_3377,In_1637,In_218);
nor U3378 (N_3378,In_1971,In_1762);
nand U3379 (N_3379,In_661,In_1823);
nand U3380 (N_3380,In_1589,In_1064);
and U3381 (N_3381,In_1747,In_923);
nor U3382 (N_3382,In_233,In_1019);
xnor U3383 (N_3383,In_758,In_1457);
nand U3384 (N_3384,In_1287,In_727);
or U3385 (N_3385,In_360,In_764);
xnor U3386 (N_3386,In_1425,In_383);
nor U3387 (N_3387,In_1875,In_50);
nor U3388 (N_3388,In_1628,In_1750);
and U3389 (N_3389,In_449,In_140);
or U3390 (N_3390,In_1655,In_1824);
and U3391 (N_3391,In_1984,In_1652);
and U3392 (N_3392,In_1614,In_601);
and U3393 (N_3393,In_1292,In_65);
nand U3394 (N_3394,In_1326,In_1484);
nor U3395 (N_3395,In_11,In_1533);
nand U3396 (N_3396,In_1915,In_348);
xnor U3397 (N_3397,In_1990,In_1204);
and U3398 (N_3398,In_1603,In_1100);
and U3399 (N_3399,In_1791,In_806);
and U3400 (N_3400,In_1527,In_582);
and U3401 (N_3401,In_1005,In_484);
and U3402 (N_3402,In_1550,In_138);
nand U3403 (N_3403,In_260,In_992);
nor U3404 (N_3404,In_174,In_1799);
nand U3405 (N_3405,In_652,In_326);
and U3406 (N_3406,In_328,In_538);
nand U3407 (N_3407,In_594,In_1932);
and U3408 (N_3408,In_1241,In_913);
nand U3409 (N_3409,In_537,In_627);
nor U3410 (N_3410,In_1510,In_762);
and U3411 (N_3411,In_923,In_565);
nand U3412 (N_3412,In_534,In_15);
or U3413 (N_3413,In_1176,In_902);
and U3414 (N_3414,In_1770,In_986);
nor U3415 (N_3415,In_1643,In_377);
nor U3416 (N_3416,In_629,In_447);
or U3417 (N_3417,In_1883,In_528);
or U3418 (N_3418,In_259,In_1351);
and U3419 (N_3419,In_1969,In_776);
and U3420 (N_3420,In_201,In_1421);
nand U3421 (N_3421,In_430,In_879);
or U3422 (N_3422,In_1855,In_1040);
nand U3423 (N_3423,In_696,In_198);
and U3424 (N_3424,In_1997,In_1874);
xor U3425 (N_3425,In_529,In_991);
nand U3426 (N_3426,In_326,In_118);
nand U3427 (N_3427,In_148,In_968);
or U3428 (N_3428,In_1420,In_1914);
and U3429 (N_3429,In_750,In_1650);
nand U3430 (N_3430,In_1657,In_878);
nor U3431 (N_3431,In_1395,In_1807);
or U3432 (N_3432,In_795,In_379);
or U3433 (N_3433,In_1676,In_1292);
nand U3434 (N_3434,In_21,In_931);
and U3435 (N_3435,In_160,In_523);
nand U3436 (N_3436,In_1542,In_318);
nand U3437 (N_3437,In_1965,In_305);
and U3438 (N_3438,In_1510,In_1018);
nand U3439 (N_3439,In_208,In_1240);
and U3440 (N_3440,In_1404,In_263);
nor U3441 (N_3441,In_1625,In_1703);
nand U3442 (N_3442,In_713,In_569);
nand U3443 (N_3443,In_213,In_1068);
and U3444 (N_3444,In_1921,In_1015);
nand U3445 (N_3445,In_1949,In_719);
and U3446 (N_3446,In_1072,In_1803);
or U3447 (N_3447,In_635,In_1744);
and U3448 (N_3448,In_52,In_767);
or U3449 (N_3449,In_1744,In_1108);
or U3450 (N_3450,In_682,In_1771);
nand U3451 (N_3451,In_593,In_365);
nand U3452 (N_3452,In_1412,In_1885);
xor U3453 (N_3453,In_951,In_1688);
nand U3454 (N_3454,In_1356,In_1888);
and U3455 (N_3455,In_257,In_1727);
nand U3456 (N_3456,In_1247,In_621);
nand U3457 (N_3457,In_1670,In_1530);
nand U3458 (N_3458,In_1584,In_471);
or U3459 (N_3459,In_100,In_1100);
nand U3460 (N_3460,In_798,In_693);
nor U3461 (N_3461,In_1238,In_1920);
nor U3462 (N_3462,In_554,In_19);
nor U3463 (N_3463,In_553,In_1965);
and U3464 (N_3464,In_1788,In_74);
nand U3465 (N_3465,In_918,In_544);
nor U3466 (N_3466,In_322,In_1632);
nand U3467 (N_3467,In_1261,In_1629);
and U3468 (N_3468,In_775,In_785);
nor U3469 (N_3469,In_1852,In_1097);
or U3470 (N_3470,In_1033,In_1421);
or U3471 (N_3471,In_1368,In_240);
or U3472 (N_3472,In_1472,In_532);
nand U3473 (N_3473,In_1768,In_1743);
nor U3474 (N_3474,In_853,In_1125);
and U3475 (N_3475,In_1571,In_1195);
or U3476 (N_3476,In_985,In_1791);
nand U3477 (N_3477,In_683,In_838);
nor U3478 (N_3478,In_1336,In_389);
and U3479 (N_3479,In_250,In_1406);
nand U3480 (N_3480,In_1296,In_1069);
or U3481 (N_3481,In_1948,In_364);
nor U3482 (N_3482,In_1440,In_824);
nor U3483 (N_3483,In_1132,In_1740);
or U3484 (N_3484,In_1528,In_395);
and U3485 (N_3485,In_431,In_1297);
nor U3486 (N_3486,In_1021,In_1986);
and U3487 (N_3487,In_1664,In_186);
nand U3488 (N_3488,In_1533,In_900);
nand U3489 (N_3489,In_83,In_174);
nand U3490 (N_3490,In_1217,In_304);
nand U3491 (N_3491,In_1844,In_1225);
nor U3492 (N_3492,In_442,In_243);
nor U3493 (N_3493,In_1700,In_1113);
and U3494 (N_3494,In_1153,In_1313);
nor U3495 (N_3495,In_574,In_1396);
nand U3496 (N_3496,In_554,In_444);
and U3497 (N_3497,In_1424,In_1104);
and U3498 (N_3498,In_201,In_1084);
and U3499 (N_3499,In_254,In_944);
or U3500 (N_3500,In_845,In_1667);
nand U3501 (N_3501,In_944,In_910);
and U3502 (N_3502,In_670,In_721);
and U3503 (N_3503,In_93,In_618);
nor U3504 (N_3504,In_1991,In_1924);
nor U3505 (N_3505,In_1116,In_172);
nor U3506 (N_3506,In_1362,In_610);
nor U3507 (N_3507,In_682,In_1908);
or U3508 (N_3508,In_1351,In_1090);
nor U3509 (N_3509,In_287,In_967);
or U3510 (N_3510,In_1440,In_856);
nor U3511 (N_3511,In_1292,In_377);
nor U3512 (N_3512,In_1369,In_85);
or U3513 (N_3513,In_1256,In_1110);
nor U3514 (N_3514,In_431,In_1294);
nor U3515 (N_3515,In_1944,In_1638);
nor U3516 (N_3516,In_691,In_1382);
and U3517 (N_3517,In_21,In_1721);
or U3518 (N_3518,In_1123,In_648);
or U3519 (N_3519,In_357,In_1611);
nand U3520 (N_3520,In_1705,In_1597);
nand U3521 (N_3521,In_1416,In_466);
nor U3522 (N_3522,In_1865,In_1568);
nand U3523 (N_3523,In_472,In_1590);
or U3524 (N_3524,In_1983,In_85);
nor U3525 (N_3525,In_1051,In_1251);
or U3526 (N_3526,In_1605,In_989);
or U3527 (N_3527,In_754,In_720);
nand U3528 (N_3528,In_1247,In_1813);
or U3529 (N_3529,In_1423,In_458);
and U3530 (N_3530,In_1909,In_1642);
or U3531 (N_3531,In_1841,In_99);
or U3532 (N_3532,In_557,In_1884);
nand U3533 (N_3533,In_1662,In_1369);
or U3534 (N_3534,In_974,In_1931);
xnor U3535 (N_3535,In_1496,In_674);
and U3536 (N_3536,In_1677,In_1958);
or U3537 (N_3537,In_743,In_1438);
or U3538 (N_3538,In_141,In_980);
nand U3539 (N_3539,In_531,In_792);
or U3540 (N_3540,In_293,In_967);
and U3541 (N_3541,In_1625,In_763);
or U3542 (N_3542,In_1252,In_452);
or U3543 (N_3543,In_420,In_385);
nor U3544 (N_3544,In_971,In_1012);
nand U3545 (N_3545,In_5,In_356);
and U3546 (N_3546,In_808,In_112);
nor U3547 (N_3547,In_655,In_17);
nand U3548 (N_3548,In_1102,In_1306);
or U3549 (N_3549,In_1856,In_1989);
and U3550 (N_3550,In_292,In_709);
and U3551 (N_3551,In_905,In_1101);
and U3552 (N_3552,In_242,In_1078);
nor U3553 (N_3553,In_840,In_144);
and U3554 (N_3554,In_963,In_1342);
and U3555 (N_3555,In_145,In_63);
and U3556 (N_3556,In_976,In_11);
or U3557 (N_3557,In_960,In_1714);
or U3558 (N_3558,In_1378,In_109);
or U3559 (N_3559,In_1740,In_1477);
or U3560 (N_3560,In_129,In_1895);
or U3561 (N_3561,In_1245,In_1667);
and U3562 (N_3562,In_802,In_404);
nor U3563 (N_3563,In_193,In_1662);
xnor U3564 (N_3564,In_154,In_1028);
and U3565 (N_3565,In_1551,In_963);
or U3566 (N_3566,In_1521,In_1671);
and U3567 (N_3567,In_1074,In_876);
nor U3568 (N_3568,In_154,In_1258);
or U3569 (N_3569,In_570,In_1406);
or U3570 (N_3570,In_1768,In_766);
and U3571 (N_3571,In_1710,In_56);
xor U3572 (N_3572,In_493,In_1919);
nand U3573 (N_3573,In_1444,In_405);
and U3574 (N_3574,In_184,In_1514);
or U3575 (N_3575,In_227,In_35);
nor U3576 (N_3576,In_1876,In_1219);
nand U3577 (N_3577,In_1833,In_713);
nand U3578 (N_3578,In_823,In_1428);
nand U3579 (N_3579,In_1572,In_896);
or U3580 (N_3580,In_1558,In_470);
and U3581 (N_3581,In_1037,In_637);
and U3582 (N_3582,In_1275,In_899);
and U3583 (N_3583,In_1752,In_1598);
or U3584 (N_3584,In_468,In_143);
nor U3585 (N_3585,In_1854,In_885);
nand U3586 (N_3586,In_323,In_786);
or U3587 (N_3587,In_1001,In_287);
nand U3588 (N_3588,In_1127,In_1811);
nor U3589 (N_3589,In_1335,In_729);
or U3590 (N_3590,In_1755,In_1930);
or U3591 (N_3591,In_1371,In_1742);
nor U3592 (N_3592,In_798,In_1671);
nor U3593 (N_3593,In_1060,In_1474);
nand U3594 (N_3594,In_1595,In_1632);
nand U3595 (N_3595,In_1889,In_1238);
or U3596 (N_3596,In_1346,In_1041);
or U3597 (N_3597,In_1390,In_170);
nand U3598 (N_3598,In_1354,In_520);
nor U3599 (N_3599,In_1946,In_1097);
or U3600 (N_3600,In_242,In_1877);
and U3601 (N_3601,In_671,In_1826);
nand U3602 (N_3602,In_436,In_1083);
nor U3603 (N_3603,In_1273,In_1401);
or U3604 (N_3604,In_491,In_56);
and U3605 (N_3605,In_1368,In_1888);
nand U3606 (N_3606,In_1609,In_478);
and U3607 (N_3607,In_1614,In_1653);
or U3608 (N_3608,In_359,In_502);
nor U3609 (N_3609,In_1061,In_1167);
and U3610 (N_3610,In_277,In_1052);
and U3611 (N_3611,In_482,In_1427);
nor U3612 (N_3612,In_138,In_957);
xor U3613 (N_3613,In_318,In_270);
and U3614 (N_3614,In_155,In_1435);
and U3615 (N_3615,In_1554,In_1577);
and U3616 (N_3616,In_909,In_505);
nor U3617 (N_3617,In_1274,In_563);
or U3618 (N_3618,In_1121,In_585);
nand U3619 (N_3619,In_481,In_1530);
nor U3620 (N_3620,In_633,In_663);
and U3621 (N_3621,In_334,In_1334);
or U3622 (N_3622,In_1361,In_1344);
xnor U3623 (N_3623,In_1368,In_1474);
or U3624 (N_3624,In_1291,In_143);
and U3625 (N_3625,In_976,In_629);
and U3626 (N_3626,In_1213,In_2);
nand U3627 (N_3627,In_1999,In_769);
nand U3628 (N_3628,In_1290,In_1327);
and U3629 (N_3629,In_390,In_1718);
or U3630 (N_3630,In_902,In_1824);
nor U3631 (N_3631,In_1368,In_1745);
nor U3632 (N_3632,In_1225,In_604);
or U3633 (N_3633,In_1084,In_816);
or U3634 (N_3634,In_353,In_1437);
or U3635 (N_3635,In_1808,In_276);
nand U3636 (N_3636,In_134,In_865);
and U3637 (N_3637,In_932,In_998);
or U3638 (N_3638,In_499,In_878);
nand U3639 (N_3639,In_1639,In_480);
or U3640 (N_3640,In_479,In_986);
nor U3641 (N_3641,In_1389,In_1640);
and U3642 (N_3642,In_191,In_1410);
or U3643 (N_3643,In_1168,In_1573);
and U3644 (N_3644,In_979,In_524);
and U3645 (N_3645,In_1771,In_1146);
or U3646 (N_3646,In_1450,In_940);
nand U3647 (N_3647,In_627,In_1703);
nand U3648 (N_3648,In_365,In_1473);
and U3649 (N_3649,In_621,In_1074);
nand U3650 (N_3650,In_919,In_952);
and U3651 (N_3651,In_475,In_474);
nor U3652 (N_3652,In_824,In_472);
and U3653 (N_3653,In_1145,In_527);
and U3654 (N_3654,In_760,In_268);
or U3655 (N_3655,In_1470,In_1234);
nor U3656 (N_3656,In_819,In_1837);
or U3657 (N_3657,In_1514,In_646);
nor U3658 (N_3658,In_1283,In_210);
nand U3659 (N_3659,In_1626,In_395);
and U3660 (N_3660,In_1562,In_1685);
nand U3661 (N_3661,In_485,In_1414);
nand U3662 (N_3662,In_9,In_902);
nand U3663 (N_3663,In_1844,In_1493);
nand U3664 (N_3664,In_518,In_51);
nand U3665 (N_3665,In_416,In_100);
nand U3666 (N_3666,In_1711,In_1497);
nand U3667 (N_3667,In_179,In_340);
or U3668 (N_3668,In_1494,In_192);
and U3669 (N_3669,In_801,In_328);
nor U3670 (N_3670,In_1744,In_816);
nand U3671 (N_3671,In_882,In_459);
xnor U3672 (N_3672,In_1758,In_1624);
nor U3673 (N_3673,In_171,In_868);
and U3674 (N_3674,In_912,In_508);
nand U3675 (N_3675,In_155,In_1804);
and U3676 (N_3676,In_254,In_666);
nor U3677 (N_3677,In_35,In_336);
and U3678 (N_3678,In_323,In_1831);
nand U3679 (N_3679,In_567,In_594);
nand U3680 (N_3680,In_150,In_1463);
nor U3681 (N_3681,In_1628,In_1704);
nand U3682 (N_3682,In_491,In_870);
nand U3683 (N_3683,In_793,In_26);
nor U3684 (N_3684,In_867,In_395);
nand U3685 (N_3685,In_1486,In_1212);
and U3686 (N_3686,In_1179,In_1314);
or U3687 (N_3687,In_180,In_406);
or U3688 (N_3688,In_1788,In_546);
nand U3689 (N_3689,In_852,In_474);
and U3690 (N_3690,In_633,In_1);
nand U3691 (N_3691,In_1161,In_1033);
and U3692 (N_3692,In_1652,In_746);
nor U3693 (N_3693,In_153,In_445);
nor U3694 (N_3694,In_308,In_1315);
or U3695 (N_3695,In_617,In_1166);
nand U3696 (N_3696,In_277,In_1386);
nand U3697 (N_3697,In_1890,In_505);
and U3698 (N_3698,In_1894,In_75);
or U3699 (N_3699,In_844,In_549);
nor U3700 (N_3700,In_1431,In_708);
nand U3701 (N_3701,In_1469,In_1993);
nand U3702 (N_3702,In_1999,In_406);
or U3703 (N_3703,In_1996,In_332);
and U3704 (N_3704,In_1678,In_1821);
and U3705 (N_3705,In_1956,In_1624);
and U3706 (N_3706,In_706,In_593);
or U3707 (N_3707,In_1680,In_806);
xor U3708 (N_3708,In_627,In_336);
nand U3709 (N_3709,In_240,In_1695);
and U3710 (N_3710,In_56,In_512);
nand U3711 (N_3711,In_990,In_752);
xnor U3712 (N_3712,In_1719,In_816);
or U3713 (N_3713,In_1154,In_372);
nand U3714 (N_3714,In_14,In_1870);
xnor U3715 (N_3715,In_184,In_1155);
and U3716 (N_3716,In_149,In_878);
nand U3717 (N_3717,In_1469,In_741);
nor U3718 (N_3718,In_1165,In_1995);
and U3719 (N_3719,In_1316,In_532);
or U3720 (N_3720,In_403,In_1000);
nand U3721 (N_3721,In_1599,In_1438);
nor U3722 (N_3722,In_558,In_1269);
or U3723 (N_3723,In_543,In_711);
nand U3724 (N_3724,In_1347,In_708);
xnor U3725 (N_3725,In_1138,In_730);
nor U3726 (N_3726,In_934,In_1528);
nor U3727 (N_3727,In_978,In_637);
nand U3728 (N_3728,In_638,In_1291);
or U3729 (N_3729,In_987,In_1753);
nor U3730 (N_3730,In_366,In_842);
nor U3731 (N_3731,In_191,In_52);
nor U3732 (N_3732,In_342,In_642);
or U3733 (N_3733,In_396,In_922);
nand U3734 (N_3734,In_162,In_1250);
or U3735 (N_3735,In_932,In_1745);
or U3736 (N_3736,In_1237,In_633);
or U3737 (N_3737,In_545,In_1229);
nor U3738 (N_3738,In_505,In_1523);
nand U3739 (N_3739,In_1922,In_588);
or U3740 (N_3740,In_1383,In_484);
and U3741 (N_3741,In_537,In_1642);
or U3742 (N_3742,In_1595,In_1998);
and U3743 (N_3743,In_1458,In_1301);
and U3744 (N_3744,In_1388,In_679);
nand U3745 (N_3745,In_1237,In_1372);
nand U3746 (N_3746,In_614,In_160);
and U3747 (N_3747,In_1067,In_271);
nand U3748 (N_3748,In_712,In_301);
nor U3749 (N_3749,In_1441,In_1002);
nand U3750 (N_3750,In_1385,In_196);
nor U3751 (N_3751,In_1744,In_1834);
and U3752 (N_3752,In_1213,In_1648);
xnor U3753 (N_3753,In_1493,In_1857);
and U3754 (N_3754,In_1569,In_895);
xor U3755 (N_3755,In_419,In_412);
nor U3756 (N_3756,In_457,In_1628);
or U3757 (N_3757,In_1914,In_1545);
or U3758 (N_3758,In_443,In_1027);
or U3759 (N_3759,In_1300,In_796);
or U3760 (N_3760,In_1645,In_370);
and U3761 (N_3761,In_1507,In_842);
or U3762 (N_3762,In_693,In_576);
nand U3763 (N_3763,In_393,In_1710);
xor U3764 (N_3764,In_1315,In_711);
xor U3765 (N_3765,In_1649,In_1832);
nor U3766 (N_3766,In_1489,In_1235);
nor U3767 (N_3767,In_692,In_1602);
nand U3768 (N_3768,In_1997,In_72);
nor U3769 (N_3769,In_706,In_184);
nand U3770 (N_3770,In_701,In_1447);
or U3771 (N_3771,In_1890,In_1393);
nand U3772 (N_3772,In_1397,In_79);
nor U3773 (N_3773,In_1027,In_1106);
nor U3774 (N_3774,In_1171,In_813);
and U3775 (N_3775,In_1021,In_470);
nand U3776 (N_3776,In_1550,In_1196);
nand U3777 (N_3777,In_1800,In_856);
or U3778 (N_3778,In_846,In_149);
or U3779 (N_3779,In_675,In_1994);
and U3780 (N_3780,In_939,In_1547);
nand U3781 (N_3781,In_1531,In_1877);
nand U3782 (N_3782,In_615,In_1521);
nand U3783 (N_3783,In_1388,In_1617);
and U3784 (N_3784,In_262,In_1940);
and U3785 (N_3785,In_291,In_1432);
xnor U3786 (N_3786,In_216,In_1565);
and U3787 (N_3787,In_1057,In_114);
or U3788 (N_3788,In_1446,In_428);
or U3789 (N_3789,In_1556,In_89);
nor U3790 (N_3790,In_1694,In_1302);
nor U3791 (N_3791,In_216,In_646);
nor U3792 (N_3792,In_1250,In_1527);
and U3793 (N_3793,In_199,In_1907);
and U3794 (N_3794,In_997,In_1930);
xnor U3795 (N_3795,In_868,In_891);
or U3796 (N_3796,In_1095,In_760);
or U3797 (N_3797,In_60,In_131);
nand U3798 (N_3798,In_1632,In_945);
or U3799 (N_3799,In_1119,In_756);
and U3800 (N_3800,In_577,In_1604);
or U3801 (N_3801,In_1213,In_934);
nor U3802 (N_3802,In_172,In_403);
or U3803 (N_3803,In_1616,In_1889);
nor U3804 (N_3804,In_7,In_304);
or U3805 (N_3805,In_415,In_336);
or U3806 (N_3806,In_460,In_1521);
nor U3807 (N_3807,In_349,In_1648);
nor U3808 (N_3808,In_280,In_82);
and U3809 (N_3809,In_1925,In_673);
or U3810 (N_3810,In_739,In_204);
and U3811 (N_3811,In_59,In_1659);
or U3812 (N_3812,In_900,In_1004);
nor U3813 (N_3813,In_177,In_58);
nor U3814 (N_3814,In_1732,In_1425);
nor U3815 (N_3815,In_204,In_1357);
nor U3816 (N_3816,In_199,In_1712);
and U3817 (N_3817,In_1703,In_358);
nor U3818 (N_3818,In_1599,In_125);
or U3819 (N_3819,In_1970,In_1719);
nor U3820 (N_3820,In_93,In_1515);
and U3821 (N_3821,In_499,In_1342);
nand U3822 (N_3822,In_1509,In_1338);
nand U3823 (N_3823,In_1602,In_1046);
xor U3824 (N_3824,In_1691,In_287);
nand U3825 (N_3825,In_1845,In_1039);
nand U3826 (N_3826,In_1422,In_1556);
nor U3827 (N_3827,In_35,In_797);
nand U3828 (N_3828,In_678,In_1703);
nor U3829 (N_3829,In_1381,In_1299);
or U3830 (N_3830,In_461,In_555);
xor U3831 (N_3831,In_879,In_938);
and U3832 (N_3832,In_782,In_386);
xnor U3833 (N_3833,In_264,In_421);
or U3834 (N_3834,In_225,In_314);
nand U3835 (N_3835,In_1403,In_429);
or U3836 (N_3836,In_727,In_18);
nand U3837 (N_3837,In_437,In_134);
nand U3838 (N_3838,In_1090,In_1765);
or U3839 (N_3839,In_1846,In_828);
or U3840 (N_3840,In_943,In_1208);
or U3841 (N_3841,In_1176,In_1013);
nor U3842 (N_3842,In_1812,In_409);
or U3843 (N_3843,In_920,In_102);
nor U3844 (N_3844,In_254,In_408);
and U3845 (N_3845,In_790,In_177);
nor U3846 (N_3846,In_767,In_1137);
and U3847 (N_3847,In_170,In_1087);
and U3848 (N_3848,In_869,In_1539);
and U3849 (N_3849,In_364,In_1148);
nor U3850 (N_3850,In_57,In_227);
or U3851 (N_3851,In_717,In_1783);
or U3852 (N_3852,In_813,In_7);
nand U3853 (N_3853,In_1100,In_307);
nand U3854 (N_3854,In_859,In_1339);
and U3855 (N_3855,In_1698,In_333);
nand U3856 (N_3856,In_180,In_111);
nor U3857 (N_3857,In_960,In_55);
nor U3858 (N_3858,In_172,In_223);
or U3859 (N_3859,In_844,In_1447);
xor U3860 (N_3860,In_271,In_143);
or U3861 (N_3861,In_1040,In_209);
or U3862 (N_3862,In_485,In_1568);
and U3863 (N_3863,In_14,In_794);
and U3864 (N_3864,In_1655,In_1549);
and U3865 (N_3865,In_1221,In_615);
nand U3866 (N_3866,In_1562,In_421);
nand U3867 (N_3867,In_541,In_165);
nor U3868 (N_3868,In_1120,In_1150);
or U3869 (N_3869,In_1896,In_1543);
and U3870 (N_3870,In_413,In_81);
nand U3871 (N_3871,In_791,In_741);
nor U3872 (N_3872,In_1301,In_1883);
and U3873 (N_3873,In_1789,In_167);
nor U3874 (N_3874,In_1255,In_1482);
nand U3875 (N_3875,In_1571,In_490);
nand U3876 (N_3876,In_364,In_1243);
or U3877 (N_3877,In_1627,In_198);
nor U3878 (N_3878,In_1797,In_1114);
and U3879 (N_3879,In_121,In_743);
xnor U3880 (N_3880,In_969,In_1013);
and U3881 (N_3881,In_248,In_262);
and U3882 (N_3882,In_1478,In_410);
or U3883 (N_3883,In_1278,In_373);
nand U3884 (N_3884,In_1179,In_728);
and U3885 (N_3885,In_1310,In_1014);
or U3886 (N_3886,In_919,In_1260);
nor U3887 (N_3887,In_33,In_89);
or U3888 (N_3888,In_278,In_304);
nand U3889 (N_3889,In_129,In_549);
or U3890 (N_3890,In_1918,In_647);
or U3891 (N_3891,In_1051,In_1400);
nand U3892 (N_3892,In_525,In_75);
xor U3893 (N_3893,In_382,In_1927);
nand U3894 (N_3894,In_1400,In_37);
nor U3895 (N_3895,In_705,In_991);
xnor U3896 (N_3896,In_1110,In_1961);
nor U3897 (N_3897,In_1688,In_1288);
nor U3898 (N_3898,In_474,In_823);
and U3899 (N_3899,In_374,In_673);
nor U3900 (N_3900,In_1652,In_54);
xnor U3901 (N_3901,In_1242,In_229);
xor U3902 (N_3902,In_1262,In_1421);
nor U3903 (N_3903,In_573,In_1571);
nand U3904 (N_3904,In_970,In_653);
and U3905 (N_3905,In_1899,In_251);
nand U3906 (N_3906,In_1227,In_442);
or U3907 (N_3907,In_630,In_1684);
nand U3908 (N_3908,In_1213,In_978);
xor U3909 (N_3909,In_1966,In_424);
nor U3910 (N_3910,In_834,In_190);
nor U3911 (N_3911,In_279,In_40);
nor U3912 (N_3912,In_855,In_637);
nor U3913 (N_3913,In_228,In_1919);
and U3914 (N_3914,In_984,In_117);
and U3915 (N_3915,In_569,In_1192);
and U3916 (N_3916,In_197,In_1622);
or U3917 (N_3917,In_802,In_815);
xnor U3918 (N_3918,In_740,In_910);
nand U3919 (N_3919,In_1567,In_1556);
and U3920 (N_3920,In_179,In_351);
xor U3921 (N_3921,In_1371,In_1702);
and U3922 (N_3922,In_1524,In_1272);
nand U3923 (N_3923,In_1308,In_785);
nor U3924 (N_3924,In_760,In_1315);
nand U3925 (N_3925,In_632,In_389);
nand U3926 (N_3926,In_1234,In_864);
and U3927 (N_3927,In_1085,In_1050);
nor U3928 (N_3928,In_1530,In_877);
nand U3929 (N_3929,In_303,In_972);
nor U3930 (N_3930,In_567,In_445);
or U3931 (N_3931,In_813,In_538);
nor U3932 (N_3932,In_38,In_237);
nor U3933 (N_3933,In_1332,In_1100);
or U3934 (N_3934,In_897,In_180);
nor U3935 (N_3935,In_1199,In_71);
and U3936 (N_3936,In_1932,In_400);
nand U3937 (N_3937,In_352,In_1728);
nand U3938 (N_3938,In_1544,In_208);
or U3939 (N_3939,In_1,In_1210);
nor U3940 (N_3940,In_1565,In_130);
nor U3941 (N_3941,In_319,In_421);
nand U3942 (N_3942,In_1944,In_1232);
or U3943 (N_3943,In_542,In_1755);
or U3944 (N_3944,In_463,In_809);
nand U3945 (N_3945,In_873,In_1777);
nand U3946 (N_3946,In_1338,In_167);
and U3947 (N_3947,In_1306,In_798);
xnor U3948 (N_3948,In_506,In_1863);
xor U3949 (N_3949,In_1571,In_598);
or U3950 (N_3950,In_1679,In_960);
xor U3951 (N_3951,In_1362,In_1482);
nor U3952 (N_3952,In_882,In_548);
nand U3953 (N_3953,In_4,In_842);
nand U3954 (N_3954,In_712,In_1235);
nor U3955 (N_3955,In_1076,In_833);
or U3956 (N_3956,In_555,In_438);
nor U3957 (N_3957,In_396,In_308);
xnor U3958 (N_3958,In_477,In_1799);
and U3959 (N_3959,In_1624,In_544);
nor U3960 (N_3960,In_1353,In_1594);
nand U3961 (N_3961,In_1289,In_707);
xor U3962 (N_3962,In_16,In_818);
nor U3963 (N_3963,In_1118,In_49);
nand U3964 (N_3964,In_1772,In_1819);
nand U3965 (N_3965,In_357,In_1963);
and U3966 (N_3966,In_126,In_1147);
or U3967 (N_3967,In_702,In_283);
or U3968 (N_3968,In_1696,In_464);
nand U3969 (N_3969,In_1828,In_1102);
and U3970 (N_3970,In_315,In_1178);
nand U3971 (N_3971,In_237,In_371);
xnor U3972 (N_3972,In_1231,In_1433);
or U3973 (N_3973,In_663,In_640);
and U3974 (N_3974,In_675,In_1006);
nor U3975 (N_3975,In_918,In_1184);
nand U3976 (N_3976,In_1085,In_1400);
nor U3977 (N_3977,In_53,In_788);
or U3978 (N_3978,In_1627,In_1000);
nand U3979 (N_3979,In_1150,In_1913);
nor U3980 (N_3980,In_1204,In_1645);
nand U3981 (N_3981,In_1874,In_1285);
or U3982 (N_3982,In_1685,In_966);
xor U3983 (N_3983,In_664,In_1328);
xnor U3984 (N_3984,In_310,In_1387);
and U3985 (N_3985,In_870,In_153);
and U3986 (N_3986,In_1869,In_186);
or U3987 (N_3987,In_141,In_1516);
or U3988 (N_3988,In_130,In_1839);
nor U3989 (N_3989,In_186,In_1672);
and U3990 (N_3990,In_825,In_1378);
nand U3991 (N_3991,In_1856,In_211);
nand U3992 (N_3992,In_210,In_275);
nand U3993 (N_3993,In_210,In_1075);
nand U3994 (N_3994,In_1797,In_491);
and U3995 (N_3995,In_888,In_96);
nand U3996 (N_3996,In_1635,In_656);
nor U3997 (N_3997,In_1217,In_1937);
nand U3998 (N_3998,In_1809,In_308);
and U3999 (N_3999,In_142,In_1262);
nand U4000 (N_4000,In_1102,In_1301);
or U4001 (N_4001,In_1082,In_4);
nor U4002 (N_4002,In_627,In_969);
nor U4003 (N_4003,In_114,In_1994);
nand U4004 (N_4004,In_1753,In_1354);
nor U4005 (N_4005,In_1782,In_252);
and U4006 (N_4006,In_1458,In_1637);
nand U4007 (N_4007,In_1476,In_1851);
xnor U4008 (N_4008,In_1300,In_780);
or U4009 (N_4009,In_1492,In_94);
or U4010 (N_4010,In_969,In_191);
and U4011 (N_4011,In_1374,In_1324);
or U4012 (N_4012,In_571,In_1339);
xor U4013 (N_4013,In_485,In_1762);
xnor U4014 (N_4014,In_309,In_1009);
nand U4015 (N_4015,In_1769,In_1140);
and U4016 (N_4016,In_1772,In_63);
and U4017 (N_4017,In_708,In_313);
nor U4018 (N_4018,In_1,In_1693);
nand U4019 (N_4019,In_286,In_71);
nand U4020 (N_4020,In_842,In_213);
or U4021 (N_4021,In_934,In_496);
nor U4022 (N_4022,In_891,In_1454);
and U4023 (N_4023,In_1978,In_1669);
or U4024 (N_4024,In_51,In_1326);
nor U4025 (N_4025,In_1063,In_166);
or U4026 (N_4026,In_440,In_727);
nor U4027 (N_4027,In_627,In_318);
or U4028 (N_4028,In_612,In_815);
nand U4029 (N_4029,In_1704,In_643);
nand U4030 (N_4030,In_1358,In_840);
nor U4031 (N_4031,In_765,In_143);
nor U4032 (N_4032,In_300,In_1365);
or U4033 (N_4033,In_284,In_1130);
nor U4034 (N_4034,In_914,In_466);
nor U4035 (N_4035,In_1913,In_633);
and U4036 (N_4036,In_1687,In_820);
xnor U4037 (N_4037,In_312,In_1501);
nor U4038 (N_4038,In_400,In_1323);
or U4039 (N_4039,In_729,In_1024);
nand U4040 (N_4040,In_467,In_1467);
or U4041 (N_4041,In_1932,In_907);
and U4042 (N_4042,In_394,In_986);
nor U4043 (N_4043,In_968,In_72);
or U4044 (N_4044,In_17,In_1830);
xor U4045 (N_4045,In_1327,In_1627);
nand U4046 (N_4046,In_50,In_1852);
or U4047 (N_4047,In_1390,In_533);
or U4048 (N_4048,In_233,In_516);
nand U4049 (N_4049,In_1202,In_1388);
and U4050 (N_4050,In_1191,In_1345);
nor U4051 (N_4051,In_415,In_1096);
xor U4052 (N_4052,In_1695,In_1558);
nand U4053 (N_4053,In_772,In_895);
nor U4054 (N_4054,In_1363,In_1548);
xnor U4055 (N_4055,In_1318,In_1289);
nor U4056 (N_4056,In_1348,In_543);
or U4057 (N_4057,In_55,In_1735);
or U4058 (N_4058,In_1546,In_1362);
xor U4059 (N_4059,In_1034,In_522);
nand U4060 (N_4060,In_441,In_112);
or U4061 (N_4061,In_942,In_1065);
or U4062 (N_4062,In_544,In_114);
or U4063 (N_4063,In_1283,In_1232);
nand U4064 (N_4064,In_195,In_994);
or U4065 (N_4065,In_1159,In_677);
or U4066 (N_4066,In_1808,In_552);
nand U4067 (N_4067,In_579,In_522);
xor U4068 (N_4068,In_683,In_1612);
nand U4069 (N_4069,In_1073,In_34);
nand U4070 (N_4070,In_1589,In_117);
nor U4071 (N_4071,In_478,In_1801);
nand U4072 (N_4072,In_409,In_1705);
and U4073 (N_4073,In_136,In_503);
and U4074 (N_4074,In_1996,In_733);
and U4075 (N_4075,In_1680,In_613);
nand U4076 (N_4076,In_1081,In_1532);
or U4077 (N_4077,In_247,In_1864);
and U4078 (N_4078,In_1634,In_1007);
or U4079 (N_4079,In_1820,In_1631);
or U4080 (N_4080,In_180,In_1580);
nand U4081 (N_4081,In_1514,In_651);
or U4082 (N_4082,In_952,In_831);
and U4083 (N_4083,In_1453,In_230);
nand U4084 (N_4084,In_643,In_1099);
nor U4085 (N_4085,In_952,In_489);
or U4086 (N_4086,In_1866,In_336);
nor U4087 (N_4087,In_1673,In_308);
and U4088 (N_4088,In_949,In_1165);
nand U4089 (N_4089,In_1415,In_619);
and U4090 (N_4090,In_905,In_1186);
and U4091 (N_4091,In_997,In_1879);
or U4092 (N_4092,In_1452,In_994);
and U4093 (N_4093,In_775,In_1809);
and U4094 (N_4094,In_856,In_1618);
nor U4095 (N_4095,In_471,In_150);
and U4096 (N_4096,In_57,In_1288);
or U4097 (N_4097,In_304,In_1503);
and U4098 (N_4098,In_1706,In_126);
nor U4099 (N_4099,In_547,In_70);
nor U4100 (N_4100,In_1435,In_171);
nor U4101 (N_4101,In_86,In_1909);
or U4102 (N_4102,In_316,In_1);
or U4103 (N_4103,In_1113,In_1413);
or U4104 (N_4104,In_1688,In_1034);
or U4105 (N_4105,In_1978,In_1391);
and U4106 (N_4106,In_187,In_1161);
and U4107 (N_4107,In_1261,In_1333);
xnor U4108 (N_4108,In_789,In_116);
and U4109 (N_4109,In_312,In_148);
or U4110 (N_4110,In_1888,In_19);
and U4111 (N_4111,In_264,In_778);
or U4112 (N_4112,In_660,In_1545);
xor U4113 (N_4113,In_620,In_1274);
nand U4114 (N_4114,In_1943,In_416);
nand U4115 (N_4115,In_280,In_462);
and U4116 (N_4116,In_1199,In_1608);
and U4117 (N_4117,In_977,In_1582);
and U4118 (N_4118,In_520,In_1943);
nor U4119 (N_4119,In_1890,In_442);
and U4120 (N_4120,In_1722,In_1515);
nor U4121 (N_4121,In_505,In_760);
and U4122 (N_4122,In_1543,In_898);
or U4123 (N_4123,In_1616,In_373);
nor U4124 (N_4124,In_758,In_593);
or U4125 (N_4125,In_790,In_924);
nand U4126 (N_4126,In_1346,In_174);
and U4127 (N_4127,In_147,In_942);
or U4128 (N_4128,In_1834,In_984);
nand U4129 (N_4129,In_811,In_1882);
nor U4130 (N_4130,In_1469,In_803);
and U4131 (N_4131,In_1669,In_486);
nand U4132 (N_4132,In_443,In_875);
nand U4133 (N_4133,In_1392,In_187);
nand U4134 (N_4134,In_440,In_36);
xor U4135 (N_4135,In_1507,In_1052);
or U4136 (N_4136,In_727,In_1808);
and U4137 (N_4137,In_1909,In_810);
nor U4138 (N_4138,In_439,In_1625);
or U4139 (N_4139,In_1428,In_924);
and U4140 (N_4140,In_1163,In_629);
or U4141 (N_4141,In_716,In_1290);
and U4142 (N_4142,In_722,In_724);
and U4143 (N_4143,In_677,In_1993);
or U4144 (N_4144,In_167,In_337);
nor U4145 (N_4145,In_541,In_1385);
or U4146 (N_4146,In_216,In_1286);
or U4147 (N_4147,In_1668,In_802);
nor U4148 (N_4148,In_446,In_46);
or U4149 (N_4149,In_1139,In_810);
or U4150 (N_4150,In_1584,In_1494);
nor U4151 (N_4151,In_1998,In_1551);
nand U4152 (N_4152,In_449,In_1624);
nand U4153 (N_4153,In_1381,In_1543);
nand U4154 (N_4154,In_1655,In_831);
nor U4155 (N_4155,In_1453,In_1329);
nor U4156 (N_4156,In_1878,In_1289);
or U4157 (N_4157,In_342,In_821);
and U4158 (N_4158,In_1948,In_1504);
and U4159 (N_4159,In_709,In_115);
nand U4160 (N_4160,In_696,In_937);
nor U4161 (N_4161,In_1427,In_313);
nor U4162 (N_4162,In_877,In_121);
and U4163 (N_4163,In_1916,In_1243);
nor U4164 (N_4164,In_977,In_1482);
nor U4165 (N_4165,In_346,In_239);
and U4166 (N_4166,In_741,In_238);
xnor U4167 (N_4167,In_1138,In_1449);
nand U4168 (N_4168,In_1622,In_206);
nor U4169 (N_4169,In_523,In_1008);
nand U4170 (N_4170,In_1786,In_1638);
nand U4171 (N_4171,In_1830,In_222);
nand U4172 (N_4172,In_1339,In_1160);
nor U4173 (N_4173,In_1794,In_115);
nand U4174 (N_4174,In_884,In_1339);
or U4175 (N_4175,In_1320,In_681);
or U4176 (N_4176,In_1069,In_701);
nor U4177 (N_4177,In_179,In_118);
or U4178 (N_4178,In_1014,In_1648);
nand U4179 (N_4179,In_749,In_189);
or U4180 (N_4180,In_1076,In_1518);
and U4181 (N_4181,In_1115,In_849);
or U4182 (N_4182,In_1322,In_47);
or U4183 (N_4183,In_1832,In_1614);
or U4184 (N_4184,In_427,In_266);
nand U4185 (N_4185,In_1864,In_972);
and U4186 (N_4186,In_1287,In_998);
nand U4187 (N_4187,In_1379,In_51);
and U4188 (N_4188,In_455,In_526);
nor U4189 (N_4189,In_151,In_896);
nand U4190 (N_4190,In_1733,In_1064);
or U4191 (N_4191,In_859,In_326);
nor U4192 (N_4192,In_177,In_1721);
nand U4193 (N_4193,In_1346,In_296);
and U4194 (N_4194,In_356,In_519);
nand U4195 (N_4195,In_1658,In_235);
or U4196 (N_4196,In_1310,In_1189);
or U4197 (N_4197,In_150,In_260);
and U4198 (N_4198,In_1446,In_1467);
or U4199 (N_4199,In_28,In_1988);
nor U4200 (N_4200,In_949,In_171);
nand U4201 (N_4201,In_988,In_1170);
nor U4202 (N_4202,In_1457,In_1609);
or U4203 (N_4203,In_1881,In_1293);
and U4204 (N_4204,In_209,In_619);
nor U4205 (N_4205,In_275,In_315);
nand U4206 (N_4206,In_1460,In_1728);
xnor U4207 (N_4207,In_1069,In_918);
or U4208 (N_4208,In_1404,In_1392);
nor U4209 (N_4209,In_26,In_1931);
nor U4210 (N_4210,In_1,In_1621);
nor U4211 (N_4211,In_1480,In_1660);
nor U4212 (N_4212,In_553,In_1234);
nand U4213 (N_4213,In_188,In_1499);
nor U4214 (N_4214,In_1259,In_734);
or U4215 (N_4215,In_575,In_1694);
nor U4216 (N_4216,In_648,In_1387);
and U4217 (N_4217,In_600,In_608);
or U4218 (N_4218,In_236,In_1490);
nor U4219 (N_4219,In_1129,In_1227);
or U4220 (N_4220,In_1468,In_793);
and U4221 (N_4221,In_1921,In_1924);
and U4222 (N_4222,In_1716,In_1973);
nor U4223 (N_4223,In_1883,In_920);
and U4224 (N_4224,In_932,In_419);
or U4225 (N_4225,In_348,In_1966);
nand U4226 (N_4226,In_300,In_1073);
nor U4227 (N_4227,In_1171,In_309);
nand U4228 (N_4228,In_216,In_1797);
and U4229 (N_4229,In_1525,In_1615);
nor U4230 (N_4230,In_716,In_426);
or U4231 (N_4231,In_546,In_1640);
and U4232 (N_4232,In_177,In_744);
and U4233 (N_4233,In_158,In_634);
or U4234 (N_4234,In_117,In_520);
and U4235 (N_4235,In_442,In_14);
xnor U4236 (N_4236,In_1598,In_43);
nor U4237 (N_4237,In_1486,In_469);
nand U4238 (N_4238,In_786,In_1151);
and U4239 (N_4239,In_597,In_350);
xnor U4240 (N_4240,In_1517,In_1157);
or U4241 (N_4241,In_1105,In_1359);
and U4242 (N_4242,In_1027,In_1235);
nand U4243 (N_4243,In_495,In_1143);
and U4244 (N_4244,In_621,In_1886);
and U4245 (N_4245,In_1180,In_704);
nor U4246 (N_4246,In_311,In_1421);
or U4247 (N_4247,In_1160,In_1786);
or U4248 (N_4248,In_1981,In_1916);
and U4249 (N_4249,In_324,In_1259);
nand U4250 (N_4250,In_1328,In_514);
or U4251 (N_4251,In_131,In_1484);
and U4252 (N_4252,In_450,In_1335);
nand U4253 (N_4253,In_658,In_610);
or U4254 (N_4254,In_698,In_1289);
nand U4255 (N_4255,In_759,In_735);
nand U4256 (N_4256,In_978,In_1100);
and U4257 (N_4257,In_1513,In_787);
xor U4258 (N_4258,In_63,In_1925);
or U4259 (N_4259,In_306,In_1535);
nor U4260 (N_4260,In_807,In_960);
or U4261 (N_4261,In_1936,In_933);
xnor U4262 (N_4262,In_788,In_1513);
nor U4263 (N_4263,In_118,In_1172);
nand U4264 (N_4264,In_1094,In_746);
and U4265 (N_4265,In_379,In_1177);
nand U4266 (N_4266,In_811,In_1183);
and U4267 (N_4267,In_987,In_734);
nor U4268 (N_4268,In_1136,In_687);
or U4269 (N_4269,In_1368,In_1613);
xor U4270 (N_4270,In_1557,In_1519);
and U4271 (N_4271,In_458,In_1699);
or U4272 (N_4272,In_1082,In_1518);
xnor U4273 (N_4273,In_1243,In_439);
and U4274 (N_4274,In_548,In_1050);
and U4275 (N_4275,In_1347,In_1710);
or U4276 (N_4276,In_895,In_480);
or U4277 (N_4277,In_1995,In_62);
nand U4278 (N_4278,In_818,In_498);
and U4279 (N_4279,In_790,In_1068);
nand U4280 (N_4280,In_22,In_674);
nor U4281 (N_4281,In_75,In_982);
or U4282 (N_4282,In_1089,In_1110);
and U4283 (N_4283,In_513,In_1051);
or U4284 (N_4284,In_1172,In_708);
nand U4285 (N_4285,In_792,In_667);
nand U4286 (N_4286,In_1117,In_769);
and U4287 (N_4287,In_1870,In_1504);
xnor U4288 (N_4288,In_253,In_1052);
nand U4289 (N_4289,In_763,In_1277);
and U4290 (N_4290,In_1086,In_391);
or U4291 (N_4291,In_1870,In_1591);
or U4292 (N_4292,In_979,In_1751);
xor U4293 (N_4293,In_1313,In_1905);
and U4294 (N_4294,In_375,In_25);
xnor U4295 (N_4295,In_1232,In_148);
and U4296 (N_4296,In_1731,In_882);
nor U4297 (N_4297,In_1228,In_938);
nand U4298 (N_4298,In_1519,In_1523);
xor U4299 (N_4299,In_1484,In_782);
xnor U4300 (N_4300,In_1088,In_1269);
or U4301 (N_4301,In_1155,In_1068);
nand U4302 (N_4302,In_319,In_1425);
or U4303 (N_4303,In_1409,In_1411);
and U4304 (N_4304,In_605,In_1020);
nor U4305 (N_4305,In_1806,In_1890);
nor U4306 (N_4306,In_475,In_1886);
nand U4307 (N_4307,In_1225,In_1595);
nand U4308 (N_4308,In_1517,In_351);
or U4309 (N_4309,In_1642,In_99);
xor U4310 (N_4310,In_239,In_1374);
nor U4311 (N_4311,In_723,In_526);
nand U4312 (N_4312,In_313,In_4);
nand U4313 (N_4313,In_605,In_1212);
nand U4314 (N_4314,In_1407,In_1110);
and U4315 (N_4315,In_575,In_1511);
nor U4316 (N_4316,In_366,In_327);
or U4317 (N_4317,In_820,In_1950);
or U4318 (N_4318,In_909,In_1068);
nor U4319 (N_4319,In_1266,In_1662);
xor U4320 (N_4320,In_1432,In_528);
and U4321 (N_4321,In_1983,In_639);
and U4322 (N_4322,In_561,In_607);
or U4323 (N_4323,In_767,In_1589);
nor U4324 (N_4324,In_496,In_537);
nand U4325 (N_4325,In_1333,In_1052);
xor U4326 (N_4326,In_1087,In_939);
nor U4327 (N_4327,In_1853,In_750);
and U4328 (N_4328,In_1446,In_1506);
xor U4329 (N_4329,In_454,In_23);
and U4330 (N_4330,In_1226,In_600);
nand U4331 (N_4331,In_1039,In_631);
and U4332 (N_4332,In_1836,In_1418);
nor U4333 (N_4333,In_1564,In_313);
and U4334 (N_4334,In_422,In_1384);
or U4335 (N_4335,In_1891,In_531);
nand U4336 (N_4336,In_1036,In_1901);
nand U4337 (N_4337,In_972,In_1597);
nor U4338 (N_4338,In_1540,In_249);
or U4339 (N_4339,In_793,In_1761);
nor U4340 (N_4340,In_648,In_1916);
nor U4341 (N_4341,In_1473,In_324);
nor U4342 (N_4342,In_1433,In_1700);
or U4343 (N_4343,In_1518,In_88);
nand U4344 (N_4344,In_1199,In_99);
nand U4345 (N_4345,In_832,In_1144);
or U4346 (N_4346,In_1740,In_473);
and U4347 (N_4347,In_740,In_117);
and U4348 (N_4348,In_1000,In_1754);
nand U4349 (N_4349,In_1179,In_1701);
nand U4350 (N_4350,In_899,In_499);
or U4351 (N_4351,In_214,In_433);
or U4352 (N_4352,In_1514,In_248);
nand U4353 (N_4353,In_233,In_1898);
nor U4354 (N_4354,In_305,In_1054);
and U4355 (N_4355,In_919,In_85);
xnor U4356 (N_4356,In_62,In_1957);
nor U4357 (N_4357,In_1198,In_1061);
and U4358 (N_4358,In_487,In_336);
and U4359 (N_4359,In_880,In_538);
nand U4360 (N_4360,In_5,In_1254);
xor U4361 (N_4361,In_658,In_390);
nor U4362 (N_4362,In_288,In_629);
xnor U4363 (N_4363,In_985,In_1107);
nor U4364 (N_4364,In_1587,In_452);
nand U4365 (N_4365,In_936,In_1476);
or U4366 (N_4366,In_1215,In_1060);
nand U4367 (N_4367,In_1744,In_349);
nand U4368 (N_4368,In_570,In_1190);
nand U4369 (N_4369,In_340,In_1353);
xnor U4370 (N_4370,In_1621,In_646);
nand U4371 (N_4371,In_955,In_205);
or U4372 (N_4372,In_751,In_1385);
nand U4373 (N_4373,In_249,In_1259);
and U4374 (N_4374,In_404,In_1032);
or U4375 (N_4375,In_874,In_763);
xor U4376 (N_4376,In_914,In_231);
nor U4377 (N_4377,In_1925,In_303);
nand U4378 (N_4378,In_466,In_270);
or U4379 (N_4379,In_1944,In_1455);
nor U4380 (N_4380,In_28,In_245);
or U4381 (N_4381,In_986,In_1027);
nor U4382 (N_4382,In_1580,In_1312);
nor U4383 (N_4383,In_332,In_41);
nor U4384 (N_4384,In_1389,In_1842);
nor U4385 (N_4385,In_1368,In_1006);
nor U4386 (N_4386,In_1698,In_937);
and U4387 (N_4387,In_1320,In_771);
nor U4388 (N_4388,In_74,In_1092);
or U4389 (N_4389,In_77,In_654);
nand U4390 (N_4390,In_947,In_644);
nor U4391 (N_4391,In_392,In_1530);
nor U4392 (N_4392,In_999,In_1792);
or U4393 (N_4393,In_1741,In_571);
nor U4394 (N_4394,In_225,In_1034);
and U4395 (N_4395,In_1659,In_254);
nor U4396 (N_4396,In_789,In_246);
nor U4397 (N_4397,In_1819,In_47);
and U4398 (N_4398,In_1707,In_1796);
xor U4399 (N_4399,In_1635,In_1507);
xnor U4400 (N_4400,In_1627,In_798);
nand U4401 (N_4401,In_535,In_1918);
nor U4402 (N_4402,In_476,In_1119);
or U4403 (N_4403,In_1370,In_686);
nor U4404 (N_4404,In_1356,In_1709);
or U4405 (N_4405,In_683,In_1272);
nand U4406 (N_4406,In_534,In_1694);
nor U4407 (N_4407,In_1,In_95);
xnor U4408 (N_4408,In_1662,In_1779);
nor U4409 (N_4409,In_1782,In_1360);
and U4410 (N_4410,In_434,In_260);
nor U4411 (N_4411,In_1051,In_504);
xor U4412 (N_4412,In_548,In_907);
and U4413 (N_4413,In_130,In_1188);
nand U4414 (N_4414,In_1423,In_1513);
or U4415 (N_4415,In_410,In_1373);
and U4416 (N_4416,In_1045,In_216);
or U4417 (N_4417,In_124,In_1854);
nand U4418 (N_4418,In_1228,In_1311);
nor U4419 (N_4419,In_1573,In_1951);
nor U4420 (N_4420,In_1931,In_1588);
nand U4421 (N_4421,In_1669,In_1597);
and U4422 (N_4422,In_145,In_67);
nand U4423 (N_4423,In_1272,In_840);
nand U4424 (N_4424,In_663,In_1473);
and U4425 (N_4425,In_1628,In_210);
nor U4426 (N_4426,In_458,In_1557);
nor U4427 (N_4427,In_1664,In_1672);
or U4428 (N_4428,In_1532,In_1281);
nand U4429 (N_4429,In_357,In_1267);
nand U4430 (N_4430,In_1757,In_1338);
and U4431 (N_4431,In_810,In_1007);
nand U4432 (N_4432,In_1292,In_725);
and U4433 (N_4433,In_1174,In_909);
nor U4434 (N_4434,In_1167,In_1433);
or U4435 (N_4435,In_25,In_130);
nand U4436 (N_4436,In_166,In_228);
nand U4437 (N_4437,In_1391,In_1323);
xnor U4438 (N_4438,In_1735,In_1186);
or U4439 (N_4439,In_1241,In_995);
and U4440 (N_4440,In_85,In_343);
nor U4441 (N_4441,In_32,In_813);
or U4442 (N_4442,In_272,In_1440);
and U4443 (N_4443,In_1853,In_1768);
xnor U4444 (N_4444,In_1116,In_141);
or U4445 (N_4445,In_1996,In_606);
or U4446 (N_4446,In_710,In_920);
or U4447 (N_4447,In_93,In_1339);
or U4448 (N_4448,In_1499,In_554);
nor U4449 (N_4449,In_613,In_1765);
and U4450 (N_4450,In_1780,In_1085);
nand U4451 (N_4451,In_1275,In_1122);
or U4452 (N_4452,In_558,In_1745);
or U4453 (N_4453,In_1218,In_367);
xnor U4454 (N_4454,In_1215,In_244);
nand U4455 (N_4455,In_5,In_117);
and U4456 (N_4456,In_701,In_1424);
and U4457 (N_4457,In_586,In_1271);
nand U4458 (N_4458,In_58,In_332);
nor U4459 (N_4459,In_929,In_684);
nor U4460 (N_4460,In_1505,In_547);
and U4461 (N_4461,In_609,In_1489);
nor U4462 (N_4462,In_844,In_247);
and U4463 (N_4463,In_115,In_1892);
and U4464 (N_4464,In_183,In_550);
or U4465 (N_4465,In_1223,In_1645);
nand U4466 (N_4466,In_396,In_1219);
nand U4467 (N_4467,In_387,In_957);
nand U4468 (N_4468,In_1866,In_1550);
xnor U4469 (N_4469,In_487,In_28);
nor U4470 (N_4470,In_119,In_669);
nand U4471 (N_4471,In_418,In_377);
xor U4472 (N_4472,In_863,In_1874);
or U4473 (N_4473,In_1463,In_375);
nand U4474 (N_4474,In_813,In_1715);
or U4475 (N_4475,In_1369,In_424);
nor U4476 (N_4476,In_413,In_1174);
and U4477 (N_4477,In_201,In_1686);
and U4478 (N_4478,In_309,In_824);
and U4479 (N_4479,In_1299,In_0);
or U4480 (N_4480,In_1527,In_668);
or U4481 (N_4481,In_957,In_267);
xnor U4482 (N_4482,In_1550,In_1743);
nand U4483 (N_4483,In_1725,In_1189);
nand U4484 (N_4484,In_1863,In_1603);
nor U4485 (N_4485,In_1328,In_1685);
nand U4486 (N_4486,In_1792,In_1285);
and U4487 (N_4487,In_701,In_1753);
and U4488 (N_4488,In_1020,In_459);
nor U4489 (N_4489,In_1190,In_1296);
nand U4490 (N_4490,In_251,In_1719);
nand U4491 (N_4491,In_1686,In_1719);
xor U4492 (N_4492,In_1655,In_1092);
nor U4493 (N_4493,In_1485,In_73);
or U4494 (N_4494,In_94,In_703);
or U4495 (N_4495,In_1136,In_779);
nor U4496 (N_4496,In_793,In_1835);
or U4497 (N_4497,In_1343,In_491);
nor U4498 (N_4498,In_1511,In_283);
or U4499 (N_4499,In_314,In_150);
and U4500 (N_4500,In_769,In_1028);
and U4501 (N_4501,In_833,In_135);
and U4502 (N_4502,In_633,In_1855);
or U4503 (N_4503,In_151,In_1261);
or U4504 (N_4504,In_716,In_246);
or U4505 (N_4505,In_289,In_778);
or U4506 (N_4506,In_917,In_261);
nor U4507 (N_4507,In_1532,In_68);
xnor U4508 (N_4508,In_1939,In_137);
xor U4509 (N_4509,In_429,In_135);
and U4510 (N_4510,In_628,In_1312);
and U4511 (N_4511,In_1311,In_1271);
nor U4512 (N_4512,In_909,In_1813);
or U4513 (N_4513,In_626,In_799);
or U4514 (N_4514,In_734,In_1758);
or U4515 (N_4515,In_374,In_977);
and U4516 (N_4516,In_1904,In_930);
and U4517 (N_4517,In_649,In_1300);
and U4518 (N_4518,In_1764,In_729);
or U4519 (N_4519,In_1733,In_1960);
nor U4520 (N_4520,In_1489,In_1124);
nand U4521 (N_4521,In_846,In_7);
or U4522 (N_4522,In_106,In_575);
nand U4523 (N_4523,In_42,In_1956);
and U4524 (N_4524,In_1737,In_1121);
or U4525 (N_4525,In_1333,In_1629);
nand U4526 (N_4526,In_1505,In_830);
nand U4527 (N_4527,In_151,In_1460);
and U4528 (N_4528,In_1053,In_260);
or U4529 (N_4529,In_1054,In_256);
xor U4530 (N_4530,In_711,In_1597);
xor U4531 (N_4531,In_741,In_271);
and U4532 (N_4532,In_1209,In_1207);
nor U4533 (N_4533,In_1093,In_216);
and U4534 (N_4534,In_1147,In_1361);
nor U4535 (N_4535,In_185,In_1791);
and U4536 (N_4536,In_314,In_1611);
nor U4537 (N_4537,In_1694,In_52);
xnor U4538 (N_4538,In_1965,In_308);
and U4539 (N_4539,In_1299,In_484);
or U4540 (N_4540,In_655,In_1948);
nand U4541 (N_4541,In_1714,In_863);
and U4542 (N_4542,In_1001,In_1501);
and U4543 (N_4543,In_325,In_111);
nor U4544 (N_4544,In_943,In_251);
and U4545 (N_4545,In_631,In_83);
and U4546 (N_4546,In_264,In_1148);
or U4547 (N_4547,In_651,In_986);
nand U4548 (N_4548,In_102,In_1808);
or U4549 (N_4549,In_195,In_1831);
and U4550 (N_4550,In_1795,In_384);
nor U4551 (N_4551,In_799,In_740);
or U4552 (N_4552,In_758,In_1652);
nor U4553 (N_4553,In_312,In_306);
nor U4554 (N_4554,In_1683,In_1968);
nand U4555 (N_4555,In_945,In_558);
and U4556 (N_4556,In_1348,In_136);
xor U4557 (N_4557,In_1355,In_932);
nand U4558 (N_4558,In_970,In_181);
nor U4559 (N_4559,In_331,In_1660);
and U4560 (N_4560,In_424,In_397);
nor U4561 (N_4561,In_414,In_1796);
xnor U4562 (N_4562,In_450,In_1481);
nand U4563 (N_4563,In_1758,In_987);
or U4564 (N_4564,In_564,In_945);
and U4565 (N_4565,In_755,In_1928);
and U4566 (N_4566,In_1583,In_572);
nand U4567 (N_4567,In_1771,In_1130);
and U4568 (N_4568,In_1868,In_1252);
nand U4569 (N_4569,In_1364,In_46);
and U4570 (N_4570,In_1214,In_73);
nand U4571 (N_4571,In_695,In_1018);
or U4572 (N_4572,In_1823,In_260);
nor U4573 (N_4573,In_1885,In_995);
nand U4574 (N_4574,In_1731,In_1989);
nor U4575 (N_4575,In_1693,In_1429);
xnor U4576 (N_4576,In_1708,In_1501);
xnor U4577 (N_4577,In_1527,In_1565);
or U4578 (N_4578,In_1173,In_464);
xnor U4579 (N_4579,In_393,In_1604);
nor U4580 (N_4580,In_186,In_1593);
or U4581 (N_4581,In_1849,In_1431);
and U4582 (N_4582,In_1623,In_1318);
xor U4583 (N_4583,In_1847,In_463);
and U4584 (N_4584,In_1630,In_1969);
nor U4585 (N_4585,In_718,In_1872);
nand U4586 (N_4586,In_1294,In_641);
and U4587 (N_4587,In_1703,In_1661);
and U4588 (N_4588,In_1661,In_518);
and U4589 (N_4589,In_1528,In_762);
nor U4590 (N_4590,In_1249,In_1203);
and U4591 (N_4591,In_1821,In_1771);
nor U4592 (N_4592,In_289,In_1593);
or U4593 (N_4593,In_1936,In_1157);
nand U4594 (N_4594,In_602,In_434);
and U4595 (N_4595,In_1992,In_987);
nand U4596 (N_4596,In_487,In_394);
xnor U4597 (N_4597,In_474,In_365);
nor U4598 (N_4598,In_1515,In_986);
xnor U4599 (N_4599,In_1336,In_63);
or U4600 (N_4600,In_1739,In_1677);
and U4601 (N_4601,In_666,In_562);
or U4602 (N_4602,In_1412,In_1474);
or U4603 (N_4603,In_638,In_292);
and U4604 (N_4604,In_209,In_1998);
xnor U4605 (N_4605,In_672,In_1102);
and U4606 (N_4606,In_662,In_986);
nor U4607 (N_4607,In_1003,In_1389);
and U4608 (N_4608,In_1913,In_1088);
xor U4609 (N_4609,In_1139,In_1236);
nor U4610 (N_4610,In_826,In_347);
nand U4611 (N_4611,In_929,In_1656);
nor U4612 (N_4612,In_771,In_129);
and U4613 (N_4613,In_1207,In_1663);
and U4614 (N_4614,In_467,In_1089);
nand U4615 (N_4615,In_544,In_1606);
and U4616 (N_4616,In_458,In_475);
and U4617 (N_4617,In_1250,In_1743);
nand U4618 (N_4618,In_1365,In_411);
nor U4619 (N_4619,In_1683,In_1980);
nor U4620 (N_4620,In_1324,In_173);
or U4621 (N_4621,In_1370,In_725);
or U4622 (N_4622,In_928,In_56);
nor U4623 (N_4623,In_1897,In_1688);
nor U4624 (N_4624,In_1831,In_216);
nand U4625 (N_4625,In_153,In_895);
nand U4626 (N_4626,In_411,In_1195);
nand U4627 (N_4627,In_123,In_93);
xnor U4628 (N_4628,In_1475,In_1100);
nand U4629 (N_4629,In_1041,In_656);
xor U4630 (N_4630,In_716,In_92);
nor U4631 (N_4631,In_655,In_516);
nor U4632 (N_4632,In_1885,In_223);
nor U4633 (N_4633,In_1329,In_1195);
nand U4634 (N_4634,In_464,In_1643);
and U4635 (N_4635,In_882,In_1912);
nor U4636 (N_4636,In_1355,In_667);
or U4637 (N_4637,In_457,In_14);
and U4638 (N_4638,In_1555,In_1490);
nor U4639 (N_4639,In_1380,In_1428);
or U4640 (N_4640,In_630,In_319);
and U4641 (N_4641,In_1182,In_39);
xor U4642 (N_4642,In_1103,In_886);
and U4643 (N_4643,In_1005,In_1275);
nor U4644 (N_4644,In_1181,In_8);
nand U4645 (N_4645,In_452,In_889);
and U4646 (N_4646,In_1751,In_505);
nor U4647 (N_4647,In_1630,In_396);
and U4648 (N_4648,In_752,In_1185);
and U4649 (N_4649,In_979,In_118);
nor U4650 (N_4650,In_916,In_1027);
nor U4651 (N_4651,In_1542,In_483);
or U4652 (N_4652,In_1136,In_1143);
and U4653 (N_4653,In_1303,In_119);
nor U4654 (N_4654,In_135,In_554);
or U4655 (N_4655,In_1945,In_546);
xnor U4656 (N_4656,In_412,In_488);
nand U4657 (N_4657,In_118,In_835);
and U4658 (N_4658,In_360,In_1569);
or U4659 (N_4659,In_727,In_1784);
and U4660 (N_4660,In_872,In_1124);
or U4661 (N_4661,In_1230,In_745);
nand U4662 (N_4662,In_71,In_461);
and U4663 (N_4663,In_469,In_1441);
or U4664 (N_4664,In_30,In_670);
or U4665 (N_4665,In_1999,In_1354);
or U4666 (N_4666,In_1697,In_850);
nand U4667 (N_4667,In_1405,In_590);
nand U4668 (N_4668,In_248,In_1525);
and U4669 (N_4669,In_828,In_1044);
nor U4670 (N_4670,In_764,In_1909);
nand U4671 (N_4671,In_1412,In_380);
or U4672 (N_4672,In_1361,In_853);
nand U4673 (N_4673,In_715,In_1930);
or U4674 (N_4674,In_468,In_715);
and U4675 (N_4675,In_1054,In_1765);
and U4676 (N_4676,In_758,In_824);
nor U4677 (N_4677,In_1896,In_873);
nand U4678 (N_4678,In_571,In_628);
or U4679 (N_4679,In_1387,In_1132);
or U4680 (N_4680,In_1501,In_91);
and U4681 (N_4681,In_812,In_378);
nand U4682 (N_4682,In_458,In_1620);
or U4683 (N_4683,In_1739,In_779);
or U4684 (N_4684,In_1213,In_1596);
and U4685 (N_4685,In_1684,In_842);
nor U4686 (N_4686,In_1795,In_784);
or U4687 (N_4687,In_299,In_1637);
and U4688 (N_4688,In_333,In_1135);
and U4689 (N_4689,In_1429,In_1270);
and U4690 (N_4690,In_1908,In_1424);
nor U4691 (N_4691,In_1289,In_932);
nand U4692 (N_4692,In_1673,In_459);
or U4693 (N_4693,In_1988,In_1812);
or U4694 (N_4694,In_994,In_347);
nor U4695 (N_4695,In_1724,In_63);
and U4696 (N_4696,In_1255,In_996);
nand U4697 (N_4697,In_22,In_721);
nor U4698 (N_4698,In_1235,In_1741);
and U4699 (N_4699,In_350,In_1801);
or U4700 (N_4700,In_312,In_1197);
or U4701 (N_4701,In_897,In_767);
or U4702 (N_4702,In_596,In_1022);
and U4703 (N_4703,In_790,In_1695);
nor U4704 (N_4704,In_1306,In_252);
and U4705 (N_4705,In_351,In_105);
and U4706 (N_4706,In_1345,In_1934);
nand U4707 (N_4707,In_234,In_898);
and U4708 (N_4708,In_1057,In_887);
and U4709 (N_4709,In_990,In_1606);
nand U4710 (N_4710,In_1521,In_139);
nand U4711 (N_4711,In_806,In_1305);
nand U4712 (N_4712,In_10,In_391);
and U4713 (N_4713,In_1189,In_873);
and U4714 (N_4714,In_649,In_911);
or U4715 (N_4715,In_117,In_1335);
nor U4716 (N_4716,In_1533,In_67);
and U4717 (N_4717,In_1999,In_983);
nor U4718 (N_4718,In_1832,In_1920);
or U4719 (N_4719,In_1748,In_1367);
nand U4720 (N_4720,In_131,In_597);
nand U4721 (N_4721,In_1259,In_579);
or U4722 (N_4722,In_770,In_121);
xor U4723 (N_4723,In_89,In_1723);
or U4724 (N_4724,In_1990,In_1111);
nor U4725 (N_4725,In_745,In_1243);
nand U4726 (N_4726,In_959,In_973);
and U4727 (N_4727,In_192,In_729);
or U4728 (N_4728,In_1795,In_1609);
nor U4729 (N_4729,In_1653,In_1955);
or U4730 (N_4730,In_1394,In_940);
xor U4731 (N_4731,In_1271,In_1981);
nand U4732 (N_4732,In_61,In_777);
nand U4733 (N_4733,In_1174,In_217);
and U4734 (N_4734,In_92,In_130);
nand U4735 (N_4735,In_479,In_1426);
and U4736 (N_4736,In_1761,In_920);
nor U4737 (N_4737,In_1322,In_813);
nor U4738 (N_4738,In_221,In_826);
nor U4739 (N_4739,In_292,In_882);
and U4740 (N_4740,In_959,In_101);
and U4741 (N_4741,In_97,In_914);
or U4742 (N_4742,In_1165,In_62);
nor U4743 (N_4743,In_1120,In_1366);
and U4744 (N_4744,In_561,In_762);
or U4745 (N_4745,In_1051,In_1792);
nor U4746 (N_4746,In_491,In_738);
nor U4747 (N_4747,In_1613,In_143);
and U4748 (N_4748,In_994,In_1292);
and U4749 (N_4749,In_167,In_418);
nand U4750 (N_4750,In_1220,In_1816);
and U4751 (N_4751,In_1252,In_693);
and U4752 (N_4752,In_1964,In_1450);
or U4753 (N_4753,In_1608,In_1105);
or U4754 (N_4754,In_70,In_1795);
nand U4755 (N_4755,In_816,In_1251);
nor U4756 (N_4756,In_742,In_118);
and U4757 (N_4757,In_177,In_219);
or U4758 (N_4758,In_180,In_1657);
nor U4759 (N_4759,In_262,In_779);
xnor U4760 (N_4760,In_1008,In_1126);
and U4761 (N_4761,In_533,In_1418);
and U4762 (N_4762,In_1606,In_484);
or U4763 (N_4763,In_1656,In_1785);
or U4764 (N_4764,In_1705,In_90);
or U4765 (N_4765,In_916,In_1640);
nand U4766 (N_4766,In_1632,In_1638);
and U4767 (N_4767,In_719,In_392);
nand U4768 (N_4768,In_1066,In_137);
or U4769 (N_4769,In_1415,In_829);
nor U4770 (N_4770,In_1816,In_954);
and U4771 (N_4771,In_2,In_753);
nand U4772 (N_4772,In_145,In_836);
nand U4773 (N_4773,In_217,In_738);
or U4774 (N_4774,In_1188,In_1403);
nand U4775 (N_4775,In_1682,In_743);
nand U4776 (N_4776,In_273,In_435);
or U4777 (N_4777,In_218,In_1172);
or U4778 (N_4778,In_1880,In_1690);
or U4779 (N_4779,In_1173,In_1679);
and U4780 (N_4780,In_1369,In_1063);
nor U4781 (N_4781,In_1743,In_1265);
xnor U4782 (N_4782,In_409,In_1553);
nor U4783 (N_4783,In_745,In_1449);
nand U4784 (N_4784,In_541,In_950);
nor U4785 (N_4785,In_1622,In_1763);
and U4786 (N_4786,In_766,In_1855);
and U4787 (N_4787,In_729,In_1007);
and U4788 (N_4788,In_1463,In_208);
and U4789 (N_4789,In_957,In_103);
nand U4790 (N_4790,In_1262,In_1855);
nor U4791 (N_4791,In_1686,In_432);
and U4792 (N_4792,In_1417,In_559);
xnor U4793 (N_4793,In_1020,In_1651);
nor U4794 (N_4794,In_824,In_1053);
and U4795 (N_4795,In_1461,In_1536);
nand U4796 (N_4796,In_448,In_1133);
xor U4797 (N_4797,In_580,In_377);
or U4798 (N_4798,In_501,In_1780);
nor U4799 (N_4799,In_105,In_1522);
or U4800 (N_4800,In_1140,In_1251);
and U4801 (N_4801,In_1485,In_830);
or U4802 (N_4802,In_31,In_67);
or U4803 (N_4803,In_1388,In_1513);
nor U4804 (N_4804,In_963,In_1683);
nor U4805 (N_4805,In_456,In_60);
nor U4806 (N_4806,In_667,In_365);
and U4807 (N_4807,In_1480,In_44);
xnor U4808 (N_4808,In_527,In_541);
nand U4809 (N_4809,In_850,In_1360);
nor U4810 (N_4810,In_269,In_14);
nor U4811 (N_4811,In_951,In_1308);
or U4812 (N_4812,In_1463,In_1932);
nand U4813 (N_4813,In_723,In_1833);
and U4814 (N_4814,In_232,In_463);
nand U4815 (N_4815,In_1397,In_408);
or U4816 (N_4816,In_1668,In_1746);
or U4817 (N_4817,In_273,In_1911);
or U4818 (N_4818,In_527,In_1813);
or U4819 (N_4819,In_719,In_1561);
nand U4820 (N_4820,In_1081,In_1477);
nor U4821 (N_4821,In_335,In_1013);
and U4822 (N_4822,In_1978,In_1353);
nor U4823 (N_4823,In_866,In_1198);
nor U4824 (N_4824,In_196,In_1062);
nor U4825 (N_4825,In_1975,In_9);
nand U4826 (N_4826,In_1974,In_281);
nand U4827 (N_4827,In_1499,In_1254);
nor U4828 (N_4828,In_1432,In_1596);
nand U4829 (N_4829,In_1395,In_1519);
or U4830 (N_4830,In_197,In_1399);
or U4831 (N_4831,In_212,In_657);
nor U4832 (N_4832,In_481,In_364);
and U4833 (N_4833,In_637,In_884);
xor U4834 (N_4834,In_1016,In_571);
or U4835 (N_4835,In_1366,In_664);
nand U4836 (N_4836,In_1689,In_631);
nor U4837 (N_4837,In_1437,In_816);
nand U4838 (N_4838,In_207,In_717);
and U4839 (N_4839,In_393,In_1138);
nor U4840 (N_4840,In_1811,In_1707);
or U4841 (N_4841,In_113,In_690);
nand U4842 (N_4842,In_1374,In_1900);
and U4843 (N_4843,In_847,In_1578);
or U4844 (N_4844,In_1108,In_864);
or U4845 (N_4845,In_1187,In_247);
nor U4846 (N_4846,In_432,In_1190);
nor U4847 (N_4847,In_133,In_1936);
nor U4848 (N_4848,In_1951,In_625);
or U4849 (N_4849,In_1916,In_529);
or U4850 (N_4850,In_810,In_284);
nor U4851 (N_4851,In_464,In_1680);
and U4852 (N_4852,In_1000,In_1277);
nor U4853 (N_4853,In_1005,In_1973);
xnor U4854 (N_4854,In_183,In_1587);
or U4855 (N_4855,In_1119,In_1264);
nor U4856 (N_4856,In_1270,In_1378);
xnor U4857 (N_4857,In_208,In_1694);
nand U4858 (N_4858,In_1706,In_1521);
and U4859 (N_4859,In_932,In_736);
and U4860 (N_4860,In_1027,In_871);
or U4861 (N_4861,In_1119,In_1863);
nor U4862 (N_4862,In_1996,In_1014);
nor U4863 (N_4863,In_673,In_1608);
nand U4864 (N_4864,In_723,In_1931);
and U4865 (N_4865,In_1734,In_899);
and U4866 (N_4866,In_64,In_842);
nand U4867 (N_4867,In_1255,In_1224);
nand U4868 (N_4868,In_390,In_1401);
nor U4869 (N_4869,In_1889,In_1715);
and U4870 (N_4870,In_1094,In_922);
nor U4871 (N_4871,In_1121,In_1352);
and U4872 (N_4872,In_1347,In_629);
xnor U4873 (N_4873,In_193,In_32);
nand U4874 (N_4874,In_1898,In_1176);
or U4875 (N_4875,In_1029,In_1430);
nand U4876 (N_4876,In_1257,In_306);
or U4877 (N_4877,In_705,In_132);
or U4878 (N_4878,In_510,In_1950);
nor U4879 (N_4879,In_1106,In_1772);
nand U4880 (N_4880,In_1880,In_743);
nand U4881 (N_4881,In_905,In_1240);
and U4882 (N_4882,In_1421,In_434);
nand U4883 (N_4883,In_268,In_1974);
nor U4884 (N_4884,In_993,In_1996);
xnor U4885 (N_4885,In_262,In_1331);
nand U4886 (N_4886,In_1192,In_1020);
and U4887 (N_4887,In_288,In_1239);
or U4888 (N_4888,In_287,In_1138);
or U4889 (N_4889,In_742,In_1029);
and U4890 (N_4890,In_1563,In_693);
and U4891 (N_4891,In_667,In_1684);
and U4892 (N_4892,In_716,In_1641);
or U4893 (N_4893,In_900,In_993);
xor U4894 (N_4894,In_1686,In_1229);
nor U4895 (N_4895,In_719,In_139);
nand U4896 (N_4896,In_1529,In_199);
nor U4897 (N_4897,In_1554,In_888);
nand U4898 (N_4898,In_1026,In_370);
or U4899 (N_4899,In_531,In_400);
and U4900 (N_4900,In_641,In_701);
nor U4901 (N_4901,In_1307,In_1823);
or U4902 (N_4902,In_869,In_1724);
nand U4903 (N_4903,In_731,In_516);
nor U4904 (N_4904,In_93,In_1841);
nor U4905 (N_4905,In_1516,In_1954);
xnor U4906 (N_4906,In_1588,In_1900);
or U4907 (N_4907,In_738,In_117);
nor U4908 (N_4908,In_1003,In_332);
and U4909 (N_4909,In_383,In_590);
nor U4910 (N_4910,In_1972,In_1753);
or U4911 (N_4911,In_713,In_226);
nand U4912 (N_4912,In_1303,In_926);
nand U4913 (N_4913,In_1214,In_1929);
nor U4914 (N_4914,In_947,In_1649);
and U4915 (N_4915,In_1667,In_216);
or U4916 (N_4916,In_633,In_342);
nor U4917 (N_4917,In_917,In_115);
nand U4918 (N_4918,In_1596,In_1983);
nand U4919 (N_4919,In_516,In_1477);
or U4920 (N_4920,In_888,In_1108);
nor U4921 (N_4921,In_515,In_259);
and U4922 (N_4922,In_356,In_823);
nand U4923 (N_4923,In_917,In_1140);
or U4924 (N_4924,In_1596,In_72);
nand U4925 (N_4925,In_86,In_116);
or U4926 (N_4926,In_350,In_699);
nand U4927 (N_4927,In_459,In_418);
nor U4928 (N_4928,In_1618,In_718);
and U4929 (N_4929,In_1593,In_792);
nand U4930 (N_4930,In_1012,In_1491);
nand U4931 (N_4931,In_307,In_1019);
nand U4932 (N_4932,In_462,In_1055);
nand U4933 (N_4933,In_1366,In_351);
nor U4934 (N_4934,In_1984,In_1043);
nand U4935 (N_4935,In_796,In_1717);
nor U4936 (N_4936,In_1548,In_271);
and U4937 (N_4937,In_688,In_877);
nand U4938 (N_4938,In_323,In_1358);
nand U4939 (N_4939,In_1125,In_1932);
nand U4940 (N_4940,In_193,In_796);
nand U4941 (N_4941,In_1036,In_338);
nor U4942 (N_4942,In_1560,In_1932);
nor U4943 (N_4943,In_1253,In_1224);
nand U4944 (N_4944,In_1140,In_830);
nor U4945 (N_4945,In_1458,In_285);
xnor U4946 (N_4946,In_1214,In_823);
nor U4947 (N_4947,In_434,In_1716);
nand U4948 (N_4948,In_72,In_1622);
nand U4949 (N_4949,In_452,In_971);
nor U4950 (N_4950,In_1920,In_1268);
nand U4951 (N_4951,In_1904,In_1022);
or U4952 (N_4952,In_523,In_699);
and U4953 (N_4953,In_654,In_376);
and U4954 (N_4954,In_280,In_1253);
and U4955 (N_4955,In_1855,In_1609);
xor U4956 (N_4956,In_979,In_1020);
or U4957 (N_4957,In_370,In_1774);
nand U4958 (N_4958,In_1303,In_1350);
and U4959 (N_4959,In_303,In_1801);
nand U4960 (N_4960,In_597,In_1021);
and U4961 (N_4961,In_285,In_1418);
or U4962 (N_4962,In_1700,In_804);
xor U4963 (N_4963,In_1979,In_960);
xnor U4964 (N_4964,In_1613,In_505);
xor U4965 (N_4965,In_1731,In_671);
and U4966 (N_4966,In_1019,In_634);
nand U4967 (N_4967,In_1831,In_1954);
nor U4968 (N_4968,In_1902,In_1294);
or U4969 (N_4969,In_270,In_437);
nand U4970 (N_4970,In_801,In_218);
or U4971 (N_4971,In_1608,In_1233);
nor U4972 (N_4972,In_1029,In_158);
nand U4973 (N_4973,In_1660,In_1412);
nor U4974 (N_4974,In_1230,In_1043);
or U4975 (N_4975,In_284,In_1000);
or U4976 (N_4976,In_873,In_39);
nand U4977 (N_4977,In_1049,In_1332);
or U4978 (N_4978,In_875,In_1547);
or U4979 (N_4979,In_246,In_1978);
nand U4980 (N_4980,In_814,In_152);
and U4981 (N_4981,In_1178,In_746);
xor U4982 (N_4982,In_150,In_1740);
nor U4983 (N_4983,In_6,In_142);
or U4984 (N_4984,In_1431,In_1151);
nand U4985 (N_4985,In_543,In_897);
nor U4986 (N_4986,In_1053,In_919);
or U4987 (N_4987,In_313,In_1137);
xnor U4988 (N_4988,In_1946,In_763);
nand U4989 (N_4989,In_635,In_1398);
xnor U4990 (N_4990,In_944,In_1753);
nor U4991 (N_4991,In_429,In_1376);
or U4992 (N_4992,In_865,In_285);
nor U4993 (N_4993,In_1166,In_515);
nor U4994 (N_4994,In_1173,In_302);
nor U4995 (N_4995,In_1217,In_1929);
xor U4996 (N_4996,In_1389,In_103);
and U4997 (N_4997,In_1056,In_682);
nand U4998 (N_4998,In_458,In_1864);
and U4999 (N_4999,In_441,In_984);
nor U5000 (N_5000,N_335,N_2206);
or U5001 (N_5001,N_3235,N_4970);
nor U5002 (N_5002,N_4078,N_4533);
nand U5003 (N_5003,N_3281,N_3871);
and U5004 (N_5004,N_60,N_4832);
and U5005 (N_5005,N_3991,N_2633);
nor U5006 (N_5006,N_419,N_4587);
xor U5007 (N_5007,N_909,N_4354);
and U5008 (N_5008,N_3835,N_1364);
or U5009 (N_5009,N_1560,N_4611);
or U5010 (N_5010,N_4346,N_3628);
and U5011 (N_5011,N_4080,N_1758);
nor U5012 (N_5012,N_2954,N_3095);
xnor U5013 (N_5013,N_2910,N_740);
and U5014 (N_5014,N_1318,N_3968);
and U5015 (N_5015,N_1368,N_1936);
or U5016 (N_5016,N_3294,N_2014);
and U5017 (N_5017,N_4675,N_3403);
and U5018 (N_5018,N_2827,N_1021);
or U5019 (N_5019,N_1717,N_754);
nor U5020 (N_5020,N_130,N_1213);
or U5021 (N_5021,N_3076,N_4215);
and U5022 (N_5022,N_4695,N_1703);
and U5023 (N_5023,N_3543,N_4418);
or U5024 (N_5024,N_2375,N_2933);
and U5025 (N_5025,N_4086,N_3614);
nor U5026 (N_5026,N_2184,N_2571);
and U5027 (N_5027,N_3387,N_1518);
xor U5028 (N_5028,N_1523,N_488);
and U5029 (N_5029,N_4170,N_230);
nand U5030 (N_5030,N_1533,N_4706);
nor U5031 (N_5031,N_4121,N_2779);
nor U5032 (N_5032,N_1556,N_3106);
nand U5033 (N_5033,N_644,N_2890);
and U5034 (N_5034,N_4775,N_4136);
nor U5035 (N_5035,N_530,N_2222);
nor U5036 (N_5036,N_1952,N_1883);
nand U5037 (N_5037,N_464,N_2036);
nor U5038 (N_5038,N_2413,N_1946);
nor U5039 (N_5039,N_14,N_839);
or U5040 (N_5040,N_1100,N_225);
or U5041 (N_5041,N_2677,N_66);
nand U5042 (N_5042,N_1082,N_371);
and U5043 (N_5043,N_2336,N_1462);
nand U5044 (N_5044,N_2983,N_4253);
nand U5045 (N_5045,N_1696,N_4765);
or U5046 (N_5046,N_4804,N_3083);
nor U5047 (N_5047,N_2021,N_2869);
nor U5048 (N_5048,N_435,N_1410);
or U5049 (N_5049,N_1067,N_3735);
or U5050 (N_5050,N_4490,N_2703);
or U5051 (N_5051,N_3572,N_2050);
nand U5052 (N_5052,N_1215,N_980);
xnor U5053 (N_5053,N_1610,N_4925);
or U5054 (N_5054,N_3715,N_1422);
nor U5055 (N_5055,N_1712,N_3452);
and U5056 (N_5056,N_2360,N_3092);
nand U5057 (N_5057,N_1894,N_905);
or U5058 (N_5058,N_291,N_4727);
xnor U5059 (N_5059,N_2108,N_1643);
and U5060 (N_5060,N_3872,N_3649);
or U5061 (N_5061,N_3493,N_1976);
or U5062 (N_5062,N_3336,N_2187);
and U5063 (N_5063,N_4333,N_3373);
or U5064 (N_5064,N_2028,N_3656);
nand U5065 (N_5065,N_760,N_4338);
or U5066 (N_5066,N_3667,N_2864);
nor U5067 (N_5067,N_1730,N_182);
or U5068 (N_5068,N_3044,N_2225);
and U5069 (N_5069,N_4374,N_3950);
or U5070 (N_5070,N_1110,N_4563);
or U5071 (N_5071,N_611,N_1459);
or U5072 (N_5072,N_4380,N_3003);
nor U5073 (N_5073,N_3560,N_1474);
or U5074 (N_5074,N_2971,N_3623);
or U5075 (N_5075,N_609,N_3248);
nor U5076 (N_5076,N_4502,N_1022);
nand U5077 (N_5077,N_2536,N_4305);
or U5078 (N_5078,N_3783,N_3876);
nand U5079 (N_5079,N_910,N_4123);
and U5080 (N_5080,N_3957,N_332);
and U5081 (N_5081,N_2938,N_3392);
nor U5082 (N_5082,N_1287,N_1588);
or U5083 (N_5083,N_1958,N_1158);
and U5084 (N_5084,N_2806,N_2425);
nand U5085 (N_5085,N_391,N_1253);
nand U5086 (N_5086,N_4439,N_2907);
and U5087 (N_5087,N_527,N_895);
or U5088 (N_5088,N_1688,N_2404);
or U5089 (N_5089,N_1687,N_2932);
xnor U5090 (N_5090,N_4024,N_4169);
nand U5091 (N_5091,N_276,N_2766);
xnor U5092 (N_5092,N_3145,N_56);
and U5093 (N_5093,N_505,N_1385);
xor U5094 (N_5094,N_3507,N_2196);
nor U5095 (N_5095,N_545,N_1152);
nand U5096 (N_5096,N_1695,N_3684);
nand U5097 (N_5097,N_4441,N_1365);
xnor U5098 (N_5098,N_4552,N_3974);
and U5099 (N_5099,N_2317,N_1845);
or U5100 (N_5100,N_852,N_3492);
nor U5101 (N_5101,N_1141,N_451);
nor U5102 (N_5102,N_625,N_3444);
nand U5103 (N_5103,N_3247,N_1757);
xor U5104 (N_5104,N_3554,N_637);
xor U5105 (N_5105,N_3813,N_3326);
and U5106 (N_5106,N_1162,N_1200);
or U5107 (N_5107,N_2666,N_2331);
and U5108 (N_5108,N_4782,N_283);
nand U5109 (N_5109,N_1642,N_359);
nand U5110 (N_5110,N_503,N_4800);
nor U5111 (N_5111,N_2884,N_3439);
nand U5112 (N_5112,N_3243,N_2001);
nand U5113 (N_5113,N_1995,N_378);
and U5114 (N_5114,N_390,N_783);
xor U5115 (N_5115,N_4688,N_1906);
or U5116 (N_5116,N_1148,N_3435);
or U5117 (N_5117,N_2032,N_2318);
or U5118 (N_5118,N_3450,N_701);
nand U5119 (N_5119,N_1443,N_1137);
nand U5120 (N_5120,N_2307,N_2248);
nand U5121 (N_5121,N_3581,N_395);
nand U5122 (N_5122,N_2922,N_1825);
nand U5123 (N_5123,N_4684,N_4151);
or U5124 (N_5124,N_2093,N_2727);
nand U5125 (N_5125,N_1028,N_3255);
and U5126 (N_5126,N_2981,N_2111);
xnor U5127 (N_5127,N_4081,N_2661);
nor U5128 (N_5128,N_2247,N_953);
or U5129 (N_5129,N_549,N_878);
or U5130 (N_5130,N_747,N_937);
or U5131 (N_5131,N_2641,N_1615);
xor U5132 (N_5132,N_3696,N_875);
xnor U5133 (N_5133,N_1093,N_3756);
and U5134 (N_5134,N_2623,N_3812);
and U5135 (N_5135,N_2059,N_3595);
nand U5136 (N_5136,N_4031,N_1829);
or U5137 (N_5137,N_1744,N_1786);
and U5138 (N_5138,N_612,N_1759);
xnor U5139 (N_5139,N_3998,N_4340);
nand U5140 (N_5140,N_2923,N_1500);
xnor U5141 (N_5141,N_1037,N_69);
nand U5142 (N_5142,N_4993,N_4063);
or U5143 (N_5143,N_3993,N_3527);
xnor U5144 (N_5144,N_536,N_18);
and U5145 (N_5145,N_3863,N_2557);
xor U5146 (N_5146,N_2878,N_1236);
xnor U5147 (N_5147,N_1899,N_4022);
nor U5148 (N_5148,N_4279,N_2485);
or U5149 (N_5149,N_4382,N_2700);
or U5150 (N_5150,N_1671,N_227);
or U5151 (N_5151,N_3068,N_3348);
or U5152 (N_5152,N_4754,N_4846);
and U5153 (N_5153,N_257,N_4485);
nand U5154 (N_5154,N_4983,N_3563);
or U5155 (N_5155,N_4069,N_1078);
and U5156 (N_5156,N_4852,N_1961);
and U5157 (N_5157,N_4650,N_983);
or U5158 (N_5158,N_2670,N_1809);
nor U5159 (N_5159,N_2467,N_935);
or U5160 (N_5160,N_3385,N_1423);
nor U5161 (N_5161,N_3358,N_4486);
and U5162 (N_5162,N_3807,N_1822);
nor U5163 (N_5163,N_1724,N_4957);
or U5164 (N_5164,N_116,N_886);
nand U5165 (N_5165,N_3246,N_3569);
xnor U5166 (N_5166,N_434,N_2889);
or U5167 (N_5167,N_3006,N_3074);
or U5168 (N_5168,N_1404,N_109);
nor U5169 (N_5169,N_4634,N_328);
or U5170 (N_5170,N_985,N_2117);
or U5171 (N_5171,N_4239,N_2495);
or U5172 (N_5172,N_2064,N_2537);
nor U5173 (N_5173,N_4373,N_3308);
nand U5174 (N_5174,N_1699,N_471);
nand U5175 (N_5175,N_982,N_1354);
and U5176 (N_5176,N_2015,N_4434);
or U5177 (N_5177,N_2646,N_2601);
nand U5178 (N_5178,N_2740,N_3672);
nand U5179 (N_5179,N_2063,N_4958);
nand U5180 (N_5180,N_845,N_2514);
nand U5181 (N_5181,N_1979,N_3830);
and U5182 (N_5182,N_3153,N_3458);
nor U5183 (N_5183,N_2974,N_58);
and U5184 (N_5184,N_3191,N_2385);
nand U5185 (N_5185,N_946,N_581);
nand U5186 (N_5186,N_3056,N_745);
or U5187 (N_5187,N_896,N_816);
nor U5188 (N_5188,N_4256,N_2316);
nand U5189 (N_5189,N_3982,N_4990);
nor U5190 (N_5190,N_2739,N_41);
and U5191 (N_5191,N_240,N_2272);
nor U5192 (N_5192,N_3662,N_1366);
or U5193 (N_5193,N_829,N_4351);
xor U5194 (N_5194,N_2065,N_3639);
or U5195 (N_5195,N_258,N_50);
nor U5196 (N_5196,N_254,N_2873);
nor U5197 (N_5197,N_3967,N_3604);
or U5198 (N_5198,N_924,N_2851);
nor U5199 (N_5199,N_2148,N_4898);
nand U5200 (N_5200,N_1277,N_3949);
xor U5201 (N_5201,N_3596,N_4263);
nand U5202 (N_5202,N_3529,N_2928);
nor U5203 (N_5203,N_3360,N_3169);
xor U5204 (N_5204,N_649,N_1700);
xnor U5205 (N_5205,N_734,N_4007);
nor U5206 (N_5206,N_1004,N_1174);
and U5207 (N_5207,N_3988,N_3794);
nand U5208 (N_5208,N_718,N_3291);
nand U5209 (N_5209,N_3231,N_432);
nor U5210 (N_5210,N_166,N_2203);
and U5211 (N_5211,N_2708,N_1993);
nor U5212 (N_5212,N_4411,N_696);
nand U5213 (N_5213,N_674,N_3111);
xnor U5214 (N_5214,N_4937,N_1994);
xnor U5215 (N_5215,N_2023,N_4058);
nor U5216 (N_5216,N_1967,N_4896);
nand U5217 (N_5217,N_1559,N_408);
nand U5218 (N_5218,N_3061,N_2378);
or U5219 (N_5219,N_4692,N_3587);
or U5220 (N_5220,N_2657,N_2113);
nand U5221 (N_5221,N_3082,N_2039);
nor U5222 (N_5222,N_2343,N_4402);
and U5223 (N_5223,N_215,N_1951);
nor U5224 (N_5224,N_202,N_2814);
nor U5225 (N_5225,N_736,N_1090);
or U5226 (N_5226,N_2783,N_3320);
nor U5227 (N_5227,N_873,N_4468);
and U5228 (N_5228,N_1864,N_791);
or U5229 (N_5229,N_2562,N_1346);
or U5230 (N_5230,N_1477,N_1298);
or U5231 (N_5231,N_4026,N_3188);
nand U5232 (N_5232,N_1733,N_1847);
nor U5233 (N_5233,N_1050,N_978);
and U5234 (N_5234,N_4674,N_2704);
nor U5235 (N_5235,N_2384,N_3112);
nor U5236 (N_5236,N_4772,N_1096);
nand U5237 (N_5237,N_3953,N_520);
nor U5238 (N_5238,N_4396,N_309);
nand U5239 (N_5239,N_2790,N_3087);
or U5240 (N_5240,N_2813,N_430);
and U5241 (N_5241,N_3409,N_3043);
nand U5242 (N_5242,N_1449,N_1187);
nand U5243 (N_5243,N_2199,N_3155);
nand U5244 (N_5244,N_1268,N_4819);
nand U5245 (N_5245,N_2699,N_4851);
nor U5246 (N_5246,N_744,N_3448);
nor U5247 (N_5247,N_385,N_1997);
or U5248 (N_5248,N_2939,N_2609);
nand U5249 (N_5249,N_4385,N_513);
or U5250 (N_5250,N_1038,N_3738);
or U5251 (N_5251,N_2638,N_1718);
and U5252 (N_5252,N_2642,N_758);
or U5253 (N_5253,N_4831,N_4590);
nor U5254 (N_5254,N_4522,N_1032);
nor U5255 (N_5255,N_3548,N_1587);
and U5256 (N_5256,N_346,N_775);
nor U5257 (N_5257,N_822,N_1930);
nor U5258 (N_5258,N_1125,N_813);
or U5259 (N_5259,N_3904,N_4391);
or U5260 (N_5260,N_337,N_2911);
and U5261 (N_5261,N_4747,N_2718);
xnor U5262 (N_5262,N_149,N_3339);
or U5263 (N_5263,N_771,N_4091);
or U5264 (N_5264,N_2845,N_3441);
xnor U5265 (N_5265,N_711,N_2521);
and U5266 (N_5266,N_2816,N_1296);
nor U5267 (N_5267,N_947,N_2269);
or U5268 (N_5268,N_2453,N_3838);
nor U5269 (N_5269,N_2150,N_1720);
or U5270 (N_5270,N_3330,N_2287);
nand U5271 (N_5271,N_4821,N_4888);
nand U5272 (N_5272,N_4792,N_2252);
and U5273 (N_5273,N_119,N_2391);
and U5274 (N_5274,N_1797,N_586);
or U5275 (N_5275,N_962,N_2879);
and U5276 (N_5276,N_957,N_1063);
or U5277 (N_5277,N_3364,N_4342);
nor U5278 (N_5278,N_659,N_154);
nand U5279 (N_5279,N_3026,N_615);
nand U5280 (N_5280,N_3005,N_4483);
nand U5281 (N_5281,N_4004,N_4273);
nand U5282 (N_5282,N_4269,N_1113);
and U5283 (N_5283,N_2305,N_2535);
or U5284 (N_5284,N_2573,N_722);
nand U5285 (N_5285,N_1992,N_406);
or U5286 (N_5286,N_3487,N_4267);
or U5287 (N_5287,N_4795,N_1424);
nor U5288 (N_5288,N_969,N_3750);
nand U5289 (N_5289,N_2842,N_3937);
nand U5290 (N_5290,N_4050,N_2198);
nor U5291 (N_5291,N_2990,N_4566);
or U5292 (N_5292,N_4619,N_427);
or U5293 (N_5293,N_4641,N_3862);
and U5294 (N_5294,N_1099,N_3668);
and U5295 (N_5295,N_2988,N_2451);
nor U5296 (N_5296,N_29,N_1458);
and U5297 (N_5297,N_1046,N_2099);
nor U5298 (N_5298,N_1824,N_1973);
or U5299 (N_5299,N_1425,N_2658);
and U5300 (N_5300,N_1095,N_3372);
nand U5301 (N_5301,N_1812,N_4099);
nor U5302 (N_5302,N_894,N_1389);
nand U5303 (N_5303,N_392,N_2811);
xnor U5304 (N_5304,N_4551,N_1059);
and U5305 (N_5305,N_4953,N_3867);
and U5306 (N_5306,N_968,N_3350);
or U5307 (N_5307,N_1432,N_572);
or U5308 (N_5308,N_893,N_640);
and U5309 (N_5309,N_2325,N_1494);
nand U5310 (N_5310,N_2242,N_790);
nor U5311 (N_5311,N_4096,N_1195);
or U5312 (N_5312,N_1060,N_4150);
nand U5313 (N_5313,N_1819,N_4968);
and U5314 (N_5314,N_3468,N_793);
nand U5315 (N_5315,N_1535,N_769);
nor U5316 (N_5316,N_4886,N_3710);
nor U5317 (N_5317,N_163,N_445);
nor U5318 (N_5318,N_4778,N_3821);
nand U5319 (N_5319,N_4447,N_1854);
and U5320 (N_5320,N_882,N_3483);
nand U5321 (N_5321,N_2430,N_17);
or U5322 (N_5322,N_3140,N_2868);
or U5323 (N_5323,N_4862,N_2957);
nor U5324 (N_5324,N_4513,N_3144);
or U5325 (N_5325,N_2625,N_3718);
nand U5326 (N_5326,N_4508,N_3340);
nand U5327 (N_5327,N_2075,N_2155);
and U5328 (N_5328,N_4055,N_370);
and U5329 (N_5329,N_4087,N_3524);
nor U5330 (N_5330,N_3546,N_4609);
or U5331 (N_5331,N_3784,N_622);
and U5332 (N_5332,N_933,N_3240);
nand U5333 (N_5333,N_1278,N_125);
nor U5334 (N_5334,N_1115,N_2082);
nor U5335 (N_5335,N_27,N_3020);
xor U5336 (N_5336,N_277,N_2559);
and U5337 (N_5337,N_1517,N_2256);
or U5338 (N_5338,N_4331,N_607);
or U5339 (N_5339,N_1889,N_2652);
and U5340 (N_5340,N_3307,N_150);
nand U5341 (N_5341,N_305,N_1878);
nand U5342 (N_5342,N_552,N_4221);
or U5343 (N_5343,N_563,N_4319);
and U5344 (N_5344,N_2607,N_2892);
and U5345 (N_5345,N_815,N_1971);
xnor U5346 (N_5346,N_2950,N_511);
xnor U5347 (N_5347,N_4006,N_3405);
nor U5348 (N_5348,N_2731,N_1495);
and U5349 (N_5349,N_1690,N_727);
and U5350 (N_5350,N_4152,N_1574);
nand U5351 (N_5351,N_1439,N_3533);
or U5352 (N_5352,N_4451,N_498);
and U5353 (N_5353,N_2751,N_2750);
nand U5354 (N_5354,N_2960,N_3895);
and U5355 (N_5355,N_3171,N_2278);
nand U5356 (N_5356,N_1913,N_749);
xor U5357 (N_5357,N_1624,N_2526);
or U5358 (N_5358,N_314,N_3592);
or U5359 (N_5359,N_2088,N_2179);
or U5360 (N_5360,N_444,N_4518);
or U5361 (N_5361,N_3707,N_2024);
or U5362 (N_5362,N_1820,N_1804);
or U5363 (N_5363,N_602,N_4876);
nand U5364 (N_5364,N_3959,N_2441);
and U5365 (N_5365,N_282,N_3086);
xor U5366 (N_5366,N_2840,N_2297);
and U5367 (N_5367,N_3397,N_2763);
nand U5368 (N_5368,N_2204,N_1303);
and U5369 (N_5369,N_2935,N_1416);
nor U5370 (N_5370,N_3841,N_88);
nor U5371 (N_5371,N_1035,N_2729);
nor U5372 (N_5372,N_192,N_4089);
and U5373 (N_5373,N_3719,N_3627);
and U5374 (N_5374,N_1515,N_1904);
and U5375 (N_5375,N_2984,N_152);
and U5376 (N_5376,N_2241,N_2645);
xor U5377 (N_5377,N_990,N_4703);
nand U5378 (N_5378,N_4435,N_1168);
and U5379 (N_5379,N_4270,N_4394);
and U5380 (N_5380,N_2566,N_3499);
nor U5381 (N_5381,N_3598,N_151);
or U5382 (N_5382,N_3190,N_591);
nor U5383 (N_5383,N_3416,N_4217);
xor U5384 (N_5384,N_2386,N_2785);
nor U5385 (N_5385,N_1903,N_1034);
nand U5386 (N_5386,N_110,N_2857);
nand U5387 (N_5387,N_401,N_4978);
nand U5388 (N_5388,N_2107,N_3424);
or U5389 (N_5389,N_2992,N_789);
and U5390 (N_5390,N_4458,N_1939);
nor U5391 (N_5391,N_2351,N_3857);
nand U5392 (N_5392,N_2273,N_2492);
and U5393 (N_5393,N_1965,N_4807);
nand U5394 (N_5394,N_3651,N_1706);
or U5395 (N_5395,N_2207,N_3067);
nor U5396 (N_5396,N_2730,N_2512);
nor U5397 (N_5397,N_4728,N_2934);
and U5398 (N_5398,N_1333,N_3525);
and U5399 (N_5399,N_1496,N_3943);
or U5400 (N_5400,N_3636,N_2650);
and U5401 (N_5401,N_1595,N_584);
nand U5402 (N_5402,N_3842,N_1437);
xnor U5403 (N_5403,N_4034,N_660);
and U5404 (N_5404,N_837,N_115);
nand U5405 (N_5405,N_928,N_2587);
nand U5406 (N_5406,N_4143,N_4226);
and U5407 (N_5407,N_3726,N_4177);
and U5408 (N_5408,N_2126,N_3365);
or U5409 (N_5409,N_2815,N_2583);
and U5410 (N_5410,N_3917,N_4500);
or U5411 (N_5411,N_189,N_3378);
and U5412 (N_5412,N_3203,N_4422);
and U5413 (N_5413,N_529,N_2765);
nor U5414 (N_5414,N_2648,N_38);
or U5415 (N_5415,N_1400,N_3304);
and U5416 (N_5416,N_2044,N_2403);
nor U5417 (N_5417,N_1390,N_340);
nor U5418 (N_5418,N_743,N_4859);
or U5419 (N_5419,N_3574,N_4989);
or U5420 (N_5420,N_3605,N_3432);
nor U5421 (N_5421,N_2267,N_2524);
nand U5422 (N_5422,N_3803,N_489);
nor U5423 (N_5423,N_4763,N_23);
nand U5424 (N_5424,N_4017,N_1608);
and U5425 (N_5425,N_4965,N_4148);
or U5426 (N_5426,N_3491,N_3211);
nand U5427 (N_5427,N_2626,N_1937);
or U5428 (N_5428,N_2525,N_4567);
and U5429 (N_5429,N_3591,N_3296);
or U5430 (N_5430,N_440,N_457);
and U5431 (N_5431,N_3096,N_2643);
nand U5432 (N_5432,N_4013,N_805);
and U5433 (N_5433,N_2544,N_1394);
and U5434 (N_5434,N_1161,N_4357);
and U5435 (N_5435,N_1285,N_1506);
and U5436 (N_5436,N_4419,N_721);
nand U5437 (N_5437,N_678,N_507);
nand U5438 (N_5438,N_2158,N_1526);
nor U5439 (N_5439,N_4963,N_4484);
nor U5440 (N_5440,N_3041,N_3576);
nand U5441 (N_5441,N_690,N_1146);
nand U5442 (N_5442,N_2320,N_4849);
and U5443 (N_5443,N_4510,N_4621);
or U5444 (N_5444,N_3028,N_3687);
xor U5445 (N_5445,N_2394,N_1739);
xnor U5446 (N_5446,N_4372,N_4463);
and U5447 (N_5447,N_3966,N_3882);
nor U5448 (N_5448,N_2837,N_3445);
and U5449 (N_5449,N_2594,N_4981);
nor U5450 (N_5450,N_2238,N_4213);
and U5451 (N_5451,N_4079,N_915);
nand U5452 (N_5452,N_1602,N_4171);
and U5453 (N_5453,N_344,N_2527);
nor U5454 (N_5454,N_4444,N_4243);
nand U5455 (N_5455,N_3221,N_1589);
or U5456 (N_5456,N_4071,N_2930);
nor U5457 (N_5457,N_4766,N_4794);
nor U5458 (N_5458,N_4731,N_2617);
and U5459 (N_5459,N_2726,N_3881);
or U5460 (N_5460,N_19,N_1694);
and U5461 (N_5461,N_4790,N_3926);
and U5462 (N_5462,N_522,N_3215);
and U5463 (N_5463,N_3367,N_1692);
nand U5464 (N_5464,N_1257,N_3801);
nand U5465 (N_5465,N_3315,N_1193);
nor U5466 (N_5466,N_841,N_2953);
nor U5467 (N_5467,N_866,N_3864);
or U5468 (N_5468,N_2339,N_1511);
nor U5469 (N_5469,N_3553,N_1293);
nor U5470 (N_5470,N_4604,N_952);
or U5471 (N_5471,N_97,N_1565);
nand U5472 (N_5472,N_4142,N_3705);
or U5473 (N_5473,N_1877,N_4139);
nor U5474 (N_5474,N_3013,N_1861);
and U5475 (N_5475,N_2639,N_3739);
nor U5476 (N_5476,N_4205,N_3342);
nand U5477 (N_5477,N_1176,N_1788);
nand U5478 (N_5478,N_2555,N_1990);
or U5479 (N_5479,N_4755,N_799);
nand U5480 (N_5480,N_122,N_1586);
and U5481 (N_5481,N_495,N_465);
and U5482 (N_5482,N_2776,N_3971);
nor U5483 (N_5483,N_3901,N_1342);
xor U5484 (N_5484,N_1566,N_468);
nand U5485 (N_5485,N_3545,N_3843);
and U5486 (N_5486,N_3147,N_4788);
nor U5487 (N_5487,N_1211,N_222);
and U5488 (N_5488,N_3230,N_501);
xnor U5489 (N_5489,N_1170,N_3979);
and U5490 (N_5490,N_2689,N_1634);
or U5491 (N_5491,N_2606,N_2274);
or U5492 (N_5492,N_2210,N_1291);
nor U5493 (N_5493,N_2946,N_4614);
nor U5494 (N_5494,N_1698,N_2258);
nand U5495 (N_5495,N_3827,N_3000);
nor U5496 (N_5496,N_3412,N_1811);
nand U5497 (N_5497,N_1598,N_3204);
or U5498 (N_5498,N_3241,N_4417);
nor U5499 (N_5499,N_1524,N_4643);
nor U5500 (N_5500,N_9,N_1133);
and U5501 (N_5501,N_4781,N_3994);
nor U5502 (N_5502,N_3497,N_3162);
or U5503 (N_5503,N_4232,N_3836);
nor U5504 (N_5504,N_1485,N_3048);
and U5505 (N_5505,N_2141,N_3960);
nor U5506 (N_5506,N_2735,N_124);
or U5507 (N_5507,N_4258,N_3757);
nand U5508 (N_5508,N_2446,N_244);
nand U5509 (N_5509,N_4218,N_706);
and U5510 (N_5510,N_1613,N_546);
nor U5511 (N_5511,N_3915,N_3894);
or U5512 (N_5512,N_105,N_1689);
or U5513 (N_5513,N_3417,N_2104);
and U5514 (N_5514,N_776,N_948);
nor U5515 (N_5515,N_3773,N_2997);
and U5516 (N_5516,N_3434,N_3314);
nor U5517 (N_5517,N_733,N_1549);
xor U5518 (N_5518,N_3679,N_1963);
xnor U5519 (N_5519,N_1341,N_4538);
nor U5520 (N_5520,N_1887,N_3728);
nor U5521 (N_5521,N_4822,N_4412);
nand U5522 (N_5522,N_1873,N_4277);
nand U5523 (N_5523,N_4835,N_4917);
and U5524 (N_5524,N_1260,N_3213);
nand U5525 (N_5525,N_906,N_3181);
or U5526 (N_5526,N_2205,N_2387);
or U5527 (N_5527,N_3116,N_1619);
nand U5528 (N_5528,N_4471,N_3879);
nand U5529 (N_5529,N_1635,N_1821);
and U5530 (N_5530,N_4237,N_1166);
nor U5531 (N_5531,N_1294,N_663);
xnor U5532 (N_5532,N_3495,N_879);
or U5533 (N_5533,N_2060,N_87);
nand U5534 (N_5534,N_1226,N_3135);
or U5535 (N_5535,N_2292,N_889);
nand U5536 (N_5536,N_1006,N_4115);
and U5537 (N_5537,N_2390,N_4686);
nor U5538 (N_5538,N_2027,N_446);
nand U5539 (N_5539,N_1466,N_2266);
nand U5540 (N_5540,N_1544,N_1014);
nor U5541 (N_5541,N_1356,N_1209);
nand U5542 (N_5542,N_3712,N_4630);
and U5543 (N_5543,N_2886,N_267);
or U5544 (N_5544,N_2157,N_3799);
nor U5545 (N_5545,N_1484,N_140);
nor U5546 (N_5546,N_474,N_162);
nor U5547 (N_5547,N_285,N_3423);
or U5548 (N_5548,N_872,N_53);
nand U5549 (N_5549,N_77,N_1892);
nor U5550 (N_5550,N_2515,N_1932);
nor U5551 (N_5551,N_1407,N_3310);
nand U5552 (N_5552,N_892,N_4247);
nor U5553 (N_5553,N_4494,N_2733);
nor U5554 (N_5554,N_4829,N_1464);
nand U5555 (N_5555,N_2159,N_400);
or U5556 (N_5556,N_2149,N_4100);
xor U5557 (N_5557,N_224,N_2288);
nand U5558 (N_5558,N_3481,N_1905);
nand U5559 (N_5559,N_2329,N_4379);
xnor U5560 (N_5560,N_4525,N_1405);
and U5561 (N_5561,N_349,N_4129);
nor U5562 (N_5562,N_1989,N_2719);
xor U5563 (N_5563,N_1107,N_2429);
and U5564 (N_5564,N_4332,N_4687);
or U5565 (N_5565,N_2826,N_515);
nand U5566 (N_5566,N_3049,N_1205);
nor U5567 (N_5567,N_850,N_598);
xor U5568 (N_5568,N_3206,N_4505);
and U5569 (N_5569,N_3720,N_3282);
or U5570 (N_5570,N_2003,N_1919);
and U5571 (N_5571,N_4661,N_557);
and U5572 (N_5572,N_3126,N_3519);
and U5573 (N_5573,N_3218,N_3375);
nor U5574 (N_5574,N_345,N_2066);
and U5575 (N_5575,N_1591,N_4934);
or U5576 (N_5576,N_966,N_3108);
nand U5577 (N_5577,N_710,N_2123);
nand U5578 (N_5578,N_2581,N_3526);
and U5579 (N_5579,N_3520,N_3201);
or U5580 (N_5580,N_2634,N_1859);
nor U5581 (N_5581,N_714,N_3535);
nand U5582 (N_5582,N_4191,N_2917);
nor U5583 (N_5583,N_4616,N_541);
nand U5584 (N_5584,N_3930,N_120);
and U5585 (N_5585,N_2102,N_699);
xnor U5586 (N_5586,N_2863,N_960);
or U5587 (N_5587,N_1127,N_4574);
and U5588 (N_5588,N_553,N_4172);
nand U5589 (N_5589,N_577,N_3077);
nor U5590 (N_5590,N_1225,N_292);
or U5591 (N_5591,N_3266,N_2942);
nand U5592 (N_5592,N_4544,N_2710);
and U5593 (N_5593,N_2070,N_2611);
nand U5594 (N_5594,N_303,N_2976);
and U5595 (N_5595,N_3611,N_1787);
or U5596 (N_5596,N_809,N_1931);
and U5597 (N_5597,N_4193,N_484);
or U5598 (N_5598,N_3438,N_1954);
or U5599 (N_5599,N_619,N_2843);
nand U5600 (N_5600,N_2952,N_3297);
nand U5601 (N_5601,N_4672,N_914);
and U5602 (N_5602,N_502,N_3708);
or U5603 (N_5603,N_4068,N_4509);
nor U5604 (N_5604,N_4104,N_3278);
nor U5605 (N_5605,N_3070,N_369);
nor U5606 (N_5606,N_926,N_3430);
and U5607 (N_5607,N_977,N_1128);
and U5608 (N_5608,N_3531,N_74);
xor U5609 (N_5609,N_3958,N_386);
nand U5610 (N_5610,N_2518,N_4931);
nand U5611 (N_5611,N_672,N_4138);
nand U5612 (N_5612,N_1490,N_1578);
nand U5613 (N_5613,N_2491,N_4927);
and U5614 (N_5614,N_1902,N_4181);
and U5615 (N_5615,N_2871,N_399);
nor U5616 (N_5616,N_4592,N_4673);
nor U5617 (N_5617,N_1147,N_2239);
nand U5618 (N_5618,N_4044,N_3575);
or U5619 (N_5619,N_1630,N_4408);
nor U5620 (N_5620,N_4711,N_4302);
and U5621 (N_5621,N_3865,N_590);
and U5622 (N_5622,N_2989,N_4815);
or U5623 (N_5623,N_770,N_4027);
and U5624 (N_5624,N_228,N_2540);
xnor U5625 (N_5625,N_3312,N_1866);
nand U5626 (N_5626,N_2615,N_1189);
nor U5627 (N_5627,N_4067,N_4797);
nand U5628 (N_5628,N_3850,N_2693);
nand U5629 (N_5629,N_3658,N_4376);
or U5630 (N_5630,N_123,N_998);
and U5631 (N_5631,N_3052,N_2333);
or U5632 (N_5632,N_1151,N_3887);
nand U5633 (N_5633,N_1839,N_2261);
nand U5634 (N_5634,N_1636,N_2428);
and U5635 (N_5635,N_4366,N_4201);
and U5636 (N_5636,N_4128,N_3946);
nand U5637 (N_5637,N_1550,N_1841);
nand U5638 (N_5638,N_2228,N_3233);
nand U5639 (N_5639,N_1637,N_1340);
nor U5640 (N_5640,N_2322,N_1953);
nor U5641 (N_5641,N_1140,N_135);
and U5642 (N_5642,N_193,N_2630);
or U5643 (N_5643,N_4793,N_278);
nand U5644 (N_5644,N_840,N_1358);
or U5645 (N_5645,N_1665,N_913);
or U5646 (N_5646,N_2590,N_1007);
or U5647 (N_5647,N_4448,N_1242);
or U5648 (N_5648,N_4875,N_3884);
and U5649 (N_5649,N_2472,N_1838);
or U5650 (N_5650,N_1601,N_3054);
and U5651 (N_5651,N_3293,N_2636);
or U5652 (N_5652,N_437,N_2564);
and U5653 (N_5653,N_2498,N_1957);
or U5654 (N_5654,N_3004,N_121);
nand U5655 (N_5655,N_3837,N_723);
or U5656 (N_5656,N_4188,N_2043);
nand U5657 (N_5657,N_784,N_2016);
or U5658 (N_5658,N_3212,N_3401);
nand U5659 (N_5659,N_562,N_1460);
nand U5660 (N_5660,N_2132,N_4691);
or U5661 (N_5661,N_1456,N_3355);
xnor U5662 (N_5662,N_2341,N_2456);
or U5663 (N_5663,N_4817,N_1326);
and U5664 (N_5664,N_25,N_4135);
and U5665 (N_5665,N_1683,N_2547);
nor U5666 (N_5666,N_2539,N_2200);
or U5667 (N_5667,N_2867,N_2276);
xnor U5668 (N_5668,N_787,N_550);
nor U5669 (N_5669,N_287,N_3831);
or U5670 (N_5670,N_3498,N_658);
xnor U5671 (N_5671,N_4701,N_1066);
nor U5672 (N_5672,N_1781,N_4349);
nand U5673 (N_5673,N_301,N_3299);
nor U5674 (N_5674,N_4437,N_4254);
or U5675 (N_5675,N_1267,N_1528);
or U5676 (N_5676,N_1678,N_3486);
and U5677 (N_5677,N_4368,N_1338);
or U5678 (N_5678,N_2046,N_4893);
or U5679 (N_5679,N_2895,N_4632);
or U5680 (N_5680,N_707,N_321);
nand U5681 (N_5681,N_2972,N_2915);
nand U5682 (N_5682,N_212,N_4863);
nand U5683 (N_5683,N_48,N_4308);
nand U5684 (N_5684,N_1981,N_3555);
and U5685 (N_5685,N_177,N_667);
and U5686 (N_5686,N_3389,N_4132);
and U5687 (N_5687,N_1235,N_2129);
xor U5688 (N_5688,N_941,N_4591);
nand U5689 (N_5689,N_315,N_82);
and U5690 (N_5690,N_3368,N_4359);
or U5691 (N_5691,N_251,N_911);
and U5692 (N_5692,N_1302,N_1986);
and U5693 (N_5693,N_2714,N_565);
nand U5694 (N_5694,N_2505,N_4045);
and U5695 (N_5695,N_2344,N_4469);
nor U5696 (N_5696,N_461,N_3889);
and U5697 (N_5697,N_3985,N_3449);
nand U5698 (N_5698,N_2612,N_4848);
or U5699 (N_5699,N_2980,N_3478);
and U5700 (N_5700,N_3539,N_180);
nand U5701 (N_5701,N_2511,N_3990);
and U5702 (N_5702,N_1876,N_2965);
or U5703 (N_5703,N_273,N_3542);
xor U5704 (N_5704,N_3473,N_3648);
and U5705 (N_5705,N_2944,N_2069);
and U5706 (N_5706,N_1780,N_467);
and U5707 (N_5707,N_499,N_1116);
or U5708 (N_5708,N_972,N_4377);
or U5709 (N_5709,N_4016,N_3079);
or U5710 (N_5710,N_1991,N_245);
nor U5711 (N_5711,N_2734,N_2306);
and U5712 (N_5712,N_4943,N_676);
nand U5713 (N_5713,N_715,N_3921);
or U5714 (N_5714,N_4597,N_3582);
and U5715 (N_5715,N_1198,N_826);
nand U5716 (N_5716,N_174,N_4329);
nor U5717 (N_5717,N_383,N_1251);
nor U5718 (N_5718,N_1988,N_2202);
or U5719 (N_5719,N_3788,N_1701);
nor U5720 (N_5720,N_3224,N_3465);
and U5721 (N_5721,N_1835,N_4195);
nor U5722 (N_5722,N_3674,N_1451);
nand U5723 (N_5723,N_2787,N_3875);
or U5724 (N_5724,N_3186,N_2692);
nand U5725 (N_5725,N_4117,N_2289);
or U5726 (N_5726,N_3910,N_3717);
xnor U5727 (N_5727,N_781,N_2510);
and U5728 (N_5728,N_3577,N_2940);
or U5729 (N_5729,N_1429,N_1433);
and U5730 (N_5730,N_4873,N_3075);
xor U5731 (N_5731,N_3663,N_3341);
or U5732 (N_5732,N_2407,N_1575);
nor U5733 (N_5733,N_2185,N_3394);
nor U5734 (N_5734,N_4720,N_1109);
nor U5735 (N_5735,N_4272,N_1398);
and U5736 (N_5736,N_1469,N_351);
nand U5737 (N_5737,N_4020,N_3538);
and U5738 (N_5738,N_2309,N_4387);
and U5739 (N_5739,N_1048,N_3846);
nand U5740 (N_5740,N_1252,N_3900);
and U5741 (N_5741,N_1309,N_698);
and U5742 (N_5742,N_555,N_211);
nor U5743 (N_5743,N_2452,N_3090);
nand U5744 (N_5744,N_1319,N_2382);
nor U5745 (N_5745,N_4183,N_237);
nand U5746 (N_5746,N_1737,N_3780);
and U5747 (N_5747,N_1516,N_4190);
nand U5748 (N_5748,N_3494,N_2908);
nand U5749 (N_5749,N_2956,N_62);
nand U5750 (N_5750,N_2115,N_71);
and U5751 (N_5751,N_1221,N_20);
nand U5752 (N_5752,N_2038,N_2829);
or U5753 (N_5753,N_2315,N_168);
or U5754 (N_5754,N_3482,N_3558);
or U5755 (N_5755,N_1360,N_4842);
or U5756 (N_5756,N_3179,N_404);
nand U5757 (N_5757,N_3257,N_1305);
nor U5758 (N_5758,N_2973,N_3376);
or U5759 (N_5759,N_3053,N_1632);
nand U5760 (N_5760,N_4360,N_2062);
xnor U5761 (N_5761,N_1438,N_3697);
xnor U5762 (N_5762,N_2323,N_1750);
and U5763 (N_5763,N_4155,N_4304);
nor U5764 (N_5764,N_797,N_2823);
or U5765 (N_5765,N_380,N_3832);
nand U5766 (N_5766,N_1807,N_2941);
nor U5767 (N_5767,N_570,N_3630);
and U5768 (N_5768,N_4603,N_3228);
nand U5769 (N_5769,N_1646,N_2475);
xor U5770 (N_5770,N_160,N_3184);
nor U5771 (N_5771,N_1542,N_1304);
nand U5772 (N_5772,N_4753,N_4532);
and U5773 (N_5773,N_1349,N_3318);
and U5774 (N_5774,N_712,N_4019);
nor U5775 (N_5775,N_12,N_463);
xnor U5776 (N_5776,N_388,N_2334);
xnor U5777 (N_5777,N_265,N_1942);
and U5778 (N_5778,N_4140,N_1212);
nand U5779 (N_5779,N_415,N_364);
and U5780 (N_5780,N_2893,N_3922);
nor U5781 (N_5781,N_4335,N_564);
xor U5782 (N_5782,N_4836,N_156);
nand U5783 (N_5783,N_1531,N_739);
or U5784 (N_5784,N_4565,N_1741);
nand U5785 (N_5785,N_1594,N_3258);
nand U5786 (N_5786,N_3039,N_2698);
nor U5787 (N_5787,N_3154,N_2875);
nand U5788 (N_5788,N_4287,N_3022);
nand U5789 (N_5789,N_2681,N_4883);
or U5790 (N_5790,N_275,N_3007);
and U5791 (N_5791,N_3964,N_2576);
nand U5792 (N_5792,N_2313,N_750);
nand U5793 (N_5793,N_832,N_3011);
and U5794 (N_5794,N_2166,N_3634);
nor U5795 (N_5795,N_2358,N_4355);
xor U5796 (N_5796,N_2328,N_3466);
xnor U5797 (N_5797,N_3325,N_3772);
nand U5798 (N_5798,N_4033,N_1826);
and U5799 (N_5799,N_1790,N_2450);
nand U5800 (N_5800,N_339,N_1434);
nand U5801 (N_5801,N_137,N_1266);
or U5802 (N_5802,N_4991,N_2250);
and U5803 (N_5803,N_3557,N_4758);
or U5804 (N_5804,N_2912,N_78);
nor U5805 (N_5805,N_4877,N_3952);
nor U5806 (N_5806,N_3180,N_2326);
nand U5807 (N_5807,N_1657,N_689);
xor U5808 (N_5808,N_1473,N_1660);
and U5809 (N_5809,N_4358,N_2487);
or U5810 (N_5810,N_4625,N_2213);
xnor U5811 (N_5811,N_4280,N_184);
and U5812 (N_5812,N_1263,N_4105);
or U5813 (N_5813,N_3819,N_4581);
nand U5814 (N_5814,N_439,N_4515);
nand U5815 (N_5815,N_1554,N_2772);
nand U5816 (N_5816,N_3504,N_4894);
or U5817 (N_5817,N_1943,N_2214);
nand U5818 (N_5818,N_2300,N_1068);
or U5819 (N_5819,N_3839,N_4834);
or U5820 (N_5820,N_2656,N_482);
nand U5821 (N_5821,N_2197,N_3149);
nor U5822 (N_5822,N_753,N_2260);
and U5823 (N_5823,N_4406,N_92);
and U5824 (N_5824,N_1020,N_4413);
nand U5825 (N_5825,N_4770,N_3676);
and U5826 (N_5826,N_2523,N_2217);
or U5827 (N_5827,N_3406,N_1852);
and U5828 (N_5828,N_3109,N_1815);
and U5829 (N_5829,N_2156,N_1453);
nor U5830 (N_5830,N_4654,N_1502);
nand U5831 (N_5831,N_2669,N_1256);
and U5832 (N_5832,N_2142,N_3174);
nand U5833 (N_5833,N_803,N_874);
nor U5834 (N_5834,N_2140,N_1367);
nor U5835 (N_5835,N_4801,N_606);
nand U5836 (N_5836,N_1069,N_3369);
nand U5837 (N_5837,N_2675,N_3777);
or U5838 (N_5838,N_2660,N_2405);
or U5839 (N_5839,N_1709,N_4840);
nand U5840 (N_5840,N_3919,N_752);
or U5841 (N_5841,N_1273,N_2308);
nor U5842 (N_5842,N_921,N_2488);
nor U5843 (N_5843,N_2774,N_4297);
nor U5844 (N_5844,N_1579,N_196);
xnor U5845 (N_5845,N_1547,N_801);
nor U5846 (N_5846,N_1171,N_677);
nand U5847 (N_5847,N_3956,N_4818);
or U5848 (N_5848,N_2432,N_725);
and U5849 (N_5849,N_4161,N_1468);
and U5850 (N_5850,N_2812,N_4111);
or U5851 (N_5851,N_2373,N_3238);
nand U5852 (N_5852,N_4539,N_1923);
or U5853 (N_5853,N_3779,N_1901);
xor U5854 (N_5854,N_2109,N_870);
or U5855 (N_5855,N_3975,N_3148);
nor U5856 (N_5856,N_1650,N_2771);
nand U5857 (N_5857,N_1801,N_4526);
or U5858 (N_5858,N_3657,N_1377);
nand U5859 (N_5859,N_3886,N_22);
nand U5860 (N_5860,N_1246,N_4443);
nand U5861 (N_5861,N_28,N_2054);
and U5862 (N_5862,N_4056,N_4750);
and U5863 (N_5863,N_788,N_838);
or U5864 (N_5864,N_4365,N_3874);
or U5865 (N_5865,N_1324,N_3151);
and U5866 (N_5866,N_4165,N_4839);
nor U5867 (N_5867,N_4986,N_2000);
nor U5868 (N_5868,N_665,N_3787);
or U5869 (N_5869,N_2847,N_298);
nor U5870 (N_5870,N_2125,N_4914);
nor U5871 (N_5871,N_4334,N_4757);
nor U5872 (N_5872,N_4920,N_3737);
xor U5873 (N_5873,N_2354,N_4321);
or U5874 (N_5874,N_4336,N_1029);
nor U5875 (N_5875,N_4464,N_3954);
xor U5876 (N_5876,N_2172,N_1498);
nor U5877 (N_5877,N_930,N_1207);
and U5878 (N_5878,N_3042,N_3584);
and U5879 (N_5879,N_4926,N_3693);
nor U5880 (N_5880,N_2809,N_1311);
nor U5881 (N_5881,N_4751,N_4210);
and U5882 (N_5882,N_450,N_4420);
and U5883 (N_5883,N_3269,N_587);
nor U5884 (N_5884,N_1402,N_3165);
and U5885 (N_5885,N_3322,N_357);
and U5886 (N_5886,N_1681,N_610);
xor U5887 (N_5887,N_2359,N_3289);
or U5888 (N_5888,N_2224,N_1157);
nor U5889 (N_5889,N_1538,N_3870);
nand U5890 (N_5890,N_3157,N_695);
nand U5891 (N_5891,N_2920,N_4895);
nand U5892 (N_5892,N_295,N_3940);
or U5893 (N_5893,N_361,N_4496);
or U5894 (N_5894,N_3856,N_3010);
or U5895 (N_5895,N_4452,N_1614);
or U5896 (N_5896,N_574,N_4003);
nor U5897 (N_5897,N_4179,N_2281);
xor U5898 (N_5898,N_2743,N_2119);
and U5899 (N_5899,N_2440,N_2434);
or U5900 (N_5900,N_1760,N_1149);
nor U5901 (N_5901,N_810,N_4960);
nand U5902 (N_5902,N_4421,N_2835);
and U5903 (N_5903,N_2543,N_1938);
or U5904 (N_5904,N_3420,N_1763);
or U5905 (N_5905,N_2777,N_2853);
nor U5906 (N_5906,N_927,N_1076);
nand U5907 (N_5907,N_2807,N_4865);
and U5908 (N_5908,N_3521,N_599);
nand U5909 (N_5909,N_4854,N_2659);
and U5910 (N_5910,N_1722,N_3970);
xnor U5911 (N_5911,N_3682,N_3609);
nand U5912 (N_5912,N_3384,N_1543);
nor U5913 (N_5913,N_90,N_2593);
nand U5914 (N_5914,N_2262,N_2520);
xnor U5915 (N_5915,N_932,N_3859);
nor U5916 (N_5916,N_547,N_1676);
xnor U5917 (N_5917,N_4617,N_3511);
nand U5918 (N_5918,N_143,N_4388);
xnor U5919 (N_5919,N_3034,N_2900);
or U5920 (N_5920,N_2087,N_4670);
nand U5921 (N_5921,N_2460,N_4969);
or U5922 (N_5922,N_2165,N_3422);
or U5923 (N_5923,N_4048,N_4998);
nand U5924 (N_5924,N_4492,N_2481);
and U5925 (N_5925,N_4095,N_4431);
nor U5926 (N_5926,N_94,N_1282);
and U5927 (N_5927,N_1056,N_213);
nor U5928 (N_5928,N_4118,N_3453);
nand U5929 (N_5929,N_1102,N_3854);
nand U5930 (N_5930,N_4189,N_1073);
or U5931 (N_5931,N_1734,N_3470);
or U5932 (N_5932,N_559,N_4487);
or U5933 (N_5933,N_645,N_4830);
nand U5934 (N_5934,N_2748,N_4322);
or U5935 (N_5935,N_2436,N_4283);
or U5936 (N_5936,N_4543,N_1909);
nor U5937 (N_5937,N_1927,N_2798);
or U5938 (N_5938,N_470,N_4903);
nand U5939 (N_5939,N_648,N_86);
nor U5940 (N_5940,N_2793,N_3029);
xor U5941 (N_5941,N_4708,N_1774);
nor U5942 (N_5942,N_37,N_4262);
nor U5943 (N_5943,N_178,N_1248);
nor U5944 (N_5944,N_3158,N_2499);
or U5945 (N_5945,N_4197,N_694);
and U5946 (N_5946,N_2722,N_2578);
and U5947 (N_5947,N_1228,N_617);
or U5948 (N_5948,N_4785,N_4204);
and U5949 (N_5949,N_327,N_945);
and U5950 (N_5950,N_4729,N_3429);
or U5951 (N_5951,N_424,N_4791);
and U5952 (N_5952,N_1329,N_157);
nor U5953 (N_5953,N_4046,N_2736);
nor U5954 (N_5954,N_1627,N_792);
or U5955 (N_5955,N_3986,N_1893);
and U5956 (N_5956,N_2226,N_3586);
xor U5957 (N_5957,N_2012,N_4461);
and U5958 (N_5958,N_4808,N_3579);
nand U5959 (N_5959,N_449,N_2321);
and U5960 (N_5960,N_2042,N_358);
xor U5961 (N_5961,N_1924,N_317);
nand U5962 (N_5962,N_3050,N_3008);
and U5963 (N_5963,N_4924,N_4162);
nor U5964 (N_5964,N_4915,N_4363);
or U5965 (N_5965,N_2061,N_864);
and U5966 (N_5966,N_4049,N_834);
nand U5967 (N_5967,N_2246,N_3911);
or U5968 (N_5968,N_4954,N_1415);
xnor U5969 (N_5969,N_269,N_1977);
nand U5970 (N_5970,N_4600,N_247);
nor U5971 (N_5971,N_1570,N_3176);
or U5972 (N_5972,N_4110,N_190);
xnor U5973 (N_5973,N_4939,N_4000);
xor U5974 (N_5974,N_2839,N_1672);
or U5975 (N_5975,N_3214,N_1705);
or U5976 (N_5976,N_2454,N_2484);
or U5977 (N_5977,N_4252,N_2780);
or U5978 (N_5978,N_1738,N_4514);
xor U5979 (N_5979,N_4288,N_4009);
or U5980 (N_5980,N_3484,N_4010);
or U5981 (N_5981,N_2804,N_3670);
and U5982 (N_5982,N_1571,N_3192);
xnor U5983 (N_5983,N_579,N_2684);
or U5984 (N_5984,N_131,N_1911);
and U5985 (N_5985,N_1160,N_4916);
nor U5986 (N_5986,N_2852,N_3327);
xnor U5987 (N_5987,N_3347,N_1512);
or U5988 (N_5988,N_3552,N_908);
and U5989 (N_5989,N_1998,N_3085);
xnor U5990 (N_5990,N_2230,N_1896);
nand U5991 (N_5991,N_4216,N_158);
nor U5992 (N_5992,N_4482,N_3222);
or U5993 (N_5993,N_3345,N_859);
nand U5994 (N_5994,N_4072,N_4820);
nand U5995 (N_5995,N_1716,N_1295);
nor U5996 (N_5996,N_2996,N_4457);
and U5997 (N_5997,N_634,N_2169);
nor U5998 (N_5998,N_4882,N_3883);
nand U5999 (N_5999,N_353,N_627);
nand U6000 (N_6000,N_1103,N_3600);
and U6001 (N_6001,N_3374,N_2676);
or U6002 (N_6002,N_3125,N_3568);
nor U6003 (N_6003,N_558,N_3066);
nor U6004 (N_6004,N_3063,N_1803);
or U6005 (N_6005,N_1978,N_347);
or U6006 (N_6006,N_4608,N_3237);
nor U6007 (N_6007,N_4381,N_4311);
and U6008 (N_6008,N_1843,N_4912);
or U6009 (N_6009,N_4192,N_4679);
nand U6010 (N_6010,N_4474,N_918);
and U6011 (N_6011,N_3691,N_4362);
nor U6012 (N_6012,N_1752,N_3506);
and U6013 (N_6013,N_2255,N_4768);
nand U6014 (N_6014,N_4541,N_593);
nor U6015 (N_6015,N_1658,N_226);
nor U6016 (N_6016,N_2483,N_3030);
nand U6017 (N_6017,N_2810,N_2951);
xor U6018 (N_6018,N_1230,N_2654);
nor U6019 (N_6019,N_1009,N_3418);
nor U6020 (N_6020,N_4635,N_473);
nand U6021 (N_6021,N_923,N_4227);
nor U6022 (N_6022,N_2859,N_3544);
and U6023 (N_6023,N_1751,N_2744);
nand U6024 (N_6024,N_582,N_4032);
xor U6025 (N_6025,N_1783,N_2178);
nand U6026 (N_6026,N_2975,N_4628);
and U6027 (N_6027,N_3516,N_2567);
nand U6028 (N_6028,N_4966,N_1045);
nand U6029 (N_6029,N_311,N_1849);
or U6030 (N_6030,N_3267,N_2961);
xor U6031 (N_6031,N_3072,N_3277);
nand U6032 (N_6032,N_1131,N_778);
and U6033 (N_6033,N_4658,N_4542);
and U6034 (N_6034,N_3379,N_1710);
or U6035 (N_6035,N_3594,N_4739);
or U6036 (N_6036,N_2604,N_3767);
nand U6037 (N_6037,N_1638,N_1888);
xnor U6038 (N_6038,N_2122,N_4352);
nor U6039 (N_6039,N_2775,N_571);
nand U6040 (N_6040,N_64,N_1631);
and U6041 (N_6041,N_2399,N_3972);
nor U6042 (N_6042,N_2098,N_453);
or U6043 (N_6043,N_4740,N_3256);
and U6044 (N_6044,N_4325,N_4714);
nand U6045 (N_6045,N_931,N_402);
nand U6046 (N_6046,N_4236,N_4106);
and U6047 (N_6047,N_99,N_4051);
or U6048 (N_6048,N_3661,N_1089);
nand U6049 (N_6049,N_794,N_1917);
and U6050 (N_6050,N_2401,N_620);
nor U6051 (N_6051,N_851,N_900);
nor U6052 (N_6052,N_961,N_4585);
xor U6053 (N_6053,N_2556,N_1846);
and U6054 (N_6054,N_1191,N_4184);
nor U6055 (N_6055,N_4733,N_4812);
nor U6056 (N_6056,N_3311,N_2705);
and U6057 (N_6057,N_2833,N_4948);
and U6058 (N_6058,N_4995,N_3709);
xor U6059 (N_6059,N_1159,N_1332);
xnor U6060 (N_6060,N_4599,N_3771);
nor U6061 (N_6061,N_4816,N_3407);
nor U6062 (N_6062,N_2560,N_4847);
or U6063 (N_6063,N_3793,N_1860);
nand U6064 (N_6064,N_3460,N_1241);
and U6065 (N_6065,N_4198,N_1656);
and U6066 (N_6066,N_1507,N_481);
nand U6067 (N_6067,N_4449,N_1334);
nand U6068 (N_6068,N_819,N_2671);
nor U6069 (N_6069,N_2904,N_3501);
nand U6070 (N_6070,N_3300,N_2296);
or U6071 (N_6071,N_2694,N_2834);
nand U6072 (N_6072,N_1569,N_4680);
nand U6073 (N_6073,N_3744,N_3635);
or U6074 (N_6074,N_1345,N_3776);
and U6075 (N_6075,N_2795,N_4685);
xor U6076 (N_6076,N_3413,N_2116);
and U6077 (N_6077,N_653,N_1933);
and U6078 (N_6078,N_5,N_2836);
and U6079 (N_6079,N_3107,N_2767);
and U6080 (N_6080,N_1025,N_4062);
or U6081 (N_6081,N_3031,N_2967);
nand U6082 (N_6082,N_4235,N_4558);
xor U6083 (N_6083,N_4241,N_3139);
nand U6084 (N_6084,N_4400,N_4577);
nor U6085 (N_6085,N_3515,N_2781);
xor U6086 (N_6086,N_394,N_420);
nor U6087 (N_6087,N_1313,N_3261);
xor U6088 (N_6088,N_3731,N_1879);
or U6089 (N_6089,N_1675,N_205);
nand U6090 (N_6090,N_1670,N_3597);
nor U6091 (N_6091,N_2236,N_4416);
or U6092 (N_6092,N_2998,N_3183);
nand U6093 (N_6093,N_1031,N_2759);
nand U6094 (N_6094,N_1728,N_1017);
nor U6095 (N_6095,N_4901,N_3505);
and U6096 (N_6096,N_242,N_4664);
nor U6097 (N_6097,N_3440,N_4869);
nor U6098 (N_6098,N_4442,N_322);
nand U6099 (N_6099,N_2008,N_173);
and U6100 (N_6100,N_1855,N_2376);
nand U6101 (N_6101,N_3722,N_3902);
nor U6102 (N_6102,N_949,N_2500);
or U6103 (N_6103,N_3234,N_3748);
nor U6104 (N_6104,N_3816,N_1830);
and U6105 (N_6105,N_4919,N_4741);
nor U6106 (N_6106,N_316,N_1);
or U6107 (N_6107,N_657,N_3489);
nor U6108 (N_6108,N_3920,N_4476);
nor U6109 (N_6109,N_1435,N_4245);
nand U6110 (N_6110,N_3123,N_679);
nand U6111 (N_6111,N_3618,N_1150);
or U6112 (N_6112,N_4107,N_1508);
nor U6113 (N_6113,N_350,N_2786);
and U6114 (N_6114,N_443,N_1387);
nor U6115 (N_6115,N_3512,N_877);
and U6116 (N_6116,N_567,N_655);
or U6117 (N_6117,N_1604,N_3500);
xnor U6118 (N_6118,N_3583,N_3939);
nor U6119 (N_6119,N_2055,N_1202);
xor U6120 (N_6120,N_3292,N_3955);
nand U6121 (N_6121,N_3,N_3932);
and U6122 (N_6122,N_1975,N_4176);
nand U6123 (N_6123,N_629,N_1844);
xnor U6124 (N_6124,N_1378,N_2077);
or U6125 (N_6125,N_2295,N_1925);
nor U6126 (N_6126,N_3677,N_4959);
xnor U6127 (N_6127,N_868,N_1509);
and U6128 (N_6128,N_4345,N_1640);
nand U6129 (N_6129,N_2649,N_862);
and U6130 (N_6130,N_2551,N_2489);
nand U6131 (N_6131,N_4174,N_1736);
or U6132 (N_6132,N_256,N_3065);
nand U6133 (N_6133,N_1834,N_1143);
nand U6134 (N_6134,N_4696,N_4278);
nand U6135 (N_6135,N_2791,N_2717);
nand U6136 (N_6136,N_818,N_1551);
xnor U6137 (N_6137,N_1900,N_589);
nor U6138 (N_6138,N_863,N_1086);
nor U6139 (N_6139,N_1339,N_2019);
and U6140 (N_6140,N_1677,N_3200);
nand U6141 (N_6141,N_777,N_1104);
and U6142 (N_6142,N_2848,N_4596);
nand U6143 (N_6143,N_1987,N_4395);
nand U6144 (N_6144,N_1070,N_2298);
or U6145 (N_6145,N_323,N_4166);
nand U6146 (N_6146,N_1836,N_2286);
or U6147 (N_6147,N_4737,N_4962);
or U6148 (N_6148,N_3254,N_4175);
nand U6149 (N_6149,N_487,N_365);
and U6150 (N_6150,N_128,N_3683);
nand U6151 (N_6151,N_255,N_4240);
and U6152 (N_6152,N_4678,N_141);
or U6153 (N_6153,N_531,N_626);
nand U6154 (N_6154,N_2468,N_3800);
or U6155 (N_6155,N_2959,N_3229);
nand U6156 (N_6156,N_1397,N_2415);
xnor U6157 (N_6157,N_4040,N_1403);
nand U6158 (N_6158,N_2921,N_4549);
nand U6159 (N_6159,N_3724,N_3769);
nand U6160 (N_6160,N_4314,N_3472);
or U6161 (N_6161,N_4131,N_1224);
nor U6162 (N_6162,N_3897,N_3802);
nand U6163 (N_6163,N_1837,N_979);
and U6164 (N_6164,N_4665,N_4083);
or U6165 (N_6165,N_93,N_4716);
or U6166 (N_6166,N_1659,N_4556);
nor U6167 (N_6167,N_2849,N_4951);
nand U6168 (N_6168,N_45,N_2049);
nor U6169 (N_6169,N_2755,N_1711);
xor U6170 (N_6170,N_2310,N_4438);
or U6171 (N_6171,N_4550,N_1450);
or U6172 (N_6172,N_2193,N_3113);
or U6173 (N_6173,N_1418,N_2662);
and U6174 (N_6174,N_3905,N_2433);
and U6175 (N_6175,N_2486,N_4606);
and U6176 (N_6176,N_2478,N_3673);
or U6177 (N_6177,N_3302,N_2340);
xor U6178 (N_6178,N_4029,N_2138);
or U6179 (N_6179,N_848,N_2091);
nand U6180 (N_6180,N_556,N_2291);
nand U6181 (N_6181,N_4907,N_4053);
and U6182 (N_6182,N_3765,N_2133);
or U6183 (N_6183,N_1426,N_4012);
and U6184 (N_6184,N_3337,N_290);
and U6185 (N_6185,N_2311,N_3209);
and U6186 (N_6186,N_903,N_3664);
nor U6187 (N_6187,N_1592,N_833);
nor U6188 (N_6188,N_2120,N_3323);
or U6189 (N_6189,N_4749,N_764);
and U6190 (N_6190,N_3055,N_203);
and U6191 (N_6191,N_3346,N_3537);
nand U6192 (N_6192,N_3442,N_1142);
nor U6193 (N_6193,N_3547,N_782);
xor U6194 (N_6194,N_1106,N_3796);
and U6195 (N_6195,N_3914,N_3899);
and U6196 (N_6196,N_2683,N_3196);
nand U6197 (N_6197,N_4667,N_4721);
or U6198 (N_6198,N_3319,N_2788);
nor U6199 (N_6199,N_4112,N_3906);
xor U6200 (N_6200,N_2423,N_4219);
nor U6201 (N_6201,N_3936,N_1343);
or U6202 (N_6202,N_3071,N_692);
and U6203 (N_6203,N_2237,N_3541);
and U6204 (N_6204,N_1470,N_569);
and U6205 (N_6205,N_4964,N_3860);
or U6206 (N_6206,N_1870,N_304);
and U6207 (N_6207,N_1522,N_3866);
and U6208 (N_6208,N_4108,N_1980);
nand U6209 (N_6209,N_3232,N_1596);
xnor U6210 (N_6210,N_2580,N_2651);
nor U6211 (N_6211,N_476,N_2194);
or U6212 (N_6212,N_856,N_821);
nand U6213 (N_6213,N_4410,N_1746);
xnor U6214 (N_6214,N_2469,N_248);
and U6215 (N_6215,N_4401,N_2131);
nor U6216 (N_6216,N_624,N_3549);
nand U6217 (N_6217,N_263,N_4536);
nand U6218 (N_6218,N_3961,N_4921);
or U6219 (N_6219,N_223,N_3018);
and U6220 (N_6220,N_2135,N_4760);
and U6221 (N_6221,N_469,N_343);
and U6222 (N_6222,N_4553,N_3733);
or U6223 (N_6223,N_4202,N_3742);
nor U6224 (N_6224,N_4985,N_2948);
nor U6225 (N_6225,N_2579,N_219);
and U6226 (N_6226,N_1192,N_3536);
and U6227 (N_6227,N_847,N_2154);
or U6228 (N_6228,N_4275,N_452);
or U6229 (N_6229,N_3645,N_3948);
nand U6230 (N_6230,N_2978,N_685);
or U6231 (N_6231,N_1949,N_2186);
nand U6232 (N_6232,N_4301,N_319);
and U6233 (N_6233,N_4656,N_601);
xor U6234 (N_6234,N_751,N_4339);
and U6235 (N_6235,N_3264,N_3931);
or U6236 (N_6236,N_3762,N_1372);
nor U6237 (N_6237,N_3380,N_34);
or U6238 (N_6238,N_3792,N_302);
and U6239 (N_6239,N_4134,N_30);
nand U6240 (N_6240,N_973,N_4979);
nor U6241 (N_6241,N_1206,N_1539);
nand U6242 (N_6242,N_828,N_4528);
and U6243 (N_6243,N_881,N_4870);
xor U6244 (N_6244,N_2035,N_271);
nand U6245 (N_6245,N_1261,N_3852);
and U6246 (N_6246,N_4584,N_2445);
or U6247 (N_6247,N_4640,N_762);
or U6248 (N_6248,N_164,N_3225);
nor U6249 (N_6249,N_1884,N_2130);
nand U6250 (N_6250,N_2444,N_2706);
nand U6251 (N_6251,N_2371,N_4028);
nor U6252 (N_6252,N_504,N_594);
and U6253 (N_6253,N_3912,N_2832);
nor U6254 (N_6254,N_1190,N_4689);
or U6255 (N_6255,N_1454,N_1386);
and U6256 (N_6256,N_1071,N_1568);
and U6257 (N_6257,N_1231,N_3270);
nor U6258 (N_6258,N_519,N_3983);
nor U6259 (N_6259,N_4462,N_4293);
nor U6260 (N_6260,N_686,N_4271);
or U6261 (N_6261,N_4975,N_458);
and U6262 (N_6262,N_2709,N_4639);
nor U6263 (N_6263,N_1633,N_1134);
nor U6264 (N_6264,N_1661,N_3120);
and U6265 (N_6265,N_4580,N_4315);
nand U6266 (N_6266,N_241,N_3578);
nand U6267 (N_6267,N_3164,N_2621);
or U6268 (N_6268,N_3463,N_111);
nor U6269 (N_6269,N_2534,N_4560);
and U6270 (N_6270,N_2565,N_1510);
and U6271 (N_6271,N_4582,N_2145);
nor U6272 (N_6272,N_2741,N_3187);
and U6273 (N_6273,N_1713,N_4399);
and U6274 (N_6274,N_2570,N_1805);
nor U6275 (N_6275,N_1155,N_4892);
or U6276 (N_6276,N_1091,N_186);
nand U6277 (N_6277,N_198,N_1871);
and U6278 (N_6278,N_61,N_1457);
xor U6279 (N_6279,N_1238,N_1180);
nor U6280 (N_6280,N_3774,N_3226);
nand U6281 (N_6281,N_4127,N_3021);
or U6282 (N_6282,N_2047,N_1851);
and U6283 (N_6283,N_4286,N_155);
nor U6284 (N_6284,N_1972,N_16);
nand U6285 (N_6285,N_3134,N_2402);
and U6286 (N_6286,N_448,N_4229);
nand U6287 (N_6287,N_2620,N_1654);
nor U6288 (N_6288,N_2244,N_312);
or U6289 (N_6289,N_209,N_3059);
or U6290 (N_6290,N_436,N_4180);
and U6291 (N_6291,N_4777,N_3734);
and U6292 (N_6292,N_2410,N_2254);
xor U6293 (N_6293,N_1015,N_766);
and U6294 (N_6294,N_3873,N_2760);
nand U6295 (N_6295,N_1478,N_3344);
nor U6296 (N_6296,N_1328,N_4465);
nor U6297 (N_6297,N_1117,N_3877);
and U6298 (N_6298,N_4036,N_1664);
xnor U6299 (N_6299,N_2589,N_855);
or U6300 (N_6300,N_3166,N_2635);
and U6301 (N_6301,N_3115,N_884);
nor U6302 (N_6302,N_4375,N_2598);
xor U6303 (N_6303,N_3485,N_4900);
nor U6304 (N_6304,N_3316,N_1629);
nand U6305 (N_6305,N_98,N_1052);
and U6306 (N_6306,N_823,N_732);
or U6307 (N_6307,N_3219,N_2128);
or U6308 (N_6308,N_4936,N_995);
and U6309 (N_6309,N_2721,N_1525);
nor U6310 (N_6310,N_3947,N_2100);
xor U6311 (N_6311,N_2057,N_1761);
nor U6312 (N_6312,N_4732,N_52);
or U6313 (N_6313,N_217,N_4459);
nor U6314 (N_6314,N_3426,N_1644);
and U6315 (N_6315,N_1314,N_1244);
or U6316 (N_6316,N_3475,N_3024);
and U6317 (N_6317,N_4341,N_167);
or U6318 (N_6318,N_4576,N_1482);
nand U6319 (N_6319,N_4326,N_207);
and U6320 (N_6320,N_2822,N_4194);
or U6321 (N_6321,N_1529,N_456);
xor U6322 (N_6322,N_4122,N_4655);
and U6323 (N_6323,N_127,N_2737);
nor U6324 (N_6324,N_7,N_2337);
and U6325 (N_6325,N_1312,N_1194);
nand U6326 (N_6326,N_3565,N_3721);
or U6327 (N_6327,N_514,N_2167);
or U6328 (N_6328,N_806,N_270);
and U6329 (N_6329,N_1323,N_3060);
nor U6330 (N_6330,N_4501,N_1427);
and U6331 (N_6331,N_4324,N_1831);
nand U6332 (N_6332,N_3383,N_4950);
nand U6333 (N_6333,N_3227,N_4248);
nand U6334 (N_6334,N_3356,N_1132);
and U6335 (N_6335,N_4922,N_2665);
nand U6336 (N_6336,N_729,N_2355);
or U6337 (N_6337,N_4776,N_4548);
or U6338 (N_6338,N_47,N_2688);
and U6339 (N_6339,N_3117,N_362);
nor U6340 (N_6340,N_4257,N_4309);
and U6341 (N_6341,N_374,N_940);
nand U6342 (N_6342,N_1258,N_1216);
nand U6343 (N_6343,N_1680,N_3786);
nand U6344 (N_6344,N_1245,N_1673);
and U6345 (N_6345,N_2448,N_2619);
or U6346 (N_6346,N_3530,N_4077);
nand U6347 (N_6347,N_1072,N_1948);
and U6348 (N_6348,N_3040,N_4637);
xnor U6349 (N_6349,N_523,N_1441);
nor U6350 (N_6350,N_2270,N_1417);
or U6351 (N_6351,N_1092,N_4586);
and U6352 (N_6352,N_2110,N_2303);
nor U6353 (N_6353,N_3763,N_2824);
or U6354 (N_6354,N_1276,N_2855);
and U6355 (N_6355,N_4918,N_1651);
and U6356 (N_6356,N_2427,N_2955);
nand U6357 (N_6357,N_4059,N_1057);
nand U6358 (N_6358,N_3824,N_3185);
xor U6359 (N_6359,N_1756,N_2463);
or U6360 (N_6360,N_431,N_1002);
or U6361 (N_6361,N_3798,N_2687);
and U6362 (N_6362,N_84,N_4980);
nor U6363 (N_6363,N_652,N_2085);
or U6364 (N_6364,N_2350,N_24);
nor U6365 (N_6365,N_2945,N_2962);
nand U6366 (N_6366,N_4047,N_2096);
nor U6367 (N_6367,N_2243,N_2443);
nor U6368 (N_6368,N_3245,N_2582);
or U6369 (N_6369,N_1842,N_2603);
xnor U6370 (N_6370,N_3534,N_200);
nand U6371 (N_6371,N_4238,N_1791);
and U6372 (N_6372,N_4660,N_4885);
or U6373 (N_6373,N_4618,N_1725);
or U6374 (N_6374,N_1546,N_4428);
and U6375 (N_6375,N_1269,N_107);
and U6376 (N_6376,N_4598,N_4242);
or U6377 (N_6377,N_1669,N_1306);
and U6378 (N_6378,N_2361,N_15);
and U6379 (N_6379,N_2800,N_3023);
nand U6380 (N_6380,N_89,N_2885);
and U6381 (N_6381,N_656,N_2966);
nand U6382 (N_6382,N_1255,N_10);
and U6383 (N_6383,N_1353,N_1620);
nand U6384 (N_6384,N_3488,N_2033);
and U6385 (N_6385,N_3396,N_2293);
xor U6386 (N_6386,N_4705,N_1745);
xor U6387 (N_6387,N_1704,N_3101);
nor U6388 (N_6388,N_187,N_145);
nand U6389 (N_6389,N_1753,N_2898);
nor U6390 (N_6390,N_2663,N_3822);
xor U6391 (N_6391,N_393,N_1005);
nor U6392 (N_6392,N_405,N_3804);
xnor U6393 (N_6393,N_1748,N_4677);
xnor U6394 (N_6394,N_1599,N_3477);
and U6395 (N_6395,N_412,N_1641);
nand U6396 (N_6396,N_524,N_1918);
and U6397 (N_6397,N_785,N_3159);
xnor U6398 (N_6398,N_992,N_1440);
nand U6399 (N_6399,N_2899,N_4225);
or U6400 (N_6400,N_4130,N_3454);
nand U6401 (N_6401,N_3009,N_3567);
xor U6402 (N_6402,N_68,N_4844);
nor U6403 (N_6403,N_2163,N_774);
nand U6404 (N_6404,N_3104,N_3999);
or U6405 (N_6405,N_4060,N_2245);
nor U6406 (N_6406,N_1984,N_4070);
nand U6407 (N_6407,N_4433,N_1779);
and U6408 (N_6408,N_1321,N_477);
and U6409 (N_6409,N_2493,N_1463);
and U6410 (N_6410,N_2220,N_1881);
nand U6411 (N_6411,N_3168,N_1693);
xor U6412 (N_6412,N_4987,N_2502);
or U6413 (N_6413,N_654,N_3476);
nand U6414 (N_6414,N_1777,N_3335);
nand U6415 (N_6415,N_814,N_639);
nand U6416 (N_6416,N_1097,N_4021);
nand U6417 (N_6417,N_3795,N_4230);
and U6418 (N_6418,N_4313,N_280);
nand U6419 (N_6419,N_1325,N_3869);
xnor U6420 (N_6420,N_3461,N_2715);
and U6421 (N_6421,N_3745,N_2605);
xnor U6422 (N_6422,N_3995,N_1557);
or U6423 (N_6423,N_1966,N_4156);
or U6424 (N_6424,N_538,N_786);
nand U6425 (N_6425,N_3421,N_2506);
nand U6426 (N_6426,N_3828,N_2347);
nor U6427 (N_6427,N_4856,N_4125);
and U6428 (N_6428,N_4364,N_3760);
nor U6429 (N_6429,N_2888,N_800);
or U6430 (N_6430,N_1652,N_1428);
nor U6431 (N_6431,N_1243,N_4809);
or U6432 (N_6432,N_8,N_3094);
nor U6433 (N_6433,N_759,N_2052);
xnor U6434 (N_6434,N_2369,N_3666);
nor U6435 (N_6435,N_4479,N_1013);
xor U6436 (N_6436,N_724,N_480);
xnor U6437 (N_6437,N_3242,N_3357);
or U6438 (N_6438,N_1452,N_860);
or U6439 (N_6439,N_3398,N_1218);
nor U6440 (N_6440,N_310,N_268);
nor U6441 (N_6441,N_4088,N_1769);
nor U6442 (N_6442,N_1534,N_1049);
xor U6443 (N_6443,N_1455,N_3888);
nand U6444 (N_6444,N_861,N_3660);
or U6445 (N_6445,N_3963,N_4945);
or U6446 (N_6446,N_1023,N_466);
or U6447 (N_6447,N_2221,N_3646);
xor U6448 (N_6448,N_4767,N_540);
or U6449 (N_6449,N_4799,N_4011);
or U6450 (N_6450,N_1279,N_2865);
xnor U6451 (N_6451,N_3012,N_1227);
xnor U6452 (N_6452,N_4090,N_2876);
and U6453 (N_6453,N_4038,N_2808);
or U6454 (N_6454,N_2673,N_2090);
and U6455 (N_6455,N_4707,N_2548);
nand U6456 (N_6456,N_4961,N_3402);
nand U6457 (N_6457,N_2053,N_2986);
xor U6458 (N_6458,N_890,N_959);
or U6459 (N_6459,N_2782,N_1079);
and U6460 (N_6460,N_284,N_971);
xor U6461 (N_6461,N_1908,N_3099);
or U6462 (N_6462,N_4636,N_1008);
nor U6463 (N_6463,N_4971,N_3532);
and U6464 (N_6464,N_2201,N_3654);
nand U6465 (N_6465,N_1962,N_1123);
nor U6466 (N_6466,N_1392,N_1183);
nand U6467 (N_6467,N_3643,N_3927);
xnor U6468 (N_6468,N_2462,N_3730);
or U6469 (N_6469,N_2728,N_713);
and U6470 (N_6470,N_2345,N_681);
nand U6471 (N_6471,N_26,N_3665);
nor U6472 (N_6472,N_2896,N_1036);
xor U6473 (N_6473,N_3833,N_2585);
or U6474 (N_6474,N_294,N_691);
and U6475 (N_6475,N_1233,N_3305);
xnor U6476 (N_6476,N_475,N_1827);
nand U6477 (N_6477,N_329,N_2171);
xor U6478 (N_6478,N_967,N_2327);
nor U6479 (N_6479,N_4605,N_605);
nand U6480 (N_6480,N_3829,N_1802);
xor U6481 (N_6481,N_3768,N_1019);
nand U6482 (N_6482,N_2264,N_1262);
or U6483 (N_6483,N_235,N_1813);
or U6484 (N_6484,N_4813,N_4583);
nand U6485 (N_6485,N_3119,N_2674);
nand U6486 (N_6486,N_2458,N_4369);
nor U6487 (N_6487,N_999,N_2828);
and U6488 (N_6488,N_3122,N_3847);
and U6489 (N_6489,N_2426,N_1122);
nor U6490 (N_6490,N_113,N_3659);
or U6491 (N_6491,N_3150,N_1234);
or U6492 (N_6492,N_2013,N_2797);
and U6493 (N_6493,N_4933,N_4386);
and U6494 (N_6494,N_4199,N_1697);
nand U6495 (N_6495,N_2697,N_1828);
nor U6496 (N_6496,N_635,N_4649);
nand U6497 (N_6497,N_963,N_1322);
and U6498 (N_6498,N_2877,N_2924);
and U6499 (N_6499,N_3980,N_483);
or U6500 (N_6500,N_4405,N_2412);
or U6501 (N_6501,N_2803,N_796);
or U6502 (N_6502,N_560,N_2764);
nand U6503 (N_6503,N_3332,N_4284);
xor U6504 (N_6504,N_4041,N_2753);
nor U6505 (N_6505,N_4265,N_2994);
nand U6506 (N_6506,N_4456,N_3845);
nor U6507 (N_6507,N_4114,N_4891);
or U6508 (N_6508,N_4475,N_3309);
or U6509 (N_6509,N_3701,N_1467);
or U6510 (N_6510,N_3550,N_3692);
xor U6511 (N_6511,N_4973,N_1229);
nand U6512 (N_6512,N_2588,N_1956);
or U6513 (N_6513,N_4789,N_4407);
nand U6514 (N_6514,N_1472,N_1030);
and U6515 (N_6515,N_4378,N_2860);
or U6516 (N_6516,N_2127,N_3929);
or U6517 (N_6517,N_493,N_2284);
nand U6518 (N_6518,N_3381,N_4814);
or U6519 (N_6519,N_1555,N_4082);
nand U6520 (N_6520,N_1138,N_2963);
nor U6521 (N_6521,N_4436,N_4717);
or U6522 (N_6522,N_1080,N_4823);
nor U6523 (N_6523,N_2861,N_1552);
nand U6524 (N_6524,N_3414,N_3295);
or U6525 (N_6525,N_2473,N_2017);
nand U6526 (N_6526,N_3566,N_600);
nand U6527 (N_6527,N_2958,N_3080);
xnor U6528 (N_6528,N_2629,N_4149);
or U6529 (N_6529,N_2105,N_4826);
nand U6530 (N_6530,N_2160,N_1960);
and U6531 (N_6531,N_1742,N_4186);
nand U6532 (N_6532,N_4337,N_3400);
nand U6533 (N_6533,N_1540,N_0);
or U6534 (N_6534,N_3014,N_2048);
or U6535 (N_6535,N_4460,N_183);
xor U6536 (N_6536,N_4935,N_360);
and U6537 (N_6537,N_1058,N_4976);
nor U6538 (N_6538,N_3699,N_4930);
or U6539 (N_6539,N_3301,N_1254);
or U6540 (N_6540,N_3189,N_2076);
or U6541 (N_6541,N_4681,N_2218);
nor U6542 (N_6542,N_3202,N_4057);
and U6543 (N_6543,N_1755,N_4796);
nor U6544 (N_6544,N_1793,N_3351);
or U6545 (N_6545,N_3047,N_1890);
and U6546 (N_6546,N_944,N_4157);
nand U6547 (N_6547,N_1274,N_491);
or U6548 (N_6548,N_616,N_1940);
nor U6549 (N_6549,N_2071,N_731);
or U6550 (N_6550,N_4932,N_172);
nand U6551 (N_6551,N_901,N_1723);
nand U6552 (N_6552,N_1217,N_3855);
nand U6553 (N_6553,N_920,N_171);
xnor U6554 (N_6554,N_3073,N_2010);
nor U6555 (N_6555,N_3032,N_664);
nand U6556 (N_6556,N_1561,N_888);
xor U6557 (N_6557,N_2232,N_249);
or U6558 (N_6558,N_1055,N_4519);
and U6559 (N_6559,N_3849,N_1164);
and U6560 (N_6560,N_1026,N_4825);
xor U6561 (N_6561,N_3528,N_1573);
xnor U6562 (N_6562,N_1912,N_2841);
or U6563 (N_6563,N_3559,N_4890);
xnor U6564 (N_6564,N_1316,N_2352);
or U6565 (N_6565,N_1850,N_2389);
or U6566 (N_6566,N_1129,N_633);
nand U6567 (N_6567,N_4702,N_580);
nand U6568 (N_6568,N_4224,N_2789);
nor U6569 (N_6569,N_2507,N_3933);
or U6570 (N_6570,N_4370,N_4972);
nor U6571 (N_6571,N_2516,N_1083);
or U6572 (N_6572,N_1275,N_3138);
and U6573 (N_6573,N_1391,N_46);
or U6574 (N_6574,N_3861,N_671);
nor U6575 (N_6575,N_4743,N_4120);
xnor U6576 (N_6576,N_2991,N_1880);
and U6577 (N_6577,N_3608,N_55);
and U6578 (N_6578,N_2844,N_4724);
nor U6579 (N_6579,N_846,N_3785);
nand U6580 (N_6580,N_1875,N_44);
and U6581 (N_6581,N_3647,N_2051);
nand U6582 (N_6582,N_3334,N_2383);
xor U6583 (N_6583,N_3324,N_3132);
and U6584 (N_6584,N_1084,N_2314);
or U6585 (N_6585,N_1853,N_2538);
nand U6586 (N_6586,N_389,N_2856);
nand U6587 (N_6587,N_2742,N_1011);
and U6588 (N_6588,N_3935,N_4759);
and U6589 (N_6589,N_1144,N_618);
and U6590 (N_6590,N_3903,N_4762);
nand U6591 (N_6591,N_4259,N_1626);
and U6592 (N_6592,N_3815,N_3274);
and U6593 (N_6593,N_3641,N_4718);
nor U6594 (N_6594,N_4466,N_2817);
nor U6595 (N_6595,N_950,N_2005);
nand U6596 (N_6596,N_1065,N_2072);
and U6597 (N_6597,N_3128,N_165);
nand U6598 (N_6598,N_767,N_1726);
nand U6599 (N_6599,N_912,N_3540);
nand U6600 (N_6600,N_3751,N_2754);
and U6601 (N_6601,N_4094,N_261);
nor U6602 (N_6602,N_423,N_3814);
nand U6603 (N_6603,N_2143,N_1921);
and U6604 (N_6604,N_4039,N_3694);
nor U6605 (N_6605,N_2437,N_2164);
or U6606 (N_6606,N_2631,N_4347);
nor U6607 (N_6607,N_1201,N_3471);
or U6608 (N_6608,N_636,N_974);
nor U6609 (N_6609,N_2031,N_954);
nand U6610 (N_6610,N_279,N_4343);
nand U6611 (N_6611,N_2146,N_3561);
xnor U6612 (N_6612,N_85,N_2395);
nor U6613 (N_6613,N_4092,N_1715);
or U6614 (N_6614,N_3562,N_3625);
xor U6615 (N_6615,N_891,N_4481);
nand U6616 (N_6616,N_1310,N_1352);
nor U6617 (N_6617,N_4719,N_4344);
and U6618 (N_6618,N_4571,N_763);
nor U6619 (N_6619,N_3622,N_3129);
or U6620 (N_6620,N_2312,N_4652);
nand U6621 (N_6621,N_1667,N_1395);
nor U6622 (N_6622,N_3644,N_1520);
nand U6623 (N_6623,N_4200,N_773);
and U6624 (N_6624,N_4946,N_1219);
nor U6625 (N_6625,N_1199,N_201);
and U6626 (N_6626,N_827,N_2349);
nor U6627 (N_6627,N_4742,N_4473);
xnor U6628 (N_6628,N_4913,N_4185);
nor U6629 (N_6629,N_673,N_2546);
nand U6630 (N_6630,N_3711,N_3513);
nand U6631 (N_6631,N_4610,N_3992);
nor U6632 (N_6632,N_3131,N_3276);
or U6633 (N_6633,N_3455,N_112);
or U6634 (N_6634,N_3840,N_2338);
xor U6635 (N_6635,N_1188,N_4146);
and U6636 (N_6636,N_661,N_1785);
xnor U6637 (N_6637,N_4884,N_2919);
or U6638 (N_6638,N_2477,N_4764);
and U6639 (N_6639,N_4498,N_2380);
xor U6640 (N_6640,N_2124,N_2471);
nor U6641 (N_6641,N_2872,N_4769);
nand U6642 (N_6642,N_668,N_2549);
nor U6643 (N_6643,N_3216,N_4806);
nand U6644 (N_6644,N_4306,N_1926);
nor U6645 (N_6645,N_3503,N_4725);
nor U6646 (N_6646,N_3797,N_4902);
and U6647 (N_6647,N_4723,N_59);
and U6648 (N_6648,N_4905,N_3084);
and U6649 (N_6649,N_1580,N_642);
xor U6650 (N_6650,N_1585,N_3093);
nor U6651 (N_6651,N_2914,N_708);
or U6652 (N_6652,N_2622,N_4453);
nor U6653 (N_6653,N_4361,N_795);
or U6654 (N_6654,N_4398,N_2466);
nor U6655 (N_6655,N_2007,N_554);
nor U6656 (N_6656,N_1077,N_2794);
xnor U6657 (N_6657,N_4805,N_2846);
nand U6658 (N_6658,N_1606,N_3675);
nor U6659 (N_6659,N_4615,N_2363);
nand U6660 (N_6660,N_2411,N_2045);
or U6661 (N_6661,N_4786,N_1379);
nor U6662 (N_6662,N_4014,N_4126);
nor U6663 (N_6663,N_4281,N_934);
nand U6664 (N_6664,N_1504,N_4018);
nor U6665 (N_6665,N_1897,N_2667);
or U6666 (N_6666,N_4530,N_3620);
and U6667 (N_6667,N_3523,N_4704);
and U6668 (N_6668,N_4593,N_1351);
nor U6669 (N_6669,N_3713,N_2374);
and U6670 (N_6670,N_3178,N_4404);
and U6671 (N_6671,N_243,N_176);
and U6672 (N_6672,N_2294,N_2831);
nand U6673 (N_6673,N_2118,N_2215);
and U6674 (N_6674,N_4693,N_1363);
or U6675 (N_6675,N_3997,N_4300);
and U6676 (N_6676,N_768,N_2720);
nand U6677 (N_6677,N_300,N_136);
nand U6678 (N_6678,N_1545,N_2004);
xor U6679 (N_6679,N_880,N_1941);
and U6680 (N_6680,N_2379,N_575);
nand U6681 (N_6681,N_2712,N_4292);
or U6682 (N_6682,N_1886,N_1370);
nor U6683 (N_6683,N_3977,N_376);
nor U6684 (N_6684,N_1445,N_1727);
nand U6685 (N_6685,N_508,N_997);
and U6686 (N_6686,N_1621,N_608);
and U6687 (N_6687,N_1898,N_3755);
or U6688 (N_6688,N_2691,N_849);
nor U6689 (N_6689,N_585,N_3810);
nand U6690 (N_6690,N_197,N_3377);
and U6691 (N_6691,N_3978,N_3969);
and U6692 (N_6692,N_2882,N_3570);
xor U6693 (N_6693,N_4531,N_4940);
or U6694 (N_6694,N_4622,N_887);
nand U6695 (N_6695,N_2249,N_2285);
nor U6696 (N_6696,N_4503,N_2985);
xor U6697 (N_6697,N_1743,N_161);
nor U6698 (N_6698,N_2519,N_398);
nand U6699 (N_6699,N_336,N_3425);
nor U6700 (N_6700,N_3853,N_3479);
and U6701 (N_6701,N_3514,N_687);
and U6702 (N_6702,N_3616,N_4209);
xnor U6703 (N_6703,N_2968,N_3848);
nor U6704 (N_6704,N_3284,N_231);
nand U6705 (N_6705,N_334,N_4699);
nor U6706 (N_6706,N_2902,N_1832);
nand U6707 (N_6707,N_3027,N_630);
nand U6708 (N_6708,N_2592,N_1789);
nor U6709 (N_6709,N_1135,N_4025);
nand U6710 (N_6710,N_4282,N_4423);
or U6711 (N_6711,N_4784,N_902);
or U6712 (N_6712,N_1350,N_204);
and U6713 (N_6713,N_2901,N_703);
and U6714 (N_6714,N_299,N_4657);
or U6715 (N_6715,N_1447,N_2713);
and U6716 (N_6716,N_1863,N_2029);
or U6717 (N_6717,N_3288,N_2913);
nand U6718 (N_6718,N_1220,N_1782);
or U6719 (N_6719,N_1776,N_4527);
or U6720 (N_6720,N_57,N_429);
nand U6721 (N_6721,N_1916,N_4350);
or U6722 (N_6722,N_4291,N_1047);
xnor U6723 (N_6723,N_576,N_1431);
nor U6724 (N_6724,N_2614,N_3371);
nor U6725 (N_6725,N_512,N_4222);
nand U6726 (N_6726,N_4414,N_2725);
xnor U6727 (N_6727,N_3700,N_1024);
nor U6728 (N_6728,N_496,N_3428);
nand U6729 (N_6729,N_486,N_1548);
or U6730 (N_6730,N_4103,N_2819);
nor U6731 (N_6731,N_1996,N_3942);
nand U6732 (N_6732,N_4208,N_3170);
nand U6733 (N_6733,N_702,N_2887);
nor U6734 (N_6734,N_4564,N_2732);
and U6735 (N_6735,N_1039,N_4779);
and U6736 (N_6736,N_3885,N_1922);
xnor U6737 (N_6737,N_4811,N_3354);
nor U6738 (N_6738,N_3273,N_3638);
nor U6739 (N_6739,N_3161,N_1721);
or U6740 (N_6740,N_4289,N_4899);
nand U6741 (N_6741,N_3759,N_101);
and U6742 (N_6742,N_4594,N_3408);
or U6743 (N_6743,N_4098,N_3702);
and U6744 (N_6744,N_4397,N_4866);
nand U6745 (N_6745,N_2421,N_2596);
or U6746 (N_6746,N_1308,N_3259);
and U6747 (N_6747,N_596,N_1286);
nor U6748 (N_6748,N_3938,N_2702);
and U6749 (N_6749,N_970,N_4251);
and U6750 (N_6750,N_2679,N_3443);
xor U6751 (N_6751,N_824,N_3002);
and U6752 (N_6752,N_2561,N_2009);
nor U6753 (N_6753,N_4153,N_2610);
or U6754 (N_6754,N_4392,N_3704);
nand U6755 (N_6755,N_4403,N_4506);
nand U6756 (N_6756,N_1184,N_4250);
nor U6757 (N_6757,N_2943,N_409);
nand U6758 (N_6758,N_1762,N_500);
nand U6759 (N_6759,N_418,N_1492);
nand U6760 (N_6760,N_1765,N_680);
nand U6761 (N_6761,N_1041,N_3612);
nand U6762 (N_6762,N_4023,N_2982);
and U6763 (N_6763,N_260,N_1740);
nand U6764 (N_6764,N_1330,N_984);
and U6765 (N_6765,N_397,N_181);
or U6766 (N_6766,N_709,N_2095);
nor U6767 (N_6767,N_4547,N_1553);
or U6768 (N_6768,N_2595,N_1208);
or U6769 (N_6769,N_897,N_3820);
nor U6770 (N_6770,N_3098,N_3016);
nor U6771 (N_6771,N_548,N_4446);
xor U6772 (N_6772,N_2365,N_102);
or U6773 (N_6773,N_1297,N_4535);
and U6774 (N_6774,N_1186,N_4432);
xnor U6775 (N_6775,N_1784,N_3716);
nand U6776 (N_6776,N_4904,N_4601);
xor U6777 (N_6777,N_4074,N_867);
nor U6778 (N_6778,N_3913,N_4545);
nor U6779 (N_6779,N_3064,N_955);
and U6780 (N_6780,N_4511,N_3606);
nand U6781 (N_6781,N_976,N_2078);
xnor U6782 (N_6782,N_4524,N_1301);
nand U6783 (N_6783,N_4994,N_2757);
or U6784 (N_6784,N_3918,N_2180);
or U6785 (N_6785,N_4426,N_741);
nor U6786 (N_6786,N_4233,N_4938);
nand U6787 (N_6787,N_1600,N_4061);
nand U6788 (N_6788,N_79,N_2550);
nand U6789 (N_6789,N_1380,N_250);
and U6790 (N_6790,N_1862,N_1292);
xor U6791 (N_6791,N_4520,N_1655);
and U6792 (N_6792,N_4944,N_1868);
nand U6793 (N_6793,N_3193,N_4626);
and U6794 (N_6794,N_916,N_1421);
or U6795 (N_6795,N_3363,N_4572);
xnor U6796 (N_6796,N_4002,N_4327);
or U6797 (N_6797,N_253,N_4860);
or U6798 (N_6798,N_220,N_3741);
and U6799 (N_6799,N_603,N_4928);
nor U6800 (N_6800,N_2575,N_3142);
nand U6801 (N_6801,N_551,N_142);
nand U6802 (N_6802,N_544,N_510);
or U6803 (N_6803,N_3220,N_1970);
or U6804 (N_6804,N_33,N_246);
nor U6805 (N_6805,N_1124,N_3989);
and U6806 (N_6806,N_3386,N_2854);
nor U6807 (N_6807,N_2533,N_2964);
nor U6808 (N_6808,N_1446,N_3923);
nor U6809 (N_6809,N_3551,N_2422);
nand U6810 (N_6810,N_4534,N_2906);
nor U6811 (N_6811,N_1204,N_1653);
and U6812 (N_6812,N_854,N_943);
nor U6813 (N_6813,N_4440,N_853);
and U6814 (N_6814,N_4015,N_4085);
or U6815 (N_6815,N_234,N_2253);
or U6816 (N_6816,N_367,N_2177);
nor U6817 (N_6817,N_3880,N_666);
xnor U6818 (N_6818,N_4595,N_4043);
and U6819 (N_6819,N_1645,N_2799);
and U6820 (N_6820,N_4320,N_341);
nor U6821 (N_6821,N_2357,N_1603);
nor U6822 (N_6822,N_1359,N_2716);
nand U6823 (N_6823,N_1120,N_2192);
nor U6824 (N_6824,N_1222,N_3362);
nand U6825 (N_6825,N_63,N_4999);
xnor U6826 (N_6826,N_4037,N_83);
nand U6827 (N_6827,N_4607,N_485);
nand U6828 (N_6828,N_366,N_1867);
and U6829 (N_6829,N_2792,N_2509);
nand U6830 (N_6830,N_662,N_2479);
or U6831 (N_6831,N_2277,N_1414);
and U6832 (N_6832,N_4318,N_42);
nand U6833 (N_6833,N_103,N_208);
or U6834 (N_6834,N_4602,N_1576);
or U6835 (N_6835,N_2211,N_704);
nor U6836 (N_6836,N_2364,N_2464);
nand U6837 (N_6837,N_2746,N_4187);
nand U6838 (N_6838,N_3436,N_381);
nor U6839 (N_6839,N_2874,N_1085);
nand U6840 (N_6840,N_1491,N_1605);
and U6841 (N_6841,N_2465,N_4709);
nor U6842 (N_6842,N_2439,N_1666);
xnor U6843 (N_6843,N_4857,N_2400);
nand U6844 (N_6844,N_4093,N_4666);
xor U6845 (N_6845,N_2240,N_4744);
and U6846 (N_6846,N_1232,N_4861);
nor U6847 (N_6847,N_3124,N_2263);
nand U6848 (N_6848,N_1501,N_4864);
and U6849 (N_6849,N_719,N_3502);
nor U6850 (N_6850,N_675,N_2227);
and U6851 (N_6851,N_426,N_2377);
or U6852 (N_6852,N_221,N_2905);
or U6853 (N_6853,N_4477,N_3303);
nand U6854 (N_6854,N_621,N_1018);
nor U6855 (N_6855,N_742,N_2995);
xnor U6856 (N_6856,N_4773,N_3601);
xnor U6857 (N_6857,N_2761,N_1858);
xor U6858 (N_6858,N_1541,N_159);
or U6859 (N_6859,N_1527,N_4084);
and U6860 (N_6860,N_318,N_11);
nor U6861 (N_6861,N_4317,N_938);
nor U6862 (N_6862,N_2745,N_4734);
or U6863 (N_6863,N_313,N_735);
or U6864 (N_6864,N_3698,N_4746);
nand U6865 (N_6865,N_613,N_684);
nand U6866 (N_6866,N_883,N_3652);
nand U6867 (N_6867,N_1196,N_1597);
nand U6868 (N_6868,N_1114,N_3217);
nor U6869 (N_6869,N_3205,N_3419);
nor U6870 (N_6870,N_51,N_2637);
nor U6871 (N_6871,N_4858,N_2188);
and U6872 (N_6872,N_2497,N_2937);
nand U6873 (N_6873,N_1914,N_525);
nor U6874 (N_6874,N_936,N_3791);
or U6875 (N_6875,N_3790,N_4726);
and U6876 (N_6876,N_528,N_3451);
or U6877 (N_6877,N_2554,N_2183);
or U6878 (N_6878,N_716,N_3789);
nor U6879 (N_6879,N_1081,N_811);
nand U6880 (N_6880,N_3637,N_2424);
or U6881 (N_6881,N_4454,N_1823);
xor U6882 (N_6882,N_942,N_1584);
nor U6883 (N_6883,N_2796,N_2234);
nor U6884 (N_6884,N_425,N_2392);
or U6885 (N_6885,N_3152,N_535);
nand U6886 (N_6886,N_1471,N_1240);
nor U6887 (N_6887,N_2655,N_1119);
nor U6888 (N_6888,N_4828,N_3260);
and U6889 (N_6889,N_4266,N_490);
nand U6890 (N_6890,N_2134,N_4573);
and U6891 (N_6891,N_3761,N_3175);
or U6892 (N_6892,N_342,N_2073);
nor U6893 (N_6893,N_1010,N_4669);
nand U6894 (N_6894,N_830,N_1315);
nand U6895 (N_6895,N_4507,N_2999);
and U6896 (N_6896,N_3626,N_1662);
and U6897 (N_6897,N_148,N_1945);
nor U6898 (N_6898,N_4517,N_1272);
nor U6899 (N_6899,N_2259,N_1331);
nand U6900 (N_6900,N_3317,N_4880);
and U6901 (N_6901,N_1436,N_4671);
nor U6902 (N_6902,N_1051,N_779);
nor U6903 (N_6903,N_1481,N_3133);
or U6904 (N_6904,N_4207,N_2563);
or U6905 (N_6905,N_2480,N_2918);
or U6906 (N_6906,N_561,N_3130);
or U6907 (N_6907,N_3025,N_1362);
nor U6908 (N_6908,N_3352,N_4001);
or U6909 (N_6909,N_1130,N_4163);
and U6910 (N_6910,N_730,N_925);
nand U6911 (N_6911,N_238,N_4612);
xor U6912 (N_6912,N_188,N_2304);
nor U6913 (N_6913,N_1289,N_2408);
and U6914 (N_6914,N_1003,N_4682);
xor U6915 (N_6915,N_4589,N_578);
nor U6916 (N_6916,N_3808,N_3633);
nor U6917 (N_6917,N_3271,N_4837);
nor U6918 (N_6918,N_2212,N_4578);
xor U6919 (N_6919,N_100,N_3141);
xor U6920 (N_6920,N_3223,N_1514);
and U6921 (N_6921,N_1357,N_2925);
or U6922 (N_6922,N_4389,N_825);
and U6923 (N_6923,N_3908,N_688);
nor U6924 (N_6924,N_3250,N_3328);
nand U6925 (N_6925,N_1794,N_4035);
or U6926 (N_6926,N_3136,N_4992);
nor U6927 (N_6927,N_566,N_2784);
or U6928 (N_6928,N_3207,N_1375);
nor U6929 (N_6929,N_3480,N_3272);
and U6930 (N_6930,N_1607,N_2768);
or U6931 (N_6931,N_3706,N_3062);
or U6932 (N_6932,N_1582,N_1935);
and U6933 (N_6933,N_259,N_3725);
nor U6934 (N_6934,N_4383,N_3928);
nor U6935 (N_6935,N_798,N_588);
nor U6936 (N_6936,N_3081,N_1265);
nor U6937 (N_6937,N_3265,N_447);
and U6938 (N_6938,N_4735,N_4495);
or U6939 (N_6939,N_1648,N_4167);
nor U6940 (N_6940,N_1798,N_604);
and U6941 (N_6941,N_169,N_2929);
nor U6942 (N_6942,N_3740,N_2457);
or U6943 (N_6943,N_2282,N_3249);
or U6944 (N_6944,N_1768,N_614);
and U6945 (N_6945,N_3944,N_308);
nor U6946 (N_6946,N_2802,N_1770);
nor U6947 (N_6947,N_3239,N_2474);
nor U6948 (N_6948,N_4874,N_2591);
and U6949 (N_6949,N_2037,N_1857);
nor U6950 (N_6950,N_2897,N_146);
nand U6951 (N_6951,N_4952,N_3508);
nand U6952 (N_6952,N_1250,N_4662);
and U6953 (N_6953,N_986,N_1959);
nor U6954 (N_6954,N_4160,N_185);
nand U6955 (N_6955,N_981,N_2332);
and U6956 (N_6956,N_2040,N_4470);
nand U6957 (N_6957,N_3782,N_2724);
nand U6958 (N_6958,N_996,N_218);
nor U6959 (N_6959,N_216,N_2522);
and U6960 (N_6960,N_1156,N_3518);
nand U6961 (N_6961,N_416,N_4698);
and U6962 (N_6962,N_2092,N_2616);
xnor U6963 (N_6963,N_2569,N_3167);
and U6964 (N_6964,N_3411,N_4356);
and U6965 (N_6965,N_2275,N_2431);
or U6966 (N_6966,N_597,N_1521);
nor U6967 (N_6967,N_1766,N_4624);
nand U6968 (N_6968,N_3509,N_2011);
or U6969 (N_6969,N_1590,N_3038);
nor U6970 (N_6970,N_2455,N_3457);
and U6971 (N_6971,N_3811,N_4697);
nand U6972 (N_6972,N_384,N_3945);
nand U6973 (N_6973,N_3110,N_2568);
or U6974 (N_6974,N_330,N_1747);
and U6975 (N_6975,N_4467,N_4497);
and U6976 (N_6976,N_2770,N_2182);
and U6977 (N_6977,N_3197,N_1810);
and U6978 (N_6978,N_1767,N_3599);
or U6979 (N_6979,N_4178,N_4645);
or U6980 (N_6980,N_4908,N_3603);
nand U6981 (N_6981,N_2613,N_4942);
xor U6982 (N_6982,N_479,N_3103);
nand U6983 (N_6983,N_1182,N_1799);
and U6984 (N_6984,N_4911,N_4064);
nor U6985 (N_6985,N_1609,N_628);
xnor U6986 (N_6986,N_2041,N_3333);
nand U6987 (N_6987,N_3890,N_4557);
or U6988 (N_6988,N_4537,N_3287);
or U6989 (N_6989,N_372,N_3615);
nor U6990 (N_6990,N_2181,N_2268);
and U6991 (N_6991,N_4631,N_4909);
and U6992 (N_6992,N_3088,N_2678);
or U6993 (N_6993,N_2690,N_1337);
and U6994 (N_6994,N_2862,N_2231);
and U6995 (N_6995,N_2584,N_521);
nand U6996 (N_6996,N_988,N_2903);
nor U6997 (N_6997,N_2858,N_899);
xnor U6998 (N_6998,N_3736,N_3770);
or U6999 (N_6999,N_898,N_2608);
or U7000 (N_7000,N_4295,N_4588);
xnor U7001 (N_7001,N_2406,N_1381);
or U7002 (N_7002,N_3613,N_2342);
xnor U7003 (N_7003,N_4353,N_3746);
or U7004 (N_7004,N_907,N_592);
nor U7005 (N_7005,N_3996,N_1856);
xnor U7006 (N_7006,N_647,N_460);
or U7007 (N_7007,N_1344,N_1348);
nand U7008 (N_7008,N_331,N_2820);
or U7009 (N_7009,N_2545,N_2438);
and U7010 (N_7010,N_326,N_4642);
nor U7011 (N_7011,N_3593,N_1172);
nand U7012 (N_7012,N_4516,N_1617);
nand U7013 (N_7013,N_4109,N_534);
nand U7014 (N_7014,N_3758,N_1475);
nor U7015 (N_7015,N_2137,N_4651);
nand U7016 (N_7016,N_288,N_3669);
nand U7017 (N_7017,N_2517,N_632);
xor U7018 (N_7018,N_396,N_4889);
nor U7019 (N_7019,N_728,N_1284);
or U7020 (N_7020,N_2079,N_175);
and U7021 (N_7021,N_1062,N_2414);
and U7022 (N_7022,N_4472,N_4713);
nor U7023 (N_7023,N_3680,N_4579);
nand U7024 (N_7024,N_3817,N_1816);
nor U7025 (N_7025,N_4872,N_956);
nor U7026 (N_7026,N_2139,N_1618);
or U7027 (N_7027,N_441,N_3078);
nor U7028 (N_7028,N_1895,N_2189);
nor U7029 (N_7029,N_3427,N_3564);
or U7030 (N_7030,N_352,N_2624);
nand U7031 (N_7031,N_1001,N_4988);
or U7032 (N_7032,N_3268,N_4298);
or U7033 (N_7033,N_3163,N_1503);
and U7034 (N_7034,N_4841,N_4427);
xnor U7035 (N_7035,N_2685,N_835);
nand U7036 (N_7036,N_2353,N_1165);
or U7037 (N_7037,N_4159,N_1442);
nor U7038 (N_7038,N_2101,N_2235);
or U7039 (N_7039,N_421,N_410);
nor U7040 (N_7040,N_1327,N_4141);
nor U7041 (N_7041,N_2701,N_4627);
nand U7042 (N_7042,N_4756,N_3017);
or U7043 (N_7043,N_2916,N_4290);
nor U7044 (N_7044,N_843,N_1623);
xnor U7045 (N_7045,N_2762,N_1663);
and U7046 (N_7046,N_4638,N_1795);
and U7047 (N_7047,N_4042,N_1153);
and U7048 (N_7048,N_3580,N_4771);
or U7049 (N_7049,N_4659,N_4260);
or U7050 (N_7050,N_1145,N_80);
nand U7051 (N_7051,N_4488,N_1300);
xor U7052 (N_7052,N_73,N_2756);
nor U7053 (N_7053,N_1928,N_1264);
nor U7054 (N_7054,N_3703,N_147);
or U7055 (N_7055,N_1167,N_4613);
nor U7056 (N_7056,N_3690,N_1999);
nand U7057 (N_7057,N_2324,N_2987);
and U7058 (N_7058,N_2030,N_4147);
xnor U7059 (N_7059,N_1872,N_4559);
xor U7060 (N_7060,N_293,N_994);
or U7061 (N_7061,N_3210,N_382);
and U7062 (N_7062,N_1203,N_1686);
xnor U7063 (N_7063,N_1027,N_2949);
nand U7064 (N_7064,N_1499,N_3433);
nand U7065 (N_7065,N_802,N_2530);
nand U7066 (N_7066,N_4923,N_1376);
or U7067 (N_7067,N_3490,N_3868);
and U7068 (N_7068,N_3279,N_106);
and U7069 (N_7069,N_1668,N_2190);
or U7070 (N_7070,N_755,N_3653);
or U7071 (N_7071,N_3781,N_3404);
nor U7072 (N_7072,N_3244,N_2089);
nand U7073 (N_7073,N_2396,N_4261);
nand U7074 (N_7074,N_1628,N_2501);
and U7075 (N_7075,N_3263,N_1773);
and U7076 (N_7076,N_3102,N_2442);
xor U7077 (N_7077,N_2970,N_1406);
nand U7078 (N_7078,N_4296,N_2769);
and U7079 (N_7079,N_2494,N_670);
or U7080 (N_7080,N_3361,N_4499);
nor U7081 (N_7081,N_286,N_2707);
or U7082 (N_7082,N_2144,N_2435);
and U7083 (N_7083,N_3976,N_4633);
nand U7084 (N_7084,N_3619,N_4409);
nor U7085 (N_7085,N_2508,N_1210);
and U7086 (N_7086,N_4264,N_4736);
nor U7087 (N_7087,N_3146,N_3349);
nor U7088 (N_7088,N_2173,N_3359);
and U7089 (N_7089,N_3764,N_3909);
or U7090 (N_7090,N_3714,N_2233);
or U7091 (N_7091,N_869,N_1622);
and U7092 (N_7092,N_3388,N_2114);
xnor U7093 (N_7093,N_756,N_3749);
nand U7094 (N_7094,N_4738,N_1639);
or U7095 (N_7095,N_1947,N_2067);
nand U7096 (N_7096,N_3395,N_4523);
and U7097 (N_7097,N_4101,N_199);
and U7098 (N_7098,N_262,N_3844);
nor U7099 (N_7099,N_2459,N_4393);
or U7100 (N_7100,N_4941,N_4676);
or U7101 (N_7101,N_506,N_2749);
nor U7102 (N_7102,N_1413,N_355);
xor U7103 (N_7103,N_1411,N_4158);
and U7104 (N_7104,N_76,N_583);
nor U7105 (N_7105,N_1775,N_2496);
and U7106 (N_7106,N_2600,N_3091);
nand U7107 (N_7107,N_2476,N_4276);
nor U7108 (N_7108,N_2346,N_1105);
nor U7109 (N_7109,N_3464,N_4646);
nor U7110 (N_7110,N_1969,N_2528);
nor U7111 (N_7111,N_1136,N_1112);
nor U7112 (N_7112,N_1616,N_1735);
nor U7113 (N_7113,N_1448,N_2348);
and U7114 (N_7114,N_1537,N_4);
or U7115 (N_7115,N_1833,N_3556);
and U7116 (N_7116,N_1185,N_3892);
nand U7117 (N_7117,N_568,N_3689);
and U7118 (N_7118,N_2979,N_3035);
nor U7119 (N_7119,N_4330,N_3624);
and U7120 (N_7120,N_4868,N_1564);
nor U7121 (N_7121,N_6,N_1384);
nand U7122 (N_7122,N_650,N_3629);
xnor U7123 (N_7123,N_3390,N_1532);
and U7124 (N_7124,N_2216,N_4384);
or U7125 (N_7125,N_1754,N_4827);
nor U7126 (N_7126,N_403,N_3313);
nor U7127 (N_7127,N_236,N_2680);
nand U7128 (N_7128,N_4997,N_4196);
nor U7129 (N_7129,N_1178,N_3723);
nor U7130 (N_7130,N_1848,N_3510);
and U7131 (N_7131,N_2302,N_939);
or U7132 (N_7132,N_1111,N_2362);
and U7133 (N_7133,N_2257,N_2152);
or U7134 (N_7134,N_379,N_3951);
xnor U7135 (N_7135,N_214,N_1729);
nor U7136 (N_7136,N_958,N_1197);
xnor U7137 (N_7137,N_518,N_4246);
nand U7138 (N_7138,N_2838,N_1907);
nand U7139 (N_7139,N_2330,N_4623);
xnor U7140 (N_7140,N_3366,N_91);
xnor U7141 (N_7141,N_2830,N_2068);
or U7142 (N_7142,N_4144,N_4803);
nor U7143 (N_7143,N_67,N_3896);
and U7144 (N_7144,N_35,N_1223);
nand U7145 (N_7145,N_820,N_4303);
nand U7146 (N_7146,N_1891,N_1974);
and U7147 (N_7147,N_526,N_2825);
or U7148 (N_7148,N_1865,N_454);
or U7149 (N_7149,N_1611,N_3585);
nand U7150 (N_7150,N_4390,N_3399);
and U7151 (N_7151,N_3753,N_320);
and U7152 (N_7152,N_2695,N_3642);
or U7153 (N_7153,N_4137,N_4211);
nand U7154 (N_7154,N_4182,N_72);
nor U7155 (N_7155,N_765,N_1371);
and U7156 (N_7156,N_1771,N_3907);
or U7157 (N_7157,N_3685,N_4745);
xnor U7158 (N_7158,N_4996,N_844);
nand U7159 (N_7159,N_1955,N_4663);
nand U7160 (N_7160,N_1476,N_1075);
nand U7161 (N_7161,N_1817,N_43);
or U7162 (N_7162,N_2752,N_1396);
or U7163 (N_7163,N_951,N_2170);
xnor U7164 (N_7164,N_4956,N_494);
nor U7165 (N_7165,N_3984,N_4575);
nand U7166 (N_7166,N_1682,N_2002);
xnor U7167 (N_7167,N_2586,N_497);
and U7168 (N_7168,N_4853,N_3681);
nor U7169 (N_7169,N_3607,N_4307);
and U7170 (N_7170,N_108,N_4710);
nand U7171 (N_7171,N_4529,N_1094);
nand U7172 (N_7172,N_3732,N_3621);
nand U7173 (N_7173,N_4065,N_4255);
nand U7174 (N_7174,N_1369,N_3252);
and U7175 (N_7175,N_281,N_1175);
nor U7176 (N_7176,N_4097,N_433);
nand U7177 (N_7177,N_1283,N_2531);
nand U7178 (N_7178,N_2191,N_1563);
nand U7179 (N_7179,N_2894,N_3121);
nand U7180 (N_7180,N_2532,N_1420);
or U7181 (N_7181,N_3987,N_2993);
nand U7182 (N_7182,N_133,N_3610);
nand U7183 (N_7183,N_876,N_3280);
nand U7184 (N_7184,N_3640,N_2418);
or U7185 (N_7185,N_2891,N_808);
nand U7186 (N_7186,N_3089,N_3834);
and U7187 (N_7187,N_3290,N_1259);
nor U7188 (N_7188,N_807,N_2723);
or U7189 (N_7189,N_1869,N_4206);
and U7190 (N_7190,N_104,N_4054);
and U7191 (N_7191,N_1169,N_3631);
nor U7192 (N_7192,N_4425,N_1934);
nand U7193 (N_7193,N_4802,N_2074);
nand U7194 (N_7194,N_2147,N_4478);
and U7195 (N_7195,N_4076,N_3033);
nand U7196 (N_7196,N_2664,N_3353);
or U7197 (N_7197,N_3251,N_4722);
nand U7198 (N_7198,N_459,N_132);
and U7199 (N_7199,N_2821,N_2504);
nand U7200 (N_7200,N_4798,N_4752);
nor U7201 (N_7201,N_858,N_49);
and U7202 (N_7202,N_3097,N_1982);
nor U7203 (N_7203,N_4124,N_4203);
and U7204 (N_7204,N_229,N_2513);
nand U7205 (N_7205,N_1118,N_904);
nand U7206 (N_7206,N_1679,N_4780);
and U7207 (N_7207,N_407,N_1290);
nor U7208 (N_7208,N_3456,N_3825);
and U7209 (N_7209,N_4450,N_1929);
and U7210 (N_7210,N_638,N_3208);
or U7211 (N_7211,N_2672,N_1684);
nand U7212 (N_7212,N_377,N_3045);
nor U7213 (N_7213,N_669,N_354);
and U7214 (N_7214,N_2265,N_1497);
xnor U7215 (N_7215,N_4783,N_2881);
nor U7216 (N_7216,N_2280,N_413);
nand U7217 (N_7217,N_2208,N_836);
nor U7218 (N_7218,N_651,N_987);
nor U7219 (N_7219,N_3934,N_1043);
or U7220 (N_7220,N_1577,N_2805);
or U7221 (N_7221,N_842,N_2084);
and U7222 (N_7222,N_4887,N_4102);
nand U7223 (N_7223,N_1558,N_1731);
and U7224 (N_7224,N_780,N_338);
nor U7225 (N_7225,N_1465,N_239);
xor U7226 (N_7226,N_2219,N_772);
nand U7227 (N_7227,N_543,N_4445);
nor U7228 (N_7228,N_2209,N_4569);
or U7229 (N_7229,N_1061,N_2880);
nand U7230 (N_7230,N_4504,N_989);
nand U7231 (N_7231,N_442,N_1885);
nor U7232 (N_7232,N_2977,N_2112);
xnor U7233 (N_7233,N_1792,N_1882);
nand U7234 (N_7234,N_4715,N_3051);
and U7235 (N_7235,N_2136,N_2553);
or U7236 (N_7236,N_4268,N_1593);
or U7237 (N_7237,N_1674,N_2653);
nor U7238 (N_7238,N_3298,N_922);
and U7239 (N_7239,N_4073,N_4116);
and U7240 (N_7240,N_266,N_438);
or U7241 (N_7241,N_373,N_3306);
nand U7242 (N_7242,N_1040,N_4075);
nor U7243 (N_7243,N_1044,N_3370);
xnor U7244 (N_7244,N_2083,N_70);
nand U7245 (N_7245,N_3194,N_2121);
and U7246 (N_7246,N_462,N_4855);
xor U7247 (N_7247,N_2301,N_3415);
xor U7248 (N_7248,N_2470,N_3100);
or U7249 (N_7249,N_2080,N_3754);
nand U7250 (N_7250,N_40,N_1042);
nand U7251 (N_7251,N_4168,N_4231);
nor U7252 (N_7252,N_4712,N_4644);
or U7253 (N_7253,N_1840,N_4133);
or U7254 (N_7254,N_2627,N_2388);
nor U7255 (N_7255,N_3778,N_4683);
or U7256 (N_7256,N_2025,N_4113);
xor U7257 (N_7257,N_3469,N_1108);
and U7258 (N_7258,N_2572,N_4234);
nor U7259 (N_7259,N_31,N_3727);
xor U7260 (N_7260,N_4850,N_1562);
or U7261 (N_7261,N_2420,N_4653);
and U7262 (N_7262,N_65,N_965);
and U7263 (N_7263,N_1983,N_2370);
xor U7264 (N_7264,N_2947,N_1280);
nor U7265 (N_7265,N_2618,N_1098);
or U7266 (N_7266,N_414,N_3602);
or U7267 (N_7267,N_1088,N_705);
and U7268 (N_7268,N_2223,N_2542);
nand U7269 (N_7269,N_2168,N_964);
and U7270 (N_7270,N_4489,N_4761);
nor U7271 (N_7271,N_3809,N_4323);
or U7272 (N_7272,N_54,N_4274);
xor U7273 (N_7273,N_1702,N_411);
and U7274 (N_7274,N_179,N_3729);
nand U7275 (N_7275,N_4455,N_1430);
and U7276 (N_7276,N_3632,N_138);
or U7277 (N_7277,N_3253,N_4491);
nor U7278 (N_7278,N_1000,N_3143);
nand U7279 (N_7279,N_2909,N_2151);
or U7280 (N_7280,N_3818,N_3338);
nand U7281 (N_7281,N_2482,N_4145);
nand U7282 (N_7282,N_2644,N_144);
or U7283 (N_7283,N_761,N_2372);
and U7284 (N_7284,N_2034,N_1814);
nor U7285 (N_7285,N_1382,N_4367);
or U7286 (N_7286,N_2870,N_195);
nor U7287 (N_7287,N_3262,N_153);
xor U7288 (N_7288,N_95,N_4694);
nand U7289 (N_7289,N_4984,N_4424);
and U7290 (N_7290,N_3391,N_478);
or U7291 (N_7291,N_2602,N_4371);
or U7292 (N_7292,N_3058,N_2449);
or U7293 (N_7293,N_2778,N_170);
nor U7294 (N_7294,N_4974,N_2056);
and U7295 (N_7295,N_1393,N_36);
and U7296 (N_7296,N_542,N_2097);
nand U7297 (N_7297,N_3775,N_210);
or U7298 (N_7298,N_1408,N_3916);
or U7299 (N_7299,N_2461,N_3686);
nand U7300 (N_7300,N_1121,N_4220);
nor U7301 (N_7301,N_2094,N_3382);
and U7302 (N_7302,N_4348,N_1012);
nor U7303 (N_7303,N_1177,N_3851);
nand U7304 (N_7304,N_804,N_3747);
xnor U7305 (N_7305,N_1944,N_643);
or U7306 (N_7306,N_3393,N_2801);
xor U7307 (N_7307,N_363,N_3343);
nor U7308 (N_7308,N_114,N_1764);
nand U7309 (N_7309,N_417,N_1796);
nand U7310 (N_7310,N_4546,N_1335);
nor U7311 (N_7311,N_3410,N_1486);
or U7312 (N_7312,N_812,N_1530);
nor U7313 (N_7313,N_1247,N_2393);
xnor U7314 (N_7314,N_1915,N_2577);
and U7315 (N_7315,N_700,N_919);
nor U7316 (N_7316,N_4700,N_252);
or U7317 (N_7317,N_3858,N_3981);
or U7318 (N_7318,N_2367,N_1583);
nor U7319 (N_7319,N_81,N_3571);
xnor U7320 (N_7320,N_4787,N_117);
nand U7321 (N_7321,N_4878,N_3177);
xor U7322 (N_7322,N_3001,N_697);
and U7323 (N_7323,N_422,N_32);
nor U7324 (N_7324,N_2628,N_3199);
or U7325 (N_7325,N_1708,N_537);
nand U7326 (N_7326,N_274,N_1288);
nand U7327 (N_7327,N_929,N_2162);
and U7328 (N_7328,N_3826,N_3019);
or U7329 (N_7329,N_296,N_1320);
xor U7330 (N_7330,N_3522,N_4647);
or U7331 (N_7331,N_4929,N_129);
or U7332 (N_7332,N_191,N_1808);
xnor U7333 (N_7333,N_3650,N_1373);
nor U7334 (N_7334,N_4223,N_1567);
nor U7335 (N_7335,N_387,N_3898);
or U7336 (N_7336,N_4052,N_1749);
and U7337 (N_7337,N_1374,N_3431);
or U7338 (N_7338,N_2020,N_2279);
and U7339 (N_7339,N_1388,N_917);
xor U7340 (N_7340,N_1307,N_4415);
and U7341 (N_7341,N_1214,N_4774);
or U7342 (N_7342,N_1444,N_2319);
nor U7343 (N_7343,N_4648,N_1487);
and U7344 (N_7344,N_2006,N_2883);
nand U7345 (N_7345,N_533,N_2503);
or U7346 (N_7346,N_3655,N_472);
nand U7347 (N_7347,N_4879,N_2026);
nand U7348 (N_7348,N_134,N_3069);
and U7349 (N_7349,N_1800,N_1239);
or U7350 (N_7350,N_356,N_2176);
nor U7351 (N_7351,N_3941,N_2447);
nor U7352 (N_7352,N_1964,N_3446);
nor U7353 (N_7353,N_96,N_4748);
and U7354 (N_7354,N_2866,N_3752);
nand U7355 (N_7355,N_3182,N_1101);
and U7356 (N_7356,N_4824,N_3743);
nand U7357 (N_7357,N_991,N_4897);
and U7358 (N_7358,N_4066,N_2969);
nor U7359 (N_7359,N_1347,N_3671);
xnor U7360 (N_7360,N_1163,N_2927);
nand U7361 (N_7361,N_4493,N_194);
nand U7362 (N_7362,N_746,N_2850);
nor U7363 (N_7363,N_1064,N_2417);
or U7364 (N_7364,N_2936,N_4030);
and U7365 (N_7365,N_2081,N_1173);
or U7366 (N_7366,N_2022,N_492);
nor U7367 (N_7367,N_1409,N_1806);
nand U7368 (N_7368,N_1401,N_3172);
or U7369 (N_7369,N_2335,N_39);
xor U7370 (N_7370,N_4881,N_3823);
or U7371 (N_7371,N_1874,N_3474);
nand U7372 (N_7372,N_885,N_375);
nor U7373 (N_7373,N_325,N_738);
nor U7374 (N_7374,N_118,N_865);
xor U7375 (N_7375,N_1625,N_4154);
nand U7376 (N_7376,N_1707,N_3688);
or U7377 (N_7377,N_3173,N_3925);
or U7378 (N_7378,N_3036,N_1281);
and U7379 (N_7379,N_4562,N_2271);
or U7380 (N_7380,N_3517,N_21);
nor U7381 (N_7381,N_2682,N_1772);
or U7382 (N_7382,N_3015,N_1719);
and U7383 (N_7383,N_2490,N_2747);
or U7384 (N_7384,N_2397,N_831);
nand U7385 (N_7385,N_2161,N_2818);
or U7386 (N_7386,N_1179,N_2251);
or U7387 (N_7387,N_1299,N_1968);
xor U7388 (N_7388,N_1732,N_646);
nand U7389 (N_7389,N_4294,N_272);
nor U7390 (N_7390,N_4540,N_3878);
and U7391 (N_7391,N_1479,N_4316);
nor U7392 (N_7392,N_1513,N_1074);
nor U7393 (N_7393,N_517,N_4521);
nand U7394 (N_7394,N_2153,N_693);
nor U7395 (N_7395,N_631,N_2283);
nor U7396 (N_7396,N_3766,N_1910);
or U7397 (N_7397,N_4949,N_2103);
nand U7398 (N_7398,N_737,N_3285);
nor U7399 (N_7399,N_1612,N_3462);
and U7400 (N_7400,N_857,N_1778);
or U7401 (N_7401,N_3893,N_3037);
nand U7402 (N_7402,N_4119,N_348);
nor U7403 (N_7403,N_428,N_4568);
nor U7404 (N_7404,N_3046,N_1493);
and U7405 (N_7405,N_3437,N_1519);
nand U7406 (N_7406,N_1383,N_3589);
and U7407 (N_7407,N_2552,N_3057);
nand U7408 (N_7408,N_4212,N_2398);
or U7409 (N_7409,N_2640,N_1985);
xor U7410 (N_7410,N_4480,N_1399);
nor U7411 (N_7411,N_1649,N_2086);
nand U7412 (N_7412,N_4845,N_1818);
or U7413 (N_7413,N_2758,N_1087);
nor U7414 (N_7414,N_1317,N_3114);
or U7415 (N_7415,N_4299,N_2416);
nor U7416 (N_7416,N_3617,N_3496);
nor U7417 (N_7417,N_717,N_4164);
or U7418 (N_7418,N_13,N_2356);
and U7419 (N_7419,N_206,N_3156);
xnor U7420 (N_7420,N_2529,N_757);
nor U7421 (N_7421,N_748,N_1505);
nand U7422 (N_7422,N_2290,N_126);
and U7423 (N_7423,N_4867,N_2599);
and U7424 (N_7424,N_871,N_2668);
or U7425 (N_7425,N_2,N_4555);
and U7426 (N_7426,N_2229,N_1271);
and U7427 (N_7427,N_233,N_455);
or U7428 (N_7428,N_720,N_2696);
or U7429 (N_7429,N_3965,N_3105);
nor U7430 (N_7430,N_1181,N_307);
xor U7431 (N_7431,N_1237,N_306);
nor U7432 (N_7432,N_1489,N_3321);
or U7433 (N_7433,N_2409,N_3678);
or U7434 (N_7434,N_1053,N_3891);
nand U7435 (N_7435,N_3331,N_324);
and U7436 (N_7436,N_75,N_2195);
or U7437 (N_7437,N_4008,N_2686);
nand U7438 (N_7438,N_2106,N_2299);
nand U7439 (N_7439,N_3806,N_1572);
xnor U7440 (N_7440,N_4833,N_264);
xnor U7441 (N_7441,N_2926,N_4214);
xnor U7442 (N_7442,N_2175,N_4328);
and U7443 (N_7443,N_1480,N_2541);
nand U7444 (N_7444,N_4955,N_2597);
nand U7445 (N_7445,N_3459,N_3924);
nor U7446 (N_7446,N_3160,N_2574);
nand U7447 (N_7447,N_2381,N_4967);
nand U7448 (N_7448,N_1483,N_4690);
nor U7449 (N_7449,N_1488,N_1419);
nor U7450 (N_7450,N_1033,N_4005);
nand U7451 (N_7451,N_4871,N_297);
xor U7452 (N_7452,N_4620,N_641);
or U7453 (N_7453,N_1685,N_682);
and U7454 (N_7454,N_1336,N_4838);
or U7455 (N_7455,N_2738,N_1714);
nand U7456 (N_7456,N_1412,N_2368);
nand U7457 (N_7457,N_333,N_4310);
and U7458 (N_7458,N_2773,N_2558);
nor U7459 (N_7459,N_3236,N_4906);
nand U7460 (N_7460,N_1126,N_3588);
nand U7461 (N_7461,N_4285,N_1536);
nor U7462 (N_7462,N_509,N_573);
and U7463 (N_7463,N_539,N_3695);
and U7464 (N_7464,N_2419,N_1355);
nor U7465 (N_7465,N_3329,N_4910);
and U7466 (N_7466,N_623,N_683);
nor U7467 (N_7467,N_4173,N_3137);
or U7468 (N_7468,N_3283,N_993);
and U7469 (N_7469,N_3275,N_1647);
nand U7470 (N_7470,N_1154,N_4228);
nor U7471 (N_7471,N_1270,N_139);
or U7472 (N_7472,N_3447,N_4561);
nand U7473 (N_7473,N_4947,N_4570);
nor U7474 (N_7474,N_4312,N_4730);
nand U7475 (N_7475,N_4430,N_1691);
or U7476 (N_7476,N_1950,N_4843);
nor U7477 (N_7477,N_3973,N_2058);
nand U7478 (N_7478,N_3118,N_2632);
nand U7479 (N_7479,N_3805,N_2174);
nor U7480 (N_7480,N_4249,N_4244);
nand U7481 (N_7481,N_1016,N_3467);
or U7482 (N_7482,N_2647,N_289);
nor U7483 (N_7483,N_2931,N_3195);
or U7484 (N_7484,N_1054,N_1139);
and U7485 (N_7485,N_232,N_3590);
nand U7486 (N_7486,N_817,N_3198);
or U7487 (N_7487,N_368,N_4668);
nand U7488 (N_7488,N_1581,N_1249);
and U7489 (N_7489,N_4629,N_3127);
nor U7490 (N_7490,N_3286,N_4977);
and U7491 (N_7491,N_4512,N_3573);
or U7492 (N_7492,N_1361,N_726);
and U7493 (N_7493,N_975,N_4554);
nand U7494 (N_7494,N_2018,N_4810);
and U7495 (N_7495,N_3962,N_2711);
and U7496 (N_7496,N_516,N_4982);
or U7497 (N_7497,N_1920,N_2366);
nor U7498 (N_7498,N_1461,N_4429);
nand U7499 (N_7499,N_595,N_532);
nor U7500 (N_7500,N_4497,N_1793);
or U7501 (N_7501,N_3278,N_3924);
nor U7502 (N_7502,N_2371,N_4513);
xor U7503 (N_7503,N_988,N_2729);
or U7504 (N_7504,N_3097,N_3372);
nor U7505 (N_7505,N_953,N_2755);
nand U7506 (N_7506,N_66,N_3063);
and U7507 (N_7507,N_3428,N_2511);
xnor U7508 (N_7508,N_415,N_1586);
nor U7509 (N_7509,N_4844,N_1766);
nand U7510 (N_7510,N_3897,N_2037);
nor U7511 (N_7511,N_4555,N_2248);
xnor U7512 (N_7512,N_4140,N_1046);
or U7513 (N_7513,N_3677,N_3224);
and U7514 (N_7514,N_4127,N_3585);
or U7515 (N_7515,N_470,N_3782);
nor U7516 (N_7516,N_4948,N_3815);
nor U7517 (N_7517,N_2224,N_3037);
or U7518 (N_7518,N_4142,N_4596);
and U7519 (N_7519,N_3405,N_1813);
nand U7520 (N_7520,N_3762,N_3200);
xor U7521 (N_7521,N_2048,N_1425);
xor U7522 (N_7522,N_3222,N_4995);
or U7523 (N_7523,N_823,N_674);
nor U7524 (N_7524,N_4613,N_1085);
nand U7525 (N_7525,N_3648,N_815);
or U7526 (N_7526,N_4719,N_3754);
xnor U7527 (N_7527,N_20,N_1455);
and U7528 (N_7528,N_3108,N_527);
nand U7529 (N_7529,N_2770,N_4746);
or U7530 (N_7530,N_3911,N_2296);
and U7531 (N_7531,N_3401,N_605);
and U7532 (N_7532,N_3742,N_426);
and U7533 (N_7533,N_4338,N_1060);
and U7534 (N_7534,N_1172,N_730);
nand U7535 (N_7535,N_1139,N_4345);
and U7536 (N_7536,N_2752,N_2809);
or U7537 (N_7537,N_260,N_710);
or U7538 (N_7538,N_4385,N_4594);
or U7539 (N_7539,N_4780,N_796);
nor U7540 (N_7540,N_3160,N_1736);
or U7541 (N_7541,N_2274,N_1589);
and U7542 (N_7542,N_2127,N_4481);
and U7543 (N_7543,N_1528,N_2791);
and U7544 (N_7544,N_153,N_2174);
nor U7545 (N_7545,N_1484,N_605);
nor U7546 (N_7546,N_318,N_3071);
nand U7547 (N_7547,N_1058,N_837);
nand U7548 (N_7548,N_2569,N_3580);
nor U7549 (N_7549,N_2031,N_2800);
nor U7550 (N_7550,N_4830,N_1798);
nand U7551 (N_7551,N_1090,N_2112);
nand U7552 (N_7552,N_4220,N_1730);
and U7553 (N_7553,N_3209,N_412);
nand U7554 (N_7554,N_1803,N_378);
nor U7555 (N_7555,N_1237,N_2291);
or U7556 (N_7556,N_4355,N_428);
nand U7557 (N_7557,N_4977,N_4491);
nor U7558 (N_7558,N_2008,N_3219);
or U7559 (N_7559,N_341,N_3745);
nand U7560 (N_7560,N_3750,N_2097);
xor U7561 (N_7561,N_4178,N_215);
nor U7562 (N_7562,N_1724,N_2575);
nand U7563 (N_7563,N_3087,N_1001);
nand U7564 (N_7564,N_3592,N_774);
or U7565 (N_7565,N_948,N_2430);
or U7566 (N_7566,N_320,N_815);
or U7567 (N_7567,N_836,N_1230);
nor U7568 (N_7568,N_2921,N_256);
xor U7569 (N_7569,N_1653,N_2609);
nor U7570 (N_7570,N_2729,N_2984);
xnor U7571 (N_7571,N_4583,N_885);
nor U7572 (N_7572,N_947,N_122);
and U7573 (N_7573,N_1481,N_1380);
nand U7574 (N_7574,N_4260,N_4340);
or U7575 (N_7575,N_4356,N_4788);
and U7576 (N_7576,N_81,N_1005);
nand U7577 (N_7577,N_763,N_1301);
or U7578 (N_7578,N_1720,N_3003);
and U7579 (N_7579,N_3265,N_2567);
nand U7580 (N_7580,N_824,N_2553);
and U7581 (N_7581,N_2691,N_2280);
nand U7582 (N_7582,N_578,N_1154);
and U7583 (N_7583,N_4423,N_1403);
or U7584 (N_7584,N_3756,N_4418);
nor U7585 (N_7585,N_436,N_4020);
nor U7586 (N_7586,N_342,N_2723);
nand U7587 (N_7587,N_2890,N_1181);
nor U7588 (N_7588,N_3060,N_3200);
or U7589 (N_7589,N_1539,N_1365);
and U7590 (N_7590,N_2579,N_779);
nor U7591 (N_7591,N_2788,N_3733);
and U7592 (N_7592,N_3013,N_1431);
or U7593 (N_7593,N_3629,N_276);
or U7594 (N_7594,N_2341,N_1379);
nand U7595 (N_7595,N_4062,N_670);
nor U7596 (N_7596,N_373,N_1157);
nand U7597 (N_7597,N_3485,N_4656);
and U7598 (N_7598,N_3928,N_2425);
nand U7599 (N_7599,N_2952,N_63);
nand U7600 (N_7600,N_1532,N_3028);
xnor U7601 (N_7601,N_4659,N_300);
nor U7602 (N_7602,N_3272,N_3667);
and U7603 (N_7603,N_1273,N_4260);
nor U7604 (N_7604,N_4328,N_3797);
nor U7605 (N_7605,N_1658,N_1364);
or U7606 (N_7606,N_214,N_1570);
nand U7607 (N_7607,N_3216,N_2526);
nand U7608 (N_7608,N_735,N_3263);
nand U7609 (N_7609,N_3340,N_2373);
or U7610 (N_7610,N_4878,N_1677);
and U7611 (N_7611,N_3616,N_3651);
nand U7612 (N_7612,N_1160,N_2051);
nor U7613 (N_7613,N_4261,N_1345);
and U7614 (N_7614,N_2776,N_1195);
nand U7615 (N_7615,N_3832,N_2633);
nand U7616 (N_7616,N_2118,N_3702);
nand U7617 (N_7617,N_4640,N_2981);
nand U7618 (N_7618,N_1363,N_2291);
nor U7619 (N_7619,N_2112,N_762);
or U7620 (N_7620,N_3008,N_2897);
nand U7621 (N_7621,N_1049,N_3357);
nand U7622 (N_7622,N_4234,N_4001);
and U7623 (N_7623,N_250,N_3401);
nand U7624 (N_7624,N_2796,N_1959);
nand U7625 (N_7625,N_3779,N_2442);
nand U7626 (N_7626,N_2629,N_1460);
nor U7627 (N_7627,N_4892,N_933);
or U7628 (N_7628,N_3471,N_2530);
nor U7629 (N_7629,N_3961,N_3122);
nor U7630 (N_7630,N_3952,N_4615);
and U7631 (N_7631,N_3159,N_2189);
or U7632 (N_7632,N_2715,N_3859);
nand U7633 (N_7633,N_3564,N_2643);
xnor U7634 (N_7634,N_3596,N_4168);
and U7635 (N_7635,N_456,N_1988);
nor U7636 (N_7636,N_623,N_3219);
nor U7637 (N_7637,N_1568,N_964);
nor U7638 (N_7638,N_4466,N_3701);
nand U7639 (N_7639,N_3484,N_4046);
or U7640 (N_7640,N_414,N_1165);
xor U7641 (N_7641,N_4627,N_4529);
nand U7642 (N_7642,N_820,N_1478);
nor U7643 (N_7643,N_4439,N_1258);
and U7644 (N_7644,N_447,N_17);
nand U7645 (N_7645,N_564,N_661);
nand U7646 (N_7646,N_4870,N_3919);
nand U7647 (N_7647,N_4997,N_315);
nor U7648 (N_7648,N_4338,N_4996);
nor U7649 (N_7649,N_3647,N_310);
nand U7650 (N_7650,N_2018,N_2223);
nor U7651 (N_7651,N_809,N_1405);
or U7652 (N_7652,N_313,N_2219);
or U7653 (N_7653,N_286,N_1379);
xor U7654 (N_7654,N_1526,N_390);
nor U7655 (N_7655,N_1614,N_1649);
nor U7656 (N_7656,N_1885,N_3644);
nor U7657 (N_7657,N_2540,N_1987);
or U7658 (N_7658,N_1710,N_4569);
nor U7659 (N_7659,N_2419,N_1708);
nor U7660 (N_7660,N_2247,N_4624);
nand U7661 (N_7661,N_2326,N_4012);
or U7662 (N_7662,N_854,N_1434);
nand U7663 (N_7663,N_298,N_338);
nor U7664 (N_7664,N_1747,N_1027);
and U7665 (N_7665,N_1056,N_1572);
or U7666 (N_7666,N_2586,N_3149);
or U7667 (N_7667,N_4248,N_3504);
or U7668 (N_7668,N_1031,N_4828);
and U7669 (N_7669,N_920,N_3119);
and U7670 (N_7670,N_775,N_989);
or U7671 (N_7671,N_294,N_63);
and U7672 (N_7672,N_708,N_3253);
or U7673 (N_7673,N_437,N_717);
nor U7674 (N_7674,N_2661,N_4328);
or U7675 (N_7675,N_410,N_3973);
and U7676 (N_7676,N_181,N_51);
nor U7677 (N_7677,N_2116,N_2375);
and U7678 (N_7678,N_2066,N_822);
nand U7679 (N_7679,N_4298,N_2321);
xor U7680 (N_7680,N_3850,N_4479);
or U7681 (N_7681,N_593,N_3386);
and U7682 (N_7682,N_4716,N_3304);
nor U7683 (N_7683,N_1124,N_3916);
or U7684 (N_7684,N_1531,N_4653);
or U7685 (N_7685,N_4071,N_466);
nor U7686 (N_7686,N_4621,N_2224);
and U7687 (N_7687,N_4113,N_777);
nor U7688 (N_7688,N_314,N_3611);
and U7689 (N_7689,N_2631,N_3295);
nand U7690 (N_7690,N_2801,N_2483);
xor U7691 (N_7691,N_2998,N_4389);
nor U7692 (N_7692,N_715,N_643);
nor U7693 (N_7693,N_1367,N_1390);
and U7694 (N_7694,N_128,N_2066);
xor U7695 (N_7695,N_4658,N_2126);
nor U7696 (N_7696,N_2175,N_3376);
nand U7697 (N_7697,N_3130,N_1429);
nand U7698 (N_7698,N_3425,N_612);
nor U7699 (N_7699,N_2809,N_230);
or U7700 (N_7700,N_2937,N_408);
or U7701 (N_7701,N_173,N_677);
nor U7702 (N_7702,N_3125,N_1340);
nor U7703 (N_7703,N_2309,N_1330);
xor U7704 (N_7704,N_2425,N_4738);
nand U7705 (N_7705,N_444,N_4327);
nand U7706 (N_7706,N_1228,N_569);
or U7707 (N_7707,N_3897,N_2720);
nand U7708 (N_7708,N_4687,N_3452);
or U7709 (N_7709,N_3340,N_302);
nor U7710 (N_7710,N_1929,N_862);
nand U7711 (N_7711,N_2984,N_2673);
and U7712 (N_7712,N_4764,N_1873);
nand U7713 (N_7713,N_1220,N_574);
nand U7714 (N_7714,N_4374,N_3941);
or U7715 (N_7715,N_4525,N_799);
nand U7716 (N_7716,N_4843,N_4063);
nand U7717 (N_7717,N_1678,N_3977);
nand U7718 (N_7718,N_449,N_3760);
xor U7719 (N_7719,N_3638,N_232);
xnor U7720 (N_7720,N_4272,N_4506);
nor U7721 (N_7721,N_4758,N_687);
or U7722 (N_7722,N_2517,N_1366);
and U7723 (N_7723,N_4961,N_4838);
or U7724 (N_7724,N_4715,N_3328);
nand U7725 (N_7725,N_2543,N_4081);
nor U7726 (N_7726,N_4780,N_1081);
and U7727 (N_7727,N_177,N_318);
nand U7728 (N_7728,N_4799,N_3668);
and U7729 (N_7729,N_2812,N_2111);
and U7730 (N_7730,N_124,N_1918);
nand U7731 (N_7731,N_1365,N_1165);
nor U7732 (N_7732,N_1009,N_555);
and U7733 (N_7733,N_1173,N_2243);
nand U7734 (N_7734,N_2735,N_3376);
or U7735 (N_7735,N_864,N_3742);
nand U7736 (N_7736,N_3799,N_2942);
nand U7737 (N_7737,N_3115,N_2837);
nand U7738 (N_7738,N_1620,N_3202);
nor U7739 (N_7739,N_4792,N_304);
nand U7740 (N_7740,N_3457,N_2559);
and U7741 (N_7741,N_2760,N_588);
and U7742 (N_7742,N_575,N_4807);
and U7743 (N_7743,N_2277,N_2488);
nand U7744 (N_7744,N_2100,N_348);
nand U7745 (N_7745,N_281,N_3593);
or U7746 (N_7746,N_4645,N_1228);
nor U7747 (N_7747,N_2796,N_1446);
nand U7748 (N_7748,N_2715,N_841);
nand U7749 (N_7749,N_1568,N_2185);
xor U7750 (N_7750,N_4601,N_2757);
nand U7751 (N_7751,N_981,N_1854);
nand U7752 (N_7752,N_3372,N_3954);
nor U7753 (N_7753,N_2871,N_3001);
nand U7754 (N_7754,N_949,N_1075);
or U7755 (N_7755,N_30,N_3673);
or U7756 (N_7756,N_4194,N_2348);
nor U7757 (N_7757,N_3202,N_1341);
nor U7758 (N_7758,N_660,N_4695);
xor U7759 (N_7759,N_1414,N_4239);
nand U7760 (N_7760,N_3796,N_1007);
and U7761 (N_7761,N_4031,N_4033);
and U7762 (N_7762,N_4666,N_4915);
and U7763 (N_7763,N_4800,N_903);
and U7764 (N_7764,N_4082,N_4851);
or U7765 (N_7765,N_4847,N_4039);
nor U7766 (N_7766,N_1565,N_3646);
nand U7767 (N_7767,N_2962,N_3847);
nor U7768 (N_7768,N_464,N_4440);
and U7769 (N_7769,N_1504,N_257);
xor U7770 (N_7770,N_636,N_2832);
and U7771 (N_7771,N_4190,N_2268);
nand U7772 (N_7772,N_2921,N_2688);
or U7773 (N_7773,N_1756,N_4649);
nand U7774 (N_7774,N_4223,N_4171);
nor U7775 (N_7775,N_2289,N_3401);
and U7776 (N_7776,N_1190,N_550);
nor U7777 (N_7777,N_6,N_48);
or U7778 (N_7778,N_3650,N_1919);
or U7779 (N_7779,N_4436,N_1139);
and U7780 (N_7780,N_3357,N_361);
or U7781 (N_7781,N_2442,N_2031);
nand U7782 (N_7782,N_1133,N_4663);
xnor U7783 (N_7783,N_1382,N_2425);
nand U7784 (N_7784,N_2627,N_4491);
nand U7785 (N_7785,N_2947,N_4266);
nor U7786 (N_7786,N_1460,N_4257);
nand U7787 (N_7787,N_2622,N_326);
nor U7788 (N_7788,N_2897,N_4859);
xor U7789 (N_7789,N_1169,N_1450);
and U7790 (N_7790,N_1017,N_4863);
xor U7791 (N_7791,N_1611,N_2379);
nand U7792 (N_7792,N_4089,N_3562);
xnor U7793 (N_7793,N_4328,N_3899);
nor U7794 (N_7794,N_2109,N_288);
and U7795 (N_7795,N_2131,N_3698);
nand U7796 (N_7796,N_3999,N_150);
or U7797 (N_7797,N_2370,N_1427);
xor U7798 (N_7798,N_4468,N_3593);
nor U7799 (N_7799,N_2058,N_442);
and U7800 (N_7800,N_1971,N_4226);
nand U7801 (N_7801,N_2042,N_3561);
nand U7802 (N_7802,N_24,N_4533);
and U7803 (N_7803,N_3089,N_4158);
nand U7804 (N_7804,N_82,N_3427);
and U7805 (N_7805,N_3497,N_4223);
and U7806 (N_7806,N_1650,N_3236);
or U7807 (N_7807,N_4275,N_4954);
nand U7808 (N_7808,N_2216,N_2215);
nand U7809 (N_7809,N_4997,N_2393);
and U7810 (N_7810,N_3194,N_4502);
nand U7811 (N_7811,N_431,N_944);
nor U7812 (N_7812,N_3171,N_242);
nand U7813 (N_7813,N_4206,N_3074);
or U7814 (N_7814,N_4331,N_2189);
nand U7815 (N_7815,N_261,N_2720);
or U7816 (N_7816,N_1731,N_2555);
nor U7817 (N_7817,N_4504,N_4774);
and U7818 (N_7818,N_1186,N_4582);
nor U7819 (N_7819,N_4253,N_1553);
nand U7820 (N_7820,N_1736,N_3061);
xnor U7821 (N_7821,N_4804,N_4913);
and U7822 (N_7822,N_2016,N_4212);
nor U7823 (N_7823,N_2647,N_796);
and U7824 (N_7824,N_1239,N_4954);
and U7825 (N_7825,N_628,N_1456);
and U7826 (N_7826,N_3009,N_2752);
nor U7827 (N_7827,N_3200,N_714);
nand U7828 (N_7828,N_2995,N_3322);
or U7829 (N_7829,N_2197,N_690);
xor U7830 (N_7830,N_1679,N_4479);
nor U7831 (N_7831,N_3598,N_4097);
and U7832 (N_7832,N_3736,N_2721);
nand U7833 (N_7833,N_249,N_3216);
nor U7834 (N_7834,N_4044,N_1111);
nor U7835 (N_7835,N_4882,N_2);
xor U7836 (N_7836,N_3525,N_4371);
or U7837 (N_7837,N_4417,N_1834);
xor U7838 (N_7838,N_2834,N_3305);
and U7839 (N_7839,N_3311,N_1902);
nand U7840 (N_7840,N_1856,N_3297);
nand U7841 (N_7841,N_2683,N_4027);
nand U7842 (N_7842,N_2046,N_1750);
nor U7843 (N_7843,N_2734,N_3579);
xor U7844 (N_7844,N_3672,N_4269);
and U7845 (N_7845,N_283,N_4896);
nand U7846 (N_7846,N_2017,N_2875);
nor U7847 (N_7847,N_4123,N_2393);
and U7848 (N_7848,N_4895,N_4106);
xor U7849 (N_7849,N_3706,N_613);
nand U7850 (N_7850,N_3961,N_1604);
or U7851 (N_7851,N_474,N_3917);
nor U7852 (N_7852,N_620,N_3334);
and U7853 (N_7853,N_752,N_3275);
nor U7854 (N_7854,N_3501,N_1595);
or U7855 (N_7855,N_2836,N_1983);
and U7856 (N_7856,N_3042,N_3603);
and U7857 (N_7857,N_2990,N_1573);
nor U7858 (N_7858,N_2693,N_1026);
nor U7859 (N_7859,N_1023,N_442);
or U7860 (N_7860,N_4040,N_672);
or U7861 (N_7861,N_3397,N_1227);
and U7862 (N_7862,N_2091,N_1081);
or U7863 (N_7863,N_3737,N_277);
and U7864 (N_7864,N_4846,N_1941);
nand U7865 (N_7865,N_4759,N_2873);
and U7866 (N_7866,N_4399,N_2398);
nor U7867 (N_7867,N_2519,N_11);
nor U7868 (N_7868,N_3128,N_416);
nor U7869 (N_7869,N_2909,N_4444);
or U7870 (N_7870,N_1211,N_902);
nor U7871 (N_7871,N_1901,N_4623);
or U7872 (N_7872,N_301,N_3158);
nor U7873 (N_7873,N_4426,N_3681);
and U7874 (N_7874,N_4861,N_3428);
and U7875 (N_7875,N_4413,N_3597);
or U7876 (N_7876,N_1922,N_2506);
or U7877 (N_7877,N_1040,N_4199);
xnor U7878 (N_7878,N_2992,N_765);
nand U7879 (N_7879,N_1674,N_484);
nand U7880 (N_7880,N_3073,N_2128);
and U7881 (N_7881,N_4863,N_1629);
and U7882 (N_7882,N_4332,N_4500);
nor U7883 (N_7883,N_772,N_3535);
or U7884 (N_7884,N_3870,N_3209);
or U7885 (N_7885,N_4517,N_3047);
nand U7886 (N_7886,N_133,N_4087);
nand U7887 (N_7887,N_2794,N_4533);
nand U7888 (N_7888,N_2647,N_337);
nor U7889 (N_7889,N_3861,N_2912);
xor U7890 (N_7890,N_3972,N_1224);
or U7891 (N_7891,N_1853,N_4911);
nand U7892 (N_7892,N_3791,N_413);
and U7893 (N_7893,N_3731,N_977);
xnor U7894 (N_7894,N_1455,N_4912);
nand U7895 (N_7895,N_3471,N_4866);
and U7896 (N_7896,N_4466,N_1874);
nand U7897 (N_7897,N_2535,N_2341);
nor U7898 (N_7898,N_4549,N_1956);
or U7899 (N_7899,N_648,N_855);
nor U7900 (N_7900,N_1486,N_678);
xnor U7901 (N_7901,N_4031,N_118);
and U7902 (N_7902,N_3331,N_3406);
xor U7903 (N_7903,N_4092,N_2014);
nor U7904 (N_7904,N_6,N_433);
nand U7905 (N_7905,N_2035,N_4368);
xor U7906 (N_7906,N_2091,N_516);
nor U7907 (N_7907,N_2909,N_1671);
nor U7908 (N_7908,N_3014,N_3701);
and U7909 (N_7909,N_3721,N_608);
xor U7910 (N_7910,N_3732,N_2274);
xor U7911 (N_7911,N_4136,N_2719);
or U7912 (N_7912,N_3990,N_2237);
nand U7913 (N_7913,N_1765,N_4148);
or U7914 (N_7914,N_518,N_4678);
nor U7915 (N_7915,N_2284,N_2709);
or U7916 (N_7916,N_2910,N_772);
and U7917 (N_7917,N_1008,N_1790);
and U7918 (N_7918,N_2011,N_3942);
nand U7919 (N_7919,N_2324,N_3610);
xor U7920 (N_7920,N_2896,N_3634);
nand U7921 (N_7921,N_3866,N_3552);
or U7922 (N_7922,N_1275,N_1145);
nor U7923 (N_7923,N_4517,N_251);
and U7924 (N_7924,N_4420,N_1591);
nand U7925 (N_7925,N_2148,N_3877);
nand U7926 (N_7926,N_1483,N_2068);
nand U7927 (N_7927,N_2175,N_4381);
nor U7928 (N_7928,N_4773,N_3221);
nor U7929 (N_7929,N_4559,N_1681);
or U7930 (N_7930,N_137,N_3893);
nor U7931 (N_7931,N_1362,N_2778);
and U7932 (N_7932,N_1519,N_1655);
nor U7933 (N_7933,N_1911,N_3159);
nand U7934 (N_7934,N_3124,N_3218);
or U7935 (N_7935,N_3476,N_1640);
or U7936 (N_7936,N_4787,N_2211);
nor U7937 (N_7937,N_2927,N_4731);
nor U7938 (N_7938,N_136,N_2160);
nand U7939 (N_7939,N_1622,N_4093);
xnor U7940 (N_7940,N_2889,N_2369);
xnor U7941 (N_7941,N_613,N_1929);
xor U7942 (N_7942,N_273,N_3260);
and U7943 (N_7943,N_4931,N_1459);
or U7944 (N_7944,N_3611,N_3364);
nand U7945 (N_7945,N_1292,N_3724);
or U7946 (N_7946,N_790,N_717);
and U7947 (N_7947,N_3100,N_3462);
or U7948 (N_7948,N_4783,N_485);
xor U7949 (N_7949,N_952,N_92);
xor U7950 (N_7950,N_1728,N_3704);
nor U7951 (N_7951,N_3864,N_3254);
or U7952 (N_7952,N_68,N_3297);
or U7953 (N_7953,N_3374,N_2033);
nor U7954 (N_7954,N_1926,N_4153);
nand U7955 (N_7955,N_2294,N_4782);
nand U7956 (N_7956,N_3840,N_1897);
xor U7957 (N_7957,N_2969,N_93);
nand U7958 (N_7958,N_2505,N_1264);
and U7959 (N_7959,N_457,N_365);
or U7960 (N_7960,N_4582,N_4943);
xor U7961 (N_7961,N_138,N_122);
and U7962 (N_7962,N_4560,N_4761);
nand U7963 (N_7963,N_1150,N_4007);
nor U7964 (N_7964,N_3664,N_1698);
or U7965 (N_7965,N_1441,N_3256);
or U7966 (N_7966,N_1360,N_1506);
and U7967 (N_7967,N_2340,N_4745);
and U7968 (N_7968,N_298,N_2829);
and U7969 (N_7969,N_3706,N_1533);
and U7970 (N_7970,N_4334,N_2536);
or U7971 (N_7971,N_3680,N_1055);
nand U7972 (N_7972,N_3299,N_2938);
or U7973 (N_7973,N_3137,N_4599);
nand U7974 (N_7974,N_4852,N_2044);
nor U7975 (N_7975,N_216,N_1184);
or U7976 (N_7976,N_2525,N_1099);
xor U7977 (N_7977,N_929,N_3342);
or U7978 (N_7978,N_3987,N_2809);
nor U7979 (N_7979,N_2510,N_4546);
nor U7980 (N_7980,N_3707,N_2937);
nand U7981 (N_7981,N_2907,N_2959);
nor U7982 (N_7982,N_1193,N_3362);
or U7983 (N_7983,N_1571,N_447);
and U7984 (N_7984,N_152,N_468);
and U7985 (N_7985,N_1258,N_3522);
nor U7986 (N_7986,N_3946,N_2332);
nand U7987 (N_7987,N_2486,N_79);
and U7988 (N_7988,N_1834,N_1808);
nor U7989 (N_7989,N_2698,N_2313);
or U7990 (N_7990,N_934,N_2959);
or U7991 (N_7991,N_520,N_4209);
or U7992 (N_7992,N_2756,N_815);
and U7993 (N_7993,N_4676,N_2956);
and U7994 (N_7994,N_2921,N_3016);
or U7995 (N_7995,N_1203,N_3802);
and U7996 (N_7996,N_60,N_1341);
xor U7997 (N_7997,N_4082,N_3663);
nand U7998 (N_7998,N_4525,N_3646);
nor U7999 (N_7999,N_2320,N_4983);
nand U8000 (N_8000,N_3040,N_4901);
nor U8001 (N_8001,N_1162,N_2184);
nand U8002 (N_8002,N_1325,N_2444);
or U8003 (N_8003,N_2284,N_297);
or U8004 (N_8004,N_2316,N_2199);
nand U8005 (N_8005,N_81,N_4306);
nand U8006 (N_8006,N_2663,N_5);
or U8007 (N_8007,N_4972,N_3176);
nand U8008 (N_8008,N_2114,N_4497);
nor U8009 (N_8009,N_2054,N_1710);
or U8010 (N_8010,N_1225,N_3800);
and U8011 (N_8011,N_1869,N_1019);
nand U8012 (N_8012,N_4654,N_582);
xor U8013 (N_8013,N_1884,N_2405);
nor U8014 (N_8014,N_3830,N_4227);
and U8015 (N_8015,N_600,N_3752);
xnor U8016 (N_8016,N_4712,N_2849);
nand U8017 (N_8017,N_933,N_1975);
and U8018 (N_8018,N_4111,N_2225);
nand U8019 (N_8019,N_4346,N_4112);
or U8020 (N_8020,N_3915,N_3230);
xnor U8021 (N_8021,N_4033,N_242);
or U8022 (N_8022,N_2418,N_4348);
nor U8023 (N_8023,N_4350,N_2163);
or U8024 (N_8024,N_1907,N_2235);
nand U8025 (N_8025,N_3112,N_2069);
nand U8026 (N_8026,N_1420,N_4809);
or U8027 (N_8027,N_335,N_924);
nor U8028 (N_8028,N_4963,N_651);
xor U8029 (N_8029,N_2752,N_389);
and U8030 (N_8030,N_2474,N_2382);
and U8031 (N_8031,N_1933,N_4716);
and U8032 (N_8032,N_643,N_3311);
nand U8033 (N_8033,N_369,N_2959);
xnor U8034 (N_8034,N_953,N_2844);
nor U8035 (N_8035,N_1332,N_1657);
nor U8036 (N_8036,N_4001,N_393);
and U8037 (N_8037,N_1654,N_361);
or U8038 (N_8038,N_3349,N_1406);
nand U8039 (N_8039,N_3597,N_4825);
and U8040 (N_8040,N_2273,N_3873);
or U8041 (N_8041,N_4669,N_3303);
nor U8042 (N_8042,N_11,N_1394);
nand U8043 (N_8043,N_3700,N_4673);
or U8044 (N_8044,N_3857,N_273);
xnor U8045 (N_8045,N_1347,N_3222);
and U8046 (N_8046,N_865,N_2399);
nand U8047 (N_8047,N_4884,N_2327);
nor U8048 (N_8048,N_4519,N_3756);
or U8049 (N_8049,N_1839,N_714);
xor U8050 (N_8050,N_4582,N_4336);
and U8051 (N_8051,N_3892,N_2673);
or U8052 (N_8052,N_4154,N_384);
xor U8053 (N_8053,N_4764,N_1910);
and U8054 (N_8054,N_2600,N_1762);
nor U8055 (N_8055,N_1794,N_364);
nor U8056 (N_8056,N_4890,N_3128);
or U8057 (N_8057,N_3568,N_3683);
or U8058 (N_8058,N_124,N_4194);
or U8059 (N_8059,N_4640,N_795);
nand U8060 (N_8060,N_4065,N_2351);
or U8061 (N_8061,N_4995,N_2894);
or U8062 (N_8062,N_3171,N_285);
nor U8063 (N_8063,N_911,N_2706);
and U8064 (N_8064,N_3298,N_481);
and U8065 (N_8065,N_559,N_2788);
nand U8066 (N_8066,N_3398,N_2645);
and U8067 (N_8067,N_2378,N_836);
nor U8068 (N_8068,N_4539,N_4195);
and U8069 (N_8069,N_1187,N_3285);
xnor U8070 (N_8070,N_739,N_3576);
and U8071 (N_8071,N_83,N_187);
xor U8072 (N_8072,N_4513,N_897);
nor U8073 (N_8073,N_1770,N_2979);
and U8074 (N_8074,N_493,N_1501);
or U8075 (N_8075,N_1111,N_2918);
or U8076 (N_8076,N_4079,N_3913);
and U8077 (N_8077,N_4685,N_1564);
xor U8078 (N_8078,N_1503,N_3540);
or U8079 (N_8079,N_1167,N_3172);
xnor U8080 (N_8080,N_4565,N_4846);
and U8081 (N_8081,N_1514,N_117);
nor U8082 (N_8082,N_4250,N_3330);
or U8083 (N_8083,N_2709,N_3066);
nand U8084 (N_8084,N_2077,N_3601);
nor U8085 (N_8085,N_914,N_3541);
xor U8086 (N_8086,N_2808,N_2320);
nor U8087 (N_8087,N_749,N_762);
xnor U8088 (N_8088,N_1099,N_1944);
nand U8089 (N_8089,N_1370,N_3433);
nor U8090 (N_8090,N_1065,N_862);
xor U8091 (N_8091,N_2244,N_2799);
or U8092 (N_8092,N_146,N_3406);
or U8093 (N_8093,N_3095,N_3182);
nor U8094 (N_8094,N_830,N_469);
and U8095 (N_8095,N_1251,N_4512);
nor U8096 (N_8096,N_3988,N_852);
nand U8097 (N_8097,N_4550,N_427);
or U8098 (N_8098,N_806,N_658);
xor U8099 (N_8099,N_4216,N_2105);
and U8100 (N_8100,N_2810,N_3062);
nand U8101 (N_8101,N_3776,N_1747);
or U8102 (N_8102,N_2384,N_273);
nor U8103 (N_8103,N_1532,N_841);
xor U8104 (N_8104,N_1523,N_2233);
nand U8105 (N_8105,N_324,N_3533);
nand U8106 (N_8106,N_1024,N_1122);
and U8107 (N_8107,N_3489,N_513);
or U8108 (N_8108,N_2739,N_2538);
or U8109 (N_8109,N_1028,N_3104);
nand U8110 (N_8110,N_416,N_704);
or U8111 (N_8111,N_3241,N_1946);
nor U8112 (N_8112,N_4106,N_4984);
nor U8113 (N_8113,N_10,N_1138);
nand U8114 (N_8114,N_803,N_2967);
xnor U8115 (N_8115,N_1220,N_3655);
nor U8116 (N_8116,N_640,N_681);
or U8117 (N_8117,N_742,N_2381);
xnor U8118 (N_8118,N_3656,N_1009);
and U8119 (N_8119,N_2929,N_415);
nand U8120 (N_8120,N_3953,N_791);
nand U8121 (N_8121,N_3733,N_3095);
nor U8122 (N_8122,N_2673,N_173);
xor U8123 (N_8123,N_1595,N_1989);
and U8124 (N_8124,N_2732,N_767);
or U8125 (N_8125,N_2953,N_3574);
nand U8126 (N_8126,N_1674,N_2462);
nor U8127 (N_8127,N_1290,N_846);
nor U8128 (N_8128,N_2696,N_521);
or U8129 (N_8129,N_27,N_3101);
or U8130 (N_8130,N_252,N_4782);
nand U8131 (N_8131,N_2684,N_2981);
or U8132 (N_8132,N_4566,N_609);
or U8133 (N_8133,N_2350,N_1155);
nand U8134 (N_8134,N_3709,N_1705);
nand U8135 (N_8135,N_2681,N_4685);
nand U8136 (N_8136,N_3377,N_4429);
or U8137 (N_8137,N_2596,N_2847);
and U8138 (N_8138,N_2109,N_3430);
and U8139 (N_8139,N_2033,N_3378);
nor U8140 (N_8140,N_4515,N_1394);
nand U8141 (N_8141,N_1801,N_754);
nor U8142 (N_8142,N_4187,N_4871);
nand U8143 (N_8143,N_131,N_322);
xor U8144 (N_8144,N_4129,N_4788);
xnor U8145 (N_8145,N_2258,N_1066);
nand U8146 (N_8146,N_926,N_2520);
or U8147 (N_8147,N_4522,N_4457);
or U8148 (N_8148,N_3586,N_1990);
or U8149 (N_8149,N_2823,N_1447);
or U8150 (N_8150,N_3085,N_2557);
nor U8151 (N_8151,N_2478,N_2667);
and U8152 (N_8152,N_2639,N_1306);
or U8153 (N_8153,N_4138,N_1256);
or U8154 (N_8154,N_4017,N_3480);
nor U8155 (N_8155,N_616,N_3434);
nand U8156 (N_8156,N_396,N_3155);
nand U8157 (N_8157,N_2908,N_534);
nor U8158 (N_8158,N_3099,N_4707);
and U8159 (N_8159,N_2608,N_952);
and U8160 (N_8160,N_3471,N_1981);
nor U8161 (N_8161,N_2566,N_96);
nand U8162 (N_8162,N_1450,N_865);
and U8163 (N_8163,N_3264,N_226);
nand U8164 (N_8164,N_3147,N_4102);
nand U8165 (N_8165,N_249,N_4468);
and U8166 (N_8166,N_1085,N_2156);
or U8167 (N_8167,N_306,N_352);
nor U8168 (N_8168,N_1518,N_4868);
nand U8169 (N_8169,N_1242,N_4309);
or U8170 (N_8170,N_605,N_4046);
nand U8171 (N_8171,N_506,N_2104);
nand U8172 (N_8172,N_714,N_2931);
or U8173 (N_8173,N_978,N_1145);
and U8174 (N_8174,N_4299,N_2800);
nor U8175 (N_8175,N_3797,N_720);
nand U8176 (N_8176,N_3245,N_698);
or U8177 (N_8177,N_4214,N_2709);
nand U8178 (N_8178,N_4853,N_2206);
or U8179 (N_8179,N_1288,N_3363);
nor U8180 (N_8180,N_3905,N_1356);
or U8181 (N_8181,N_4791,N_3346);
xnor U8182 (N_8182,N_3645,N_2317);
nand U8183 (N_8183,N_3145,N_1061);
nand U8184 (N_8184,N_561,N_2088);
nand U8185 (N_8185,N_1795,N_4220);
nand U8186 (N_8186,N_3215,N_3011);
nor U8187 (N_8187,N_1534,N_3775);
xor U8188 (N_8188,N_238,N_4077);
nor U8189 (N_8189,N_3440,N_3209);
nor U8190 (N_8190,N_3465,N_3096);
and U8191 (N_8191,N_3066,N_1375);
nand U8192 (N_8192,N_501,N_1583);
and U8193 (N_8193,N_3014,N_3480);
nand U8194 (N_8194,N_4177,N_3565);
or U8195 (N_8195,N_1549,N_3718);
or U8196 (N_8196,N_2253,N_3086);
nand U8197 (N_8197,N_4221,N_2637);
xnor U8198 (N_8198,N_1443,N_1662);
nor U8199 (N_8199,N_4591,N_494);
nor U8200 (N_8200,N_2863,N_3600);
xor U8201 (N_8201,N_3801,N_3718);
and U8202 (N_8202,N_520,N_4342);
nor U8203 (N_8203,N_1725,N_1574);
nand U8204 (N_8204,N_3997,N_3740);
xnor U8205 (N_8205,N_2309,N_4571);
xor U8206 (N_8206,N_528,N_4358);
nor U8207 (N_8207,N_3164,N_4788);
nor U8208 (N_8208,N_1578,N_1616);
or U8209 (N_8209,N_1125,N_4696);
or U8210 (N_8210,N_4207,N_3101);
nand U8211 (N_8211,N_4706,N_1819);
nand U8212 (N_8212,N_3789,N_4156);
nor U8213 (N_8213,N_1,N_2620);
and U8214 (N_8214,N_2118,N_1376);
xor U8215 (N_8215,N_1917,N_2374);
and U8216 (N_8216,N_4213,N_4617);
nor U8217 (N_8217,N_1050,N_3290);
or U8218 (N_8218,N_2816,N_3266);
and U8219 (N_8219,N_2096,N_4841);
nor U8220 (N_8220,N_4602,N_1135);
nand U8221 (N_8221,N_3536,N_1678);
and U8222 (N_8222,N_4419,N_2196);
nand U8223 (N_8223,N_704,N_4484);
xor U8224 (N_8224,N_2302,N_1637);
nand U8225 (N_8225,N_206,N_1510);
and U8226 (N_8226,N_4598,N_862);
or U8227 (N_8227,N_2230,N_2722);
nand U8228 (N_8228,N_4330,N_2742);
nor U8229 (N_8229,N_1569,N_314);
nand U8230 (N_8230,N_849,N_3832);
and U8231 (N_8231,N_958,N_850);
nand U8232 (N_8232,N_706,N_4990);
xnor U8233 (N_8233,N_1191,N_2921);
nand U8234 (N_8234,N_2641,N_1292);
nand U8235 (N_8235,N_2687,N_4185);
nor U8236 (N_8236,N_6,N_1398);
xnor U8237 (N_8237,N_3117,N_1610);
and U8238 (N_8238,N_3350,N_2426);
or U8239 (N_8239,N_3251,N_417);
nor U8240 (N_8240,N_971,N_216);
nor U8241 (N_8241,N_1318,N_822);
nand U8242 (N_8242,N_1702,N_3053);
or U8243 (N_8243,N_2916,N_429);
nand U8244 (N_8244,N_2732,N_4836);
and U8245 (N_8245,N_3392,N_4116);
or U8246 (N_8246,N_918,N_628);
nor U8247 (N_8247,N_334,N_687);
and U8248 (N_8248,N_1126,N_2307);
nand U8249 (N_8249,N_4543,N_4245);
nor U8250 (N_8250,N_2601,N_35);
nor U8251 (N_8251,N_1617,N_488);
and U8252 (N_8252,N_4304,N_1074);
nor U8253 (N_8253,N_2946,N_2320);
nor U8254 (N_8254,N_4532,N_4232);
nand U8255 (N_8255,N_3308,N_3239);
or U8256 (N_8256,N_2431,N_41);
nand U8257 (N_8257,N_3122,N_412);
and U8258 (N_8258,N_1793,N_2742);
nor U8259 (N_8259,N_1837,N_1053);
xor U8260 (N_8260,N_33,N_3548);
nor U8261 (N_8261,N_3428,N_1589);
nor U8262 (N_8262,N_944,N_4806);
or U8263 (N_8263,N_3025,N_2461);
nor U8264 (N_8264,N_86,N_3469);
or U8265 (N_8265,N_3436,N_484);
nor U8266 (N_8266,N_2782,N_3385);
nand U8267 (N_8267,N_4183,N_3573);
or U8268 (N_8268,N_2977,N_513);
nand U8269 (N_8269,N_4187,N_2832);
nand U8270 (N_8270,N_597,N_3944);
nor U8271 (N_8271,N_2116,N_598);
xnor U8272 (N_8272,N_687,N_2883);
and U8273 (N_8273,N_3617,N_1990);
nand U8274 (N_8274,N_4247,N_314);
nor U8275 (N_8275,N_2642,N_1621);
nor U8276 (N_8276,N_2260,N_2424);
or U8277 (N_8277,N_1329,N_3654);
and U8278 (N_8278,N_3386,N_1074);
nor U8279 (N_8279,N_3453,N_2659);
and U8280 (N_8280,N_4924,N_2754);
and U8281 (N_8281,N_1704,N_4498);
and U8282 (N_8282,N_1674,N_3291);
and U8283 (N_8283,N_1436,N_3825);
nand U8284 (N_8284,N_4483,N_2008);
or U8285 (N_8285,N_3686,N_3252);
nor U8286 (N_8286,N_2863,N_411);
and U8287 (N_8287,N_2463,N_2341);
nand U8288 (N_8288,N_3508,N_3484);
nand U8289 (N_8289,N_4465,N_391);
nor U8290 (N_8290,N_1568,N_3290);
and U8291 (N_8291,N_2897,N_960);
and U8292 (N_8292,N_2902,N_1940);
and U8293 (N_8293,N_2238,N_2539);
nor U8294 (N_8294,N_4679,N_2845);
or U8295 (N_8295,N_54,N_3740);
or U8296 (N_8296,N_3508,N_1025);
nand U8297 (N_8297,N_3063,N_3757);
nand U8298 (N_8298,N_2815,N_1014);
nand U8299 (N_8299,N_2642,N_1059);
xnor U8300 (N_8300,N_1292,N_278);
and U8301 (N_8301,N_4138,N_3972);
and U8302 (N_8302,N_3998,N_751);
or U8303 (N_8303,N_3594,N_3689);
or U8304 (N_8304,N_1638,N_1063);
or U8305 (N_8305,N_1774,N_140);
or U8306 (N_8306,N_1827,N_2025);
nor U8307 (N_8307,N_2410,N_3632);
or U8308 (N_8308,N_280,N_3924);
xnor U8309 (N_8309,N_2157,N_3006);
or U8310 (N_8310,N_2423,N_4839);
nor U8311 (N_8311,N_2402,N_2507);
nand U8312 (N_8312,N_1987,N_2313);
or U8313 (N_8313,N_3767,N_4434);
nor U8314 (N_8314,N_4815,N_4642);
nand U8315 (N_8315,N_906,N_4434);
nor U8316 (N_8316,N_1564,N_4942);
nor U8317 (N_8317,N_2669,N_2075);
nand U8318 (N_8318,N_2053,N_1491);
nand U8319 (N_8319,N_2185,N_2408);
or U8320 (N_8320,N_2568,N_4868);
and U8321 (N_8321,N_1026,N_3351);
nor U8322 (N_8322,N_1086,N_1988);
nor U8323 (N_8323,N_3685,N_4949);
nand U8324 (N_8324,N_3096,N_3639);
and U8325 (N_8325,N_4506,N_135);
nor U8326 (N_8326,N_2046,N_1567);
xor U8327 (N_8327,N_3171,N_4915);
nand U8328 (N_8328,N_2718,N_3264);
nor U8329 (N_8329,N_1506,N_557);
xor U8330 (N_8330,N_2470,N_47);
or U8331 (N_8331,N_1630,N_2991);
and U8332 (N_8332,N_4626,N_920);
or U8333 (N_8333,N_329,N_2071);
and U8334 (N_8334,N_3955,N_1450);
nand U8335 (N_8335,N_1497,N_1013);
nand U8336 (N_8336,N_3348,N_810);
xor U8337 (N_8337,N_250,N_727);
and U8338 (N_8338,N_423,N_519);
nor U8339 (N_8339,N_2603,N_1925);
and U8340 (N_8340,N_3409,N_330);
nor U8341 (N_8341,N_2899,N_404);
nand U8342 (N_8342,N_1592,N_3963);
nor U8343 (N_8343,N_1119,N_1822);
nor U8344 (N_8344,N_122,N_2529);
and U8345 (N_8345,N_3133,N_4056);
and U8346 (N_8346,N_1586,N_2439);
nor U8347 (N_8347,N_4157,N_243);
nand U8348 (N_8348,N_2214,N_1200);
nor U8349 (N_8349,N_1565,N_671);
nand U8350 (N_8350,N_3859,N_130);
or U8351 (N_8351,N_3012,N_4172);
or U8352 (N_8352,N_1408,N_3954);
nor U8353 (N_8353,N_3096,N_2642);
nand U8354 (N_8354,N_540,N_4083);
and U8355 (N_8355,N_4145,N_3824);
nand U8356 (N_8356,N_2487,N_138);
and U8357 (N_8357,N_4964,N_3133);
nor U8358 (N_8358,N_246,N_1853);
xor U8359 (N_8359,N_4781,N_1287);
and U8360 (N_8360,N_3348,N_1398);
xnor U8361 (N_8361,N_502,N_3309);
or U8362 (N_8362,N_4899,N_407);
or U8363 (N_8363,N_4087,N_321);
xor U8364 (N_8364,N_4614,N_963);
and U8365 (N_8365,N_1270,N_575);
or U8366 (N_8366,N_1604,N_4280);
nor U8367 (N_8367,N_837,N_885);
or U8368 (N_8368,N_210,N_3157);
nand U8369 (N_8369,N_63,N_4271);
and U8370 (N_8370,N_779,N_3844);
and U8371 (N_8371,N_4088,N_3872);
and U8372 (N_8372,N_3654,N_4964);
nand U8373 (N_8373,N_4724,N_424);
or U8374 (N_8374,N_4846,N_3582);
nand U8375 (N_8375,N_4940,N_4742);
nor U8376 (N_8376,N_4023,N_1356);
nor U8377 (N_8377,N_1231,N_677);
nor U8378 (N_8378,N_2561,N_4279);
or U8379 (N_8379,N_4374,N_2821);
nor U8380 (N_8380,N_1289,N_1715);
xor U8381 (N_8381,N_625,N_255);
or U8382 (N_8382,N_3951,N_4554);
or U8383 (N_8383,N_599,N_2137);
and U8384 (N_8384,N_2742,N_216);
or U8385 (N_8385,N_2688,N_2941);
and U8386 (N_8386,N_1380,N_1143);
and U8387 (N_8387,N_1807,N_2184);
nand U8388 (N_8388,N_3906,N_4102);
nand U8389 (N_8389,N_630,N_67);
and U8390 (N_8390,N_2057,N_3734);
or U8391 (N_8391,N_144,N_3963);
nor U8392 (N_8392,N_1049,N_523);
or U8393 (N_8393,N_2965,N_38);
nand U8394 (N_8394,N_1805,N_1657);
nand U8395 (N_8395,N_4881,N_1183);
and U8396 (N_8396,N_2872,N_4031);
nand U8397 (N_8397,N_2454,N_4490);
or U8398 (N_8398,N_4150,N_988);
nand U8399 (N_8399,N_4757,N_2662);
nor U8400 (N_8400,N_4954,N_2286);
and U8401 (N_8401,N_1335,N_778);
or U8402 (N_8402,N_3532,N_166);
or U8403 (N_8403,N_1404,N_1550);
or U8404 (N_8404,N_1441,N_250);
and U8405 (N_8405,N_3125,N_3736);
and U8406 (N_8406,N_2918,N_3643);
or U8407 (N_8407,N_3113,N_105);
and U8408 (N_8408,N_1892,N_3299);
or U8409 (N_8409,N_3171,N_252);
and U8410 (N_8410,N_3059,N_1660);
nand U8411 (N_8411,N_783,N_2140);
nor U8412 (N_8412,N_497,N_2994);
nand U8413 (N_8413,N_1819,N_1873);
and U8414 (N_8414,N_3252,N_874);
or U8415 (N_8415,N_4315,N_2697);
nor U8416 (N_8416,N_3714,N_203);
or U8417 (N_8417,N_4499,N_109);
nand U8418 (N_8418,N_4603,N_1526);
nand U8419 (N_8419,N_1266,N_213);
or U8420 (N_8420,N_4009,N_3097);
and U8421 (N_8421,N_4392,N_4564);
nand U8422 (N_8422,N_2214,N_717);
nor U8423 (N_8423,N_3770,N_4527);
and U8424 (N_8424,N_4590,N_3163);
nor U8425 (N_8425,N_342,N_237);
and U8426 (N_8426,N_1337,N_2400);
nor U8427 (N_8427,N_4888,N_1316);
nand U8428 (N_8428,N_868,N_0);
nand U8429 (N_8429,N_4206,N_1801);
and U8430 (N_8430,N_2669,N_98);
nor U8431 (N_8431,N_3753,N_4048);
nor U8432 (N_8432,N_1561,N_539);
nand U8433 (N_8433,N_406,N_777);
and U8434 (N_8434,N_81,N_3137);
nand U8435 (N_8435,N_1957,N_749);
xor U8436 (N_8436,N_519,N_3671);
or U8437 (N_8437,N_3826,N_4248);
xor U8438 (N_8438,N_948,N_851);
nor U8439 (N_8439,N_1886,N_1519);
nor U8440 (N_8440,N_4835,N_1430);
and U8441 (N_8441,N_2191,N_3350);
nand U8442 (N_8442,N_1317,N_3565);
and U8443 (N_8443,N_4093,N_2810);
nand U8444 (N_8444,N_649,N_4988);
xnor U8445 (N_8445,N_3877,N_4657);
or U8446 (N_8446,N_965,N_3335);
and U8447 (N_8447,N_406,N_3787);
nor U8448 (N_8448,N_4780,N_4836);
nor U8449 (N_8449,N_2671,N_4486);
and U8450 (N_8450,N_4216,N_2909);
nor U8451 (N_8451,N_4994,N_3231);
or U8452 (N_8452,N_3701,N_4514);
and U8453 (N_8453,N_2017,N_3148);
nor U8454 (N_8454,N_1927,N_272);
nand U8455 (N_8455,N_3682,N_1393);
nor U8456 (N_8456,N_2563,N_3886);
nor U8457 (N_8457,N_1837,N_3970);
nand U8458 (N_8458,N_1099,N_4225);
nand U8459 (N_8459,N_2987,N_4096);
and U8460 (N_8460,N_3437,N_1833);
and U8461 (N_8461,N_62,N_1785);
or U8462 (N_8462,N_677,N_4678);
nand U8463 (N_8463,N_2522,N_3843);
and U8464 (N_8464,N_1072,N_3732);
and U8465 (N_8465,N_2161,N_4199);
nand U8466 (N_8466,N_313,N_3458);
nor U8467 (N_8467,N_1151,N_4708);
nand U8468 (N_8468,N_2489,N_4213);
nand U8469 (N_8469,N_4892,N_187);
or U8470 (N_8470,N_2463,N_3623);
and U8471 (N_8471,N_93,N_1605);
or U8472 (N_8472,N_3437,N_1111);
or U8473 (N_8473,N_4790,N_1453);
and U8474 (N_8474,N_1856,N_3004);
nor U8475 (N_8475,N_4104,N_1147);
nor U8476 (N_8476,N_3358,N_2571);
and U8477 (N_8477,N_1316,N_4085);
or U8478 (N_8478,N_4499,N_1818);
nand U8479 (N_8479,N_2386,N_348);
nor U8480 (N_8480,N_2094,N_3576);
nand U8481 (N_8481,N_3752,N_5);
and U8482 (N_8482,N_4658,N_3522);
nor U8483 (N_8483,N_86,N_2268);
nand U8484 (N_8484,N_3940,N_987);
nand U8485 (N_8485,N_487,N_956);
nand U8486 (N_8486,N_2189,N_2790);
and U8487 (N_8487,N_671,N_168);
nor U8488 (N_8488,N_2684,N_4575);
or U8489 (N_8489,N_3734,N_678);
nor U8490 (N_8490,N_2584,N_3225);
nand U8491 (N_8491,N_535,N_1564);
nand U8492 (N_8492,N_194,N_496);
nor U8493 (N_8493,N_3092,N_4658);
nand U8494 (N_8494,N_3798,N_3648);
or U8495 (N_8495,N_1998,N_2302);
or U8496 (N_8496,N_1263,N_1372);
nor U8497 (N_8497,N_721,N_4970);
nand U8498 (N_8498,N_995,N_1154);
or U8499 (N_8499,N_2902,N_1032);
nand U8500 (N_8500,N_4336,N_2905);
nor U8501 (N_8501,N_2402,N_1224);
or U8502 (N_8502,N_1268,N_435);
nor U8503 (N_8503,N_2392,N_4334);
and U8504 (N_8504,N_2852,N_1512);
nor U8505 (N_8505,N_3179,N_2402);
nor U8506 (N_8506,N_2200,N_3433);
xnor U8507 (N_8507,N_599,N_3423);
and U8508 (N_8508,N_3257,N_2026);
and U8509 (N_8509,N_2955,N_2167);
and U8510 (N_8510,N_2377,N_776);
or U8511 (N_8511,N_4250,N_727);
nand U8512 (N_8512,N_1685,N_149);
and U8513 (N_8513,N_2561,N_1504);
xor U8514 (N_8514,N_4235,N_775);
xnor U8515 (N_8515,N_2884,N_1336);
nor U8516 (N_8516,N_958,N_53);
nand U8517 (N_8517,N_3832,N_1259);
or U8518 (N_8518,N_4521,N_515);
nand U8519 (N_8519,N_3491,N_2052);
nor U8520 (N_8520,N_4949,N_3933);
and U8521 (N_8521,N_1566,N_3622);
and U8522 (N_8522,N_1184,N_4455);
xor U8523 (N_8523,N_972,N_1644);
xnor U8524 (N_8524,N_4997,N_3069);
and U8525 (N_8525,N_216,N_895);
and U8526 (N_8526,N_4127,N_3622);
nand U8527 (N_8527,N_2274,N_1433);
or U8528 (N_8528,N_375,N_3377);
or U8529 (N_8529,N_1364,N_4995);
or U8530 (N_8530,N_3115,N_994);
nand U8531 (N_8531,N_514,N_1284);
nor U8532 (N_8532,N_2806,N_3966);
xor U8533 (N_8533,N_3421,N_2343);
and U8534 (N_8534,N_3067,N_4130);
nand U8535 (N_8535,N_3938,N_1868);
nand U8536 (N_8536,N_3450,N_1422);
xor U8537 (N_8537,N_4468,N_2569);
nand U8538 (N_8538,N_4372,N_3812);
and U8539 (N_8539,N_702,N_1709);
xnor U8540 (N_8540,N_4989,N_4556);
nor U8541 (N_8541,N_2985,N_3044);
and U8542 (N_8542,N_302,N_4146);
and U8543 (N_8543,N_4726,N_2479);
nand U8544 (N_8544,N_2410,N_1679);
nor U8545 (N_8545,N_4803,N_389);
nand U8546 (N_8546,N_3690,N_1840);
or U8547 (N_8547,N_1776,N_1118);
and U8548 (N_8548,N_1824,N_4142);
and U8549 (N_8549,N_2688,N_2946);
xor U8550 (N_8550,N_2013,N_4768);
nand U8551 (N_8551,N_1535,N_2985);
nor U8552 (N_8552,N_2202,N_2907);
nand U8553 (N_8553,N_1607,N_4846);
and U8554 (N_8554,N_2131,N_1526);
nand U8555 (N_8555,N_3273,N_3737);
or U8556 (N_8556,N_1884,N_3251);
and U8557 (N_8557,N_3630,N_4877);
and U8558 (N_8558,N_4951,N_2065);
or U8559 (N_8559,N_3831,N_1070);
or U8560 (N_8560,N_2029,N_4366);
xor U8561 (N_8561,N_1259,N_3178);
and U8562 (N_8562,N_2014,N_4435);
and U8563 (N_8563,N_1790,N_1954);
and U8564 (N_8564,N_4166,N_1530);
nand U8565 (N_8565,N_2304,N_2609);
nand U8566 (N_8566,N_307,N_4386);
and U8567 (N_8567,N_683,N_4680);
nor U8568 (N_8568,N_3985,N_1627);
or U8569 (N_8569,N_181,N_2057);
and U8570 (N_8570,N_2486,N_2425);
xor U8571 (N_8571,N_2564,N_3776);
nand U8572 (N_8572,N_2913,N_2248);
or U8573 (N_8573,N_3840,N_499);
and U8574 (N_8574,N_1760,N_2876);
and U8575 (N_8575,N_115,N_1104);
or U8576 (N_8576,N_468,N_4121);
nor U8577 (N_8577,N_2618,N_1643);
nor U8578 (N_8578,N_3089,N_871);
and U8579 (N_8579,N_1073,N_576);
or U8580 (N_8580,N_947,N_4839);
or U8581 (N_8581,N_1133,N_3783);
and U8582 (N_8582,N_2352,N_4296);
nor U8583 (N_8583,N_2753,N_4233);
and U8584 (N_8584,N_788,N_3852);
or U8585 (N_8585,N_3306,N_1195);
or U8586 (N_8586,N_1546,N_436);
xnor U8587 (N_8587,N_3378,N_4231);
and U8588 (N_8588,N_3393,N_3060);
nor U8589 (N_8589,N_4943,N_109);
or U8590 (N_8590,N_2770,N_4319);
nor U8591 (N_8591,N_2089,N_3996);
nor U8592 (N_8592,N_2338,N_1193);
or U8593 (N_8593,N_236,N_1755);
or U8594 (N_8594,N_1950,N_1558);
nand U8595 (N_8595,N_4878,N_3172);
and U8596 (N_8596,N_2654,N_3522);
or U8597 (N_8597,N_2563,N_4312);
and U8598 (N_8598,N_670,N_304);
and U8599 (N_8599,N_2074,N_571);
or U8600 (N_8600,N_4058,N_2531);
nor U8601 (N_8601,N_3878,N_4027);
nand U8602 (N_8602,N_2192,N_2113);
xor U8603 (N_8603,N_842,N_10);
or U8604 (N_8604,N_4930,N_1541);
xor U8605 (N_8605,N_4813,N_4222);
nor U8606 (N_8606,N_881,N_3483);
nand U8607 (N_8607,N_2464,N_4271);
nand U8608 (N_8608,N_1240,N_3470);
nand U8609 (N_8609,N_2425,N_3653);
nand U8610 (N_8610,N_2878,N_752);
nand U8611 (N_8611,N_1448,N_4718);
nor U8612 (N_8612,N_4238,N_1637);
or U8613 (N_8613,N_209,N_1587);
nor U8614 (N_8614,N_2880,N_3163);
nand U8615 (N_8615,N_4973,N_810);
or U8616 (N_8616,N_895,N_3112);
and U8617 (N_8617,N_2055,N_2067);
and U8618 (N_8618,N_4925,N_4455);
nor U8619 (N_8619,N_2474,N_486);
or U8620 (N_8620,N_1233,N_768);
and U8621 (N_8621,N_3029,N_424);
nand U8622 (N_8622,N_2566,N_1408);
nand U8623 (N_8623,N_3296,N_807);
nand U8624 (N_8624,N_3028,N_2701);
nor U8625 (N_8625,N_4581,N_4391);
or U8626 (N_8626,N_2031,N_3242);
or U8627 (N_8627,N_3892,N_694);
nor U8628 (N_8628,N_1038,N_2973);
and U8629 (N_8629,N_2877,N_4197);
nor U8630 (N_8630,N_305,N_3951);
nor U8631 (N_8631,N_4520,N_3188);
nor U8632 (N_8632,N_3991,N_1395);
nand U8633 (N_8633,N_2046,N_3090);
nor U8634 (N_8634,N_596,N_3299);
and U8635 (N_8635,N_4772,N_4197);
nor U8636 (N_8636,N_2037,N_2158);
nor U8637 (N_8637,N_2525,N_2773);
and U8638 (N_8638,N_2464,N_3794);
nor U8639 (N_8639,N_1574,N_58);
and U8640 (N_8640,N_81,N_3189);
nor U8641 (N_8641,N_4580,N_4666);
nor U8642 (N_8642,N_761,N_3964);
nor U8643 (N_8643,N_575,N_2546);
and U8644 (N_8644,N_4831,N_563);
or U8645 (N_8645,N_102,N_3764);
or U8646 (N_8646,N_768,N_234);
nand U8647 (N_8647,N_496,N_918);
nand U8648 (N_8648,N_4800,N_473);
or U8649 (N_8649,N_4977,N_1574);
and U8650 (N_8650,N_358,N_4607);
xor U8651 (N_8651,N_2427,N_627);
and U8652 (N_8652,N_4568,N_4663);
nand U8653 (N_8653,N_1939,N_506);
and U8654 (N_8654,N_3288,N_4121);
or U8655 (N_8655,N_774,N_3322);
and U8656 (N_8656,N_4367,N_1844);
or U8657 (N_8657,N_2562,N_4641);
xnor U8658 (N_8658,N_1497,N_4489);
and U8659 (N_8659,N_371,N_2925);
xnor U8660 (N_8660,N_1997,N_2549);
or U8661 (N_8661,N_4331,N_171);
or U8662 (N_8662,N_4149,N_1271);
nand U8663 (N_8663,N_295,N_976);
nand U8664 (N_8664,N_1978,N_1467);
or U8665 (N_8665,N_4384,N_3969);
or U8666 (N_8666,N_4670,N_2666);
nor U8667 (N_8667,N_3758,N_611);
or U8668 (N_8668,N_4395,N_4915);
or U8669 (N_8669,N_1323,N_4623);
nand U8670 (N_8670,N_2112,N_2488);
nor U8671 (N_8671,N_999,N_358);
nand U8672 (N_8672,N_3542,N_4307);
or U8673 (N_8673,N_1756,N_1422);
and U8674 (N_8674,N_3130,N_2619);
xnor U8675 (N_8675,N_1636,N_4453);
and U8676 (N_8676,N_2488,N_2499);
xor U8677 (N_8677,N_2249,N_483);
or U8678 (N_8678,N_452,N_1620);
and U8679 (N_8679,N_3201,N_318);
or U8680 (N_8680,N_3800,N_3765);
and U8681 (N_8681,N_3161,N_3951);
nor U8682 (N_8682,N_1104,N_4714);
nand U8683 (N_8683,N_2766,N_2661);
nand U8684 (N_8684,N_2232,N_4929);
nand U8685 (N_8685,N_3911,N_3918);
nand U8686 (N_8686,N_1350,N_3225);
and U8687 (N_8687,N_1467,N_3400);
or U8688 (N_8688,N_963,N_703);
nand U8689 (N_8689,N_2725,N_2695);
nand U8690 (N_8690,N_1124,N_595);
and U8691 (N_8691,N_968,N_2942);
xor U8692 (N_8692,N_13,N_4890);
and U8693 (N_8693,N_4239,N_1614);
nand U8694 (N_8694,N_4373,N_864);
or U8695 (N_8695,N_2744,N_2159);
xnor U8696 (N_8696,N_1959,N_1452);
or U8697 (N_8697,N_1849,N_3986);
or U8698 (N_8698,N_3652,N_3280);
nand U8699 (N_8699,N_2634,N_3639);
or U8700 (N_8700,N_387,N_3133);
or U8701 (N_8701,N_3462,N_296);
or U8702 (N_8702,N_244,N_1963);
or U8703 (N_8703,N_739,N_2942);
nand U8704 (N_8704,N_3840,N_3440);
nor U8705 (N_8705,N_3683,N_633);
or U8706 (N_8706,N_4820,N_4494);
or U8707 (N_8707,N_3388,N_4889);
or U8708 (N_8708,N_576,N_3417);
nand U8709 (N_8709,N_4980,N_3643);
nor U8710 (N_8710,N_2791,N_3991);
or U8711 (N_8711,N_3418,N_1508);
nor U8712 (N_8712,N_3625,N_2924);
and U8713 (N_8713,N_175,N_2227);
nor U8714 (N_8714,N_1342,N_2122);
nor U8715 (N_8715,N_329,N_2933);
nor U8716 (N_8716,N_1906,N_1549);
and U8717 (N_8717,N_641,N_1442);
nor U8718 (N_8718,N_4179,N_3133);
nand U8719 (N_8719,N_527,N_2981);
nor U8720 (N_8720,N_2027,N_1500);
nand U8721 (N_8721,N_2864,N_603);
nand U8722 (N_8722,N_282,N_634);
nor U8723 (N_8723,N_4489,N_1521);
nand U8724 (N_8724,N_4562,N_2176);
nor U8725 (N_8725,N_4710,N_3565);
nor U8726 (N_8726,N_4993,N_3559);
nand U8727 (N_8727,N_2342,N_989);
nor U8728 (N_8728,N_3553,N_3223);
or U8729 (N_8729,N_2080,N_44);
xor U8730 (N_8730,N_3744,N_885);
and U8731 (N_8731,N_582,N_4418);
or U8732 (N_8732,N_2594,N_2465);
and U8733 (N_8733,N_3627,N_3158);
xor U8734 (N_8734,N_3685,N_3888);
nor U8735 (N_8735,N_1882,N_386);
and U8736 (N_8736,N_1268,N_823);
nor U8737 (N_8737,N_3606,N_2615);
and U8738 (N_8738,N_1802,N_914);
and U8739 (N_8739,N_1632,N_2427);
nor U8740 (N_8740,N_1567,N_2188);
nor U8741 (N_8741,N_2889,N_1912);
nor U8742 (N_8742,N_60,N_4903);
xnor U8743 (N_8743,N_3990,N_1389);
nand U8744 (N_8744,N_240,N_3191);
nand U8745 (N_8745,N_3195,N_2983);
nand U8746 (N_8746,N_1675,N_2508);
nand U8747 (N_8747,N_3830,N_4646);
xor U8748 (N_8748,N_2853,N_4918);
and U8749 (N_8749,N_2751,N_3439);
and U8750 (N_8750,N_4423,N_4579);
nor U8751 (N_8751,N_2698,N_3456);
xor U8752 (N_8752,N_1879,N_1027);
and U8753 (N_8753,N_341,N_593);
or U8754 (N_8754,N_4985,N_2694);
or U8755 (N_8755,N_1413,N_1796);
and U8756 (N_8756,N_1732,N_2533);
and U8757 (N_8757,N_4543,N_1691);
and U8758 (N_8758,N_2313,N_1302);
nand U8759 (N_8759,N_2939,N_4975);
and U8760 (N_8760,N_2063,N_4625);
nor U8761 (N_8761,N_4104,N_4746);
nor U8762 (N_8762,N_2207,N_562);
nor U8763 (N_8763,N_3783,N_1282);
xor U8764 (N_8764,N_3279,N_1747);
and U8765 (N_8765,N_863,N_3506);
nor U8766 (N_8766,N_532,N_4988);
nor U8767 (N_8767,N_3825,N_2454);
nand U8768 (N_8768,N_4582,N_3188);
xor U8769 (N_8769,N_3644,N_4363);
nand U8770 (N_8770,N_3132,N_1400);
nand U8771 (N_8771,N_1329,N_2023);
or U8772 (N_8772,N_3163,N_2978);
nand U8773 (N_8773,N_1048,N_4830);
and U8774 (N_8774,N_2538,N_210);
nand U8775 (N_8775,N_67,N_621);
and U8776 (N_8776,N_4323,N_196);
and U8777 (N_8777,N_1767,N_423);
and U8778 (N_8778,N_3771,N_1324);
nand U8779 (N_8779,N_2117,N_3833);
nand U8780 (N_8780,N_988,N_347);
or U8781 (N_8781,N_1382,N_1470);
nor U8782 (N_8782,N_4141,N_3467);
nand U8783 (N_8783,N_1491,N_3669);
and U8784 (N_8784,N_3316,N_4306);
nand U8785 (N_8785,N_1269,N_1372);
nand U8786 (N_8786,N_4176,N_3377);
and U8787 (N_8787,N_4941,N_4120);
xnor U8788 (N_8788,N_2148,N_2824);
or U8789 (N_8789,N_377,N_3894);
nor U8790 (N_8790,N_3588,N_2394);
or U8791 (N_8791,N_94,N_1438);
nor U8792 (N_8792,N_1469,N_598);
or U8793 (N_8793,N_2393,N_605);
and U8794 (N_8794,N_2449,N_2166);
or U8795 (N_8795,N_3636,N_4578);
and U8796 (N_8796,N_2715,N_775);
and U8797 (N_8797,N_190,N_2646);
nand U8798 (N_8798,N_1577,N_49);
nor U8799 (N_8799,N_3990,N_2576);
and U8800 (N_8800,N_2861,N_4234);
nor U8801 (N_8801,N_3283,N_87);
or U8802 (N_8802,N_4661,N_4484);
nor U8803 (N_8803,N_286,N_2779);
xor U8804 (N_8804,N_4918,N_1600);
or U8805 (N_8805,N_2655,N_4781);
or U8806 (N_8806,N_2780,N_4415);
xnor U8807 (N_8807,N_4360,N_3818);
nor U8808 (N_8808,N_2895,N_3703);
or U8809 (N_8809,N_942,N_4497);
xnor U8810 (N_8810,N_4193,N_797);
or U8811 (N_8811,N_4683,N_3602);
xnor U8812 (N_8812,N_1076,N_1935);
nor U8813 (N_8813,N_2314,N_1630);
nor U8814 (N_8814,N_4382,N_3318);
nor U8815 (N_8815,N_342,N_3933);
nand U8816 (N_8816,N_538,N_2210);
nand U8817 (N_8817,N_776,N_3887);
or U8818 (N_8818,N_914,N_3302);
nor U8819 (N_8819,N_4582,N_4771);
nand U8820 (N_8820,N_2936,N_2574);
or U8821 (N_8821,N_3441,N_2186);
nand U8822 (N_8822,N_4388,N_4563);
nand U8823 (N_8823,N_795,N_2218);
xnor U8824 (N_8824,N_4386,N_3606);
xor U8825 (N_8825,N_3614,N_582);
or U8826 (N_8826,N_996,N_4547);
or U8827 (N_8827,N_3482,N_963);
and U8828 (N_8828,N_581,N_3804);
nor U8829 (N_8829,N_2069,N_4478);
or U8830 (N_8830,N_3380,N_950);
or U8831 (N_8831,N_1438,N_3073);
xor U8832 (N_8832,N_836,N_2163);
or U8833 (N_8833,N_3647,N_2193);
and U8834 (N_8834,N_80,N_2953);
nand U8835 (N_8835,N_1583,N_1448);
and U8836 (N_8836,N_1512,N_2617);
and U8837 (N_8837,N_1290,N_4138);
nor U8838 (N_8838,N_1947,N_2974);
nand U8839 (N_8839,N_1927,N_1838);
nor U8840 (N_8840,N_4015,N_344);
or U8841 (N_8841,N_1511,N_889);
xor U8842 (N_8842,N_1349,N_3028);
or U8843 (N_8843,N_3978,N_4587);
nor U8844 (N_8844,N_4831,N_3153);
or U8845 (N_8845,N_3963,N_264);
or U8846 (N_8846,N_2069,N_3208);
and U8847 (N_8847,N_1511,N_2604);
nor U8848 (N_8848,N_4634,N_3112);
xnor U8849 (N_8849,N_4507,N_27);
nand U8850 (N_8850,N_358,N_4510);
nand U8851 (N_8851,N_4854,N_1517);
or U8852 (N_8852,N_691,N_2589);
nor U8853 (N_8853,N_384,N_2859);
nor U8854 (N_8854,N_924,N_1322);
nand U8855 (N_8855,N_1584,N_588);
nor U8856 (N_8856,N_3960,N_2151);
nand U8857 (N_8857,N_509,N_4888);
xor U8858 (N_8858,N_221,N_3303);
nor U8859 (N_8859,N_684,N_1190);
or U8860 (N_8860,N_1770,N_4472);
or U8861 (N_8861,N_2552,N_3799);
and U8862 (N_8862,N_2356,N_4240);
or U8863 (N_8863,N_4028,N_2440);
nand U8864 (N_8864,N_4780,N_1989);
nor U8865 (N_8865,N_4783,N_4065);
and U8866 (N_8866,N_1071,N_253);
nand U8867 (N_8867,N_1593,N_470);
and U8868 (N_8868,N_4981,N_3796);
nand U8869 (N_8869,N_2476,N_55);
nand U8870 (N_8870,N_4960,N_1753);
nand U8871 (N_8871,N_871,N_3596);
and U8872 (N_8872,N_4117,N_523);
and U8873 (N_8873,N_1216,N_4604);
and U8874 (N_8874,N_1448,N_3666);
and U8875 (N_8875,N_1032,N_4282);
nor U8876 (N_8876,N_966,N_3476);
nand U8877 (N_8877,N_606,N_42);
and U8878 (N_8878,N_4537,N_2315);
nor U8879 (N_8879,N_1083,N_2001);
and U8880 (N_8880,N_2480,N_3987);
and U8881 (N_8881,N_2959,N_2408);
or U8882 (N_8882,N_683,N_1176);
xnor U8883 (N_8883,N_4745,N_220);
or U8884 (N_8884,N_1496,N_3897);
or U8885 (N_8885,N_2138,N_1184);
or U8886 (N_8886,N_3254,N_897);
nand U8887 (N_8887,N_2192,N_2563);
nor U8888 (N_8888,N_2591,N_3539);
nor U8889 (N_8889,N_2664,N_58);
nand U8890 (N_8890,N_4659,N_4751);
or U8891 (N_8891,N_4664,N_1931);
nor U8892 (N_8892,N_426,N_1352);
and U8893 (N_8893,N_2136,N_1806);
nand U8894 (N_8894,N_472,N_1148);
or U8895 (N_8895,N_1344,N_4043);
nor U8896 (N_8896,N_3274,N_2131);
and U8897 (N_8897,N_1872,N_251);
xor U8898 (N_8898,N_4733,N_1417);
xnor U8899 (N_8899,N_4771,N_56);
nand U8900 (N_8900,N_248,N_2497);
nor U8901 (N_8901,N_719,N_134);
and U8902 (N_8902,N_64,N_4353);
nor U8903 (N_8903,N_1998,N_2705);
nor U8904 (N_8904,N_1248,N_4779);
and U8905 (N_8905,N_4907,N_4205);
or U8906 (N_8906,N_163,N_3857);
and U8907 (N_8907,N_303,N_2348);
xnor U8908 (N_8908,N_1554,N_1098);
and U8909 (N_8909,N_1320,N_4921);
xnor U8910 (N_8910,N_1581,N_661);
or U8911 (N_8911,N_2735,N_3906);
and U8912 (N_8912,N_3855,N_108);
or U8913 (N_8913,N_2426,N_1894);
nand U8914 (N_8914,N_1372,N_4490);
xor U8915 (N_8915,N_4670,N_420);
or U8916 (N_8916,N_3046,N_4202);
nand U8917 (N_8917,N_4124,N_1042);
nor U8918 (N_8918,N_3356,N_2490);
or U8919 (N_8919,N_3258,N_2717);
nor U8920 (N_8920,N_1153,N_4131);
and U8921 (N_8921,N_3366,N_564);
nor U8922 (N_8922,N_1703,N_2059);
nor U8923 (N_8923,N_1787,N_1952);
and U8924 (N_8924,N_2240,N_79);
nor U8925 (N_8925,N_1118,N_84);
or U8926 (N_8926,N_2377,N_3641);
xnor U8927 (N_8927,N_2467,N_3230);
nor U8928 (N_8928,N_1111,N_2823);
and U8929 (N_8929,N_1006,N_4701);
or U8930 (N_8930,N_43,N_1141);
nand U8931 (N_8931,N_272,N_3083);
or U8932 (N_8932,N_1809,N_3478);
nor U8933 (N_8933,N_4537,N_4798);
and U8934 (N_8934,N_833,N_3422);
nor U8935 (N_8935,N_507,N_3770);
nor U8936 (N_8936,N_1416,N_4144);
nand U8937 (N_8937,N_3398,N_2038);
or U8938 (N_8938,N_3087,N_3602);
nor U8939 (N_8939,N_3402,N_1628);
xor U8940 (N_8940,N_4138,N_3460);
nand U8941 (N_8941,N_812,N_195);
xor U8942 (N_8942,N_1075,N_3999);
xnor U8943 (N_8943,N_2146,N_676);
or U8944 (N_8944,N_592,N_4918);
and U8945 (N_8945,N_23,N_2787);
and U8946 (N_8946,N_1712,N_4086);
nand U8947 (N_8947,N_2083,N_1776);
nor U8948 (N_8948,N_3582,N_2764);
and U8949 (N_8949,N_4503,N_934);
or U8950 (N_8950,N_1887,N_3896);
and U8951 (N_8951,N_3009,N_2072);
nand U8952 (N_8952,N_2297,N_3800);
nand U8953 (N_8953,N_617,N_1096);
nor U8954 (N_8954,N_4659,N_375);
or U8955 (N_8955,N_3273,N_3455);
or U8956 (N_8956,N_3118,N_1040);
nor U8957 (N_8957,N_1016,N_2720);
or U8958 (N_8958,N_130,N_27);
nor U8959 (N_8959,N_3596,N_1024);
nor U8960 (N_8960,N_4519,N_2123);
nor U8961 (N_8961,N_1736,N_2427);
nand U8962 (N_8962,N_1052,N_1683);
xor U8963 (N_8963,N_3185,N_2566);
nor U8964 (N_8964,N_2506,N_3192);
or U8965 (N_8965,N_4671,N_3736);
nor U8966 (N_8966,N_2216,N_1927);
nand U8967 (N_8967,N_2177,N_1714);
nor U8968 (N_8968,N_3842,N_3651);
or U8969 (N_8969,N_1269,N_126);
and U8970 (N_8970,N_43,N_4869);
nor U8971 (N_8971,N_579,N_2285);
or U8972 (N_8972,N_2237,N_3963);
nand U8973 (N_8973,N_688,N_3418);
nand U8974 (N_8974,N_2906,N_1113);
nor U8975 (N_8975,N_3496,N_3661);
or U8976 (N_8976,N_2240,N_90);
or U8977 (N_8977,N_1919,N_3261);
or U8978 (N_8978,N_4854,N_3211);
or U8979 (N_8979,N_2799,N_1794);
or U8980 (N_8980,N_2086,N_634);
and U8981 (N_8981,N_4570,N_2088);
and U8982 (N_8982,N_2592,N_4720);
xor U8983 (N_8983,N_1795,N_3759);
xnor U8984 (N_8984,N_4149,N_2564);
and U8985 (N_8985,N_375,N_4512);
nor U8986 (N_8986,N_4285,N_97);
nand U8987 (N_8987,N_3925,N_2160);
nor U8988 (N_8988,N_766,N_4306);
or U8989 (N_8989,N_2189,N_603);
nand U8990 (N_8990,N_2096,N_3423);
nand U8991 (N_8991,N_4074,N_3015);
or U8992 (N_8992,N_2186,N_994);
nor U8993 (N_8993,N_2620,N_1299);
nand U8994 (N_8994,N_1575,N_2593);
xor U8995 (N_8995,N_2250,N_4715);
and U8996 (N_8996,N_3490,N_1361);
or U8997 (N_8997,N_4035,N_3531);
xor U8998 (N_8998,N_4466,N_3685);
or U8999 (N_8999,N_2099,N_2936);
nand U9000 (N_9000,N_3564,N_3341);
or U9001 (N_9001,N_4685,N_2130);
xnor U9002 (N_9002,N_1755,N_3287);
or U9003 (N_9003,N_3272,N_3756);
or U9004 (N_9004,N_2551,N_1587);
and U9005 (N_9005,N_2394,N_928);
nor U9006 (N_9006,N_923,N_3610);
or U9007 (N_9007,N_2640,N_2669);
nand U9008 (N_9008,N_2477,N_4661);
and U9009 (N_9009,N_2199,N_787);
nand U9010 (N_9010,N_3715,N_658);
nand U9011 (N_9011,N_2458,N_1678);
xnor U9012 (N_9012,N_363,N_2240);
nand U9013 (N_9013,N_3560,N_3732);
xor U9014 (N_9014,N_646,N_2947);
nor U9015 (N_9015,N_3013,N_3077);
nand U9016 (N_9016,N_27,N_2664);
and U9017 (N_9017,N_2317,N_142);
nor U9018 (N_9018,N_231,N_1946);
xor U9019 (N_9019,N_3632,N_4807);
or U9020 (N_9020,N_3039,N_3875);
or U9021 (N_9021,N_4390,N_4821);
nand U9022 (N_9022,N_111,N_4140);
nand U9023 (N_9023,N_100,N_4734);
xor U9024 (N_9024,N_515,N_4265);
nor U9025 (N_9025,N_2028,N_2984);
nor U9026 (N_9026,N_1208,N_459);
nand U9027 (N_9027,N_4063,N_1487);
nor U9028 (N_9028,N_3904,N_2261);
and U9029 (N_9029,N_949,N_2071);
and U9030 (N_9030,N_4238,N_1401);
and U9031 (N_9031,N_3550,N_1730);
and U9032 (N_9032,N_671,N_1344);
nand U9033 (N_9033,N_2840,N_527);
nand U9034 (N_9034,N_1989,N_4666);
nand U9035 (N_9035,N_4888,N_3232);
nor U9036 (N_9036,N_3686,N_2830);
and U9037 (N_9037,N_1402,N_4204);
nor U9038 (N_9038,N_1677,N_3034);
or U9039 (N_9039,N_4778,N_3711);
or U9040 (N_9040,N_2356,N_2476);
xnor U9041 (N_9041,N_3843,N_2972);
or U9042 (N_9042,N_3,N_4561);
and U9043 (N_9043,N_1629,N_2126);
nand U9044 (N_9044,N_3328,N_3895);
or U9045 (N_9045,N_4919,N_2527);
or U9046 (N_9046,N_4563,N_4381);
or U9047 (N_9047,N_1353,N_2123);
and U9048 (N_9048,N_3941,N_1208);
nor U9049 (N_9049,N_4724,N_1007);
nor U9050 (N_9050,N_4143,N_959);
or U9051 (N_9051,N_367,N_4104);
nor U9052 (N_9052,N_317,N_2718);
and U9053 (N_9053,N_2423,N_2007);
or U9054 (N_9054,N_40,N_2263);
nor U9055 (N_9055,N_4071,N_996);
nand U9056 (N_9056,N_1185,N_1515);
or U9057 (N_9057,N_1151,N_430);
nand U9058 (N_9058,N_4542,N_4913);
xnor U9059 (N_9059,N_4418,N_519);
or U9060 (N_9060,N_2723,N_1001);
and U9061 (N_9061,N_1318,N_3272);
or U9062 (N_9062,N_4016,N_3159);
nor U9063 (N_9063,N_2592,N_3858);
and U9064 (N_9064,N_2422,N_2682);
nand U9065 (N_9065,N_608,N_1305);
nor U9066 (N_9066,N_174,N_3764);
nor U9067 (N_9067,N_2950,N_2827);
and U9068 (N_9068,N_3123,N_2571);
and U9069 (N_9069,N_3305,N_2325);
nand U9070 (N_9070,N_1864,N_920);
xnor U9071 (N_9071,N_3400,N_2753);
nor U9072 (N_9072,N_1492,N_1655);
xnor U9073 (N_9073,N_2985,N_2764);
nor U9074 (N_9074,N_376,N_667);
xor U9075 (N_9075,N_2771,N_3070);
nor U9076 (N_9076,N_4908,N_103);
xnor U9077 (N_9077,N_956,N_591);
xor U9078 (N_9078,N_4180,N_1358);
xnor U9079 (N_9079,N_4429,N_3075);
or U9080 (N_9080,N_784,N_3358);
xor U9081 (N_9081,N_4982,N_795);
nand U9082 (N_9082,N_4260,N_493);
nand U9083 (N_9083,N_376,N_4173);
xnor U9084 (N_9084,N_255,N_4601);
or U9085 (N_9085,N_1594,N_2127);
nand U9086 (N_9086,N_2954,N_1791);
nor U9087 (N_9087,N_3537,N_3371);
nor U9088 (N_9088,N_2800,N_569);
and U9089 (N_9089,N_2760,N_185);
or U9090 (N_9090,N_3511,N_1984);
and U9091 (N_9091,N_1320,N_2937);
nand U9092 (N_9092,N_1064,N_4677);
and U9093 (N_9093,N_1072,N_303);
and U9094 (N_9094,N_597,N_2089);
and U9095 (N_9095,N_1578,N_2063);
or U9096 (N_9096,N_188,N_51);
and U9097 (N_9097,N_3118,N_3442);
or U9098 (N_9098,N_116,N_2962);
or U9099 (N_9099,N_1401,N_706);
and U9100 (N_9100,N_3275,N_3586);
or U9101 (N_9101,N_945,N_964);
nand U9102 (N_9102,N_870,N_3514);
nand U9103 (N_9103,N_1685,N_2498);
nand U9104 (N_9104,N_1715,N_723);
nor U9105 (N_9105,N_4732,N_3011);
or U9106 (N_9106,N_1261,N_4744);
or U9107 (N_9107,N_1135,N_4718);
or U9108 (N_9108,N_2279,N_904);
nand U9109 (N_9109,N_3257,N_1120);
nand U9110 (N_9110,N_2986,N_1441);
nand U9111 (N_9111,N_4456,N_2479);
or U9112 (N_9112,N_3625,N_82);
xor U9113 (N_9113,N_1553,N_44);
nand U9114 (N_9114,N_3687,N_3231);
and U9115 (N_9115,N_1542,N_4710);
nor U9116 (N_9116,N_3723,N_3242);
or U9117 (N_9117,N_4042,N_4706);
xnor U9118 (N_9118,N_2580,N_4446);
nand U9119 (N_9119,N_3773,N_2846);
xnor U9120 (N_9120,N_2749,N_1816);
and U9121 (N_9121,N_4264,N_3719);
nor U9122 (N_9122,N_3712,N_1791);
nand U9123 (N_9123,N_141,N_1681);
nand U9124 (N_9124,N_3075,N_1331);
and U9125 (N_9125,N_2090,N_1890);
nand U9126 (N_9126,N_1885,N_895);
and U9127 (N_9127,N_2060,N_4482);
or U9128 (N_9128,N_2376,N_1357);
nand U9129 (N_9129,N_1720,N_4314);
or U9130 (N_9130,N_1334,N_991);
nand U9131 (N_9131,N_2220,N_4240);
and U9132 (N_9132,N_4372,N_4355);
nor U9133 (N_9133,N_1593,N_2989);
nand U9134 (N_9134,N_629,N_237);
nand U9135 (N_9135,N_928,N_1067);
nand U9136 (N_9136,N_3149,N_4503);
and U9137 (N_9137,N_4618,N_4684);
nor U9138 (N_9138,N_4692,N_2010);
or U9139 (N_9139,N_2691,N_4855);
xor U9140 (N_9140,N_2920,N_2636);
nor U9141 (N_9141,N_3471,N_198);
nand U9142 (N_9142,N_1844,N_2145);
nand U9143 (N_9143,N_1729,N_490);
nand U9144 (N_9144,N_3846,N_4607);
or U9145 (N_9145,N_1768,N_701);
or U9146 (N_9146,N_3047,N_665);
nor U9147 (N_9147,N_1175,N_2481);
and U9148 (N_9148,N_1998,N_351);
and U9149 (N_9149,N_563,N_4723);
or U9150 (N_9150,N_1971,N_650);
xnor U9151 (N_9151,N_2268,N_4938);
nor U9152 (N_9152,N_4690,N_2682);
nor U9153 (N_9153,N_3048,N_4053);
or U9154 (N_9154,N_4533,N_2217);
nor U9155 (N_9155,N_321,N_4186);
nor U9156 (N_9156,N_2974,N_1971);
or U9157 (N_9157,N_2793,N_2339);
or U9158 (N_9158,N_841,N_4120);
or U9159 (N_9159,N_437,N_1956);
nand U9160 (N_9160,N_2652,N_4495);
and U9161 (N_9161,N_3784,N_2341);
nand U9162 (N_9162,N_1488,N_2143);
nor U9163 (N_9163,N_4108,N_3283);
or U9164 (N_9164,N_2857,N_4228);
nand U9165 (N_9165,N_2010,N_2035);
nand U9166 (N_9166,N_1464,N_4037);
and U9167 (N_9167,N_1904,N_4654);
and U9168 (N_9168,N_2264,N_1571);
or U9169 (N_9169,N_4750,N_4414);
and U9170 (N_9170,N_840,N_1339);
and U9171 (N_9171,N_1528,N_2935);
and U9172 (N_9172,N_3985,N_1373);
and U9173 (N_9173,N_4645,N_491);
xnor U9174 (N_9174,N_1626,N_4965);
xor U9175 (N_9175,N_2733,N_4978);
nand U9176 (N_9176,N_32,N_2391);
and U9177 (N_9177,N_1004,N_4119);
or U9178 (N_9178,N_1544,N_3498);
and U9179 (N_9179,N_3861,N_3719);
and U9180 (N_9180,N_2229,N_4134);
nand U9181 (N_9181,N_2433,N_3250);
or U9182 (N_9182,N_4695,N_4069);
nor U9183 (N_9183,N_1998,N_2345);
nand U9184 (N_9184,N_27,N_842);
and U9185 (N_9185,N_3011,N_2168);
nand U9186 (N_9186,N_1548,N_4340);
nand U9187 (N_9187,N_4305,N_6);
nor U9188 (N_9188,N_1060,N_1782);
nor U9189 (N_9189,N_3578,N_824);
and U9190 (N_9190,N_4723,N_790);
nor U9191 (N_9191,N_2022,N_1546);
and U9192 (N_9192,N_1665,N_1670);
nor U9193 (N_9193,N_4959,N_1697);
nor U9194 (N_9194,N_1831,N_1957);
xnor U9195 (N_9195,N_3929,N_557);
or U9196 (N_9196,N_847,N_17);
or U9197 (N_9197,N_2938,N_1251);
nand U9198 (N_9198,N_1373,N_1748);
nor U9199 (N_9199,N_128,N_4813);
or U9200 (N_9200,N_4218,N_3699);
or U9201 (N_9201,N_4553,N_2150);
nor U9202 (N_9202,N_4715,N_2614);
or U9203 (N_9203,N_4761,N_2830);
or U9204 (N_9204,N_4966,N_29);
xnor U9205 (N_9205,N_4345,N_1362);
or U9206 (N_9206,N_4847,N_2479);
or U9207 (N_9207,N_2998,N_1893);
and U9208 (N_9208,N_4338,N_3296);
nand U9209 (N_9209,N_3570,N_4393);
or U9210 (N_9210,N_4805,N_2176);
and U9211 (N_9211,N_1162,N_1824);
nand U9212 (N_9212,N_80,N_4137);
nor U9213 (N_9213,N_275,N_4844);
or U9214 (N_9214,N_4942,N_535);
nor U9215 (N_9215,N_62,N_1503);
nand U9216 (N_9216,N_2561,N_761);
nor U9217 (N_9217,N_1124,N_3696);
or U9218 (N_9218,N_4758,N_1425);
and U9219 (N_9219,N_3517,N_4880);
or U9220 (N_9220,N_818,N_4238);
nand U9221 (N_9221,N_3871,N_4843);
nor U9222 (N_9222,N_1210,N_2780);
or U9223 (N_9223,N_3669,N_3677);
and U9224 (N_9224,N_3946,N_523);
nand U9225 (N_9225,N_316,N_2547);
nor U9226 (N_9226,N_4736,N_285);
nand U9227 (N_9227,N_4171,N_4270);
nor U9228 (N_9228,N_1512,N_319);
or U9229 (N_9229,N_4300,N_2035);
or U9230 (N_9230,N_2299,N_1872);
nand U9231 (N_9231,N_3111,N_3440);
nand U9232 (N_9232,N_1585,N_4825);
nor U9233 (N_9233,N_1538,N_4474);
and U9234 (N_9234,N_2129,N_1328);
xnor U9235 (N_9235,N_1564,N_1724);
nand U9236 (N_9236,N_3739,N_2693);
and U9237 (N_9237,N_2016,N_941);
nor U9238 (N_9238,N_1364,N_1660);
xnor U9239 (N_9239,N_3288,N_1528);
and U9240 (N_9240,N_2264,N_3415);
or U9241 (N_9241,N_1594,N_3375);
nor U9242 (N_9242,N_3842,N_1109);
and U9243 (N_9243,N_1220,N_4797);
nand U9244 (N_9244,N_787,N_3031);
xor U9245 (N_9245,N_338,N_4661);
nand U9246 (N_9246,N_4141,N_2861);
nor U9247 (N_9247,N_3671,N_1312);
nand U9248 (N_9248,N_2170,N_3800);
or U9249 (N_9249,N_3854,N_1661);
nor U9250 (N_9250,N_2401,N_1936);
nand U9251 (N_9251,N_327,N_753);
xor U9252 (N_9252,N_3162,N_998);
xnor U9253 (N_9253,N_3486,N_3468);
nand U9254 (N_9254,N_2717,N_33);
nand U9255 (N_9255,N_2639,N_655);
xnor U9256 (N_9256,N_697,N_2553);
or U9257 (N_9257,N_4271,N_2841);
nand U9258 (N_9258,N_4772,N_418);
nor U9259 (N_9259,N_609,N_2408);
nor U9260 (N_9260,N_1760,N_301);
nand U9261 (N_9261,N_868,N_3708);
or U9262 (N_9262,N_1364,N_2711);
or U9263 (N_9263,N_134,N_136);
xnor U9264 (N_9264,N_3347,N_4881);
or U9265 (N_9265,N_2789,N_1792);
and U9266 (N_9266,N_3727,N_1698);
or U9267 (N_9267,N_2037,N_1231);
nor U9268 (N_9268,N_1283,N_3317);
and U9269 (N_9269,N_2318,N_1066);
and U9270 (N_9270,N_3853,N_1610);
or U9271 (N_9271,N_1015,N_4761);
nor U9272 (N_9272,N_2716,N_4112);
nand U9273 (N_9273,N_1722,N_2590);
or U9274 (N_9274,N_1560,N_366);
nor U9275 (N_9275,N_353,N_902);
nand U9276 (N_9276,N_4885,N_642);
or U9277 (N_9277,N_2729,N_1346);
nor U9278 (N_9278,N_2721,N_4334);
nor U9279 (N_9279,N_4441,N_3550);
and U9280 (N_9280,N_3062,N_1892);
or U9281 (N_9281,N_1855,N_2892);
nand U9282 (N_9282,N_8,N_970);
xnor U9283 (N_9283,N_3628,N_2171);
nor U9284 (N_9284,N_3933,N_993);
nor U9285 (N_9285,N_2037,N_4358);
nor U9286 (N_9286,N_829,N_3040);
nor U9287 (N_9287,N_330,N_4366);
nor U9288 (N_9288,N_41,N_522);
nand U9289 (N_9289,N_257,N_3542);
or U9290 (N_9290,N_578,N_856);
xor U9291 (N_9291,N_4228,N_1264);
or U9292 (N_9292,N_2131,N_1725);
or U9293 (N_9293,N_3081,N_3661);
nor U9294 (N_9294,N_2658,N_1372);
nor U9295 (N_9295,N_1604,N_592);
nand U9296 (N_9296,N_1773,N_3076);
nand U9297 (N_9297,N_2817,N_3104);
nand U9298 (N_9298,N_896,N_1863);
nor U9299 (N_9299,N_4431,N_4884);
and U9300 (N_9300,N_3963,N_3511);
nor U9301 (N_9301,N_800,N_2696);
nor U9302 (N_9302,N_2179,N_3037);
nand U9303 (N_9303,N_1461,N_3622);
nand U9304 (N_9304,N_4728,N_2302);
nand U9305 (N_9305,N_515,N_3863);
or U9306 (N_9306,N_1570,N_842);
or U9307 (N_9307,N_4777,N_622);
nand U9308 (N_9308,N_2413,N_3309);
nor U9309 (N_9309,N_4514,N_1272);
nand U9310 (N_9310,N_1729,N_3873);
or U9311 (N_9311,N_982,N_1050);
nand U9312 (N_9312,N_3824,N_1604);
or U9313 (N_9313,N_4486,N_830);
nor U9314 (N_9314,N_3777,N_2665);
xnor U9315 (N_9315,N_4077,N_678);
nor U9316 (N_9316,N_2051,N_298);
or U9317 (N_9317,N_1870,N_3969);
or U9318 (N_9318,N_1959,N_3563);
or U9319 (N_9319,N_4079,N_2500);
and U9320 (N_9320,N_3564,N_1670);
nor U9321 (N_9321,N_4897,N_3106);
nand U9322 (N_9322,N_524,N_4065);
and U9323 (N_9323,N_3218,N_4629);
nor U9324 (N_9324,N_3540,N_391);
and U9325 (N_9325,N_3499,N_3472);
and U9326 (N_9326,N_2904,N_849);
and U9327 (N_9327,N_4388,N_2951);
nor U9328 (N_9328,N_4076,N_3207);
and U9329 (N_9329,N_3474,N_1100);
nor U9330 (N_9330,N_2191,N_2493);
or U9331 (N_9331,N_4510,N_1891);
nand U9332 (N_9332,N_3874,N_359);
nand U9333 (N_9333,N_3501,N_2388);
xnor U9334 (N_9334,N_1727,N_1698);
nor U9335 (N_9335,N_488,N_1631);
and U9336 (N_9336,N_3183,N_51);
nand U9337 (N_9337,N_486,N_4254);
or U9338 (N_9338,N_3430,N_4971);
and U9339 (N_9339,N_333,N_4902);
or U9340 (N_9340,N_2306,N_629);
xnor U9341 (N_9341,N_4483,N_1418);
nand U9342 (N_9342,N_2226,N_937);
xor U9343 (N_9343,N_3734,N_3894);
nor U9344 (N_9344,N_4942,N_74);
nand U9345 (N_9345,N_555,N_3563);
nor U9346 (N_9346,N_2653,N_177);
or U9347 (N_9347,N_4950,N_120);
or U9348 (N_9348,N_384,N_498);
or U9349 (N_9349,N_218,N_1545);
and U9350 (N_9350,N_1141,N_2554);
nor U9351 (N_9351,N_2551,N_2524);
nand U9352 (N_9352,N_3044,N_2986);
and U9353 (N_9353,N_4276,N_3329);
nand U9354 (N_9354,N_713,N_4667);
nor U9355 (N_9355,N_2368,N_1621);
and U9356 (N_9356,N_1980,N_231);
nor U9357 (N_9357,N_2431,N_1723);
nand U9358 (N_9358,N_707,N_2998);
nand U9359 (N_9359,N_4101,N_4943);
and U9360 (N_9360,N_2733,N_2528);
or U9361 (N_9361,N_4533,N_3791);
and U9362 (N_9362,N_2134,N_4561);
nand U9363 (N_9363,N_259,N_848);
xnor U9364 (N_9364,N_2582,N_2948);
or U9365 (N_9365,N_322,N_4185);
xor U9366 (N_9366,N_2267,N_762);
or U9367 (N_9367,N_4538,N_29);
xnor U9368 (N_9368,N_1642,N_2612);
xnor U9369 (N_9369,N_4636,N_2359);
nand U9370 (N_9370,N_4495,N_4125);
or U9371 (N_9371,N_3158,N_210);
nand U9372 (N_9372,N_2429,N_937);
or U9373 (N_9373,N_3469,N_877);
xor U9374 (N_9374,N_3355,N_587);
nand U9375 (N_9375,N_4475,N_3329);
nand U9376 (N_9376,N_44,N_4797);
nand U9377 (N_9377,N_1790,N_833);
and U9378 (N_9378,N_497,N_4195);
nand U9379 (N_9379,N_3829,N_435);
xnor U9380 (N_9380,N_97,N_4926);
and U9381 (N_9381,N_3233,N_2220);
nor U9382 (N_9382,N_3515,N_2054);
nand U9383 (N_9383,N_2860,N_3199);
nor U9384 (N_9384,N_3167,N_3190);
nand U9385 (N_9385,N_26,N_798);
nand U9386 (N_9386,N_2010,N_2144);
or U9387 (N_9387,N_1817,N_1281);
nor U9388 (N_9388,N_1132,N_541);
or U9389 (N_9389,N_4345,N_76);
xnor U9390 (N_9390,N_3664,N_3096);
xor U9391 (N_9391,N_1541,N_3011);
nand U9392 (N_9392,N_2600,N_1857);
or U9393 (N_9393,N_4641,N_1991);
or U9394 (N_9394,N_2103,N_3017);
xnor U9395 (N_9395,N_2988,N_1577);
nand U9396 (N_9396,N_2389,N_2540);
and U9397 (N_9397,N_4948,N_3645);
or U9398 (N_9398,N_3504,N_3639);
or U9399 (N_9399,N_4647,N_2721);
or U9400 (N_9400,N_2958,N_649);
nor U9401 (N_9401,N_1651,N_3125);
or U9402 (N_9402,N_3356,N_2665);
nor U9403 (N_9403,N_4307,N_2862);
nor U9404 (N_9404,N_1322,N_3402);
and U9405 (N_9405,N_1297,N_2086);
and U9406 (N_9406,N_800,N_894);
or U9407 (N_9407,N_4636,N_2326);
xor U9408 (N_9408,N_428,N_1367);
nor U9409 (N_9409,N_1010,N_503);
nand U9410 (N_9410,N_3643,N_2410);
and U9411 (N_9411,N_3643,N_3314);
nor U9412 (N_9412,N_1402,N_4365);
nor U9413 (N_9413,N_3261,N_3402);
xor U9414 (N_9414,N_2890,N_1141);
or U9415 (N_9415,N_664,N_56);
nand U9416 (N_9416,N_3894,N_2082);
nand U9417 (N_9417,N_3530,N_4096);
or U9418 (N_9418,N_1499,N_2530);
xnor U9419 (N_9419,N_1140,N_588);
nand U9420 (N_9420,N_963,N_2689);
and U9421 (N_9421,N_2370,N_153);
nand U9422 (N_9422,N_2438,N_1979);
and U9423 (N_9423,N_3647,N_1501);
xor U9424 (N_9424,N_4577,N_2993);
or U9425 (N_9425,N_3358,N_778);
and U9426 (N_9426,N_865,N_2978);
nand U9427 (N_9427,N_3843,N_3275);
nor U9428 (N_9428,N_2177,N_3191);
nor U9429 (N_9429,N_2529,N_3936);
nor U9430 (N_9430,N_1582,N_1458);
nor U9431 (N_9431,N_1661,N_1512);
and U9432 (N_9432,N_788,N_32);
or U9433 (N_9433,N_43,N_4809);
xnor U9434 (N_9434,N_3043,N_255);
nand U9435 (N_9435,N_1015,N_2576);
nor U9436 (N_9436,N_2040,N_57);
nor U9437 (N_9437,N_380,N_1380);
nand U9438 (N_9438,N_3906,N_4413);
and U9439 (N_9439,N_4633,N_2229);
nor U9440 (N_9440,N_2099,N_4849);
nor U9441 (N_9441,N_2885,N_1347);
nand U9442 (N_9442,N_4998,N_30);
nand U9443 (N_9443,N_1835,N_1453);
nand U9444 (N_9444,N_3338,N_2069);
nand U9445 (N_9445,N_4248,N_4698);
or U9446 (N_9446,N_1995,N_2572);
nand U9447 (N_9447,N_192,N_3143);
xnor U9448 (N_9448,N_4891,N_4752);
nor U9449 (N_9449,N_1930,N_1942);
and U9450 (N_9450,N_2533,N_4472);
and U9451 (N_9451,N_1647,N_2754);
xnor U9452 (N_9452,N_2850,N_2504);
nor U9453 (N_9453,N_2465,N_4859);
and U9454 (N_9454,N_3998,N_4803);
or U9455 (N_9455,N_3470,N_318);
nand U9456 (N_9456,N_2781,N_3255);
nand U9457 (N_9457,N_272,N_2075);
nor U9458 (N_9458,N_1529,N_3888);
nor U9459 (N_9459,N_1306,N_2181);
or U9460 (N_9460,N_2997,N_3494);
and U9461 (N_9461,N_763,N_3305);
and U9462 (N_9462,N_8,N_3048);
and U9463 (N_9463,N_4439,N_3964);
or U9464 (N_9464,N_4985,N_4739);
nor U9465 (N_9465,N_1938,N_3872);
and U9466 (N_9466,N_459,N_3129);
and U9467 (N_9467,N_1645,N_1399);
or U9468 (N_9468,N_123,N_782);
and U9469 (N_9469,N_2657,N_2689);
or U9470 (N_9470,N_1859,N_4165);
nand U9471 (N_9471,N_1735,N_2823);
nand U9472 (N_9472,N_1939,N_2219);
nand U9473 (N_9473,N_3148,N_3602);
and U9474 (N_9474,N_4538,N_829);
nor U9475 (N_9475,N_3516,N_591);
or U9476 (N_9476,N_26,N_747);
nor U9477 (N_9477,N_271,N_2297);
nor U9478 (N_9478,N_734,N_2731);
nand U9479 (N_9479,N_2077,N_4755);
nand U9480 (N_9480,N_2984,N_2926);
nor U9481 (N_9481,N_4978,N_4713);
nor U9482 (N_9482,N_1955,N_2340);
nand U9483 (N_9483,N_873,N_1601);
or U9484 (N_9484,N_1916,N_617);
and U9485 (N_9485,N_3665,N_1896);
or U9486 (N_9486,N_2466,N_3214);
nor U9487 (N_9487,N_1888,N_2673);
nand U9488 (N_9488,N_1645,N_1667);
and U9489 (N_9489,N_1590,N_1021);
nor U9490 (N_9490,N_815,N_3052);
nor U9491 (N_9491,N_3542,N_4457);
nor U9492 (N_9492,N_316,N_335);
and U9493 (N_9493,N_4733,N_3484);
and U9494 (N_9494,N_4368,N_4243);
and U9495 (N_9495,N_2353,N_3565);
xor U9496 (N_9496,N_3374,N_1164);
nor U9497 (N_9497,N_378,N_86);
or U9498 (N_9498,N_2988,N_3918);
nand U9499 (N_9499,N_3062,N_234);
nand U9500 (N_9500,N_4401,N_1362);
nand U9501 (N_9501,N_4027,N_4507);
nor U9502 (N_9502,N_1098,N_2841);
nand U9503 (N_9503,N_2123,N_3870);
nor U9504 (N_9504,N_3906,N_2104);
or U9505 (N_9505,N_1078,N_3085);
and U9506 (N_9506,N_466,N_798);
and U9507 (N_9507,N_1674,N_3995);
nand U9508 (N_9508,N_2813,N_840);
nand U9509 (N_9509,N_3509,N_3033);
nand U9510 (N_9510,N_2127,N_4254);
nand U9511 (N_9511,N_4321,N_2629);
nor U9512 (N_9512,N_4021,N_1545);
nor U9513 (N_9513,N_2752,N_4419);
nor U9514 (N_9514,N_770,N_4618);
or U9515 (N_9515,N_4182,N_1605);
nand U9516 (N_9516,N_1347,N_133);
nor U9517 (N_9517,N_1635,N_3171);
or U9518 (N_9518,N_1904,N_1165);
nor U9519 (N_9519,N_2055,N_2120);
or U9520 (N_9520,N_4134,N_2120);
and U9521 (N_9521,N_3869,N_2767);
and U9522 (N_9522,N_4078,N_965);
nand U9523 (N_9523,N_4753,N_4091);
xnor U9524 (N_9524,N_3854,N_4602);
nor U9525 (N_9525,N_4159,N_1109);
or U9526 (N_9526,N_1736,N_1695);
nand U9527 (N_9527,N_902,N_2159);
nand U9528 (N_9528,N_2007,N_1911);
xnor U9529 (N_9529,N_1800,N_4981);
nor U9530 (N_9530,N_3210,N_1773);
nor U9531 (N_9531,N_187,N_1600);
and U9532 (N_9532,N_2980,N_1201);
nand U9533 (N_9533,N_4101,N_3442);
nand U9534 (N_9534,N_3757,N_578);
nor U9535 (N_9535,N_1743,N_3140);
or U9536 (N_9536,N_1967,N_3025);
nand U9537 (N_9537,N_3023,N_3819);
or U9538 (N_9538,N_968,N_2212);
xor U9539 (N_9539,N_291,N_3968);
nand U9540 (N_9540,N_2938,N_1014);
nor U9541 (N_9541,N_4865,N_1769);
nor U9542 (N_9542,N_2631,N_3953);
xnor U9543 (N_9543,N_536,N_1072);
or U9544 (N_9544,N_3443,N_2350);
xnor U9545 (N_9545,N_1927,N_2493);
and U9546 (N_9546,N_959,N_1317);
nor U9547 (N_9547,N_4303,N_2979);
nor U9548 (N_9548,N_3135,N_12);
nand U9549 (N_9549,N_3291,N_4325);
and U9550 (N_9550,N_1613,N_3127);
nand U9551 (N_9551,N_344,N_2800);
or U9552 (N_9552,N_2436,N_3309);
nand U9553 (N_9553,N_2444,N_4352);
and U9554 (N_9554,N_1287,N_3196);
or U9555 (N_9555,N_2216,N_594);
nor U9556 (N_9556,N_825,N_2334);
nor U9557 (N_9557,N_1939,N_4069);
xor U9558 (N_9558,N_2033,N_2113);
nand U9559 (N_9559,N_4635,N_75);
xnor U9560 (N_9560,N_4568,N_3211);
nor U9561 (N_9561,N_2024,N_2044);
and U9562 (N_9562,N_3346,N_1005);
nor U9563 (N_9563,N_487,N_617);
or U9564 (N_9564,N_4805,N_2264);
and U9565 (N_9565,N_2662,N_104);
nand U9566 (N_9566,N_525,N_472);
and U9567 (N_9567,N_2212,N_4895);
and U9568 (N_9568,N_4306,N_1120);
and U9569 (N_9569,N_2370,N_3329);
xnor U9570 (N_9570,N_1059,N_3226);
and U9571 (N_9571,N_1151,N_4756);
and U9572 (N_9572,N_3531,N_734);
and U9573 (N_9573,N_3820,N_3471);
nor U9574 (N_9574,N_2019,N_4757);
and U9575 (N_9575,N_3079,N_1805);
nand U9576 (N_9576,N_923,N_1748);
nor U9577 (N_9577,N_1646,N_4611);
nor U9578 (N_9578,N_3053,N_780);
and U9579 (N_9579,N_1889,N_2987);
nand U9580 (N_9580,N_1532,N_1438);
nor U9581 (N_9581,N_3994,N_3495);
or U9582 (N_9582,N_2585,N_1919);
nor U9583 (N_9583,N_2387,N_1052);
xnor U9584 (N_9584,N_1524,N_2037);
or U9585 (N_9585,N_2286,N_3120);
and U9586 (N_9586,N_851,N_4806);
nand U9587 (N_9587,N_394,N_3282);
nand U9588 (N_9588,N_3168,N_819);
xor U9589 (N_9589,N_3121,N_1591);
and U9590 (N_9590,N_2179,N_4557);
nor U9591 (N_9591,N_1958,N_4026);
nand U9592 (N_9592,N_2061,N_1213);
nand U9593 (N_9593,N_4864,N_2049);
xor U9594 (N_9594,N_754,N_3892);
xor U9595 (N_9595,N_995,N_1027);
or U9596 (N_9596,N_1314,N_1329);
xor U9597 (N_9597,N_139,N_4349);
nand U9598 (N_9598,N_2371,N_763);
nand U9599 (N_9599,N_3020,N_1932);
or U9600 (N_9600,N_4437,N_2745);
or U9601 (N_9601,N_3191,N_2799);
xnor U9602 (N_9602,N_1367,N_4545);
and U9603 (N_9603,N_2540,N_4432);
nor U9604 (N_9604,N_267,N_1614);
and U9605 (N_9605,N_1072,N_3139);
and U9606 (N_9606,N_4920,N_1952);
or U9607 (N_9607,N_81,N_1063);
nor U9608 (N_9608,N_3004,N_2482);
nor U9609 (N_9609,N_4162,N_3479);
and U9610 (N_9610,N_1169,N_3481);
and U9611 (N_9611,N_2737,N_4321);
nor U9612 (N_9612,N_332,N_1305);
or U9613 (N_9613,N_4627,N_1976);
nor U9614 (N_9614,N_4772,N_2024);
and U9615 (N_9615,N_1908,N_2847);
or U9616 (N_9616,N_4979,N_577);
nand U9617 (N_9617,N_776,N_1596);
nand U9618 (N_9618,N_2606,N_2194);
nor U9619 (N_9619,N_2164,N_3714);
and U9620 (N_9620,N_3698,N_2869);
nand U9621 (N_9621,N_4307,N_4125);
nand U9622 (N_9622,N_879,N_3301);
nand U9623 (N_9623,N_3288,N_1409);
or U9624 (N_9624,N_1996,N_2242);
or U9625 (N_9625,N_1201,N_218);
xnor U9626 (N_9626,N_3893,N_1596);
or U9627 (N_9627,N_4275,N_3733);
nand U9628 (N_9628,N_575,N_4309);
or U9629 (N_9629,N_4386,N_3052);
xor U9630 (N_9630,N_4650,N_1508);
and U9631 (N_9631,N_2324,N_898);
or U9632 (N_9632,N_3173,N_3707);
nand U9633 (N_9633,N_4713,N_3939);
nor U9634 (N_9634,N_728,N_2490);
nor U9635 (N_9635,N_630,N_2668);
or U9636 (N_9636,N_3104,N_614);
nand U9637 (N_9637,N_3363,N_3913);
or U9638 (N_9638,N_1763,N_2357);
and U9639 (N_9639,N_2213,N_3243);
or U9640 (N_9640,N_1827,N_4614);
or U9641 (N_9641,N_4601,N_719);
nor U9642 (N_9642,N_2544,N_2510);
or U9643 (N_9643,N_1601,N_775);
nor U9644 (N_9644,N_4164,N_2560);
nor U9645 (N_9645,N_3321,N_4438);
xor U9646 (N_9646,N_4626,N_1523);
or U9647 (N_9647,N_4615,N_2776);
nand U9648 (N_9648,N_4688,N_4145);
nand U9649 (N_9649,N_2992,N_873);
nand U9650 (N_9650,N_2309,N_2136);
nand U9651 (N_9651,N_3244,N_2970);
or U9652 (N_9652,N_3737,N_4083);
xor U9653 (N_9653,N_823,N_4805);
nand U9654 (N_9654,N_2397,N_2529);
and U9655 (N_9655,N_568,N_2759);
nor U9656 (N_9656,N_1969,N_229);
xor U9657 (N_9657,N_4349,N_1324);
nand U9658 (N_9658,N_4414,N_1138);
nor U9659 (N_9659,N_4120,N_3177);
and U9660 (N_9660,N_1831,N_3402);
nor U9661 (N_9661,N_4639,N_3414);
and U9662 (N_9662,N_802,N_3763);
and U9663 (N_9663,N_332,N_1865);
nand U9664 (N_9664,N_1771,N_2687);
or U9665 (N_9665,N_3000,N_2848);
nand U9666 (N_9666,N_4916,N_1491);
xor U9667 (N_9667,N_517,N_1603);
or U9668 (N_9668,N_3378,N_3371);
and U9669 (N_9669,N_4156,N_3774);
xnor U9670 (N_9670,N_4173,N_1299);
and U9671 (N_9671,N_1818,N_2286);
xnor U9672 (N_9672,N_4862,N_2018);
or U9673 (N_9673,N_414,N_2871);
and U9674 (N_9674,N_4685,N_4802);
and U9675 (N_9675,N_3922,N_2536);
nor U9676 (N_9676,N_2221,N_4252);
xor U9677 (N_9677,N_1242,N_1827);
xnor U9678 (N_9678,N_3717,N_247);
nand U9679 (N_9679,N_2989,N_4434);
nand U9680 (N_9680,N_139,N_2725);
nor U9681 (N_9681,N_1683,N_253);
nand U9682 (N_9682,N_2835,N_363);
and U9683 (N_9683,N_3143,N_4285);
nor U9684 (N_9684,N_88,N_1413);
nor U9685 (N_9685,N_2871,N_638);
nor U9686 (N_9686,N_4583,N_432);
nand U9687 (N_9687,N_821,N_2442);
or U9688 (N_9688,N_4233,N_3796);
and U9689 (N_9689,N_4985,N_2049);
or U9690 (N_9690,N_1303,N_81);
xnor U9691 (N_9691,N_4953,N_691);
nor U9692 (N_9692,N_4063,N_4741);
nor U9693 (N_9693,N_1708,N_4755);
nor U9694 (N_9694,N_3729,N_1623);
and U9695 (N_9695,N_4684,N_634);
nand U9696 (N_9696,N_3936,N_2157);
and U9697 (N_9697,N_3820,N_3856);
or U9698 (N_9698,N_4919,N_3270);
nor U9699 (N_9699,N_4151,N_63);
nor U9700 (N_9700,N_2676,N_1446);
nand U9701 (N_9701,N_1361,N_4860);
nand U9702 (N_9702,N_1249,N_3914);
nor U9703 (N_9703,N_4382,N_898);
nor U9704 (N_9704,N_3388,N_4983);
and U9705 (N_9705,N_3068,N_2195);
xor U9706 (N_9706,N_126,N_1700);
nand U9707 (N_9707,N_4615,N_1543);
nand U9708 (N_9708,N_2977,N_3467);
or U9709 (N_9709,N_2883,N_3049);
nand U9710 (N_9710,N_1363,N_3408);
nor U9711 (N_9711,N_4819,N_3089);
nor U9712 (N_9712,N_848,N_1700);
nand U9713 (N_9713,N_1694,N_578);
nand U9714 (N_9714,N_4495,N_4826);
or U9715 (N_9715,N_1913,N_3831);
and U9716 (N_9716,N_4873,N_4800);
and U9717 (N_9717,N_3815,N_1032);
nand U9718 (N_9718,N_2115,N_1937);
or U9719 (N_9719,N_4850,N_1851);
or U9720 (N_9720,N_1248,N_4275);
or U9721 (N_9721,N_2382,N_3959);
and U9722 (N_9722,N_3320,N_4272);
nor U9723 (N_9723,N_663,N_3284);
nand U9724 (N_9724,N_523,N_4063);
nor U9725 (N_9725,N_4118,N_3899);
or U9726 (N_9726,N_1628,N_3761);
or U9727 (N_9727,N_3051,N_4176);
nand U9728 (N_9728,N_1468,N_466);
nor U9729 (N_9729,N_449,N_4320);
nand U9730 (N_9730,N_3651,N_549);
and U9731 (N_9731,N_4122,N_3332);
nor U9732 (N_9732,N_3829,N_2953);
or U9733 (N_9733,N_1039,N_969);
or U9734 (N_9734,N_4907,N_2520);
or U9735 (N_9735,N_13,N_765);
nand U9736 (N_9736,N_2540,N_2350);
and U9737 (N_9737,N_734,N_4051);
nor U9738 (N_9738,N_4945,N_1891);
nand U9739 (N_9739,N_3387,N_531);
or U9740 (N_9740,N_3067,N_2601);
nand U9741 (N_9741,N_705,N_3686);
xor U9742 (N_9742,N_3617,N_1593);
nand U9743 (N_9743,N_959,N_4779);
or U9744 (N_9744,N_3039,N_2242);
and U9745 (N_9745,N_4463,N_4004);
nor U9746 (N_9746,N_3255,N_2190);
nor U9747 (N_9747,N_3552,N_2037);
and U9748 (N_9748,N_1578,N_3925);
and U9749 (N_9749,N_1154,N_1193);
nor U9750 (N_9750,N_1431,N_593);
nand U9751 (N_9751,N_2748,N_3841);
nand U9752 (N_9752,N_1770,N_2933);
nand U9753 (N_9753,N_2484,N_4278);
and U9754 (N_9754,N_1190,N_2718);
nand U9755 (N_9755,N_2228,N_3768);
nand U9756 (N_9756,N_2528,N_3649);
or U9757 (N_9757,N_2957,N_2706);
or U9758 (N_9758,N_483,N_1490);
and U9759 (N_9759,N_266,N_0);
or U9760 (N_9760,N_4823,N_4504);
or U9761 (N_9761,N_4736,N_2479);
and U9762 (N_9762,N_1247,N_2654);
xor U9763 (N_9763,N_1109,N_3939);
or U9764 (N_9764,N_2133,N_1463);
and U9765 (N_9765,N_2371,N_3564);
or U9766 (N_9766,N_3310,N_2047);
nor U9767 (N_9767,N_2937,N_761);
nor U9768 (N_9768,N_4380,N_2522);
and U9769 (N_9769,N_2851,N_2348);
and U9770 (N_9770,N_4202,N_1751);
and U9771 (N_9771,N_827,N_3041);
nor U9772 (N_9772,N_2665,N_483);
and U9773 (N_9773,N_4245,N_1550);
and U9774 (N_9774,N_3985,N_4773);
xnor U9775 (N_9775,N_4231,N_2671);
and U9776 (N_9776,N_4802,N_4464);
or U9777 (N_9777,N_290,N_246);
nand U9778 (N_9778,N_525,N_4995);
and U9779 (N_9779,N_3025,N_2641);
nand U9780 (N_9780,N_3017,N_137);
nand U9781 (N_9781,N_3933,N_2386);
nand U9782 (N_9782,N_362,N_1501);
or U9783 (N_9783,N_3621,N_1391);
and U9784 (N_9784,N_2857,N_1972);
and U9785 (N_9785,N_4053,N_2354);
nand U9786 (N_9786,N_4909,N_1013);
nand U9787 (N_9787,N_4539,N_4642);
and U9788 (N_9788,N_331,N_282);
or U9789 (N_9789,N_1849,N_2900);
nor U9790 (N_9790,N_2375,N_2466);
xor U9791 (N_9791,N_71,N_3672);
nor U9792 (N_9792,N_439,N_3172);
nand U9793 (N_9793,N_3787,N_1407);
nand U9794 (N_9794,N_1164,N_387);
xnor U9795 (N_9795,N_3645,N_243);
nor U9796 (N_9796,N_222,N_2938);
xor U9797 (N_9797,N_1360,N_2434);
nor U9798 (N_9798,N_2634,N_132);
nor U9799 (N_9799,N_3089,N_4590);
nor U9800 (N_9800,N_4835,N_2875);
nand U9801 (N_9801,N_1635,N_564);
xor U9802 (N_9802,N_2962,N_1288);
xnor U9803 (N_9803,N_3589,N_1843);
and U9804 (N_9804,N_3983,N_4477);
xnor U9805 (N_9805,N_373,N_4301);
nand U9806 (N_9806,N_2170,N_4908);
and U9807 (N_9807,N_2350,N_2381);
nand U9808 (N_9808,N_1723,N_2970);
nor U9809 (N_9809,N_2646,N_2343);
nor U9810 (N_9810,N_4831,N_2279);
nor U9811 (N_9811,N_3473,N_3899);
xor U9812 (N_9812,N_4004,N_970);
nor U9813 (N_9813,N_27,N_4298);
and U9814 (N_9814,N_1686,N_4470);
nor U9815 (N_9815,N_4434,N_1115);
or U9816 (N_9816,N_1129,N_723);
and U9817 (N_9817,N_2640,N_1721);
nand U9818 (N_9818,N_2804,N_1030);
and U9819 (N_9819,N_4397,N_904);
or U9820 (N_9820,N_4372,N_732);
nor U9821 (N_9821,N_131,N_4268);
nand U9822 (N_9822,N_4320,N_4216);
xnor U9823 (N_9823,N_2919,N_4606);
or U9824 (N_9824,N_3299,N_3816);
xnor U9825 (N_9825,N_933,N_1893);
nor U9826 (N_9826,N_4986,N_260);
and U9827 (N_9827,N_1653,N_687);
or U9828 (N_9828,N_4235,N_4898);
xnor U9829 (N_9829,N_2351,N_3058);
nor U9830 (N_9830,N_3716,N_2169);
or U9831 (N_9831,N_1070,N_1226);
and U9832 (N_9832,N_2125,N_344);
or U9833 (N_9833,N_3022,N_2333);
or U9834 (N_9834,N_4984,N_4046);
nor U9835 (N_9835,N_885,N_3602);
or U9836 (N_9836,N_4273,N_1502);
and U9837 (N_9837,N_4919,N_4999);
nand U9838 (N_9838,N_4677,N_4033);
nand U9839 (N_9839,N_2072,N_4649);
or U9840 (N_9840,N_39,N_948);
or U9841 (N_9841,N_2954,N_3852);
nand U9842 (N_9842,N_984,N_3452);
nor U9843 (N_9843,N_3934,N_3863);
and U9844 (N_9844,N_957,N_731);
or U9845 (N_9845,N_2790,N_689);
or U9846 (N_9846,N_2562,N_493);
nor U9847 (N_9847,N_1052,N_3002);
or U9848 (N_9848,N_639,N_3430);
nand U9849 (N_9849,N_2836,N_1309);
nand U9850 (N_9850,N_202,N_2000);
and U9851 (N_9851,N_4117,N_97);
and U9852 (N_9852,N_4407,N_3619);
xnor U9853 (N_9853,N_3666,N_4761);
and U9854 (N_9854,N_488,N_3517);
nand U9855 (N_9855,N_2308,N_1165);
xor U9856 (N_9856,N_425,N_340);
or U9857 (N_9857,N_1452,N_2496);
nand U9858 (N_9858,N_4610,N_787);
nand U9859 (N_9859,N_3101,N_3180);
nand U9860 (N_9860,N_3249,N_4387);
or U9861 (N_9861,N_1903,N_3832);
nor U9862 (N_9862,N_4513,N_1646);
nand U9863 (N_9863,N_3208,N_3959);
nor U9864 (N_9864,N_4255,N_2887);
or U9865 (N_9865,N_3098,N_4661);
nor U9866 (N_9866,N_4860,N_3746);
nor U9867 (N_9867,N_4,N_2440);
or U9868 (N_9868,N_2506,N_129);
xnor U9869 (N_9869,N_1044,N_1294);
nand U9870 (N_9870,N_4774,N_159);
nor U9871 (N_9871,N_2494,N_4601);
nand U9872 (N_9872,N_3447,N_4545);
nor U9873 (N_9873,N_4161,N_1148);
xnor U9874 (N_9874,N_66,N_1944);
or U9875 (N_9875,N_433,N_4886);
nor U9876 (N_9876,N_4508,N_3);
nor U9877 (N_9877,N_2210,N_3886);
or U9878 (N_9878,N_832,N_88);
nor U9879 (N_9879,N_3498,N_130);
nor U9880 (N_9880,N_4798,N_4140);
and U9881 (N_9881,N_4174,N_3453);
and U9882 (N_9882,N_3106,N_1672);
or U9883 (N_9883,N_10,N_581);
nand U9884 (N_9884,N_4234,N_271);
nor U9885 (N_9885,N_2680,N_2519);
and U9886 (N_9886,N_1661,N_1920);
nand U9887 (N_9887,N_2301,N_1753);
and U9888 (N_9888,N_2261,N_4050);
and U9889 (N_9889,N_2743,N_1309);
or U9890 (N_9890,N_1356,N_3053);
and U9891 (N_9891,N_1613,N_1954);
nand U9892 (N_9892,N_4398,N_2274);
and U9893 (N_9893,N_2335,N_2213);
xor U9894 (N_9894,N_2698,N_4793);
or U9895 (N_9895,N_212,N_2294);
nor U9896 (N_9896,N_4144,N_3740);
nand U9897 (N_9897,N_157,N_2530);
or U9898 (N_9898,N_2779,N_1613);
or U9899 (N_9899,N_2842,N_1569);
or U9900 (N_9900,N_1393,N_3934);
nor U9901 (N_9901,N_2171,N_3419);
or U9902 (N_9902,N_125,N_3417);
nand U9903 (N_9903,N_2506,N_2412);
and U9904 (N_9904,N_1878,N_2294);
nand U9905 (N_9905,N_230,N_4174);
nand U9906 (N_9906,N_4805,N_1157);
nand U9907 (N_9907,N_1234,N_1832);
xnor U9908 (N_9908,N_3071,N_2100);
or U9909 (N_9909,N_3417,N_1675);
nor U9910 (N_9910,N_1513,N_3915);
and U9911 (N_9911,N_1618,N_980);
xor U9912 (N_9912,N_880,N_4406);
nor U9913 (N_9913,N_1138,N_2652);
nor U9914 (N_9914,N_4062,N_1441);
or U9915 (N_9915,N_1397,N_3764);
or U9916 (N_9916,N_389,N_935);
and U9917 (N_9917,N_4333,N_2594);
nand U9918 (N_9918,N_2783,N_1015);
nand U9919 (N_9919,N_3013,N_3438);
and U9920 (N_9920,N_995,N_4451);
or U9921 (N_9921,N_3111,N_3996);
and U9922 (N_9922,N_3846,N_3778);
or U9923 (N_9923,N_4747,N_2874);
nor U9924 (N_9924,N_828,N_3572);
and U9925 (N_9925,N_3873,N_4687);
and U9926 (N_9926,N_78,N_3463);
or U9927 (N_9927,N_708,N_4419);
nand U9928 (N_9928,N_4114,N_169);
and U9929 (N_9929,N_3821,N_3701);
and U9930 (N_9930,N_761,N_159);
nor U9931 (N_9931,N_889,N_579);
nor U9932 (N_9932,N_407,N_3981);
and U9933 (N_9933,N_4570,N_3913);
xor U9934 (N_9934,N_1699,N_66);
nand U9935 (N_9935,N_4742,N_1241);
nand U9936 (N_9936,N_2730,N_4548);
nor U9937 (N_9937,N_4369,N_1529);
nand U9938 (N_9938,N_4536,N_4394);
or U9939 (N_9939,N_221,N_2532);
nor U9940 (N_9940,N_4030,N_3166);
nor U9941 (N_9941,N_4594,N_741);
or U9942 (N_9942,N_4029,N_1552);
and U9943 (N_9943,N_2380,N_602);
or U9944 (N_9944,N_673,N_541);
and U9945 (N_9945,N_550,N_1734);
and U9946 (N_9946,N_4128,N_2219);
or U9947 (N_9947,N_1235,N_2777);
or U9948 (N_9948,N_3848,N_1642);
nand U9949 (N_9949,N_4674,N_3207);
nor U9950 (N_9950,N_2127,N_2368);
and U9951 (N_9951,N_4659,N_3426);
and U9952 (N_9952,N_2678,N_1959);
or U9953 (N_9953,N_2055,N_3366);
and U9954 (N_9954,N_1747,N_1786);
and U9955 (N_9955,N_3608,N_1420);
and U9956 (N_9956,N_1015,N_3156);
xor U9957 (N_9957,N_498,N_1352);
and U9958 (N_9958,N_2892,N_2258);
and U9959 (N_9959,N_4853,N_1716);
nor U9960 (N_9960,N_4876,N_907);
nor U9961 (N_9961,N_4818,N_1236);
or U9962 (N_9962,N_3437,N_835);
or U9963 (N_9963,N_3264,N_403);
nand U9964 (N_9964,N_540,N_2253);
nor U9965 (N_9965,N_318,N_1472);
or U9966 (N_9966,N_839,N_927);
and U9967 (N_9967,N_3527,N_226);
or U9968 (N_9968,N_4272,N_4358);
nand U9969 (N_9969,N_2555,N_4096);
nand U9970 (N_9970,N_4370,N_1515);
nor U9971 (N_9971,N_1176,N_2082);
or U9972 (N_9972,N_2215,N_4017);
nor U9973 (N_9973,N_4168,N_2683);
nor U9974 (N_9974,N_2090,N_2720);
or U9975 (N_9975,N_3835,N_3364);
nor U9976 (N_9976,N_708,N_357);
or U9977 (N_9977,N_1456,N_1385);
and U9978 (N_9978,N_1320,N_4978);
or U9979 (N_9979,N_721,N_4071);
and U9980 (N_9980,N_2933,N_4576);
nor U9981 (N_9981,N_2453,N_1879);
nor U9982 (N_9982,N_1619,N_680);
and U9983 (N_9983,N_3680,N_2214);
and U9984 (N_9984,N_1919,N_490);
nor U9985 (N_9985,N_1040,N_2793);
nand U9986 (N_9986,N_4602,N_650);
nand U9987 (N_9987,N_4439,N_4893);
and U9988 (N_9988,N_1425,N_1569);
or U9989 (N_9989,N_1369,N_592);
or U9990 (N_9990,N_3116,N_1114);
or U9991 (N_9991,N_3990,N_2049);
nand U9992 (N_9992,N_3031,N_4618);
xor U9993 (N_9993,N_3654,N_2366);
and U9994 (N_9994,N_1078,N_545);
nor U9995 (N_9995,N_99,N_916);
nand U9996 (N_9996,N_2280,N_3513);
and U9997 (N_9997,N_4950,N_626);
nor U9998 (N_9998,N_1320,N_2970);
or U9999 (N_9999,N_1510,N_2148);
nor U10000 (N_10000,N_5898,N_7404);
nand U10001 (N_10001,N_6915,N_5423);
nand U10002 (N_10002,N_6165,N_9591);
nand U10003 (N_10003,N_5402,N_5712);
and U10004 (N_10004,N_5366,N_9836);
nand U10005 (N_10005,N_8580,N_5939);
nor U10006 (N_10006,N_5320,N_8631);
nand U10007 (N_10007,N_5624,N_6827);
and U10008 (N_10008,N_7325,N_7954);
xnor U10009 (N_10009,N_7651,N_8805);
or U10010 (N_10010,N_6509,N_9873);
and U10011 (N_10011,N_8473,N_5830);
nand U10012 (N_10012,N_8526,N_5225);
and U10013 (N_10013,N_5273,N_8585);
nand U10014 (N_10014,N_8405,N_7435);
nand U10015 (N_10015,N_5767,N_5504);
and U10016 (N_10016,N_8141,N_7291);
nand U10017 (N_10017,N_6271,N_8480);
xor U10018 (N_10018,N_5622,N_7851);
or U10019 (N_10019,N_5936,N_8911);
and U10020 (N_10020,N_6201,N_9973);
nand U10021 (N_10021,N_6280,N_8926);
xor U10022 (N_10022,N_5294,N_6313);
nand U10023 (N_10023,N_9530,N_9070);
or U10024 (N_10024,N_9512,N_6823);
and U10025 (N_10025,N_9649,N_7332);
or U10026 (N_10026,N_6939,N_7159);
and U10027 (N_10027,N_5647,N_8668);
or U10028 (N_10028,N_7657,N_8536);
or U10029 (N_10029,N_5508,N_5006);
nor U10030 (N_10030,N_8535,N_6183);
nand U10031 (N_10031,N_9273,N_8037);
or U10032 (N_10032,N_8324,N_5568);
or U10033 (N_10033,N_8080,N_8571);
and U10034 (N_10034,N_6391,N_9449);
or U10035 (N_10035,N_6738,N_9738);
nor U10036 (N_10036,N_9984,N_6488);
and U10037 (N_10037,N_5535,N_8666);
and U10038 (N_10038,N_7192,N_7044);
nand U10039 (N_10039,N_8837,N_8913);
or U10040 (N_10040,N_5334,N_8378);
nor U10041 (N_10041,N_8552,N_7683);
or U10042 (N_10042,N_6261,N_5292);
nand U10043 (N_10043,N_5884,N_9233);
nand U10044 (N_10044,N_8295,N_6906);
nand U10045 (N_10045,N_6769,N_7284);
nor U10046 (N_10046,N_6722,N_9025);
or U10047 (N_10047,N_8395,N_5408);
or U10048 (N_10048,N_8776,N_5598);
nor U10049 (N_10049,N_6188,N_7925);
nand U10050 (N_10050,N_6283,N_5077);
or U10051 (N_10051,N_9138,N_7521);
nor U10052 (N_10052,N_9995,N_6500);
or U10053 (N_10053,N_8732,N_9797);
and U10054 (N_10054,N_9952,N_8073);
nand U10055 (N_10055,N_5527,N_8112);
and U10056 (N_10056,N_8312,N_7956);
nand U10057 (N_10057,N_7005,N_7022);
or U10058 (N_10058,N_5432,N_5836);
and U10059 (N_10059,N_8787,N_7275);
nand U10060 (N_10060,N_6403,N_7273);
xnor U10061 (N_10061,N_5957,N_7343);
nor U10062 (N_10062,N_9764,N_6886);
nand U10063 (N_10063,N_7002,N_9661);
xnor U10064 (N_10064,N_7514,N_7142);
and U10065 (N_10065,N_9859,N_8968);
nor U10066 (N_10066,N_6426,N_8916);
and U10067 (N_10067,N_8772,N_8649);
nor U10068 (N_10068,N_9168,N_6756);
xnor U10069 (N_10069,N_6636,N_8306);
nand U10070 (N_10070,N_9595,N_8276);
nand U10071 (N_10071,N_6366,N_6585);
and U10072 (N_10072,N_8903,N_6067);
nor U10073 (N_10073,N_8232,N_5361);
nor U10074 (N_10074,N_9183,N_9906);
or U10075 (N_10075,N_6536,N_5411);
xnor U10076 (N_10076,N_5026,N_9151);
nor U10077 (N_10077,N_7049,N_9035);
nor U10078 (N_10078,N_8368,N_8716);
and U10079 (N_10079,N_8163,N_7035);
xor U10080 (N_10080,N_7759,N_7852);
xor U10081 (N_10081,N_9781,N_7638);
nand U10082 (N_10082,N_8385,N_5515);
nand U10083 (N_10083,N_6332,N_8231);
nor U10084 (N_10084,N_5671,N_9248);
nand U10085 (N_10085,N_8981,N_8660);
or U10086 (N_10086,N_9976,N_8407);
nor U10087 (N_10087,N_7277,N_7983);
and U10088 (N_10088,N_6777,N_7562);
or U10089 (N_10089,N_9135,N_6846);
and U10090 (N_10090,N_7179,N_9754);
or U10091 (N_10091,N_5639,N_7635);
nand U10092 (N_10092,N_5770,N_5253);
nand U10093 (N_10093,N_5759,N_5742);
nor U10094 (N_10094,N_8778,N_9324);
nor U10095 (N_10095,N_6760,N_9852);
nand U10096 (N_10096,N_8083,N_8203);
nor U10097 (N_10097,N_9706,N_6184);
or U10098 (N_10098,N_6033,N_5463);
and U10099 (N_10099,N_8710,N_8410);
nor U10100 (N_10100,N_9089,N_5344);
or U10101 (N_10101,N_5016,N_5410);
and U10102 (N_10102,N_9721,N_6074);
nor U10103 (N_10103,N_5843,N_8643);
and U10104 (N_10104,N_9670,N_8010);
or U10105 (N_10105,N_6304,N_6057);
nand U10106 (N_10106,N_5701,N_7898);
or U10107 (N_10107,N_7783,N_5386);
and U10108 (N_10108,N_7381,N_8792);
xnor U10109 (N_10109,N_8576,N_9621);
or U10110 (N_10110,N_8977,N_7459);
or U10111 (N_10111,N_8542,N_6264);
or U10112 (N_10112,N_9300,N_5905);
and U10113 (N_10113,N_9014,N_5125);
nor U10114 (N_10114,N_9407,N_5858);
nand U10115 (N_10115,N_9559,N_9175);
and U10116 (N_10116,N_8558,N_5157);
xor U10117 (N_10117,N_5699,N_8985);
and U10118 (N_10118,N_5660,N_6737);
nor U10119 (N_10119,N_9839,N_9954);
and U10120 (N_10120,N_5771,N_8097);
and U10121 (N_10121,N_6808,N_6071);
or U10122 (N_10122,N_9096,N_9685);
or U10123 (N_10123,N_7344,N_5246);
nor U10124 (N_10124,N_6592,N_8744);
nand U10125 (N_10125,N_5618,N_7437);
or U10126 (N_10126,N_7556,N_7874);
nor U10127 (N_10127,N_7861,N_8548);
nor U10128 (N_10128,N_5669,N_8109);
nand U10129 (N_10129,N_5638,N_8415);
nor U10130 (N_10130,N_5749,N_9130);
nor U10131 (N_10131,N_5807,N_5585);
and U10132 (N_10132,N_8742,N_5126);
or U10133 (N_10133,N_9226,N_6819);
xnor U10134 (N_10134,N_6344,N_7242);
nor U10135 (N_10135,N_7014,N_9520);
nor U10136 (N_10136,N_5740,N_9101);
and U10137 (N_10137,N_7485,N_7848);
and U10138 (N_10138,N_6387,N_8884);
and U10139 (N_10139,N_6618,N_9994);
nand U10140 (N_10140,N_8628,N_8507);
or U10141 (N_10141,N_5043,N_6217);
and U10142 (N_10142,N_7228,N_5391);
and U10143 (N_10143,N_8294,N_9056);
nor U10144 (N_10144,N_5708,N_6407);
and U10145 (N_10145,N_8618,N_9467);
or U10146 (N_10146,N_7553,N_9710);
or U10147 (N_10147,N_6853,N_5162);
nor U10148 (N_10148,N_5730,N_9869);
and U10149 (N_10149,N_7055,N_6900);
and U10150 (N_10150,N_7483,N_5722);
or U10151 (N_10151,N_8070,N_7705);
nand U10152 (N_10152,N_7924,N_9214);
nor U10153 (N_10153,N_7955,N_5227);
and U10154 (N_10154,N_9480,N_9321);
nor U10155 (N_10155,N_8960,N_6158);
nand U10156 (N_10156,N_9374,N_7109);
and U10157 (N_10157,N_9156,N_5626);
and U10158 (N_10158,N_9126,N_9526);
nor U10159 (N_10159,N_9543,N_5677);
nor U10160 (N_10160,N_6685,N_8088);
nor U10161 (N_10161,N_5780,N_5909);
or U10162 (N_10162,N_8767,N_5890);
and U10163 (N_10163,N_6087,N_5746);
xor U10164 (N_10164,N_7588,N_6671);
nand U10165 (N_10165,N_7658,N_5089);
nand U10166 (N_10166,N_9609,N_8586);
and U10167 (N_10167,N_8713,N_9337);
nor U10168 (N_10168,N_8734,N_5500);
or U10169 (N_10169,N_7775,N_8557);
nand U10170 (N_10170,N_8430,N_8756);
or U10171 (N_10171,N_5260,N_7021);
nand U10172 (N_10172,N_7127,N_6386);
nor U10173 (N_10173,N_6883,N_6098);
nand U10174 (N_10174,N_8028,N_6953);
or U10175 (N_10175,N_9692,N_9680);
or U10176 (N_10176,N_7555,N_5002);
nand U10177 (N_10177,N_9004,N_7686);
or U10178 (N_10178,N_9483,N_7152);
or U10179 (N_10179,N_9338,N_7252);
and U10180 (N_10180,N_8174,N_7356);
nand U10181 (N_10181,N_8326,N_8269);
or U10182 (N_10182,N_6935,N_5897);
nor U10183 (N_10183,N_6330,N_7517);
nand U10184 (N_10184,N_8371,N_6113);
nand U10185 (N_10185,N_8244,N_5584);
and U10186 (N_10186,N_7372,N_5078);
and U10187 (N_10187,N_8741,N_5529);
nor U10188 (N_10188,N_8945,N_5203);
nand U10189 (N_10189,N_6754,N_6944);
or U10190 (N_10190,N_8328,N_8384);
or U10191 (N_10191,N_9511,N_8450);
xor U10192 (N_10192,N_5088,N_9644);
and U10193 (N_10193,N_7479,N_7505);
and U10194 (N_10194,N_9770,N_8360);
xor U10195 (N_10195,N_8357,N_5952);
xor U10196 (N_10196,N_5844,N_9768);
nor U10197 (N_10197,N_9345,N_8991);
nor U10198 (N_10198,N_9555,N_7977);
nor U10199 (N_10199,N_7672,N_8655);
xor U10200 (N_10200,N_7026,N_7173);
or U10201 (N_10201,N_8501,N_6502);
nand U10202 (N_10202,N_5766,N_5921);
and U10203 (N_10203,N_9411,N_6894);
and U10204 (N_10204,N_8892,N_7432);
nand U10205 (N_10205,N_8342,N_5044);
nand U10206 (N_10206,N_5847,N_5673);
nor U10207 (N_10207,N_5631,N_5062);
and U10208 (N_10208,N_6416,N_9794);
or U10209 (N_10209,N_7659,N_6861);
nor U10210 (N_10210,N_7218,N_8252);
nand U10211 (N_10211,N_5978,N_8305);
and U10212 (N_10212,N_5916,N_8139);
xnor U10213 (N_10213,N_7605,N_8162);
xnor U10214 (N_10214,N_9748,N_7897);
xor U10215 (N_10215,N_9729,N_9416);
or U10216 (N_10216,N_6520,N_6637);
nor U10217 (N_10217,N_8086,N_9351);
and U10218 (N_10218,N_8504,N_7757);
nor U10219 (N_10219,N_7393,N_8952);
nand U10220 (N_10220,N_6784,N_6958);
nor U10221 (N_10221,N_7177,N_8498);
nand U10222 (N_10222,N_7311,N_9785);
nor U10223 (N_10223,N_9594,N_9572);
nand U10224 (N_10224,N_7374,N_9563);
xor U10225 (N_10225,N_6718,N_6879);
nand U10226 (N_10226,N_5656,N_8486);
xor U10227 (N_10227,N_5054,N_8370);
nand U10228 (N_10228,N_8137,N_6736);
or U10229 (N_10229,N_6952,N_9801);
nand U10230 (N_10230,N_8191,N_5946);
and U10231 (N_10231,N_7515,N_6367);
nand U10232 (N_10232,N_8811,N_9016);
or U10233 (N_10233,N_9390,N_9971);
nand U10234 (N_10234,N_8158,N_9205);
nor U10235 (N_10235,N_8715,N_5851);
nor U10236 (N_10236,N_9335,N_9931);
nand U10237 (N_10237,N_6447,N_9082);
nand U10238 (N_10238,N_6216,N_8213);
and U10239 (N_10239,N_6762,N_6845);
or U10240 (N_10240,N_6035,N_6405);
and U10241 (N_10241,N_7737,N_5537);
or U10242 (N_10242,N_6936,N_7592);
nand U10243 (N_10243,N_7265,N_6943);
and U10244 (N_10244,N_9499,N_8914);
xor U10245 (N_10245,N_6663,N_9157);
nand U10246 (N_10246,N_6088,N_9777);
or U10247 (N_10247,N_7742,N_7357);
nand U10248 (N_10248,N_7354,N_7087);
nor U10249 (N_10249,N_7774,N_9241);
nor U10250 (N_10250,N_8878,N_7497);
nand U10251 (N_10251,N_6634,N_5630);
nor U10252 (N_10252,N_9421,N_7153);
and U10253 (N_10253,N_9478,N_7348);
nor U10254 (N_10254,N_5961,N_9492);
and U10255 (N_10255,N_9534,N_7476);
or U10256 (N_10256,N_9033,N_5892);
nand U10257 (N_10257,N_8671,N_9367);
and U10258 (N_10258,N_6335,N_7099);
and U10259 (N_10259,N_5931,N_8506);
and U10260 (N_10260,N_7887,N_9034);
nor U10261 (N_10261,N_6907,N_7091);
and U10262 (N_10262,N_8856,N_6695);
or U10263 (N_10263,N_7712,N_7602);
nand U10264 (N_10264,N_6550,N_8390);
or U10265 (N_10265,N_9115,N_6160);
or U10266 (N_10266,N_8531,N_5238);
nor U10267 (N_10267,N_5610,N_6253);
and U10268 (N_10268,N_9602,N_7254);
xnor U10269 (N_10269,N_7560,N_5676);
nor U10270 (N_10270,N_7756,N_8169);
or U10271 (N_10271,N_9845,N_7798);
and U10272 (N_10272,N_8271,N_6558);
xor U10273 (N_10273,N_7895,N_9514);
or U10274 (N_10274,N_5335,N_5325);
and U10275 (N_10275,N_9074,N_6013);
nand U10276 (N_10276,N_7030,N_5517);
xor U10277 (N_10277,N_9604,N_5367);
nor U10278 (N_10278,N_6123,N_8565);
nor U10279 (N_10279,N_7965,N_8898);
xnor U10280 (N_10280,N_6593,N_5095);
nand U10281 (N_10281,N_8115,N_8893);
nand U10282 (N_10282,N_9732,N_5231);
nor U10283 (N_10283,N_8561,N_8841);
nor U10284 (N_10284,N_9872,N_5982);
xnor U10285 (N_10285,N_6290,N_8662);
or U10286 (N_10286,N_8608,N_6034);
xnor U10287 (N_10287,N_8197,N_6638);
nand U10288 (N_10288,N_9395,N_6022);
nand U10289 (N_10289,N_8211,N_7542);
nand U10290 (N_10290,N_9036,N_5101);
xor U10291 (N_10291,N_9160,N_8796);
or U10292 (N_10292,N_8095,N_9122);
nand U10293 (N_10293,N_9786,N_6857);
nand U10294 (N_10294,N_7201,N_9718);
nor U10295 (N_10295,N_6453,N_9775);
or U10296 (N_10296,N_8301,N_9981);
or U10297 (N_10297,N_6969,N_8052);
nor U10298 (N_10298,N_8094,N_9114);
nor U10299 (N_10299,N_5655,N_9857);
and U10300 (N_10300,N_7629,N_6246);
and U10301 (N_10301,N_7362,N_8079);
nand U10302 (N_10302,N_5969,N_8014);
and U10303 (N_10303,N_6941,N_7386);
nor U10304 (N_10304,N_5204,N_8067);
nor U10305 (N_10305,N_6309,N_6462);
and U10306 (N_10306,N_9593,N_9784);
or U10307 (N_10307,N_5663,N_5450);
and U10308 (N_10308,N_6270,N_9856);
nand U10309 (N_10309,N_7175,N_5876);
or U10310 (N_10310,N_6122,N_5802);
xnor U10311 (N_10311,N_9366,N_9540);
xor U10312 (N_10312,N_6968,N_7586);
or U10313 (N_10313,N_9332,N_8569);
xnor U10314 (N_10314,N_8516,N_9057);
nand U10315 (N_10315,N_6965,N_6373);
xor U10316 (N_10316,N_9454,N_8277);
or U10317 (N_10317,N_7241,N_9817);
nor U10318 (N_10318,N_7624,N_8427);
nor U10319 (N_10319,N_5181,N_8147);
or U10320 (N_10320,N_7538,N_9271);
nor U10321 (N_10321,N_6006,N_9686);
or U10322 (N_10322,N_5865,N_8915);
nor U10323 (N_10323,N_7917,N_6901);
nand U10324 (N_10324,N_7680,N_8381);
and U10325 (N_10325,N_7844,N_8566);
nand U10326 (N_10326,N_7569,N_5154);
nor U10327 (N_10327,N_5736,N_8989);
nor U10328 (N_10328,N_5400,N_6202);
nor U10329 (N_10329,N_5454,N_6241);
nand U10330 (N_10330,N_6070,N_6279);
and U10331 (N_10331,N_5464,N_9296);
nand U10332 (N_10332,N_5904,N_8352);
and U10333 (N_10333,N_5670,N_9422);
or U10334 (N_10334,N_8829,N_6112);
or U10335 (N_10335,N_9245,N_6099);
or U10336 (N_10336,N_5321,N_8921);
and U10337 (N_10337,N_7987,N_6037);
nor U10338 (N_10338,N_5922,N_6404);
nand U10339 (N_10339,N_6859,N_8283);
and U10340 (N_10340,N_9268,N_8265);
or U10341 (N_10341,N_6233,N_5314);
nand U10342 (N_10342,N_7707,N_5903);
nor U10343 (N_10343,N_8515,N_8600);
xor U10344 (N_10344,N_7663,N_7670);
nor U10345 (N_10345,N_5439,N_8555);
or U10346 (N_10346,N_9368,N_5451);
xnor U10347 (N_10347,N_6889,N_6480);
nor U10348 (N_10348,N_5490,N_9923);
nand U10349 (N_10349,N_5561,N_6009);
nor U10350 (N_10350,N_8857,N_9633);
and U10351 (N_10351,N_6972,N_8383);
nand U10352 (N_10352,N_7527,N_5689);
nand U10353 (N_10353,N_6337,N_7306);
nor U10354 (N_10354,N_8821,N_7340);
nand U10355 (N_10355,N_9556,N_8118);
and U10356 (N_10356,N_9714,N_8938);
and U10357 (N_10357,N_8361,N_8809);
nor U10358 (N_10358,N_7655,N_6244);
and U10359 (N_10359,N_7984,N_7610);
or U10360 (N_10360,N_7979,N_5359);
nand U10361 (N_10361,N_5681,N_7346);
or U10362 (N_10362,N_7056,N_7577);
nor U10363 (N_10363,N_6951,N_9146);
or U10364 (N_10364,N_6862,N_5236);
and U10365 (N_10365,N_9145,N_9805);
nand U10366 (N_10366,N_6641,N_5661);
nand U10367 (N_10367,N_8359,N_6397);
nor U10368 (N_10368,N_6564,N_6997);
and U10369 (N_10369,N_8847,N_5682);
nand U10370 (N_10370,N_7564,N_8138);
and U10371 (N_10371,N_9796,N_5710);
nand U10372 (N_10372,N_8661,N_9711);
or U10373 (N_10373,N_7631,N_8044);
or U10374 (N_10374,N_6927,N_9547);
and U10375 (N_10375,N_6491,N_8177);
and U10376 (N_10376,N_6154,N_7143);
and U10377 (N_10377,N_6227,N_7043);
nor U10378 (N_10378,N_7788,N_8313);
xor U10379 (N_10379,N_8433,N_6798);
or U10380 (N_10380,N_8492,N_5816);
and U10381 (N_10381,N_6025,N_7991);
xor U10382 (N_10382,N_7807,N_5139);
or U10383 (N_10383,N_6041,N_6702);
or U10384 (N_10384,N_5243,N_8988);
or U10385 (N_10385,N_5199,N_6733);
nor U10386 (N_10386,N_6414,N_7268);
nand U10387 (N_10387,N_7383,N_9278);
and U10388 (N_10388,N_6501,N_9780);
and U10389 (N_10389,N_6306,N_6623);
and U10390 (N_10390,N_6323,N_7523);
and U10391 (N_10391,N_8338,N_7941);
nor U10392 (N_10392,N_5611,N_5857);
and U10393 (N_10393,N_9200,N_6069);
or U10394 (N_10394,N_7040,N_6785);
nand U10395 (N_10395,N_7571,N_7008);
or U10396 (N_10396,N_8794,N_6434);
nand U10397 (N_10397,N_5316,N_7349);
xnor U10398 (N_10398,N_7596,N_9837);
xnor U10399 (N_10399,N_6869,N_7981);
xnor U10400 (N_10400,N_7978,N_9531);
nand U10401 (N_10401,N_5440,N_6913);
nand U10402 (N_10402,N_8899,N_5853);
nor U10403 (N_10403,N_6223,N_6989);
nor U10404 (N_10404,N_5113,N_9590);
or U10405 (N_10405,N_8309,N_8148);
and U10406 (N_10406,N_8454,N_8534);
or U10407 (N_10407,N_5473,N_6175);
and U10408 (N_10408,N_7454,N_5972);
nor U10409 (N_10409,N_5553,N_7801);
or U10410 (N_10410,N_9106,N_8520);
xor U10411 (N_10411,N_7846,N_9677);
xor U10412 (N_10412,N_8860,N_6127);
and U10413 (N_10413,N_7666,N_6342);
and U10414 (N_10414,N_8564,N_8285);
nor U10415 (N_10415,N_5901,N_7760);
and U10416 (N_10416,N_6720,N_5239);
or U10417 (N_10417,N_8701,N_7029);
xor U10418 (N_10418,N_7235,N_8425);
and U10419 (N_10419,N_6432,N_5188);
or U10420 (N_10420,N_7964,N_7295);
nand U10421 (N_10421,N_8582,N_9398);
nor U10422 (N_10422,N_8084,N_8196);
xnor U10423 (N_10423,N_5118,N_9588);
xnor U10424 (N_10424,N_6855,N_9210);
xor U10425 (N_10425,N_9452,N_9155);
and U10426 (N_10426,N_9538,N_9829);
or U10427 (N_10427,N_5434,N_8245);
and U10428 (N_10428,N_7949,N_8749);
nand U10429 (N_10429,N_6884,N_9149);
or U10430 (N_10430,N_8961,N_8472);
nand U10431 (N_10431,N_5397,N_6640);
nor U10432 (N_10432,N_5202,N_6131);
or U10433 (N_10433,N_5613,N_7758);
and U10434 (N_10434,N_7085,N_6851);
nor U10435 (N_10435,N_7723,N_8999);
or U10436 (N_10436,N_6818,N_6679);
nor U10437 (N_10437,N_9958,N_8268);
nor U10438 (N_10438,N_8474,N_9095);
nand U10439 (N_10439,N_8842,N_6716);
nor U10440 (N_10440,N_9725,N_5412);
or U10441 (N_10441,N_9884,N_6826);
nand U10442 (N_10442,N_9447,N_6990);
nor U10443 (N_10443,N_8752,N_6214);
xor U10444 (N_10444,N_8559,N_7628);
nand U10445 (N_10445,N_9341,N_7989);
nor U10446 (N_10446,N_6003,N_6780);
nand U10447 (N_10447,N_9651,N_6504);
nand U10448 (N_10448,N_9654,N_9440);
and U10449 (N_10449,N_9652,N_7077);
and U10450 (N_10450,N_5237,N_5284);
or U10451 (N_10451,N_9026,N_6800);
xor U10452 (N_10452,N_7208,N_5538);
nand U10453 (N_10453,N_7111,N_5667);
nand U10454 (N_10454,N_5606,N_5407);
nor U10455 (N_10455,N_8834,N_9254);
xor U10456 (N_10456,N_8704,N_6940);
nor U10457 (N_10457,N_9825,N_9349);
nor U10458 (N_10458,N_5045,N_7431);
and U10459 (N_10459,N_5801,N_9892);
nand U10460 (N_10460,N_9433,N_5652);
nor U10461 (N_10461,N_6143,N_7271);
nand U10462 (N_10462,N_8895,N_6456);
and U10463 (N_10463,N_7168,N_6863);
and U10464 (N_10464,N_8615,N_8619);
xnor U10465 (N_10465,N_7122,N_8868);
and U10466 (N_10466,N_6840,N_9667);
nand U10467 (N_10467,N_8060,N_9935);
and U10468 (N_10468,N_5992,N_8270);
and U10469 (N_10469,N_7997,N_7973);
or U10470 (N_10470,N_7699,N_5342);
xnor U10471 (N_10471,N_6082,N_9678);
nor U10472 (N_10472,N_9740,N_7191);
or U10473 (N_10473,N_8578,N_8397);
and U10474 (N_10474,N_5988,N_9250);
nor U10475 (N_10475,N_8172,N_5594);
nand U10476 (N_10476,N_9075,N_9955);
and U10477 (N_10477,N_5797,N_5184);
xor U10478 (N_10478,N_6834,N_5696);
nor U10479 (N_10479,N_7512,N_8765);
nor U10480 (N_10480,N_5443,N_7442);
nand U10481 (N_10481,N_7833,N_7802);
nor U10482 (N_10482,N_7425,N_9355);
nand U10483 (N_10483,N_7752,N_8388);
or U10484 (N_10484,N_6522,N_9989);
nand U10485 (N_10485,N_7229,N_6905);
and U10486 (N_10486,N_5629,N_5825);
nand U10487 (N_10487,N_9133,N_7713);
nand U10488 (N_10488,N_5793,N_9871);
xnor U10489 (N_10489,N_9207,N_9119);
or U10490 (N_10490,N_9013,N_7953);
nor U10491 (N_10491,N_8862,N_8062);
or U10492 (N_10492,N_9039,N_6329);
xnor U10493 (N_10493,N_6556,N_8702);
nor U10494 (N_10494,N_7970,N_7183);
nor U10495 (N_10495,N_6612,N_7767);
xor U10496 (N_10496,N_7006,N_9097);
and U10497 (N_10497,N_6530,N_7826);
xnor U10498 (N_10498,N_7836,N_7509);
or U10499 (N_10499,N_9282,N_5530);
or U10500 (N_10500,N_8250,N_7656);
nor U10501 (N_10501,N_7104,N_8613);
nand U10502 (N_10502,N_7821,N_7793);
and U10503 (N_10503,N_8403,N_9635);
or U10504 (N_10504,N_8077,N_8743);
nor U10505 (N_10505,N_9808,N_6212);
and U10506 (N_10506,N_9410,N_8646);
or U10507 (N_10507,N_8836,N_6059);
nor U10508 (N_10508,N_8761,N_9311);
and U10509 (N_10509,N_6413,N_5798);
and U10510 (N_10510,N_9877,N_6169);
nand U10511 (N_10511,N_9170,N_8828);
and U10512 (N_10512,N_9788,N_9011);
nor U10513 (N_10513,N_6820,N_8350);
and U10514 (N_10514,N_7028,N_7722);
nand U10515 (N_10515,N_5910,N_7715);
nor U10516 (N_10516,N_9589,N_9596);
nand U10517 (N_10517,N_8050,N_8645);
nand U10518 (N_10518,N_6608,N_8670);
or U10519 (N_10519,N_9949,N_7999);
and U10520 (N_10520,N_5487,N_5233);
and U10521 (N_10521,N_8007,N_8399);
nand U10522 (N_10522,N_7450,N_5595);
nor U10523 (N_10523,N_7041,N_9838);
or U10524 (N_10524,N_8820,N_9629);
or U10525 (N_10525,N_8344,N_6433);
nand U10526 (N_10526,N_6492,N_9045);
nand U10527 (N_10527,N_8194,N_9319);
and U10528 (N_10528,N_5385,N_8438);
nor U10529 (N_10529,N_6828,N_5186);
xnor U10530 (N_10530,N_7345,N_9578);
and U10531 (N_10531,N_9018,N_8103);
or U10532 (N_10532,N_6847,N_5923);
or U10533 (N_10533,N_7779,N_9079);
xor U10534 (N_10534,N_8008,N_6963);
or U10535 (N_10535,N_9587,N_5037);
nor U10536 (N_10536,N_7888,N_7169);
or U10537 (N_10537,N_6801,N_9361);
and U10538 (N_10538,N_6412,N_5588);
xnor U10539 (N_10539,N_8426,N_9966);
nor U10540 (N_10540,N_6930,N_5688);
and U10541 (N_10541,N_6740,N_9929);
nand U10542 (N_10542,N_9350,N_7012);
and U10543 (N_10543,N_5330,N_7632);
nor U10544 (N_10544,N_8192,N_5761);
and U10545 (N_10545,N_6029,N_8993);
xnor U10546 (N_10546,N_8807,N_5729);
and U10547 (N_10547,N_6186,N_5861);
or U10548 (N_10548,N_5305,N_6476);
or U10549 (N_10549,N_9123,N_7777);
nor U10550 (N_10550,N_6288,N_5286);
nand U10551 (N_10551,N_5963,N_7734);
nand U10552 (N_10552,N_9102,N_9462);
xnor U10553 (N_10553,N_8747,N_5480);
xor U10554 (N_10554,N_6892,N_5545);
and U10555 (N_10555,N_8046,N_5945);
and U10556 (N_10556,N_8240,N_7210);
and U10557 (N_10557,N_7580,N_5250);
or U10558 (N_10558,N_7667,N_5634);
nand U10559 (N_10559,N_5651,N_7901);
xnor U10560 (N_10560,N_6483,N_8524);
and U10561 (N_10561,N_6683,N_5229);
nor U10562 (N_10562,N_9585,N_7186);
nand U10563 (N_10563,N_7245,N_8036);
nor U10564 (N_10564,N_5781,N_9864);
or U10565 (N_10565,N_8880,N_6804);
nor U10566 (N_10566,N_5031,N_8461);
nor U10567 (N_10567,N_7859,N_9281);
or U10568 (N_10568,N_5213,N_6409);
nor U10569 (N_10569,N_7118,N_5547);
nor U10570 (N_10570,N_5422,N_6277);
nand U10571 (N_10571,N_9072,N_8708);
nor U10572 (N_10572,N_6726,N_8614);
nor U10573 (N_10573,N_9807,N_5557);
nor U10574 (N_10574,N_8266,N_5068);
and U10575 (N_10575,N_7766,N_6163);
nor U10576 (N_10576,N_8248,N_7320);
nand U10577 (N_10577,N_9258,N_6810);
xor U10578 (N_10578,N_6377,N_8341);
nand U10579 (N_10579,N_7661,N_7335);
or U10580 (N_10580,N_9299,N_9854);
nor U10581 (N_10581,N_5970,N_9608);
and U10582 (N_10582,N_8258,N_7815);
and U10583 (N_10583,N_8042,N_5525);
and U10584 (N_10584,N_6945,N_5441);
nand U10585 (N_10585,N_6717,N_9498);
or U10586 (N_10586,N_8372,N_5519);
nand U10587 (N_10587,N_9021,N_5999);
nand U10588 (N_10588,N_7379,N_8065);
nand U10589 (N_10589,N_9795,N_5262);
and U10590 (N_10590,N_7504,N_9674);
nor U10591 (N_10591,N_8358,N_7135);
nor U10592 (N_10592,N_7967,N_6417);
nor U10593 (N_10593,N_6466,N_8105);
nor U10594 (N_10594,N_6027,N_6966);
nand U10595 (N_10595,N_6515,N_5476);
nand U10596 (N_10596,N_7297,N_9752);
nor U10597 (N_10597,N_9178,N_8303);
or U10598 (N_10598,N_6100,N_9793);
nor U10599 (N_10599,N_9548,N_9461);
xor U10600 (N_10600,N_6644,N_9519);
nor U10601 (N_10601,N_9662,N_9309);
nand U10602 (N_10602,N_9235,N_7176);
and U10603 (N_10603,N_6693,N_5339);
or U10604 (N_10604,N_5586,N_9848);
xnor U10605 (N_10605,N_6727,N_6506);
nor U10606 (N_10606,N_7544,N_5326);
or U10607 (N_10607,N_5570,N_8373);
nand U10608 (N_10608,N_6157,N_8562);
nor U10609 (N_10609,N_7598,N_6529);
nand U10610 (N_10610,N_6420,N_8210);
nor U10611 (N_10611,N_6971,N_7637);
nand U10612 (N_10612,N_6097,N_5217);
nor U10613 (N_10613,N_8310,N_6162);
nand U10614 (N_10614,N_6371,N_8200);
nand U10615 (N_10615,N_8687,N_6898);
nand U10616 (N_10616,N_9583,N_6995);
nand U10617 (N_10617,N_9998,N_9750);
or U10618 (N_10618,N_9019,N_9516);
xor U10619 (N_10619,N_7231,N_6334);
or U10620 (N_10620,N_8748,N_8465);
nor U10621 (N_10621,N_9342,N_8574);
and U10622 (N_10622,N_5300,N_8085);
xor U10623 (N_10623,N_8331,N_7636);
nor U10624 (N_10624,N_7187,N_8019);
xnor U10625 (N_10625,N_6017,N_7330);
and U10626 (N_10626,N_9500,N_5442);
and U10627 (N_10627,N_8499,N_6379);
and U10628 (N_10628,N_8457,N_5200);
and U10629 (N_10629,N_9001,N_8236);
or U10630 (N_10630,N_6803,N_5140);
or U10631 (N_10631,N_5057,N_8293);
or U10632 (N_10632,N_7405,N_9694);
and U10633 (N_10633,N_9179,N_5070);
xnor U10634 (N_10634,N_5474,N_7975);
and U10635 (N_10635,N_8161,N_8414);
and U10636 (N_10636,N_6036,N_7764);
or U10637 (N_10637,N_6055,N_9551);
nor U10638 (N_10638,N_6365,N_9163);
or U10639 (N_10639,N_5348,N_9835);
xor U10640 (N_10640,N_5278,N_5261);
xor U10641 (N_10641,N_8238,N_6984);
and U10642 (N_10642,N_8779,N_7502);
xnor U10643 (N_10643,N_6660,N_6832);
nand U10644 (N_10644,N_7948,N_5971);
and U10645 (N_10645,N_6293,N_9288);
nor U10646 (N_10646,N_7535,N_5299);
nor U10647 (N_10647,N_5085,N_7792);
or U10648 (N_10648,N_5871,N_5919);
and U10649 (N_10649,N_7438,N_8688);
nand U10650 (N_10650,N_5449,N_8812);
xor U10651 (N_10651,N_8973,N_6200);
or U10652 (N_10652,N_7264,N_8967);
or U10653 (N_10653,N_9806,N_6696);
nor U10654 (N_10654,N_7371,N_5244);
and U10655 (N_10655,N_9223,N_6400);
nor U10656 (N_10656,N_7178,N_5715);
and U10657 (N_10657,N_9790,N_7448);
or U10658 (N_10658,N_6690,N_6830);
and U10659 (N_10659,N_6723,N_7524);
and U10660 (N_10660,N_5683,N_7740);
nor U10661 (N_10661,N_5364,N_6878);
and U10662 (N_10662,N_9053,N_5150);
and U10663 (N_10663,N_6311,N_6666);
nand U10664 (N_10664,N_7702,N_9222);
and U10665 (N_10665,N_8594,N_6908);
xnor U10666 (N_10666,N_9137,N_6471);
nand U10667 (N_10667,N_6424,N_5055);
nor U10668 (N_10668,N_9023,N_5920);
and U10669 (N_10669,N_9192,N_9765);
xnor U10670 (N_10670,N_7828,N_9081);
nor U10671 (N_10671,N_8782,N_6135);
nor U10672 (N_10672,N_5384,N_8302);
nand U10673 (N_10673,N_6553,N_5378);
and U10674 (N_10674,N_8165,N_6291);
nand U10675 (N_10675,N_6252,N_6174);
or U10676 (N_10676,N_9294,N_9727);
or U10677 (N_10677,N_6662,N_6194);
or U10678 (N_10678,N_6136,N_9465);
nor U10679 (N_10679,N_8648,N_6750);
or U10680 (N_10680,N_8402,N_6419);
nor U10681 (N_10681,N_8193,N_8863);
and U10682 (N_10682,N_9592,N_9459);
or U10683 (N_10683,N_8612,N_9818);
or U10684 (N_10684,N_8259,N_8260);
or U10685 (N_10685,N_7400,N_9660);
and U10686 (N_10686,N_8209,N_8607);
and U10687 (N_10687,N_9515,N_8286);
nand U10688 (N_10688,N_5311,N_9535);
and U10689 (N_10689,N_7105,N_9204);
and U10690 (N_10690,N_5705,N_7182);
or U10691 (N_10691,N_5990,N_8032);
xnor U10692 (N_10692,N_6742,N_8435);
and U10693 (N_10693,N_5755,N_5735);
and U10694 (N_10694,N_6729,N_5465);
nor U10695 (N_10695,N_8589,N_5427);
or U10696 (N_10696,N_7200,N_9190);
nand U10697 (N_10697,N_8553,N_7677);
xnor U10698 (N_10698,N_6496,N_5521);
or U10699 (N_10699,N_7139,N_6235);
and U10700 (N_10700,N_9951,N_5119);
or U10701 (N_10701,N_5565,N_6873);
nand U10702 (N_10702,N_9505,N_8030);
nor U10703 (N_10703,N_6998,N_9327);
nand U10704 (N_10704,N_5349,N_6340);
nand U10705 (N_10705,N_7107,N_8307);
nand U10706 (N_10706,N_7212,N_9708);
and U10707 (N_10707,N_5533,N_8773);
nand U10708 (N_10708,N_9925,N_7093);
nor U10709 (N_10709,N_6833,N_8322);
or U10710 (N_10710,N_7986,N_7475);
or U10711 (N_10711,N_8160,N_9755);
nor U10712 (N_10712,N_9716,N_7414);
and U10713 (N_10713,N_7591,N_6469);
and U10714 (N_10714,N_8815,N_6594);
and U10715 (N_10715,N_8737,N_8449);
or U10716 (N_10716,N_8530,N_6178);
and U10717 (N_10717,N_6147,N_5297);
xnor U10718 (N_10718,N_8131,N_7327);
nand U10719 (N_10719,N_6150,N_9453);
nor U10720 (N_10720,N_8997,N_5593);
nand U10721 (N_10721,N_6516,N_7649);
nand U10722 (N_10722,N_8634,N_7939);
nand U10723 (N_10723,N_5174,N_9833);
nor U10724 (N_10724,N_6771,N_9975);
and U10725 (N_10725,N_8549,N_8849);
and U10726 (N_10726,N_9247,N_5028);
nand U10727 (N_10727,N_7185,N_6020);
nor U10728 (N_10728,N_8944,N_7078);
nor U10729 (N_10729,N_6470,N_8386);
and U10730 (N_10730,N_9231,N_9103);
nor U10731 (N_10731,N_7156,N_7451);
nor U10732 (N_10732,N_6468,N_6396);
or U10733 (N_10733,N_6778,N_9980);
nor U10734 (N_10734,N_8468,N_5024);
nor U10735 (N_10735,N_8803,N_6275);
or U10736 (N_10736,N_6042,N_9141);
nand U10737 (N_10737,N_7539,N_8347);
nand U10738 (N_10738,N_8343,N_9220);
or U10739 (N_10739,N_6706,N_7455);
or U10740 (N_10740,N_7336,N_9632);
or U10741 (N_10741,N_7388,N_9862);
nand U10742 (N_10742,N_8218,N_7958);
xor U10743 (N_10743,N_6495,N_9295);
nand U10744 (N_10744,N_9712,N_7224);
or U10745 (N_10745,N_6355,N_7549);
or U10746 (N_10746,N_7120,N_7247);
nor U10747 (N_10747,N_7938,N_9972);
xor U10748 (N_10748,N_7220,N_7326);
and U10749 (N_10749,N_7972,N_9606);
and U10750 (N_10750,N_7170,N_7392);
nand U10751 (N_10751,N_7731,N_8883);
xnor U10752 (N_10752,N_8832,N_6195);
and U10753 (N_10753,N_6046,N_5350);
and U10754 (N_10754,N_9227,N_8484);
and U10755 (N_10755,N_5210,N_9739);
and U10756 (N_10756,N_5636,N_5725);
nand U10757 (N_10757,N_9030,N_8049);
nor U10758 (N_10758,N_5009,N_7487);
nand U10759 (N_10759,N_9704,N_7492);
nand U10760 (N_10760,N_6472,N_7389);
xnor U10761 (N_10761,N_7974,N_8408);
nor U10762 (N_10762,N_7710,N_9312);
or U10763 (N_10763,N_7630,N_6177);
or U10764 (N_10764,N_7398,N_6452);
or U10765 (N_10765,N_6015,N_9683);
xor U10766 (N_10766,N_8233,N_9792);
nand U10767 (N_10767,N_9724,N_8695);
nor U10768 (N_10768,N_7020,N_9663);
nand U10769 (N_10769,N_6449,N_5520);
nor U10770 (N_10770,N_9152,N_6591);
nand U10771 (N_10771,N_9586,N_9743);
xor U10772 (N_10772,N_6341,N_9529);
and U10773 (N_10773,N_6645,N_8318);
nor U10774 (N_10774,N_9782,N_7684);
and U10775 (N_10775,N_7929,N_8547);
nor U10776 (N_10776,N_7469,N_7697);
xnor U10777 (N_10777,N_8226,N_8690);
and U10778 (N_10778,N_9687,N_7119);
nand U10779 (N_10779,N_7599,N_7402);
nor U10780 (N_10780,N_6446,N_7930);
and U10781 (N_10781,N_7013,N_8003);
nand U10782 (N_10782,N_9919,N_7337);
or U10783 (N_10783,N_6839,N_5352);
nand U10784 (N_10784,N_6008,N_9198);
and U10785 (N_10785,N_6316,N_6393);
or U10786 (N_10786,N_6667,N_5600);
nor U10787 (N_10787,N_9307,N_9067);
or U10788 (N_10788,N_6066,N_5191);
or U10789 (N_10789,N_8718,N_9427);
and U10790 (N_10790,N_8482,N_9783);
or U10791 (N_10791,N_6615,N_9920);
or U10792 (N_10792,N_8145,N_7647);
and U10793 (N_10793,N_6234,N_9484);
nand U10794 (N_10794,N_5911,N_6314);
nor U10795 (N_10795,N_8904,N_9940);
and U10796 (N_10796,N_9328,N_8298);
xnor U10797 (N_10797,N_6230,N_7106);
xnor U10798 (N_10798,N_6392,N_9565);
nand U10799 (N_10799,N_5887,N_6319);
and U10800 (N_10800,N_9489,N_8455);
nand U10801 (N_10801,N_6688,N_6642);
or U10802 (N_10802,N_8592,N_7994);
xnor U10803 (N_10803,N_7239,N_5828);
and U10804 (N_10804,N_9153,N_6240);
or U10805 (N_10805,N_8966,N_8714);
nor U10806 (N_10806,N_6352,N_9229);
and U10807 (N_10807,N_9614,N_6116);
nor U10808 (N_10808,N_6381,N_6364);
and U10809 (N_10809,N_6743,N_7768);
or U10810 (N_10810,N_6677,N_7117);
nand U10811 (N_10811,N_9992,N_8235);
and U10812 (N_10812,N_6628,N_6583);
nor U10813 (N_10813,N_8140,N_9208);
or U10814 (N_10814,N_7081,N_7470);
xor U10815 (N_10815,N_6507,N_5518);
xnor U10816 (N_10816,N_8365,N_6909);
or U10817 (N_10817,N_6336,N_7669);
nor U10818 (N_10818,N_6653,N_8229);
nand U10819 (N_10819,N_7314,N_8420);
and U10820 (N_10820,N_9702,N_5419);
nor U10821 (N_10821,N_8120,N_8640);
nor U10822 (N_10822,N_6614,N_9435);
and U10823 (N_10823,N_7076,N_5234);
and U10824 (N_10824,N_5840,N_9382);
nand U10825 (N_10825,N_9622,N_5343);
nor U10826 (N_10826,N_5123,N_7568);
nand U10827 (N_10827,N_5007,N_9507);
or U10828 (N_10828,N_5144,N_9539);
xor U10829 (N_10829,N_7806,N_9945);
and U10830 (N_10830,N_8345,N_9701);
nand U10831 (N_10831,N_9394,N_6301);
or U10832 (N_10832,N_6513,N_6134);
or U10833 (N_10833,N_8959,N_8791);
and U10834 (N_10834,N_6802,N_5888);
nor U10835 (N_10835,N_8142,N_7209);
or U10836 (N_10836,N_5372,N_8146);
or U10837 (N_10837,N_5959,N_5882);
and U10838 (N_10838,N_8861,N_6655);
or U10839 (N_10839,N_7563,N_5193);
nand U10840 (N_10840,N_5270,N_6598);
and U10841 (N_10841,N_9084,N_9314);
nor U10842 (N_10842,N_6665,N_7960);
xor U10843 (N_10843,N_7126,N_9824);
nor U10844 (N_10844,N_5979,N_5587);
nand U10845 (N_10845,N_6812,N_5731);
nand U10846 (N_10846,N_5691,N_6825);
nand U10847 (N_10847,N_9914,N_8056);
nor U10848 (N_10848,N_8725,N_5015);
nor U10849 (N_10849,N_6153,N_5134);
nand U10850 (N_10850,N_9402,N_6893);
xor U10851 (N_10851,N_6877,N_9567);
or U10852 (N_10852,N_9444,N_5485);
and U10853 (N_10853,N_5941,N_8675);
and U10854 (N_10854,N_7654,N_6575);
nor U10855 (N_10855,N_7907,N_8321);
nand U10856 (N_10856,N_5267,N_8987);
nand U10857 (N_10857,N_7063,N_5685);
and U10858 (N_10858,N_5281,N_8709);
nand U10859 (N_10859,N_8497,N_7782);
nand U10860 (N_10860,N_7433,N_6659);
nand U10861 (N_10861,N_8072,N_9196);
nand U10862 (N_10862,N_5051,N_9946);
xnor U10863 (N_10863,N_7808,N_8389);
nand U10864 (N_10864,N_5522,N_5214);
nor U10865 (N_10865,N_9990,N_8319);
or U10866 (N_10866,N_7350,N_6375);
nor U10867 (N_10867,N_7082,N_9513);
nand U10868 (N_10868,N_8760,N_8366);
nor U10869 (N_10869,N_5686,N_6681);
nor U10870 (N_10870,N_6692,N_9876);
or U10871 (N_10871,N_7843,N_6043);
nor U10872 (N_10872,N_5388,N_8102);
or U10873 (N_10873,N_7959,N_5257);
nand U10874 (N_10874,N_7207,N_9883);
nor U10875 (N_10875,N_9330,N_9849);
or U10876 (N_10876,N_9028,N_7460);
nand U10877 (N_10877,N_7363,N_8325);
or U10878 (N_10878,N_5328,N_9728);
or U10879 (N_10879,N_7461,N_7309);
xnor U10880 (N_10880,N_6238,N_5481);
or U10881 (N_10881,N_9006,N_8736);
and U10882 (N_10882,N_5989,N_6543);
nand U10883 (N_10883,N_6656,N_9042);
xor U10884 (N_10884,N_9336,N_8024);
and U10885 (N_10885,N_6652,N_7597);
nand U10886 (N_10886,N_8920,N_6300);
nand U10887 (N_10887,N_8132,N_9934);
or U10888 (N_10888,N_6239,N_5396);
nand U10889 (N_10889,N_9401,N_9568);
nor U10890 (N_10890,N_9154,N_6005);
nand U10891 (N_10891,N_8099,N_8416);
xor U10892 (N_10892,N_6431,N_9044);
nand U10893 (N_10893,N_6946,N_9763);
and U10894 (N_10894,N_8897,N_8273);
xor U10895 (N_10895,N_7166,N_7822);
nand U10896 (N_10896,N_8135,N_7545);
nand U10897 (N_10897,N_9655,N_5641);
xnor U10898 (N_10898,N_7270,N_9071);
nand U10899 (N_10899,N_5401,N_9537);
nor U10900 (N_10900,N_8917,N_8935);
and U10901 (N_10901,N_5614,N_7033);
nor U10902 (N_10902,N_7957,N_7045);
and U10903 (N_10903,N_7625,N_8717);
and U10904 (N_10904,N_5182,N_8282);
or U10905 (N_10905,N_7007,N_8933);
and U10906 (N_10906,N_8107,N_7612);
and U10907 (N_10907,N_8947,N_8296);
nor U10908 (N_10908,N_6486,N_6028);
or U10909 (N_10909,N_6620,N_5220);
nand U10910 (N_10910,N_6579,N_9458);
and U10911 (N_10911,N_9206,N_5030);
or U10912 (N_10912,N_9570,N_5083);
and U10913 (N_10913,N_7394,N_5360);
and U10914 (N_10914,N_8104,N_8314);
xor U10915 (N_10915,N_6527,N_6870);
and U10916 (N_10916,N_9358,N_9916);
xor U10917 (N_10917,N_8630,N_5764);
nand U10918 (N_10918,N_7706,N_8387);
nor U10919 (N_10919,N_5650,N_9054);
xor U10920 (N_10920,N_5993,N_6782);
nand U10921 (N_10921,N_7369,N_5559);
or U10922 (N_10922,N_7364,N_8508);
nor U10923 (N_10923,N_7700,N_9734);
and U10924 (N_10924,N_5620,N_7634);
nor U10925 (N_10925,N_5569,N_8061);
nand U10926 (N_10926,N_8186,N_9486);
and U10927 (N_10927,N_6650,N_8221);
nand U10928 (N_10928,N_7057,N_5453);
or U10929 (N_10929,N_8879,N_5168);
nor U10930 (N_10930,N_8641,N_6937);
nand U10931 (N_10931,N_7279,N_9365);
and U10932 (N_10932,N_5052,N_9488);
and U10933 (N_10933,N_7711,N_7472);
and U10934 (N_10934,N_5455,N_6700);
xor U10935 (N_10935,N_9917,N_9090);
or U10936 (N_10936,N_5609,N_6757);
xnor U10937 (N_10937,N_7305,N_5206);
nor U10938 (N_10938,N_9303,N_5324);
nand U10939 (N_10939,N_5394,N_7036);
or U10940 (N_10940,N_6263,N_9012);
nand U10941 (N_10941,N_5205,N_6586);
or U10942 (N_10942,N_6064,N_9610);
nand U10943 (N_10943,N_7985,N_8144);
or U10944 (N_10944,N_8125,N_6831);
and U10945 (N_10945,N_6824,N_6203);
and U10946 (N_10946,N_8826,N_5841);
or U10947 (N_10947,N_5466,N_8624);
nor U10948 (N_10948,N_7024,N_6190);
or U10949 (N_10949,N_9166,N_8902);
or U10950 (N_10950,N_5032,N_6450);
nand U10951 (N_10951,N_7094,N_7912);
nand U10952 (N_10952,N_9943,N_7891);
or U10953 (N_10953,N_7728,N_6120);
or U10954 (N_10954,N_7195,N_9317);
nor U10955 (N_10955,N_5033,N_5404);
xnor U10956 (N_10956,N_7359,N_7430);
nand U10957 (N_10957,N_6821,N_6458);
xor U10958 (N_10958,N_9283,N_7233);
and U10959 (N_10959,N_9027,N_6746);
nor U10960 (N_10960,N_6101,N_6872);
and U10961 (N_10961,N_5483,N_5472);
or U10962 (N_10962,N_7916,N_9131);
nor U10963 (N_10963,N_6479,N_7709);
and U10964 (N_10964,N_6254,N_8733);
nand U10965 (N_10965,N_9117,N_8040);
and U10966 (N_10966,N_6661,N_9830);
nor U10967 (N_10967,N_9939,N_7131);
nand U10968 (N_10968,N_5674,N_9648);
nand U10969 (N_10969,N_9383,N_9631);
nand U10970 (N_10970,N_5940,N_8035);
nand U10971 (N_10971,N_5251,N_8154);
nor U10972 (N_10972,N_7847,N_9550);
or U10973 (N_10973,N_8189,N_9379);
nor U10974 (N_10974,N_5684,N_7595);
nor U10975 (N_10975,N_7589,N_7908);
nor U10976 (N_10976,N_6347,N_6533);
xnor U10977 (N_10977,N_9905,N_6730);
xor U10978 (N_10978,N_6932,N_8057);
xnor U10979 (N_10979,N_9533,N_7730);
nand U10980 (N_10980,N_6350,N_6464);
nor U10981 (N_10981,N_9475,N_6047);
and U10982 (N_10982,N_6444,N_5815);
and U10983 (N_10983,N_9194,N_5425);
xnor U10984 (N_10984,N_6903,N_6390);
nor U10985 (N_10985,N_5929,N_7047);
nor U10986 (N_10986,N_9251,N_6372);
nand U10987 (N_10987,N_8242,N_6532);
or U10988 (N_10988,N_6711,N_7017);
or U10989 (N_10989,N_6574,N_5597);
nand U10990 (N_10990,N_6370,N_9647);
and U10991 (N_10991,N_9320,N_7290);
and U10992 (N_10992,N_7163,N_9184);
nor U10993 (N_10993,N_7260,N_5331);
xnor U10994 (N_10994,N_8279,N_8595);
nor U10995 (N_10995,N_7579,N_7375);
or U10996 (N_10996,N_5293,N_8775);
nor U10997 (N_10997,N_5703,N_7456);
and U10998 (N_10998,N_9148,N_5194);
and U10999 (N_10999,N_7787,N_9456);
and U11000 (N_11000,N_5779,N_8644);
nand U11001 (N_11001,N_8602,N_8071);
xor U11002 (N_11002,N_9124,N_5128);
and U11003 (N_11003,N_5303,N_8937);
and U11004 (N_11004,N_9259,N_5819);
nand U11005 (N_11005,N_6109,N_6753);
and U11006 (N_11006,N_5716,N_5582);
nand U11007 (N_11007,N_9024,N_7370);
nor U11008 (N_11008,N_9381,N_7572);
and U11009 (N_11009,N_7838,N_7165);
nand U11010 (N_11010,N_5365,N_8694);
or U11011 (N_11011,N_6888,N_7411);
and U11012 (N_11012,N_9544,N_5356);
or U11013 (N_11013,N_8738,N_7583);
nand U11014 (N_11014,N_5493,N_5501);
nor U11015 (N_11015,N_6698,N_7434);
or U11016 (N_11016,N_9600,N_7796);
nor U11017 (N_11017,N_5122,N_9658);
nand U11018 (N_11018,N_5924,N_8206);
nor U11019 (N_11019,N_7877,N_9938);
or U11020 (N_11020,N_6975,N_5942);
nand U11021 (N_11021,N_8409,N_9560);
and U11022 (N_11022,N_5477,N_5209);
and U11023 (N_11023,N_7590,N_7420);
nor U11024 (N_11024,N_6841,N_8875);
xnor U11025 (N_11025,N_8632,N_7067);
and U11026 (N_11026,N_5000,N_6192);
and U11027 (N_11027,N_7214,N_6299);
xor U11028 (N_11028,N_7009,N_8833);
xnor U11029 (N_11029,N_9187,N_9274);
and U11030 (N_11030,N_8106,N_7501);
and U11031 (N_11031,N_5950,N_8663);
nor U11032 (N_11032,N_9431,N_9255);
xor U11033 (N_11033,N_8919,N_8176);
xor U11034 (N_11034,N_7814,N_8428);
or U11035 (N_11035,N_5165,N_9466);
and U11036 (N_11036,N_9641,N_7452);
nand U11037 (N_11037,N_9087,N_7162);
or U11038 (N_11038,N_8523,N_7771);
and U11039 (N_11039,N_5822,N_6208);
nand U11040 (N_11040,N_5488,N_6443);
nor U11041 (N_11041,N_6146,N_5794);
or U11042 (N_11042,N_5824,N_6249);
or U11043 (N_11043,N_6410,N_8337);
and U11044 (N_11044,N_7914,N_7377);
and U11045 (N_11045,N_7408,N_7516);
nand U11046 (N_11046,N_6076,N_6494);
nor U11047 (N_11047,N_5130,N_8957);
nand U11048 (N_11048,N_9627,N_6302);
nand U11049 (N_11049,N_8224,N_8393);
and U11050 (N_11050,N_8441,N_8887);
and U11051 (N_11051,N_9289,N_9010);
nor U11052 (N_11052,N_7620,N_5413);
or U11053 (N_11053,N_7436,N_8223);
or U11054 (N_11054,N_6061,N_8858);
and U11055 (N_11055,N_5560,N_8667);
or U11056 (N_11056,N_5373,N_8155);
or U11057 (N_11057,N_9086,N_7735);
or U11058 (N_11058,N_9360,N_5001);
and U11059 (N_11059,N_7188,N_6813);
nor U11060 (N_11060,N_7171,N_8272);
and U11061 (N_11061,N_5713,N_5893);
nand U11062 (N_11062,N_9915,N_8068);
or U11063 (N_11063,N_8654,N_8164);
nor U11064 (N_11064,N_9601,N_9017);
nor U11065 (N_11065,N_7409,N_9002);
and U11066 (N_11066,N_9699,N_6108);
nand U11067 (N_11067,N_7982,N_7084);
nand U11068 (N_11068,N_7333,N_9182);
nor U11069 (N_11069,N_5060,N_5256);
nand U11070 (N_11070,N_6259,N_9470);
and U11071 (N_11071,N_8039,N_7226);
nand U11072 (N_11072,N_6599,N_7831);
or U11073 (N_11073,N_6562,N_7221);
or U11074 (N_11074,N_6408,N_7875);
xnor U11075 (N_11075,N_5259,N_7611);
or U11076 (N_11076,N_6021,N_9893);
and U11077 (N_11077,N_8627,N_5272);
nand U11078 (N_11078,N_8621,N_9898);
or U11079 (N_11079,N_5637,N_5856);
or U11080 (N_11080,N_9688,N_8528);
or U11081 (N_11081,N_9493,N_5189);
and U11082 (N_11082,N_7031,N_8522);
and U11083 (N_11083,N_9953,N_5049);
or U11084 (N_11084,N_9766,N_9363);
xor U11085 (N_11085,N_9172,N_5754);
nor U11086 (N_11086,N_6333,N_8584);
nor U11087 (N_11087,N_7525,N_9639);
nand U11088 (N_11088,N_8986,N_8510);
or U11089 (N_11089,N_7754,N_7307);
xnor U11090 (N_11090,N_8678,N_7190);
nand U11091 (N_11091,N_7871,N_8601);
and U11092 (N_11092,N_5116,N_7467);
nor U11093 (N_11093,N_9668,N_8943);
nand U11094 (N_11094,N_8906,N_7429);
nor U11095 (N_11095,N_8063,N_6610);
xor U11096 (N_11096,N_8797,N_6875);
nor U11097 (N_11097,N_7222,N_6274);
nand U11098 (N_11098,N_8525,N_8839);
and U11099 (N_11099,N_6461,N_7263);
nand U11100 (N_11100,N_6016,N_7819);
or U11101 (N_11101,N_7189,N_5692);
or U11102 (N_11102,N_5675,N_9216);
nand U11103 (N_11103,N_5242,N_8963);
or U11104 (N_11104,N_5280,N_5750);
nor U11105 (N_11105,N_6376,N_8041);
nand U11106 (N_11106,N_8819,N_6767);
nor U11107 (N_11107,N_8822,N_8058);
nor U11108 (N_11108,N_7227,N_8537);
or U11109 (N_11109,N_5589,N_6080);
xnor U11110 (N_11110,N_9771,N_5063);
and U11111 (N_11111,N_5215,N_6382);
xor U11112 (N_11112,N_9904,N_8679);
and U11113 (N_11113,N_8965,N_5839);
or U11114 (N_11114,N_7048,N_5041);
and U11115 (N_11115,N_6083,N_6477);
nor U11116 (N_11116,N_8228,N_8940);
xnor U11117 (N_11117,N_7751,N_5039);
or U11118 (N_11118,N_8489,N_6773);
nor U11119 (N_11119,N_7652,N_7360);
and U11120 (N_11120,N_6619,N_7011);
nor U11121 (N_11121,N_5263,N_9306);
or U11122 (N_11122,N_7927,N_9490);
or U11123 (N_11123,N_9809,N_8278);
xnor U11124 (N_11124,N_5823,N_9827);
or U11125 (N_11125,N_9371,N_5207);
xor U11126 (N_11126,N_5985,N_9896);
nand U11127 (N_11127,N_8156,N_7721);
nor U11128 (N_11128,N_6626,N_6149);
and U11129 (N_11129,N_8800,N_7727);
and U11130 (N_11130,N_8227,N_9947);
and U11131 (N_11131,N_6474,N_8394);
nand U11132 (N_11132,N_7406,N_8413);
nand U11133 (N_11133,N_5818,N_8327);
nand U11134 (N_11134,N_8124,N_7141);
xnor U11135 (N_11135,N_7992,N_9158);
or U11136 (N_11136,N_9313,N_9136);
and U11137 (N_11137,N_7718,N_7541);
nor U11138 (N_11138,N_7096,N_8262);
nand U11139 (N_11139,N_9962,N_6713);
nor U11140 (N_11140,N_5532,N_6012);
or U11141 (N_11141,N_6442,N_9731);
nor U11142 (N_11142,N_6960,N_7996);
or U11143 (N_11143,N_8533,N_6205);
or U11144 (N_11144,N_8505,N_9999);
or U11145 (N_11145,N_7678,N_9703);
and U11146 (N_11146,N_8459,N_6457);
nor U11147 (N_11147,N_9298,N_5058);
and U11148 (N_11148,N_7147,N_6728);
nand U11149 (N_11149,N_8551,N_9476);
nand U11150 (N_11150,N_5456,N_9749);
nand U11151 (N_11151,N_6985,N_5266);
or U11152 (N_11152,N_9209,N_6256);
or U11153 (N_11153,N_9225,N_5741);
nor U11154 (N_11154,N_9050,N_6220);
nor U11155 (N_11155,N_8799,N_6747);
and U11156 (N_11156,N_5486,N_5448);
xor U11157 (N_11157,N_5109,N_5577);
and U11158 (N_11158,N_7466,N_6427);
nand U11159 (N_11159,N_6176,N_5081);
nand U11160 (N_11160,N_6670,N_8101);
nor U11161 (N_11161,N_9850,N_6260);
and U11162 (N_11162,N_8728,N_9063);
or U11163 (N_11163,N_9853,N_8100);
and U11164 (N_11164,N_7181,N_5811);
nor U11165 (N_11165,N_5345,N_7397);
and U11166 (N_11166,N_8658,N_5265);
nand U11167 (N_11167,N_5837,N_9523);
nand U11168 (N_11168,N_5951,N_5291);
nand U11169 (N_11169,N_5277,N_6010);
nor U11170 (N_11170,N_6473,N_5879);
or U11171 (N_11171,N_5645,N_6856);
or U11172 (N_11172,N_5424,N_7331);
nor U11173 (N_11173,N_5581,N_6838);
xnor U11174 (N_11174,N_8339,N_9628);
and U11175 (N_11175,N_6092,N_7234);
and U11176 (N_11176,N_9950,N_5268);
or U11177 (N_11177,N_8188,N_6567);
and U11178 (N_11178,N_5496,N_8418);
nand U11179 (N_11179,N_9878,N_8804);
nand U11180 (N_11180,N_8496,N_8568);
nand U11181 (N_11181,N_9275,N_5874);
and U11182 (N_11182,N_5141,N_7717);
nor U11183 (N_11183,N_7255,N_8629);
xnor U11184 (N_11184,N_6978,N_8406);
nor U11185 (N_11185,N_9617,N_9760);
nand U11186 (N_11186,N_6836,N_7352);
nand U11187 (N_11187,N_6126,N_8814);
nand U11188 (N_11188,N_6031,N_9455);
nor U11189 (N_11189,N_8817,N_9880);
or U11190 (N_11190,N_9083,N_6639);
nand U11191 (N_11191,N_7744,N_5333);
or U11192 (N_11192,N_5974,N_7641);
nand U11193 (N_11193,N_6363,N_9468);
nand U11194 (N_11194,N_5087,N_5127);
and U11195 (N_11195,N_9624,N_5375);
xnor U11196 (N_11196,N_8864,N_5092);
nor U11197 (N_11197,N_5160,N_5928);
and U11198 (N_11198,N_5734,N_9104);
nor U11199 (N_11199,N_5875,N_8456);
nand U11200 (N_11200,N_6448,N_7528);
xor U11201 (N_11201,N_5310,N_7773);
and U11202 (N_11202,N_7130,N_7816);
nand U11203 (N_11203,N_6322,N_7259);
or U11204 (N_11204,N_8419,N_9804);
nand U11205 (N_11205,N_5552,N_7387);
or U11206 (N_11206,N_7698,N_8682);
xnor U11207 (N_11207,N_6540,N_7879);
nand U11208 (N_11208,N_5420,N_5079);
nor U11209 (N_11209,N_7919,N_9887);
nor U11210 (N_11210,N_6815,N_8932);
nor U11211 (N_11211,N_5657,N_8853);
and U11212 (N_11212,N_8927,N_6191);
xor U11213 (N_11213,N_8757,N_8948);
and U11214 (N_11214,N_8076,N_8751);
nand U11215 (N_11215,N_6439,N_7230);
or U11216 (N_11216,N_7809,N_6369);
or U11217 (N_11217,N_6219,N_5446);
or U11218 (N_11218,N_5395,N_7892);
and U11219 (N_11219,N_7289,N_7180);
and U11220 (N_11220,N_9979,N_9942);
nand U11221 (N_11221,N_9380,N_9326);
nand U11222 (N_11222,N_9346,N_5680);
nor U11223 (N_11223,N_5789,N_7532);
and U11224 (N_11224,N_8222,N_6791);
nor U11225 (N_11225,N_6499,N_5800);
or U11226 (N_11226,N_6973,N_9816);
nor U11227 (N_11227,N_9269,N_9308);
nand U11228 (N_11228,N_8953,N_8026);
nor U11229 (N_11229,N_9690,N_9637);
and U11230 (N_11230,N_8544,N_5539);
or U11231 (N_11231,N_7494,N_5809);
nor U11232 (N_11232,N_9420,N_5102);
or U11233 (N_11233,N_9125,N_7750);
and U11234 (N_11234,N_7695,N_7042);
nand U11235 (N_11235,N_8114,N_8349);
or U11236 (N_11236,N_7857,N_5870);
and U11237 (N_11237,N_7942,N_6498);
xnor U11238 (N_11238,N_6478,N_8133);
or U11239 (N_11239,N_6436,N_9897);
and U11240 (N_11240,N_5608,N_8494);
and U11241 (N_11241,N_9669,N_6912);
and U11242 (N_11242,N_7010,N_5902);
nor U11243 (N_11243,N_6772,N_8978);
nor U11244 (N_11244,N_8092,N_7484);
xor U11245 (N_11245,N_9316,N_9237);
nand U11246 (N_11246,N_8855,N_9436);
xnor U11247 (N_11247,N_9536,N_5619);
nor U11248 (N_11248,N_7946,N_8925);
nor U11249 (N_11249,N_8000,N_8726);
nand U11250 (N_11250,N_6482,N_5064);
and U11251 (N_11251,N_9956,N_7140);
nor U11252 (N_11252,N_6056,N_6415);
and U11253 (N_11253,N_6701,N_9143);
or U11254 (N_11254,N_7444,N_9290);
or U11255 (N_11255,N_7855,N_9088);
and U11256 (N_11256,N_7976,N_8976);
and U11257 (N_11257,N_9344,N_9171);
nand U11258 (N_11258,N_5768,N_6763);
and U11259 (N_11259,N_7146,N_5494);
nand U11260 (N_11260,N_7215,N_7116);
and U11261 (N_11261,N_6198,N_8824);
nand U11262 (N_11262,N_9870,N_8043);
nand U11263 (N_11263,N_8798,N_6011);
xor U11264 (N_11264,N_7679,N_9509);
or U11265 (N_11265,N_5491,N_5752);
nand U11266 (N_11266,N_8025,N_8074);
nor U11267 (N_11267,N_9517,N_9675);
or U11268 (N_11268,N_7566,N_7547);
and U11269 (N_11269,N_6265,N_6051);
or U11270 (N_11270,N_9469,N_5129);
xnor U11271 (N_11271,N_7800,N_6546);
xnor U11272 (N_11272,N_7246,N_7519);
and U11273 (N_11273,N_8635,N_5603);
nand U11274 (N_11274,N_6114,N_5240);
or U11275 (N_11275,N_7781,N_6267);
nand U11276 (N_11276,N_8598,N_6970);
nand U11277 (N_11277,N_9009,N_7866);
nor U11278 (N_11278,N_7884,N_9831);
nor U11279 (N_11279,N_9315,N_8184);
and U11280 (N_11280,N_7493,N_6475);
and U11281 (N_11281,N_6602,N_9238);
or U11282 (N_11282,N_9108,N_9861);
and U11283 (N_11283,N_5099,N_5309);
or U11284 (N_11284,N_7749,N_5813);
or U11285 (N_11285,N_6680,N_7906);
or U11286 (N_11286,N_7691,N_6531);
nor U11287 (N_11287,N_5137,N_7761);
nand U11288 (N_11288,N_5812,N_9046);
nand U11289 (N_11289,N_9773,N_7440);
nor U11290 (N_11290,N_7944,N_8876);
nand U11291 (N_11291,N_5666,N_9891);
or U11292 (N_11292,N_6353,N_9477);
or U11293 (N_11293,N_6435,N_7593);
nor U11294 (N_11294,N_9252,N_9697);
or U11295 (N_11295,N_6914,N_6327);
or U11296 (N_11296,N_9285,N_9964);
nand U11297 (N_11297,N_6566,N_7743);
nor U11298 (N_11298,N_6356,N_8178);
nor U11299 (N_11299,N_7931,N_6576);
nand U11300 (N_11300,N_6864,N_9176);
nand U11301 (N_11301,N_5862,N_9863);
xnor U11302 (N_11302,N_5966,N_5390);
and U11303 (N_11303,N_8838,N_7551);
nand U11304 (N_11304,N_9844,N_7724);
xnor U11305 (N_11305,N_5693,N_8478);
nand U11306 (N_11306,N_8888,N_6755);
xnor U11307 (N_11307,N_7317,N_9473);
or U11308 (N_11308,N_8055,N_5208);
or U11309 (N_11309,N_7053,N_9941);
nor U11310 (N_11310,N_5223,N_8891);
nand U11311 (N_11311,N_5076,N_9541);
nor U11312 (N_11312,N_7900,N_5414);
nand U11313 (N_11313,N_6052,N_5460);
and U11314 (N_11314,N_6933,N_7550);
nor U11315 (N_11315,N_8950,N_6207);
or U11316 (N_11316,N_5918,N_5791);
nand U11317 (N_11317,N_9527,N_6607);
nor U11318 (N_11318,N_6865,N_5556);
or U11319 (N_11319,N_6523,N_5170);
nand U11320 (N_11320,N_5308,N_7995);
nand U11321 (N_11321,N_5183,N_8583);
nand U11322 (N_11322,N_6285,N_8596);
and U11323 (N_11323,N_7065,N_9599);
or U11324 (N_11324,N_7883,N_8284);
nor U11325 (N_11325,N_5984,N_8587);
nor U11326 (N_11326,N_8128,N_5571);
or U11327 (N_11327,N_6094,N_6613);
or U11328 (N_11328,N_6437,N_7240);
nand U11329 (N_11329,N_8375,N_7419);
or U11330 (N_11330,N_7250,N_8354);
nand U11331 (N_11331,N_7971,N_7399);
nor U11332 (N_11332,N_5086,N_8346);
and U11333 (N_11333,N_9922,N_5672);
and U11334 (N_11334,N_5932,N_6954);
xnor U11335 (N_11335,N_9902,N_7575);
and U11336 (N_11336,N_5298,N_8784);
nand U11337 (N_11337,N_8724,N_8539);
nand U11338 (N_11338,N_9219,N_6887);
nand U11339 (N_11339,N_8922,N_6565);
nand U11340 (N_11340,N_9230,N_5817);
xor U11341 (N_11341,N_6899,N_9546);
or U11342 (N_11342,N_7368,N_8719);
or U11343 (N_11343,N_8529,N_9846);
nor U11344 (N_11344,N_9908,N_5994);
nor U11345 (N_11345,N_5148,N_8777);
or U11346 (N_11346,N_8064,N_7536);
or U11347 (N_11347,N_5176,N_7054);
nor U11348 (N_11348,N_5329,N_7614);
nand U11349 (N_11349,N_8936,N_9638);
xnor U11350 (N_11350,N_6282,N_9616);
nand U11351 (N_11351,N_5135,N_8755);
or U11352 (N_11352,N_9291,N_9847);
nor U11353 (N_11353,N_7893,N_9626);
nor U11354 (N_11354,N_6213,N_5687);
nand U11355 (N_11355,N_5881,N_8181);
nand U11356 (N_11356,N_6225,N_6658);
nor U11357 (N_11357,N_5889,N_7510);
and U11358 (N_11358,N_7578,N_6339);
xor U11359 (N_11359,N_6060,N_5778);
or U11360 (N_11360,N_9978,N_8823);
and U11361 (N_11361,N_6725,N_5724);
nor U11362 (N_11362,N_6318,N_5644);
or U11363 (N_11363,N_5986,N_7840);
xnor U11364 (N_11364,N_7223,N_6044);
and U11365 (N_11365,N_9375,N_9331);
xor U11366 (N_11366,N_5164,N_8554);
nand U11367 (N_11367,N_6977,N_8503);
nor U11368 (N_11368,N_5461,N_6251);
or U11369 (N_11369,N_7441,N_8786);
or U11370 (N_11370,N_6632,N_9988);
or U11371 (N_11371,N_6896,N_9265);
nand U11372 (N_11372,N_7071,N_8159);
nor U11373 (N_11373,N_7692,N_5369);
nand U11374 (N_11374,N_6817,N_5376);
xnor U11375 (N_11375,N_7615,N_6243);
or U11376 (N_11376,N_9936,N_7269);
and U11377 (N_11377,N_9751,N_6654);
or U11378 (N_11378,N_6924,N_8123);
nor U11379 (N_11379,N_9418,N_5774);
nand U11380 (N_11380,N_7617,N_9803);
nand U11381 (N_11381,N_5020,N_6361);
or U11382 (N_11382,N_8545,N_8638);
nor U11383 (N_11383,N_9580,N_5695);
or U11384 (N_11384,N_9020,N_6004);
nor U11385 (N_11385,N_5226,N_9270);
nand U11386 (N_11386,N_7407,N_5546);
or U11387 (N_11387,N_9177,N_9618);
nand U11388 (N_11388,N_9693,N_5290);
nand U11389 (N_11389,N_8275,N_7108);
nor U11390 (N_11390,N_6928,N_9868);
or U11391 (N_11391,N_8854,N_7574);
or U11392 (N_11392,N_5100,N_6152);
xor U11393 (N_11393,N_5906,N_8173);
xnor U11394 (N_11394,N_6018,N_6890);
or U11395 (N_11395,N_7825,N_9362);
nor U11396 (N_11396,N_5855,N_7613);
nand U11397 (N_11397,N_7341,N_7038);
nand U11398 (N_11398,N_5665,N_8720);
nor U11399 (N_11399,N_5926,N_7882);
and U11400 (N_11400,N_5131,N_8871);
and U11401 (N_11401,N_5908,N_8243);
or U11402 (N_11402,N_6310,N_7913);
or U11403 (N_11403,N_8930,N_9620);
nor U11404 (N_11404,N_5498,N_8411);
nand U11405 (N_11405,N_5967,N_7449);
xor U11406 (N_11406,N_5785,N_8802);
or U11407 (N_11407,N_5017,N_8400);
and U11408 (N_11408,N_5852,N_7272);
or U11409 (N_11409,N_9495,N_8984);
nor U11410 (N_11410,N_8954,N_7447);
nand U11411 (N_11411,N_8845,N_7100);
or U11412 (N_11412,N_6806,N_7785);
and U11413 (N_11413,N_7581,N_8651);
nor U11414 (N_11414,N_5185,N_6493);
or U11415 (N_11415,N_7763,N_5698);
and U11416 (N_11416,N_6582,N_7193);
and U11417 (N_11417,N_9386,N_5471);
or U11418 (N_11418,N_6624,N_5235);
xnor U11419 (N_11419,N_9756,N_5947);
or U11420 (N_11420,N_8166,N_5012);
and U11421 (N_11421,N_5803,N_8300);
and U11422 (N_11422,N_7426,N_5934);
nor U11423 (N_11423,N_7347,N_9049);
and U11424 (N_11424,N_6631,N_5772);
nand U11425 (N_11425,N_8969,N_6885);
and U11426 (N_11426,N_7791,N_8290);
or U11427 (N_11427,N_7339,N_5526);
nand U11428 (N_11428,N_5010,N_6993);
and U11429 (N_11429,N_5827,N_5158);
or U11430 (N_11430,N_9457,N_8412);
xor U11431 (N_11431,N_6774,N_8126);
xor U11432 (N_11432,N_9705,N_5065);
nand U11433 (N_11433,N_7194,N_8460);
nor U11434 (N_11434,N_5640,N_9746);
or U11435 (N_11435,N_8806,N_5433);
or U11436 (N_11436,N_7626,N_9673);
nand U11437 (N_11437,N_6089,N_7850);
or U11438 (N_11438,N_7199,N_7004);
nor U11439 (N_11439,N_8900,N_9413);
or U11440 (N_11440,N_9051,N_8626);
nor U11441 (N_11441,N_9246,N_8983);
nor U11442 (N_11442,N_9506,N_5445);
nand U11443 (N_11443,N_5706,N_8230);
xor U11444 (N_11444,N_8110,N_6748);
nor U11445 (N_11445,N_7790,N_6151);
nor U11446 (N_11446,N_8982,N_6983);
nand U11447 (N_11447,N_7001,N_7794);
and U11448 (N_11448,N_9261,N_8005);
nor U11449 (N_11449,N_6406,N_7134);
or U11450 (N_11450,N_7424,N_8483);
or U11451 (N_11451,N_9834,N_8391);
nand U11452 (N_11452,N_7923,N_9100);
or U11453 (N_11453,N_6168,N_6422);
nor U11454 (N_11454,N_7253,N_9093);
or U11455 (N_11455,N_7112,N_9695);
nand U11456 (N_11456,N_7876,N_5201);
nand U11457 (N_11457,N_7498,N_9968);
nand U11458 (N_11458,N_9997,N_7310);
nor U11459 (N_11459,N_8616,N_6272);
or U11460 (N_11460,N_5503,N_6664);
nand U11461 (N_11461,N_7046,N_9603);
nand U11462 (N_11462,N_9522,N_8471);
xnor U11463 (N_11463,N_7739,N_8971);
nand U11464 (N_11464,N_6394,N_7061);
or U11465 (N_11465,N_7863,N_7507);
and U11466 (N_11466,N_6600,N_5459);
or U11467 (N_11467,N_7534,N_6130);
and U11468 (N_11468,N_9719,N_5949);
nand U11469 (N_11469,N_9557,N_6570);
nor U11470 (N_11470,N_5664,N_7439);
nand U11471 (N_11471,N_5763,N_7633);
nand U11472 (N_11472,N_5523,N_8604);
xnor U11473 (N_11473,N_5953,N_6222);
nor U11474 (N_11474,N_8048,N_8846);
and U11475 (N_11475,N_7103,N_7016);
nor U11476 (N_11476,N_6343,N_7160);
or U11477 (N_11477,N_8452,N_5612);
xnor U11478 (N_11478,N_8946,N_9165);
nand U11479 (N_11479,N_6647,N_5061);
nor U11480 (N_11480,N_7548,N_9441);
nand U11481 (N_11481,N_8264,N_5727);
and U11482 (N_11482,N_9888,N_9558);
nand U11483 (N_11483,N_7911,N_8677);
nor U11484 (N_11484,N_9650,N_7862);
nor U11485 (N_11485,N_8541,N_9134);
nor U11486 (N_11486,N_9127,N_8909);
and U11487 (N_11487,N_7745,N_8487);
and U11488 (N_11488,N_7232,N_5436);
nand U11489 (N_11489,N_6621,N_6787);
nand U11490 (N_11490,N_7945,N_8013);
and U11491 (N_11491,N_6019,N_6674);
or U11492 (N_11492,N_9043,N_6321);
nor U11493 (N_11493,N_7559,N_5976);
nand U11494 (N_11494,N_9256,N_9524);
and U11495 (N_11495,N_6451,N_6128);
or U11496 (N_11496,N_9388,N_7158);
or U11497 (N_11497,N_7257,N_9774);
nor U11498 (N_11498,N_7365,N_5221);
nor U11499 (N_11499,N_6580,N_6678);
nand U11500 (N_11500,N_7427,N_9722);
xor U11501 (N_11501,N_5381,N_5437);
and U11502 (N_11502,N_8835,N_8336);
nor U11503 (N_11503,N_9501,N_9073);
xnor U11504 (N_11504,N_8018,N_8844);
or U11505 (N_11505,N_6445,N_5495);
nand U11506 (N_11506,N_9353,N_9354);
xor U11507 (N_11507,N_7865,N_5869);
nor U11508 (N_11508,N_9180,N_5831);
nor U11509 (N_11509,N_5826,N_9111);
nor U11510 (N_11510,N_8081,N_8006);
xnor U11511 (N_11511,N_8882,N_7558);
nor U11512 (N_11512,N_7701,N_9232);
nand U11513 (N_11513,N_8703,N_5332);
nand U11514 (N_11514,N_7921,N_5760);
xnor U11515 (N_11515,N_6776,N_8637);
nor U11516 (N_11516,N_5098,N_8964);
and U11517 (N_11517,N_5502,N_5383);
or U11518 (N_11518,N_5212,N_6947);
or U11519 (N_11519,N_7092,N_5860);
or U11520 (N_11520,N_6629,N_7518);
nand U11521 (N_11521,N_7219,N_7812);
or U11522 (N_11522,N_8121,N_8610);
nand U11523 (N_11523,N_5387,N_5340);
nand U11524 (N_11524,N_9867,N_7963);
xnor U11525 (N_11525,N_8750,N_8573);
xnor U11526 (N_11526,N_8780,N_9957);
xor U11527 (N_11527,N_6844,N_8665);
or U11528 (N_11528,N_6273,N_8401);
or U11529 (N_11529,N_8869,N_5008);
and U11530 (N_11530,N_5468,N_6182);
nand U11531 (N_11531,N_5124,N_9762);
xor U11532 (N_11532,N_6315,N_7725);
nand U11533 (N_11533,N_9132,N_7059);
and U11534 (N_11534,N_8622,N_5218);
and U11535 (N_11535,N_9284,N_5574);
or U11536 (N_11536,N_5172,N_6544);
nor U11537 (N_11537,N_5913,N_8208);
or U11538 (N_11538,N_6528,N_8021);
or U11539 (N_11539,N_8698,N_8873);
nand U11540 (N_11540,N_8491,N_7293);
and U11541 (N_11541,N_8910,N_7113);
and U11542 (N_11542,N_5093,N_7936);
xnor U11543 (N_11543,N_6646,N_6133);
nand U11544 (N_11544,N_9581,N_6229);
or U11545 (N_11545,N_8502,N_5452);
nand U11546 (N_11546,N_9623,N_9564);
nor U11547 (N_11547,N_7552,N_6278);
nor U11548 (N_11548,N_6584,N_7765);
and U11549 (N_11549,N_7950,N_5514);
nand U11550 (N_11550,N_9323,N_5714);
xnor U11551 (N_11551,N_8444,N_7064);
and U11552 (N_11552,N_7820,N_5604);
and U11553 (N_11553,N_5254,N_7174);
nor U11554 (N_11554,N_6441,N_8150);
nand U11555 (N_11555,N_5509,N_9612);
or U11556 (N_11556,N_8923,N_5592);
nor U11557 (N_11557,N_9211,N_5492);
and U11558 (N_11558,N_6167,N_9357);
and U11559 (N_11559,N_6761,N_6994);
nand U11560 (N_11560,N_5751,N_9048);
and U11561 (N_11561,N_6232,N_7940);
and U11562 (N_11562,N_5849,N_8527);
nand U11563 (N_11563,N_6276,N_9681);
or U11564 (N_11564,N_5247,N_9400);
nand U11565 (N_11565,N_6850,N_7606);
or U11566 (N_11566,N_5105,N_7358);
and U11567 (N_11567,N_5374,N_5023);
nand U11568 (N_11568,N_8234,N_9910);
nand U11569 (N_11569,N_8122,N_6781);
nand U11570 (N_11570,N_8253,N_9318);
and U11571 (N_11571,N_5621,N_8202);
and U11572 (N_11572,N_9504,N_9895);
nand U11573 (N_11573,N_9619,N_7531);
or U11574 (N_11574,N_5753,N_6248);
nand U11575 (N_11575,N_7060,N_9937);
or U11576 (N_11576,N_7585,N_7671);
nand U11577 (N_11577,N_6789,N_5883);
xor U11578 (N_11578,N_6548,N_6351);
xnor U11579 (N_11579,N_9965,N_8711);
nor U11580 (N_11580,N_8918,N_6876);
and U11581 (N_11581,N_6258,N_8217);
nand U11582 (N_11582,N_5551,N_7052);
and U11583 (N_11583,N_8992,N_6589);
nor U11584 (N_11584,N_6526,N_5507);
nand U11585 (N_11585,N_9359,N_7910);
nand U11586 (N_11586,N_9041,N_6399);
or U11587 (N_11587,N_8905,N_9276);
or U11588 (N_11588,N_5796,N_8766);
nor U11589 (N_11589,N_6111,N_6866);
and U11590 (N_11590,N_5003,N_7072);
nor U11591 (N_11591,N_8237,N_7417);
nand U11592 (N_11592,N_7184,N_7546);
and U11593 (N_11593,N_9215,N_5848);
nor U11594 (N_11594,N_7243,N_7748);
and U11595 (N_11595,N_6922,N_6354);
nand U11596 (N_11596,N_7732,N_8872);
and U11597 (N_11597,N_9293,N_8681);
nand U11598 (N_11598,N_8190,N_5885);
or U11599 (N_11599,N_5745,N_6980);
nand U11600 (N_11600,N_9634,N_5541);
and U11601 (N_11601,N_7353,N_8830);
and U11602 (N_11602,N_8697,N_9494);
nand U11603 (N_11603,N_9147,N_7421);
and U11604 (N_11604,N_8980,N_8129);
and U11605 (N_11605,N_8995,N_8722);
nand U11606 (N_11606,N_6053,N_7687);
xor U11607 (N_11607,N_5625,N_6262);
or U11608 (N_11608,N_5649,N_9234);
and U11609 (N_11609,N_8075,N_6714);
and U11610 (N_11610,N_5995,N_7813);
nand U11611 (N_11611,N_6799,N_6139);
nand U11612 (N_11612,N_7600,N_5739);
or U11613 (N_11613,N_7811,N_7829);
and U11614 (N_11614,N_8597,N_9865);
and U11615 (N_11615,N_9340,N_7462);
nand U11616 (N_11616,N_7988,N_8929);
nor U11617 (N_11617,N_9107,N_8422);
nor U11618 (N_11618,N_6145,N_8572);
xor U11619 (N_11619,N_7051,N_6749);
nor U11620 (N_11620,N_5925,N_9573);
nor U11621 (N_11621,N_8942,N_9959);
and U11622 (N_11622,N_6459,N_9428);
nor U11623 (N_11623,N_9091,N_5632);
nand U11624 (N_11624,N_7202,N_6849);
and U11625 (N_11625,N_7458,N_6517);
or U11626 (N_11626,N_7083,N_7934);
nand U11627 (N_11627,N_5777,N_7755);
nand U11628 (N_11628,N_7854,N_8705);
nand U11629 (N_11629,N_7315,N_5563);
nand U11630 (N_11630,N_5071,N_7896);
xnor U11631 (N_11631,N_9960,N_7301);
nand U11632 (N_11632,N_6554,N_5528);
xor U11633 (N_11633,N_6401,N_7937);
and U11634 (N_11634,N_6512,N_5915);
or U11635 (N_11635,N_9378,N_9426);
or U11636 (N_11636,N_6874,N_8355);
nor U11637 (N_11637,N_5161,N_9890);
or U11638 (N_11638,N_6045,N_9497);
and U11639 (N_11639,N_6545,N_7329);
nand U11640 (N_11640,N_7784,N_5564);
nor U11641 (N_11641,N_7769,N_6440);
nor U11642 (N_11642,N_9052,N_8683);
or U11643 (N_11643,N_5484,N_5418);
xnor U11644 (N_11644,N_7500,N_5765);
nor U11645 (N_11645,N_5363,N_7157);
nor U11646 (N_11646,N_7928,N_6595);
and U11647 (N_11647,N_6180,N_5558);
and U11648 (N_11648,N_5398,N_9144);
nand U11649 (N_11649,N_6084,N_8116);
xor U11650 (N_11650,N_9672,N_9263);
and U11651 (N_11651,N_5805,N_8066);
nand U11652 (N_11652,N_5018,N_6796);
xor U11653 (N_11653,N_9387,N_5769);
xor U11654 (N_11654,N_7213,N_5075);
and U11655 (N_11655,N_8311,N_6578);
or U11656 (N_11656,N_6284,N_6118);
and U11657 (N_11657,N_8029,N_8546);
nor U11658 (N_11658,N_5338,N_7823);
nor U11659 (N_11659,N_9812,N_6269);
nand U11660 (N_11660,N_8175,N_5591);
or U11661 (N_11661,N_8434,N_5258);
nand U11662 (N_11662,N_5368,N_5958);
nand U11663 (N_11663,N_7380,N_9244);
or U11664 (N_11664,N_5011,N_5899);
nor U11665 (N_11665,N_6395,N_9776);
xnor U11666 (N_11666,N_7933,N_5337);
nand U11667 (N_11667,N_6024,N_7899);
nand U11668 (N_11668,N_9726,N_6161);
nor U11669 (N_11669,N_8241,N_8590);
nor U11670 (N_11670,N_7003,N_6317);
or U11671 (N_11671,N_8685,N_6481);
xnor U11672 (N_11672,N_8763,N_7688);
or U11673 (N_11673,N_8901,N_7570);
and U11674 (N_11674,N_6852,N_5973);
nand U11675 (N_11675,N_5738,N_7465);
nor U11676 (N_11676,N_6081,N_9823);
or U11677 (N_11677,N_8431,N_9415);
nor U11678 (N_11678,N_6625,N_7097);
and U11679 (N_11679,N_7708,N_9199);
nor U11680 (N_11680,N_6768,N_6904);
or U11681 (N_11681,N_9613,N_6807);
nand U11682 (N_11682,N_7582,N_9439);
xor U11683 (N_11683,N_6950,N_8513);
nand U11684 (N_11684,N_8451,N_9185);
and U11685 (N_11685,N_6929,N_9735);
or U11686 (N_11686,N_8297,N_7050);
and U11687 (N_11687,N_7453,N_9707);
nor U11688 (N_11688,N_5718,N_5190);
nor U11689 (N_11689,N_6129,N_8870);
and U11690 (N_11690,N_5997,N_6255);
and U11691 (N_11691,N_9193,N_9224);
nor U11692 (N_11692,N_6297,N_7248);
nand U11693 (N_11693,N_9913,N_5426);
nor U11694 (N_11694,N_7920,N_5829);
nand U11695 (N_11695,N_7496,N_9882);
nor U11696 (N_11696,N_5795,N_5478);
nand U11697 (N_11697,N_8215,N_6228);
xnor U11698 (N_11698,N_8700,N_9164);
and U11699 (N_11699,N_5409,N_7124);
xnor U11700 (N_11700,N_5489,N_5864);
nand U11701 (N_11701,N_6058,N_7244);
nand U11702 (N_11702,N_6287,N_9485);
and U11703 (N_11703,N_5573,N_8442);
nor U11704 (N_11704,N_9993,N_8908);
and U11705 (N_11705,N_9502,N_5748);
nor U11706 (N_11706,N_8866,N_9828);
nand U11707 (N_11707,N_6423,N_5732);
and U11708 (N_11708,N_5642,N_5171);
or U11709 (N_11709,N_6979,N_8183);
or U11710 (N_11710,N_6156,N_8113);
nor U11711 (N_11711,N_7266,N_6721);
nand U11712 (N_11712,N_5318,N_6956);
and U11713 (N_11713,N_5073,N_9272);
nor U11714 (N_11714,N_6552,N_8479);
and U11715 (N_11715,N_5562,N_5550);
xnor U11716 (N_11716,N_9717,N_9779);
xor U11717 (N_11717,N_7382,N_6119);
nor U11718 (N_11718,N_9399,N_7644);
or U11719 (N_11719,N_7286,N_5991);
or U11720 (N_11720,N_5534,N_8045);
nor U11721 (N_11721,N_5163,N_6561);
or U11722 (N_11722,N_6231,N_8153);
nand U11723 (N_11723,N_6411,N_5249);
nand U11724 (N_11724,N_6179,N_7351);
and U11725 (N_11725,N_5930,N_9239);
nor U11726 (N_11726,N_6622,N_8570);
nor U11727 (N_11727,N_5322,N_6294);
nand U11728 (N_11728,N_9875,N_6144);
or U11729 (N_11729,N_9900,N_9003);
nand U11730 (N_11730,N_5747,N_5835);
and U11731 (N_11731,N_8287,N_5097);
xor U11732 (N_11732,N_9819,N_8652);
and U11733 (N_11733,N_9720,N_7089);
xor U11734 (N_11734,N_8239,N_7491);
nand U11735 (N_11735,N_5599,N_7274);
and U11736 (N_11736,N_9080,N_5264);
or U11737 (N_11737,N_6689,N_7015);
nor U11738 (N_11738,N_5998,N_6104);
or U11739 (N_11739,N_7423,N_9881);
nand U11740 (N_11740,N_7488,N_5834);
nand U11741 (N_11741,N_5720,N_7133);
nand U11742 (N_11742,N_8495,N_8180);
and U11743 (N_11743,N_7839,N_9963);
nand U11744 (N_11744,N_8593,N_6957);
nand U11745 (N_11745,N_6062,N_8016);
xnor U11746 (N_11746,N_5954,N_7853);
and U11747 (N_11747,N_9159,N_8783);
and U11748 (N_11748,N_9078,N_8398);
and U11749 (N_11749,N_6961,N_5602);
nor U11750 (N_11750,N_7886,N_9325);
nor U11751 (N_11751,N_5863,N_8001);
nand U11752 (N_11752,N_6704,N_6992);
or U11753 (N_11753,N_9569,N_8781);
and U11754 (N_11754,N_5187,N_9909);
xor U11755 (N_11755,N_5996,N_9113);
nand U11756 (N_11756,N_5914,N_9542);
nand U11757 (N_11757,N_7499,N_9723);
nand U11758 (N_11758,N_9753,N_9759);
xor U11759 (N_11759,N_9197,N_6616);
nand U11760 (N_11760,N_5590,N_5362);
nand U11761 (N_11761,N_8848,N_6770);
nor U11762 (N_11762,N_5438,N_8712);
xor U11763 (N_11763,N_6955,N_5933);
nor U11764 (N_11764,N_9369,N_6669);
and U11765 (N_11765,N_6172,N_5121);
nor U11766 (N_11766,N_6384,N_5252);
xor U11767 (N_11767,N_5776,N_8605);
xor U11768 (N_11768,N_8657,N_6096);
nor U11769 (N_11769,N_8874,N_6848);
xor U11770 (N_11770,N_7998,N_9279);
or U11771 (N_11771,N_5196,N_8512);
nand U11772 (N_11772,N_5050,N_6038);
xnor U11773 (N_11773,N_8611,N_9851);
or U11774 (N_11774,N_5482,N_9047);
and U11775 (N_11775,N_9302,N_9491);
nand U11776 (N_11776,N_7990,N_5912);
nor U11777 (N_11777,N_7415,N_8362);
nor U11778 (N_11778,N_6489,N_7694);
nor U11779 (N_11779,N_5658,N_5034);
or U11780 (N_11780,N_7121,N_5389);
nor U11781 (N_11781,N_7878,N_7280);
nor U11782 (N_11782,N_7073,N_5854);
or U11783 (N_11783,N_8639,N_6719);
and U11784 (N_11784,N_9657,N_6759);
xor U11785 (N_11785,N_7276,N_5497);
and U11786 (N_11786,N_9611,N_7594);
and U11787 (N_11787,N_5066,N_8540);
nor U11788 (N_11788,N_6775,N_7416);
nand U11789 (N_11789,N_9924,N_8519);
nor U11790 (N_11790,N_7237,N_9802);
nor U11791 (N_11791,N_5067,N_5955);
and U11792 (N_11792,N_6535,N_6581);
or U11793 (N_11793,N_6617,N_9811);
nand U11794 (N_11794,N_9521,N_7885);
and U11795 (N_11795,N_6538,N_6712);
or U11796 (N_11796,N_8051,N_9348);
nor U11797 (N_11797,N_9029,N_9709);
nand U11798 (N_11798,N_6510,N_5654);
xor U11799 (N_11799,N_5868,N_7039);
and U11800 (N_11800,N_9140,N_9671);
nor U11801 (N_11801,N_8436,N_5230);
nand U11802 (N_11802,N_6751,N_6181);
or U11803 (N_11803,N_9597,N_7019);
xor U11804 (N_11804,N_9577,N_8363);
nand U11805 (N_11805,N_5513,N_9077);
xnor U11806 (N_11806,N_7845,N_6988);
xor U11807 (N_11807,N_9471,N_5211);
and U11808 (N_11808,N_7642,N_5578);
or U11809 (N_11809,N_5145,N_5744);
nor U11810 (N_11810,N_7300,N_5511);
or U11811 (N_11811,N_8291,N_5623);
nand U11812 (N_11812,N_7880,N_7601);
and U11813 (N_11813,N_7915,N_7457);
or U11814 (N_11814,N_6603,N_7261);
or U11815 (N_11815,N_9730,N_9645);
or U11816 (N_11816,N_9814,N_5354);
nor U11817 (N_11817,N_7267,N_5304);
nor U11818 (N_11818,N_9116,N_8488);
or U11819 (N_11819,N_7145,N_7716);
and U11820 (N_11820,N_9310,N_8974);
nand U11821 (N_11821,N_5787,N_7478);
or U11822 (N_11822,N_6204,N_9479);
nor U11823 (N_11823,N_6455,N_5635);
nor U11824 (N_11824,N_6684,N_8423);
nor U11825 (N_11825,N_9297,N_5895);
nor U11826 (N_11826,N_5806,N_5607);
nand U11827 (N_11827,N_7834,N_6209);
and U11828 (N_11828,N_9761,N_7993);
nand U11829 (N_11829,N_7366,N_8774);
xor U11830 (N_11830,N_5859,N_5721);
nand U11831 (N_11831,N_7786,N_9967);
nor U11832 (N_11832,N_9799,N_6657);
or U11833 (N_11833,N_6976,N_5040);
xor U11834 (N_11834,N_9181,N_6557);
nand U11835 (N_11835,N_8928,N_9162);
and U11836 (N_11836,N_7926,N_8924);
nor U11837 (N_11837,N_9424,N_9787);
nand U11838 (N_11838,N_7074,N_5627);
nor U11839 (N_11839,N_7150,N_5762);
xnor U11840 (N_11840,N_7619,N_6383);
and U11841 (N_11841,N_5694,N_9607);
and U11842 (N_11842,N_8379,N_8134);
or U11843 (N_11843,N_5907,N_8477);
or U11844 (N_11844,N_6374,N_8462);
nor U11845 (N_11845,N_9376,N_7646);
or U11846 (N_11846,N_5005,N_8334);
or U11847 (N_11847,N_6324,N_6357);
nor U11848 (N_11848,N_8171,N_7148);
nor U11849 (N_11849,N_6790,N_5353);
nand U11850 (N_11850,N_9482,N_5021);
nand U11851 (N_11851,N_9031,N_6001);
and U11852 (N_11852,N_9826,N_8111);
and U11853 (N_11853,N_7803,N_8979);
or U11854 (N_11854,N_8769,N_5248);
nand U11855 (N_11855,N_7486,N_7968);
nor U11856 (N_11856,N_8886,N_9121);
nor U11857 (N_11857,N_9532,N_5510);
or U11858 (N_11858,N_9926,N_5479);
nand U11859 (N_11859,N_7144,N_8207);
and U11860 (N_11860,N_6465,N_8199);
nor U11861 (N_11861,N_9889,N_6703);
nor U11862 (N_11862,N_9448,N_7287);
and U11863 (N_11863,N_6298,N_7894);
nand U11864 (N_11864,N_5147,N_6164);
or U11865 (N_11865,N_5393,N_9059);
or U11866 (N_11866,N_9221,N_7138);
nand U11867 (N_11867,N_6115,N_8464);
nand U11868 (N_11868,N_7872,N_6920);
nand U11869 (N_11869,N_7281,N_5775);
nor U11870 (N_11870,N_9347,N_7947);
nand U11871 (N_11871,N_9894,N_6843);
nor U11872 (N_11872,N_7428,N_8377);
nand U11873 (N_11873,N_9377,N_7197);
nand U11874 (N_11874,N_6125,N_7154);
nor U11875 (N_11875,N_7741,N_9474);
or U11876 (N_11876,N_7206,N_7489);
or U11877 (N_11877,N_6604,N_8740);
or U11878 (N_11878,N_7481,N_5810);
nand U11879 (N_11879,N_7025,N_6518);
and U11880 (N_11880,N_9858,N_5153);
nor U11881 (N_11881,N_9842,N_5115);
nand U11882 (N_11882,N_8367,N_5758);
nand U11883 (N_11883,N_8642,N_9202);
and U11884 (N_11884,N_9874,N_5846);
and U11885 (N_11885,N_7909,N_5198);
and U11886 (N_11886,N_7125,N_6910);
xnor U11887 (N_11887,N_7918,N_5149);
nor U11888 (N_11888,N_8004,N_5117);
nor U11889 (N_11889,N_9630,N_7778);
or U11890 (N_11890,N_9574,N_7753);
xnor U11891 (N_11891,N_9446,N_7302);
nand U11892 (N_11892,N_8246,N_8620);
or U11893 (N_11893,N_9518,N_9286);
or U11894 (N_11894,N_5136,N_7943);
and U11895 (N_11895,N_7789,N_7881);
nor U11896 (N_11896,N_8429,N_9189);
and U11897 (N_11897,N_5417,N_6792);
xor U11898 (N_11898,N_8650,N_5499);
nand U11899 (N_11899,N_9292,N_8852);
nand U11900 (N_11900,N_9068,N_5447);
and U11901 (N_11901,N_6039,N_6745);
and U11902 (N_11902,N_6577,N_6609);
and U11903 (N_11903,N_7088,N_9986);
or U11904 (N_11904,N_8168,N_9676);
xor U11905 (N_11905,N_5358,N_7873);
and U11906 (N_11906,N_6305,N_7367);
or U11907 (N_11907,N_7323,N_5633);
nor U11908 (N_11908,N_8308,N_9969);
nand U11909 (N_11909,N_9918,N_8518);
and U11910 (N_11910,N_5943,N_6237);
and U11911 (N_11911,N_9582,N_8466);
or U11912 (N_11912,N_8054,N_5279);
or U11913 (N_11913,N_7905,N_5180);
nand U11914 (N_11914,N_7835,N_9062);
nand U11915 (N_11915,N_6485,N_5935);
nand U11916 (N_11916,N_9015,N_5142);
xor U11917 (N_11917,N_6708,N_8392);
nand U11918 (N_11918,N_9744,N_6764);
or U11919 (N_11919,N_5617,N_7471);
and U11920 (N_11920,N_5782,N_9886);
xnor U11921 (N_11921,N_7495,N_8421);
nand U11922 (N_11922,N_9879,N_9384);
nor U11923 (N_11923,N_8396,N_6926);
nand U11924 (N_11924,N_7128,N_8730);
xnor U11925 (N_11925,N_9571,N_5821);
xnor U11926 (N_11926,N_8330,N_7477);
nor U11927 (N_11927,N_8249,N_9810);
and U11928 (N_11928,N_9715,N_5296);
nor U11929 (N_11929,N_8376,N_6786);
xor U11930 (N_11930,N_8521,N_5096);
nor U11931 (N_11931,N_8955,N_8440);
and U11932 (N_11932,N_8664,N_5756);
nor U11933 (N_11933,N_9821,N_9264);
nor U11934 (N_11934,N_6155,N_8723);
xor U11935 (N_11935,N_7098,N_5072);
nand U11936 (N_11936,N_5962,N_7738);
and U11937 (N_11937,N_7932,N_8941);
xnor U11938 (N_11938,N_8404,N_6362);
nor U11939 (N_11939,N_8493,N_6547);
xor U11940 (N_11940,N_6326,N_8069);
nor U11941 (N_11941,N_6307,N_6868);
nor U11942 (N_11942,N_7018,N_9201);
nor U11943 (N_11943,N_9928,N_5719);
nor U11944 (N_11944,N_7537,N_8448);
and U11945 (N_11945,N_6797,N_6268);
xor U11946 (N_11946,N_6739,N_6539);
nand U11947 (N_11947,N_8785,N_5428);
nand U11948 (N_11948,N_8850,N_7216);
or U11949 (N_11949,N_9393,N_9414);
and U11950 (N_11950,N_6196,N_6880);
nand U11951 (N_11951,N_8721,N_5377);
or U11952 (N_11952,N_5728,N_9472);
nor U11953 (N_11953,N_9432,N_7696);
and U11954 (N_11954,N_6871,N_8727);
or U11955 (N_11955,N_7837,N_9094);
nand U11956 (N_11956,N_5219,N_9236);
or U11957 (N_11957,N_5717,N_8998);
or U11958 (N_11958,N_8149,N_6206);
or U11959 (N_11959,N_6897,N_9403);
nor U11960 (N_11960,N_6173,N_5917);
or U11961 (N_11961,N_5965,N_9545);
or U11962 (N_11962,N_5084,N_5524);
xor U11963 (N_11963,N_9277,N_5159);
nor U11964 (N_11964,N_7322,N_6707);
xor U11965 (N_11965,N_9065,N_6325);
xor U11966 (N_11966,N_6573,N_8753);
or U11967 (N_11967,N_9008,N_9304);
nand U11968 (N_11968,N_7070,N_9109);
xor U11969 (N_11969,N_9260,N_5421);
nand U11970 (N_11970,N_5659,N_6430);
xor U11971 (N_11971,N_5403,N_7736);
and U11972 (N_11972,N_5245,N_9985);
and U11973 (N_11973,N_9636,N_8676);
nor U11974 (N_11974,N_6078,N_6072);
or U11975 (N_11975,N_6986,N_8759);
xnor U11976 (N_11976,N_7650,N_5108);
nand U11977 (N_11977,N_5866,N_8304);
or U11978 (N_11978,N_8201,N_9167);
nand U11979 (N_11979,N_9689,N_5458);
nand U11980 (N_11980,N_5576,N_9139);
and U11981 (N_11981,N_6709,N_5516);
or U11982 (N_11982,N_9195,N_5799);
xor U11983 (N_11983,N_8267,N_6643);
xnor U11984 (N_11984,N_5960,N_6050);
nand U11985 (N_11985,N_9737,N_6000);
nand U11986 (N_11986,N_6142,N_5531);
and U11987 (N_11987,N_9412,N_5467);
xor U11988 (N_11988,N_5269,N_8476);
and U11989 (N_11989,N_9408,N_7324);
or U11990 (N_11990,N_9758,N_6902);
nand U11991 (N_11991,N_7685,N_7622);
nor U11992 (N_11992,N_7618,N_8931);
nand U11993 (N_11993,N_8653,N_8768);
and U11994 (N_11994,N_8467,N_6124);
nand U11995 (N_11995,N_9434,N_8151);
or U11996 (N_11996,N_6388,N_7482);
nand U11997 (N_11997,N_6734,N_9430);
nand U11998 (N_11998,N_6982,N_6421);
and U11999 (N_11999,N_6672,N_8090);
nor U12000 (N_12000,N_5702,N_7856);
nand U12001 (N_12001,N_9549,N_7376);
and U12002 (N_12002,N_7149,N_5241);
nand U12003 (N_12003,N_7312,N_6368);
nand U12004 (N_12004,N_9129,N_9022);
nand U12005 (N_12005,N_7533,N_8509);
nor U12006 (N_12006,N_6597,N_7443);
nand U12007 (N_12007,N_9443,N_7587);
and U12008 (N_12008,N_6454,N_9451);
nand U12009 (N_12009,N_7520,N_6588);
or U12010 (N_12010,N_7817,N_6934);
nand U12011 (N_12011,N_9696,N_6881);
nor U12012 (N_12012,N_9679,N_7604);
nand U12013 (N_12013,N_7868,N_6682);
and U12014 (N_12014,N_9425,N_7704);
and U12015 (N_12015,N_9508,N_7860);
nor U12016 (N_12016,N_5167,N_6289);
nand U12017 (N_12017,N_7403,N_8470);
or U12018 (N_12018,N_9217,N_8912);
nand U12019 (N_12019,N_8939,N_6346);
or U12020 (N_12020,N_8119,N_5302);
and U12021 (N_12021,N_9098,N_7258);
and U12022 (N_12022,N_9242,N_6467);
xor U12023 (N_12023,N_7316,N_6921);
and U12024 (N_12024,N_8214,N_5579);
nand U12025 (N_12025,N_6551,N_6497);
and U12026 (N_12026,N_9203,N_6425);
or U12027 (N_12027,N_8475,N_5014);
nor U12028 (N_12028,N_8684,N_9757);
or U12029 (N_12029,N_5429,N_5029);
nor U12030 (N_12030,N_8179,N_7238);
or U12031 (N_12031,N_6093,N_8575);
or U12032 (N_12032,N_9745,N_8532);
nor U12033 (N_12033,N_9460,N_7508);
or U12034 (N_12034,N_6132,N_8012);
and U12035 (N_12035,N_9463,N_6068);
or U12036 (N_12036,N_9982,N_7729);
or U12037 (N_12037,N_5371,N_6429);
and U12038 (N_12038,N_7770,N_9405);
or U12039 (N_12039,N_9561,N_5306);
nor U12040 (N_12040,N_9903,N_9322);
nand U12041 (N_12041,N_8329,N_5274);
or U12042 (N_12042,N_6858,N_6811);
and U12043 (N_12043,N_9983,N_9927);
and U12044 (N_12044,N_5723,N_7690);
nand U12045 (N_12045,N_8831,N_7236);
xnor U12046 (N_12046,N_5838,N_9996);
and U12047 (N_12047,N_8696,N_9037);
and U12048 (N_12048,N_9257,N_7318);
nor U12049 (N_12049,N_6193,N_9243);
nand U12050 (N_12050,N_9747,N_8020);
nand U12051 (N_12051,N_9213,N_6245);
nand U12052 (N_12052,N_8699,N_5575);
and U12053 (N_12053,N_8255,N_5216);
xor U12054 (N_12054,N_5289,N_7211);
xor U12055 (N_12055,N_6788,N_5927);
nand U12056 (N_12056,N_5036,N_8808);
and U12057 (N_12057,N_7529,N_5937);
xor U12058 (N_12058,N_7288,N_7396);
xor U12059 (N_12059,N_8002,N_8380);
nor U12060 (N_12060,N_8059,N_5475);
and U12061 (N_12061,N_7962,N_7623);
or U12062 (N_12062,N_8463,N_6795);
nor U12063 (N_12063,N_7922,N_8446);
and U12064 (N_12064,N_8108,N_9553);
nor U12065 (N_12065,N_5733,N_5462);
nand U12066 (N_12066,N_6312,N_5643);
nand U12067 (N_12067,N_6560,N_6668);
or U12068 (N_12068,N_5307,N_5111);
or U12069 (N_12069,N_7129,N_5146);
nor U12070 (N_12070,N_5399,N_6925);
nand U12071 (N_12071,N_9552,N_8152);
or U12072 (N_12072,N_5346,N_7621);
nand U12073 (N_12073,N_9373,N_7298);
and U12074 (N_12074,N_9932,N_8606);
and U12075 (N_12075,N_6221,N_7132);
nand U12076 (N_12076,N_8167,N_9496);
nand U12077 (N_12077,N_7776,N_5103);
or U12078 (N_12078,N_5977,N_6686);
and U12079 (N_12079,N_6842,N_6242);
or U12080 (N_12080,N_5894,N_8754);
and U12081 (N_12081,N_7378,N_7151);
or U12082 (N_12082,N_7682,N_6077);
and U12083 (N_12083,N_8351,N_7204);
or U12084 (N_12084,N_6063,N_7864);
and U12085 (N_12085,N_5282,N_6673);
xor U12086 (N_12086,N_6328,N_9566);
nand U12087 (N_12087,N_9579,N_7101);
nand U12088 (N_12088,N_6054,N_8348);
nand U12089 (N_12089,N_7530,N_8136);
nor U12090 (N_12090,N_7299,N_7075);
and U12091 (N_12091,N_7468,N_8316);
or U12092 (N_12092,N_9064,N_7639);
xnor U12093 (N_12093,N_7303,N_5232);
nand U12094 (N_12094,N_8934,N_6590);
nand U12095 (N_12095,N_8825,N_8289);
and U12096 (N_12096,N_7935,N_8707);
or U12097 (N_12097,N_5900,N_6106);
nor U12098 (N_12098,N_6648,N_8689);
or U12099 (N_12099,N_9741,N_7334);
nand U12100 (N_12100,N_9840,N_6691);
or U12101 (N_12101,N_6487,N_5074);
and U12102 (N_12102,N_8673,N_5430);
nand U12103 (N_12103,N_7858,N_8729);
and U12104 (N_12104,N_5628,N_6537);
nand U12105 (N_12105,N_8975,N_9396);
nand U12106 (N_12106,N_6286,N_5287);
nand U12107 (N_12107,N_6048,N_7418);
and U12108 (N_12108,N_9640,N_5540);
nand U12109 (N_12109,N_9970,N_6923);
nand U12110 (N_12110,N_8859,N_9058);
or U12111 (N_12111,N_7401,N_8771);
xnor U12112 (N_12112,N_5173,N_5110);
nand U12113 (N_12113,N_8053,N_9191);
or U12114 (N_12114,N_5566,N_6793);
and U12115 (N_12115,N_9392,N_5178);
nand U12116 (N_12116,N_8577,N_7086);
nor U12117 (N_12117,N_8288,N_6197);
nor U12118 (N_12118,N_8591,N_7557);
and U12119 (N_12119,N_7567,N_7115);
nand U12120 (N_12120,N_7066,N_5080);
nor U12121 (N_12121,N_5896,N_6938);
xor U12122 (N_12122,N_9736,N_6996);
nor U12123 (N_12123,N_7961,N_5956);
nand U12124 (N_12124,N_8735,N_8579);
and U12125 (N_12125,N_8500,N_5027);
xor U12126 (N_12126,N_9815,N_6247);
or U12127 (N_12127,N_6484,N_9713);
or U12128 (N_12128,N_5975,N_6065);
nor U12129 (N_12129,N_9228,N_7123);
nand U12130 (N_12130,N_7714,N_5288);
and U12131 (N_12131,N_9733,N_8560);
and U12132 (N_12132,N_7172,N_9007);
or U12133 (N_12133,N_8972,N_8204);
nand U12134 (N_12134,N_9218,N_5983);
nand U12135 (N_12135,N_8323,N_7037);
or U12136 (N_12136,N_6534,N_9372);
nor U12137 (N_12137,N_6837,N_7526);
xnor U12138 (N_12138,N_8317,N_7095);
and U12139 (N_12139,N_8469,N_5035);
or U12140 (N_12140,N_6942,N_6348);
and U12141 (N_12141,N_9301,N_7867);
and U12142 (N_12142,N_5114,N_6814);
or U12143 (N_12143,N_9267,N_9598);
or U12144 (N_12144,N_5549,N_8292);
and U12145 (N_12145,N_7155,N_9417);
or U12146 (N_12146,N_6292,N_5025);
nand U12147 (N_12147,N_6389,N_8216);
or U12148 (N_12148,N_7000,N_6715);
xnor U12149 (N_12149,N_8865,N_5004);
nand U12150 (N_12150,N_9305,N_5315);
xnor U12151 (N_12151,N_5469,N_9912);
nand U12152 (N_12152,N_6503,N_5783);
and U12153 (N_12153,N_7747,N_8091);
and U12154 (N_12154,N_8567,N_6002);
or U12155 (N_12155,N_8706,N_9092);
nand U12156 (N_12156,N_7412,N_7422);
or U12157 (N_12157,N_8082,N_5653);
nor U12158 (N_12158,N_9161,N_9503);
and U12159 (N_12159,N_5405,N_8840);
nand U12160 (N_12160,N_7951,N_5347);
or U12161 (N_12161,N_8353,N_5222);
nor U12162 (N_12162,N_6627,N_9253);
xnor U12163 (N_12163,N_9684,N_8017);
nand U12164 (N_12164,N_7640,N_6724);
nand U12165 (N_12165,N_9174,N_9666);
nand U12166 (N_12166,N_8453,N_9772);
nand U12167 (N_12167,N_7603,N_5175);
and U12168 (N_12168,N_5379,N_6308);
and U12169 (N_12169,N_7902,N_6090);
xor U12170 (N_12170,N_6967,N_5773);
nand U12171 (N_12171,N_7818,N_5790);
xor U12172 (N_12172,N_7561,N_5275);
nor U12173 (N_12173,N_9885,N_7080);
and U12174 (N_12174,N_6601,N_5276);
nor U12175 (N_12175,N_6281,N_6987);
or U12176 (N_12176,N_7463,N_6809);
and U12177 (N_12177,N_7565,N_6250);
or U12178 (N_12178,N_5543,N_8656);
nor U12179 (N_12179,N_6766,N_7167);
nand U12180 (N_12180,N_6605,N_9961);
nand U12181 (N_12181,N_7890,N_8813);
nor U12182 (N_12182,N_5370,N_5662);
and U12183 (N_12183,N_5195,N_7296);
nor U12184 (N_12184,N_5707,N_7511);
and U12185 (N_12185,N_5542,N_8543);
nor U12186 (N_12186,N_8157,N_5104);
and U12187 (N_12187,N_5808,N_5980);
and U12188 (N_12188,N_5554,N_8437);
nand U12189 (N_12189,N_5056,N_5415);
nand U12190 (N_12190,N_8810,N_5406);
or U12191 (N_12191,N_6428,N_7980);
nand U12192 (N_12192,N_6758,N_5155);
nor U12193 (N_12193,N_7355,N_9930);
nor U12194 (N_12194,N_5107,N_5106);
nand U12195 (N_12195,N_8623,N_8205);
or U12196 (N_12196,N_7446,N_6741);
or U12197 (N_12197,N_6148,N_9038);
and U12198 (N_12198,N_9060,N_5886);
or U12199 (N_12199,N_9510,N_5832);
and U12200 (N_12200,N_9334,N_8098);
and U12201 (N_12201,N_6891,N_6079);
nor U12202 (N_12202,N_8481,N_6981);
or U12203 (N_12203,N_8625,N_6611);
and U12204 (N_12204,N_6170,N_7464);
or U12205 (N_12205,N_7256,N_9791);
nand U12206 (N_12206,N_9000,N_5512);
nor U12207 (N_12207,N_9105,N_6030);
nand U12208 (N_12208,N_7648,N_6697);
nand U12209 (N_12209,N_8093,N_6596);
or U12210 (N_12210,N_5878,N_6105);
or U12211 (N_12211,N_6917,N_5877);
nand U12212 (N_12212,N_9528,N_7810);
nor U12213 (N_12213,N_9822,N_5380);
xnor U12214 (N_12214,N_6508,N_8263);
or U12215 (N_12215,N_6524,N_8827);
and U12216 (N_12216,N_6103,N_5042);
nand U12217 (N_12217,N_6295,N_9445);
nand U12218 (N_12218,N_7304,N_7772);
nor U12219 (N_12219,N_8633,N_8636);
and U12220 (N_12220,N_8220,N_9901);
and U12221 (N_12221,N_7114,N_8511);
nor U12222 (N_12222,N_5431,N_5143);
and U12223 (N_12223,N_8443,N_6735);
or U12224 (N_12224,N_7780,N_5327);
nor U12225 (N_12225,N_6542,N_6999);
nor U12226 (N_12226,N_6117,N_6835);
and U12227 (N_12227,N_7110,N_9240);
and U12228 (N_12228,N_8225,N_5082);
nand U12229 (N_12229,N_5646,N_8907);
and U12230 (N_12230,N_6359,N_6744);
nor U12231 (N_12231,N_6521,N_6805);
nand U12232 (N_12232,N_8127,N_5382);
and U12233 (N_12233,N_7249,N_7513);
and U12234 (N_12234,N_6460,N_8958);
nand U12235 (N_12235,N_9605,N_8556);
xnor U12236 (N_12236,N_5301,N_6687);
and U12237 (N_12237,N_8356,N_5700);
nor U12238 (N_12238,N_7969,N_7616);
xor U12239 (N_12239,N_6710,N_7576);
and U12240 (N_12240,N_5548,N_5968);
nand U12241 (N_12241,N_5094,N_6918);
or U12242 (N_12242,N_8603,N_7849);
or U12243 (N_12243,N_9576,N_7136);
or U12244 (N_12244,N_6514,N_5948);
xor U12245 (N_12245,N_8299,N_5697);
or U12246 (N_12246,N_8881,N_9142);
nor U12247 (N_12247,N_6519,N_7385);
and U12248 (N_12248,N_5179,N_8490);
nor U12249 (N_12249,N_9061,N_5820);
or U12250 (N_12250,N_6187,N_6159);
or U12251 (N_12251,N_9800,N_7321);
xnor U12252 (N_12252,N_9643,N_5132);
xor U12253 (N_12253,N_6138,N_8009);
nand U12254 (N_12254,N_7308,N_7490);
or U12255 (N_12255,N_6338,N_9442);
and U12256 (N_12256,N_5555,N_5668);
nand U12257 (N_12257,N_9120,N_9487);
nand U12258 (N_12258,N_5435,N_9525);
xnor U12259 (N_12259,N_9974,N_5392);
nor U12260 (N_12260,N_9575,N_7023);
nor U12261 (N_12261,N_5177,N_8078);
nor U12262 (N_12262,N_6073,N_7540);
nand U12263 (N_12263,N_6121,N_9391);
or U12264 (N_12264,N_8693,N_5506);
nor U12265 (N_12265,N_7653,N_9481);
or U12266 (N_12266,N_6974,N_6075);
nor U12267 (N_12267,N_5351,N_7137);
nor U12268 (N_12268,N_6349,N_6171);
nor U12269 (N_12269,N_7319,N_9437);
or U12270 (N_12270,N_5709,N_5046);
nand U12271 (N_12271,N_8432,N_7665);
nor U12272 (N_12272,N_9691,N_5271);
nand U12273 (N_12273,N_5048,N_7795);
and U12274 (N_12274,N_8015,N_7283);
nand U12275 (N_12275,N_5788,N_7797);
nor U12276 (N_12276,N_9040,N_8023);
and U12277 (N_12277,N_9099,N_8257);
and U12278 (N_12278,N_5616,N_9069);
or U12279 (N_12279,N_9767,N_7395);
and U12280 (N_12280,N_8170,N_8745);
xnor U12281 (N_12281,N_8795,N_6210);
nand U12282 (N_12282,N_8647,N_6137);
or U12283 (N_12283,N_5152,N_5255);
or U12284 (N_12284,N_9813,N_6563);
and U12285 (N_12285,N_5138,N_8550);
or U12286 (N_12286,N_8790,N_8281);
nor U12287 (N_12287,N_8247,N_6040);
or U12288 (N_12288,N_6882,N_8758);
nor U12289 (N_12289,N_6085,N_6931);
and U12290 (N_12290,N_8659,N_8692);
xnor U12291 (N_12291,N_5850,N_9843);
nand U12292 (N_12292,N_8033,N_9173);
nor U12293 (N_12293,N_6991,N_8691);
nor U12294 (N_12294,N_8256,N_5022);
nor U12295 (N_12295,N_6402,N_5845);
and U12296 (N_12296,N_6345,N_5156);
nand U12297 (N_12297,N_5596,N_9933);
nand U12298 (N_12298,N_9128,N_7390);
nor U12299 (N_12299,N_6699,N_5678);
or U12300 (N_12300,N_9921,N_5019);
nor U12301 (N_12301,N_8762,N_6779);
nor U12302 (N_12302,N_7217,N_7842);
nor U12303 (N_12303,N_7068,N_9625);
xnor U12304 (N_12304,N_6086,N_7746);
and U12305 (N_12305,N_8212,N_8096);
or U12306 (N_12306,N_6023,N_5842);
xnor U12307 (N_12307,N_8022,N_5047);
or U12308 (N_12308,N_5053,N_7799);
or U12309 (N_12309,N_6569,N_5090);
nand U12310 (N_12310,N_6215,N_7675);
or U12311 (N_12311,N_8818,N_6895);
xor U12312 (N_12312,N_7522,N_6505);
nand U12313 (N_12313,N_8731,N_7681);
nand U12314 (N_12314,N_5151,N_5355);
and U12315 (N_12315,N_9682,N_7034);
nand U12316 (N_12316,N_7196,N_9409);
or U12317 (N_12317,N_9841,N_9266);
and U12318 (N_12318,N_6948,N_8333);
and U12319 (N_12319,N_8458,N_9249);
or U12320 (N_12320,N_9343,N_8485);
nand U12321 (N_12321,N_9450,N_6854);
nor U12322 (N_12322,N_5981,N_7824);
and U12323 (N_12323,N_8788,N_5737);
and U12324 (N_12324,N_8789,N_6555);
xor U12325 (N_12325,N_8143,N_8280);
nand U12326 (N_12326,N_7410,N_8680);
and U12327 (N_12327,N_6360,N_8514);
nand U12328 (N_12328,N_6525,N_6568);
nand U12329 (N_12329,N_8672,N_5833);
nor U12330 (N_12330,N_8251,N_5192);
nor U12331 (N_12331,N_7102,N_8956);
or U12332 (N_12332,N_8538,N_6606);
or U12333 (N_12333,N_7689,N_9118);
xor U12334 (N_12334,N_5319,N_6964);
or U12335 (N_12335,N_6962,N_7225);
nor U12336 (N_12336,N_6822,N_8843);
nand U12337 (N_12337,N_8087,N_6418);
and U12338 (N_12338,N_5704,N_7643);
or U12339 (N_12339,N_9339,N_6026);
and U12340 (N_12340,N_6783,N_8047);
xnor U12341 (N_12341,N_9419,N_7673);
nor U12342 (N_12342,N_5323,N_7164);
xor U12343 (N_12343,N_6765,N_9700);
nand U12344 (N_12344,N_7660,N_6211);
or U12345 (N_12345,N_9110,N_9364);
nand U12346 (N_12346,N_5792,N_9659);
nor U12347 (N_12347,N_9642,N_7966);
nand U12348 (N_12348,N_9855,N_5804);
and U12349 (N_12349,N_5069,N_9085);
or U12350 (N_12350,N_8951,N_6919);
and U12351 (N_12351,N_7328,N_5757);
xnor U12352 (N_12352,N_5814,N_7607);
xnor U12353 (N_12353,N_5285,N_5228);
nor U12354 (N_12354,N_6049,N_8793);
nor U12355 (N_12355,N_9076,N_8990);
nor U12356 (N_12356,N_5567,N_9212);
xnor U12357 (N_12357,N_6296,N_7069);
or U12358 (N_12358,N_5891,N_6380);
nand U12359 (N_12359,N_8816,N_5295);
nor U12360 (N_12360,N_9188,N_7474);
xor U12361 (N_12361,N_6358,N_5317);
nor U12362 (N_12362,N_5572,N_9333);
and U12363 (N_12363,N_7870,N_6257);
or U12364 (N_12364,N_7205,N_9423);
nor U12365 (N_12365,N_9911,N_5336);
nor U12366 (N_12366,N_8517,N_8195);
or U12367 (N_12367,N_9653,N_6911);
or U12368 (N_12368,N_5357,N_7473);
or U12369 (N_12369,N_6463,N_9389);
or U12370 (N_12370,N_6916,N_5601);
and U12371 (N_12371,N_8417,N_8739);
and U12372 (N_12372,N_7703,N_7904);
or U12373 (N_12373,N_9169,N_8382);
or U12374 (N_12374,N_6959,N_9280);
and U12375 (N_12375,N_7903,N_8117);
or U12376 (N_12376,N_7506,N_6226);
nand U12377 (N_12377,N_8182,N_7373);
nor U12378 (N_12378,N_9356,N_7278);
and U12379 (N_12379,N_6320,N_7090);
nor U12380 (N_12380,N_9789,N_5648);
nor U12381 (N_12381,N_5013,N_9987);
and U12382 (N_12382,N_7338,N_6633);
and U12383 (N_12383,N_8364,N_8996);
xnor U12384 (N_12384,N_9370,N_6816);
nand U12385 (N_12385,N_8340,N_7720);
or U12386 (N_12386,N_7762,N_5166);
and U12387 (N_12387,N_9820,N_8563);
or U12388 (N_12388,N_7285,N_7573);
or U12389 (N_12389,N_8332,N_5091);
or U12390 (N_12390,N_8764,N_7554);
and U12391 (N_12391,N_9287,N_7693);
nand U12392 (N_12392,N_8851,N_7726);
or U12393 (N_12393,N_9150,N_9112);
xnor U12394 (N_12394,N_6676,N_7027);
nand U12395 (N_12395,N_7543,N_6651);
xor U12396 (N_12396,N_8219,N_6649);
and U12397 (N_12397,N_5536,N_5938);
nor U12398 (N_12398,N_8038,N_8617);
nor U12399 (N_12399,N_6224,N_8669);
nor U12400 (N_12400,N_5987,N_5711);
or U12401 (N_12401,N_6095,N_8885);
and U12402 (N_12402,N_6731,N_6166);
nand U12403 (N_12403,N_9404,N_9554);
xor U12404 (N_12404,N_6675,N_9352);
nor U12405 (N_12405,N_9832,N_5580);
xnor U12406 (N_12406,N_8254,N_9055);
nor U12407 (N_12407,N_9562,N_8890);
and U12408 (N_12408,N_5784,N_7733);
and U12409 (N_12409,N_5679,N_8320);
or U12410 (N_12410,N_8424,N_9977);
nand U12411 (N_12411,N_9615,N_7832);
and U12412 (N_12412,N_7203,N_9665);
and U12413 (N_12413,N_6867,N_9464);
and U12414 (N_12414,N_5470,N_7342);
nor U12415 (N_12415,N_9899,N_8896);
or U12416 (N_12416,N_6630,N_5283);
or U12417 (N_12417,N_7058,N_9907);
and U12418 (N_12418,N_6694,N_7413);
nand U12419 (N_12419,N_9798,N_9032);
and U12420 (N_12420,N_7251,N_8746);
nand U12421 (N_12421,N_8801,N_5743);
or U12422 (N_12422,N_6303,N_7645);
and U12423 (N_12423,N_9944,N_6587);
and U12424 (N_12424,N_6218,N_8599);
nand U12425 (N_12425,N_6107,N_6438);
nor U12426 (N_12426,N_5505,N_5444);
and U12427 (N_12427,N_9406,N_8588);
and U12428 (N_12428,N_8970,N_6398);
nor U12429 (N_12429,N_8011,N_6141);
nor U12430 (N_12430,N_5690,N_8187);
or U12431 (N_12431,N_7889,N_5880);
xor U12432 (N_12432,N_6949,N_5133);
and U12433 (N_12433,N_9991,N_5112);
nand U12434 (N_12434,N_6140,N_7445);
xnor U12435 (N_12435,N_8889,N_5341);
nand U12436 (N_12436,N_6378,N_6110);
nor U12437 (N_12437,N_5726,N_5605);
nor U12438 (N_12438,N_8609,N_8374);
and U12439 (N_12439,N_9698,N_7313);
and U12440 (N_12440,N_8034,N_5944);
and U12441 (N_12441,N_6794,N_7804);
nand U12442 (N_12442,N_6014,N_9860);
and U12443 (N_12443,N_8770,N_7361);
nor U12444 (N_12444,N_8674,N_8447);
and U12445 (N_12445,N_6199,N_5583);
nor U12446 (N_12446,N_8877,N_7830);
or U12447 (N_12447,N_6829,N_6236);
xnor U12448 (N_12448,N_8027,N_5544);
nand U12449 (N_12449,N_9005,N_7391);
or U12450 (N_12450,N_8185,N_6549);
or U12451 (N_12451,N_7584,N_6032);
xnor U12452 (N_12452,N_9186,N_8031);
nand U12453 (N_12453,N_8089,N_6860);
and U12454 (N_12454,N_9948,N_9584);
or U12455 (N_12455,N_6511,N_7664);
xnor U12456 (N_12456,N_7609,N_9329);
or U12457 (N_12457,N_7282,N_9742);
nor U12458 (N_12458,N_9664,N_7503);
or U12459 (N_12459,N_7668,N_7032);
and U12460 (N_12460,N_5313,N_6185);
or U12461 (N_12461,N_8261,N_8274);
nor U12462 (N_12462,N_5867,N_7869);
or U12463 (N_12463,N_7805,N_7262);
and U12464 (N_12464,N_5964,N_8581);
nand U12465 (N_12465,N_8439,N_8867);
nand U12466 (N_12466,N_8315,N_5120);
xnor U12467 (N_12467,N_9397,N_9646);
nand U12468 (N_12468,N_5873,N_7292);
and U12469 (N_12469,N_8962,N_7161);
or U12470 (N_12470,N_6189,N_5197);
and U12471 (N_12471,N_7662,N_9066);
or U12472 (N_12472,N_6752,N_7294);
and U12473 (N_12473,N_8686,N_7384);
nor U12474 (N_12474,N_6635,N_6266);
nand U12475 (N_12475,N_9656,N_7952);
or U12476 (N_12476,N_9438,N_5872);
and U12477 (N_12477,N_7062,N_5457);
and U12478 (N_12478,N_6559,N_6102);
or U12479 (N_12479,N_8130,N_6732);
and U12480 (N_12480,N_7608,N_7079);
xnor U12481 (N_12481,N_9769,N_8994);
and U12482 (N_12482,N_9778,N_5038);
nor U12483 (N_12483,N_6490,N_7198);
or U12484 (N_12484,N_6091,N_7827);
xnor U12485 (N_12485,N_5059,N_7627);
nor U12486 (N_12486,N_6572,N_6705);
nand U12487 (N_12487,N_6541,N_7719);
or U12488 (N_12488,N_5416,N_6571);
nor U12489 (N_12489,N_6331,N_5786);
xor U12490 (N_12490,N_8369,N_7480);
xor U12491 (N_12491,N_8335,N_6007);
xor U12492 (N_12492,N_5224,N_8198);
xnor U12493 (N_12493,N_5312,N_8949);
or U12494 (N_12494,N_7674,N_7676);
nor U12495 (N_12495,N_5615,N_6385);
or U12496 (N_12496,N_7841,N_8445);
nor U12497 (N_12497,N_9429,N_9866);
and U12498 (N_12498,N_5169,N_9262);
nand U12499 (N_12499,N_8894,N_9385);
nand U12500 (N_12500,N_7349,N_9636);
or U12501 (N_12501,N_8643,N_6871);
nor U12502 (N_12502,N_9543,N_5379);
and U12503 (N_12503,N_5788,N_9929);
nand U12504 (N_12504,N_6886,N_8808);
or U12505 (N_12505,N_7155,N_9995);
nor U12506 (N_12506,N_8081,N_7322);
or U12507 (N_12507,N_5563,N_9921);
or U12508 (N_12508,N_8650,N_5974);
nand U12509 (N_12509,N_9249,N_9107);
and U12510 (N_12510,N_6463,N_5438);
nand U12511 (N_12511,N_8347,N_9471);
nand U12512 (N_12512,N_5727,N_9509);
and U12513 (N_12513,N_9374,N_6487);
or U12514 (N_12514,N_5501,N_9897);
xnor U12515 (N_12515,N_8919,N_7248);
or U12516 (N_12516,N_8994,N_9160);
and U12517 (N_12517,N_9817,N_9128);
or U12518 (N_12518,N_5837,N_5403);
nand U12519 (N_12519,N_8668,N_8881);
or U12520 (N_12520,N_6649,N_9232);
and U12521 (N_12521,N_9335,N_5746);
and U12522 (N_12522,N_8703,N_6552);
nor U12523 (N_12523,N_5221,N_5095);
and U12524 (N_12524,N_7070,N_5629);
and U12525 (N_12525,N_5430,N_7074);
or U12526 (N_12526,N_7784,N_7593);
xnor U12527 (N_12527,N_6658,N_9937);
nor U12528 (N_12528,N_9578,N_8049);
xor U12529 (N_12529,N_9363,N_5466);
nor U12530 (N_12530,N_7693,N_7868);
and U12531 (N_12531,N_7150,N_7994);
or U12532 (N_12532,N_9800,N_5130);
and U12533 (N_12533,N_5793,N_6471);
nor U12534 (N_12534,N_9753,N_7284);
or U12535 (N_12535,N_9434,N_9802);
nor U12536 (N_12536,N_5155,N_9395);
and U12537 (N_12537,N_8753,N_8146);
and U12538 (N_12538,N_7093,N_7352);
nor U12539 (N_12539,N_8305,N_7193);
xnor U12540 (N_12540,N_9335,N_5515);
and U12541 (N_12541,N_5865,N_9102);
nor U12542 (N_12542,N_8797,N_8314);
nor U12543 (N_12543,N_8471,N_7386);
or U12544 (N_12544,N_7301,N_5582);
nand U12545 (N_12545,N_9214,N_6366);
nand U12546 (N_12546,N_5193,N_5602);
or U12547 (N_12547,N_6053,N_8470);
nand U12548 (N_12548,N_8417,N_8016);
or U12549 (N_12549,N_5972,N_6773);
and U12550 (N_12550,N_5799,N_8023);
nand U12551 (N_12551,N_6064,N_5272);
and U12552 (N_12552,N_6504,N_8321);
and U12553 (N_12553,N_7050,N_5614);
nand U12554 (N_12554,N_7592,N_5666);
and U12555 (N_12555,N_9337,N_5153);
or U12556 (N_12556,N_8867,N_5784);
nand U12557 (N_12557,N_6657,N_6249);
or U12558 (N_12558,N_7529,N_7027);
or U12559 (N_12559,N_7038,N_9860);
and U12560 (N_12560,N_7316,N_9596);
and U12561 (N_12561,N_5886,N_8621);
and U12562 (N_12562,N_6065,N_5856);
nor U12563 (N_12563,N_6339,N_7905);
or U12564 (N_12564,N_7933,N_5000);
or U12565 (N_12565,N_9664,N_7843);
and U12566 (N_12566,N_7628,N_9251);
nor U12567 (N_12567,N_6988,N_9868);
nand U12568 (N_12568,N_6738,N_5343);
nor U12569 (N_12569,N_8793,N_7643);
nand U12570 (N_12570,N_5872,N_5627);
nor U12571 (N_12571,N_8231,N_7452);
nand U12572 (N_12572,N_6756,N_6916);
nand U12573 (N_12573,N_7364,N_7889);
or U12574 (N_12574,N_5904,N_8974);
xnor U12575 (N_12575,N_6377,N_8566);
or U12576 (N_12576,N_7558,N_7092);
nand U12577 (N_12577,N_9409,N_8386);
and U12578 (N_12578,N_5775,N_6048);
and U12579 (N_12579,N_9738,N_5868);
xnor U12580 (N_12580,N_8653,N_5524);
nand U12581 (N_12581,N_6937,N_7047);
nand U12582 (N_12582,N_8268,N_6543);
or U12583 (N_12583,N_5624,N_6548);
nor U12584 (N_12584,N_5134,N_6455);
nand U12585 (N_12585,N_8272,N_6927);
nand U12586 (N_12586,N_8980,N_5630);
nand U12587 (N_12587,N_8255,N_6796);
nand U12588 (N_12588,N_5145,N_7246);
xnor U12589 (N_12589,N_5908,N_5655);
nor U12590 (N_12590,N_8738,N_6041);
nand U12591 (N_12591,N_9097,N_9206);
and U12592 (N_12592,N_6020,N_8660);
nand U12593 (N_12593,N_8525,N_7893);
and U12594 (N_12594,N_6057,N_7629);
xor U12595 (N_12595,N_5230,N_7234);
nor U12596 (N_12596,N_7799,N_5109);
nor U12597 (N_12597,N_5895,N_9185);
xor U12598 (N_12598,N_6036,N_8298);
and U12599 (N_12599,N_9399,N_9915);
nor U12600 (N_12600,N_8876,N_9400);
or U12601 (N_12601,N_8279,N_5886);
nor U12602 (N_12602,N_9730,N_6166);
xnor U12603 (N_12603,N_9253,N_7505);
or U12604 (N_12604,N_5455,N_8862);
or U12605 (N_12605,N_7666,N_6655);
xnor U12606 (N_12606,N_6491,N_5427);
nand U12607 (N_12607,N_5345,N_5795);
and U12608 (N_12608,N_9796,N_5029);
xor U12609 (N_12609,N_8537,N_7512);
xor U12610 (N_12610,N_7340,N_9862);
nor U12611 (N_12611,N_9224,N_7353);
xnor U12612 (N_12612,N_7081,N_6623);
nand U12613 (N_12613,N_5797,N_6680);
or U12614 (N_12614,N_6552,N_8427);
or U12615 (N_12615,N_9932,N_8117);
and U12616 (N_12616,N_7055,N_7463);
xor U12617 (N_12617,N_7995,N_8666);
nor U12618 (N_12618,N_5888,N_9659);
nand U12619 (N_12619,N_9501,N_8607);
and U12620 (N_12620,N_7324,N_8793);
nand U12621 (N_12621,N_5917,N_5083);
nor U12622 (N_12622,N_8287,N_7187);
nand U12623 (N_12623,N_9960,N_8907);
nor U12624 (N_12624,N_7438,N_6086);
and U12625 (N_12625,N_5925,N_5497);
and U12626 (N_12626,N_6289,N_7357);
nand U12627 (N_12627,N_5525,N_9295);
nand U12628 (N_12628,N_6281,N_7768);
nand U12629 (N_12629,N_7667,N_6775);
and U12630 (N_12630,N_7864,N_5440);
or U12631 (N_12631,N_8628,N_7215);
nand U12632 (N_12632,N_7559,N_6172);
or U12633 (N_12633,N_7131,N_7502);
xor U12634 (N_12634,N_7728,N_5930);
nand U12635 (N_12635,N_7586,N_6242);
and U12636 (N_12636,N_5116,N_7647);
nor U12637 (N_12637,N_5769,N_8159);
nor U12638 (N_12638,N_8961,N_9427);
nand U12639 (N_12639,N_6327,N_7171);
and U12640 (N_12640,N_5625,N_6018);
and U12641 (N_12641,N_5232,N_9389);
and U12642 (N_12642,N_6162,N_9257);
and U12643 (N_12643,N_6481,N_5053);
nand U12644 (N_12644,N_9809,N_9261);
and U12645 (N_12645,N_9012,N_6623);
nand U12646 (N_12646,N_5657,N_6131);
nand U12647 (N_12647,N_7883,N_7926);
nor U12648 (N_12648,N_8341,N_6572);
or U12649 (N_12649,N_8710,N_9438);
nand U12650 (N_12650,N_6039,N_5802);
and U12651 (N_12651,N_7776,N_7243);
and U12652 (N_12652,N_9924,N_6349);
nor U12653 (N_12653,N_6233,N_9604);
xnor U12654 (N_12654,N_8667,N_5770);
or U12655 (N_12655,N_9030,N_6412);
nor U12656 (N_12656,N_6684,N_9807);
or U12657 (N_12657,N_7628,N_5706);
nor U12658 (N_12658,N_5061,N_8532);
nor U12659 (N_12659,N_5720,N_8143);
or U12660 (N_12660,N_6791,N_8372);
or U12661 (N_12661,N_9038,N_7714);
nor U12662 (N_12662,N_5611,N_5570);
nor U12663 (N_12663,N_8695,N_7748);
and U12664 (N_12664,N_9008,N_6438);
nor U12665 (N_12665,N_5906,N_5899);
or U12666 (N_12666,N_9881,N_8850);
and U12667 (N_12667,N_5474,N_8832);
or U12668 (N_12668,N_6173,N_9658);
nand U12669 (N_12669,N_5401,N_8977);
nand U12670 (N_12670,N_8652,N_9258);
xnor U12671 (N_12671,N_9168,N_8911);
xnor U12672 (N_12672,N_9302,N_8833);
or U12673 (N_12673,N_5012,N_5536);
or U12674 (N_12674,N_7309,N_9475);
nor U12675 (N_12675,N_9794,N_5597);
and U12676 (N_12676,N_7276,N_8654);
and U12677 (N_12677,N_5156,N_7642);
or U12678 (N_12678,N_6460,N_5251);
or U12679 (N_12679,N_8921,N_5783);
and U12680 (N_12680,N_6881,N_5037);
xnor U12681 (N_12681,N_6622,N_5907);
and U12682 (N_12682,N_9955,N_5831);
nand U12683 (N_12683,N_6504,N_8355);
xnor U12684 (N_12684,N_6771,N_5613);
nand U12685 (N_12685,N_9031,N_7301);
or U12686 (N_12686,N_6649,N_5198);
and U12687 (N_12687,N_9215,N_5390);
xor U12688 (N_12688,N_5546,N_9494);
nor U12689 (N_12689,N_8407,N_7572);
xor U12690 (N_12690,N_5931,N_9580);
and U12691 (N_12691,N_7823,N_6764);
and U12692 (N_12692,N_5886,N_5190);
and U12693 (N_12693,N_7018,N_7681);
nand U12694 (N_12694,N_6758,N_8236);
nand U12695 (N_12695,N_8166,N_9450);
nor U12696 (N_12696,N_6454,N_6523);
or U12697 (N_12697,N_8456,N_8300);
nand U12698 (N_12698,N_5265,N_6633);
or U12699 (N_12699,N_9436,N_5956);
nand U12700 (N_12700,N_6212,N_7246);
and U12701 (N_12701,N_7316,N_6200);
or U12702 (N_12702,N_8373,N_8973);
and U12703 (N_12703,N_8127,N_6239);
nor U12704 (N_12704,N_6439,N_9535);
or U12705 (N_12705,N_9823,N_7405);
or U12706 (N_12706,N_8108,N_5111);
xnor U12707 (N_12707,N_5784,N_8339);
nand U12708 (N_12708,N_6248,N_8859);
nand U12709 (N_12709,N_7539,N_9823);
nor U12710 (N_12710,N_9902,N_5311);
nand U12711 (N_12711,N_7290,N_6270);
and U12712 (N_12712,N_8392,N_5174);
nor U12713 (N_12713,N_6253,N_9431);
or U12714 (N_12714,N_7447,N_8509);
or U12715 (N_12715,N_5474,N_8073);
xor U12716 (N_12716,N_9167,N_8048);
nor U12717 (N_12717,N_8706,N_9337);
nand U12718 (N_12718,N_5954,N_9076);
and U12719 (N_12719,N_9713,N_5238);
nand U12720 (N_12720,N_9880,N_7560);
nand U12721 (N_12721,N_8006,N_6218);
xor U12722 (N_12722,N_9286,N_5387);
and U12723 (N_12723,N_8561,N_7799);
nor U12724 (N_12724,N_5070,N_8869);
or U12725 (N_12725,N_8302,N_8262);
and U12726 (N_12726,N_9508,N_8868);
or U12727 (N_12727,N_8970,N_9696);
nand U12728 (N_12728,N_6766,N_6748);
or U12729 (N_12729,N_9947,N_5828);
nor U12730 (N_12730,N_5581,N_8861);
xor U12731 (N_12731,N_5784,N_6923);
or U12732 (N_12732,N_5586,N_7025);
nand U12733 (N_12733,N_5519,N_5996);
nor U12734 (N_12734,N_9864,N_8009);
or U12735 (N_12735,N_9713,N_8206);
or U12736 (N_12736,N_8146,N_5622);
nor U12737 (N_12737,N_7761,N_6360);
and U12738 (N_12738,N_6454,N_8769);
nor U12739 (N_12739,N_9493,N_5616);
or U12740 (N_12740,N_7414,N_5940);
nand U12741 (N_12741,N_5081,N_7413);
or U12742 (N_12742,N_9610,N_8160);
nand U12743 (N_12743,N_9750,N_6204);
nor U12744 (N_12744,N_5948,N_8199);
nand U12745 (N_12745,N_6688,N_9719);
xnor U12746 (N_12746,N_8928,N_8457);
and U12747 (N_12747,N_5032,N_6492);
nand U12748 (N_12748,N_8040,N_5190);
nand U12749 (N_12749,N_5964,N_5116);
and U12750 (N_12750,N_6052,N_6603);
nor U12751 (N_12751,N_5504,N_6804);
nand U12752 (N_12752,N_7836,N_9911);
nor U12753 (N_12753,N_5415,N_8075);
and U12754 (N_12754,N_7970,N_5027);
and U12755 (N_12755,N_5712,N_8357);
and U12756 (N_12756,N_5912,N_6082);
nor U12757 (N_12757,N_7370,N_7615);
or U12758 (N_12758,N_7878,N_7750);
nand U12759 (N_12759,N_9816,N_7419);
or U12760 (N_12760,N_5235,N_6311);
or U12761 (N_12761,N_8074,N_7059);
or U12762 (N_12762,N_6009,N_7266);
nor U12763 (N_12763,N_7166,N_6151);
and U12764 (N_12764,N_9497,N_8457);
nand U12765 (N_12765,N_6711,N_8422);
nand U12766 (N_12766,N_5360,N_6271);
and U12767 (N_12767,N_8025,N_6199);
or U12768 (N_12768,N_8173,N_7748);
nand U12769 (N_12769,N_9836,N_8753);
or U12770 (N_12770,N_7471,N_8581);
and U12771 (N_12771,N_5682,N_7370);
or U12772 (N_12772,N_5686,N_9900);
nor U12773 (N_12773,N_5770,N_6361);
and U12774 (N_12774,N_7219,N_9591);
nand U12775 (N_12775,N_6476,N_7837);
nor U12776 (N_12776,N_5817,N_6829);
or U12777 (N_12777,N_9229,N_5797);
or U12778 (N_12778,N_9653,N_5378);
nor U12779 (N_12779,N_7392,N_7999);
nand U12780 (N_12780,N_8675,N_8659);
nand U12781 (N_12781,N_5265,N_8190);
nor U12782 (N_12782,N_9678,N_7614);
nand U12783 (N_12783,N_8396,N_5498);
nand U12784 (N_12784,N_6572,N_9721);
and U12785 (N_12785,N_9499,N_5892);
or U12786 (N_12786,N_9400,N_7342);
nor U12787 (N_12787,N_7229,N_8008);
or U12788 (N_12788,N_6778,N_9399);
nor U12789 (N_12789,N_5123,N_5063);
xor U12790 (N_12790,N_8034,N_5793);
nand U12791 (N_12791,N_5066,N_7442);
nor U12792 (N_12792,N_7991,N_9259);
and U12793 (N_12793,N_9706,N_7069);
nand U12794 (N_12794,N_5353,N_9486);
and U12795 (N_12795,N_9705,N_5857);
or U12796 (N_12796,N_8465,N_8929);
nand U12797 (N_12797,N_5275,N_9810);
or U12798 (N_12798,N_5999,N_9930);
or U12799 (N_12799,N_8776,N_5815);
or U12800 (N_12800,N_7807,N_8717);
nand U12801 (N_12801,N_9412,N_8689);
xor U12802 (N_12802,N_8899,N_9581);
nor U12803 (N_12803,N_9354,N_8802);
or U12804 (N_12804,N_7868,N_5419);
nor U12805 (N_12805,N_7138,N_7687);
or U12806 (N_12806,N_6095,N_5585);
nor U12807 (N_12807,N_8344,N_8611);
nand U12808 (N_12808,N_5039,N_5859);
and U12809 (N_12809,N_8146,N_9903);
or U12810 (N_12810,N_7940,N_8763);
nor U12811 (N_12811,N_6822,N_8630);
or U12812 (N_12812,N_7055,N_5744);
nor U12813 (N_12813,N_9900,N_6288);
nor U12814 (N_12814,N_5233,N_5447);
xor U12815 (N_12815,N_7495,N_9226);
nand U12816 (N_12816,N_7074,N_9636);
and U12817 (N_12817,N_7161,N_6045);
and U12818 (N_12818,N_9499,N_6061);
or U12819 (N_12819,N_5480,N_9229);
or U12820 (N_12820,N_6648,N_7501);
and U12821 (N_12821,N_7159,N_7201);
and U12822 (N_12822,N_9309,N_8544);
and U12823 (N_12823,N_9852,N_6843);
or U12824 (N_12824,N_6267,N_6069);
xnor U12825 (N_12825,N_7639,N_5883);
and U12826 (N_12826,N_5108,N_5665);
or U12827 (N_12827,N_7773,N_8199);
and U12828 (N_12828,N_5487,N_7339);
nor U12829 (N_12829,N_5866,N_6396);
nand U12830 (N_12830,N_9773,N_8297);
and U12831 (N_12831,N_8187,N_5549);
or U12832 (N_12832,N_9936,N_6483);
nand U12833 (N_12833,N_8355,N_9380);
or U12834 (N_12834,N_5431,N_9322);
nor U12835 (N_12835,N_7464,N_5731);
or U12836 (N_12836,N_9543,N_5303);
or U12837 (N_12837,N_9144,N_7358);
nand U12838 (N_12838,N_8207,N_6745);
or U12839 (N_12839,N_6369,N_5484);
nor U12840 (N_12840,N_8854,N_9334);
xor U12841 (N_12841,N_6354,N_8922);
nor U12842 (N_12842,N_7556,N_9740);
nor U12843 (N_12843,N_5028,N_7251);
or U12844 (N_12844,N_8573,N_8193);
nor U12845 (N_12845,N_7159,N_8287);
nor U12846 (N_12846,N_7672,N_6286);
xnor U12847 (N_12847,N_7528,N_6733);
and U12848 (N_12848,N_6656,N_7684);
nor U12849 (N_12849,N_8323,N_7797);
nand U12850 (N_12850,N_6808,N_5414);
nand U12851 (N_12851,N_9542,N_6882);
or U12852 (N_12852,N_8905,N_7421);
and U12853 (N_12853,N_7829,N_7406);
and U12854 (N_12854,N_6393,N_6339);
nand U12855 (N_12855,N_5080,N_5157);
and U12856 (N_12856,N_5513,N_9757);
and U12857 (N_12857,N_8172,N_5697);
xor U12858 (N_12858,N_6990,N_5984);
or U12859 (N_12859,N_7628,N_5728);
xnor U12860 (N_12860,N_5376,N_6177);
nor U12861 (N_12861,N_5268,N_9165);
nand U12862 (N_12862,N_6936,N_8209);
or U12863 (N_12863,N_6175,N_6586);
nand U12864 (N_12864,N_9340,N_5240);
nand U12865 (N_12865,N_7819,N_9452);
or U12866 (N_12866,N_8647,N_8311);
and U12867 (N_12867,N_7108,N_7062);
and U12868 (N_12868,N_8748,N_7880);
xnor U12869 (N_12869,N_7394,N_6860);
or U12870 (N_12870,N_8954,N_6144);
nor U12871 (N_12871,N_9558,N_6438);
and U12872 (N_12872,N_8632,N_7677);
xor U12873 (N_12873,N_9541,N_5607);
nand U12874 (N_12874,N_5244,N_6932);
nand U12875 (N_12875,N_9273,N_8791);
nor U12876 (N_12876,N_7558,N_8935);
and U12877 (N_12877,N_8348,N_9600);
or U12878 (N_12878,N_5161,N_6192);
or U12879 (N_12879,N_6952,N_6472);
and U12880 (N_12880,N_7112,N_7717);
and U12881 (N_12881,N_7943,N_8942);
xor U12882 (N_12882,N_9779,N_8883);
or U12883 (N_12883,N_9350,N_6504);
nor U12884 (N_12884,N_5018,N_7987);
or U12885 (N_12885,N_5247,N_6715);
or U12886 (N_12886,N_5675,N_6757);
or U12887 (N_12887,N_6178,N_5320);
and U12888 (N_12888,N_5331,N_6024);
nand U12889 (N_12889,N_7503,N_8892);
nand U12890 (N_12890,N_6236,N_9131);
xnor U12891 (N_12891,N_7048,N_7579);
and U12892 (N_12892,N_5238,N_7008);
or U12893 (N_12893,N_7456,N_7605);
nand U12894 (N_12894,N_6344,N_8996);
nand U12895 (N_12895,N_9879,N_8731);
and U12896 (N_12896,N_9433,N_9717);
and U12897 (N_12897,N_5381,N_9112);
and U12898 (N_12898,N_6209,N_9688);
and U12899 (N_12899,N_7845,N_7326);
or U12900 (N_12900,N_7988,N_7364);
nor U12901 (N_12901,N_5413,N_8917);
nand U12902 (N_12902,N_6059,N_6589);
or U12903 (N_12903,N_8875,N_9299);
or U12904 (N_12904,N_9160,N_5731);
xnor U12905 (N_12905,N_5385,N_8715);
and U12906 (N_12906,N_9172,N_6398);
nand U12907 (N_12907,N_8362,N_5830);
and U12908 (N_12908,N_7695,N_8592);
or U12909 (N_12909,N_6991,N_9974);
and U12910 (N_12910,N_8300,N_8141);
or U12911 (N_12911,N_5251,N_5170);
nor U12912 (N_12912,N_6040,N_6471);
nand U12913 (N_12913,N_6415,N_5104);
and U12914 (N_12914,N_8573,N_8181);
nand U12915 (N_12915,N_9585,N_8521);
and U12916 (N_12916,N_9990,N_6624);
or U12917 (N_12917,N_5091,N_5207);
nand U12918 (N_12918,N_5944,N_9111);
or U12919 (N_12919,N_9194,N_7814);
or U12920 (N_12920,N_5807,N_5911);
and U12921 (N_12921,N_6123,N_5903);
nor U12922 (N_12922,N_9262,N_6193);
or U12923 (N_12923,N_5965,N_9228);
and U12924 (N_12924,N_7881,N_5964);
or U12925 (N_12925,N_7362,N_9395);
nand U12926 (N_12926,N_6215,N_6171);
nor U12927 (N_12927,N_8919,N_6431);
and U12928 (N_12928,N_8795,N_6531);
or U12929 (N_12929,N_6377,N_8876);
and U12930 (N_12930,N_9653,N_5942);
or U12931 (N_12931,N_8468,N_8121);
nand U12932 (N_12932,N_9228,N_8322);
nor U12933 (N_12933,N_6542,N_5278);
nor U12934 (N_12934,N_7640,N_9605);
and U12935 (N_12935,N_6393,N_9505);
and U12936 (N_12936,N_8826,N_8985);
nor U12937 (N_12937,N_7739,N_8789);
and U12938 (N_12938,N_5784,N_8981);
or U12939 (N_12939,N_6193,N_6759);
or U12940 (N_12940,N_6994,N_5249);
xnor U12941 (N_12941,N_8344,N_5681);
xor U12942 (N_12942,N_9361,N_7392);
and U12943 (N_12943,N_5211,N_5986);
and U12944 (N_12944,N_9534,N_6401);
nor U12945 (N_12945,N_8050,N_7483);
or U12946 (N_12946,N_5995,N_9317);
nor U12947 (N_12947,N_6256,N_7121);
nand U12948 (N_12948,N_8481,N_6382);
or U12949 (N_12949,N_6302,N_5873);
nand U12950 (N_12950,N_8930,N_6467);
and U12951 (N_12951,N_8138,N_7588);
nand U12952 (N_12952,N_5518,N_9926);
and U12953 (N_12953,N_8193,N_9702);
and U12954 (N_12954,N_9043,N_6708);
or U12955 (N_12955,N_5800,N_5937);
nand U12956 (N_12956,N_7108,N_5866);
nand U12957 (N_12957,N_6755,N_5461);
xor U12958 (N_12958,N_5687,N_7049);
or U12959 (N_12959,N_7096,N_9658);
nor U12960 (N_12960,N_7976,N_5745);
nor U12961 (N_12961,N_9294,N_7197);
xor U12962 (N_12962,N_5657,N_5136);
or U12963 (N_12963,N_8965,N_5995);
and U12964 (N_12964,N_9713,N_5597);
or U12965 (N_12965,N_9747,N_6545);
or U12966 (N_12966,N_9818,N_9880);
or U12967 (N_12967,N_7181,N_9823);
and U12968 (N_12968,N_6033,N_9696);
and U12969 (N_12969,N_5962,N_5284);
nor U12970 (N_12970,N_9532,N_7246);
and U12971 (N_12971,N_7706,N_7082);
and U12972 (N_12972,N_6745,N_6024);
or U12973 (N_12973,N_8174,N_8407);
or U12974 (N_12974,N_5704,N_9114);
nor U12975 (N_12975,N_8216,N_9139);
or U12976 (N_12976,N_6463,N_9817);
or U12977 (N_12977,N_6973,N_7444);
xor U12978 (N_12978,N_9814,N_7414);
and U12979 (N_12979,N_9248,N_5157);
nor U12980 (N_12980,N_6905,N_9660);
and U12981 (N_12981,N_8857,N_8135);
or U12982 (N_12982,N_9304,N_7694);
and U12983 (N_12983,N_5943,N_8065);
xnor U12984 (N_12984,N_8521,N_8171);
nor U12985 (N_12985,N_8803,N_7724);
and U12986 (N_12986,N_7953,N_9984);
nand U12987 (N_12987,N_7135,N_9032);
xnor U12988 (N_12988,N_6253,N_9410);
nor U12989 (N_12989,N_9994,N_9220);
nor U12990 (N_12990,N_7172,N_6134);
and U12991 (N_12991,N_5356,N_5928);
nand U12992 (N_12992,N_6031,N_6228);
or U12993 (N_12993,N_9890,N_9744);
nand U12994 (N_12994,N_8356,N_5796);
nor U12995 (N_12995,N_5588,N_6332);
nand U12996 (N_12996,N_5174,N_5346);
nor U12997 (N_12997,N_7489,N_8499);
and U12998 (N_12998,N_9922,N_8336);
and U12999 (N_12999,N_9723,N_7036);
and U13000 (N_13000,N_8452,N_7369);
nand U13001 (N_13001,N_9322,N_7033);
xnor U13002 (N_13002,N_7268,N_8864);
xnor U13003 (N_13003,N_8568,N_8769);
nor U13004 (N_13004,N_7574,N_6244);
nor U13005 (N_13005,N_8669,N_7108);
and U13006 (N_13006,N_5066,N_5737);
or U13007 (N_13007,N_5474,N_5195);
nand U13008 (N_13008,N_6779,N_9793);
or U13009 (N_13009,N_7288,N_9235);
nor U13010 (N_13010,N_5730,N_6780);
nor U13011 (N_13011,N_6118,N_8503);
and U13012 (N_13012,N_8141,N_7728);
or U13013 (N_13013,N_5003,N_6758);
nand U13014 (N_13014,N_9612,N_6529);
nor U13015 (N_13015,N_9934,N_9961);
or U13016 (N_13016,N_7197,N_8212);
and U13017 (N_13017,N_7334,N_8134);
or U13018 (N_13018,N_8188,N_9740);
nand U13019 (N_13019,N_8893,N_7427);
nor U13020 (N_13020,N_8245,N_7546);
and U13021 (N_13021,N_8541,N_9519);
nor U13022 (N_13022,N_5896,N_9027);
nor U13023 (N_13023,N_8887,N_7215);
nand U13024 (N_13024,N_8263,N_6381);
and U13025 (N_13025,N_6576,N_5079);
or U13026 (N_13026,N_5715,N_9967);
and U13027 (N_13027,N_7643,N_8507);
nand U13028 (N_13028,N_5553,N_5521);
and U13029 (N_13029,N_6692,N_7863);
and U13030 (N_13030,N_9233,N_9666);
nand U13031 (N_13031,N_8126,N_7755);
nand U13032 (N_13032,N_7566,N_8724);
or U13033 (N_13033,N_6224,N_8830);
and U13034 (N_13034,N_6715,N_5861);
nor U13035 (N_13035,N_5577,N_8350);
xor U13036 (N_13036,N_6643,N_7065);
and U13037 (N_13037,N_7688,N_7129);
or U13038 (N_13038,N_6148,N_5896);
nor U13039 (N_13039,N_6440,N_6599);
and U13040 (N_13040,N_9635,N_6064);
xnor U13041 (N_13041,N_5492,N_8822);
nand U13042 (N_13042,N_9631,N_7826);
nor U13043 (N_13043,N_9748,N_7546);
or U13044 (N_13044,N_5620,N_7376);
nor U13045 (N_13045,N_8596,N_9738);
and U13046 (N_13046,N_8757,N_5387);
and U13047 (N_13047,N_7029,N_9823);
xnor U13048 (N_13048,N_7626,N_7356);
nand U13049 (N_13049,N_9335,N_5883);
nand U13050 (N_13050,N_5298,N_8376);
nand U13051 (N_13051,N_5691,N_9724);
nand U13052 (N_13052,N_5828,N_7694);
and U13053 (N_13053,N_9100,N_8834);
xnor U13054 (N_13054,N_9122,N_5164);
xnor U13055 (N_13055,N_8640,N_7120);
nand U13056 (N_13056,N_9204,N_5069);
xor U13057 (N_13057,N_7191,N_8952);
nand U13058 (N_13058,N_8842,N_6761);
and U13059 (N_13059,N_5620,N_8159);
and U13060 (N_13060,N_7156,N_8154);
or U13061 (N_13061,N_7516,N_8639);
nor U13062 (N_13062,N_5932,N_8137);
xnor U13063 (N_13063,N_5863,N_5024);
nand U13064 (N_13064,N_7254,N_5354);
or U13065 (N_13065,N_6436,N_8974);
nor U13066 (N_13066,N_7223,N_9320);
or U13067 (N_13067,N_5106,N_9872);
xnor U13068 (N_13068,N_9867,N_5641);
nor U13069 (N_13069,N_5938,N_7120);
nor U13070 (N_13070,N_5331,N_6131);
or U13071 (N_13071,N_5791,N_8364);
xor U13072 (N_13072,N_8140,N_9606);
nand U13073 (N_13073,N_7561,N_7351);
nand U13074 (N_13074,N_6049,N_6838);
or U13075 (N_13075,N_9703,N_7723);
and U13076 (N_13076,N_5163,N_8086);
nor U13077 (N_13077,N_7110,N_9381);
nand U13078 (N_13078,N_6232,N_6052);
or U13079 (N_13079,N_5806,N_5018);
or U13080 (N_13080,N_8720,N_6943);
nor U13081 (N_13081,N_9186,N_6719);
and U13082 (N_13082,N_8434,N_8236);
xor U13083 (N_13083,N_6725,N_7235);
nor U13084 (N_13084,N_7006,N_6558);
nand U13085 (N_13085,N_6321,N_8392);
or U13086 (N_13086,N_9123,N_8851);
nor U13087 (N_13087,N_8489,N_5125);
or U13088 (N_13088,N_7757,N_5703);
and U13089 (N_13089,N_6855,N_8427);
nor U13090 (N_13090,N_8782,N_6245);
nand U13091 (N_13091,N_9668,N_7556);
nand U13092 (N_13092,N_7627,N_5038);
nand U13093 (N_13093,N_7845,N_7706);
nand U13094 (N_13094,N_7408,N_6947);
or U13095 (N_13095,N_9443,N_6054);
nor U13096 (N_13096,N_7264,N_6502);
and U13097 (N_13097,N_9929,N_6066);
nand U13098 (N_13098,N_9067,N_8587);
xnor U13099 (N_13099,N_9060,N_7504);
xor U13100 (N_13100,N_8665,N_7928);
nand U13101 (N_13101,N_9456,N_8271);
nor U13102 (N_13102,N_6355,N_6224);
xor U13103 (N_13103,N_6253,N_9052);
or U13104 (N_13104,N_6730,N_7797);
xnor U13105 (N_13105,N_6885,N_6591);
xnor U13106 (N_13106,N_9383,N_8442);
nor U13107 (N_13107,N_8091,N_9815);
and U13108 (N_13108,N_9978,N_5591);
nor U13109 (N_13109,N_6677,N_8668);
or U13110 (N_13110,N_7646,N_5049);
or U13111 (N_13111,N_7073,N_5225);
nor U13112 (N_13112,N_7271,N_6089);
nor U13113 (N_13113,N_8255,N_7652);
nand U13114 (N_13114,N_6670,N_8615);
nand U13115 (N_13115,N_8314,N_7416);
or U13116 (N_13116,N_9968,N_5327);
and U13117 (N_13117,N_6206,N_9315);
nor U13118 (N_13118,N_6617,N_6333);
nor U13119 (N_13119,N_5516,N_6164);
xor U13120 (N_13120,N_7347,N_6122);
xnor U13121 (N_13121,N_7922,N_6139);
and U13122 (N_13122,N_9477,N_9279);
nand U13123 (N_13123,N_8647,N_9946);
and U13124 (N_13124,N_9332,N_7062);
nor U13125 (N_13125,N_7435,N_6593);
xor U13126 (N_13126,N_8753,N_7117);
and U13127 (N_13127,N_8769,N_5445);
nand U13128 (N_13128,N_9323,N_9599);
and U13129 (N_13129,N_9035,N_7069);
or U13130 (N_13130,N_7418,N_5200);
nor U13131 (N_13131,N_9119,N_7013);
nor U13132 (N_13132,N_9573,N_8378);
nor U13133 (N_13133,N_6660,N_6860);
or U13134 (N_13134,N_9675,N_7254);
or U13135 (N_13135,N_7447,N_6080);
xnor U13136 (N_13136,N_8658,N_5856);
nor U13137 (N_13137,N_9382,N_6366);
xnor U13138 (N_13138,N_6263,N_6247);
or U13139 (N_13139,N_6788,N_5758);
or U13140 (N_13140,N_6672,N_7246);
or U13141 (N_13141,N_9685,N_9852);
nand U13142 (N_13142,N_9353,N_9925);
and U13143 (N_13143,N_6060,N_8205);
and U13144 (N_13144,N_5484,N_6084);
nand U13145 (N_13145,N_6113,N_9574);
xor U13146 (N_13146,N_9551,N_9990);
nand U13147 (N_13147,N_9914,N_5405);
or U13148 (N_13148,N_5470,N_6762);
nand U13149 (N_13149,N_6140,N_5004);
nand U13150 (N_13150,N_7842,N_7671);
nor U13151 (N_13151,N_9501,N_8914);
nand U13152 (N_13152,N_6647,N_6145);
nor U13153 (N_13153,N_7983,N_6021);
xor U13154 (N_13154,N_6315,N_5241);
nand U13155 (N_13155,N_5244,N_6234);
nor U13156 (N_13156,N_8518,N_8672);
or U13157 (N_13157,N_7051,N_9958);
nand U13158 (N_13158,N_8018,N_7370);
xnor U13159 (N_13159,N_6791,N_9457);
nand U13160 (N_13160,N_9292,N_7059);
or U13161 (N_13161,N_8277,N_5286);
nor U13162 (N_13162,N_5198,N_9246);
or U13163 (N_13163,N_7911,N_9398);
and U13164 (N_13164,N_7001,N_7005);
or U13165 (N_13165,N_8731,N_5598);
or U13166 (N_13166,N_8787,N_7630);
nor U13167 (N_13167,N_5193,N_6316);
nand U13168 (N_13168,N_9518,N_8919);
nor U13169 (N_13169,N_8019,N_5603);
and U13170 (N_13170,N_8275,N_8538);
nor U13171 (N_13171,N_9926,N_8063);
nand U13172 (N_13172,N_7761,N_6309);
or U13173 (N_13173,N_6288,N_9451);
nor U13174 (N_13174,N_5062,N_9313);
and U13175 (N_13175,N_7957,N_5849);
nor U13176 (N_13176,N_9897,N_8792);
or U13177 (N_13177,N_5092,N_8296);
and U13178 (N_13178,N_7081,N_5094);
nor U13179 (N_13179,N_9281,N_5764);
nand U13180 (N_13180,N_7074,N_8125);
nand U13181 (N_13181,N_8589,N_6965);
nor U13182 (N_13182,N_9342,N_9774);
nand U13183 (N_13183,N_9947,N_5573);
nor U13184 (N_13184,N_5918,N_6095);
and U13185 (N_13185,N_5648,N_6359);
or U13186 (N_13186,N_9064,N_8143);
nand U13187 (N_13187,N_8070,N_7414);
or U13188 (N_13188,N_6100,N_6530);
and U13189 (N_13189,N_9237,N_8191);
nor U13190 (N_13190,N_6857,N_6957);
or U13191 (N_13191,N_8786,N_6266);
nand U13192 (N_13192,N_9789,N_6545);
or U13193 (N_13193,N_8971,N_6340);
nand U13194 (N_13194,N_5384,N_8273);
and U13195 (N_13195,N_8433,N_9564);
nand U13196 (N_13196,N_5977,N_6239);
nand U13197 (N_13197,N_8237,N_6021);
and U13198 (N_13198,N_8952,N_9389);
nand U13199 (N_13199,N_9257,N_9834);
nor U13200 (N_13200,N_6121,N_7876);
nor U13201 (N_13201,N_7849,N_9275);
nand U13202 (N_13202,N_8744,N_5084);
nor U13203 (N_13203,N_8739,N_9157);
nor U13204 (N_13204,N_8656,N_5934);
nand U13205 (N_13205,N_7772,N_5870);
or U13206 (N_13206,N_8633,N_9980);
or U13207 (N_13207,N_9691,N_5072);
or U13208 (N_13208,N_9229,N_8089);
xor U13209 (N_13209,N_7648,N_9170);
and U13210 (N_13210,N_8552,N_5606);
nand U13211 (N_13211,N_8372,N_6501);
or U13212 (N_13212,N_7301,N_6107);
nor U13213 (N_13213,N_7602,N_8602);
nor U13214 (N_13214,N_7653,N_7000);
nor U13215 (N_13215,N_9630,N_7812);
or U13216 (N_13216,N_9542,N_9876);
or U13217 (N_13217,N_9627,N_9620);
or U13218 (N_13218,N_5647,N_8554);
xor U13219 (N_13219,N_8381,N_8080);
nand U13220 (N_13220,N_5624,N_9511);
and U13221 (N_13221,N_5536,N_6714);
and U13222 (N_13222,N_6481,N_6880);
nor U13223 (N_13223,N_9323,N_9479);
or U13224 (N_13224,N_6570,N_8905);
and U13225 (N_13225,N_8629,N_7956);
or U13226 (N_13226,N_8948,N_8771);
and U13227 (N_13227,N_8468,N_7144);
nand U13228 (N_13228,N_6850,N_8882);
or U13229 (N_13229,N_6757,N_6562);
and U13230 (N_13230,N_6694,N_8623);
and U13231 (N_13231,N_5508,N_9086);
nand U13232 (N_13232,N_9746,N_8220);
and U13233 (N_13233,N_6644,N_8148);
xor U13234 (N_13234,N_8126,N_9064);
and U13235 (N_13235,N_9054,N_6582);
or U13236 (N_13236,N_6027,N_7627);
and U13237 (N_13237,N_7315,N_7393);
nor U13238 (N_13238,N_8773,N_6542);
nand U13239 (N_13239,N_9626,N_7496);
nand U13240 (N_13240,N_5150,N_8197);
nand U13241 (N_13241,N_7938,N_9379);
and U13242 (N_13242,N_6893,N_5608);
or U13243 (N_13243,N_6648,N_6338);
and U13244 (N_13244,N_6165,N_8457);
nor U13245 (N_13245,N_6029,N_8214);
and U13246 (N_13246,N_9263,N_9008);
nor U13247 (N_13247,N_6466,N_7920);
nand U13248 (N_13248,N_7848,N_8080);
nand U13249 (N_13249,N_9711,N_8887);
and U13250 (N_13250,N_7036,N_7328);
and U13251 (N_13251,N_6438,N_9516);
nand U13252 (N_13252,N_7732,N_5506);
and U13253 (N_13253,N_6338,N_7943);
and U13254 (N_13254,N_7885,N_5523);
or U13255 (N_13255,N_7522,N_7662);
and U13256 (N_13256,N_7991,N_8608);
or U13257 (N_13257,N_5566,N_9073);
and U13258 (N_13258,N_8046,N_8862);
nand U13259 (N_13259,N_6484,N_6502);
nand U13260 (N_13260,N_5715,N_9543);
or U13261 (N_13261,N_8797,N_9592);
and U13262 (N_13262,N_5451,N_6902);
and U13263 (N_13263,N_8258,N_8150);
and U13264 (N_13264,N_6946,N_6692);
and U13265 (N_13265,N_5253,N_5756);
nor U13266 (N_13266,N_6581,N_5460);
and U13267 (N_13267,N_8800,N_8865);
nand U13268 (N_13268,N_6193,N_7414);
nor U13269 (N_13269,N_5599,N_9292);
or U13270 (N_13270,N_5938,N_5044);
nand U13271 (N_13271,N_5407,N_7385);
and U13272 (N_13272,N_5221,N_6888);
nand U13273 (N_13273,N_6395,N_5583);
nand U13274 (N_13274,N_6829,N_5377);
xnor U13275 (N_13275,N_6326,N_6224);
and U13276 (N_13276,N_9503,N_7840);
and U13277 (N_13277,N_8028,N_5110);
nand U13278 (N_13278,N_8938,N_9325);
nand U13279 (N_13279,N_7605,N_8621);
nand U13280 (N_13280,N_7907,N_6069);
nor U13281 (N_13281,N_9286,N_9938);
nor U13282 (N_13282,N_7301,N_8312);
nor U13283 (N_13283,N_5578,N_6726);
or U13284 (N_13284,N_9967,N_6083);
nor U13285 (N_13285,N_9661,N_6297);
nor U13286 (N_13286,N_7844,N_8892);
or U13287 (N_13287,N_7487,N_5446);
nand U13288 (N_13288,N_6629,N_6873);
xnor U13289 (N_13289,N_6789,N_7634);
xor U13290 (N_13290,N_7773,N_8480);
and U13291 (N_13291,N_6269,N_7337);
and U13292 (N_13292,N_6316,N_5340);
and U13293 (N_13293,N_9038,N_8499);
xor U13294 (N_13294,N_9727,N_8148);
nor U13295 (N_13295,N_6755,N_7228);
or U13296 (N_13296,N_6193,N_6644);
or U13297 (N_13297,N_7773,N_8078);
xor U13298 (N_13298,N_5786,N_6803);
nand U13299 (N_13299,N_9802,N_6104);
and U13300 (N_13300,N_8146,N_7932);
and U13301 (N_13301,N_5484,N_5247);
or U13302 (N_13302,N_6940,N_7212);
nand U13303 (N_13303,N_6848,N_5971);
or U13304 (N_13304,N_8174,N_9626);
and U13305 (N_13305,N_8620,N_9470);
nor U13306 (N_13306,N_6321,N_5014);
xor U13307 (N_13307,N_5299,N_9965);
or U13308 (N_13308,N_8318,N_9372);
xor U13309 (N_13309,N_6007,N_7930);
or U13310 (N_13310,N_7354,N_7615);
nand U13311 (N_13311,N_8093,N_9645);
or U13312 (N_13312,N_5435,N_9288);
or U13313 (N_13313,N_9639,N_6176);
or U13314 (N_13314,N_5318,N_9292);
nor U13315 (N_13315,N_5692,N_8370);
or U13316 (N_13316,N_9078,N_9019);
or U13317 (N_13317,N_7659,N_5136);
and U13318 (N_13318,N_8449,N_5383);
or U13319 (N_13319,N_8021,N_6266);
nand U13320 (N_13320,N_6014,N_8498);
nor U13321 (N_13321,N_9398,N_7567);
nand U13322 (N_13322,N_9677,N_7580);
and U13323 (N_13323,N_7199,N_6143);
nand U13324 (N_13324,N_8704,N_8458);
or U13325 (N_13325,N_5567,N_6798);
or U13326 (N_13326,N_6549,N_9340);
and U13327 (N_13327,N_8020,N_5734);
nor U13328 (N_13328,N_6054,N_8268);
nand U13329 (N_13329,N_6901,N_6117);
nand U13330 (N_13330,N_5624,N_6058);
or U13331 (N_13331,N_7734,N_9554);
nor U13332 (N_13332,N_8935,N_8445);
nand U13333 (N_13333,N_7509,N_8746);
and U13334 (N_13334,N_5599,N_9884);
nand U13335 (N_13335,N_9868,N_6848);
nor U13336 (N_13336,N_9792,N_6014);
nand U13337 (N_13337,N_7313,N_9733);
and U13338 (N_13338,N_5747,N_6831);
nor U13339 (N_13339,N_7197,N_5803);
or U13340 (N_13340,N_9993,N_6209);
nor U13341 (N_13341,N_6548,N_7755);
nor U13342 (N_13342,N_8536,N_7252);
nand U13343 (N_13343,N_5553,N_5322);
nor U13344 (N_13344,N_7386,N_8617);
or U13345 (N_13345,N_5865,N_9381);
nor U13346 (N_13346,N_8251,N_9869);
and U13347 (N_13347,N_6173,N_9886);
and U13348 (N_13348,N_9775,N_5593);
or U13349 (N_13349,N_8854,N_8755);
xnor U13350 (N_13350,N_5215,N_9529);
and U13351 (N_13351,N_8204,N_9671);
nand U13352 (N_13352,N_6398,N_8355);
and U13353 (N_13353,N_5892,N_5412);
nor U13354 (N_13354,N_7501,N_6509);
nor U13355 (N_13355,N_5656,N_8485);
and U13356 (N_13356,N_9679,N_7471);
nand U13357 (N_13357,N_7034,N_7565);
nor U13358 (N_13358,N_5625,N_9291);
or U13359 (N_13359,N_9119,N_9363);
and U13360 (N_13360,N_7284,N_7014);
nand U13361 (N_13361,N_6940,N_8825);
or U13362 (N_13362,N_9754,N_8591);
nand U13363 (N_13363,N_6020,N_8270);
or U13364 (N_13364,N_8253,N_8136);
or U13365 (N_13365,N_8328,N_9128);
or U13366 (N_13366,N_6175,N_7107);
nor U13367 (N_13367,N_6200,N_9585);
nor U13368 (N_13368,N_8131,N_7008);
and U13369 (N_13369,N_9138,N_9609);
nor U13370 (N_13370,N_9582,N_6943);
nor U13371 (N_13371,N_9021,N_9551);
or U13372 (N_13372,N_9291,N_5632);
or U13373 (N_13373,N_9191,N_7029);
xor U13374 (N_13374,N_9776,N_9399);
nor U13375 (N_13375,N_5151,N_5420);
nor U13376 (N_13376,N_6087,N_5328);
or U13377 (N_13377,N_7200,N_6451);
nor U13378 (N_13378,N_6103,N_6499);
and U13379 (N_13379,N_7738,N_9472);
nor U13380 (N_13380,N_7760,N_8356);
or U13381 (N_13381,N_9927,N_6630);
and U13382 (N_13382,N_9293,N_7063);
nor U13383 (N_13383,N_5831,N_5655);
nor U13384 (N_13384,N_7142,N_5010);
or U13385 (N_13385,N_5197,N_7693);
nor U13386 (N_13386,N_8135,N_5552);
or U13387 (N_13387,N_8084,N_9720);
nand U13388 (N_13388,N_7928,N_7366);
xor U13389 (N_13389,N_6035,N_5398);
nor U13390 (N_13390,N_9351,N_5800);
xnor U13391 (N_13391,N_9112,N_8182);
nand U13392 (N_13392,N_9378,N_6175);
nor U13393 (N_13393,N_8340,N_9777);
and U13394 (N_13394,N_7572,N_8707);
or U13395 (N_13395,N_9978,N_9778);
nand U13396 (N_13396,N_6513,N_8305);
or U13397 (N_13397,N_8369,N_9030);
and U13398 (N_13398,N_8806,N_5812);
and U13399 (N_13399,N_7710,N_8224);
nor U13400 (N_13400,N_8733,N_9537);
nor U13401 (N_13401,N_9279,N_8958);
nor U13402 (N_13402,N_8779,N_5100);
nor U13403 (N_13403,N_8170,N_5896);
xor U13404 (N_13404,N_6557,N_9515);
or U13405 (N_13405,N_9216,N_7754);
xnor U13406 (N_13406,N_6273,N_5640);
nor U13407 (N_13407,N_6058,N_6325);
nor U13408 (N_13408,N_7756,N_5792);
nor U13409 (N_13409,N_5347,N_6833);
or U13410 (N_13410,N_8857,N_5499);
nand U13411 (N_13411,N_5877,N_8737);
nor U13412 (N_13412,N_6451,N_9123);
or U13413 (N_13413,N_7885,N_8549);
and U13414 (N_13414,N_6636,N_5256);
nand U13415 (N_13415,N_9766,N_5441);
nand U13416 (N_13416,N_6889,N_8872);
or U13417 (N_13417,N_7604,N_7075);
nor U13418 (N_13418,N_6489,N_6207);
nor U13419 (N_13419,N_9314,N_9615);
or U13420 (N_13420,N_7266,N_7839);
nand U13421 (N_13421,N_9628,N_9750);
nor U13422 (N_13422,N_5802,N_7512);
xor U13423 (N_13423,N_5332,N_7027);
nand U13424 (N_13424,N_6169,N_8474);
nand U13425 (N_13425,N_8094,N_6847);
nand U13426 (N_13426,N_8660,N_8481);
xor U13427 (N_13427,N_5106,N_6111);
or U13428 (N_13428,N_5458,N_6353);
xor U13429 (N_13429,N_9886,N_6440);
and U13430 (N_13430,N_8357,N_5867);
nand U13431 (N_13431,N_7816,N_9880);
nand U13432 (N_13432,N_9846,N_7994);
or U13433 (N_13433,N_8775,N_6072);
or U13434 (N_13434,N_7908,N_8235);
nor U13435 (N_13435,N_6725,N_9453);
and U13436 (N_13436,N_9887,N_5364);
nor U13437 (N_13437,N_9878,N_6446);
and U13438 (N_13438,N_5951,N_5752);
or U13439 (N_13439,N_5255,N_8685);
nor U13440 (N_13440,N_6078,N_9297);
nor U13441 (N_13441,N_7770,N_5723);
and U13442 (N_13442,N_6381,N_7969);
nor U13443 (N_13443,N_8984,N_9749);
nand U13444 (N_13444,N_9328,N_5446);
and U13445 (N_13445,N_7553,N_5221);
and U13446 (N_13446,N_6760,N_7893);
nor U13447 (N_13447,N_8193,N_9910);
and U13448 (N_13448,N_6094,N_6607);
and U13449 (N_13449,N_8962,N_7944);
or U13450 (N_13450,N_7388,N_6679);
or U13451 (N_13451,N_7871,N_5191);
nor U13452 (N_13452,N_7079,N_5250);
and U13453 (N_13453,N_9325,N_9765);
nor U13454 (N_13454,N_7367,N_5442);
or U13455 (N_13455,N_5157,N_9416);
nor U13456 (N_13456,N_8344,N_6155);
and U13457 (N_13457,N_7769,N_6073);
or U13458 (N_13458,N_9425,N_7057);
xnor U13459 (N_13459,N_8025,N_8183);
xor U13460 (N_13460,N_6409,N_9677);
nor U13461 (N_13461,N_5788,N_5640);
or U13462 (N_13462,N_6878,N_9434);
and U13463 (N_13463,N_9460,N_8466);
or U13464 (N_13464,N_9915,N_6106);
nand U13465 (N_13465,N_6499,N_6754);
and U13466 (N_13466,N_7545,N_7449);
xnor U13467 (N_13467,N_9084,N_8673);
and U13468 (N_13468,N_5490,N_5369);
and U13469 (N_13469,N_7556,N_7600);
xnor U13470 (N_13470,N_8092,N_9597);
or U13471 (N_13471,N_8690,N_8095);
nand U13472 (N_13472,N_6000,N_6208);
nor U13473 (N_13473,N_5636,N_7374);
and U13474 (N_13474,N_6117,N_8566);
xnor U13475 (N_13475,N_9330,N_8627);
and U13476 (N_13476,N_9231,N_7690);
xnor U13477 (N_13477,N_9384,N_8408);
or U13478 (N_13478,N_6955,N_6322);
and U13479 (N_13479,N_9818,N_6022);
nor U13480 (N_13480,N_6745,N_7837);
and U13481 (N_13481,N_7676,N_7748);
or U13482 (N_13482,N_6280,N_9983);
xor U13483 (N_13483,N_9401,N_5475);
nand U13484 (N_13484,N_5478,N_9871);
nand U13485 (N_13485,N_6589,N_5822);
nor U13486 (N_13486,N_5845,N_7541);
or U13487 (N_13487,N_8160,N_5486);
nand U13488 (N_13488,N_8099,N_8191);
xnor U13489 (N_13489,N_6711,N_7700);
nand U13490 (N_13490,N_9068,N_5442);
or U13491 (N_13491,N_9788,N_9900);
xor U13492 (N_13492,N_5237,N_5033);
or U13493 (N_13493,N_6243,N_6649);
nor U13494 (N_13494,N_7789,N_9485);
nor U13495 (N_13495,N_5601,N_9177);
or U13496 (N_13496,N_5529,N_8243);
and U13497 (N_13497,N_9053,N_6903);
or U13498 (N_13498,N_8628,N_6168);
nor U13499 (N_13499,N_5742,N_9387);
nor U13500 (N_13500,N_9807,N_7811);
and U13501 (N_13501,N_5519,N_6370);
or U13502 (N_13502,N_9942,N_6082);
nand U13503 (N_13503,N_9625,N_7256);
or U13504 (N_13504,N_6597,N_8705);
nand U13505 (N_13505,N_7657,N_5222);
and U13506 (N_13506,N_5411,N_9497);
nand U13507 (N_13507,N_9547,N_6009);
and U13508 (N_13508,N_5660,N_7392);
nand U13509 (N_13509,N_8771,N_8995);
and U13510 (N_13510,N_9176,N_9600);
and U13511 (N_13511,N_8406,N_8669);
or U13512 (N_13512,N_8491,N_9329);
or U13513 (N_13513,N_5918,N_6082);
xor U13514 (N_13514,N_7637,N_8453);
nand U13515 (N_13515,N_5240,N_7364);
or U13516 (N_13516,N_8325,N_7516);
or U13517 (N_13517,N_6142,N_9379);
xor U13518 (N_13518,N_5026,N_9628);
nor U13519 (N_13519,N_9408,N_7075);
and U13520 (N_13520,N_7239,N_5255);
and U13521 (N_13521,N_5468,N_6973);
nand U13522 (N_13522,N_8687,N_6671);
or U13523 (N_13523,N_5459,N_9221);
or U13524 (N_13524,N_6245,N_6269);
nor U13525 (N_13525,N_8769,N_6614);
nand U13526 (N_13526,N_6806,N_6317);
and U13527 (N_13527,N_9081,N_7225);
or U13528 (N_13528,N_8570,N_9942);
nor U13529 (N_13529,N_5991,N_6829);
nand U13530 (N_13530,N_5530,N_6473);
nor U13531 (N_13531,N_9993,N_9218);
or U13532 (N_13532,N_5830,N_8497);
or U13533 (N_13533,N_9467,N_8436);
and U13534 (N_13534,N_8561,N_9350);
or U13535 (N_13535,N_5570,N_7096);
nand U13536 (N_13536,N_7438,N_9895);
nor U13537 (N_13537,N_9644,N_8483);
and U13538 (N_13538,N_6151,N_5821);
or U13539 (N_13539,N_7647,N_9915);
or U13540 (N_13540,N_5355,N_8485);
nor U13541 (N_13541,N_7706,N_6303);
and U13542 (N_13542,N_8723,N_9000);
xor U13543 (N_13543,N_9144,N_9506);
nand U13544 (N_13544,N_5246,N_7769);
nor U13545 (N_13545,N_8886,N_7827);
xor U13546 (N_13546,N_6926,N_8159);
nor U13547 (N_13547,N_8300,N_6858);
and U13548 (N_13548,N_7564,N_8730);
and U13549 (N_13549,N_8571,N_6106);
and U13550 (N_13550,N_8998,N_8877);
or U13551 (N_13551,N_6072,N_5806);
nand U13552 (N_13552,N_6994,N_5937);
or U13553 (N_13553,N_9066,N_9512);
nor U13554 (N_13554,N_8502,N_8860);
nor U13555 (N_13555,N_7273,N_6897);
or U13556 (N_13556,N_6350,N_8031);
nand U13557 (N_13557,N_7861,N_7549);
xnor U13558 (N_13558,N_7582,N_6750);
nand U13559 (N_13559,N_5614,N_9233);
and U13560 (N_13560,N_8267,N_7974);
and U13561 (N_13561,N_8623,N_8641);
nor U13562 (N_13562,N_7998,N_8657);
xor U13563 (N_13563,N_7168,N_7768);
nand U13564 (N_13564,N_7056,N_9628);
or U13565 (N_13565,N_5260,N_7733);
and U13566 (N_13566,N_5717,N_9456);
nand U13567 (N_13567,N_5584,N_9712);
or U13568 (N_13568,N_8781,N_5198);
nand U13569 (N_13569,N_7836,N_5905);
or U13570 (N_13570,N_5511,N_6405);
nand U13571 (N_13571,N_8650,N_9025);
or U13572 (N_13572,N_7584,N_8197);
nor U13573 (N_13573,N_5997,N_8350);
nor U13574 (N_13574,N_6966,N_5080);
or U13575 (N_13575,N_6726,N_5928);
and U13576 (N_13576,N_9190,N_8116);
nand U13577 (N_13577,N_8964,N_7471);
xor U13578 (N_13578,N_5262,N_9006);
nor U13579 (N_13579,N_5586,N_8777);
xnor U13580 (N_13580,N_8122,N_7892);
nor U13581 (N_13581,N_8092,N_8087);
or U13582 (N_13582,N_5377,N_8700);
or U13583 (N_13583,N_7717,N_8552);
and U13584 (N_13584,N_9746,N_5117);
nand U13585 (N_13585,N_9991,N_6017);
nand U13586 (N_13586,N_9675,N_8180);
and U13587 (N_13587,N_9220,N_5591);
or U13588 (N_13588,N_6981,N_5236);
or U13589 (N_13589,N_6887,N_6484);
or U13590 (N_13590,N_8014,N_8158);
nor U13591 (N_13591,N_5199,N_9609);
xnor U13592 (N_13592,N_5218,N_6174);
nor U13593 (N_13593,N_5130,N_9640);
and U13594 (N_13594,N_5510,N_5503);
nor U13595 (N_13595,N_5222,N_5006);
nor U13596 (N_13596,N_7094,N_8838);
nor U13597 (N_13597,N_8678,N_6437);
and U13598 (N_13598,N_7802,N_9900);
nor U13599 (N_13599,N_5666,N_9142);
nand U13600 (N_13600,N_5305,N_8468);
or U13601 (N_13601,N_7230,N_6912);
nand U13602 (N_13602,N_9857,N_7149);
or U13603 (N_13603,N_9827,N_5685);
nor U13604 (N_13604,N_5694,N_6884);
nand U13605 (N_13605,N_6871,N_7925);
nand U13606 (N_13606,N_5301,N_7693);
or U13607 (N_13607,N_5608,N_5492);
nor U13608 (N_13608,N_8769,N_9498);
or U13609 (N_13609,N_5272,N_6058);
nor U13610 (N_13610,N_6484,N_5040);
and U13611 (N_13611,N_8501,N_7546);
or U13612 (N_13612,N_7591,N_7202);
nand U13613 (N_13613,N_8418,N_9841);
nand U13614 (N_13614,N_7613,N_6588);
nor U13615 (N_13615,N_5457,N_6366);
and U13616 (N_13616,N_7828,N_8459);
nand U13617 (N_13617,N_5284,N_7903);
nand U13618 (N_13618,N_5607,N_9623);
and U13619 (N_13619,N_9286,N_5504);
and U13620 (N_13620,N_8370,N_6773);
or U13621 (N_13621,N_6619,N_8525);
nand U13622 (N_13622,N_5880,N_8776);
nand U13623 (N_13623,N_8232,N_6901);
or U13624 (N_13624,N_6306,N_7096);
and U13625 (N_13625,N_7543,N_5512);
or U13626 (N_13626,N_9162,N_5567);
xnor U13627 (N_13627,N_8660,N_7544);
or U13628 (N_13628,N_7216,N_7321);
and U13629 (N_13629,N_6891,N_5221);
and U13630 (N_13630,N_8890,N_5800);
xor U13631 (N_13631,N_6890,N_6430);
and U13632 (N_13632,N_9610,N_8417);
nor U13633 (N_13633,N_7126,N_5649);
nor U13634 (N_13634,N_8401,N_8993);
and U13635 (N_13635,N_9033,N_6685);
nand U13636 (N_13636,N_8918,N_5454);
or U13637 (N_13637,N_7393,N_9432);
nand U13638 (N_13638,N_6689,N_6787);
or U13639 (N_13639,N_9469,N_5447);
nor U13640 (N_13640,N_8897,N_9012);
and U13641 (N_13641,N_5002,N_6847);
or U13642 (N_13642,N_9744,N_8663);
nand U13643 (N_13643,N_9235,N_9806);
nor U13644 (N_13644,N_7816,N_5190);
nand U13645 (N_13645,N_9279,N_5136);
xnor U13646 (N_13646,N_6934,N_8719);
or U13647 (N_13647,N_9160,N_7322);
nand U13648 (N_13648,N_8278,N_6913);
nand U13649 (N_13649,N_7028,N_5377);
nor U13650 (N_13650,N_7218,N_8244);
or U13651 (N_13651,N_9090,N_6788);
nor U13652 (N_13652,N_8011,N_5046);
or U13653 (N_13653,N_9806,N_7803);
and U13654 (N_13654,N_8097,N_9544);
nand U13655 (N_13655,N_8626,N_8276);
nor U13656 (N_13656,N_9549,N_8649);
or U13657 (N_13657,N_5242,N_6659);
or U13658 (N_13658,N_8194,N_8455);
and U13659 (N_13659,N_7856,N_7756);
and U13660 (N_13660,N_6759,N_9559);
nand U13661 (N_13661,N_9234,N_6026);
nor U13662 (N_13662,N_9122,N_9591);
and U13663 (N_13663,N_9044,N_7600);
nor U13664 (N_13664,N_9747,N_5365);
and U13665 (N_13665,N_5477,N_9648);
xnor U13666 (N_13666,N_9894,N_9182);
nor U13667 (N_13667,N_9917,N_6424);
nor U13668 (N_13668,N_6362,N_7068);
nor U13669 (N_13669,N_8102,N_8558);
nand U13670 (N_13670,N_8198,N_8380);
or U13671 (N_13671,N_7949,N_5361);
nor U13672 (N_13672,N_6902,N_6637);
nand U13673 (N_13673,N_6620,N_9058);
and U13674 (N_13674,N_9524,N_6396);
and U13675 (N_13675,N_9798,N_5066);
or U13676 (N_13676,N_5861,N_5410);
and U13677 (N_13677,N_9543,N_6294);
or U13678 (N_13678,N_9365,N_5935);
or U13679 (N_13679,N_7223,N_5318);
nor U13680 (N_13680,N_5913,N_5827);
xor U13681 (N_13681,N_8674,N_7918);
and U13682 (N_13682,N_5757,N_7715);
xnor U13683 (N_13683,N_7562,N_7360);
nor U13684 (N_13684,N_6377,N_9351);
nor U13685 (N_13685,N_7938,N_7397);
xnor U13686 (N_13686,N_6985,N_9228);
nand U13687 (N_13687,N_7569,N_6996);
nand U13688 (N_13688,N_7281,N_7613);
nor U13689 (N_13689,N_9000,N_5564);
and U13690 (N_13690,N_6389,N_7401);
xor U13691 (N_13691,N_5279,N_8418);
nand U13692 (N_13692,N_6808,N_9476);
and U13693 (N_13693,N_9422,N_9072);
nand U13694 (N_13694,N_7753,N_9692);
xnor U13695 (N_13695,N_8882,N_7023);
xnor U13696 (N_13696,N_5553,N_8517);
nor U13697 (N_13697,N_9170,N_9005);
and U13698 (N_13698,N_9569,N_9761);
xnor U13699 (N_13699,N_6048,N_5688);
nand U13700 (N_13700,N_8356,N_6204);
nand U13701 (N_13701,N_8048,N_5867);
nand U13702 (N_13702,N_5107,N_9941);
or U13703 (N_13703,N_9289,N_9752);
nor U13704 (N_13704,N_6953,N_7370);
nor U13705 (N_13705,N_7494,N_9655);
and U13706 (N_13706,N_8777,N_9519);
nor U13707 (N_13707,N_5281,N_7653);
nand U13708 (N_13708,N_9500,N_9932);
or U13709 (N_13709,N_6526,N_5602);
nor U13710 (N_13710,N_9055,N_7571);
and U13711 (N_13711,N_7315,N_9247);
and U13712 (N_13712,N_5616,N_8002);
or U13713 (N_13713,N_7793,N_9300);
nand U13714 (N_13714,N_5562,N_6798);
and U13715 (N_13715,N_5314,N_7764);
nand U13716 (N_13716,N_5776,N_6605);
or U13717 (N_13717,N_8868,N_6331);
nand U13718 (N_13718,N_8558,N_9527);
xor U13719 (N_13719,N_8154,N_8336);
or U13720 (N_13720,N_9708,N_8296);
nor U13721 (N_13721,N_7617,N_5570);
or U13722 (N_13722,N_7308,N_7248);
and U13723 (N_13723,N_8127,N_6644);
nor U13724 (N_13724,N_9366,N_7455);
nand U13725 (N_13725,N_7565,N_9205);
and U13726 (N_13726,N_5635,N_8769);
nand U13727 (N_13727,N_9000,N_9882);
or U13728 (N_13728,N_8324,N_6549);
nor U13729 (N_13729,N_5075,N_8450);
nor U13730 (N_13730,N_5642,N_8482);
nand U13731 (N_13731,N_8270,N_9694);
nand U13732 (N_13732,N_6928,N_6380);
or U13733 (N_13733,N_8239,N_7144);
nand U13734 (N_13734,N_7191,N_9791);
or U13735 (N_13735,N_5176,N_7647);
or U13736 (N_13736,N_8319,N_9368);
or U13737 (N_13737,N_9384,N_6726);
and U13738 (N_13738,N_9991,N_5804);
nor U13739 (N_13739,N_5138,N_6104);
or U13740 (N_13740,N_7500,N_9807);
nand U13741 (N_13741,N_5827,N_6791);
or U13742 (N_13742,N_7481,N_6189);
nand U13743 (N_13743,N_7276,N_5560);
and U13744 (N_13744,N_5868,N_9332);
or U13745 (N_13745,N_9831,N_6697);
nand U13746 (N_13746,N_6076,N_8764);
or U13747 (N_13747,N_8115,N_5306);
xor U13748 (N_13748,N_5509,N_5856);
or U13749 (N_13749,N_7825,N_9004);
or U13750 (N_13750,N_5542,N_5341);
or U13751 (N_13751,N_5433,N_8225);
nand U13752 (N_13752,N_5385,N_8428);
nand U13753 (N_13753,N_6061,N_7625);
nor U13754 (N_13754,N_9524,N_9860);
nor U13755 (N_13755,N_5803,N_6169);
nand U13756 (N_13756,N_9793,N_5899);
xor U13757 (N_13757,N_9004,N_7904);
nor U13758 (N_13758,N_9401,N_5253);
and U13759 (N_13759,N_5647,N_5976);
nor U13760 (N_13760,N_7640,N_6156);
and U13761 (N_13761,N_6005,N_6573);
or U13762 (N_13762,N_9236,N_8414);
or U13763 (N_13763,N_7933,N_6961);
nor U13764 (N_13764,N_7204,N_6857);
nand U13765 (N_13765,N_5734,N_9723);
nor U13766 (N_13766,N_5572,N_5831);
nor U13767 (N_13767,N_9696,N_9900);
nand U13768 (N_13768,N_9730,N_8098);
nor U13769 (N_13769,N_9755,N_5354);
nand U13770 (N_13770,N_8171,N_6147);
or U13771 (N_13771,N_5783,N_5907);
xor U13772 (N_13772,N_5468,N_9700);
and U13773 (N_13773,N_6087,N_5266);
nand U13774 (N_13774,N_8487,N_7482);
or U13775 (N_13775,N_8106,N_5515);
and U13776 (N_13776,N_7534,N_7823);
xnor U13777 (N_13777,N_5320,N_9142);
nand U13778 (N_13778,N_9926,N_9614);
and U13779 (N_13779,N_7854,N_7198);
nand U13780 (N_13780,N_8790,N_5853);
or U13781 (N_13781,N_5752,N_5799);
or U13782 (N_13782,N_9516,N_5935);
nor U13783 (N_13783,N_7814,N_7642);
and U13784 (N_13784,N_9093,N_9351);
nor U13785 (N_13785,N_8761,N_6761);
and U13786 (N_13786,N_8595,N_5286);
xnor U13787 (N_13787,N_8867,N_9429);
or U13788 (N_13788,N_9052,N_6757);
or U13789 (N_13789,N_8779,N_7417);
or U13790 (N_13790,N_9778,N_5745);
nor U13791 (N_13791,N_7466,N_5521);
and U13792 (N_13792,N_6999,N_8263);
xor U13793 (N_13793,N_9011,N_8055);
xor U13794 (N_13794,N_9228,N_9909);
nor U13795 (N_13795,N_5307,N_7711);
nor U13796 (N_13796,N_6461,N_6354);
nor U13797 (N_13797,N_7840,N_9882);
and U13798 (N_13798,N_8716,N_9940);
nand U13799 (N_13799,N_8784,N_6577);
and U13800 (N_13800,N_9120,N_5235);
nand U13801 (N_13801,N_8597,N_7789);
or U13802 (N_13802,N_8155,N_7324);
nor U13803 (N_13803,N_7955,N_6759);
and U13804 (N_13804,N_5575,N_8311);
or U13805 (N_13805,N_5911,N_8549);
or U13806 (N_13806,N_7085,N_9444);
nor U13807 (N_13807,N_5024,N_6444);
or U13808 (N_13808,N_7725,N_9320);
and U13809 (N_13809,N_8813,N_5809);
or U13810 (N_13810,N_7571,N_6789);
nor U13811 (N_13811,N_6507,N_7599);
nand U13812 (N_13812,N_8695,N_6442);
or U13813 (N_13813,N_6976,N_5756);
or U13814 (N_13814,N_9170,N_9550);
nand U13815 (N_13815,N_9145,N_5468);
nor U13816 (N_13816,N_7282,N_9131);
or U13817 (N_13817,N_9487,N_9204);
xor U13818 (N_13818,N_6887,N_6676);
nor U13819 (N_13819,N_9169,N_9767);
and U13820 (N_13820,N_7587,N_5959);
and U13821 (N_13821,N_8355,N_8675);
or U13822 (N_13822,N_7246,N_9044);
and U13823 (N_13823,N_5773,N_9364);
or U13824 (N_13824,N_7143,N_8385);
nand U13825 (N_13825,N_9014,N_5860);
xor U13826 (N_13826,N_5703,N_5733);
nand U13827 (N_13827,N_9842,N_6287);
nand U13828 (N_13828,N_5134,N_7264);
nor U13829 (N_13829,N_6569,N_7246);
and U13830 (N_13830,N_9213,N_8710);
and U13831 (N_13831,N_5799,N_7334);
and U13832 (N_13832,N_9396,N_8351);
xor U13833 (N_13833,N_5827,N_8013);
xor U13834 (N_13834,N_8483,N_5100);
nor U13835 (N_13835,N_8727,N_7758);
or U13836 (N_13836,N_5677,N_7603);
nor U13837 (N_13837,N_7848,N_7975);
nor U13838 (N_13838,N_6223,N_7887);
and U13839 (N_13839,N_9985,N_7279);
nand U13840 (N_13840,N_5125,N_8032);
nor U13841 (N_13841,N_9065,N_8612);
nor U13842 (N_13842,N_8089,N_8040);
and U13843 (N_13843,N_6983,N_7020);
nor U13844 (N_13844,N_7634,N_9834);
xor U13845 (N_13845,N_8111,N_7904);
nor U13846 (N_13846,N_7361,N_8839);
xnor U13847 (N_13847,N_9684,N_6139);
nand U13848 (N_13848,N_7700,N_7522);
and U13849 (N_13849,N_6905,N_7277);
and U13850 (N_13850,N_5088,N_6524);
nor U13851 (N_13851,N_5944,N_7391);
or U13852 (N_13852,N_6557,N_9338);
xor U13853 (N_13853,N_9794,N_7919);
and U13854 (N_13854,N_6198,N_7401);
nand U13855 (N_13855,N_8381,N_6556);
and U13856 (N_13856,N_6175,N_9843);
nand U13857 (N_13857,N_8535,N_7921);
and U13858 (N_13858,N_8265,N_8280);
or U13859 (N_13859,N_8765,N_9962);
nor U13860 (N_13860,N_7080,N_8884);
nand U13861 (N_13861,N_5237,N_8288);
nor U13862 (N_13862,N_6772,N_9084);
or U13863 (N_13863,N_8558,N_7612);
nor U13864 (N_13864,N_6734,N_5384);
nor U13865 (N_13865,N_9711,N_5341);
and U13866 (N_13866,N_5070,N_6481);
xnor U13867 (N_13867,N_5232,N_7921);
nor U13868 (N_13868,N_9872,N_9544);
and U13869 (N_13869,N_5443,N_8276);
nand U13870 (N_13870,N_7757,N_9868);
nand U13871 (N_13871,N_8205,N_6370);
nor U13872 (N_13872,N_9861,N_9532);
nand U13873 (N_13873,N_7259,N_5362);
and U13874 (N_13874,N_8249,N_6635);
or U13875 (N_13875,N_9840,N_9571);
nand U13876 (N_13876,N_8889,N_6746);
or U13877 (N_13877,N_8390,N_5954);
and U13878 (N_13878,N_5608,N_7394);
or U13879 (N_13879,N_7254,N_6499);
or U13880 (N_13880,N_5247,N_6161);
nor U13881 (N_13881,N_7598,N_9362);
or U13882 (N_13882,N_8113,N_9867);
and U13883 (N_13883,N_8314,N_5038);
or U13884 (N_13884,N_9438,N_9920);
or U13885 (N_13885,N_5750,N_9451);
xor U13886 (N_13886,N_7846,N_8702);
and U13887 (N_13887,N_6883,N_7562);
and U13888 (N_13888,N_9598,N_9384);
nand U13889 (N_13889,N_7846,N_8800);
nor U13890 (N_13890,N_7145,N_7674);
and U13891 (N_13891,N_6130,N_5926);
nor U13892 (N_13892,N_6254,N_7748);
or U13893 (N_13893,N_7959,N_5418);
or U13894 (N_13894,N_7453,N_6067);
or U13895 (N_13895,N_6418,N_8712);
nor U13896 (N_13896,N_6681,N_8274);
xnor U13897 (N_13897,N_6180,N_6461);
or U13898 (N_13898,N_8579,N_7771);
nand U13899 (N_13899,N_6180,N_5453);
or U13900 (N_13900,N_7180,N_9806);
and U13901 (N_13901,N_8552,N_7278);
or U13902 (N_13902,N_9403,N_5909);
nor U13903 (N_13903,N_5379,N_6951);
nor U13904 (N_13904,N_9638,N_5421);
and U13905 (N_13905,N_5027,N_8428);
or U13906 (N_13906,N_6891,N_7402);
or U13907 (N_13907,N_5018,N_9081);
or U13908 (N_13908,N_6803,N_9094);
nor U13909 (N_13909,N_6340,N_8732);
nor U13910 (N_13910,N_5657,N_8200);
and U13911 (N_13911,N_8933,N_8428);
nor U13912 (N_13912,N_5862,N_7509);
nand U13913 (N_13913,N_6483,N_6584);
nand U13914 (N_13914,N_9562,N_7225);
or U13915 (N_13915,N_8714,N_5859);
or U13916 (N_13916,N_8761,N_8896);
and U13917 (N_13917,N_9827,N_9385);
and U13918 (N_13918,N_6979,N_6881);
or U13919 (N_13919,N_8472,N_5340);
or U13920 (N_13920,N_5698,N_6709);
or U13921 (N_13921,N_8692,N_9305);
nor U13922 (N_13922,N_7150,N_9162);
nand U13923 (N_13923,N_6894,N_7237);
nor U13924 (N_13924,N_8212,N_9026);
and U13925 (N_13925,N_7959,N_5705);
or U13926 (N_13926,N_7701,N_6423);
or U13927 (N_13927,N_8414,N_8572);
nor U13928 (N_13928,N_8996,N_9289);
or U13929 (N_13929,N_5837,N_5336);
nand U13930 (N_13930,N_8586,N_8967);
nor U13931 (N_13931,N_9643,N_5764);
or U13932 (N_13932,N_8098,N_5862);
xnor U13933 (N_13933,N_7942,N_5017);
nor U13934 (N_13934,N_5969,N_5374);
nor U13935 (N_13935,N_5654,N_7933);
nand U13936 (N_13936,N_8883,N_5190);
nand U13937 (N_13937,N_8857,N_6464);
and U13938 (N_13938,N_9803,N_6621);
or U13939 (N_13939,N_5400,N_5728);
nor U13940 (N_13940,N_8546,N_9171);
or U13941 (N_13941,N_5497,N_6968);
nor U13942 (N_13942,N_8443,N_9055);
or U13943 (N_13943,N_8022,N_9532);
or U13944 (N_13944,N_7398,N_9748);
and U13945 (N_13945,N_9671,N_5389);
nand U13946 (N_13946,N_8012,N_9816);
nor U13947 (N_13947,N_9459,N_5441);
and U13948 (N_13948,N_7234,N_7724);
and U13949 (N_13949,N_9528,N_8037);
nor U13950 (N_13950,N_6097,N_8867);
nor U13951 (N_13951,N_7729,N_5759);
nor U13952 (N_13952,N_5441,N_5067);
nor U13953 (N_13953,N_5879,N_6488);
or U13954 (N_13954,N_9262,N_8336);
nand U13955 (N_13955,N_6219,N_5093);
nor U13956 (N_13956,N_9479,N_5044);
nand U13957 (N_13957,N_9224,N_8064);
and U13958 (N_13958,N_8565,N_9041);
xnor U13959 (N_13959,N_6394,N_6656);
and U13960 (N_13960,N_9455,N_7271);
or U13961 (N_13961,N_9963,N_7060);
or U13962 (N_13962,N_9900,N_9633);
or U13963 (N_13963,N_8960,N_8897);
nand U13964 (N_13964,N_9678,N_9711);
or U13965 (N_13965,N_9389,N_5345);
nor U13966 (N_13966,N_5473,N_8440);
and U13967 (N_13967,N_9155,N_5360);
nand U13968 (N_13968,N_9886,N_5448);
xor U13969 (N_13969,N_7666,N_5499);
xor U13970 (N_13970,N_7593,N_6624);
and U13971 (N_13971,N_5021,N_7340);
and U13972 (N_13972,N_7152,N_8670);
or U13973 (N_13973,N_8099,N_9200);
nor U13974 (N_13974,N_8785,N_7599);
and U13975 (N_13975,N_9839,N_8616);
nor U13976 (N_13976,N_9132,N_5350);
or U13977 (N_13977,N_6906,N_9818);
or U13978 (N_13978,N_7019,N_6367);
and U13979 (N_13979,N_9610,N_9854);
and U13980 (N_13980,N_7085,N_9359);
or U13981 (N_13981,N_6074,N_8917);
or U13982 (N_13982,N_8612,N_6560);
xnor U13983 (N_13983,N_5025,N_9901);
nor U13984 (N_13984,N_5649,N_7198);
and U13985 (N_13985,N_7664,N_8262);
or U13986 (N_13986,N_7624,N_6150);
xor U13987 (N_13987,N_8121,N_5051);
nand U13988 (N_13988,N_6918,N_5896);
nor U13989 (N_13989,N_6257,N_9521);
nor U13990 (N_13990,N_8929,N_6707);
nand U13991 (N_13991,N_9240,N_7337);
xor U13992 (N_13992,N_9875,N_8609);
or U13993 (N_13993,N_6715,N_9148);
and U13994 (N_13994,N_5885,N_7900);
and U13995 (N_13995,N_7504,N_5555);
and U13996 (N_13996,N_9351,N_7371);
nor U13997 (N_13997,N_9584,N_7023);
nand U13998 (N_13998,N_9154,N_7904);
xor U13999 (N_13999,N_8146,N_8013);
nand U14000 (N_14000,N_5571,N_6168);
nor U14001 (N_14001,N_6916,N_9172);
and U14002 (N_14002,N_5005,N_7084);
nor U14003 (N_14003,N_9395,N_9467);
or U14004 (N_14004,N_5956,N_5422);
or U14005 (N_14005,N_9786,N_8476);
nand U14006 (N_14006,N_5089,N_9360);
nand U14007 (N_14007,N_6206,N_9062);
nand U14008 (N_14008,N_7473,N_9731);
and U14009 (N_14009,N_5218,N_9227);
xor U14010 (N_14010,N_6767,N_7373);
xnor U14011 (N_14011,N_5765,N_6831);
nand U14012 (N_14012,N_5740,N_7449);
nand U14013 (N_14013,N_6152,N_5792);
xnor U14014 (N_14014,N_6522,N_6727);
nand U14015 (N_14015,N_7080,N_8719);
xnor U14016 (N_14016,N_5017,N_5554);
nand U14017 (N_14017,N_7127,N_9699);
xnor U14018 (N_14018,N_8524,N_7414);
and U14019 (N_14019,N_8997,N_5340);
and U14020 (N_14020,N_6734,N_6003);
or U14021 (N_14021,N_6118,N_5861);
and U14022 (N_14022,N_8062,N_8488);
or U14023 (N_14023,N_9383,N_5032);
nand U14024 (N_14024,N_9346,N_8379);
nor U14025 (N_14025,N_6426,N_6456);
nand U14026 (N_14026,N_8294,N_9503);
and U14027 (N_14027,N_7353,N_8692);
and U14028 (N_14028,N_5694,N_8635);
or U14029 (N_14029,N_6347,N_8411);
and U14030 (N_14030,N_8715,N_7257);
and U14031 (N_14031,N_5234,N_5034);
nand U14032 (N_14032,N_8426,N_7854);
and U14033 (N_14033,N_9280,N_9443);
nor U14034 (N_14034,N_9991,N_8447);
nor U14035 (N_14035,N_7010,N_6847);
nor U14036 (N_14036,N_5541,N_5615);
and U14037 (N_14037,N_7797,N_6411);
and U14038 (N_14038,N_9004,N_9891);
and U14039 (N_14039,N_7148,N_5804);
nand U14040 (N_14040,N_6647,N_5830);
or U14041 (N_14041,N_6758,N_9015);
and U14042 (N_14042,N_7625,N_5912);
and U14043 (N_14043,N_7765,N_5257);
and U14044 (N_14044,N_8532,N_9676);
nor U14045 (N_14045,N_9489,N_6122);
or U14046 (N_14046,N_8063,N_9344);
or U14047 (N_14047,N_6190,N_6815);
or U14048 (N_14048,N_8309,N_6872);
nor U14049 (N_14049,N_9441,N_5142);
or U14050 (N_14050,N_7723,N_9891);
xor U14051 (N_14051,N_7818,N_8390);
xnor U14052 (N_14052,N_9670,N_6598);
or U14053 (N_14053,N_5579,N_8631);
nor U14054 (N_14054,N_5657,N_9786);
and U14055 (N_14055,N_9547,N_5732);
nand U14056 (N_14056,N_8411,N_9058);
or U14057 (N_14057,N_9305,N_6399);
and U14058 (N_14058,N_6170,N_7895);
and U14059 (N_14059,N_5351,N_7651);
or U14060 (N_14060,N_7928,N_5246);
nor U14061 (N_14061,N_5305,N_5093);
nor U14062 (N_14062,N_8728,N_6546);
nand U14063 (N_14063,N_7186,N_6321);
nand U14064 (N_14064,N_9893,N_6120);
nor U14065 (N_14065,N_6440,N_6628);
xor U14066 (N_14066,N_6724,N_8169);
nor U14067 (N_14067,N_5583,N_6908);
and U14068 (N_14068,N_7347,N_6831);
xor U14069 (N_14069,N_6931,N_6036);
or U14070 (N_14070,N_5354,N_7370);
nor U14071 (N_14071,N_8722,N_7340);
nand U14072 (N_14072,N_6560,N_5457);
nor U14073 (N_14073,N_5944,N_5129);
nand U14074 (N_14074,N_7058,N_6403);
and U14075 (N_14075,N_8599,N_7292);
nor U14076 (N_14076,N_6562,N_5359);
nand U14077 (N_14077,N_7953,N_9152);
or U14078 (N_14078,N_5165,N_6439);
and U14079 (N_14079,N_5792,N_8425);
nand U14080 (N_14080,N_6759,N_5140);
nor U14081 (N_14081,N_8398,N_5681);
xnor U14082 (N_14082,N_9705,N_6635);
nor U14083 (N_14083,N_7771,N_8412);
nand U14084 (N_14084,N_6904,N_6542);
and U14085 (N_14085,N_5886,N_8420);
nor U14086 (N_14086,N_7933,N_5674);
nor U14087 (N_14087,N_8787,N_8760);
or U14088 (N_14088,N_5119,N_5919);
nand U14089 (N_14089,N_7163,N_5327);
nand U14090 (N_14090,N_6849,N_6635);
and U14091 (N_14091,N_7074,N_7733);
and U14092 (N_14092,N_9769,N_6579);
nor U14093 (N_14093,N_5793,N_7850);
nand U14094 (N_14094,N_7007,N_5930);
nor U14095 (N_14095,N_7749,N_5010);
nor U14096 (N_14096,N_9747,N_8687);
and U14097 (N_14097,N_7444,N_8592);
nand U14098 (N_14098,N_6093,N_7157);
or U14099 (N_14099,N_8336,N_8606);
nand U14100 (N_14100,N_9693,N_6622);
nand U14101 (N_14101,N_7671,N_9829);
or U14102 (N_14102,N_8693,N_6581);
nand U14103 (N_14103,N_7443,N_7028);
nand U14104 (N_14104,N_5538,N_6348);
nor U14105 (N_14105,N_9650,N_9048);
nor U14106 (N_14106,N_9853,N_8917);
and U14107 (N_14107,N_8021,N_8336);
and U14108 (N_14108,N_5442,N_8854);
nand U14109 (N_14109,N_9766,N_8751);
or U14110 (N_14110,N_9150,N_6112);
nor U14111 (N_14111,N_8601,N_7559);
nor U14112 (N_14112,N_7056,N_9831);
xnor U14113 (N_14113,N_6782,N_5089);
nor U14114 (N_14114,N_6064,N_9811);
nor U14115 (N_14115,N_9749,N_8978);
nand U14116 (N_14116,N_6932,N_7156);
and U14117 (N_14117,N_9181,N_5560);
nand U14118 (N_14118,N_8315,N_7278);
and U14119 (N_14119,N_6964,N_6882);
xnor U14120 (N_14120,N_6653,N_8869);
and U14121 (N_14121,N_7940,N_8842);
nand U14122 (N_14122,N_6396,N_8539);
and U14123 (N_14123,N_5524,N_6769);
nor U14124 (N_14124,N_5064,N_9052);
nand U14125 (N_14125,N_5558,N_8051);
xor U14126 (N_14126,N_7484,N_8419);
nor U14127 (N_14127,N_6231,N_9204);
or U14128 (N_14128,N_7025,N_8375);
and U14129 (N_14129,N_7197,N_9501);
and U14130 (N_14130,N_9602,N_9331);
nand U14131 (N_14131,N_9947,N_5947);
or U14132 (N_14132,N_7102,N_6711);
nor U14133 (N_14133,N_7701,N_5257);
and U14134 (N_14134,N_8756,N_5846);
nand U14135 (N_14135,N_8390,N_9223);
or U14136 (N_14136,N_7431,N_8528);
nor U14137 (N_14137,N_5867,N_5949);
nor U14138 (N_14138,N_8890,N_9504);
or U14139 (N_14139,N_5869,N_7005);
nand U14140 (N_14140,N_5729,N_5366);
or U14141 (N_14141,N_6510,N_9156);
nand U14142 (N_14142,N_7844,N_6029);
xor U14143 (N_14143,N_6598,N_5456);
or U14144 (N_14144,N_6921,N_8749);
nand U14145 (N_14145,N_8651,N_5235);
and U14146 (N_14146,N_7999,N_6294);
nand U14147 (N_14147,N_7849,N_8479);
or U14148 (N_14148,N_8394,N_6307);
nand U14149 (N_14149,N_6928,N_8188);
or U14150 (N_14150,N_6952,N_8745);
or U14151 (N_14151,N_7802,N_6371);
nor U14152 (N_14152,N_6584,N_8594);
nand U14153 (N_14153,N_8725,N_8866);
nand U14154 (N_14154,N_8220,N_7573);
and U14155 (N_14155,N_9034,N_8568);
xor U14156 (N_14156,N_6937,N_5245);
nand U14157 (N_14157,N_8601,N_7675);
or U14158 (N_14158,N_5953,N_5382);
nor U14159 (N_14159,N_8534,N_6515);
nand U14160 (N_14160,N_9572,N_8635);
nor U14161 (N_14161,N_7833,N_5093);
nand U14162 (N_14162,N_7069,N_6209);
nand U14163 (N_14163,N_8129,N_6379);
or U14164 (N_14164,N_5003,N_5804);
nor U14165 (N_14165,N_6546,N_8312);
or U14166 (N_14166,N_7510,N_6289);
nor U14167 (N_14167,N_5562,N_6305);
nand U14168 (N_14168,N_8430,N_7643);
or U14169 (N_14169,N_7377,N_7682);
nor U14170 (N_14170,N_6265,N_5214);
or U14171 (N_14171,N_7880,N_9462);
or U14172 (N_14172,N_5714,N_8847);
nor U14173 (N_14173,N_7064,N_7329);
or U14174 (N_14174,N_8876,N_7027);
and U14175 (N_14175,N_6360,N_9355);
or U14176 (N_14176,N_5220,N_5389);
nor U14177 (N_14177,N_7912,N_7056);
xor U14178 (N_14178,N_7293,N_8089);
nand U14179 (N_14179,N_6847,N_8534);
and U14180 (N_14180,N_9849,N_5217);
xnor U14181 (N_14181,N_6394,N_6171);
or U14182 (N_14182,N_9431,N_7036);
and U14183 (N_14183,N_9692,N_7309);
nand U14184 (N_14184,N_9925,N_7408);
nand U14185 (N_14185,N_7504,N_9537);
xor U14186 (N_14186,N_9423,N_9233);
nor U14187 (N_14187,N_6238,N_9182);
or U14188 (N_14188,N_9223,N_5829);
and U14189 (N_14189,N_5677,N_9599);
and U14190 (N_14190,N_9708,N_7982);
nor U14191 (N_14191,N_7850,N_5899);
nor U14192 (N_14192,N_6297,N_5906);
or U14193 (N_14193,N_9607,N_5907);
or U14194 (N_14194,N_6978,N_8257);
nand U14195 (N_14195,N_9371,N_6008);
or U14196 (N_14196,N_6321,N_5974);
nand U14197 (N_14197,N_5613,N_6172);
and U14198 (N_14198,N_6352,N_5487);
nor U14199 (N_14199,N_7774,N_9620);
nand U14200 (N_14200,N_6460,N_6730);
or U14201 (N_14201,N_9908,N_6281);
nand U14202 (N_14202,N_5524,N_6997);
nand U14203 (N_14203,N_6108,N_8465);
nand U14204 (N_14204,N_9944,N_8686);
nor U14205 (N_14205,N_5827,N_7392);
or U14206 (N_14206,N_8007,N_5206);
nand U14207 (N_14207,N_9706,N_5713);
nand U14208 (N_14208,N_7212,N_9794);
or U14209 (N_14209,N_6397,N_6380);
and U14210 (N_14210,N_7330,N_6464);
nand U14211 (N_14211,N_7000,N_7792);
or U14212 (N_14212,N_8025,N_5534);
nand U14213 (N_14213,N_9524,N_5192);
nand U14214 (N_14214,N_6952,N_8076);
and U14215 (N_14215,N_6954,N_6075);
and U14216 (N_14216,N_9947,N_5144);
nor U14217 (N_14217,N_9250,N_8323);
and U14218 (N_14218,N_9965,N_9760);
and U14219 (N_14219,N_8725,N_8300);
nor U14220 (N_14220,N_7587,N_6048);
nor U14221 (N_14221,N_6891,N_5503);
nor U14222 (N_14222,N_7009,N_6365);
nor U14223 (N_14223,N_6685,N_6844);
xnor U14224 (N_14224,N_8538,N_8350);
nor U14225 (N_14225,N_7161,N_6415);
or U14226 (N_14226,N_5857,N_5044);
and U14227 (N_14227,N_5630,N_7909);
or U14228 (N_14228,N_5918,N_5973);
or U14229 (N_14229,N_9029,N_5622);
nand U14230 (N_14230,N_9156,N_7392);
and U14231 (N_14231,N_8068,N_9959);
nand U14232 (N_14232,N_8169,N_9780);
or U14233 (N_14233,N_8233,N_6120);
nor U14234 (N_14234,N_5340,N_8915);
nor U14235 (N_14235,N_9046,N_9236);
nand U14236 (N_14236,N_6174,N_9082);
nand U14237 (N_14237,N_5727,N_7405);
nand U14238 (N_14238,N_5071,N_7678);
or U14239 (N_14239,N_6823,N_8477);
and U14240 (N_14240,N_6845,N_6127);
or U14241 (N_14241,N_8731,N_5746);
or U14242 (N_14242,N_6352,N_9856);
and U14243 (N_14243,N_5774,N_9766);
and U14244 (N_14244,N_6697,N_5435);
nand U14245 (N_14245,N_9552,N_5451);
nor U14246 (N_14246,N_6599,N_7893);
and U14247 (N_14247,N_9572,N_5375);
and U14248 (N_14248,N_9178,N_9606);
nor U14249 (N_14249,N_9395,N_9873);
xor U14250 (N_14250,N_6699,N_6861);
or U14251 (N_14251,N_7502,N_8982);
nor U14252 (N_14252,N_8798,N_9637);
or U14253 (N_14253,N_8855,N_5358);
nor U14254 (N_14254,N_6988,N_6469);
xor U14255 (N_14255,N_9846,N_6451);
xnor U14256 (N_14256,N_6516,N_9630);
and U14257 (N_14257,N_5804,N_5201);
xor U14258 (N_14258,N_8682,N_6297);
or U14259 (N_14259,N_9728,N_6133);
or U14260 (N_14260,N_8155,N_5944);
and U14261 (N_14261,N_5873,N_6851);
and U14262 (N_14262,N_6025,N_9847);
or U14263 (N_14263,N_9216,N_5138);
xor U14264 (N_14264,N_9460,N_6681);
or U14265 (N_14265,N_5416,N_8493);
xor U14266 (N_14266,N_5228,N_7189);
xor U14267 (N_14267,N_5746,N_8472);
and U14268 (N_14268,N_5869,N_6555);
nand U14269 (N_14269,N_8778,N_8683);
nor U14270 (N_14270,N_8899,N_7101);
nand U14271 (N_14271,N_6087,N_6730);
nor U14272 (N_14272,N_5920,N_9841);
nand U14273 (N_14273,N_8141,N_6888);
or U14274 (N_14274,N_9264,N_9063);
nand U14275 (N_14275,N_5841,N_9909);
and U14276 (N_14276,N_5810,N_8402);
and U14277 (N_14277,N_7443,N_8432);
nor U14278 (N_14278,N_6671,N_8626);
nand U14279 (N_14279,N_8072,N_9603);
and U14280 (N_14280,N_5004,N_7705);
nor U14281 (N_14281,N_9801,N_7392);
or U14282 (N_14282,N_7912,N_6623);
nand U14283 (N_14283,N_7388,N_8244);
and U14284 (N_14284,N_5958,N_9143);
xor U14285 (N_14285,N_5751,N_6991);
and U14286 (N_14286,N_9387,N_9257);
and U14287 (N_14287,N_8859,N_9105);
nor U14288 (N_14288,N_6688,N_6359);
or U14289 (N_14289,N_7753,N_9434);
and U14290 (N_14290,N_6036,N_9455);
or U14291 (N_14291,N_8104,N_9118);
nor U14292 (N_14292,N_5141,N_7139);
nand U14293 (N_14293,N_5311,N_5045);
and U14294 (N_14294,N_7488,N_5509);
xnor U14295 (N_14295,N_5776,N_6841);
nor U14296 (N_14296,N_7682,N_6678);
or U14297 (N_14297,N_7086,N_5230);
or U14298 (N_14298,N_9824,N_6893);
and U14299 (N_14299,N_7913,N_9781);
nor U14300 (N_14300,N_6520,N_9329);
nor U14301 (N_14301,N_7919,N_9589);
or U14302 (N_14302,N_6922,N_7078);
nor U14303 (N_14303,N_6977,N_6500);
or U14304 (N_14304,N_5626,N_5062);
or U14305 (N_14305,N_9514,N_5110);
nor U14306 (N_14306,N_9551,N_9762);
and U14307 (N_14307,N_9855,N_8181);
nand U14308 (N_14308,N_5928,N_5319);
and U14309 (N_14309,N_6348,N_8159);
nand U14310 (N_14310,N_7849,N_7418);
nand U14311 (N_14311,N_6462,N_7402);
xor U14312 (N_14312,N_6819,N_6140);
nor U14313 (N_14313,N_6710,N_8131);
nor U14314 (N_14314,N_8332,N_5760);
nor U14315 (N_14315,N_7773,N_8244);
xnor U14316 (N_14316,N_6963,N_8915);
and U14317 (N_14317,N_8990,N_8180);
nor U14318 (N_14318,N_6454,N_5281);
nor U14319 (N_14319,N_7314,N_7343);
and U14320 (N_14320,N_7508,N_8825);
or U14321 (N_14321,N_9999,N_9941);
or U14322 (N_14322,N_5820,N_7963);
nand U14323 (N_14323,N_8106,N_8374);
or U14324 (N_14324,N_7355,N_9742);
and U14325 (N_14325,N_8923,N_8161);
nor U14326 (N_14326,N_7647,N_6809);
xor U14327 (N_14327,N_7934,N_5792);
and U14328 (N_14328,N_9748,N_9557);
nor U14329 (N_14329,N_6263,N_9059);
and U14330 (N_14330,N_8338,N_9542);
nor U14331 (N_14331,N_8084,N_7655);
and U14332 (N_14332,N_8673,N_7987);
nand U14333 (N_14333,N_9871,N_6802);
nand U14334 (N_14334,N_9555,N_6291);
nor U14335 (N_14335,N_6032,N_7647);
nor U14336 (N_14336,N_8721,N_9397);
nand U14337 (N_14337,N_6989,N_5520);
or U14338 (N_14338,N_5231,N_8860);
or U14339 (N_14339,N_6247,N_7535);
or U14340 (N_14340,N_5680,N_5817);
nor U14341 (N_14341,N_5218,N_6907);
and U14342 (N_14342,N_5444,N_7831);
nand U14343 (N_14343,N_8412,N_5634);
and U14344 (N_14344,N_8417,N_8765);
nand U14345 (N_14345,N_8224,N_9821);
nand U14346 (N_14346,N_9293,N_6064);
nand U14347 (N_14347,N_5347,N_9949);
nor U14348 (N_14348,N_7748,N_9997);
and U14349 (N_14349,N_5858,N_5333);
and U14350 (N_14350,N_8962,N_5590);
nand U14351 (N_14351,N_6874,N_6747);
or U14352 (N_14352,N_8124,N_8558);
nand U14353 (N_14353,N_7792,N_8952);
nor U14354 (N_14354,N_9339,N_6691);
nor U14355 (N_14355,N_6027,N_5737);
nand U14356 (N_14356,N_9780,N_7740);
xnor U14357 (N_14357,N_6624,N_7464);
nand U14358 (N_14358,N_7765,N_5956);
nor U14359 (N_14359,N_8245,N_7725);
or U14360 (N_14360,N_9276,N_9742);
nand U14361 (N_14361,N_9285,N_6662);
nor U14362 (N_14362,N_8342,N_8804);
or U14363 (N_14363,N_8290,N_8488);
and U14364 (N_14364,N_7629,N_9853);
nand U14365 (N_14365,N_9450,N_8072);
and U14366 (N_14366,N_9821,N_7415);
nor U14367 (N_14367,N_8714,N_8541);
nand U14368 (N_14368,N_8482,N_7877);
nand U14369 (N_14369,N_9051,N_5994);
nor U14370 (N_14370,N_9493,N_5892);
nand U14371 (N_14371,N_9540,N_9150);
nor U14372 (N_14372,N_6165,N_8905);
and U14373 (N_14373,N_5918,N_6516);
nand U14374 (N_14374,N_9890,N_7511);
and U14375 (N_14375,N_9598,N_5813);
xor U14376 (N_14376,N_6344,N_7357);
or U14377 (N_14377,N_6396,N_5201);
nand U14378 (N_14378,N_7677,N_9186);
and U14379 (N_14379,N_8524,N_6465);
nand U14380 (N_14380,N_9086,N_6978);
and U14381 (N_14381,N_6502,N_8092);
or U14382 (N_14382,N_7183,N_6826);
and U14383 (N_14383,N_5396,N_5588);
nor U14384 (N_14384,N_7128,N_5643);
nand U14385 (N_14385,N_8172,N_9883);
or U14386 (N_14386,N_8740,N_5139);
nor U14387 (N_14387,N_9342,N_5863);
xnor U14388 (N_14388,N_9801,N_9421);
or U14389 (N_14389,N_6625,N_6678);
or U14390 (N_14390,N_7895,N_6673);
and U14391 (N_14391,N_8136,N_6192);
nand U14392 (N_14392,N_6086,N_9125);
nand U14393 (N_14393,N_8966,N_6028);
nand U14394 (N_14394,N_6090,N_6906);
xor U14395 (N_14395,N_9056,N_9613);
nand U14396 (N_14396,N_9608,N_9114);
xor U14397 (N_14397,N_6336,N_6649);
or U14398 (N_14398,N_7187,N_6155);
nand U14399 (N_14399,N_8711,N_9930);
nand U14400 (N_14400,N_9654,N_6425);
and U14401 (N_14401,N_5055,N_8725);
or U14402 (N_14402,N_6099,N_6688);
nand U14403 (N_14403,N_8631,N_6592);
nor U14404 (N_14404,N_8439,N_7237);
or U14405 (N_14405,N_7668,N_8264);
and U14406 (N_14406,N_6810,N_6800);
or U14407 (N_14407,N_7812,N_5315);
or U14408 (N_14408,N_9561,N_8177);
nand U14409 (N_14409,N_8937,N_7786);
or U14410 (N_14410,N_5698,N_8503);
xnor U14411 (N_14411,N_5425,N_5146);
nand U14412 (N_14412,N_7604,N_6335);
nand U14413 (N_14413,N_9371,N_9299);
nor U14414 (N_14414,N_5104,N_8339);
nand U14415 (N_14415,N_7865,N_7331);
xor U14416 (N_14416,N_9940,N_7556);
or U14417 (N_14417,N_6360,N_5795);
and U14418 (N_14418,N_6406,N_7416);
nand U14419 (N_14419,N_6758,N_7491);
and U14420 (N_14420,N_8362,N_6409);
or U14421 (N_14421,N_6929,N_5891);
or U14422 (N_14422,N_9054,N_5303);
xnor U14423 (N_14423,N_7069,N_6671);
and U14424 (N_14424,N_6949,N_9472);
nand U14425 (N_14425,N_7321,N_8060);
and U14426 (N_14426,N_8089,N_5462);
and U14427 (N_14427,N_9728,N_7190);
nand U14428 (N_14428,N_9674,N_6918);
and U14429 (N_14429,N_9840,N_5705);
nor U14430 (N_14430,N_8708,N_5805);
nand U14431 (N_14431,N_7254,N_8400);
nor U14432 (N_14432,N_9794,N_9674);
or U14433 (N_14433,N_8411,N_8876);
nor U14434 (N_14434,N_9490,N_9111);
and U14435 (N_14435,N_9526,N_5200);
xor U14436 (N_14436,N_9345,N_6877);
nand U14437 (N_14437,N_8530,N_9291);
or U14438 (N_14438,N_9250,N_6299);
nand U14439 (N_14439,N_9460,N_9255);
or U14440 (N_14440,N_9185,N_5844);
and U14441 (N_14441,N_8508,N_8433);
nor U14442 (N_14442,N_8105,N_9217);
or U14443 (N_14443,N_7853,N_6353);
nand U14444 (N_14444,N_5937,N_9137);
and U14445 (N_14445,N_6416,N_7659);
or U14446 (N_14446,N_7788,N_8417);
xor U14447 (N_14447,N_8590,N_8028);
and U14448 (N_14448,N_5532,N_7600);
nor U14449 (N_14449,N_9244,N_9236);
xor U14450 (N_14450,N_9742,N_7075);
nor U14451 (N_14451,N_7396,N_9694);
nor U14452 (N_14452,N_9569,N_7277);
xnor U14453 (N_14453,N_6725,N_8326);
nor U14454 (N_14454,N_8197,N_8053);
nor U14455 (N_14455,N_7037,N_5566);
or U14456 (N_14456,N_5218,N_6504);
nor U14457 (N_14457,N_5298,N_8816);
or U14458 (N_14458,N_5774,N_7637);
nor U14459 (N_14459,N_8295,N_5717);
nor U14460 (N_14460,N_8259,N_5880);
xor U14461 (N_14461,N_9994,N_5803);
nand U14462 (N_14462,N_7706,N_8827);
nor U14463 (N_14463,N_8086,N_9637);
nand U14464 (N_14464,N_6824,N_7161);
nor U14465 (N_14465,N_8559,N_6268);
or U14466 (N_14466,N_5783,N_7181);
nor U14467 (N_14467,N_6863,N_9669);
nor U14468 (N_14468,N_6876,N_6188);
xnor U14469 (N_14469,N_8335,N_6686);
and U14470 (N_14470,N_8217,N_6607);
nor U14471 (N_14471,N_9584,N_5751);
or U14472 (N_14472,N_9405,N_6236);
xor U14473 (N_14473,N_7798,N_8480);
nor U14474 (N_14474,N_7403,N_5836);
and U14475 (N_14475,N_9571,N_6194);
xnor U14476 (N_14476,N_7858,N_9318);
or U14477 (N_14477,N_5940,N_9465);
and U14478 (N_14478,N_6526,N_5201);
xnor U14479 (N_14479,N_9964,N_9701);
or U14480 (N_14480,N_9986,N_7087);
nand U14481 (N_14481,N_8876,N_5470);
or U14482 (N_14482,N_7514,N_8335);
nor U14483 (N_14483,N_9735,N_7223);
and U14484 (N_14484,N_9606,N_5322);
nand U14485 (N_14485,N_9449,N_6356);
nor U14486 (N_14486,N_7192,N_6823);
and U14487 (N_14487,N_5096,N_5295);
and U14488 (N_14488,N_8367,N_6386);
xor U14489 (N_14489,N_6183,N_7739);
xor U14490 (N_14490,N_9911,N_8652);
xnor U14491 (N_14491,N_5632,N_5951);
and U14492 (N_14492,N_8398,N_6772);
nor U14493 (N_14493,N_8503,N_7529);
and U14494 (N_14494,N_5610,N_7217);
nor U14495 (N_14495,N_7594,N_7528);
nor U14496 (N_14496,N_8255,N_8098);
nand U14497 (N_14497,N_5506,N_5269);
nand U14498 (N_14498,N_7941,N_7648);
and U14499 (N_14499,N_8883,N_7445);
nand U14500 (N_14500,N_6686,N_7943);
or U14501 (N_14501,N_8378,N_6129);
nor U14502 (N_14502,N_5112,N_6713);
nor U14503 (N_14503,N_5384,N_6422);
nor U14504 (N_14504,N_8184,N_9647);
and U14505 (N_14505,N_6533,N_6763);
or U14506 (N_14506,N_8274,N_9444);
nand U14507 (N_14507,N_9174,N_8795);
or U14508 (N_14508,N_7130,N_6334);
nor U14509 (N_14509,N_5650,N_8708);
nand U14510 (N_14510,N_6249,N_5381);
nor U14511 (N_14511,N_5522,N_8192);
xnor U14512 (N_14512,N_9622,N_5388);
and U14513 (N_14513,N_6318,N_9300);
nor U14514 (N_14514,N_9593,N_7467);
and U14515 (N_14515,N_7081,N_6862);
nor U14516 (N_14516,N_9726,N_7802);
nor U14517 (N_14517,N_7131,N_5795);
nor U14518 (N_14518,N_9898,N_8614);
and U14519 (N_14519,N_5633,N_8724);
nor U14520 (N_14520,N_5767,N_8215);
nand U14521 (N_14521,N_9564,N_6441);
and U14522 (N_14522,N_9866,N_9404);
nor U14523 (N_14523,N_8035,N_8881);
nand U14524 (N_14524,N_5429,N_8177);
nand U14525 (N_14525,N_6691,N_5920);
nand U14526 (N_14526,N_7566,N_5389);
nand U14527 (N_14527,N_6746,N_6655);
and U14528 (N_14528,N_5473,N_6610);
xnor U14529 (N_14529,N_6858,N_8984);
nand U14530 (N_14530,N_9211,N_8027);
or U14531 (N_14531,N_7316,N_9112);
nand U14532 (N_14532,N_9861,N_6557);
nor U14533 (N_14533,N_5050,N_8424);
or U14534 (N_14534,N_6850,N_5080);
xor U14535 (N_14535,N_9917,N_9147);
and U14536 (N_14536,N_7518,N_6774);
or U14537 (N_14537,N_7780,N_9776);
nand U14538 (N_14538,N_8581,N_8874);
xor U14539 (N_14539,N_9254,N_8322);
and U14540 (N_14540,N_7130,N_8880);
and U14541 (N_14541,N_7116,N_9335);
and U14542 (N_14542,N_5017,N_5813);
nand U14543 (N_14543,N_8149,N_8816);
nor U14544 (N_14544,N_5519,N_9260);
nand U14545 (N_14545,N_8704,N_5486);
nor U14546 (N_14546,N_6617,N_6741);
or U14547 (N_14547,N_5392,N_8888);
and U14548 (N_14548,N_6498,N_6965);
and U14549 (N_14549,N_7188,N_6252);
nand U14550 (N_14550,N_8440,N_7691);
xnor U14551 (N_14551,N_6496,N_9232);
or U14552 (N_14552,N_9169,N_6807);
xor U14553 (N_14553,N_7348,N_7522);
xnor U14554 (N_14554,N_8371,N_8571);
and U14555 (N_14555,N_7931,N_6830);
nor U14556 (N_14556,N_7289,N_8642);
nor U14557 (N_14557,N_5364,N_7869);
nand U14558 (N_14558,N_9457,N_6510);
nand U14559 (N_14559,N_7081,N_8593);
or U14560 (N_14560,N_9411,N_9395);
and U14561 (N_14561,N_7386,N_8144);
nand U14562 (N_14562,N_8336,N_7036);
or U14563 (N_14563,N_7041,N_5939);
or U14564 (N_14564,N_9547,N_9485);
nand U14565 (N_14565,N_5651,N_6094);
and U14566 (N_14566,N_7690,N_6223);
nand U14567 (N_14567,N_9626,N_6503);
nand U14568 (N_14568,N_9048,N_8276);
and U14569 (N_14569,N_6745,N_8409);
and U14570 (N_14570,N_7858,N_9436);
and U14571 (N_14571,N_7183,N_8621);
xnor U14572 (N_14572,N_6091,N_9534);
or U14573 (N_14573,N_6617,N_9693);
nand U14574 (N_14574,N_6770,N_5279);
and U14575 (N_14575,N_7377,N_8250);
and U14576 (N_14576,N_9200,N_6736);
and U14577 (N_14577,N_7741,N_7586);
nor U14578 (N_14578,N_5628,N_8825);
or U14579 (N_14579,N_6370,N_8615);
nor U14580 (N_14580,N_8365,N_8392);
or U14581 (N_14581,N_9929,N_7516);
or U14582 (N_14582,N_5198,N_6586);
and U14583 (N_14583,N_5918,N_7293);
nand U14584 (N_14584,N_6463,N_6073);
and U14585 (N_14585,N_7393,N_9972);
and U14586 (N_14586,N_7708,N_6722);
or U14587 (N_14587,N_7999,N_6940);
or U14588 (N_14588,N_9306,N_6381);
or U14589 (N_14589,N_6522,N_6664);
or U14590 (N_14590,N_8277,N_7579);
nor U14591 (N_14591,N_5465,N_5123);
and U14592 (N_14592,N_6728,N_5504);
or U14593 (N_14593,N_5849,N_7662);
or U14594 (N_14594,N_5805,N_8768);
or U14595 (N_14595,N_6999,N_7429);
or U14596 (N_14596,N_6276,N_5859);
or U14597 (N_14597,N_8777,N_7870);
or U14598 (N_14598,N_6873,N_6399);
and U14599 (N_14599,N_7919,N_5672);
nand U14600 (N_14600,N_8926,N_6436);
or U14601 (N_14601,N_8035,N_6958);
nand U14602 (N_14602,N_9625,N_5440);
and U14603 (N_14603,N_5541,N_9333);
and U14604 (N_14604,N_8858,N_5523);
or U14605 (N_14605,N_9496,N_7264);
xor U14606 (N_14606,N_6186,N_6750);
nand U14607 (N_14607,N_7195,N_9587);
and U14608 (N_14608,N_6988,N_6473);
nor U14609 (N_14609,N_9577,N_9741);
or U14610 (N_14610,N_8971,N_5658);
and U14611 (N_14611,N_5824,N_8801);
nand U14612 (N_14612,N_6719,N_9983);
nor U14613 (N_14613,N_7555,N_5160);
xor U14614 (N_14614,N_9797,N_6582);
or U14615 (N_14615,N_9179,N_7653);
nor U14616 (N_14616,N_6302,N_9785);
and U14617 (N_14617,N_8688,N_5828);
xnor U14618 (N_14618,N_8313,N_9771);
nor U14619 (N_14619,N_7035,N_9344);
xor U14620 (N_14620,N_7743,N_6860);
nand U14621 (N_14621,N_9458,N_5536);
and U14622 (N_14622,N_5407,N_8861);
nor U14623 (N_14623,N_8425,N_8062);
or U14624 (N_14624,N_9876,N_5691);
and U14625 (N_14625,N_7055,N_5505);
or U14626 (N_14626,N_9014,N_9269);
nor U14627 (N_14627,N_7341,N_5730);
or U14628 (N_14628,N_7212,N_6194);
nand U14629 (N_14629,N_9259,N_5001);
nand U14630 (N_14630,N_6503,N_9390);
and U14631 (N_14631,N_9545,N_5865);
nor U14632 (N_14632,N_5634,N_9654);
and U14633 (N_14633,N_7105,N_8415);
and U14634 (N_14634,N_6334,N_7500);
and U14635 (N_14635,N_6349,N_8722);
and U14636 (N_14636,N_9489,N_9629);
or U14637 (N_14637,N_8595,N_5670);
nand U14638 (N_14638,N_5561,N_5351);
xor U14639 (N_14639,N_7053,N_5854);
and U14640 (N_14640,N_9122,N_9247);
and U14641 (N_14641,N_6212,N_9919);
or U14642 (N_14642,N_7740,N_8059);
and U14643 (N_14643,N_8004,N_8135);
nor U14644 (N_14644,N_7545,N_8138);
nand U14645 (N_14645,N_5483,N_8959);
or U14646 (N_14646,N_6714,N_5334);
nor U14647 (N_14647,N_5212,N_6725);
and U14648 (N_14648,N_7146,N_8407);
xor U14649 (N_14649,N_5753,N_7401);
or U14650 (N_14650,N_5510,N_9039);
and U14651 (N_14651,N_6675,N_5279);
nor U14652 (N_14652,N_7581,N_6270);
nor U14653 (N_14653,N_8032,N_5007);
and U14654 (N_14654,N_8785,N_6347);
nand U14655 (N_14655,N_7511,N_5628);
nand U14656 (N_14656,N_9452,N_8336);
or U14657 (N_14657,N_8232,N_7485);
nor U14658 (N_14658,N_7438,N_7956);
nand U14659 (N_14659,N_7854,N_6817);
or U14660 (N_14660,N_9495,N_7792);
xor U14661 (N_14661,N_7478,N_9620);
or U14662 (N_14662,N_8871,N_7055);
and U14663 (N_14663,N_7633,N_5587);
xnor U14664 (N_14664,N_5015,N_8311);
nor U14665 (N_14665,N_5204,N_5814);
or U14666 (N_14666,N_5671,N_6702);
and U14667 (N_14667,N_8283,N_9161);
nand U14668 (N_14668,N_6111,N_7337);
nor U14669 (N_14669,N_9055,N_7330);
nand U14670 (N_14670,N_5732,N_5513);
or U14671 (N_14671,N_5336,N_5290);
nor U14672 (N_14672,N_8288,N_9587);
nor U14673 (N_14673,N_7839,N_9230);
nor U14674 (N_14674,N_6372,N_7431);
and U14675 (N_14675,N_5952,N_7435);
and U14676 (N_14676,N_8001,N_9819);
nor U14677 (N_14677,N_5615,N_7186);
nand U14678 (N_14678,N_6107,N_6242);
or U14679 (N_14679,N_6063,N_5387);
and U14680 (N_14680,N_9877,N_9220);
or U14681 (N_14681,N_9075,N_9180);
nand U14682 (N_14682,N_8953,N_8591);
nor U14683 (N_14683,N_8651,N_5074);
nor U14684 (N_14684,N_9799,N_9275);
or U14685 (N_14685,N_7366,N_6831);
and U14686 (N_14686,N_9540,N_5629);
nor U14687 (N_14687,N_9066,N_8928);
and U14688 (N_14688,N_6219,N_7395);
or U14689 (N_14689,N_9360,N_5316);
nor U14690 (N_14690,N_7789,N_7920);
nand U14691 (N_14691,N_5805,N_8319);
xor U14692 (N_14692,N_7096,N_6713);
nand U14693 (N_14693,N_7546,N_7681);
and U14694 (N_14694,N_7906,N_8584);
nor U14695 (N_14695,N_5178,N_6587);
and U14696 (N_14696,N_6893,N_6954);
and U14697 (N_14697,N_8116,N_5743);
and U14698 (N_14698,N_9909,N_8635);
nor U14699 (N_14699,N_6925,N_7172);
nand U14700 (N_14700,N_9554,N_8914);
or U14701 (N_14701,N_5073,N_9951);
nor U14702 (N_14702,N_5113,N_5937);
nor U14703 (N_14703,N_5412,N_9911);
and U14704 (N_14704,N_6076,N_7919);
or U14705 (N_14705,N_6002,N_6395);
or U14706 (N_14706,N_5877,N_6919);
and U14707 (N_14707,N_6518,N_6490);
and U14708 (N_14708,N_5744,N_7590);
or U14709 (N_14709,N_6508,N_7587);
nand U14710 (N_14710,N_6493,N_9055);
or U14711 (N_14711,N_7261,N_7774);
and U14712 (N_14712,N_9196,N_5976);
nor U14713 (N_14713,N_8897,N_6078);
nor U14714 (N_14714,N_5683,N_7597);
nand U14715 (N_14715,N_8013,N_6518);
and U14716 (N_14716,N_9157,N_5548);
nand U14717 (N_14717,N_8092,N_5533);
or U14718 (N_14718,N_6178,N_9552);
xnor U14719 (N_14719,N_9165,N_5345);
or U14720 (N_14720,N_6682,N_7425);
and U14721 (N_14721,N_9326,N_9282);
and U14722 (N_14722,N_6140,N_8528);
or U14723 (N_14723,N_5949,N_8053);
nor U14724 (N_14724,N_9466,N_6037);
nand U14725 (N_14725,N_6291,N_7299);
nand U14726 (N_14726,N_7341,N_5748);
nor U14727 (N_14727,N_7733,N_7903);
xnor U14728 (N_14728,N_5042,N_9401);
nor U14729 (N_14729,N_8751,N_5627);
or U14730 (N_14730,N_9169,N_9054);
nand U14731 (N_14731,N_7589,N_8969);
nor U14732 (N_14732,N_8570,N_7842);
and U14733 (N_14733,N_8086,N_8640);
nor U14734 (N_14734,N_6700,N_9085);
nand U14735 (N_14735,N_6505,N_7404);
nand U14736 (N_14736,N_5769,N_8485);
nor U14737 (N_14737,N_7135,N_8450);
and U14738 (N_14738,N_6494,N_5262);
nor U14739 (N_14739,N_8926,N_8658);
or U14740 (N_14740,N_6666,N_6256);
or U14741 (N_14741,N_7982,N_7377);
xnor U14742 (N_14742,N_6150,N_6410);
and U14743 (N_14743,N_6146,N_5051);
nand U14744 (N_14744,N_8448,N_8361);
nor U14745 (N_14745,N_5985,N_7402);
nor U14746 (N_14746,N_8556,N_8956);
or U14747 (N_14747,N_8753,N_8887);
xnor U14748 (N_14748,N_7934,N_8846);
nor U14749 (N_14749,N_7628,N_8795);
xor U14750 (N_14750,N_6384,N_9659);
or U14751 (N_14751,N_8589,N_6030);
xnor U14752 (N_14752,N_5575,N_6421);
nor U14753 (N_14753,N_6587,N_9303);
and U14754 (N_14754,N_9499,N_6269);
and U14755 (N_14755,N_6699,N_6103);
or U14756 (N_14756,N_7135,N_9930);
or U14757 (N_14757,N_9976,N_9584);
nor U14758 (N_14758,N_9426,N_5078);
and U14759 (N_14759,N_9984,N_5359);
or U14760 (N_14760,N_9738,N_8624);
nor U14761 (N_14761,N_7138,N_5154);
xor U14762 (N_14762,N_6284,N_8899);
or U14763 (N_14763,N_6370,N_9155);
nand U14764 (N_14764,N_5128,N_6545);
xor U14765 (N_14765,N_6202,N_7714);
nor U14766 (N_14766,N_8582,N_6300);
nand U14767 (N_14767,N_6942,N_6429);
nand U14768 (N_14768,N_5720,N_5691);
or U14769 (N_14769,N_6478,N_9979);
or U14770 (N_14770,N_8064,N_7580);
xnor U14771 (N_14771,N_9705,N_8580);
nand U14772 (N_14772,N_7218,N_5604);
nand U14773 (N_14773,N_7327,N_6807);
and U14774 (N_14774,N_9837,N_8929);
and U14775 (N_14775,N_6526,N_6466);
nor U14776 (N_14776,N_6825,N_5982);
nor U14777 (N_14777,N_8228,N_7480);
and U14778 (N_14778,N_6784,N_8197);
nand U14779 (N_14779,N_5517,N_9276);
nand U14780 (N_14780,N_6842,N_8962);
and U14781 (N_14781,N_5045,N_9692);
or U14782 (N_14782,N_5621,N_6508);
or U14783 (N_14783,N_6089,N_5478);
and U14784 (N_14784,N_5662,N_8629);
or U14785 (N_14785,N_6082,N_7952);
and U14786 (N_14786,N_8571,N_7580);
and U14787 (N_14787,N_7712,N_9667);
nor U14788 (N_14788,N_7193,N_5657);
nor U14789 (N_14789,N_5754,N_5049);
and U14790 (N_14790,N_6914,N_8099);
and U14791 (N_14791,N_6254,N_7467);
nand U14792 (N_14792,N_6013,N_6455);
and U14793 (N_14793,N_8673,N_8725);
or U14794 (N_14794,N_6362,N_7909);
xnor U14795 (N_14795,N_5553,N_8260);
nand U14796 (N_14796,N_5950,N_7506);
xnor U14797 (N_14797,N_6874,N_9799);
or U14798 (N_14798,N_6576,N_8707);
nor U14799 (N_14799,N_9706,N_5517);
or U14800 (N_14800,N_9565,N_9484);
and U14801 (N_14801,N_6445,N_7973);
nand U14802 (N_14802,N_5985,N_8937);
or U14803 (N_14803,N_6942,N_7496);
or U14804 (N_14804,N_8666,N_5425);
nand U14805 (N_14805,N_7616,N_7091);
nand U14806 (N_14806,N_8914,N_7697);
xor U14807 (N_14807,N_5040,N_5808);
xnor U14808 (N_14808,N_8201,N_8883);
nor U14809 (N_14809,N_7029,N_9849);
nand U14810 (N_14810,N_7842,N_6148);
nor U14811 (N_14811,N_8206,N_5649);
and U14812 (N_14812,N_8735,N_9358);
nor U14813 (N_14813,N_9089,N_5106);
or U14814 (N_14814,N_7899,N_7649);
nand U14815 (N_14815,N_7765,N_6098);
and U14816 (N_14816,N_6860,N_6393);
nor U14817 (N_14817,N_5941,N_8550);
nand U14818 (N_14818,N_6240,N_5071);
and U14819 (N_14819,N_7435,N_7031);
xnor U14820 (N_14820,N_6598,N_8270);
xor U14821 (N_14821,N_8825,N_9997);
and U14822 (N_14822,N_5445,N_6006);
and U14823 (N_14823,N_8011,N_7489);
xnor U14824 (N_14824,N_8063,N_6995);
or U14825 (N_14825,N_9354,N_6535);
nor U14826 (N_14826,N_5169,N_8569);
nand U14827 (N_14827,N_6952,N_6241);
nor U14828 (N_14828,N_7485,N_8794);
or U14829 (N_14829,N_5901,N_5352);
nand U14830 (N_14830,N_5874,N_9438);
or U14831 (N_14831,N_9420,N_6263);
nor U14832 (N_14832,N_8867,N_6181);
nand U14833 (N_14833,N_7442,N_7257);
and U14834 (N_14834,N_5121,N_8992);
and U14835 (N_14835,N_5388,N_6345);
nor U14836 (N_14836,N_9314,N_5694);
nor U14837 (N_14837,N_5938,N_5159);
xor U14838 (N_14838,N_7269,N_8122);
nor U14839 (N_14839,N_9108,N_5993);
or U14840 (N_14840,N_9069,N_9926);
and U14841 (N_14841,N_9601,N_8938);
and U14842 (N_14842,N_5097,N_5934);
nor U14843 (N_14843,N_6847,N_6717);
and U14844 (N_14844,N_6312,N_9191);
or U14845 (N_14845,N_7519,N_7231);
and U14846 (N_14846,N_9434,N_9039);
and U14847 (N_14847,N_8272,N_5003);
nand U14848 (N_14848,N_9338,N_6236);
nor U14849 (N_14849,N_8402,N_7265);
nand U14850 (N_14850,N_8565,N_5104);
or U14851 (N_14851,N_6380,N_7397);
nand U14852 (N_14852,N_7627,N_8022);
xor U14853 (N_14853,N_7721,N_5165);
nand U14854 (N_14854,N_6261,N_7718);
nor U14855 (N_14855,N_7598,N_7714);
nand U14856 (N_14856,N_9060,N_9396);
or U14857 (N_14857,N_9883,N_9508);
nor U14858 (N_14858,N_8567,N_5133);
or U14859 (N_14859,N_8730,N_8393);
or U14860 (N_14860,N_6813,N_7372);
or U14861 (N_14861,N_6982,N_8135);
or U14862 (N_14862,N_9247,N_6913);
and U14863 (N_14863,N_5571,N_9245);
xnor U14864 (N_14864,N_6266,N_5229);
and U14865 (N_14865,N_9890,N_7767);
nand U14866 (N_14866,N_5755,N_9561);
nor U14867 (N_14867,N_6185,N_5343);
and U14868 (N_14868,N_7245,N_6082);
nand U14869 (N_14869,N_6501,N_7091);
or U14870 (N_14870,N_9702,N_9468);
nor U14871 (N_14871,N_9196,N_8542);
or U14872 (N_14872,N_7132,N_5803);
nand U14873 (N_14873,N_9585,N_5606);
nor U14874 (N_14874,N_9452,N_8659);
or U14875 (N_14875,N_8832,N_9422);
nand U14876 (N_14876,N_6038,N_7130);
and U14877 (N_14877,N_8975,N_9300);
nand U14878 (N_14878,N_5205,N_7553);
nand U14879 (N_14879,N_6960,N_6767);
or U14880 (N_14880,N_7184,N_9383);
and U14881 (N_14881,N_6408,N_6035);
or U14882 (N_14882,N_6128,N_9693);
or U14883 (N_14883,N_8224,N_6736);
nand U14884 (N_14884,N_5173,N_9999);
and U14885 (N_14885,N_5400,N_6475);
and U14886 (N_14886,N_9309,N_7922);
nand U14887 (N_14887,N_6654,N_8840);
and U14888 (N_14888,N_8233,N_9357);
nand U14889 (N_14889,N_9674,N_6134);
nor U14890 (N_14890,N_6427,N_7829);
xor U14891 (N_14891,N_7565,N_8529);
or U14892 (N_14892,N_9787,N_6086);
nor U14893 (N_14893,N_6080,N_5285);
or U14894 (N_14894,N_7186,N_9856);
or U14895 (N_14895,N_9666,N_9522);
nor U14896 (N_14896,N_8681,N_6008);
nor U14897 (N_14897,N_8868,N_8719);
nand U14898 (N_14898,N_8699,N_5739);
nand U14899 (N_14899,N_5408,N_7664);
and U14900 (N_14900,N_5367,N_8418);
and U14901 (N_14901,N_5444,N_9454);
or U14902 (N_14902,N_7529,N_9623);
nor U14903 (N_14903,N_8941,N_8924);
or U14904 (N_14904,N_7167,N_5612);
nand U14905 (N_14905,N_9557,N_5850);
nor U14906 (N_14906,N_8509,N_5880);
and U14907 (N_14907,N_5981,N_6354);
and U14908 (N_14908,N_7899,N_8073);
and U14909 (N_14909,N_8674,N_6498);
or U14910 (N_14910,N_7227,N_9416);
nand U14911 (N_14911,N_5751,N_8933);
or U14912 (N_14912,N_6952,N_9550);
or U14913 (N_14913,N_7119,N_5266);
xor U14914 (N_14914,N_7723,N_7794);
xnor U14915 (N_14915,N_6238,N_9919);
and U14916 (N_14916,N_6785,N_6178);
xnor U14917 (N_14917,N_7553,N_9578);
nor U14918 (N_14918,N_7277,N_6304);
nand U14919 (N_14919,N_5662,N_9753);
nor U14920 (N_14920,N_6790,N_7417);
xnor U14921 (N_14921,N_6048,N_5722);
and U14922 (N_14922,N_5348,N_7847);
and U14923 (N_14923,N_8453,N_5462);
nand U14924 (N_14924,N_7746,N_5932);
and U14925 (N_14925,N_7362,N_5338);
nand U14926 (N_14926,N_9523,N_7970);
nor U14927 (N_14927,N_8629,N_8891);
nor U14928 (N_14928,N_7737,N_8525);
and U14929 (N_14929,N_9433,N_7429);
nor U14930 (N_14930,N_7810,N_7015);
and U14931 (N_14931,N_8300,N_7559);
nor U14932 (N_14932,N_9671,N_8572);
xnor U14933 (N_14933,N_9973,N_5881);
nand U14934 (N_14934,N_8776,N_6535);
nor U14935 (N_14935,N_7951,N_6284);
nand U14936 (N_14936,N_5578,N_9361);
and U14937 (N_14937,N_9409,N_6221);
and U14938 (N_14938,N_7957,N_5035);
nor U14939 (N_14939,N_5284,N_6247);
xnor U14940 (N_14940,N_9458,N_6172);
nor U14941 (N_14941,N_5312,N_6893);
nor U14942 (N_14942,N_7840,N_5969);
xnor U14943 (N_14943,N_9334,N_7252);
or U14944 (N_14944,N_8572,N_6587);
and U14945 (N_14945,N_6145,N_9584);
and U14946 (N_14946,N_7089,N_8332);
nor U14947 (N_14947,N_6527,N_8092);
xor U14948 (N_14948,N_5415,N_6370);
or U14949 (N_14949,N_5691,N_5123);
or U14950 (N_14950,N_8501,N_8830);
or U14951 (N_14951,N_5436,N_7029);
nor U14952 (N_14952,N_9233,N_9518);
nor U14953 (N_14953,N_5886,N_9477);
nor U14954 (N_14954,N_5581,N_7690);
nor U14955 (N_14955,N_9291,N_9299);
or U14956 (N_14956,N_9497,N_6561);
nand U14957 (N_14957,N_5194,N_6717);
xnor U14958 (N_14958,N_8886,N_6990);
xnor U14959 (N_14959,N_8990,N_8553);
and U14960 (N_14960,N_8639,N_5382);
and U14961 (N_14961,N_7182,N_6208);
or U14962 (N_14962,N_8793,N_8218);
or U14963 (N_14963,N_6006,N_5229);
xor U14964 (N_14964,N_6935,N_5457);
nand U14965 (N_14965,N_5846,N_6232);
nand U14966 (N_14966,N_6418,N_5200);
nand U14967 (N_14967,N_9420,N_5553);
and U14968 (N_14968,N_7828,N_8298);
or U14969 (N_14969,N_8012,N_6180);
nor U14970 (N_14970,N_5808,N_6317);
nand U14971 (N_14971,N_8886,N_6606);
nor U14972 (N_14972,N_9342,N_9660);
nand U14973 (N_14973,N_8083,N_5723);
nor U14974 (N_14974,N_5459,N_7096);
nor U14975 (N_14975,N_6640,N_7893);
nand U14976 (N_14976,N_9574,N_8381);
nand U14977 (N_14977,N_6243,N_6540);
or U14978 (N_14978,N_7656,N_9244);
and U14979 (N_14979,N_6563,N_8179);
nor U14980 (N_14980,N_7573,N_9393);
and U14981 (N_14981,N_5502,N_6978);
and U14982 (N_14982,N_7947,N_7900);
or U14983 (N_14983,N_5436,N_6106);
or U14984 (N_14984,N_7722,N_6618);
nand U14985 (N_14985,N_8906,N_8590);
nor U14986 (N_14986,N_7017,N_9926);
nand U14987 (N_14987,N_6229,N_6717);
nor U14988 (N_14988,N_9115,N_8943);
nand U14989 (N_14989,N_8784,N_8405);
nor U14990 (N_14990,N_8874,N_6353);
nand U14991 (N_14991,N_5553,N_9292);
and U14992 (N_14992,N_9980,N_6453);
nor U14993 (N_14993,N_7214,N_9222);
nor U14994 (N_14994,N_9569,N_9647);
and U14995 (N_14995,N_9362,N_8934);
and U14996 (N_14996,N_9664,N_5118);
xnor U14997 (N_14997,N_5121,N_5186);
or U14998 (N_14998,N_8672,N_7270);
nor U14999 (N_14999,N_9152,N_6498);
nand U15000 (N_15000,N_12746,N_13504);
nor U15001 (N_15001,N_13321,N_14658);
and U15002 (N_15002,N_12984,N_10134);
nand U15003 (N_15003,N_12235,N_12737);
nor U15004 (N_15004,N_13425,N_12453);
nand U15005 (N_15005,N_12097,N_14756);
nand U15006 (N_15006,N_10261,N_11018);
and U15007 (N_15007,N_11110,N_13974);
and U15008 (N_15008,N_13348,N_11282);
xor U15009 (N_15009,N_10317,N_13331);
nand U15010 (N_15010,N_14456,N_14612);
or U15011 (N_15011,N_12704,N_10325);
and U15012 (N_15012,N_11284,N_14614);
nor U15013 (N_15013,N_14771,N_13773);
xor U15014 (N_15014,N_11427,N_14097);
and U15015 (N_15015,N_10593,N_13806);
xnor U15016 (N_15016,N_11590,N_12364);
and U15017 (N_15017,N_10814,N_13696);
and U15018 (N_15018,N_10313,N_11154);
nand U15019 (N_15019,N_14810,N_10648);
nand U15020 (N_15020,N_13505,N_11687);
and U15021 (N_15021,N_13841,N_10847);
and U15022 (N_15022,N_14419,N_13038);
nor U15023 (N_15023,N_13647,N_11725);
nor U15024 (N_15024,N_10180,N_14371);
nand U15025 (N_15025,N_11360,N_13768);
and U15026 (N_15026,N_10217,N_12058);
or U15027 (N_15027,N_10609,N_10703);
nor U15028 (N_15028,N_13492,N_14285);
and U15029 (N_15029,N_10541,N_14414);
nor U15030 (N_15030,N_12509,N_13958);
nand U15031 (N_15031,N_12233,N_14970);
and U15032 (N_15032,N_12572,N_13774);
nand U15033 (N_15033,N_10408,N_14298);
and U15034 (N_15034,N_14493,N_13084);
or U15035 (N_15035,N_11376,N_12836);
xor U15036 (N_15036,N_14837,N_11966);
nor U15037 (N_15037,N_13398,N_14642);
xnor U15038 (N_15038,N_12371,N_10674);
nor U15039 (N_15039,N_11795,N_14832);
and U15040 (N_15040,N_12851,N_12803);
xnor U15041 (N_15041,N_13883,N_11079);
nand U15042 (N_15042,N_10719,N_13093);
nand U15043 (N_15043,N_12996,N_10548);
nor U15044 (N_15044,N_11092,N_14113);
nand U15045 (N_15045,N_11512,N_10105);
or U15046 (N_15046,N_10854,N_14941);
and U15047 (N_15047,N_13360,N_13596);
and U15048 (N_15048,N_11542,N_14668);
or U15049 (N_15049,N_13961,N_10468);
nand U15050 (N_15050,N_11367,N_11569);
nor U15051 (N_15051,N_13821,N_10725);
xor U15052 (N_15052,N_10666,N_10615);
or U15053 (N_15053,N_14227,N_12722);
nand U15054 (N_15054,N_14813,N_14348);
and U15055 (N_15055,N_12585,N_14959);
nor U15056 (N_15056,N_11767,N_13133);
nor U15057 (N_15057,N_12669,N_14099);
xor U15058 (N_15058,N_12170,N_14039);
or U15059 (N_15059,N_12063,N_13902);
nand U15060 (N_15060,N_10106,N_13631);
and U15061 (N_15061,N_13490,N_10439);
and U15062 (N_15062,N_14715,N_12577);
or U15063 (N_15063,N_13769,N_14996);
xor U15064 (N_15064,N_10855,N_14648);
nor U15065 (N_15065,N_11188,N_12910);
nor U15066 (N_15066,N_14987,N_10170);
and U15067 (N_15067,N_13470,N_13016);
or U15068 (N_15068,N_12379,N_14461);
or U15069 (N_15069,N_13651,N_10024);
and U15070 (N_15070,N_14901,N_13298);
nor U15071 (N_15071,N_11967,N_14569);
nand U15072 (N_15072,N_14939,N_11475);
nand U15073 (N_15073,N_14302,N_14381);
and U15074 (N_15074,N_14253,N_10090);
and U15075 (N_15075,N_13823,N_13280);
nand U15076 (N_15076,N_14033,N_11239);
and U15077 (N_15077,N_11441,N_14281);
or U15078 (N_15078,N_12751,N_12539);
nor U15079 (N_15079,N_14591,N_14586);
nor U15080 (N_15080,N_11036,N_13882);
nand U15081 (N_15081,N_13231,N_13799);
or U15082 (N_15082,N_10019,N_10571);
or U15083 (N_15083,N_13738,N_10359);
nand U15084 (N_15084,N_14952,N_10418);
nor U15085 (N_15085,N_13600,N_13842);
or U15086 (N_15086,N_13538,N_10536);
and U15087 (N_15087,N_10311,N_14573);
xor U15088 (N_15088,N_13199,N_12191);
xor U15089 (N_15089,N_11143,N_11405);
and U15090 (N_15090,N_11872,N_10561);
xnor U15091 (N_15091,N_10691,N_10128);
nor U15092 (N_15092,N_11813,N_14183);
nor U15093 (N_15093,N_12426,N_12439);
xor U15094 (N_15094,N_13818,N_10492);
nor U15095 (N_15095,N_12523,N_14712);
and U15096 (N_15096,N_13182,N_14580);
and U15097 (N_15097,N_13756,N_14009);
nor U15098 (N_15098,N_12346,N_13075);
nand U15099 (N_15099,N_11107,N_10628);
or U15100 (N_15100,N_14861,N_11127);
nor U15101 (N_15101,N_13764,N_10419);
xor U15102 (N_15102,N_12874,N_13173);
nor U15103 (N_15103,N_14080,N_10812);
and U15104 (N_15104,N_14136,N_13071);
nor U15105 (N_15105,N_13645,N_11684);
xor U15106 (N_15106,N_11365,N_14839);
and U15107 (N_15107,N_10328,N_10566);
and U15108 (N_15108,N_13443,N_13664);
nor U15109 (N_15109,N_14283,N_14339);
xor U15110 (N_15110,N_11488,N_14583);
nor U15111 (N_15111,N_10281,N_10277);
nor U15112 (N_15112,N_12457,N_11979);
or U15113 (N_15113,N_13900,N_13397);
nor U15114 (N_15114,N_13185,N_13175);
nand U15115 (N_15115,N_11274,N_10808);
or U15116 (N_15116,N_14278,N_11716);
or U15117 (N_15117,N_12425,N_11269);
or U15118 (N_15118,N_12220,N_14868);
and U15119 (N_15119,N_10710,N_11503);
or U15120 (N_15120,N_10035,N_13471);
nor U15121 (N_15121,N_11290,N_14149);
nand U15122 (N_15122,N_14858,N_10339);
and U15123 (N_15123,N_11436,N_13116);
nand U15124 (N_15124,N_14847,N_11950);
nor U15125 (N_15125,N_11611,N_10165);
nor U15126 (N_15126,N_14507,N_13221);
nor U15127 (N_15127,N_10078,N_13389);
and U15128 (N_15128,N_11189,N_14654);
or U15129 (N_15129,N_14958,N_11869);
and U15130 (N_15130,N_14264,N_10255);
nand U15131 (N_15131,N_11997,N_14155);
nor U15132 (N_15132,N_10399,N_14174);
and U15133 (N_15133,N_11840,N_11697);
nor U15134 (N_15134,N_10163,N_13580);
or U15135 (N_15135,N_14686,N_14262);
nand U15136 (N_15136,N_14675,N_11844);
nor U15137 (N_15137,N_13922,N_12416);
nor U15138 (N_15138,N_14191,N_14116);
or U15139 (N_15139,N_10770,N_10517);
nand U15140 (N_15140,N_10214,N_14060);
and U15141 (N_15141,N_10712,N_12989);
nand U15142 (N_15142,N_11070,N_10154);
or U15143 (N_15143,N_11901,N_13551);
or U15144 (N_15144,N_12405,N_10899);
and U15145 (N_15145,N_13478,N_10864);
xnor U15146 (N_15146,N_11007,N_13669);
and U15147 (N_15147,N_10156,N_12437);
and U15148 (N_15148,N_10876,N_14392);
nor U15149 (N_15149,N_12979,N_10025);
nand U15150 (N_15150,N_11013,N_11287);
or U15151 (N_15151,N_11774,N_13181);
xnor U15152 (N_15152,N_14092,N_12449);
or U15153 (N_15153,N_13826,N_13853);
nor U15154 (N_15154,N_14611,N_14446);
xnor U15155 (N_15155,N_13299,N_14535);
and U15156 (N_15156,N_10365,N_14023);
and U15157 (N_15157,N_10810,N_13254);
or U15158 (N_15158,N_11064,N_13092);
nand U15159 (N_15159,N_14000,N_13160);
and U15160 (N_15160,N_10423,N_12525);
nor U15161 (N_15161,N_12933,N_10693);
xor U15162 (N_15162,N_13088,N_10452);
nand U15163 (N_15163,N_10148,N_10006);
nor U15164 (N_15164,N_11927,N_12810);
and U15165 (N_15165,N_12360,N_10370);
and U15166 (N_15166,N_13165,N_14528);
and U15167 (N_15167,N_11656,N_13134);
nand U15168 (N_15168,N_12090,N_11125);
nand U15169 (N_15169,N_11004,N_13214);
and U15170 (N_15170,N_13909,N_14126);
or U15171 (N_15171,N_11120,N_10574);
and U15172 (N_15172,N_12712,N_12532);
and U15173 (N_15173,N_10977,N_14002);
nand U15174 (N_15174,N_11778,N_14277);
or U15175 (N_15175,N_10224,N_10935);
nor U15176 (N_15176,N_12383,N_14900);
or U15177 (N_15177,N_13447,N_14971);
and U15178 (N_15178,N_14106,N_12269);
and U15179 (N_15179,N_12276,N_11499);
nor U15180 (N_15180,N_13969,N_12195);
nor U15181 (N_15181,N_12628,N_14230);
nor U15182 (N_15182,N_11743,N_10320);
and U15183 (N_15183,N_13822,N_12403);
nor U15184 (N_15184,N_14754,N_14440);
xnor U15185 (N_15185,N_12842,N_11052);
and U15186 (N_15186,N_12375,N_11679);
nor U15187 (N_15187,N_10434,N_12132);
and U15188 (N_15188,N_11345,N_12871);
or U15189 (N_15189,N_11853,N_14484);
nor U15190 (N_15190,N_10984,N_13627);
or U15191 (N_15191,N_10777,N_11948);
nor U15192 (N_15192,N_11889,N_10260);
and U15193 (N_15193,N_12978,N_10064);
and U15194 (N_15194,N_14396,N_11447);
and U15195 (N_15195,N_11226,N_13310);
nand U15196 (N_15196,N_10075,N_10914);
nor U15197 (N_15197,N_12588,N_12126);
or U15198 (N_15198,N_11119,N_14275);
or U15199 (N_15199,N_14318,N_10690);
nor U15200 (N_15200,N_14076,N_10385);
or U15201 (N_15201,N_12596,N_10733);
or U15202 (N_15202,N_14259,N_14038);
or U15203 (N_15203,N_14180,N_12666);
or U15204 (N_15204,N_14869,N_14347);
nor U15205 (N_15205,N_12255,N_10512);
or U15206 (N_15206,N_13949,N_14773);
or U15207 (N_15207,N_14101,N_14159);
or U15208 (N_15208,N_14423,N_12561);
nand U15209 (N_15209,N_11547,N_12782);
and U15210 (N_15210,N_13386,N_14991);
nand U15211 (N_15211,N_12505,N_14804);
nor U15212 (N_15212,N_10034,N_13058);
or U15213 (N_15213,N_13211,N_11208);
nor U15214 (N_15214,N_14359,N_11662);
and U15215 (N_15215,N_12319,N_14747);
nor U15216 (N_15216,N_14037,N_12321);
nand U15217 (N_15217,N_10881,N_13915);
nor U15218 (N_15218,N_10098,N_13128);
nand U15219 (N_15219,N_10240,N_13012);
nand U15220 (N_15220,N_14560,N_12277);
nor U15221 (N_15221,N_11893,N_13438);
nand U15222 (N_15222,N_11255,N_12312);
nor U15223 (N_15223,N_14305,N_14833);
nand U15224 (N_15224,N_12273,N_12774);
nand U15225 (N_15225,N_11409,N_11157);
nand U15226 (N_15226,N_10023,N_10369);
and U15227 (N_15227,N_10605,N_11969);
nor U15228 (N_15228,N_14376,N_10737);
xnor U15229 (N_15229,N_14388,N_12584);
and U15230 (N_15230,N_13779,N_12677);
or U15231 (N_15231,N_10254,N_12600);
nor U15232 (N_15232,N_12189,N_11701);
or U15233 (N_15233,N_11404,N_11056);
xnor U15234 (N_15234,N_10781,N_12470);
and U15235 (N_15235,N_10110,N_12920);
and U15236 (N_15236,N_13145,N_11775);
nor U15237 (N_15237,N_12023,N_12680);
nand U15238 (N_15238,N_13771,N_10069);
xor U15239 (N_15239,N_12099,N_12245);
or U15240 (N_15240,N_14481,N_11112);
nand U15241 (N_15241,N_12185,N_13695);
and U15242 (N_15242,N_13390,N_10179);
nor U15243 (N_15243,N_10947,N_14718);
nor U15244 (N_15244,N_10403,N_10883);
and U15245 (N_15245,N_14225,N_13255);
nand U15246 (N_15246,N_12860,N_14766);
nor U15247 (N_15247,N_13451,N_14759);
and U15248 (N_15248,N_12694,N_13010);
nor U15249 (N_15249,N_14947,N_12864);
nor U15250 (N_15250,N_14843,N_10396);
and U15251 (N_15251,N_13617,N_10870);
nand U15252 (N_15252,N_12696,N_11084);
nor U15253 (N_15253,N_11122,N_13813);
or U15254 (N_15254,N_14962,N_10546);
and U15255 (N_15255,N_13983,N_14834);
nor U15256 (N_15256,N_13239,N_11814);
and U15257 (N_15257,N_10558,N_12804);
and U15258 (N_15258,N_13632,N_10981);
or U15259 (N_15259,N_10708,N_13159);
or U15260 (N_15260,N_12299,N_14653);
nand U15261 (N_15261,N_10203,N_10695);
nand U15262 (N_15262,N_10324,N_13805);
nand U15263 (N_15263,N_10701,N_13735);
and U15264 (N_15264,N_13743,N_10259);
or U15265 (N_15265,N_12018,N_13024);
xor U15266 (N_15266,N_12930,N_10169);
and U15267 (N_15267,N_14995,N_11080);
and U15268 (N_15268,N_13474,N_12314);
or U15269 (N_15269,N_14755,N_10125);
and U15270 (N_15270,N_14503,N_11248);
nor U15271 (N_15271,N_14245,N_14244);
nand U15272 (N_15272,N_12041,N_11314);
nor U15273 (N_15273,N_12318,N_11012);
or U15274 (N_15274,N_11414,N_13599);
nor U15275 (N_15275,N_11210,N_12144);
nor U15276 (N_15276,N_13869,N_13069);
and U15277 (N_15277,N_14306,N_14935);
xnor U15278 (N_15278,N_10803,N_13021);
nor U15279 (N_15279,N_14851,N_12762);
nand U15280 (N_15280,N_13237,N_13573);
or U15281 (N_15281,N_10092,N_10960);
or U15282 (N_15282,N_12711,N_13213);
nand U15283 (N_15283,N_14108,N_14240);
and U15284 (N_15284,N_11257,N_11552);
or U15285 (N_15285,N_12633,N_12905);
nor U15286 (N_15286,N_13685,N_10208);
xor U15287 (N_15287,N_12950,N_13056);
and U15288 (N_15288,N_12637,N_11635);
xor U15289 (N_15289,N_12334,N_11164);
xor U15290 (N_15290,N_10962,N_12591);
nor U15291 (N_15291,N_13448,N_13475);
xor U15292 (N_15292,N_14955,N_14067);
or U15293 (N_15293,N_10166,N_14413);
nand U15294 (N_15294,N_11995,N_13520);
xnor U15295 (N_15295,N_11060,N_11477);
nor U15296 (N_15296,N_11977,N_12858);
nor U15297 (N_15297,N_14053,N_14466);
nor U15298 (N_15298,N_11779,N_10964);
and U15299 (N_15299,N_12395,N_12770);
xnor U15300 (N_15300,N_12355,N_10652);
and U15301 (N_15301,N_13163,N_11909);
xnor U15302 (N_15302,N_12899,N_12545);
nor U15303 (N_15303,N_13709,N_13997);
or U15304 (N_15304,N_13650,N_14160);
nand U15305 (N_15305,N_10307,N_14171);
and U15306 (N_15306,N_13962,N_12567);
nor U15307 (N_15307,N_11249,N_10620);
or U15308 (N_15308,N_11571,N_11088);
xnor U15309 (N_15309,N_12323,N_13320);
xnor U15310 (N_15310,N_11200,N_13592);
nor U15311 (N_15311,N_13750,N_14814);
nor U15312 (N_15312,N_14494,N_13993);
nor U15313 (N_15313,N_11289,N_11683);
nand U15314 (N_15314,N_13081,N_11742);
and U15315 (N_15315,N_10212,N_13571);
and U15316 (N_15316,N_11196,N_10045);
nand U15317 (N_15317,N_12384,N_12703);
nand U15318 (N_15318,N_13780,N_10826);
nand U15319 (N_15319,N_14777,N_14937);
nand U15320 (N_15320,N_14742,N_10298);
nor U15321 (N_15321,N_14677,N_11628);
and U15322 (N_15322,N_13238,N_10435);
and U15323 (N_15323,N_10626,N_13905);
and U15324 (N_15324,N_12004,N_12106);
xor U15325 (N_15325,N_11584,N_13115);
or U15326 (N_15326,N_13266,N_13910);
and U15327 (N_15327,N_11008,N_10951);
or U15328 (N_15328,N_14320,N_12214);
nand U15329 (N_15329,N_14966,N_12915);
nor U15330 (N_15330,N_10150,N_14650);
nand U15331 (N_15331,N_10677,N_13665);
or U15332 (N_15332,N_14566,N_11476);
and U15333 (N_15333,N_12262,N_11241);
nand U15334 (N_15334,N_12209,N_10675);
nor U15335 (N_15335,N_14042,N_14316);
or U15336 (N_15336,N_12216,N_13361);
nor U15337 (N_15337,N_10241,N_13858);
and U15338 (N_15338,N_14062,N_13370);
or U15339 (N_15339,N_13710,N_12192);
xnor U15340 (N_15340,N_11858,N_12678);
or U15341 (N_15341,N_14871,N_12186);
xor U15342 (N_15342,N_12908,N_13112);
or U15343 (N_15343,N_10731,N_13542);
or U15344 (N_15344,N_12648,N_13096);
nor U15345 (N_15345,N_11891,N_10372);
and U15346 (N_15346,N_12503,N_11462);
nor U15347 (N_15347,N_14378,N_10787);
nor U15348 (N_15348,N_13989,N_12753);
nand U15349 (N_15349,N_13688,N_13122);
nor U15350 (N_15350,N_11837,N_13378);
nor U15351 (N_15351,N_13809,N_11279);
and U15352 (N_15352,N_13296,N_11726);
nand U15353 (N_15353,N_14899,N_11090);
nor U15354 (N_15354,N_12227,N_11473);
nand U15355 (N_15355,N_14064,N_12446);
or U15356 (N_15356,N_14075,N_14228);
nor U15357 (N_15357,N_12408,N_10687);
and U15358 (N_15358,N_14252,N_10697);
nand U15359 (N_15359,N_10384,N_13792);
and U15360 (N_15360,N_14107,N_10478);
or U15361 (N_15361,N_14865,N_14189);
or U15362 (N_15362,N_13123,N_11002);
xnor U15363 (N_15363,N_14404,N_13666);
or U15364 (N_15364,N_11236,N_13765);
nor U15365 (N_15365,N_14809,N_11001);
xnor U15366 (N_15366,N_11597,N_12983);
nand U15367 (N_15367,N_12060,N_10642);
or U15368 (N_15368,N_10856,N_10314);
nor U15369 (N_15369,N_12636,N_10665);
or U15370 (N_15370,N_13844,N_11850);
or U15371 (N_15371,N_14104,N_12533);
and U15372 (N_15372,N_11579,N_13379);
nand U15373 (N_15373,N_10604,N_13498);
and U15374 (N_15374,N_12242,N_13547);
nand U15375 (N_15375,N_12530,N_14957);
and U15376 (N_15376,N_14243,N_13790);
nor U15377 (N_15377,N_14472,N_13946);
or U15378 (N_15378,N_12118,N_14515);
xnor U15379 (N_15379,N_14273,N_13248);
nand U15380 (N_15380,N_10650,N_14844);
nor U15381 (N_15381,N_11788,N_11460);
nand U15382 (N_15382,N_10268,N_10059);
xor U15383 (N_15383,N_11881,N_12007);
nand U15384 (N_15384,N_10042,N_11222);
and U15385 (N_15385,N_14087,N_13775);
nand U15386 (N_15386,N_14830,N_14723);
xnor U15387 (N_15387,N_14735,N_10748);
nand U15388 (N_15388,N_14911,N_12026);
nand U15389 (N_15389,N_14822,N_14625);
or U15390 (N_15390,N_13350,N_11372);
or U15391 (N_15391,N_11528,N_11161);
and U15392 (N_15392,N_12849,N_13391);
nand U15393 (N_15393,N_13875,N_10705);
nor U15394 (N_15394,N_13945,N_12166);
nor U15395 (N_15395,N_11972,N_10361);
and U15396 (N_15396,N_10337,N_12368);
xnor U15397 (N_15397,N_10430,N_12499);
and U15398 (N_15398,N_14695,N_11042);
nand U15399 (N_15399,N_13870,N_10636);
and U15400 (N_15400,N_12875,N_12671);
and U15401 (N_15401,N_13080,N_11232);
or U15402 (N_15402,N_14634,N_12517);
or U15403 (N_15403,N_14465,N_10751);
nor U15404 (N_15404,N_14750,N_11915);
or U15405 (N_15405,N_12386,N_14694);
nor U15406 (N_15406,N_14676,N_10834);
nand U15407 (N_15407,N_12583,N_11212);
and U15408 (N_15408,N_10872,N_10722);
and U15409 (N_15409,N_10406,N_10200);
and U15410 (N_15410,N_11906,N_12834);
and U15411 (N_15411,N_10011,N_12404);
and U15412 (N_15412,N_10462,N_11809);
nand U15413 (N_15413,N_10581,N_14795);
nor U15414 (N_15414,N_10638,N_12767);
or U15415 (N_15415,N_12841,N_11659);
nand U15416 (N_15416,N_12549,N_11336);
nor U15417 (N_15417,N_10511,N_14436);
nor U15418 (N_15418,N_13724,N_14998);
or U15419 (N_15419,N_10103,N_12623);
and U15420 (N_15420,N_14597,N_11914);
nand U15421 (N_15421,N_13423,N_14687);
nand U15422 (N_15422,N_13459,N_13405);
nand U15423 (N_15423,N_11507,N_11911);
xnor U15424 (N_15424,N_12709,N_10889);
or U15425 (N_15425,N_14391,N_13003);
or U15426 (N_15426,N_13281,N_10842);
nor U15427 (N_15427,N_10461,N_13440);
and U15428 (N_15428,N_12706,N_13876);
nand U15429 (N_15429,N_13183,N_11424);
nand U15430 (N_15430,N_11066,N_11759);
nand U15431 (N_15431,N_14944,N_12045);
and U15432 (N_15432,N_14195,N_13387);
or U15433 (N_15433,N_14315,N_13245);
xor U15434 (N_15434,N_14117,N_11855);
nor U15435 (N_15435,N_11686,N_11691);
and U15436 (N_15436,N_10031,N_13434);
nand U15437 (N_15437,N_12761,N_11570);
and U15438 (N_15438,N_12800,N_11259);
and U15439 (N_15439,N_11213,N_13218);
and U15440 (N_15440,N_10058,N_13225);
or U15441 (N_15441,N_11403,N_14527);
nand U15442 (N_15442,N_14217,N_10679);
nand U15443 (N_15443,N_10432,N_14112);
nand U15444 (N_15444,N_10721,N_12613);
xor U15445 (N_15445,N_13687,N_12645);
nor U15446 (N_15446,N_13531,N_12487);
nand U15447 (N_15447,N_12484,N_10657);
and U15448 (N_15448,N_14521,N_10617);
nand U15449 (N_15449,N_11332,N_11832);
nand U15450 (N_15450,N_12982,N_11163);
and U15451 (N_15451,N_14519,N_14655);
and U15452 (N_15452,N_11639,N_12024);
or U15453 (N_15453,N_11334,N_13286);
and U15454 (N_15454,N_14887,N_10482);
nand U15455 (N_15455,N_11760,N_14874);
nor U15456 (N_15456,N_10640,N_11823);
nand U15457 (N_15457,N_12272,N_10716);
and U15458 (N_15458,N_10734,N_10197);
xnor U15459 (N_15459,N_13359,N_11587);
or U15460 (N_15460,N_10258,N_12458);
nor U15461 (N_15461,N_13584,N_11339);
or U15462 (N_15462,N_11934,N_11310);
nor U15463 (N_15463,N_13548,N_12868);
xnor U15464 (N_15464,N_13493,N_14725);
nor U15465 (N_15465,N_12749,N_13344);
and U15466 (N_15466,N_14096,N_13814);
nor U15467 (N_15467,N_10211,N_10472);
or U15468 (N_15468,N_13736,N_13219);
nor U15469 (N_15469,N_10530,N_12759);
nor U15470 (N_15470,N_12612,N_12382);
or U15471 (N_15471,N_14644,N_10185);
or U15472 (N_15472,N_13457,N_13143);
nor U15473 (N_15473,N_13267,N_11791);
or U15474 (N_15474,N_11884,N_11704);
xnor U15475 (N_15475,N_10644,N_11737);
nand U15476 (N_15476,N_12856,N_12054);
nor U15477 (N_15477,N_14088,N_10285);
nor U15478 (N_15478,N_13412,N_12268);
nand U15479 (N_15479,N_11993,N_12158);
nor U15480 (N_15480,N_11385,N_11793);
and U15481 (N_15481,N_14078,N_12328);
xnor U15482 (N_15482,N_12504,N_12631);
xnor U15483 (N_15483,N_14226,N_10991);
nor U15484 (N_15484,N_11594,N_10460);
nor U15485 (N_15485,N_10678,N_13034);
nand U15486 (N_15486,N_14319,N_11373);
nand U15487 (N_15487,N_11482,N_13996);
nand U15488 (N_15488,N_11751,N_14688);
or U15489 (N_15489,N_13382,N_14736);
nor U15490 (N_15490,N_11452,N_13461);
nor U15491 (N_15491,N_12196,N_11451);
nor U15492 (N_15492,N_14438,N_11947);
xnor U15493 (N_15493,N_12267,N_14460);
nor U15494 (N_15494,N_14094,N_11899);
and U15495 (N_15495,N_10442,N_11538);
nor U15496 (N_15496,N_12768,N_10393);
or U15497 (N_15497,N_12422,N_10220);
or U15498 (N_15498,N_13722,N_14334);
nor U15499 (N_15499,N_11626,N_12164);
or U15500 (N_15500,N_14125,N_10114);
nor U15501 (N_15501,N_13323,N_13845);
and U15502 (N_15502,N_14137,N_10953);
xor U15503 (N_15503,N_10565,N_13393);
and U15504 (N_15504,N_14969,N_14506);
xnor U15505 (N_15505,N_13485,N_13014);
or U15506 (N_15506,N_14201,N_10882);
nand U15507 (N_15507,N_11184,N_13643);
nand U15508 (N_15508,N_11370,N_14550);
and U15509 (N_15509,N_10395,N_11199);
nor U15510 (N_15510,N_12056,N_13274);
or U15511 (N_15511,N_13694,N_10465);
nor U15512 (N_15512,N_11666,N_11917);
nor U15513 (N_15513,N_14474,N_13109);
and U15514 (N_15514,N_14282,N_12789);
nor U15515 (N_15515,N_13168,N_12564);
nand U15516 (N_15516,N_11739,N_10862);
nand U15517 (N_15517,N_10137,N_10264);
or U15518 (N_15518,N_13186,N_14170);
nor U15519 (N_15519,N_13897,N_13037);
nor U15520 (N_15520,N_13878,N_12413);
nand U15521 (N_15521,N_10199,N_11640);
or U15522 (N_15522,N_11117,N_12315);
nor U15523 (N_15523,N_12901,N_12345);
or U15524 (N_15524,N_14565,N_13659);
and U15525 (N_15525,N_14545,N_13881);
nor U15526 (N_15526,N_13424,N_12531);
nand U15527 (N_15527,N_10651,N_11900);
xor U15528 (N_15528,N_14229,N_14205);
or U15529 (N_15529,N_12673,N_12253);
nand U15530 (N_15530,N_13884,N_12990);
or U15531 (N_15531,N_13874,N_12365);
nand U15532 (N_15532,N_12931,N_12254);
and U15533 (N_15533,N_12785,N_13973);
nor U15534 (N_15534,N_13394,N_11892);
xnor U15535 (N_15535,N_13369,N_13064);
or U15536 (N_15536,N_13820,N_13342);
or U15537 (N_15537,N_10742,N_11961);
nor U15538 (N_15538,N_11733,N_13777);
nand U15539 (N_15539,N_10857,N_12427);
or U15540 (N_15540,N_10004,N_13510);
or U15541 (N_15541,N_13250,N_14661);
or U15542 (N_15542,N_10972,N_12125);
or U15543 (N_15543,N_11142,N_11515);
and U15544 (N_15544,N_11946,N_12009);
nor U15545 (N_15545,N_14393,N_13700);
or U15546 (N_15546,N_14857,N_10443);
and U15547 (N_15547,N_13911,N_10002);
or U15548 (N_15548,N_12865,N_12392);
nor U15549 (N_15549,N_12434,N_10043);
nand U15550 (N_15550,N_12942,N_10863);
nor U15551 (N_15551,N_11722,N_10771);
or U15552 (N_15552,N_12559,N_11433);
nand U15553 (N_15553,N_13355,N_11419);
nand U15554 (N_15554,N_10957,N_10557);
nor U15555 (N_15555,N_12483,N_10252);
or U15556 (N_15556,N_11342,N_14985);
or U15557 (N_15557,N_13469,N_11102);
and U15558 (N_15558,N_14697,N_12225);
or U15559 (N_15559,N_12124,N_12248);
and U15560 (N_15560,N_10080,N_13200);
nand U15561 (N_15561,N_10850,N_13385);
or U15562 (N_15562,N_11087,N_12218);
xor U15563 (N_15563,N_12755,N_12515);
or U15564 (N_15564,N_11902,N_14890);
nand U15565 (N_15565,N_12701,N_11252);
nand U15566 (N_15566,N_10917,N_14726);
and U15567 (N_15567,N_14210,N_12347);
nand U15568 (N_15568,N_11502,N_12547);
xnor U15569 (N_15569,N_14961,N_14300);
nand U15570 (N_15570,N_12553,N_13029);
nor U15571 (N_15571,N_11307,N_12037);
and U15572 (N_15572,N_13932,N_12965);
nor U15573 (N_15573,N_11471,N_12327);
or U15574 (N_15574,N_10845,N_12435);
and U15575 (N_15575,N_11811,N_13339);
nor U15576 (N_15576,N_13303,N_10547);
nand U15577 (N_15577,N_13912,N_11612);
and U15578 (N_15578,N_11416,N_11582);
xnor U15579 (N_15579,N_13770,N_12608);
nand U15580 (N_15580,N_14891,N_13811);
or U15581 (N_15581,N_10162,N_10242);
or U15582 (N_15582,N_11341,N_10323);
and U15583 (N_15583,N_12174,N_10014);
nand U15584 (N_15584,N_11525,N_11159);
and U15585 (N_15585,N_10378,N_12175);
nor U15586 (N_15586,N_13570,N_13972);
nand U15587 (N_15587,N_13333,N_11463);
nand U15588 (N_15588,N_11930,N_11329);
xor U15589 (N_15589,N_11177,N_14853);
nor U15590 (N_15590,N_14983,N_11058);
and U15591 (N_15591,N_10858,N_12096);
xor U15592 (N_15592,N_11218,N_10552);
or U15593 (N_15593,N_11192,N_14325);
and U15594 (N_15594,N_13164,N_11908);
or U15595 (N_15595,N_11077,N_14906);
xnor U15596 (N_15596,N_13578,N_12872);
and U15597 (N_15597,N_12257,N_13918);
and U15598 (N_15598,N_14314,N_14841);
or U15599 (N_15599,N_14596,N_14888);
nand U15600 (N_15600,N_11261,N_10877);
xor U15601 (N_15601,N_13935,N_12279);
and U15602 (N_15602,N_10730,N_12656);
nand U15603 (N_15603,N_11040,N_10283);
or U15604 (N_15604,N_12433,N_14133);
and U15605 (N_15605,N_12676,N_10469);
nand U15606 (N_15606,N_12679,N_14458);
xor U15607 (N_15607,N_12005,N_12008);
or U15608 (N_15608,N_11954,N_10489);
nor U15609 (N_15609,N_13887,N_14635);
nor U15610 (N_15610,N_10945,N_12727);
and U15611 (N_15611,N_14208,N_12469);
or U15612 (N_15612,N_10331,N_14979);
nand U15613 (N_15613,N_11031,N_13442);
nand U15614 (N_15614,N_13324,N_11381);
and U15615 (N_15615,N_12888,N_10373);
nor U15616 (N_15616,N_13772,N_13258);
xnor U15617 (N_15617,N_13049,N_12716);
nor U15618 (N_15618,N_13207,N_11091);
nand U15619 (N_15619,N_13721,N_12919);
nand U15620 (N_15620,N_14729,N_10822);
nor U15621 (N_15621,N_13692,N_13533);
nor U15622 (N_15622,N_14202,N_12265);
nor U15623 (N_15623,N_10946,N_13923);
nand U15624 (N_15624,N_12857,N_12649);
xor U15625 (N_15625,N_14114,N_11757);
and U15626 (N_15626,N_12536,N_12662);
and U15627 (N_15627,N_14190,N_11715);
nor U15628 (N_15628,N_12027,N_12454);
nand U15629 (N_15629,N_11953,N_13302);
and U15630 (N_15630,N_14641,N_13732);
and U15631 (N_15631,N_13970,N_14331);
and U15632 (N_15632,N_13226,N_14618);
or U15633 (N_15633,N_13971,N_14951);
nor U15634 (N_15634,N_12014,N_10458);
xnor U15635 (N_15635,N_13094,N_10447);
nand U15636 (N_15636,N_12845,N_12667);
or U15637 (N_15637,N_10391,N_14708);
xnor U15638 (N_15638,N_11874,N_10251);
xnor U15639 (N_15639,N_13301,N_14512);
or U15640 (N_15640,N_11896,N_11727);
xor U15641 (N_15641,N_14848,N_12997);
xnor U15642 (N_15642,N_13744,N_14990);
and U15643 (N_15643,N_10499,N_12194);
nand U15644 (N_15644,N_11233,N_11692);
and U15645 (N_15645,N_12792,N_12975);
or U15646 (N_15646,N_13616,N_13784);
nor U15647 (N_15647,N_12301,N_11677);
and U15648 (N_15648,N_12145,N_13890);
nor U15649 (N_15649,N_13515,N_13135);
and U15650 (N_15650,N_14602,N_14369);
and U15651 (N_15651,N_11592,N_14247);
or U15652 (N_15652,N_14907,N_10487);
or U15653 (N_15653,N_13047,N_12535);
nand U15654 (N_15654,N_13951,N_14713);
nand U15655 (N_15655,N_12855,N_14885);
and U15656 (N_15656,N_13283,N_14238);
or U15657 (N_15657,N_12123,N_13942);
or U15658 (N_15658,N_11147,N_12605);
xor U15659 (N_15659,N_10383,N_11556);
or U15660 (N_15660,N_13896,N_10569);
or U15661 (N_15661,N_11732,N_12167);
and U15662 (N_15662,N_10757,N_12366);
nor U15663 (N_15663,N_11877,N_13693);
or U15664 (N_15664,N_11568,N_12438);
nand U15665 (N_15665,N_12720,N_14919);
nand U15666 (N_15666,N_13835,N_10714);
nor U15667 (N_15667,N_11989,N_11806);
and U15668 (N_15668,N_13567,N_12862);
xnor U15669 (N_15669,N_12743,N_14821);
and U15670 (N_15670,N_12897,N_13227);
nor U15671 (N_15671,N_12620,N_10983);
nor U15672 (N_15672,N_13535,N_11945);
and U15673 (N_15673,N_11608,N_10871);
nor U15674 (N_15674,N_14379,N_13854);
nand U15675 (N_15675,N_13407,N_10115);
and U15676 (N_15676,N_14831,N_14198);
or U15677 (N_15677,N_11942,N_12491);
nand U15678 (N_15678,N_12969,N_14589);
and U15679 (N_15679,N_14442,N_12622);
or U15680 (N_15680,N_11134,N_13543);
nor U15681 (N_15681,N_11637,N_12529);
nand U15682 (N_15682,N_11609,N_11375);
nor U15683 (N_15683,N_12304,N_10927);
and U15684 (N_15684,N_12156,N_11183);
xor U15685 (N_15685,N_10590,N_11994);
and U15686 (N_15686,N_12548,N_12414);
nand U15687 (N_15687,N_13289,N_11644);
xnor U15688 (N_15688,N_10698,N_13708);
nand U15689 (N_15689,N_14102,N_11368);
nor U15690 (N_15690,N_11519,N_11027);
or U15691 (N_15691,N_13667,N_13648);
nand U15692 (N_15692,N_11411,N_10262);
and U15693 (N_15693,N_10614,N_14105);
nor U15694 (N_15694,N_13605,N_12157);
and U15695 (N_15695,N_14035,N_10732);
and U15696 (N_15696,N_14050,N_14924);
and U15697 (N_15697,N_13048,N_10121);
and U15698 (N_15698,N_12870,N_13497);
and U15699 (N_15699,N_11053,N_14850);
or U15700 (N_15700,N_11219,N_13454);
and U15701 (N_15701,N_12876,N_14680);
nand U15702 (N_15702,N_10723,N_13730);
and U15703 (N_15703,N_12788,N_10752);
nor U15704 (N_15704,N_10133,N_10783);
nand U15705 (N_15705,N_12957,N_11023);
and U15706 (N_15706,N_11730,N_11746);
and U15707 (N_15707,N_14554,N_13947);
or U15708 (N_15708,N_13193,N_14516);
nor U15709 (N_15709,N_14931,N_11313);
nand U15710 (N_15710,N_13396,N_14293);
and U15711 (N_15711,N_13417,N_11240);
nor U15712 (N_15712,N_13975,N_11819);
nand U15713 (N_15713,N_13082,N_11540);
nor U15714 (N_15714,N_13967,N_10142);
or U15715 (N_15715,N_12471,N_14016);
and U15716 (N_15716,N_14151,N_14864);
or U15717 (N_15717,N_10194,N_11798);
nand U15718 (N_15718,N_11539,N_14578);
nor U15719 (N_15719,N_12610,N_14989);
or U15720 (N_15720,N_12479,N_14194);
nand U15721 (N_15721,N_14204,N_14324);
xnor U15722 (N_15722,N_14296,N_13742);
xor U15723 (N_15723,N_14141,N_10046);
nand U15724 (N_15724,N_11010,N_11245);
xnor U15725 (N_15725,N_11173,N_11005);
or U15726 (N_15726,N_11516,N_13817);
or U15727 (N_15727,N_10294,N_12153);
nand U15728 (N_15728,N_14917,N_14337);
and U15729 (N_15729,N_12077,N_11936);
xnor U15730 (N_15730,N_11158,N_14854);
and U15731 (N_15731,N_12230,N_11931);
and U15732 (N_15732,N_11565,N_12351);
nand U15733 (N_15733,N_10794,N_11772);
nor U15734 (N_15734,N_12331,N_14904);
and U15735 (N_15735,N_12786,N_10488);
and U15736 (N_15736,N_14256,N_14760);
nand U15737 (N_15737,N_13372,N_12339);
nand U15738 (N_15738,N_13803,N_13435);
nand U15739 (N_15739,N_11718,N_11415);
or U15740 (N_15740,N_10321,N_14679);
nand U15741 (N_15741,N_14724,N_11215);
and U15742 (N_15742,N_10067,N_13711);
or U15743 (N_15743,N_11402,N_14284);
nand U15744 (N_15744,N_12114,N_12831);
nand U15745 (N_15745,N_12108,N_13198);
nand U15746 (N_15746,N_10779,N_11794);
or U15747 (N_15747,N_12001,N_10790);
or U15748 (N_15748,N_11103,N_10118);
nor U15749 (N_15749,N_10713,N_10147);
and U15750 (N_15750,N_14399,N_12117);
and U15751 (N_15751,N_14445,N_10422);
and U15752 (N_15752,N_12038,N_11000);
nor U15753 (N_15753,N_10760,N_13131);
and U15754 (N_15754,N_13789,N_14251);
nand U15755 (N_15755,N_11393,N_10146);
nor U15756 (N_15756,N_14003,N_10318);
and U15757 (N_15757,N_13994,N_11316);
and U15758 (N_15758,N_12168,N_13727);
and U15759 (N_15759,N_10597,N_14090);
or U15760 (N_15760,N_10966,N_14524);
nor U15761 (N_15761,N_12302,N_14912);
and U15762 (N_15762,N_13251,N_12146);
nand U15763 (N_15763,N_12330,N_14153);
nand U15764 (N_15764,N_12951,N_10726);
nand U15765 (N_15765,N_13558,N_12094);
or U15766 (N_15766,N_14568,N_11465);
xnor U15767 (N_15767,N_12450,N_12593);
nand U15768 (N_15768,N_12943,N_10689);
or U15769 (N_15769,N_14895,N_14373);
nor U15770 (N_15770,N_11981,N_14509);
and U15771 (N_15771,N_13574,N_13495);
nand U15772 (N_15772,N_10649,N_11258);
nor U15773 (N_15773,N_12296,N_11944);
or U15774 (N_15774,N_11109,N_11111);
and U15775 (N_15775,N_12205,N_12873);
nor U15776 (N_15776,N_12565,N_14139);
and U15777 (N_15777,N_14328,N_13169);
nand U15778 (N_15778,N_11765,N_14669);
and U15779 (N_15779,N_12967,N_14172);
nand U15780 (N_15780,N_14405,N_12907);
nor U15781 (N_15781,N_12030,N_13326);
nor U15782 (N_15782,N_12359,N_14239);
nor U15783 (N_15783,N_14066,N_12073);
or U15784 (N_15784,N_12820,N_14860);
or U15785 (N_15785,N_11302,N_13276);
nor U15786 (N_15786,N_12340,N_12754);
and U15787 (N_15787,N_13740,N_12546);
or U15788 (N_15788,N_14930,N_10225);
or U15789 (N_15789,N_12280,N_11595);
and U15790 (N_15790,N_12651,N_11446);
nor U15791 (N_15791,N_11822,N_13126);
and U15792 (N_15792,N_14617,N_14690);
nand U15793 (N_15793,N_10428,N_11277);
and U15794 (N_15794,N_10269,N_12805);
nand U15795 (N_15795,N_13672,N_13174);
and U15796 (N_15796,N_13801,N_11216);
or U15797 (N_15797,N_13812,N_14714);
nor U15798 (N_15798,N_11141,N_12376);
and U15799 (N_15799,N_11286,N_11466);
xor U15800 (N_15800,N_13091,N_14666);
and U15801 (N_15801,N_13819,N_14175);
nor U15802 (N_15802,N_12459,N_13432);
nor U15803 (N_15803,N_13880,N_14345);
or U15804 (N_15804,N_10645,N_10491);
nor U15805 (N_15805,N_14815,N_11484);
or U15806 (N_15806,N_10886,N_10117);
or U15807 (N_15807,N_13824,N_14704);
nor U15808 (N_15808,N_12432,N_10345);
xor U15809 (N_15809,N_14146,N_11789);
nor U15810 (N_15810,N_12204,N_13422);
nor U15811 (N_15811,N_10222,N_13356);
nand U15812 (N_15812,N_11443,N_13057);
nand U15813 (N_15813,N_11802,N_12763);
and U15814 (N_15814,N_11095,N_10191);
xor U15815 (N_15815,N_13886,N_11160);
nor U15816 (N_15816,N_12428,N_14123);
or U15817 (N_15817,N_11940,N_13146);
nor U15818 (N_15818,N_14605,N_13121);
xor U15819 (N_15819,N_14375,N_10380);
and U15820 (N_15820,N_14761,N_14789);
and U15821 (N_15821,N_12717,N_10329);
nor U15822 (N_15822,N_10056,N_14462);
or U15823 (N_15823,N_11176,N_14628);
nand U15824 (N_15824,N_10610,N_12136);
xnor U15825 (N_15825,N_10607,N_11022);
and U15826 (N_15826,N_11133,N_12187);
or U15827 (N_15827,N_14044,N_12349);
nor U15828 (N_15828,N_13800,N_13089);
and U15829 (N_15829,N_13409,N_11964);
and U15830 (N_15830,N_12138,N_12658);
and U15831 (N_15831,N_13428,N_13260);
nor U15832 (N_15832,N_13941,N_11044);
xnor U15833 (N_15833,N_12243,N_12088);
or U15834 (N_15834,N_14196,N_12830);
or U15835 (N_15835,N_12971,N_10159);
or U15836 (N_15836,N_12955,N_11267);
and U15837 (N_15837,N_10410,N_12766);
nand U15838 (N_15838,N_11581,N_12906);
or U15839 (N_15839,N_10843,N_14091);
nor U15840 (N_15840,N_13102,N_13313);
nand U15841 (N_15841,N_10122,N_12537);
xnor U15842 (N_15842,N_11904,N_10762);
or U15843 (N_15843,N_13395,N_13242);
and U15844 (N_15844,N_12250,N_11231);
and U15845 (N_15845,N_10084,N_10213);
nor U15846 (N_15846,N_11729,N_13527);
nor U15847 (N_15847,N_14338,N_12641);
or U15848 (N_15848,N_14006,N_14775);
and U15849 (N_15849,N_13463,N_13843);
or U15850 (N_15850,N_10140,N_11992);
nand U15851 (N_15851,N_13928,N_10736);
and U15852 (N_15852,N_12311,N_13078);
nand U15853 (N_15853,N_10219,N_14501);
nor U15854 (N_15854,N_13892,N_14467);
and U15855 (N_15855,N_13456,N_11501);
or U15856 (N_15856,N_14476,N_10161);
or U15857 (N_15857,N_11591,N_11836);
nor U15858 (N_15858,N_14406,N_12738);
or U15859 (N_15859,N_12541,N_11898);
or U15860 (N_15860,N_14469,N_14692);
nor U15861 (N_15861,N_14898,N_12934);
nand U15862 (N_15862,N_10635,N_10038);
or U15863 (N_15863,N_10233,N_10588);
nor U15864 (N_15864,N_13621,N_14313);
and U15865 (N_15865,N_14185,N_11654);
or U15866 (N_15866,N_13610,N_11305);
nand U15867 (N_15867,N_11824,N_10746);
nand U15868 (N_15868,N_12105,N_10151);
or U15869 (N_15869,N_14942,N_10943);
or U15870 (N_15870,N_14015,N_12329);
nor U15871 (N_15871,N_11071,N_10680);
nor U15872 (N_15872,N_14743,N_12173);
nor U15873 (N_15873,N_10755,N_10388);
nand U15874 (N_15874,N_14052,N_10920);
and U15875 (N_15875,N_11457,N_14993);
nor U15876 (N_15876,N_13829,N_13560);
and U15877 (N_15877,N_14478,N_13446);
and U15878 (N_15878,N_14757,N_13483);
or U15879 (N_15879,N_12815,N_13747);
or U15880 (N_15880,N_11721,N_10377);
nand U15881 (N_15881,N_10659,N_14557);
and U15882 (N_15882,N_14177,N_12072);
or U15883 (N_15883,N_10425,N_12625);
or U15884 (N_15884,N_14774,N_10400);
and U15885 (N_15885,N_11985,N_14200);
nand U15886 (N_15886,N_14975,N_11291);
or U15887 (N_15887,N_12927,N_13999);
nand U15888 (N_15888,N_10525,N_13150);
nor U15889 (N_15889,N_11317,N_12829);
or U15890 (N_15890,N_11195,N_13715);
or U15891 (N_15891,N_13371,N_11668);
and U15892 (N_15892,N_10888,N_12476);
nand U15893 (N_15893,N_10065,N_11524);
nand U15894 (N_15894,N_11182,N_13005);
or U15895 (N_15895,N_10915,N_12291);
and U15896 (N_15896,N_10001,N_14425);
nand U15897 (N_15897,N_11113,N_11939);
nor U15898 (N_15898,N_10894,N_11299);
nand U15899 (N_15899,N_13476,N_11207);
nor U15900 (N_15900,N_12199,N_11672);
and U15901 (N_15901,N_11527,N_10579);
nor U15902 (N_15902,N_12913,N_10263);
or U15903 (N_15903,N_11846,N_13297);
nor U15904 (N_15904,N_10559,N_11999);
nand U15905 (N_15905,N_11051,N_12356);
nor U15906 (N_15906,N_12387,N_13726);
nand U15907 (N_15907,N_11167,N_13240);
or U15908 (N_15908,N_10444,N_11175);
or U15909 (N_15909,N_14357,N_13794);
nor U15910 (N_15910,N_12215,N_10348);
nor U15911 (N_15911,N_12611,N_12650);
xnor U15912 (N_15912,N_10315,N_14218);
or U15913 (N_15913,N_13604,N_12674);
nand U15914 (N_15914,N_11104,N_11275);
and U15915 (N_15915,N_14385,N_10533);
and U15916 (N_15916,N_10618,N_13921);
nor U15917 (N_15917,N_10193,N_14459);
or U15918 (N_15918,N_14927,N_12391);
nand U15919 (N_15919,N_10349,N_12543);
or U15920 (N_15920,N_14659,N_14418);
and U15921 (N_15921,N_13241,N_10270);
and U15922 (N_15922,N_10824,N_12956);
nand U15923 (N_15923,N_11713,N_14709);
or U15924 (N_15924,N_13452,N_11497);
and U15925 (N_15925,N_14386,N_13127);
and U15926 (N_15926,N_12061,N_13234);
nand U15927 (N_15927,N_11340,N_13635);
and U15928 (N_15928,N_13906,N_14308);
or U15929 (N_15929,N_14130,N_11839);
or U15930 (N_15930,N_10089,N_13011);
or U15931 (N_15931,N_10573,N_10699);
nand U15932 (N_15932,N_11242,N_11919);
xor U15933 (N_15933,N_12861,N_13095);
or U15934 (N_15934,N_11688,N_12343);
nand U15935 (N_15935,N_11922,N_12015);
and U15936 (N_15936,N_14918,N_10231);
nand U15937 (N_15937,N_14954,N_12322);
nor U15938 (N_15938,N_14808,N_11234);
or U15939 (N_15939,N_12807,N_14981);
nor U15940 (N_15940,N_11563,N_13053);
nor U15941 (N_15941,N_10516,N_13172);
nor U15942 (N_15942,N_14681,N_12892);
or U15943 (N_15943,N_12828,N_12151);
nand U15944 (N_15944,N_13035,N_14823);
nand U15945 (N_15945,N_11244,N_14950);
xnor U15946 (N_15946,N_10849,N_10996);
or U15947 (N_15947,N_14372,N_10586);
and U15948 (N_15948,N_11315,N_12497);
nand U15949 (N_15949,N_12406,N_13837);
and U15950 (N_15950,N_13006,N_13114);
nor U15951 (N_15951,N_14179,N_14311);
or U15952 (N_15952,N_10906,N_12290);
xor U15953 (N_15953,N_13786,N_10094);
or U15954 (N_15954,N_12236,N_14246);
nor U15955 (N_15955,N_11548,N_11588);
and U15956 (N_15956,N_11555,N_12465);
xnor U15957 (N_15957,N_13223,N_12635);
or U15958 (N_15958,N_14652,N_11632);
nand U15959 (N_15959,N_14209,N_12455);
or U15960 (N_15960,N_13891,N_12019);
and U15961 (N_15961,N_11646,N_11545);
or U15962 (N_15962,N_13215,N_12200);
nand U15963 (N_15963,N_14144,N_11185);
and U15964 (N_15964,N_11521,N_12796);
and U15965 (N_15965,N_13676,N_10087);
and U15966 (N_15966,N_14693,N_10807);
nand U15967 (N_15967,N_14128,N_14640);
xnor U15968 (N_15968,N_11965,N_10113);
xnor U15969 (N_15969,N_11272,N_11629);
xor U15970 (N_15970,N_10560,N_10503);
nor U15971 (N_15971,N_10013,N_14684);
and U15972 (N_15972,N_10431,N_11144);
or U15973 (N_15973,N_10008,N_10515);
and U15974 (N_15974,N_10696,N_12131);
xnor U15975 (N_15975,N_10669,N_13413);
nor U15976 (N_15976,N_14214,N_12238);
or U15977 (N_15977,N_14036,N_12372);
xnor U15978 (N_15978,N_14193,N_11198);
nand U15979 (N_15979,N_10132,N_14082);
or U15980 (N_15980,N_11880,N_11225);
nand U15981 (N_15981,N_11374,N_14054);
and U15982 (N_15982,N_14657,N_11752);
nor U15983 (N_15983,N_12878,N_14019);
xnor U15984 (N_15984,N_14601,N_12973);
and U15985 (N_15985,N_10660,N_13960);
nor U15986 (N_15986,N_12573,N_14336);
nand U15987 (N_15987,N_10234,N_13834);
nor U15988 (N_15988,N_11875,N_13861);
nor U15989 (N_15989,N_12630,N_12357);
xnor U15990 (N_15990,N_13166,N_13178);
nand U15991 (N_15991,N_11303,N_14258);
nand U15992 (N_15992,N_10608,N_10932);
nand U15993 (N_15993,N_10685,N_14923);
or U15994 (N_15994,N_14797,N_14913);
nor U15995 (N_15995,N_11014,N_14570);
and U15996 (N_15996,N_14909,N_10707);
nand U15997 (N_15997,N_13427,N_14525);
nor U15998 (N_15998,N_12691,N_10880);
nand U15999 (N_15999,N_10667,N_12937);
nor U16000 (N_16000,N_11506,N_12684);
nor U16001 (N_16001,N_12006,N_13028);
and U16002 (N_16002,N_13783,N_13282);
or U16003 (N_16003,N_12811,N_10027);
nand U16004 (N_16004,N_11361,N_11250);
and U16005 (N_16005,N_14606,N_14366);
and U16006 (N_16006,N_11057,N_13607);
or U16007 (N_16007,N_12980,N_13187);
nand U16008 (N_16008,N_14877,N_13099);
nor U16009 (N_16009,N_12832,N_14541);
and U16010 (N_16010,N_11298,N_13608);
xor U16011 (N_16011,N_13956,N_13136);
xor U16012 (N_16012,N_12394,N_14409);
nor U16013 (N_16013,N_11155,N_13927);
nor U16014 (N_16014,N_12380,N_11223);
or U16015 (N_16015,N_12985,N_14489);
and U16016 (N_16016,N_11702,N_14178);
nand U16017 (N_16017,N_14518,N_10931);
or U16018 (N_16018,N_14818,N_12777);
nor U16019 (N_16019,N_10338,N_13952);
xor U16020 (N_16020,N_13980,N_11838);
xor U16021 (N_16021,N_13025,N_13455);
and U16022 (N_16022,N_10684,N_10476);
nand U16023 (N_16023,N_11074,N_10653);
nand U16024 (N_16024,N_13380,N_14028);
xor U16025 (N_16025,N_12784,N_14443);
nor U16026 (N_16026,N_14363,N_12619);
or U16027 (N_16027,N_11178,N_12057);
nor U16028 (N_16028,N_10918,N_11808);
and U16029 (N_16029,N_10160,N_14976);
nand U16030 (N_16030,N_13113,N_10356);
xnor U16031 (N_16031,N_10138,N_13522);
xnor U16032 (N_16032,N_13966,N_11514);
nor U16033 (N_16033,N_11204,N_14482);
nand U16034 (N_16034,N_13177,N_10671);
xnor U16035 (N_16035,N_11674,N_11032);
and U16036 (N_16036,N_14633,N_12519);
or U16037 (N_16037,N_13839,N_13467);
xor U16038 (N_16038,N_14410,N_13020);
nand U16039 (N_16039,N_11755,N_14368);
nor U16040 (N_16040,N_14145,N_13987);
nor U16041 (N_16041,N_13618,N_14491);
nand U16042 (N_16042,N_10830,N_11856);
and U16043 (N_16043,N_13196,N_10717);
nor U16044 (N_16044,N_11828,N_12947);
xor U16045 (N_16045,N_12765,N_12473);
or U16046 (N_16046,N_13489,N_13595);
and U16047 (N_16047,N_11835,N_14588);
and U16048 (N_16048,N_10279,N_14672);
and U16049 (N_16049,N_11651,N_14608);
xor U16050 (N_16050,N_11882,N_14870);
and U16051 (N_16051,N_14475,N_12522);
or U16052 (N_16052,N_13449,N_10041);
nand U16053 (N_16053,N_11038,N_11598);
nor U16054 (N_16054,N_14424,N_12084);
xnor U16055 (N_16055,N_12409,N_13167);
and U16056 (N_16056,N_13259,N_11362);
nor U16057 (N_16057,N_13363,N_12154);
xor U16058 (N_16058,N_12467,N_12211);
or U16059 (N_16059,N_10037,N_14343);
nand U16060 (N_16060,N_11391,N_11975);
and U16061 (N_16061,N_12002,N_10866);
and U16062 (N_16062,N_10415,N_11863);
nand U16063 (N_16063,N_13411,N_12721);
nor U16064 (N_16064,N_14727,N_11283);
and U16065 (N_16065,N_11321,N_10119);
or U16066 (N_16066,N_11309,N_14925);
and U16067 (N_16067,N_12261,N_13275);
or U16068 (N_16068,N_13760,N_14157);
nor U16069 (N_16069,N_11437,N_13261);
nor U16070 (N_16070,N_11387,N_10099);
or U16071 (N_16071,N_13086,N_10768);
and U16072 (N_16072,N_13059,N_13745);
xnor U16073 (N_16073,N_11055,N_11870);
and U16074 (N_16074,N_10544,N_10414);
or U16075 (N_16075,N_11817,N_14093);
and U16076 (N_16076,N_11820,N_11352);
nor U16077 (N_16077,N_10390,N_10289);
nand U16078 (N_16078,N_14582,N_13270);
or U16079 (N_16079,N_11599,N_11504);
and U16080 (N_16080,N_11601,N_11395);
and U16081 (N_16081,N_10950,N_13357);
xnor U16082 (N_16082,N_13725,N_13249);
nand U16083 (N_16083,N_13741,N_11785);
or U16084 (N_16084,N_14594,N_12699);
nor U16085 (N_16085,N_10641,N_11312);
nor U16086 (N_16086,N_12127,N_10958);
and U16087 (N_16087,N_11456,N_11201);
nand U16088 (N_16088,N_12902,N_14294);
and U16089 (N_16089,N_13068,N_13306);
and U16090 (N_16090,N_13609,N_12953);
nor U16091 (N_16091,N_14786,N_12180);
nor U16092 (N_16092,N_11720,N_13899);
or U16093 (N_16093,N_10471,N_14717);
nor U16094 (N_16094,N_14945,N_10360);
nand U16095 (N_16095,N_12051,N_14929);
and U16096 (N_16096,N_12163,N_10181);
or U16097 (N_16097,N_13662,N_11887);
and U16098 (N_16098,N_12589,N_10589);
nor U16099 (N_16099,N_13516,N_11991);
or U16100 (N_16100,N_14086,N_11146);
nor U16101 (N_16101,N_10860,N_12115);
and U16102 (N_16102,N_14622,N_14173);
nand U16103 (N_16103,N_10498,N_14656);
or U16104 (N_16104,N_12133,N_10724);
or U16105 (N_16105,N_10799,N_11671);
xnor U16106 (N_16106,N_10093,N_12431);
nor U16107 (N_16107,N_10483,N_10567);
or U16108 (N_16108,N_13111,N_10047);
nor U16109 (N_16109,N_14769,N_12029);
or U16110 (N_16110,N_10326,N_11422);
or U16111 (N_16111,N_10036,N_12398);
and U16112 (N_16112,N_14441,N_10521);
or U16113 (N_16113,N_14119,N_11567);
or U16114 (N_16114,N_10741,N_12137);
nor U16115 (N_16115,N_13677,N_12500);
nand U16116 (N_16116,N_13322,N_12686);
nor U16117 (N_16117,N_12866,N_10009);
and U16118 (N_16118,N_11624,N_11168);
nand U16119 (N_16119,N_14312,N_11025);
nor U16120 (N_16120,N_10923,N_11827);
nor U16121 (N_16121,N_12640,N_11068);
or U16122 (N_16122,N_13314,N_11293);
nor U16123 (N_16123,N_12232,N_12419);
nor U16124 (N_16124,N_10273,N_14025);
nor U16125 (N_16125,N_11406,N_13257);
and U16126 (N_16126,N_12445,N_12016);
nand U16127 (N_16127,N_10619,N_14517);
nor U16128 (N_16128,N_13450,N_10885);
xnor U16129 (N_16129,N_10743,N_12884);
or U16130 (N_16130,N_14271,N_13191);
nand U16131 (N_16131,N_13623,N_10791);
or U16132 (N_16132,N_14829,N_13591);
nand U16133 (N_16133,N_11600,N_10613);
and U16134 (N_16134,N_11695,N_12582);
and U16135 (N_16135,N_10291,N_11398);
nand U16136 (N_16136,N_11363,N_12569);
and U16137 (N_16137,N_12512,N_13577);
and U16138 (N_16138,N_10352,N_14257);
and U16139 (N_16139,N_13914,N_11660);
nor U16140 (N_16140,N_13889,N_13502);
nand U16141 (N_16141,N_14297,N_14477);
nand U16142 (N_16142,N_14061,N_11933);
nor U16143 (N_16143,N_13045,N_11017);
or U16144 (N_16144,N_10778,N_12182);
nand U16145 (N_16145,N_11394,N_11617);
nor U16146 (N_16146,N_14897,N_14593);
or U16147 (N_16147,N_11082,N_14856);
nor U16148 (N_16148,N_14342,N_14621);
or U16149 (N_16149,N_14737,N_12139);
or U16150 (N_16150,N_11694,N_10852);
or U16151 (N_16151,N_13365,N_11115);
nor U16152 (N_16152,N_14673,N_11783);
nand U16153 (N_16153,N_11531,N_10928);
and U16154 (N_16154,N_14543,N_10551);
nor U16155 (N_16155,N_13565,N_12551);
nand U16156 (N_16156,N_14110,N_13400);
and U16157 (N_16157,N_10000,N_13697);
nor U16158 (N_16158,N_12481,N_10949);
and U16159 (N_16159,N_10284,N_12813);
or U16160 (N_16160,N_12020,N_10606);
xor U16161 (N_16161,N_10944,N_12179);
nand U16162 (N_16162,N_14626,N_14046);
xnor U16163 (N_16163,N_13879,N_14496);
nand U16164 (N_16164,N_12659,N_12165);
nand U16165 (N_16165,N_14455,N_11744);
and U16166 (N_16166,N_13597,N_14488);
nor U16167 (N_16167,N_10238,N_12606);
nor U16168 (N_16168,N_12335,N_14274);
nor U16169 (N_16169,N_12033,N_13151);
xor U16170 (N_16170,N_13023,N_12436);
nor U16171 (N_16171,N_13924,N_10786);
and U16172 (N_16172,N_14533,N_10050);
and U16173 (N_16173,N_10459,N_14852);
and U16174 (N_16174,N_13468,N_14551);
nand U16175 (N_16175,N_13236,N_12881);
or U16176 (N_16176,N_10910,N_12287);
nor U16177 (N_16177,N_13293,N_10246);
and U16178 (N_16178,N_12838,N_11825);
or U16179 (N_16179,N_12134,N_10421);
and U16180 (N_16180,N_12827,N_10186);
and U16181 (N_16181,N_14710,N_13317);
and U16182 (N_16182,N_10965,N_12444);
and U16183 (N_16183,N_11351,N_14479);
nor U16184 (N_16184,N_11518,N_14862);
and U16185 (N_16185,N_11432,N_13501);
nand U16186 (N_16186,N_12713,N_13147);
nor U16187 (N_16187,N_13561,N_10022);
nor U16188 (N_16188,N_11099,N_12183);
nand U16189 (N_16189,N_13653,N_13229);
or U16190 (N_16190,N_13766,N_14083);
and U16191 (N_16191,N_14699,N_13707);
nor U16192 (N_16192,N_12687,N_14920);
nor U16193 (N_16193,N_13401,N_10303);
and U16194 (N_16194,N_13279,N_14184);
and U16195 (N_16195,N_11800,N_10859);
and U16196 (N_16196,N_12863,N_10639);
nor U16197 (N_16197,N_11630,N_14546);
or U16198 (N_16198,N_11166,N_13195);
nand U16199 (N_16199,N_11636,N_14248);
nor U16200 (N_16200,N_10837,N_12067);
nor U16201 (N_16201,N_10744,N_12050);
nor U16202 (N_16202,N_13060,N_12886);
nor U16203 (N_16203,N_11682,N_11006);
nor U16204 (N_16204,N_11280,N_12049);
nand U16205 (N_16205,N_14740,N_11382);
and U16206 (N_16206,N_10759,N_11429);
nor U16207 (N_16207,N_11706,N_13273);
nor U16208 (N_16208,N_11100,N_13431);
or U16209 (N_16209,N_12472,N_13278);
and U16210 (N_16210,N_11513,N_11011);
nor U16211 (N_16211,N_14896,N_14722);
and U16212 (N_16212,N_12229,N_10535);
xnor U16213 (N_16213,N_13670,N_14361);
and U16214 (N_16214,N_13828,N_11123);
nand U16215 (N_16215,N_12652,N_13804);
and U16216 (N_16216,N_13534,N_12966);
or U16217 (N_16217,N_11575,N_13349);
or U16218 (N_16218,N_10209,N_10780);
nor U16219 (N_16219,N_11171,N_10343);
or U16220 (N_16220,N_10149,N_14236);
and U16221 (N_16221,N_14905,N_10555);
nor U16222 (N_16222,N_11543,N_14374);
and U16223 (N_16223,N_10844,N_14303);
and U16224 (N_16224,N_14835,N_11648);
xnor U16225 (N_16225,N_11464,N_14129);
or U16226 (N_16226,N_13119,N_11956);
or U16227 (N_16227,N_10835,N_11458);
or U16228 (N_16228,N_12607,N_13364);
and U16229 (N_16229,N_11205,N_14728);
and U16230 (N_16230,N_12690,N_13155);
or U16231 (N_16231,N_11621,N_12011);
nor U16232 (N_16232,N_10509,N_10861);
nand U16233 (N_16233,N_14531,N_13576);
or U16234 (N_16234,N_13124,N_14234);
and U16235 (N_16235,N_13197,N_12017);
nor U16236 (N_16236,N_12632,N_14365);
xnor U16237 (N_16237,N_10585,N_13866);
or U16238 (N_16238,N_14383,N_14801);
or U16239 (N_16239,N_14428,N_11530);
nand U16240 (N_16240,N_14421,N_12122);
and U16241 (N_16241,N_14928,N_13626);
or U16242 (N_16242,N_13399,N_11627);
nor U16243 (N_16243,N_12231,N_14738);
nand U16244 (N_16244,N_14796,N_11921);
nand U16245 (N_16245,N_11399,N_10819);
and U16246 (N_16246,N_14156,N_12485);
or U16247 (N_16247,N_10367,N_14212);
nand U16248 (N_16248,N_14408,N_11913);
nor U16249 (N_16249,N_10887,N_10890);
and U16250 (N_16250,N_11285,N_13329);
or U16251 (N_16251,N_11132,N_12032);
xnor U16252 (N_16252,N_11358,N_13564);
nor U16253 (N_16253,N_14344,N_14563);
nand U16254 (N_16254,N_10838,N_14514);
and U16255 (N_16255,N_11998,N_13327);
xor U16256 (N_16256,N_11487,N_14572);
xnor U16257 (N_16257,N_13157,N_10496);
nor U16258 (N_16258,N_13308,N_13954);
and U16259 (N_16259,N_12140,N_10490);
and U16260 (N_16260,N_14609,N_12377);
and U16261 (N_16261,N_12542,N_12511);
nor U16262 (N_16262,N_14547,N_13105);
or U16263 (N_16263,N_11740,N_10207);
nand U16264 (N_16264,N_14384,N_12555);
or U16265 (N_16265,N_10709,N_12926);
nand U16266 (N_16266,N_14782,N_13673);
and U16267 (N_16267,N_13351,N_12848);
nor U16268 (N_16268,N_14431,N_12760);
nor U16269 (N_16269,N_11769,N_13209);
nand U16270 (N_16270,N_14836,N_10392);
or U16271 (N_16271,N_13986,N_10300);
xnor U16272 (N_16272,N_13335,N_11152);
nand U16273 (N_16273,N_13554,N_12824);
nand U16274 (N_16274,N_10672,N_12521);
and U16275 (N_16275,N_10553,N_10077);
nand U16276 (N_16276,N_14322,N_11876);
xor U16277 (N_16277,N_13244,N_12594);
or U16278 (N_16278,N_11379,N_12806);
nand U16279 (N_16279,N_13658,N_12341);
nor U16280 (N_16280,N_12954,N_11449);
or U16281 (N_16281,N_14370,N_13040);
or U16282 (N_16282,N_14207,N_12949);
nand U16283 (N_16283,N_12981,N_12941);
or U16284 (N_16284,N_14707,N_13085);
and U16285 (N_16285,N_14564,N_10086);
and U16286 (N_16286,N_12234,N_12303);
nor U16287 (N_16287,N_13039,N_13815);
or U16288 (N_16288,N_13204,N_10600);
nor U16289 (N_16289,N_12634,N_13444);
xnor U16290 (N_16290,N_13579,N_14846);
and U16291 (N_16291,N_14387,N_14646);
xnor U16292 (N_16292,N_10839,N_13305);
or U16293 (N_16293,N_13067,N_12142);
and U16294 (N_16294,N_11812,N_11453);
nand U16295 (N_16295,N_12787,N_14691);
nor U16296 (N_16296,N_13097,N_13062);
or U16297 (N_16297,N_12169,N_12665);
and U16298 (N_16298,N_13066,N_11019);
and U16299 (N_16299,N_12928,N_12826);
nor U16300 (N_16300,N_14992,N_13894);
nand U16301 (N_16301,N_13642,N_13464);
nand U16302 (N_16302,N_14875,N_13004);
or U16303 (N_16303,N_14651,N_10683);
nand U16304 (N_16304,N_11327,N_10467);
and U16305 (N_16305,N_11988,N_12728);
or U16306 (N_16306,N_14817,N_10055);
nand U16307 (N_16307,N_10486,N_11978);
or U16308 (N_16308,N_13706,N_11857);
or U16309 (N_16309,N_14352,N_14349);
and U16310 (N_16310,N_12821,N_11736);
or U16311 (N_16311,N_12940,N_11221);
or U16312 (N_16312,N_10522,N_13519);
nor U16313 (N_16313,N_10076,N_12363);
and U16314 (N_16314,N_14059,N_13352);
nor U16315 (N_16315,N_11698,N_12354);
nand U16316 (N_16316,N_14664,N_10998);
or U16317 (N_16317,N_14235,N_12440);
nor U16318 (N_16318,N_10633,N_11486);
nor U16319 (N_16319,N_11905,N_13499);
nand U16320 (N_16320,N_11509,N_12793);
nor U16321 (N_16321,N_11918,N_11045);
xor U16322 (N_16322,N_12781,N_13210);
or U16323 (N_16323,N_12725,N_10952);
and U16324 (N_16324,N_14576,N_11337);
or U16325 (N_16325,N_14508,N_14982);
nor U16326 (N_16326,N_14397,N_13309);
and U16327 (N_16327,N_13362,N_13496);
nand U16328 (N_16328,N_13537,N_12369);
and U16329 (N_16329,N_11748,N_13838);
or U16330 (N_16330,N_11522,N_11645);
nor U16331 (N_16331,N_14803,N_11193);
nand U16332 (N_16332,N_14270,N_12557);
or U16333 (N_16333,N_11371,N_10473);
and U16334 (N_16334,N_12278,N_14581);
or U16335 (N_16335,N_10292,N_14994);
nand U16336 (N_16336,N_14403,N_13850);
or U16337 (N_16337,N_11150,N_10896);
nand U16338 (N_16338,N_10416,N_10248);
and U16339 (N_16339,N_13341,N_13729);
or U16340 (N_16340,N_11661,N_13655);
and U16341 (N_16341,N_11349,N_10554);
or U16342 (N_16342,N_11553,N_14882);
xnor U16343 (N_16343,N_13514,N_13684);
or U16344 (N_16344,N_14162,N_11747);
and U16345 (N_16345,N_10420,N_10130);
xnor U16346 (N_16346,N_13795,N_10761);
nor U16347 (N_16347,N_11357,N_14537);
or U16348 (N_16348,N_14329,N_11890);
nor U16349 (N_16349,N_11472,N_11072);
nand U16350 (N_16350,N_13539,N_14631);
and U16351 (N_16351,N_14649,N_12352);
xnor U16352 (N_16352,N_14886,N_11843);
and U16353 (N_16353,N_14330,N_13139);
nand U16354 (N_16354,N_10053,N_12771);
or U16355 (N_16355,N_11920,N_12526);
or U16356 (N_16356,N_14826,N_13827);
and U16357 (N_16357,N_11888,N_10772);
nor U16358 (N_16358,N_12442,N_11474);
and U16359 (N_16359,N_14499,N_11816);
or U16360 (N_16360,N_14977,N_11481);
nor U16361 (N_16361,N_10527,N_11401);
and U16362 (N_16362,N_12808,N_11826);
nor U16363 (N_16363,N_12150,N_11728);
and U16364 (N_16364,N_11508,N_14453);
and U16365 (N_16365,N_12925,N_13796);
nand U16366 (N_16366,N_11235,N_10363);
and U16367 (N_16367,N_11383,N_14685);
nand U16368 (N_16368,N_14480,N_14963);
or U16369 (N_16369,N_11054,N_10030);
xnor U16370 (N_16370,N_13699,N_14607);
or U16371 (N_16371,N_12797,N_14530);
xor U16372 (N_16372,N_12524,N_14223);
nand U16373 (N_16373,N_13787,N_13683);
xor U16374 (N_16374,N_13586,N_11041);
and U16375 (N_16375,N_10568,N_12289);
nor U16376 (N_16376,N_10987,N_11420);
or U16377 (N_16377,N_14452,N_13929);
nor U16378 (N_16378,N_11444,N_14549);
or U16379 (N_16379,N_14705,N_14287);
nand U16380 (N_16380,N_13019,N_12681);
nand U16381 (N_16381,N_10956,N_12264);
or U16382 (N_16382,N_12081,N_14505);
nor U16383 (N_16383,N_13140,N_13158);
xnor U16384 (N_16384,N_11593,N_13998);
nand U16385 (N_16385,N_14949,N_14776);
nor U16386 (N_16386,N_11680,N_13737);
nor U16387 (N_16387,N_11450,N_14999);
or U16388 (N_16388,N_10335,N_11311);
and U16389 (N_16389,N_13402,N_10545);
nor U16390 (N_16390,N_14301,N_13559);
nand U16391 (N_16391,N_11069,N_14304);
nor U16392 (N_16392,N_11925,N_11021);
and U16393 (N_16393,N_11035,N_10959);
or U16394 (N_16394,N_12012,N_14536);
and U16395 (N_16395,N_13530,N_14049);
nor U16396 (N_16396,N_10514,N_10229);
or U16397 (N_16397,N_14394,N_11719);
nor U16398 (N_16398,N_14932,N_14008);
or U16399 (N_16399,N_14490,N_13917);
nand U16400 (N_16400,N_12295,N_12285);
and U16401 (N_16401,N_14069,N_10978);
nand U16402 (N_16402,N_14401,N_10939);
and U16403 (N_16403,N_12963,N_11724);
nand U16404 (N_16404,N_11771,N_13681);
nor U16405 (N_16405,N_11924,N_10908);
and U16406 (N_16406,N_13055,N_12320);
or U16407 (N_16407,N_10454,N_14186);
nor U16408 (N_16408,N_12750,N_14665);
or U16409 (N_16409,N_11408,N_12891);
and U16410 (N_16410,N_11664,N_10594);
nor U16411 (N_16411,N_11523,N_10310);
or U16412 (N_16412,N_12042,N_10327);
nand U16413 (N_16413,N_10930,N_10789);
or U16414 (N_16414,N_12922,N_11505);
and U16415 (N_16415,N_12065,N_10223);
and U16416 (N_16416,N_11322,N_11937);
and U16417 (N_16417,N_14584,N_12617);
nor U16418 (N_16418,N_13436,N_14295);
and U16419 (N_16419,N_12566,N_14806);
nand U16420 (N_16420,N_10354,N_14768);
nor U16421 (N_16421,N_11955,N_13441);
nand U16422 (N_16422,N_13752,N_14636);
nand U16423 (N_16423,N_13336,N_13536);
and U16424 (N_16424,N_10655,N_14211);
nor U16425 (N_16425,N_12109,N_10249);
and U16426 (N_16426,N_11190,N_12309);
nor U16427 (N_16427,N_11421,N_12429);
nand U16428 (N_16428,N_12602,N_11354);
xor U16429 (N_16429,N_10942,N_12887);
nor U16430 (N_16430,N_13903,N_11089);
xnor U16431 (N_16431,N_11318,N_12397);
nor U16432 (N_16432,N_13682,N_12141);
and U16433 (N_16433,N_10750,N_11952);
nor U16434 (N_16434,N_10074,N_10773);
or U16435 (N_16435,N_11842,N_12477);
nor U16436 (N_16436,N_12336,N_10401);
nand U16437 (N_16437,N_10276,N_14152);
or U16438 (N_16438,N_13594,N_14731);
xor U16439 (N_16439,N_12914,N_12995);
and U16440 (N_16440,N_11170,N_14956);
xor U16441 (N_16441,N_12653,N_10028);
and U16442 (N_16442,N_11603,N_12147);
and U16443 (N_16443,N_13491,N_13521);
xor U16444 (N_16444,N_11197,N_11356);
nor U16445 (N_16445,N_10253,N_13083);
xor U16446 (N_16446,N_11413,N_14468);
nor U16447 (N_16447,N_14783,N_13384);
nor U16448 (N_16448,N_11288,N_12100);
and U16449 (N_16449,N_14377,N_14389);
or U16450 (N_16450,N_14017,N_11191);
and U16451 (N_16451,N_11738,N_10237);
nand U16452 (N_16452,N_10938,N_14451);
xor U16453 (N_16453,N_14463,N_10484);
or U16454 (N_16454,N_13985,N_13634);
nand U16455 (N_16455,N_10735,N_10929);
nand U16456 (N_16456,N_11776,N_11319);
nand U16457 (N_16457,N_13018,N_10519);
nor U16458 (N_16458,N_11033,N_10096);
or U16459 (N_16459,N_12670,N_11209);
nor U16460 (N_16460,N_11669,N_11766);
nand U16461 (N_16461,N_10305,N_10825);
nand U16462 (N_16462,N_13862,N_12402);
nor U16463 (N_16463,N_12575,N_11663);
nor U16464 (N_16464,N_12626,N_14417);
nand U16465 (N_16465,N_10057,N_11335);
nor U16466 (N_16466,N_11745,N_12736);
nand U16467 (N_16467,N_10353,N_13232);
and U16468 (N_16468,N_11410,N_13857);
nor U16469 (N_16469,N_13939,N_11987);
nand U16470 (N_16470,N_12714,N_12853);
and U16471 (N_16471,N_10616,N_11276);
nor U16472 (N_16472,N_11535,N_14267);
and U16473 (N_16473,N_12451,N_12488);
and U16474 (N_16474,N_10919,N_11065);
or U16475 (N_16475,N_10572,N_13180);
xor U16476 (N_16476,N_10564,N_14432);
nand U16477 (N_16477,N_13030,N_14063);
or U16478 (N_16478,N_14188,N_13460);
and U16479 (N_16479,N_10351,N_13762);
nor U16480 (N_16480,N_10152,N_13074);
nor U16481 (N_16481,N_12388,N_14749);
and U16482 (N_16482,N_13933,N_13638);
and U16483 (N_16483,N_13846,N_11735);
nor U16484 (N_16484,N_14199,N_14811);
nor U16485 (N_16485,N_12932,N_12748);
nor U16486 (N_16486,N_12839,N_10424);
nand U16487 (N_16487,N_12912,N_14450);
nand U16488 (N_16488,N_14279,N_12120);
xnor U16489 (N_16489,N_12128,N_11262);
and U16490 (N_16490,N_14307,N_12756);
nand U16491 (N_16491,N_11971,N_12079);
or U16492 (N_16492,N_12361,N_14335);
or U16493 (N_16493,N_13763,N_14571);
and U16494 (N_16494,N_10177,N_12251);
and U16495 (N_16495,N_13420,N_12046);
nor U16496 (N_16496,N_11763,N_11883);
or U16497 (N_16497,N_10173,N_10358);
nand U16498 (N_16498,N_10457,N_14182);
or U16499 (N_16499,N_13860,N_12224);
and U16500 (N_16500,N_12071,N_12468);
xor U16501 (N_16501,N_11847,N_14997);
xnor U16502 (N_16502,N_13556,N_13714);
and U16503 (N_16503,N_11831,N_10647);
nand U16504 (N_16504,N_14147,N_13224);
nand U16505 (N_16505,N_14510,N_13354);
nand U16506 (N_16506,N_10398,N_11764);
and U16507 (N_16507,N_12021,N_10769);
and U16508 (N_16508,N_12478,N_14483);
and U16509 (N_16509,N_12850,N_14286);
nand U16510 (N_16510,N_14880,N_10127);
nand U16511 (N_16511,N_13825,N_14934);
nand U16512 (N_16512,N_10532,N_11061);
or U16513 (N_16513,N_11049,N_11602);
or U16514 (N_16514,N_14914,N_12025);
xnor U16515 (N_16515,N_12962,N_12087);
and U16516 (N_16516,N_11331,N_14683);
xnor U16517 (N_16517,N_14556,N_14029);
and U16518 (N_16518,N_11710,N_14739);
or U16519 (N_16519,N_10664,N_14696);
and U16520 (N_16520,N_12859,N_12909);
or U16521 (N_16521,N_10611,N_10878);
nand U16522 (N_16522,N_13494,N_11400);
or U16523 (N_16523,N_10739,N_10206);
nor U16524 (N_16524,N_14820,N_12086);
or U16525 (N_16525,N_10417,N_10784);
nor U16526 (N_16526,N_12654,N_10720);
nand U16527 (N_16527,N_14520,N_11294);
xnor U16528 (N_16528,N_14894,N_10005);
and U16529 (N_16529,N_13877,N_14005);
nand U16530 (N_16530,N_11479,N_10925);
nand U16531 (N_16531,N_14068,N_11203);
or U16532 (N_16532,N_14333,N_11643);
nand U16533 (N_16533,N_11251,N_14577);
and U16534 (N_16534,N_13506,N_11114);
or U16535 (N_16535,N_13895,N_10196);
nand U16536 (N_16536,N_12833,N_13624);
nand U16537 (N_16537,N_11614,N_13614);
nand U16538 (N_16538,N_14426,N_12895);
or U16539 (N_16539,N_13154,N_12644);
and U16540 (N_16540,N_11741,N_12112);
and U16541 (N_16541,N_14960,N_11938);
or U16542 (N_16542,N_14122,N_13269);
or U16543 (N_16543,N_12904,N_12936);
and U16544 (N_16544,N_11848,N_12317);
nor U16545 (N_16545,N_13500,N_10296);
and U16546 (N_16546,N_13953,N_11454);
xnor U16547 (N_16547,N_10449,N_10989);
nand U16548 (N_16548,N_13702,N_13767);
and U16549 (N_16549,N_11709,N_13698);
nand U16550 (N_16550,N_11431,N_12400);
nand U16551 (N_16551,N_13753,N_11187);
nor U16552 (N_16552,N_12107,N_11407);
or U16553 (N_16553,N_11796,N_10562);
or U16554 (N_16554,N_13426,N_12818);
and U16555 (N_16555,N_11678,N_14624);
nor U16556 (N_16556,N_11448,N_12333);
nor U16557 (N_16557,N_11753,N_10629);
nand U16558 (N_16558,N_12809,N_12660);
and U16559 (N_16559,N_13318,N_14630);
xor U16560 (N_16560,N_11397,N_14434);
nor U16561 (N_16561,N_13991,N_13017);
xnor U16562 (N_16562,N_14380,N_13026);
nor U16563 (N_16563,N_14026,N_10729);
and U16564 (N_16564,N_10818,N_10788);
and U16565 (N_16565,N_12241,N_12162);
xnor U16566 (N_16566,N_10330,N_13849);
or U16567 (N_16567,N_14689,N_11273);
nand U16568 (N_16568,N_14884,N_10676);
or U16569 (N_16569,N_13256,N_13637);
nand U16570 (N_16570,N_14486,N_13285);
and U16571 (N_16571,N_14574,N_11983);
or U16572 (N_16572,N_12177,N_13042);
xor U16573 (N_16573,N_14142,N_13808);
or U16574 (N_16574,N_11864,N_10230);
or U16575 (N_16575,N_14448,N_13022);
and U16576 (N_16576,N_11982,N_10052);
or U16577 (N_16577,N_11137,N_14232);
nand U16578 (N_16578,N_10218,N_12460);
and U16579 (N_16579,N_10523,N_14784);
and U16580 (N_16580,N_12424,N_12110);
xnor U16581 (N_16581,N_11098,N_12510);
and U16582 (N_16582,N_13976,N_13674);
and U16583 (N_16583,N_10831,N_12968);
or U16584 (N_16584,N_13713,N_14077);
and U16585 (N_16585,N_10210,N_11386);
nor U16586 (N_16586,N_10905,N_10969);
nand U16587 (N_16587,N_10040,N_13507);
or U16588 (N_16588,N_14751,N_12035);
and U16589 (N_16589,N_11557,N_11647);
nor U16590 (N_16590,N_14447,N_11047);
xnor U16591 (N_16591,N_11849,N_12707);
nand U16592 (N_16592,N_12938,N_10963);
nand U16593 (N_16593,N_13968,N_12731);
or U16594 (N_16594,N_12417,N_12324);
nand U16595 (N_16595,N_14964,N_11690);
and U16596 (N_16596,N_10967,N_13189);
nand U16597 (N_16597,N_13781,N_10507);
or U16598 (N_16598,N_10109,N_10411);
nand U16599 (N_16599,N_13661,N_10921);
and U16600 (N_16600,N_14045,N_11253);
nand U16601 (N_16601,N_14241,N_14323);
nor U16602 (N_16602,N_11075,N_11377);
nand U16603 (N_16603,N_14893,N_10841);
or U16604 (N_16604,N_13484,N_10387);
xnor U16605 (N_16605,N_12801,N_11344);
or U16606 (N_16606,N_12091,N_11673);
nand U16607 (N_16607,N_14260,N_10245);
or U16608 (N_16608,N_11585,N_13509);
xor U16609 (N_16609,N_11655,N_12724);
nor U16610 (N_16610,N_13701,N_12496);
nor U16611 (N_16611,N_11264,N_12399);
or U16612 (N_16612,N_14933,N_12348);
nor U16613 (N_16613,N_13027,N_12742);
and U16614 (N_16614,N_13979,N_10088);
or U16615 (N_16615,N_10100,N_11818);
nor U16616 (N_16616,N_10583,N_13938);
and U16617 (N_16617,N_10048,N_11046);
nor U16618 (N_16618,N_11968,N_10587);
xnor U16619 (N_16619,N_11353,N_14341);
or U16620 (N_16620,N_10776,N_11435);
or U16621 (N_16621,N_12534,N_14161);
nor U16622 (N_16622,N_11355,N_10990);
or U16623 (N_16623,N_14206,N_13612);
nor U16624 (N_16624,N_11929,N_13926);
and U16625 (N_16625,N_14288,N_13532);
xnor U16626 (N_16626,N_11984,N_13751);
or U16627 (N_16627,N_13553,N_13032);
or U16628 (N_16628,N_10178,N_12518);
or U16629 (N_16629,N_11923,N_12411);
and U16630 (N_16630,N_13948,N_14502);
nor U16631 (N_16631,N_10909,N_10145);
nor U16632 (N_16632,N_14643,N_14449);
nand U16633 (N_16633,N_13481,N_11532);
and U16634 (N_16634,N_13585,N_10542);
nor U16635 (N_16635,N_13919,N_12447);
xnor U16636 (N_16636,N_12700,N_13410);
nor U16637 (N_16637,N_13000,N_12597);
or U16638 (N_16638,N_12560,N_13107);
nand U16639 (N_16639,N_12203,N_11613);
or U16640 (N_16640,N_12260,N_12814);
nand U16641 (N_16641,N_14433,N_13581);
nor U16642 (N_16642,N_12745,N_13663);
and U16643 (N_16643,N_12374,N_12964);
xor U16644 (N_16644,N_13712,N_11649);
and U16645 (N_16645,N_13517,N_14522);
nor U16646 (N_16646,N_11804,N_14154);
nor U16647 (N_16647,N_10694,N_14878);
nor U16648 (N_16648,N_14487,N_10322);
nand U16649 (N_16649,N_13130,N_14048);
nor U16650 (N_16650,N_13330,N_10143);
xnor U16651 (N_16651,N_13036,N_13633);
nor U16652 (N_16652,N_12562,N_11015);
xor U16653 (N_16653,N_10438,N_12083);
and U16654 (N_16654,N_11610,N_12689);
nor U16655 (N_16655,N_14639,N_12883);
or U16656 (N_16656,N_12207,N_14150);
nor U16657 (N_16657,N_13704,N_14280);
nand U16658 (N_16658,N_13264,N_13920);
nor U16659 (N_16659,N_12752,N_12275);
or U16660 (N_16660,N_10836,N_11867);
and U16661 (N_16661,N_11810,N_10975);
or U16662 (N_16662,N_11974,N_10205);
nand U16663 (N_16663,N_11067,N_12854);
nand U16664 (N_16664,N_11325,N_10368);
and U16665 (N_16665,N_11105,N_13832);
or U16666 (N_16666,N_11871,N_13603);
nor U16667 (N_16667,N_10018,N_10937);
and U16668 (N_16668,N_14040,N_11623);
or U16669 (N_16669,N_14539,N_13925);
and U16670 (N_16670,N_14792,N_13002);
nand U16671 (N_16671,N_14131,N_11300);
and U16672 (N_16672,N_13287,N_10274);
xor U16673 (N_16673,N_10828,N_10747);
and U16674 (N_16674,N_11330,N_13797);
or U16675 (N_16675,N_12286,N_13073);
and U16676 (N_16676,N_11076,N_12880);
or U16677 (N_16677,N_10718,N_13156);
nor U16678 (N_16678,N_12263,N_13408);
or U16679 (N_16679,N_11179,N_11708);
nand U16680 (N_16680,N_14047,N_12293);
and U16681 (N_16681,N_13831,N_14073);
and U16682 (N_16682,N_14250,N_10603);
or U16683 (N_16683,N_10381,N_12420);
nand U16684 (N_16684,N_10728,N_14948);
nand U16685 (N_16685,N_13873,N_10510);
and U16686 (N_16686,N_13466,N_13959);
nor U16687 (N_16687,N_13513,N_11260);
nor U16688 (N_16688,N_12802,N_10167);
or U16689 (N_16689,N_10832,N_12992);
nand U16690 (N_16690,N_11492,N_14127);
and U16691 (N_16691,N_10202,N_12381);
and U16692 (N_16692,N_14351,N_12944);
and U16693 (N_16693,N_12991,N_13007);
or U16694 (N_16694,N_12493,N_11128);
nand U16695 (N_16695,N_11202,N_12240);
and U16696 (N_16696,N_12430,N_13840);
nand U16697 (N_16697,N_12609,N_14638);
xor U16698 (N_16698,N_11879,N_12682);
nor U16699 (N_16699,N_14327,N_10405);
nor U16700 (N_16700,N_14770,N_11801);
nand U16701 (N_16701,N_12661,N_12732);
or U16702 (N_16702,N_11423,N_10010);
or U16703 (N_16703,N_14013,N_13518);
nand U16704 (N_16704,N_10441,N_12013);
or U16705 (N_16705,N_12198,N_10188);
and U16706 (N_16706,N_12618,N_10898);
nand U16707 (N_16707,N_13106,N_13957);
and U16708 (N_16708,N_10033,N_14915);
nor U16709 (N_16709,N_13893,N_13557);
or U16710 (N_16710,N_14192,N_13170);
nand U16711 (N_16711,N_12066,N_14310);
and U16712 (N_16712,N_10848,N_11130);
nor U16713 (N_16713,N_12294,N_10575);
nand U16714 (N_16714,N_14021,N_12595);
nor U16715 (N_16715,N_10500,N_13277);
or U16716 (N_16716,N_11962,N_12494);
and U16717 (N_16717,N_14647,N_11096);
nand U16718 (N_16718,N_14595,N_12924);
nor U16719 (N_16719,N_11605,N_13644);
or U16720 (N_16720,N_11990,N_11153);
or U16721 (N_16721,N_14748,N_10187);
nand U16722 (N_16722,N_12098,N_11676);
nand U16723 (N_16723,N_11773,N_14164);
or U16724 (N_16724,N_13343,N_10362);
nor U16725 (N_16725,N_14056,N_14504);
or U16726 (N_16726,N_14353,N_13307);
nand U16727 (N_16727,N_12095,N_10994);
nor U16728 (N_16728,N_11986,N_10809);
or U16729 (N_16729,N_14098,N_12031);
nand U16730 (N_16730,N_12089,N_10686);
xnor U16731 (N_16731,N_11016,N_10039);
and U16732 (N_16732,N_12258,N_11750);
and U16733 (N_16733,N_12516,N_13566);
nor U16734 (N_16734,N_14734,N_14758);
or U16735 (N_16735,N_14603,N_12816);
xnor U16736 (N_16736,N_10216,N_13041);
nor U16737 (N_16737,N_10884,N_14840);
and U16738 (N_16738,N_11517,N_14010);
or U16739 (N_16739,N_11907,N_14867);
and U16740 (N_16740,N_10997,N_10407);
and U16741 (N_16741,N_11174,N_14168);
nand U16742 (N_16742,N_10062,N_12744);
and U16743 (N_16743,N_12159,N_14089);
nor U16744 (N_16744,N_12879,N_12514);
and U16745 (N_16745,N_11028,N_12903);
nor U16746 (N_16746,N_13524,N_11761);
nor U16747 (N_16747,N_11970,N_14513);
nor U16748 (N_16748,N_13479,N_13978);
nand U16749 (N_16749,N_11976,N_11717);
xor U16750 (N_16750,N_10534,N_14269);
and U16751 (N_16751,N_11792,N_14395);
nand U16752 (N_16752,N_11943,N_13117);
xnor U16753 (N_16753,N_13718,N_11797);
nand U16754 (N_16754,N_14711,N_11126);
nor U16755 (N_16755,N_14763,N_14070);
nand U16756 (N_16756,N_12977,N_11050);
nor U16757 (N_16757,N_10174,N_14390);
and U16758 (N_16758,N_13076,N_13943);
and U16759 (N_16759,N_13439,N_13690);
or U16760 (N_16760,N_14242,N_10334);
or U16761 (N_16761,N_14354,N_13646);
xnor U16762 (N_16762,N_13982,N_14579);
nand U16763 (N_16763,N_11841,N_11149);
and U16764 (N_16764,N_12373,N_11606);
nand U16765 (N_16765,N_13749,N_12353);
and U16766 (N_16766,N_12629,N_11430);
or U16767 (N_16767,N_11346,N_13366);
nand U16768 (N_16768,N_14973,N_11498);
nand U16769 (N_16769,N_13934,N_10172);
nor U16770 (N_16770,N_11131,N_14587);
or U16771 (N_16771,N_10820,N_10867);
and U16772 (N_16772,N_14721,N_10688);
nand U16773 (N_16773,N_10265,N_10793);
or U16774 (N_16774,N_10336,N_13138);
xor U16775 (N_16775,N_11805,N_13552);
and U16776 (N_16776,N_10782,N_13201);
xnor U16777 (N_16777,N_12958,N_12130);
nand U16778 (N_16778,N_13582,N_14321);
nor U16779 (N_16779,N_12148,N_10980);
or U16780 (N_16780,N_11951,N_10992);
or U16781 (N_16781,N_10738,N_13110);
and U16782 (N_16782,N_10448,N_11490);
and U16783 (N_16783,N_10903,N_10141);
and U16784 (N_16784,N_12490,N_10800);
or U16785 (N_16785,N_14255,N_10333);
and U16786 (N_16786,N_13142,N_14980);
and U16787 (N_16787,N_14526,N_11712);
and U16788 (N_16788,N_13788,N_10907);
nor U16789 (N_16789,N_11833,N_11024);
or U16790 (N_16790,N_14001,N_10021);
nor U16791 (N_16791,N_14812,N_14616);
xor U16792 (N_16792,N_12508,N_14892);
and U16793 (N_16793,N_13070,N_14946);
nand U16794 (N_16794,N_12734,N_12779);
and U16795 (N_16795,N_13746,N_10176);
or U16796 (N_16796,N_10082,N_10226);
nand U16797 (N_16797,N_14645,N_10256);
nand U16798 (N_16798,N_12378,N_12976);
nand U16799 (N_16799,N_11638,N_13913);
or U16800 (N_16800,N_10529,N_11469);
nand U16801 (N_16801,N_10479,N_11491);
and U16802 (N_16802,N_14943,N_11256);
nand U16803 (N_16803,N_14922,N_10221);
nand U16804 (N_16804,N_13686,N_10155);
xnor U16805 (N_16805,N_14140,N_11094);
nand U16806 (N_16806,N_10602,N_12935);
nand U16807 (N_16807,N_11658,N_10267);
or U16808 (N_16808,N_10993,N_13590);
nor U16809 (N_16809,N_13445,N_12580);
nand U16810 (N_16810,N_14309,N_11121);
xnor U16811 (N_16811,N_13546,N_11932);
and U16812 (N_16812,N_10355,N_10816);
or U16813 (N_16813,N_12837,N_12149);
and U16814 (N_16814,N_13216,N_14018);
and U16815 (N_16815,N_13087,N_12160);
or U16816 (N_16816,N_14599,N_11520);
nor U16817 (N_16817,N_13748,N_11780);
nand U16818 (N_16818,N_12344,N_14412);
xor U16819 (N_16819,N_10124,N_10879);
nor U16820 (N_16820,N_10112,N_14169);
nor U16821 (N_16821,N_10049,N_13868);
nor U16822 (N_16822,N_10157,N_10985);
nand U16823 (N_16823,N_11455,N_10973);
xnor U16824 (N_16824,N_11083,N_10797);
or U16825 (N_16825,N_14166,N_10375);
nor U16826 (N_16826,N_12894,N_10250);
nand U16827 (N_16827,N_11705,N_12412);
xnor U16828 (N_16828,N_14263,N_12259);
xor U16829 (N_16829,N_14495,N_11026);
nand U16830 (N_16830,N_12988,N_12869);
and U16831 (N_16831,N_12078,N_13044);
nor U16832 (N_16832,N_13680,N_11292);
nor U16833 (N_16833,N_13406,N_12044);
nand U16834 (N_16834,N_10466,N_13793);
and U16835 (N_16835,N_11959,N_12994);
or U16836 (N_16836,N_12155,N_14788);
nor U16837 (N_16837,N_10955,N_11101);
nand U16838 (N_16838,N_10244,N_14590);
xnor U16839 (N_16839,N_12844,N_13433);
nand U16840 (N_16840,N_10916,N_14752);
and U16841 (N_16841,N_14824,N_12401);
nor U16842 (N_16842,N_11439,N_11392);
and U16843 (N_16843,N_12614,N_12300);
nand U16844 (N_16844,N_10426,N_13473);
and U16845 (N_16845,N_10865,N_10539);
or U16846 (N_16846,N_11426,N_14020);
and U16847 (N_16847,N_10227,N_14921);
or U16848 (N_16848,N_12668,N_14007);
and U16849 (N_16849,N_10504,N_14592);
nand U16850 (N_16850,N_14926,N_13205);
and U16851 (N_16851,N_14876,N_11139);
nand U16852 (N_16852,N_13194,N_10158);
and U16853 (N_16853,N_10116,N_14261);
nand U16854 (N_16854,N_10851,N_10933);
and U16855 (N_16855,N_10236,N_11758);
and U16856 (N_16856,N_10302,N_14272);
nor U16857 (N_16857,N_14299,N_12705);
and U16858 (N_16858,N_14249,N_10595);
nand U16859 (N_16859,N_12172,N_12102);
xnor U16860 (N_16860,N_13304,N_14439);
or U16861 (N_16861,N_14032,N_10257);
xor U16862 (N_16862,N_11496,N_10576);
and U16863 (N_16863,N_10168,N_10774);
nand U16864 (N_16864,N_10016,N_13583);
nand U16865 (N_16865,N_10763,N_13009);
and U16866 (N_16866,N_10350,N_12080);
and U16867 (N_16867,N_12672,N_14148);
nor U16868 (N_16868,N_12893,N_13628);
nand U16869 (N_16869,N_14043,N_14291);
or U16870 (N_16870,N_10656,N_11116);
nor U16871 (N_16871,N_10139,N_10833);
nor U16872 (N_16872,N_12221,N_13132);
or U16873 (N_16873,N_13179,N_10312);
or U16874 (N_16874,N_11494,N_12113);
nand U16875 (N_16875,N_10097,N_14213);
or U16876 (N_16876,N_14030,N_10183);
or U16877 (N_16877,N_10754,N_12590);
and U16878 (N_16878,N_12482,N_11657);
xor U16879 (N_16879,N_13392,N_10347);
or U16880 (N_16880,N_13488,N_10612);
and U16881 (N_16881,N_13791,N_11438);
and U16882 (N_16882,N_11980,N_11228);
nor U16883 (N_16883,N_14181,N_13776);
xnor U16884 (N_16884,N_12698,N_11425);
and U16885 (N_16885,N_13015,N_10003);
or U16886 (N_16886,N_11412,N_13312);
and U16887 (N_16887,N_12847,N_10846);
or U16888 (N_16888,N_13063,N_14276);
nand U16889 (N_16889,N_11333,N_10402);
nor U16890 (N_16890,N_12563,N_13125);
and U16891 (N_16891,N_13598,N_14358);
and U16892 (N_16892,N_12578,N_11326);
or U16893 (N_16893,N_10806,N_10986);
or U16894 (N_16894,N_13246,N_12729);
nand U16895 (N_16895,N_11912,N_10239);
nor U16896 (N_16896,N_13778,N_11596);
nor U16897 (N_16897,N_11172,N_10190);
nor U16898 (N_16898,N_14085,N_10184);
nor U16899 (N_16899,N_10282,N_12281);
xor U16900 (N_16900,N_12210,N_10366);
nand U16901 (N_16901,N_12407,N_13262);
nor U16902 (N_16902,N_10913,N_10968);
nor U16903 (N_16903,N_10485,N_10875);
or U16904 (N_16904,N_12305,N_10344);
or U16905 (N_16905,N_11003,N_10427);
nand U16906 (N_16906,N_12456,N_14538);
and U16907 (N_16907,N_14872,N_13184);
nor U16908 (N_16908,N_11777,N_13418);
and U16909 (N_16909,N_14220,N_12639);
xnor U16910 (N_16910,N_10775,N_14266);
and U16911 (N_16911,N_14745,N_13907);
nand U16912 (N_16912,N_11480,N_10715);
and U16913 (N_16913,N_12647,N_11246);
or U16914 (N_16914,N_12615,N_10129);
xnor U16915 (N_16915,N_10026,N_10404);
or U16916 (N_16916,N_14471,N_10495);
nand U16917 (N_16917,N_13588,N_11799);
nor U16918 (N_16918,N_11266,N_10904);
and U16919 (N_16919,N_14072,N_14362);
xnor U16920 (N_16920,N_11468,N_10706);
nand U16921 (N_16921,N_14158,N_10627);
nand U16922 (N_16922,N_12986,N_12775);
and U16923 (N_16923,N_14807,N_12817);
or U16924 (N_16924,N_12769,N_12178);
and U16925 (N_16925,N_13268,N_10243);
or U16926 (N_16926,N_10549,N_10450);
or U16927 (N_16927,N_13830,N_14828);
and U16928 (N_16928,N_14938,N_13901);
nand U16929 (N_16929,N_11583,N_11734);
or U16930 (N_16930,N_12222,N_12772);
nor U16931 (N_16931,N_14613,N_14529);
xor U16932 (N_16932,N_11873,N_13851);
and U16933 (N_16933,N_12741,N_10123);
nand U16934 (N_16934,N_11895,N_10293);
nor U16935 (N_16935,N_10480,N_14265);
nand U16936 (N_16936,N_12825,N_13660);
or U16937 (N_16937,N_11573,N_12390);
nor U16938 (N_16938,N_12794,N_10924);
nand U16939 (N_16939,N_11271,N_10271);
or U16940 (N_16940,N_10753,N_11723);
or U16941 (N_16941,N_12093,N_10804);
or U16942 (N_16942,N_12486,N_12685);
or U16943 (N_16943,N_13072,N_11926);
nor U16944 (N_16944,N_11886,N_10974);
and U16945 (N_16945,N_12692,N_12252);
or U16946 (N_16946,N_10538,N_12579);
nor U16947 (N_16947,N_11650,N_10455);
nand U16948 (N_16948,N_13848,N_10912);
nand U16949 (N_16949,N_13381,N_12987);
xor U16950 (N_16950,N_14978,N_11320);
nor U16951 (N_16951,N_11224,N_10815);
and U16952 (N_16952,N_13816,N_10144);
nor U16953 (N_16953,N_14268,N_11642);
nor U16954 (N_16954,N_13334,N_12898);
and U16955 (N_16955,N_11461,N_10247);
nor U16956 (N_16956,N_13429,N_12896);
nand U16957 (N_16957,N_12598,N_14610);
nand U16958 (N_16958,N_14074,N_14233);
nand U16959 (N_16959,N_12337,N_11129);
nand U16960 (N_16960,N_11633,N_14544);
or U16961 (N_16961,N_13328,N_12135);
nor U16962 (N_16962,N_11237,N_13640);
nor U16963 (N_16963,N_10670,N_11136);
or U16964 (N_16964,N_12688,N_14988);
xor U16965 (N_16965,N_13008,N_13222);
nand U16966 (N_16966,N_12739,N_10357);
and U16967 (N_16967,N_14027,N_11973);
nor U16968 (N_16968,N_12961,N_14011);
and U16969 (N_16969,N_14805,N_11063);
xnor U16970 (N_16970,N_14224,N_11770);
nand U16971 (N_16971,N_11625,N_13885);
nor U16972 (N_16972,N_11510,N_10893);
nand U16973 (N_16973,N_12308,N_12627);
and U16974 (N_16974,N_10897,N_11700);
nor U16975 (N_16975,N_13188,N_11459);
and U16976 (N_16976,N_13377,N_13955);
nor U16977 (N_16977,N_12843,N_12790);
or U16978 (N_16978,N_14132,N_11186);
nand U16979 (N_16979,N_14124,N_13528);
xnor U16980 (N_16980,N_10662,N_11389);
or U16981 (N_16981,N_10634,N_14623);
and U16982 (N_16982,N_10988,N_11062);
nand U16983 (N_16983,N_10582,N_13802);
nor U16984 (N_16984,N_11243,N_12675);
and U16985 (N_16985,N_13368,N_11860);
xor U16986 (N_16986,N_10453,N_14540);
xnor U16987 (N_16987,N_12480,N_10661);
nand U16988 (N_16988,N_12441,N_10131);
or U16989 (N_16989,N_12193,N_11304);
or U16990 (N_16990,N_12506,N_14109);
nand U16991 (N_16991,N_14084,N_13104);
and U16992 (N_16992,N_13782,N_13208);
and U16993 (N_16993,N_13563,N_13376);
or U16994 (N_16994,N_12544,N_12616);
and U16995 (N_16995,N_10827,N_12812);
and U16996 (N_16996,N_13611,N_13734);
or U16997 (N_16997,N_11897,N_10584);
or U16998 (N_16998,N_13050,N_11572);
and U16999 (N_16999,N_12036,N_14402);
or U17000 (N_17000,N_12683,N_10126);
xnor U17001 (N_17001,N_13144,N_14497);
nand U17002 (N_17002,N_10895,N_14772);
or U17003 (N_17003,N_10306,N_14500);
or U17004 (N_17004,N_10798,N_12498);
nor U17005 (N_17005,N_12452,N_11560);
nor U17006 (N_17006,N_13587,N_12501);
and U17007 (N_17007,N_11541,N_13944);
xor U17008 (N_17008,N_12929,N_13100);
nand U17009 (N_17009,N_12798,N_14986);
xnor U17010 (N_17010,N_12778,N_13503);
and U17011 (N_17011,N_13689,N_13051);
nand U17012 (N_17012,N_11229,N_14081);
and U17013 (N_17013,N_13992,N_14422);
and U17014 (N_17014,N_10386,N_14400);
nor U17015 (N_17015,N_13415,N_11194);
nor U17016 (N_17016,N_13937,N_11165);
and U17017 (N_17017,N_14794,N_14014);
nor U17018 (N_17018,N_12715,N_11108);
nor U17019 (N_17019,N_10456,N_13192);
nor U17020 (N_17020,N_12520,N_10198);
nand U17021 (N_17021,N_13525,N_13990);
xor U17022 (N_17022,N_13622,N_14787);
nor U17023 (N_17023,N_13705,N_11380);
and U17024 (N_17024,N_14730,N_14290);
nand U17025 (N_17025,N_11148,N_11211);
nand U17026 (N_17026,N_11941,N_14548);
or U17027 (N_17027,N_11928,N_11586);
or U17028 (N_17028,N_13202,N_13319);
and U17029 (N_17029,N_10668,N_13758);
or U17030 (N_17030,N_12047,N_12601);
or U17031 (N_17031,N_14670,N_12952);
nand U17032 (N_17032,N_14332,N_11558);
or U17033 (N_17033,N_13511,N_13512);
and U17034 (N_17034,N_13731,N_10433);
and U17035 (N_17035,N_12695,N_14702);
nand U17036 (N_17036,N_12283,N_13477);
nor U17037 (N_17037,N_12764,N_13052);
nand U17038 (N_17038,N_13421,N_13465);
or U17039 (N_17039,N_10801,N_10029);
nor U17040 (N_17040,N_10961,N_12747);
nand U17041 (N_17041,N_13482,N_14444);
nor U17042 (N_17042,N_11470,N_11135);
or U17043 (N_17043,N_13964,N_14532);
or U17044 (N_17044,N_11546,N_11689);
xnor U17045 (N_17045,N_12900,N_13523);
and U17046 (N_17046,N_10012,N_12576);
xnor U17047 (N_17047,N_13678,N_14427);
and U17048 (N_17048,N_14559,N_10101);
and U17049 (N_17049,N_13755,N_10528);
nand U17050 (N_17050,N_12326,N_14415);
or U17051 (N_17051,N_14041,N_11619);
nor U17052 (N_17052,N_11830,N_11369);
or U17053 (N_17053,N_10364,N_12733);
and U17054 (N_17054,N_13541,N_13294);
xnor U17055 (N_17055,N_10948,N_13916);
and U17056 (N_17056,N_10195,N_11564);
nor U17057 (N_17057,N_14873,N_14356);
xnor U17058 (N_17058,N_14889,N_14845);
and U17059 (N_17059,N_11169,N_13615);
nor U17060 (N_17060,N_14703,N_14435);
xor U17061 (N_17061,N_13703,N_12022);
nor U17062 (N_17062,N_10232,N_14407);
nor U17063 (N_17063,N_13462,N_10869);
or U17064 (N_17064,N_10228,N_13679);
or U17065 (N_17065,N_12332,N_10192);
nand U17066 (N_17066,N_11534,N_14765);
or U17067 (N_17067,N_13416,N_12723);
nand U17068 (N_17068,N_12918,N_14360);
or U17069 (N_17069,N_10745,N_12161);
or U17070 (N_17070,N_11343,N_10481);
and U17071 (N_17071,N_10971,N_12076);
nand U17072 (N_17072,N_12819,N_11073);
or U17073 (N_17073,N_11390,N_10494);
or U17074 (N_17074,N_12550,N_14733);
nand U17075 (N_17075,N_10290,N_14163);
nand U17076 (N_17076,N_10692,N_12184);
or U17077 (N_17077,N_11550,N_10319);
nor U17078 (N_17078,N_10936,N_13054);
nand U17079 (N_17079,N_11378,N_13759);
or U17080 (N_17080,N_11030,N_14629);
xor U17081 (N_17081,N_13855,N_13575);
xor U17082 (N_17082,N_12271,N_14780);
xnor U17083 (N_17083,N_12423,N_13807);
nand U17084 (N_17084,N_11181,N_11861);
or U17085 (N_17085,N_10389,N_11878);
xnor U17086 (N_17086,N_11577,N_10470);
nor U17087 (N_17087,N_11641,N_12697);
and U17088 (N_17088,N_12208,N_11533);
nand U17089 (N_17089,N_13950,N_14953);
or U17090 (N_17090,N_12219,N_14778);
or U17091 (N_17091,N_14138,N_10622);
or U17092 (N_17092,N_12069,N_11301);
and U17093 (N_17093,N_14012,N_12350);
or U17094 (N_17094,N_11854,N_13602);
nand U17095 (N_17095,N_10301,N_10970);
and U17096 (N_17096,N_11885,N_12217);
and U17097 (N_17097,N_10032,N_14790);
or U17098 (N_17098,N_12492,N_12974);
or U17099 (N_17099,N_10506,N_13316);
and U17100 (N_17100,N_12310,N_12119);
and U17101 (N_17101,N_12462,N_13550);
nor U17102 (N_17102,N_11693,N_12297);
nand U17103 (N_17103,N_12643,N_10182);
nor U17104 (N_17104,N_12558,N_14698);
nand U17105 (N_17105,N_12513,N_10308);
or U17106 (N_17106,N_14492,N_14558);
nor U17107 (N_17107,N_11589,N_13325);
xor U17108 (N_17108,N_11308,N_12040);
and U17109 (N_17109,N_10654,N_13190);
nor U17110 (N_17110,N_11903,N_10598);
nand U17111 (N_17111,N_11699,N_14429);
and U17112 (N_17112,N_14552,N_10266);
nor U17113 (N_17113,N_13315,N_14753);
and U17114 (N_17114,N_14454,N_11428);
and U17115 (N_17115,N_12568,N_10204);
and U17116 (N_17116,N_10711,N_12244);
nand U17117 (N_17117,N_14967,N_10901);
and U17118 (N_17118,N_14167,N_13137);
and U17119 (N_17119,N_11782,N_11217);
xor U17120 (N_17120,N_12780,N_14855);
nor U17121 (N_17121,N_12710,N_11230);
and U17122 (N_17122,N_10702,N_11670);
xor U17123 (N_17123,N_10153,N_14031);
nand U17124 (N_17124,N_14292,N_10175);
and U17125 (N_17125,N_14910,N_11665);
nand U17126 (N_17126,N_12367,N_14620);
nor U17127 (N_17127,N_10591,N_14671);
nand U17128 (N_17128,N_13977,N_12718);
xnor U17129 (N_17129,N_13981,N_10136);
nand U17130 (N_17130,N_12188,N_10792);
and U17131 (N_17131,N_10811,N_10508);
nor U17132 (N_17132,N_10624,N_11845);
or U17133 (N_17133,N_11762,N_12495);
nor U17134 (N_17134,N_12554,N_12292);
or U17135 (N_17135,N_10813,N_10475);
nand U17136 (N_17136,N_12338,N_10060);
nor U17137 (N_17137,N_12298,N_12466);
or U17138 (N_17138,N_12882,N_13383);
xor U17139 (N_17139,N_12574,N_14798);
nor U17140 (N_17140,N_11566,N_11297);
xor U17141 (N_17141,N_14511,N_12502);
or U17142 (N_17142,N_14340,N_11085);
or U17143 (N_17143,N_10394,N_12726);
and U17144 (N_17144,N_12799,N_10374);
xor U17145 (N_17145,N_14667,N_14065);
or U17146 (N_17146,N_14827,N_11620);
and U17147 (N_17147,N_13717,N_11703);
xnor U17148 (N_17148,N_13374,N_14779);
or U17149 (N_17149,N_10531,N_10340);
nor U17150 (N_17150,N_13077,N_14057);
nand U17151 (N_17151,N_11756,N_12959);
nor U17152 (N_17152,N_13657,N_11489);
nor U17153 (N_17153,N_14111,N_11768);
and U17154 (N_17154,N_10054,N_13430);
xor U17155 (N_17155,N_12948,N_14575);
xnor U17156 (N_17156,N_13545,N_11442);
and U17157 (N_17157,N_10085,N_11037);
nor U17158 (N_17158,N_10902,N_10764);
nor U17159 (N_17159,N_13472,N_10429);
xnor U17160 (N_17160,N_14682,N_14974);
or U17161 (N_17161,N_13930,N_12642);
xnor U17162 (N_17162,N_11554,N_14143);
nand U17163 (N_17163,N_12034,N_11562);
xor U17164 (N_17164,N_11815,N_10497);
nand U17165 (N_17165,N_10941,N_12396);
and U17166 (N_17166,N_12646,N_12074);
nand U17167 (N_17167,N_13033,N_12415);
or U17168 (N_17168,N_14662,N_13728);
xor U17169 (N_17169,N_10072,N_14600);
or U17170 (N_17170,N_12085,N_12237);
nor U17171 (N_17171,N_14916,N_13562);
or U17172 (N_17172,N_12823,N_11675);
xnor U17173 (N_17173,N_12103,N_10520);
nor U17174 (N_17174,N_14561,N_14411);
or U17175 (N_17175,N_10501,N_11681);
or U17176 (N_17176,N_13300,N_10104);
xnor U17177 (N_17177,N_12528,N_14838);
xnor U17178 (N_17178,N_13931,N_13723);
and U17179 (N_17179,N_10646,N_12052);
and U17180 (N_17180,N_14799,N_10446);
nor U17181 (N_17181,N_13103,N_14883);
nor U17182 (N_17182,N_13865,N_13220);
xor U17183 (N_17183,N_12039,N_13458);
nand U17184 (N_17184,N_11366,N_11384);
or U17185 (N_17185,N_12540,N_14762);
or U17186 (N_17186,N_11622,N_10563);
nand U17187 (N_17187,N_12852,N_13061);
and U17188 (N_17188,N_14764,N_12246);
nand U17189 (N_17189,N_14802,N_10051);
nand U17190 (N_17190,N_12527,N_10342);
nand U17191 (N_17191,N_13149,N_14254);
xnor U17192 (N_17192,N_11124,N_11328);
xor U17193 (N_17193,N_14165,N_13419);
nor U17194 (N_17194,N_14719,N_11561);
nor U17195 (N_17195,N_12213,N_11511);
nand U17196 (N_17196,N_14051,N_11214);
nand U17197 (N_17197,N_14355,N_13486);
nor U17198 (N_17198,N_12840,N_12624);
or U17199 (N_17199,N_12418,N_10477);
nor U17200 (N_17200,N_12795,N_13414);
nor U17201 (N_17201,N_12358,N_13757);
nand U17202 (N_17202,N_11949,N_10758);
and U17203 (N_17203,N_10976,N_14781);
nand U17204 (N_17204,N_12092,N_13639);
and U17205 (N_17205,N_13403,N_13101);
and U17206 (N_17206,N_13001,N_10091);
nand U17207 (N_17207,N_10796,N_12410);
and U17208 (N_17208,N_10637,N_11020);
nor U17209 (N_17209,N_14842,N_10081);
nor U17210 (N_17210,N_12587,N_14732);
nor U17211 (N_17211,N_10823,N_10765);
nand U17212 (N_17212,N_13675,N_10868);
and U17213 (N_17213,N_12972,N_13988);
nor U17214 (N_17214,N_13291,N_11960);
or U17215 (N_17215,N_13606,N_10275);
nand U17216 (N_17216,N_10570,N_13347);
nand U17217 (N_17217,N_10513,N_12256);
and U17218 (N_17218,N_13247,N_10900);
or U17219 (N_17219,N_11483,N_10940);
nand U17220 (N_17220,N_11667,N_12055);
nand U17221 (N_17221,N_14103,N_12316);
and U17222 (N_17222,N_12791,N_12911);
or U17223 (N_17223,N_10379,N_13984);
nor U17224 (N_17224,N_10111,N_11478);
xnor U17225 (N_17225,N_12448,N_12939);
nand U17226 (N_17226,N_10537,N_14034);
nand U17227 (N_17227,N_11278,N_11634);
xnor U17228 (N_17228,N_11862,N_14585);
xnor U17229 (N_17229,N_13337,N_14058);
or U17230 (N_17230,N_14663,N_14849);
or U17231 (N_17231,N_14022,N_11445);
or U17232 (N_17232,N_11263,N_10295);
nand U17233 (N_17233,N_14100,N_10063);
and U17234 (N_17234,N_10071,N_11238);
or U17235 (N_17235,N_12313,N_13761);
xnor U17236 (N_17236,N_10440,N_14741);
and U17237 (N_17237,N_11029,N_12758);
and U17238 (N_17238,N_13375,N_12342);
and U17239 (N_17239,N_13171,N_14367);
and U17240 (N_17240,N_14326,N_13480);
and U17241 (N_17241,N_10740,N_13636);
nand U17242 (N_17242,N_12890,N_12270);
nand U17243 (N_17243,N_11009,N_10954);
xnor U17244 (N_17244,N_12101,N_10493);
and U17245 (N_17245,N_14350,N_12730);
or U17246 (N_17246,N_14767,N_11296);
nand U17247 (N_17247,N_11034,N_10979);
and U17248 (N_17248,N_13338,N_14903);
and U17249 (N_17249,N_13437,N_11388);
or U17250 (N_17250,N_12070,N_13345);
nor U17251 (N_17251,N_11868,N_12489);
nor U17252 (N_17252,N_11495,N_14187);
and U17253 (N_17253,N_12461,N_14473);
or U17254 (N_17254,N_13243,N_14464);
nand U17255 (N_17255,N_11227,N_10095);
nand U17256 (N_17256,N_11996,N_14800);
and U17257 (N_17257,N_11493,N_10007);
xnor U17258 (N_17258,N_12946,N_13716);
xnor U17259 (N_17259,N_12916,N_10309);
nor U17260 (N_17260,N_13863,N_13836);
and U17261 (N_17261,N_10682,N_13013);
or U17262 (N_17262,N_12507,N_14095);
and U17263 (N_17263,N_12307,N_11731);
and U17264 (N_17264,N_11829,N_14485);
nand U17265 (N_17265,N_13340,N_11537);
nor U17266 (N_17266,N_10474,N_10681);
and U17267 (N_17267,N_14746,N_13217);
xnor U17268 (N_17268,N_12581,N_10829);
nor U17269 (N_17269,N_10601,N_10821);
xor U17270 (N_17270,N_11910,N_12603);
or U17271 (N_17271,N_11865,N_14120);
and U17272 (N_17272,N_10982,N_14221);
nand U17273 (N_17273,N_13271,N_10874);
and U17274 (N_17274,N_13152,N_11039);
and U17275 (N_17275,N_12443,N_13569);
and U17276 (N_17276,N_12421,N_14627);
and U17277 (N_17277,N_10934,N_13798);
and U17278 (N_17278,N_11485,N_12570);
xnor U17279 (N_17279,N_12663,N_13252);
xnor U17280 (N_17280,N_14785,N_13568);
nor U17281 (N_17281,N_13649,N_11338);
or U17282 (N_17282,N_10278,N_10749);
nor U17283 (N_17283,N_11551,N_12274);
nand U17284 (N_17284,N_13641,N_12463);
or U17285 (N_17285,N_10540,N_13613);
or U17286 (N_17286,N_12693,N_12000);
and U17287 (N_17287,N_13904,N_13292);
nor U17288 (N_17288,N_10592,N_11851);
and U17289 (N_17289,N_11418,N_12599);
and U17290 (N_17290,N_14176,N_13549);
nand U17291 (N_17291,N_11048,N_11059);
or U17292 (N_17292,N_13118,N_10802);
nor U17293 (N_17293,N_10596,N_11859);
and U17294 (N_17294,N_13852,N_14237);
nor U17295 (N_17295,N_13046,N_13963);
or U17296 (N_17296,N_11434,N_11852);
nand U17297 (N_17297,N_10840,N_12266);
and U17298 (N_17298,N_10766,N_10805);
nand U17299 (N_17299,N_11364,N_10287);
nor U17300 (N_17300,N_11324,N_12393);
nor U17301 (N_17301,N_13833,N_14071);
nor U17302 (N_17302,N_11306,N_11097);
and U17303 (N_17303,N_10171,N_12960);
nand U17304 (N_17304,N_12719,N_11086);
nand U17305 (N_17305,N_10346,N_12249);
or U17306 (N_17306,N_10201,N_11578);
or U17307 (N_17307,N_12325,N_14965);
nand U17308 (N_17308,N_11781,N_10700);
xnor U17309 (N_17309,N_14879,N_13965);
and U17310 (N_17310,N_10623,N_10556);
and U17311 (N_17311,N_13995,N_11866);
nand U17312 (N_17312,N_12846,N_10107);
or U17313 (N_17313,N_11078,N_10341);
nand U17314 (N_17314,N_11604,N_13601);
or U17315 (N_17315,N_10663,N_13652);
nor U17316 (N_17316,N_12247,N_11151);
nand U17317 (N_17317,N_10382,N_12923);
or U17318 (N_17318,N_10795,N_13629);
nand U17319 (N_17319,N_13346,N_10332);
and U17320 (N_17320,N_13872,N_14881);
nand U17321 (N_17321,N_12740,N_10297);
nand U17322 (N_17322,N_11323,N_13856);
or U17323 (N_17323,N_10316,N_12889);
nand U17324 (N_17324,N_13555,N_14619);
or U17325 (N_17325,N_10577,N_14716);
nor U17326 (N_17326,N_11254,N_13284);
and U17327 (N_17327,N_10061,N_13847);
nand U17328 (N_17328,N_13619,N_12282);
or U17329 (N_17329,N_12075,N_13253);
and U17330 (N_17330,N_14216,N_12116);
xnor U17331 (N_17331,N_10189,N_12464);
or U17332 (N_17332,N_14420,N_11529);
or U17333 (N_17333,N_13508,N_12993);
nand U17334 (N_17334,N_13108,N_12592);
and U17335 (N_17335,N_13161,N_10286);
and U17336 (N_17336,N_14701,N_13487);
xor U17337 (N_17337,N_10108,N_11935);
nor U17338 (N_17338,N_13671,N_11631);
nand U17339 (N_17339,N_13295,N_13754);
and U17340 (N_17340,N_10673,N_13120);
and U17341 (N_17341,N_12062,N_12003);
nor U17342 (N_17342,N_13898,N_10632);
nand U17343 (N_17343,N_13290,N_11754);
nor U17344 (N_17344,N_12757,N_14567);
or U17345 (N_17345,N_12702,N_11958);
and U17346 (N_17346,N_11544,N_11350);
or U17347 (N_17347,N_11652,N_13311);
nor U17348 (N_17348,N_12288,N_13668);
nand U17349 (N_17349,N_10853,N_12571);
nor U17350 (N_17350,N_10068,N_11118);
nor U17351 (N_17351,N_13593,N_14674);
or U17352 (N_17352,N_11180,N_13908);
nor U17353 (N_17353,N_14720,N_12206);
or U17354 (N_17354,N_13153,N_11348);
or U17355 (N_17355,N_12885,N_10280);
xor U17356 (N_17356,N_12586,N_10505);
and U17357 (N_17357,N_12043,N_12362);
nor U17358 (N_17358,N_12776,N_10621);
and U17359 (N_17359,N_11140,N_14555);
xor U17360 (N_17360,N_12181,N_14197);
nand U17361 (N_17361,N_12389,N_12867);
and U17362 (N_17362,N_11536,N_11696);
nand U17363 (N_17363,N_10409,N_10102);
and U17364 (N_17364,N_10658,N_12708);
xor U17365 (N_17365,N_14416,N_14940);
and U17366 (N_17366,N_12945,N_14055);
or U17367 (N_17367,N_13176,N_13141);
xnor U17368 (N_17368,N_13230,N_11803);
nor U17369 (N_17369,N_13162,N_12921);
and U17370 (N_17370,N_12226,N_11957);
or U17371 (N_17371,N_10756,N_11270);
and U17372 (N_17372,N_10891,N_14382);
or U17373 (N_17373,N_14470,N_10070);
nor U17374 (N_17374,N_12970,N_11268);
or U17375 (N_17375,N_12121,N_13720);
nand U17376 (N_17376,N_11707,N_11162);
nand U17377 (N_17377,N_12048,N_12998);
or U17378 (N_17378,N_11916,N_13589);
and U17379 (N_17379,N_14863,N_11417);
and U17380 (N_17380,N_14816,N_10044);
and U17381 (N_17381,N_14542,N_10578);
xor U17382 (N_17382,N_12538,N_13654);
nor U17383 (N_17383,N_11580,N_14706);
or U17384 (N_17384,N_14222,N_14215);
nor U17385 (N_17385,N_12999,N_13785);
nand U17386 (N_17386,N_14902,N_12638);
nand U17387 (N_17387,N_11821,N_12783);
nor U17388 (N_17388,N_11156,N_12385);
nand U17389 (N_17389,N_10995,N_13936);
or U17390 (N_17390,N_11574,N_13656);
xnor U17391 (N_17391,N_11615,N_11714);
nand U17392 (N_17392,N_10464,N_14637);
nand U17393 (N_17393,N_13388,N_12239);
xor U17394 (N_17394,N_14118,N_12171);
nor U17395 (N_17395,N_11281,N_13719);
xnor U17396 (N_17396,N_12068,N_14135);
or U17397 (N_17397,N_14498,N_12657);
and U17398 (N_17398,N_12053,N_14678);
nand U17399 (N_17399,N_12059,N_12202);
nand U17400 (N_17400,N_11093,N_14024);
and U17401 (N_17401,N_10083,N_12604);
and U17402 (N_17402,N_12474,N_11500);
nor U17403 (N_17403,N_14968,N_12917);
or U17404 (N_17404,N_14908,N_10215);
and U17405 (N_17405,N_11549,N_12212);
or U17406 (N_17406,N_12064,N_13940);
and U17407 (N_17407,N_13572,N_10922);
nand U17408 (N_17408,N_13206,N_11787);
nor U17409 (N_17409,N_14203,N_12190);
or U17410 (N_17410,N_12082,N_10412);
and U17411 (N_17411,N_13031,N_10020);
and U17412 (N_17412,N_13859,N_14523);
nor U17413 (N_17413,N_14660,N_14457);
nand U17414 (N_17414,N_12143,N_11616);
or U17415 (N_17415,N_13620,N_10445);
and U17416 (N_17416,N_13212,N_12475);
or U17417 (N_17417,N_14115,N_10580);
nor U17418 (N_17418,N_11607,N_11618);
nand U17419 (N_17419,N_12664,N_12197);
nand U17420 (N_17420,N_14972,N_11786);
or U17421 (N_17421,N_11526,N_10135);
or U17422 (N_17422,N_10073,N_14437);
and U17423 (N_17423,N_11081,N_10727);
and U17424 (N_17424,N_10304,N_13871);
nand U17425 (N_17425,N_13630,N_10502);
and U17426 (N_17426,N_10817,N_13867);
and U17427 (N_17427,N_13526,N_10079);
nand U17428 (N_17428,N_13148,N_13625);
nor U17429 (N_17429,N_10785,N_12552);
or U17430 (N_17430,N_10524,N_13332);
nand U17431 (N_17431,N_13228,N_10767);
nand U17432 (N_17432,N_10397,N_10437);
and U17433 (N_17433,N_11467,N_11295);
or U17434 (N_17434,N_13810,N_10543);
nor U17435 (N_17435,N_13353,N_11265);
nand U17436 (N_17436,N_14231,N_13263);
and U17437 (N_17437,N_11138,N_14791);
nand U17438 (N_17438,N_11396,N_11834);
nor U17439 (N_17439,N_13529,N_11206);
nand U17440 (N_17440,N_14859,N_12104);
xor U17441 (N_17441,N_14793,N_13739);
nand U17442 (N_17442,N_10015,N_14866);
xor U17443 (N_17443,N_12621,N_12370);
nor U17444 (N_17444,N_10371,N_12152);
nand U17445 (N_17445,N_14346,N_14364);
or U17446 (N_17446,N_10704,N_13098);
and U17447 (N_17447,N_10066,N_10288);
nand U17448 (N_17448,N_14134,N_10911);
and U17449 (N_17449,N_13404,N_14825);
or U17450 (N_17450,N_12877,N_10892);
xor U17451 (N_17451,N_14398,N_10463);
or U17452 (N_17452,N_12010,N_11145);
and U17453 (N_17453,N_13090,N_11894);
or U17454 (N_17454,N_13288,N_12111);
nand U17455 (N_17455,N_10451,N_14121);
nor U17456 (N_17456,N_13733,N_13453);
or U17457 (N_17457,N_10164,N_10599);
nand U17458 (N_17458,N_12284,N_12228);
and U17459 (N_17459,N_10518,N_14317);
or U17460 (N_17460,N_11784,N_11106);
xor U17461 (N_17461,N_12028,N_11749);
nand U17462 (N_17462,N_14984,N_11559);
nand U17463 (N_17463,N_14004,N_10120);
nor U17464 (N_17464,N_11711,N_14219);
xnor U17465 (N_17465,N_10235,N_13065);
and U17466 (N_17466,N_11220,N_10873);
nand U17467 (N_17467,N_13043,N_10413);
or U17468 (N_17468,N_12556,N_11576);
xnor U17469 (N_17469,N_13691,N_13888);
or U17470 (N_17470,N_10630,N_12306);
nand U17471 (N_17471,N_13864,N_10625);
nor U17472 (N_17472,N_10526,N_14604);
or U17473 (N_17473,N_12822,N_11440);
or U17474 (N_17474,N_14744,N_14553);
xor U17475 (N_17475,N_10631,N_13373);
and U17476 (N_17476,N_11807,N_11043);
nand U17477 (N_17477,N_12201,N_11653);
or U17478 (N_17478,N_13544,N_10376);
and U17479 (N_17479,N_14936,N_14534);
or U17480 (N_17480,N_13079,N_14819);
or U17481 (N_17481,N_14289,N_13203);
nand U17482 (N_17482,N_14598,N_13272);
and U17483 (N_17483,N_10017,N_10436);
nor U17484 (N_17484,N_12735,N_14079);
nand U17485 (N_17485,N_14615,N_11685);
nand U17486 (N_17486,N_10272,N_14430);
nor U17487 (N_17487,N_11790,N_12835);
xnor U17488 (N_17488,N_12223,N_10299);
and U17489 (N_17489,N_14632,N_10926);
or U17490 (N_17490,N_10999,N_11247);
and U17491 (N_17491,N_13540,N_11359);
and U17492 (N_17492,N_10643,N_13129);
nor U17493 (N_17493,N_13235,N_13367);
nand U17494 (N_17494,N_13233,N_10550);
nand U17495 (N_17495,N_12773,N_12655);
nor U17496 (N_17496,N_13358,N_12129);
nor U17497 (N_17497,N_11963,N_12176);
and U17498 (N_17498,N_14700,N_14562);
xor U17499 (N_17499,N_11347,N_13265);
nand U17500 (N_17500,N_11181,N_12846);
and U17501 (N_17501,N_10540,N_11276);
or U17502 (N_17502,N_14935,N_14286);
nor U17503 (N_17503,N_10246,N_10392);
nand U17504 (N_17504,N_11185,N_13682);
nor U17505 (N_17505,N_11948,N_13338);
nand U17506 (N_17506,N_13081,N_12612);
or U17507 (N_17507,N_10082,N_12389);
and U17508 (N_17508,N_13752,N_14811);
nand U17509 (N_17509,N_11903,N_12998);
and U17510 (N_17510,N_14979,N_14902);
and U17511 (N_17511,N_12869,N_10418);
nand U17512 (N_17512,N_14582,N_14395);
or U17513 (N_17513,N_13933,N_14010);
and U17514 (N_17514,N_10349,N_14596);
and U17515 (N_17515,N_10623,N_13939);
xor U17516 (N_17516,N_10842,N_11702);
or U17517 (N_17517,N_14062,N_13023);
nor U17518 (N_17518,N_13368,N_10080);
and U17519 (N_17519,N_11242,N_11810);
nor U17520 (N_17520,N_14773,N_12848);
or U17521 (N_17521,N_12630,N_14103);
or U17522 (N_17522,N_12900,N_13080);
nand U17523 (N_17523,N_10542,N_13970);
nand U17524 (N_17524,N_13644,N_11150);
and U17525 (N_17525,N_12371,N_10835);
or U17526 (N_17526,N_12939,N_12384);
or U17527 (N_17527,N_12872,N_13285);
or U17528 (N_17528,N_10750,N_14546);
nand U17529 (N_17529,N_13524,N_14035);
xor U17530 (N_17530,N_12393,N_14956);
nand U17531 (N_17531,N_11872,N_11324);
and U17532 (N_17532,N_11656,N_11304);
or U17533 (N_17533,N_13202,N_14478);
or U17534 (N_17534,N_11632,N_13931);
and U17535 (N_17535,N_10811,N_10513);
nor U17536 (N_17536,N_10494,N_14357);
nand U17537 (N_17537,N_13677,N_11461);
or U17538 (N_17538,N_10918,N_13906);
and U17539 (N_17539,N_13001,N_13185);
xor U17540 (N_17540,N_12016,N_13208);
nand U17541 (N_17541,N_13733,N_13634);
nand U17542 (N_17542,N_11429,N_11863);
and U17543 (N_17543,N_13247,N_11974);
nor U17544 (N_17544,N_12125,N_13154);
xnor U17545 (N_17545,N_10536,N_14525);
nor U17546 (N_17546,N_12313,N_10800);
or U17547 (N_17547,N_14273,N_13758);
or U17548 (N_17548,N_14456,N_10595);
nand U17549 (N_17549,N_14762,N_12869);
nand U17550 (N_17550,N_13247,N_10438);
nand U17551 (N_17551,N_13685,N_14749);
and U17552 (N_17552,N_10813,N_14941);
nand U17553 (N_17553,N_13789,N_14354);
nand U17554 (N_17554,N_12289,N_14093);
nor U17555 (N_17555,N_10884,N_10335);
xor U17556 (N_17556,N_13668,N_13718);
nor U17557 (N_17557,N_13690,N_11473);
nand U17558 (N_17558,N_13846,N_10481);
nor U17559 (N_17559,N_14807,N_13678);
xnor U17560 (N_17560,N_12702,N_11830);
xor U17561 (N_17561,N_10247,N_11591);
nand U17562 (N_17562,N_12887,N_13894);
nor U17563 (N_17563,N_12989,N_11617);
and U17564 (N_17564,N_11336,N_10940);
and U17565 (N_17565,N_11103,N_10800);
xor U17566 (N_17566,N_11214,N_14513);
nor U17567 (N_17567,N_12942,N_12936);
xor U17568 (N_17568,N_10698,N_11998);
nor U17569 (N_17569,N_10998,N_10644);
and U17570 (N_17570,N_14344,N_11786);
nor U17571 (N_17571,N_10415,N_11669);
nor U17572 (N_17572,N_13644,N_13097);
nor U17573 (N_17573,N_12936,N_10699);
xnor U17574 (N_17574,N_12286,N_12119);
or U17575 (N_17575,N_11181,N_14310);
and U17576 (N_17576,N_13568,N_12224);
nand U17577 (N_17577,N_11754,N_12814);
and U17578 (N_17578,N_10465,N_11284);
and U17579 (N_17579,N_11685,N_13070);
xor U17580 (N_17580,N_10823,N_12238);
or U17581 (N_17581,N_14509,N_11026);
or U17582 (N_17582,N_11251,N_13077);
nor U17583 (N_17583,N_12353,N_10222);
and U17584 (N_17584,N_13803,N_14436);
nor U17585 (N_17585,N_11589,N_12348);
and U17586 (N_17586,N_10133,N_12309);
nor U17587 (N_17587,N_10782,N_10770);
and U17588 (N_17588,N_13017,N_11038);
nand U17589 (N_17589,N_14545,N_12003);
or U17590 (N_17590,N_10845,N_13545);
and U17591 (N_17591,N_11316,N_11811);
nor U17592 (N_17592,N_11990,N_11524);
nor U17593 (N_17593,N_13078,N_12556);
nand U17594 (N_17594,N_14734,N_10790);
and U17595 (N_17595,N_10583,N_10792);
nor U17596 (N_17596,N_14536,N_13596);
or U17597 (N_17597,N_13141,N_13445);
and U17598 (N_17598,N_14235,N_13222);
and U17599 (N_17599,N_13407,N_12449);
nand U17600 (N_17600,N_12779,N_14355);
xor U17601 (N_17601,N_11189,N_10780);
nor U17602 (N_17602,N_14160,N_12668);
or U17603 (N_17603,N_12713,N_10947);
and U17604 (N_17604,N_12640,N_11570);
nor U17605 (N_17605,N_10631,N_11800);
nor U17606 (N_17606,N_11427,N_10539);
xnor U17607 (N_17607,N_12460,N_11019);
nor U17608 (N_17608,N_12159,N_13295);
xor U17609 (N_17609,N_10010,N_11703);
or U17610 (N_17610,N_10543,N_14859);
nand U17611 (N_17611,N_14262,N_14449);
nand U17612 (N_17612,N_10109,N_13965);
nor U17613 (N_17613,N_12943,N_12395);
or U17614 (N_17614,N_13891,N_10200);
nand U17615 (N_17615,N_14923,N_13951);
and U17616 (N_17616,N_13826,N_14049);
and U17617 (N_17617,N_11121,N_14582);
or U17618 (N_17618,N_13457,N_12413);
xor U17619 (N_17619,N_11222,N_11819);
and U17620 (N_17620,N_12986,N_11947);
xor U17621 (N_17621,N_14574,N_10598);
or U17622 (N_17622,N_14027,N_10307);
or U17623 (N_17623,N_14938,N_13031);
nor U17624 (N_17624,N_14884,N_10320);
and U17625 (N_17625,N_13745,N_13784);
nor U17626 (N_17626,N_11604,N_12635);
and U17627 (N_17627,N_13325,N_14225);
xor U17628 (N_17628,N_11859,N_10383);
nor U17629 (N_17629,N_12973,N_13736);
xor U17630 (N_17630,N_10323,N_10135);
and U17631 (N_17631,N_14599,N_14295);
xor U17632 (N_17632,N_12479,N_12406);
xnor U17633 (N_17633,N_11438,N_13644);
or U17634 (N_17634,N_14067,N_11555);
or U17635 (N_17635,N_12070,N_11361);
xnor U17636 (N_17636,N_14826,N_10904);
nor U17637 (N_17637,N_12731,N_13361);
nor U17638 (N_17638,N_14835,N_12472);
and U17639 (N_17639,N_10866,N_12866);
or U17640 (N_17640,N_11007,N_13841);
or U17641 (N_17641,N_13622,N_13719);
nand U17642 (N_17642,N_11645,N_13952);
and U17643 (N_17643,N_14950,N_10506);
or U17644 (N_17644,N_13154,N_11766);
nand U17645 (N_17645,N_11100,N_10899);
or U17646 (N_17646,N_14837,N_10864);
nand U17647 (N_17647,N_13464,N_13019);
and U17648 (N_17648,N_11522,N_11917);
and U17649 (N_17649,N_13906,N_14377);
xnor U17650 (N_17650,N_11054,N_10656);
nand U17651 (N_17651,N_11203,N_12838);
and U17652 (N_17652,N_12404,N_12107);
nor U17653 (N_17653,N_10828,N_14788);
nand U17654 (N_17654,N_12699,N_13579);
xnor U17655 (N_17655,N_12731,N_13648);
nand U17656 (N_17656,N_12515,N_11372);
nor U17657 (N_17657,N_14890,N_12134);
and U17658 (N_17658,N_12679,N_14542);
nor U17659 (N_17659,N_14938,N_10160);
or U17660 (N_17660,N_14599,N_12090);
nand U17661 (N_17661,N_10195,N_10778);
xor U17662 (N_17662,N_13235,N_13334);
nand U17663 (N_17663,N_11758,N_10723);
nand U17664 (N_17664,N_11350,N_10478);
or U17665 (N_17665,N_10133,N_12759);
nor U17666 (N_17666,N_13806,N_14628);
xnor U17667 (N_17667,N_13936,N_13185);
and U17668 (N_17668,N_11341,N_14922);
or U17669 (N_17669,N_13282,N_11106);
or U17670 (N_17670,N_11695,N_13990);
and U17671 (N_17671,N_13468,N_10109);
nor U17672 (N_17672,N_12966,N_13607);
nor U17673 (N_17673,N_11692,N_12168);
nor U17674 (N_17674,N_13603,N_14089);
and U17675 (N_17675,N_12647,N_11919);
and U17676 (N_17676,N_12860,N_10545);
or U17677 (N_17677,N_13881,N_13160);
and U17678 (N_17678,N_10930,N_12698);
or U17679 (N_17679,N_10100,N_13644);
and U17680 (N_17680,N_11671,N_11453);
nor U17681 (N_17681,N_14805,N_10443);
and U17682 (N_17682,N_13471,N_13883);
nor U17683 (N_17683,N_11407,N_13353);
nor U17684 (N_17684,N_14226,N_10728);
or U17685 (N_17685,N_10892,N_13117);
nor U17686 (N_17686,N_13378,N_10005);
and U17687 (N_17687,N_13041,N_11639);
or U17688 (N_17688,N_13105,N_13275);
nand U17689 (N_17689,N_10013,N_11235);
nand U17690 (N_17690,N_13142,N_11168);
or U17691 (N_17691,N_13833,N_13353);
nand U17692 (N_17692,N_14014,N_12521);
nand U17693 (N_17693,N_12198,N_13948);
nor U17694 (N_17694,N_11002,N_12635);
and U17695 (N_17695,N_10579,N_13599);
nor U17696 (N_17696,N_12145,N_12610);
or U17697 (N_17697,N_11839,N_12932);
and U17698 (N_17698,N_11184,N_11539);
nor U17699 (N_17699,N_13533,N_14317);
nand U17700 (N_17700,N_11618,N_12438);
or U17701 (N_17701,N_10362,N_11241);
and U17702 (N_17702,N_10450,N_14532);
nor U17703 (N_17703,N_10317,N_11445);
or U17704 (N_17704,N_10772,N_10653);
xor U17705 (N_17705,N_14073,N_11414);
and U17706 (N_17706,N_10014,N_14763);
nor U17707 (N_17707,N_13005,N_12367);
or U17708 (N_17708,N_12603,N_14318);
and U17709 (N_17709,N_14891,N_12678);
nor U17710 (N_17710,N_13112,N_13887);
and U17711 (N_17711,N_11024,N_10472);
xor U17712 (N_17712,N_12889,N_12267);
nor U17713 (N_17713,N_11581,N_10293);
and U17714 (N_17714,N_12681,N_10241);
nor U17715 (N_17715,N_11554,N_13131);
nand U17716 (N_17716,N_14768,N_10962);
and U17717 (N_17717,N_11925,N_14242);
nand U17718 (N_17718,N_13853,N_14124);
nor U17719 (N_17719,N_10411,N_10649);
and U17720 (N_17720,N_11566,N_14192);
and U17721 (N_17721,N_11021,N_11852);
nor U17722 (N_17722,N_11042,N_14653);
nor U17723 (N_17723,N_14420,N_14531);
nand U17724 (N_17724,N_11337,N_12121);
nand U17725 (N_17725,N_11875,N_13049);
and U17726 (N_17726,N_14050,N_11600);
xnor U17727 (N_17727,N_14548,N_13970);
nor U17728 (N_17728,N_12302,N_10751);
nor U17729 (N_17729,N_13224,N_11804);
and U17730 (N_17730,N_14354,N_11995);
nand U17731 (N_17731,N_10382,N_13393);
nand U17732 (N_17732,N_12892,N_12787);
nor U17733 (N_17733,N_10006,N_14679);
or U17734 (N_17734,N_11585,N_12040);
nand U17735 (N_17735,N_14571,N_10968);
and U17736 (N_17736,N_13906,N_14450);
or U17737 (N_17737,N_12332,N_11834);
or U17738 (N_17738,N_12204,N_13858);
nor U17739 (N_17739,N_10046,N_14513);
and U17740 (N_17740,N_11702,N_11989);
nor U17741 (N_17741,N_13083,N_10873);
and U17742 (N_17742,N_11056,N_12768);
nand U17743 (N_17743,N_10170,N_14033);
or U17744 (N_17744,N_13886,N_12990);
and U17745 (N_17745,N_12110,N_14367);
or U17746 (N_17746,N_13558,N_12717);
and U17747 (N_17747,N_11743,N_14635);
or U17748 (N_17748,N_10182,N_13034);
nor U17749 (N_17749,N_10951,N_13720);
or U17750 (N_17750,N_10403,N_12818);
xnor U17751 (N_17751,N_14143,N_13888);
xnor U17752 (N_17752,N_11040,N_11349);
and U17753 (N_17753,N_13610,N_10247);
or U17754 (N_17754,N_11394,N_10672);
nor U17755 (N_17755,N_10549,N_10596);
nor U17756 (N_17756,N_14942,N_13385);
xor U17757 (N_17757,N_10009,N_13125);
xnor U17758 (N_17758,N_13308,N_11015);
or U17759 (N_17759,N_14407,N_11415);
and U17760 (N_17760,N_13194,N_10433);
or U17761 (N_17761,N_13858,N_11285);
or U17762 (N_17762,N_10773,N_12440);
xnor U17763 (N_17763,N_10989,N_13854);
and U17764 (N_17764,N_11995,N_14112);
nor U17765 (N_17765,N_14664,N_14355);
or U17766 (N_17766,N_12797,N_14722);
nor U17767 (N_17767,N_14051,N_12232);
nand U17768 (N_17768,N_13292,N_11913);
and U17769 (N_17769,N_14705,N_11035);
and U17770 (N_17770,N_13200,N_12601);
xnor U17771 (N_17771,N_11629,N_13076);
nand U17772 (N_17772,N_14069,N_14450);
and U17773 (N_17773,N_10023,N_10505);
nand U17774 (N_17774,N_10401,N_10991);
or U17775 (N_17775,N_12839,N_10706);
xor U17776 (N_17776,N_13666,N_13417);
nor U17777 (N_17777,N_10575,N_14622);
and U17778 (N_17778,N_12415,N_14215);
or U17779 (N_17779,N_14186,N_12740);
and U17780 (N_17780,N_11798,N_12145);
nand U17781 (N_17781,N_11701,N_10242);
and U17782 (N_17782,N_14824,N_13747);
and U17783 (N_17783,N_10704,N_12307);
nor U17784 (N_17784,N_14887,N_13813);
nor U17785 (N_17785,N_13203,N_11847);
xnor U17786 (N_17786,N_11783,N_12868);
nor U17787 (N_17787,N_11666,N_14306);
xor U17788 (N_17788,N_10853,N_10894);
nand U17789 (N_17789,N_14379,N_10285);
or U17790 (N_17790,N_13752,N_10310);
nor U17791 (N_17791,N_10395,N_11670);
and U17792 (N_17792,N_10777,N_11652);
xor U17793 (N_17793,N_10767,N_13215);
nor U17794 (N_17794,N_13519,N_13400);
and U17795 (N_17795,N_10804,N_10603);
nand U17796 (N_17796,N_14555,N_12844);
nor U17797 (N_17797,N_14932,N_11843);
nor U17798 (N_17798,N_13986,N_10062);
or U17799 (N_17799,N_11580,N_10257);
nor U17800 (N_17800,N_12140,N_12565);
and U17801 (N_17801,N_14638,N_12546);
nor U17802 (N_17802,N_13508,N_10264);
and U17803 (N_17803,N_11153,N_11835);
or U17804 (N_17804,N_10425,N_10192);
and U17805 (N_17805,N_14623,N_11810);
nand U17806 (N_17806,N_13833,N_14468);
nand U17807 (N_17807,N_10256,N_12169);
or U17808 (N_17808,N_13232,N_12536);
or U17809 (N_17809,N_14813,N_14479);
nor U17810 (N_17810,N_13764,N_12549);
and U17811 (N_17811,N_14399,N_10815);
nand U17812 (N_17812,N_12119,N_12118);
and U17813 (N_17813,N_14162,N_14638);
or U17814 (N_17814,N_13051,N_12093);
xnor U17815 (N_17815,N_10433,N_14934);
nor U17816 (N_17816,N_10276,N_11029);
or U17817 (N_17817,N_12048,N_10042);
and U17818 (N_17818,N_14898,N_13641);
nor U17819 (N_17819,N_11958,N_11796);
and U17820 (N_17820,N_14696,N_13638);
nand U17821 (N_17821,N_14805,N_10855);
and U17822 (N_17822,N_13566,N_11227);
nor U17823 (N_17823,N_12668,N_12302);
nor U17824 (N_17824,N_14421,N_13687);
or U17825 (N_17825,N_14558,N_12139);
and U17826 (N_17826,N_11432,N_14917);
or U17827 (N_17827,N_13699,N_11062);
nor U17828 (N_17828,N_12150,N_13718);
xor U17829 (N_17829,N_10002,N_10858);
xnor U17830 (N_17830,N_12097,N_12081);
nand U17831 (N_17831,N_10881,N_12341);
nand U17832 (N_17832,N_11247,N_13475);
or U17833 (N_17833,N_14590,N_10746);
and U17834 (N_17834,N_10245,N_11475);
nand U17835 (N_17835,N_10282,N_12920);
and U17836 (N_17836,N_10268,N_11021);
xor U17837 (N_17837,N_11570,N_14711);
nor U17838 (N_17838,N_12628,N_13755);
or U17839 (N_17839,N_10858,N_11607);
or U17840 (N_17840,N_11033,N_12279);
nor U17841 (N_17841,N_10554,N_13547);
nor U17842 (N_17842,N_11088,N_12329);
and U17843 (N_17843,N_14324,N_12125);
and U17844 (N_17844,N_12867,N_14087);
nor U17845 (N_17845,N_12425,N_11826);
nand U17846 (N_17846,N_11617,N_14904);
nor U17847 (N_17847,N_13941,N_10362);
nor U17848 (N_17848,N_14540,N_11424);
and U17849 (N_17849,N_12640,N_12251);
or U17850 (N_17850,N_12833,N_12428);
or U17851 (N_17851,N_12505,N_13851);
and U17852 (N_17852,N_14729,N_12261);
or U17853 (N_17853,N_14712,N_10258);
or U17854 (N_17854,N_10007,N_13500);
or U17855 (N_17855,N_11022,N_10306);
or U17856 (N_17856,N_14088,N_11303);
nor U17857 (N_17857,N_14562,N_13743);
and U17858 (N_17858,N_11743,N_11939);
nand U17859 (N_17859,N_10107,N_14615);
nor U17860 (N_17860,N_12488,N_12371);
nand U17861 (N_17861,N_13002,N_12250);
or U17862 (N_17862,N_12521,N_11946);
nor U17863 (N_17863,N_14425,N_13482);
xor U17864 (N_17864,N_13638,N_11798);
or U17865 (N_17865,N_11351,N_12139);
xnor U17866 (N_17866,N_10481,N_12831);
nor U17867 (N_17867,N_14474,N_11302);
nand U17868 (N_17868,N_11768,N_12367);
xnor U17869 (N_17869,N_13065,N_13539);
nand U17870 (N_17870,N_11336,N_10550);
nor U17871 (N_17871,N_12742,N_13569);
or U17872 (N_17872,N_13966,N_12966);
xor U17873 (N_17873,N_14087,N_13243);
nor U17874 (N_17874,N_12117,N_14203);
and U17875 (N_17875,N_11243,N_10763);
and U17876 (N_17876,N_12054,N_14858);
and U17877 (N_17877,N_10485,N_11546);
or U17878 (N_17878,N_12937,N_14482);
or U17879 (N_17879,N_11954,N_10468);
nand U17880 (N_17880,N_10435,N_13160);
nand U17881 (N_17881,N_13087,N_12339);
or U17882 (N_17882,N_12459,N_10972);
nand U17883 (N_17883,N_13548,N_13828);
and U17884 (N_17884,N_13749,N_10373);
or U17885 (N_17885,N_13058,N_14969);
xor U17886 (N_17886,N_13405,N_13907);
and U17887 (N_17887,N_11143,N_13369);
nand U17888 (N_17888,N_13714,N_14943);
or U17889 (N_17889,N_11593,N_10440);
or U17890 (N_17890,N_11176,N_14676);
xor U17891 (N_17891,N_14287,N_10520);
nand U17892 (N_17892,N_13351,N_10042);
nor U17893 (N_17893,N_10377,N_12528);
and U17894 (N_17894,N_11501,N_11601);
nor U17895 (N_17895,N_12897,N_10836);
nor U17896 (N_17896,N_10469,N_14804);
nor U17897 (N_17897,N_10711,N_13496);
or U17898 (N_17898,N_12584,N_11061);
and U17899 (N_17899,N_13275,N_14133);
nand U17900 (N_17900,N_10983,N_13445);
nand U17901 (N_17901,N_10878,N_11693);
nand U17902 (N_17902,N_11095,N_13277);
nand U17903 (N_17903,N_14819,N_14959);
xnor U17904 (N_17904,N_14655,N_10540);
or U17905 (N_17905,N_14414,N_11997);
nor U17906 (N_17906,N_11827,N_10007);
nor U17907 (N_17907,N_13233,N_10469);
nand U17908 (N_17908,N_13093,N_13869);
nand U17909 (N_17909,N_14062,N_14429);
nor U17910 (N_17910,N_13987,N_12380);
nand U17911 (N_17911,N_10390,N_10553);
and U17912 (N_17912,N_14905,N_14470);
and U17913 (N_17913,N_13202,N_11389);
or U17914 (N_17914,N_13466,N_10713);
xnor U17915 (N_17915,N_14598,N_14021);
nand U17916 (N_17916,N_10004,N_13605);
nor U17917 (N_17917,N_13581,N_14729);
and U17918 (N_17918,N_12091,N_14593);
and U17919 (N_17919,N_12628,N_11898);
nand U17920 (N_17920,N_13800,N_13735);
nor U17921 (N_17921,N_12029,N_12047);
nor U17922 (N_17922,N_10846,N_14321);
nor U17923 (N_17923,N_10316,N_13560);
or U17924 (N_17924,N_10541,N_12918);
nand U17925 (N_17925,N_13726,N_13044);
or U17926 (N_17926,N_10010,N_12415);
and U17927 (N_17927,N_12591,N_14209);
nor U17928 (N_17928,N_13427,N_12427);
xor U17929 (N_17929,N_12859,N_11762);
nand U17930 (N_17930,N_10526,N_14951);
and U17931 (N_17931,N_10020,N_12770);
nand U17932 (N_17932,N_10554,N_11511);
nand U17933 (N_17933,N_12393,N_10272);
nand U17934 (N_17934,N_11312,N_13051);
and U17935 (N_17935,N_12926,N_13302);
nand U17936 (N_17936,N_13071,N_12701);
nand U17937 (N_17937,N_10333,N_14270);
or U17938 (N_17938,N_14033,N_12291);
nand U17939 (N_17939,N_12078,N_10696);
or U17940 (N_17940,N_11584,N_13383);
nand U17941 (N_17941,N_10808,N_12891);
or U17942 (N_17942,N_12033,N_12019);
and U17943 (N_17943,N_11748,N_13463);
nand U17944 (N_17944,N_11795,N_11864);
or U17945 (N_17945,N_11954,N_12496);
or U17946 (N_17946,N_13477,N_14414);
or U17947 (N_17947,N_11881,N_12554);
or U17948 (N_17948,N_11304,N_14100);
nand U17949 (N_17949,N_10208,N_14375);
nand U17950 (N_17950,N_11731,N_14944);
and U17951 (N_17951,N_13866,N_14517);
nand U17952 (N_17952,N_12020,N_12811);
nor U17953 (N_17953,N_11712,N_10024);
xnor U17954 (N_17954,N_11528,N_11328);
and U17955 (N_17955,N_11859,N_14809);
nor U17956 (N_17956,N_10493,N_11537);
and U17957 (N_17957,N_11729,N_14943);
or U17958 (N_17958,N_11092,N_12884);
nor U17959 (N_17959,N_13580,N_12670);
nand U17960 (N_17960,N_11536,N_13090);
and U17961 (N_17961,N_14729,N_12127);
or U17962 (N_17962,N_14406,N_14606);
xor U17963 (N_17963,N_12787,N_10123);
xor U17964 (N_17964,N_12931,N_11194);
nor U17965 (N_17965,N_10461,N_14130);
nand U17966 (N_17966,N_14393,N_11944);
nor U17967 (N_17967,N_13531,N_11732);
nor U17968 (N_17968,N_12675,N_14630);
nor U17969 (N_17969,N_10099,N_13071);
xor U17970 (N_17970,N_11200,N_10143);
nand U17971 (N_17971,N_13713,N_12425);
nor U17972 (N_17972,N_12052,N_11562);
nand U17973 (N_17973,N_11817,N_10230);
and U17974 (N_17974,N_10430,N_11727);
nor U17975 (N_17975,N_11358,N_11317);
and U17976 (N_17976,N_14630,N_12473);
nand U17977 (N_17977,N_10783,N_12609);
xor U17978 (N_17978,N_12582,N_12153);
nand U17979 (N_17979,N_14065,N_11812);
xnor U17980 (N_17980,N_10568,N_10290);
nor U17981 (N_17981,N_13601,N_13694);
and U17982 (N_17982,N_10959,N_12172);
nand U17983 (N_17983,N_11313,N_11985);
or U17984 (N_17984,N_11561,N_13588);
nor U17985 (N_17985,N_11556,N_12495);
xor U17986 (N_17986,N_12663,N_12721);
nor U17987 (N_17987,N_13138,N_12016);
nand U17988 (N_17988,N_13873,N_10300);
nand U17989 (N_17989,N_10544,N_12924);
nand U17990 (N_17990,N_10345,N_10025);
or U17991 (N_17991,N_13395,N_10965);
xnor U17992 (N_17992,N_11126,N_14855);
and U17993 (N_17993,N_11679,N_10575);
and U17994 (N_17994,N_10761,N_11227);
nor U17995 (N_17995,N_12516,N_13148);
nand U17996 (N_17996,N_10640,N_12875);
nand U17997 (N_17997,N_13996,N_12788);
and U17998 (N_17998,N_13285,N_13995);
or U17999 (N_17999,N_10480,N_14749);
and U18000 (N_18000,N_11600,N_11930);
nor U18001 (N_18001,N_10752,N_11692);
nor U18002 (N_18002,N_14312,N_10596);
or U18003 (N_18003,N_10549,N_10063);
nand U18004 (N_18004,N_13129,N_14158);
nand U18005 (N_18005,N_14355,N_11950);
or U18006 (N_18006,N_11739,N_14495);
or U18007 (N_18007,N_10406,N_11499);
or U18008 (N_18008,N_12001,N_13403);
and U18009 (N_18009,N_10010,N_14812);
nor U18010 (N_18010,N_10690,N_11758);
or U18011 (N_18011,N_11542,N_14069);
or U18012 (N_18012,N_12043,N_12875);
or U18013 (N_18013,N_13672,N_12681);
or U18014 (N_18014,N_10620,N_11882);
or U18015 (N_18015,N_11937,N_11792);
xnor U18016 (N_18016,N_11075,N_12153);
nand U18017 (N_18017,N_13842,N_11644);
or U18018 (N_18018,N_13269,N_12557);
nand U18019 (N_18019,N_13965,N_13487);
nor U18020 (N_18020,N_12205,N_10564);
or U18021 (N_18021,N_12363,N_13473);
and U18022 (N_18022,N_11982,N_13234);
or U18023 (N_18023,N_12365,N_11724);
or U18024 (N_18024,N_12955,N_13892);
nand U18025 (N_18025,N_11606,N_13025);
and U18026 (N_18026,N_10649,N_14578);
and U18027 (N_18027,N_10357,N_13432);
and U18028 (N_18028,N_10060,N_12810);
or U18029 (N_18029,N_12981,N_12124);
nand U18030 (N_18030,N_12256,N_11904);
nand U18031 (N_18031,N_10590,N_14695);
nor U18032 (N_18032,N_12577,N_10738);
nand U18033 (N_18033,N_10707,N_10991);
nand U18034 (N_18034,N_10366,N_13665);
nand U18035 (N_18035,N_13527,N_14520);
nand U18036 (N_18036,N_12770,N_10090);
nand U18037 (N_18037,N_12486,N_12452);
or U18038 (N_18038,N_11220,N_12731);
nand U18039 (N_18039,N_12718,N_12664);
or U18040 (N_18040,N_14033,N_13052);
nor U18041 (N_18041,N_12329,N_10933);
nor U18042 (N_18042,N_10769,N_13440);
nand U18043 (N_18043,N_10631,N_13816);
nand U18044 (N_18044,N_10256,N_12972);
or U18045 (N_18045,N_10269,N_12931);
nand U18046 (N_18046,N_12825,N_11358);
nand U18047 (N_18047,N_13966,N_14477);
or U18048 (N_18048,N_13078,N_14923);
and U18049 (N_18049,N_12249,N_12877);
and U18050 (N_18050,N_13223,N_11303);
nand U18051 (N_18051,N_14832,N_14794);
nor U18052 (N_18052,N_10443,N_12855);
or U18053 (N_18053,N_13212,N_12315);
nand U18054 (N_18054,N_11546,N_10446);
xor U18055 (N_18055,N_13179,N_10044);
xnor U18056 (N_18056,N_14204,N_13225);
and U18057 (N_18057,N_12082,N_11452);
nand U18058 (N_18058,N_10921,N_13001);
nor U18059 (N_18059,N_14526,N_12518);
or U18060 (N_18060,N_12418,N_12832);
or U18061 (N_18061,N_12674,N_12207);
nand U18062 (N_18062,N_13840,N_11954);
nand U18063 (N_18063,N_10538,N_13605);
xnor U18064 (N_18064,N_12427,N_14860);
nor U18065 (N_18065,N_13191,N_10134);
or U18066 (N_18066,N_14623,N_12963);
nor U18067 (N_18067,N_12618,N_10945);
and U18068 (N_18068,N_11642,N_10516);
nand U18069 (N_18069,N_10437,N_11242);
or U18070 (N_18070,N_10734,N_11218);
or U18071 (N_18071,N_12351,N_13589);
nand U18072 (N_18072,N_10295,N_10923);
nor U18073 (N_18073,N_10858,N_14114);
nor U18074 (N_18074,N_10780,N_12100);
and U18075 (N_18075,N_10581,N_13976);
nand U18076 (N_18076,N_14872,N_14622);
nand U18077 (N_18077,N_10020,N_10760);
or U18078 (N_18078,N_11345,N_10073);
or U18079 (N_18079,N_13759,N_13880);
or U18080 (N_18080,N_13402,N_12447);
nand U18081 (N_18081,N_12740,N_14145);
nand U18082 (N_18082,N_11122,N_10613);
nand U18083 (N_18083,N_11647,N_13818);
nand U18084 (N_18084,N_14945,N_11099);
xnor U18085 (N_18085,N_11872,N_14931);
nor U18086 (N_18086,N_14297,N_14174);
and U18087 (N_18087,N_11174,N_14778);
and U18088 (N_18088,N_13288,N_14080);
nand U18089 (N_18089,N_11984,N_10899);
nand U18090 (N_18090,N_12670,N_14518);
and U18091 (N_18091,N_14449,N_10158);
and U18092 (N_18092,N_12785,N_14059);
nor U18093 (N_18093,N_11177,N_10714);
nor U18094 (N_18094,N_12456,N_11478);
xor U18095 (N_18095,N_11612,N_13875);
nor U18096 (N_18096,N_11166,N_13892);
and U18097 (N_18097,N_12054,N_14355);
nor U18098 (N_18098,N_13820,N_13285);
and U18099 (N_18099,N_11157,N_10249);
nor U18100 (N_18100,N_13113,N_12077);
xor U18101 (N_18101,N_10605,N_11004);
or U18102 (N_18102,N_13121,N_11275);
or U18103 (N_18103,N_11749,N_14724);
and U18104 (N_18104,N_12957,N_11461);
nor U18105 (N_18105,N_12771,N_14852);
and U18106 (N_18106,N_12661,N_13528);
nor U18107 (N_18107,N_10110,N_14494);
and U18108 (N_18108,N_10777,N_10357);
nand U18109 (N_18109,N_13039,N_13193);
nand U18110 (N_18110,N_14253,N_10480);
nand U18111 (N_18111,N_13677,N_10888);
and U18112 (N_18112,N_10856,N_12496);
nor U18113 (N_18113,N_14458,N_11914);
or U18114 (N_18114,N_14190,N_10431);
or U18115 (N_18115,N_14897,N_14263);
nand U18116 (N_18116,N_11865,N_13803);
nor U18117 (N_18117,N_14542,N_14412);
or U18118 (N_18118,N_14401,N_14735);
nor U18119 (N_18119,N_10165,N_13145);
xor U18120 (N_18120,N_13540,N_11497);
or U18121 (N_18121,N_14380,N_12950);
xor U18122 (N_18122,N_12541,N_11690);
or U18123 (N_18123,N_13944,N_12857);
xor U18124 (N_18124,N_14143,N_12467);
nand U18125 (N_18125,N_11532,N_11481);
nand U18126 (N_18126,N_14980,N_11800);
nor U18127 (N_18127,N_13124,N_11868);
nor U18128 (N_18128,N_13384,N_11217);
and U18129 (N_18129,N_14580,N_10101);
nand U18130 (N_18130,N_11881,N_10030);
and U18131 (N_18131,N_13278,N_14554);
nor U18132 (N_18132,N_10316,N_10367);
and U18133 (N_18133,N_11853,N_14826);
and U18134 (N_18134,N_13826,N_14211);
or U18135 (N_18135,N_12239,N_11933);
xnor U18136 (N_18136,N_10066,N_10436);
nor U18137 (N_18137,N_10652,N_10680);
and U18138 (N_18138,N_12262,N_13035);
nand U18139 (N_18139,N_13450,N_11844);
and U18140 (N_18140,N_11040,N_11516);
nand U18141 (N_18141,N_13139,N_10485);
or U18142 (N_18142,N_14850,N_12595);
nor U18143 (N_18143,N_14477,N_12457);
or U18144 (N_18144,N_14185,N_14559);
and U18145 (N_18145,N_13984,N_10036);
and U18146 (N_18146,N_11389,N_13069);
and U18147 (N_18147,N_11270,N_12355);
nand U18148 (N_18148,N_13755,N_13950);
or U18149 (N_18149,N_13871,N_12172);
or U18150 (N_18150,N_11147,N_12423);
or U18151 (N_18151,N_10548,N_11288);
or U18152 (N_18152,N_11617,N_12873);
nor U18153 (N_18153,N_10364,N_10499);
nor U18154 (N_18154,N_14763,N_13939);
nor U18155 (N_18155,N_10198,N_14043);
or U18156 (N_18156,N_11917,N_14162);
and U18157 (N_18157,N_11852,N_13498);
xor U18158 (N_18158,N_10936,N_10869);
nor U18159 (N_18159,N_13953,N_13859);
nor U18160 (N_18160,N_14145,N_10628);
and U18161 (N_18161,N_11268,N_14143);
nand U18162 (N_18162,N_12112,N_13747);
nor U18163 (N_18163,N_14305,N_10279);
nand U18164 (N_18164,N_14040,N_13421);
nor U18165 (N_18165,N_10465,N_14134);
nor U18166 (N_18166,N_13285,N_10715);
or U18167 (N_18167,N_12608,N_10343);
or U18168 (N_18168,N_12698,N_11163);
or U18169 (N_18169,N_12539,N_14712);
nor U18170 (N_18170,N_13571,N_10963);
xor U18171 (N_18171,N_11457,N_11622);
nand U18172 (N_18172,N_12599,N_11231);
nand U18173 (N_18173,N_11581,N_11749);
xor U18174 (N_18174,N_11076,N_11703);
xor U18175 (N_18175,N_10672,N_13178);
nand U18176 (N_18176,N_13197,N_10902);
xnor U18177 (N_18177,N_13800,N_11163);
and U18178 (N_18178,N_13762,N_13197);
or U18179 (N_18179,N_14039,N_10027);
nand U18180 (N_18180,N_11951,N_12682);
or U18181 (N_18181,N_13570,N_10775);
or U18182 (N_18182,N_14416,N_12329);
nor U18183 (N_18183,N_13728,N_14120);
nand U18184 (N_18184,N_13856,N_12169);
nand U18185 (N_18185,N_13895,N_11886);
or U18186 (N_18186,N_14013,N_11644);
and U18187 (N_18187,N_11341,N_11432);
nand U18188 (N_18188,N_10653,N_12493);
and U18189 (N_18189,N_14005,N_10855);
and U18190 (N_18190,N_10359,N_11470);
nand U18191 (N_18191,N_10330,N_12407);
and U18192 (N_18192,N_11251,N_12138);
and U18193 (N_18193,N_10648,N_13046);
and U18194 (N_18194,N_12318,N_11717);
or U18195 (N_18195,N_10446,N_10946);
and U18196 (N_18196,N_14836,N_12575);
xnor U18197 (N_18197,N_12555,N_11758);
nand U18198 (N_18198,N_14355,N_12238);
and U18199 (N_18199,N_12166,N_13856);
xnor U18200 (N_18200,N_13099,N_14656);
nand U18201 (N_18201,N_12239,N_11799);
or U18202 (N_18202,N_11881,N_14415);
or U18203 (N_18203,N_12154,N_13664);
nor U18204 (N_18204,N_14528,N_10382);
or U18205 (N_18205,N_11647,N_11170);
and U18206 (N_18206,N_12743,N_13207);
xor U18207 (N_18207,N_11966,N_12779);
nor U18208 (N_18208,N_13088,N_12955);
or U18209 (N_18209,N_10570,N_11769);
or U18210 (N_18210,N_12463,N_10608);
nand U18211 (N_18211,N_14817,N_10128);
and U18212 (N_18212,N_11444,N_14468);
or U18213 (N_18213,N_11858,N_14618);
and U18214 (N_18214,N_12063,N_11040);
nand U18215 (N_18215,N_11693,N_10162);
nand U18216 (N_18216,N_14376,N_11352);
or U18217 (N_18217,N_14312,N_13525);
or U18218 (N_18218,N_11022,N_14015);
nor U18219 (N_18219,N_12401,N_10308);
xnor U18220 (N_18220,N_12709,N_14298);
nand U18221 (N_18221,N_10544,N_11707);
or U18222 (N_18222,N_10773,N_14853);
or U18223 (N_18223,N_11208,N_11330);
xnor U18224 (N_18224,N_13815,N_12658);
nand U18225 (N_18225,N_12819,N_12836);
nor U18226 (N_18226,N_14247,N_14762);
or U18227 (N_18227,N_12273,N_14585);
or U18228 (N_18228,N_14429,N_12119);
or U18229 (N_18229,N_11762,N_10645);
xnor U18230 (N_18230,N_13480,N_10485);
nor U18231 (N_18231,N_11036,N_11881);
nand U18232 (N_18232,N_11963,N_12971);
or U18233 (N_18233,N_11324,N_12724);
nor U18234 (N_18234,N_10518,N_10480);
and U18235 (N_18235,N_10440,N_11851);
xor U18236 (N_18236,N_11465,N_10464);
nand U18237 (N_18237,N_11873,N_10728);
and U18238 (N_18238,N_10759,N_13762);
nor U18239 (N_18239,N_11563,N_12496);
and U18240 (N_18240,N_14704,N_11050);
and U18241 (N_18241,N_13781,N_11625);
nand U18242 (N_18242,N_13718,N_11327);
nor U18243 (N_18243,N_14590,N_12889);
or U18244 (N_18244,N_14896,N_14889);
and U18245 (N_18245,N_12612,N_13441);
nand U18246 (N_18246,N_12745,N_12638);
or U18247 (N_18247,N_11902,N_13422);
and U18248 (N_18248,N_14278,N_13693);
xnor U18249 (N_18249,N_13081,N_12952);
or U18250 (N_18250,N_14704,N_13495);
xnor U18251 (N_18251,N_13390,N_10855);
or U18252 (N_18252,N_12782,N_11288);
and U18253 (N_18253,N_12970,N_12808);
or U18254 (N_18254,N_11666,N_12457);
and U18255 (N_18255,N_11603,N_12806);
nor U18256 (N_18256,N_14153,N_13752);
or U18257 (N_18257,N_11968,N_12942);
nand U18258 (N_18258,N_13108,N_14158);
or U18259 (N_18259,N_10235,N_12937);
or U18260 (N_18260,N_10236,N_12871);
nor U18261 (N_18261,N_12993,N_12531);
nand U18262 (N_18262,N_10950,N_10938);
or U18263 (N_18263,N_10938,N_10966);
and U18264 (N_18264,N_11105,N_12682);
nor U18265 (N_18265,N_12488,N_12892);
and U18266 (N_18266,N_10874,N_10304);
nand U18267 (N_18267,N_14440,N_12264);
or U18268 (N_18268,N_12680,N_11836);
nor U18269 (N_18269,N_12584,N_14074);
nor U18270 (N_18270,N_13305,N_10926);
xor U18271 (N_18271,N_14173,N_11051);
xnor U18272 (N_18272,N_11159,N_11746);
or U18273 (N_18273,N_10772,N_11459);
nor U18274 (N_18274,N_10077,N_13722);
nor U18275 (N_18275,N_14488,N_10377);
or U18276 (N_18276,N_14381,N_12316);
and U18277 (N_18277,N_10303,N_14465);
or U18278 (N_18278,N_14017,N_12787);
or U18279 (N_18279,N_12320,N_14652);
xor U18280 (N_18280,N_10148,N_14882);
or U18281 (N_18281,N_14366,N_10876);
nor U18282 (N_18282,N_12199,N_10721);
nor U18283 (N_18283,N_13146,N_11796);
nand U18284 (N_18284,N_11167,N_11024);
nand U18285 (N_18285,N_14987,N_13543);
nand U18286 (N_18286,N_12733,N_13495);
xnor U18287 (N_18287,N_13483,N_13341);
and U18288 (N_18288,N_14389,N_12167);
nor U18289 (N_18289,N_12641,N_12049);
and U18290 (N_18290,N_13086,N_12316);
nor U18291 (N_18291,N_10908,N_11512);
and U18292 (N_18292,N_12585,N_13810);
or U18293 (N_18293,N_14477,N_13982);
or U18294 (N_18294,N_12065,N_13517);
nor U18295 (N_18295,N_14011,N_11434);
or U18296 (N_18296,N_14351,N_11693);
nor U18297 (N_18297,N_11047,N_12399);
nand U18298 (N_18298,N_12030,N_14982);
xnor U18299 (N_18299,N_11285,N_11792);
nand U18300 (N_18300,N_13657,N_14096);
or U18301 (N_18301,N_14535,N_10885);
nand U18302 (N_18302,N_10339,N_10190);
or U18303 (N_18303,N_13180,N_14846);
xor U18304 (N_18304,N_11956,N_10702);
xnor U18305 (N_18305,N_13980,N_12347);
and U18306 (N_18306,N_10908,N_12708);
nor U18307 (N_18307,N_13999,N_11331);
nor U18308 (N_18308,N_14722,N_10981);
and U18309 (N_18309,N_10705,N_10764);
or U18310 (N_18310,N_12887,N_14030);
nor U18311 (N_18311,N_12935,N_10663);
or U18312 (N_18312,N_10735,N_10782);
xor U18313 (N_18313,N_12084,N_12978);
or U18314 (N_18314,N_10237,N_12957);
nor U18315 (N_18315,N_10880,N_10688);
or U18316 (N_18316,N_12597,N_11610);
nor U18317 (N_18317,N_14532,N_11116);
xnor U18318 (N_18318,N_10253,N_13221);
nand U18319 (N_18319,N_13247,N_14268);
or U18320 (N_18320,N_11048,N_12052);
nor U18321 (N_18321,N_10390,N_10454);
nand U18322 (N_18322,N_14871,N_10342);
nand U18323 (N_18323,N_12103,N_10056);
and U18324 (N_18324,N_11075,N_10986);
and U18325 (N_18325,N_14480,N_10588);
or U18326 (N_18326,N_14100,N_13758);
xnor U18327 (N_18327,N_12731,N_11190);
or U18328 (N_18328,N_11908,N_13644);
nand U18329 (N_18329,N_13734,N_10057);
or U18330 (N_18330,N_13296,N_10240);
nand U18331 (N_18331,N_11281,N_12317);
and U18332 (N_18332,N_13782,N_14398);
nand U18333 (N_18333,N_11631,N_13590);
nand U18334 (N_18334,N_10443,N_11754);
and U18335 (N_18335,N_10378,N_14212);
and U18336 (N_18336,N_14461,N_14656);
or U18337 (N_18337,N_12691,N_13363);
nand U18338 (N_18338,N_10586,N_14983);
xnor U18339 (N_18339,N_12561,N_11181);
or U18340 (N_18340,N_13245,N_14822);
xnor U18341 (N_18341,N_13237,N_14338);
nor U18342 (N_18342,N_11563,N_12518);
or U18343 (N_18343,N_12038,N_14307);
xnor U18344 (N_18344,N_11194,N_13354);
nor U18345 (N_18345,N_12841,N_12263);
or U18346 (N_18346,N_10412,N_14861);
and U18347 (N_18347,N_12746,N_14913);
and U18348 (N_18348,N_10602,N_12554);
or U18349 (N_18349,N_14707,N_13458);
nor U18350 (N_18350,N_11415,N_14586);
nand U18351 (N_18351,N_14748,N_12831);
and U18352 (N_18352,N_11573,N_10237);
nor U18353 (N_18353,N_10475,N_10133);
and U18354 (N_18354,N_12636,N_13530);
or U18355 (N_18355,N_11669,N_14350);
and U18356 (N_18356,N_11942,N_14411);
or U18357 (N_18357,N_12056,N_12479);
xor U18358 (N_18358,N_12699,N_10668);
and U18359 (N_18359,N_13390,N_14638);
or U18360 (N_18360,N_13748,N_10070);
nand U18361 (N_18361,N_12763,N_11181);
nor U18362 (N_18362,N_12215,N_14195);
nand U18363 (N_18363,N_13008,N_12033);
nor U18364 (N_18364,N_11663,N_10680);
or U18365 (N_18365,N_11560,N_13307);
and U18366 (N_18366,N_12439,N_12066);
nor U18367 (N_18367,N_11718,N_14202);
and U18368 (N_18368,N_11429,N_10785);
xnor U18369 (N_18369,N_10265,N_10471);
and U18370 (N_18370,N_14043,N_13454);
nor U18371 (N_18371,N_10362,N_13579);
and U18372 (N_18372,N_14628,N_11356);
nand U18373 (N_18373,N_14716,N_13814);
nor U18374 (N_18374,N_14241,N_10210);
and U18375 (N_18375,N_13473,N_14008);
and U18376 (N_18376,N_13889,N_11569);
and U18377 (N_18377,N_14869,N_14808);
and U18378 (N_18378,N_12293,N_14019);
nor U18379 (N_18379,N_14783,N_13660);
or U18380 (N_18380,N_11236,N_10740);
nor U18381 (N_18381,N_12912,N_13641);
nand U18382 (N_18382,N_12374,N_14345);
nand U18383 (N_18383,N_14611,N_14906);
or U18384 (N_18384,N_13586,N_10160);
nor U18385 (N_18385,N_12160,N_14045);
or U18386 (N_18386,N_10229,N_13056);
nand U18387 (N_18387,N_10172,N_13708);
or U18388 (N_18388,N_13037,N_11852);
nand U18389 (N_18389,N_13310,N_12565);
and U18390 (N_18390,N_11332,N_13832);
nor U18391 (N_18391,N_10242,N_11920);
xnor U18392 (N_18392,N_14966,N_12498);
or U18393 (N_18393,N_10459,N_10322);
or U18394 (N_18394,N_11120,N_13604);
and U18395 (N_18395,N_14894,N_13560);
or U18396 (N_18396,N_14723,N_13697);
xnor U18397 (N_18397,N_11795,N_11561);
nand U18398 (N_18398,N_10510,N_11975);
or U18399 (N_18399,N_14368,N_14534);
xor U18400 (N_18400,N_11748,N_10754);
and U18401 (N_18401,N_11844,N_13577);
and U18402 (N_18402,N_13756,N_13610);
or U18403 (N_18403,N_13769,N_11930);
nor U18404 (N_18404,N_12225,N_11253);
xnor U18405 (N_18405,N_11022,N_12450);
nand U18406 (N_18406,N_13335,N_13247);
nor U18407 (N_18407,N_10414,N_13351);
nand U18408 (N_18408,N_12168,N_13047);
nand U18409 (N_18409,N_13514,N_11131);
nor U18410 (N_18410,N_11650,N_12996);
and U18411 (N_18411,N_10522,N_12087);
or U18412 (N_18412,N_10293,N_14350);
and U18413 (N_18413,N_12338,N_12022);
nor U18414 (N_18414,N_10207,N_12833);
or U18415 (N_18415,N_10840,N_11315);
nand U18416 (N_18416,N_12579,N_13500);
nor U18417 (N_18417,N_14133,N_14979);
nand U18418 (N_18418,N_13208,N_14938);
or U18419 (N_18419,N_10377,N_11136);
and U18420 (N_18420,N_10520,N_11891);
nor U18421 (N_18421,N_14577,N_11937);
nand U18422 (N_18422,N_10932,N_14889);
or U18423 (N_18423,N_12383,N_10764);
nor U18424 (N_18424,N_13919,N_13325);
and U18425 (N_18425,N_13034,N_12534);
nand U18426 (N_18426,N_12851,N_11555);
nand U18427 (N_18427,N_14670,N_13043);
xnor U18428 (N_18428,N_10211,N_13117);
and U18429 (N_18429,N_12337,N_10803);
nand U18430 (N_18430,N_14938,N_10711);
nand U18431 (N_18431,N_14928,N_14568);
nand U18432 (N_18432,N_14093,N_14873);
and U18433 (N_18433,N_14779,N_12000);
xor U18434 (N_18434,N_10493,N_11728);
or U18435 (N_18435,N_10039,N_12461);
xnor U18436 (N_18436,N_14343,N_12247);
or U18437 (N_18437,N_13988,N_13620);
nor U18438 (N_18438,N_13583,N_13479);
nor U18439 (N_18439,N_13198,N_12537);
nand U18440 (N_18440,N_14890,N_13834);
or U18441 (N_18441,N_13245,N_11672);
or U18442 (N_18442,N_10141,N_11790);
or U18443 (N_18443,N_12649,N_13788);
nand U18444 (N_18444,N_12199,N_13384);
nor U18445 (N_18445,N_10871,N_13215);
or U18446 (N_18446,N_12247,N_12044);
xnor U18447 (N_18447,N_13584,N_11164);
nand U18448 (N_18448,N_10602,N_14980);
or U18449 (N_18449,N_11390,N_12753);
nor U18450 (N_18450,N_11218,N_12848);
and U18451 (N_18451,N_13307,N_11173);
nand U18452 (N_18452,N_13244,N_12783);
or U18453 (N_18453,N_14849,N_12959);
or U18454 (N_18454,N_10309,N_12400);
or U18455 (N_18455,N_10912,N_11912);
and U18456 (N_18456,N_12245,N_10208);
nand U18457 (N_18457,N_12326,N_12095);
nor U18458 (N_18458,N_10815,N_10767);
and U18459 (N_18459,N_14585,N_14842);
xor U18460 (N_18460,N_13532,N_11387);
xor U18461 (N_18461,N_12019,N_14701);
or U18462 (N_18462,N_14271,N_12207);
or U18463 (N_18463,N_12368,N_13134);
xnor U18464 (N_18464,N_10671,N_10727);
nor U18465 (N_18465,N_11453,N_14061);
nand U18466 (N_18466,N_14629,N_12605);
nand U18467 (N_18467,N_11528,N_12695);
and U18468 (N_18468,N_12303,N_14741);
and U18469 (N_18469,N_14097,N_13693);
nor U18470 (N_18470,N_12809,N_14250);
nor U18471 (N_18471,N_10449,N_12527);
and U18472 (N_18472,N_14664,N_11515);
or U18473 (N_18473,N_10447,N_10348);
nor U18474 (N_18474,N_10037,N_14119);
or U18475 (N_18475,N_10332,N_12353);
xnor U18476 (N_18476,N_11240,N_14391);
and U18477 (N_18477,N_12849,N_12502);
and U18478 (N_18478,N_12787,N_11006);
and U18479 (N_18479,N_11606,N_11834);
xor U18480 (N_18480,N_11869,N_14425);
xnor U18481 (N_18481,N_12393,N_10011);
nand U18482 (N_18482,N_13115,N_13053);
nor U18483 (N_18483,N_14931,N_11455);
nor U18484 (N_18484,N_12622,N_14869);
nor U18485 (N_18485,N_13455,N_11450);
nand U18486 (N_18486,N_11872,N_10000);
and U18487 (N_18487,N_12610,N_14364);
nor U18488 (N_18488,N_14808,N_14792);
or U18489 (N_18489,N_10201,N_11074);
nor U18490 (N_18490,N_11935,N_11589);
nand U18491 (N_18491,N_10435,N_11198);
xnor U18492 (N_18492,N_11632,N_10380);
nand U18493 (N_18493,N_13555,N_12858);
nor U18494 (N_18494,N_12049,N_10717);
nand U18495 (N_18495,N_11540,N_11928);
or U18496 (N_18496,N_10516,N_10974);
nor U18497 (N_18497,N_10758,N_10383);
xnor U18498 (N_18498,N_13703,N_10272);
or U18499 (N_18499,N_14268,N_10788);
nor U18500 (N_18500,N_14782,N_14999);
or U18501 (N_18501,N_14401,N_14728);
xnor U18502 (N_18502,N_12830,N_12069);
and U18503 (N_18503,N_11080,N_10493);
or U18504 (N_18504,N_14097,N_11239);
or U18505 (N_18505,N_10808,N_13642);
xor U18506 (N_18506,N_10436,N_14809);
or U18507 (N_18507,N_13898,N_10246);
or U18508 (N_18508,N_12836,N_14726);
and U18509 (N_18509,N_14722,N_14250);
or U18510 (N_18510,N_10727,N_14057);
or U18511 (N_18511,N_10544,N_10326);
nor U18512 (N_18512,N_13238,N_14176);
nand U18513 (N_18513,N_10262,N_10728);
nor U18514 (N_18514,N_11596,N_13434);
nor U18515 (N_18515,N_11580,N_11689);
xnor U18516 (N_18516,N_10545,N_13078);
xor U18517 (N_18517,N_11931,N_14248);
or U18518 (N_18518,N_12984,N_12637);
nand U18519 (N_18519,N_12442,N_10650);
nor U18520 (N_18520,N_12392,N_14858);
and U18521 (N_18521,N_10514,N_12673);
or U18522 (N_18522,N_13333,N_12095);
nor U18523 (N_18523,N_13815,N_14652);
nor U18524 (N_18524,N_14067,N_14781);
and U18525 (N_18525,N_10866,N_14005);
or U18526 (N_18526,N_12452,N_12954);
nor U18527 (N_18527,N_13526,N_12374);
and U18528 (N_18528,N_11448,N_14200);
nor U18529 (N_18529,N_14322,N_13907);
nand U18530 (N_18530,N_14794,N_12269);
nor U18531 (N_18531,N_14220,N_10582);
or U18532 (N_18532,N_11064,N_12441);
nor U18533 (N_18533,N_11359,N_13963);
or U18534 (N_18534,N_14814,N_11021);
nand U18535 (N_18535,N_12874,N_10522);
and U18536 (N_18536,N_11316,N_14940);
or U18537 (N_18537,N_11076,N_10528);
xor U18538 (N_18538,N_12542,N_10383);
nand U18539 (N_18539,N_10283,N_10089);
and U18540 (N_18540,N_14117,N_10981);
nor U18541 (N_18541,N_13304,N_12646);
nor U18542 (N_18542,N_12816,N_12840);
xor U18543 (N_18543,N_14716,N_10176);
nor U18544 (N_18544,N_14299,N_12324);
nor U18545 (N_18545,N_11325,N_13409);
or U18546 (N_18546,N_14454,N_13520);
or U18547 (N_18547,N_12845,N_13760);
or U18548 (N_18548,N_12785,N_12265);
xnor U18549 (N_18549,N_13552,N_10289);
nor U18550 (N_18550,N_11427,N_13995);
and U18551 (N_18551,N_12201,N_14133);
nand U18552 (N_18552,N_10281,N_13226);
nand U18553 (N_18553,N_13138,N_14841);
or U18554 (N_18554,N_14261,N_11467);
and U18555 (N_18555,N_14567,N_10276);
or U18556 (N_18556,N_11737,N_11566);
and U18557 (N_18557,N_14437,N_10532);
or U18558 (N_18558,N_11342,N_11857);
nand U18559 (N_18559,N_12432,N_12046);
nor U18560 (N_18560,N_10957,N_13875);
or U18561 (N_18561,N_10104,N_13999);
and U18562 (N_18562,N_11985,N_12044);
and U18563 (N_18563,N_12744,N_13332);
or U18564 (N_18564,N_11750,N_14593);
xnor U18565 (N_18565,N_11392,N_11606);
and U18566 (N_18566,N_14006,N_11077);
nand U18567 (N_18567,N_14662,N_12655);
and U18568 (N_18568,N_14091,N_12361);
or U18569 (N_18569,N_10442,N_14559);
nand U18570 (N_18570,N_11785,N_12614);
nand U18571 (N_18571,N_13082,N_13429);
and U18572 (N_18572,N_10647,N_13900);
nor U18573 (N_18573,N_12789,N_10632);
nor U18574 (N_18574,N_11048,N_10367);
or U18575 (N_18575,N_10875,N_10714);
or U18576 (N_18576,N_12443,N_14828);
nor U18577 (N_18577,N_13102,N_14699);
nor U18578 (N_18578,N_12481,N_11257);
xor U18579 (N_18579,N_11750,N_12053);
and U18580 (N_18580,N_11185,N_11918);
and U18581 (N_18581,N_10902,N_11381);
nand U18582 (N_18582,N_11960,N_10516);
nand U18583 (N_18583,N_13866,N_11053);
nand U18584 (N_18584,N_14250,N_14831);
or U18585 (N_18585,N_14822,N_11644);
nor U18586 (N_18586,N_10884,N_10178);
or U18587 (N_18587,N_12284,N_14900);
nor U18588 (N_18588,N_12971,N_13750);
and U18589 (N_18589,N_11292,N_13827);
xnor U18590 (N_18590,N_12329,N_12904);
nor U18591 (N_18591,N_13505,N_11607);
nand U18592 (N_18592,N_14641,N_14367);
or U18593 (N_18593,N_11887,N_14966);
or U18594 (N_18594,N_12123,N_13041);
and U18595 (N_18595,N_13936,N_12578);
or U18596 (N_18596,N_12214,N_13922);
or U18597 (N_18597,N_12287,N_10292);
nor U18598 (N_18598,N_13185,N_14452);
or U18599 (N_18599,N_12954,N_12152);
or U18600 (N_18600,N_10508,N_11818);
and U18601 (N_18601,N_14621,N_14372);
and U18602 (N_18602,N_10782,N_13721);
nor U18603 (N_18603,N_12804,N_10041);
and U18604 (N_18604,N_12730,N_11064);
and U18605 (N_18605,N_13948,N_11562);
and U18606 (N_18606,N_11030,N_14160);
and U18607 (N_18607,N_11068,N_11733);
or U18608 (N_18608,N_10657,N_13642);
nand U18609 (N_18609,N_11983,N_10291);
and U18610 (N_18610,N_13773,N_13281);
or U18611 (N_18611,N_12743,N_10087);
and U18612 (N_18612,N_13621,N_10741);
xor U18613 (N_18613,N_12481,N_13305);
nand U18614 (N_18614,N_11354,N_14492);
or U18615 (N_18615,N_10911,N_13251);
xor U18616 (N_18616,N_12071,N_14345);
nand U18617 (N_18617,N_14305,N_10188);
and U18618 (N_18618,N_12093,N_14060);
xor U18619 (N_18619,N_11607,N_14136);
and U18620 (N_18620,N_11826,N_13133);
nand U18621 (N_18621,N_12194,N_13451);
nand U18622 (N_18622,N_13862,N_10246);
and U18623 (N_18623,N_12935,N_10692);
or U18624 (N_18624,N_13339,N_12680);
and U18625 (N_18625,N_10193,N_14685);
nand U18626 (N_18626,N_14046,N_14291);
nand U18627 (N_18627,N_11974,N_10703);
nor U18628 (N_18628,N_10587,N_12954);
nand U18629 (N_18629,N_12791,N_13024);
or U18630 (N_18630,N_10766,N_14193);
and U18631 (N_18631,N_13096,N_11316);
nand U18632 (N_18632,N_14288,N_10231);
nor U18633 (N_18633,N_11920,N_10590);
nor U18634 (N_18634,N_11593,N_12230);
nand U18635 (N_18635,N_14554,N_14050);
and U18636 (N_18636,N_12532,N_14234);
nand U18637 (N_18637,N_11414,N_11931);
and U18638 (N_18638,N_11412,N_10403);
or U18639 (N_18639,N_13271,N_13305);
nand U18640 (N_18640,N_11034,N_14107);
and U18641 (N_18641,N_12930,N_13807);
or U18642 (N_18642,N_14381,N_12217);
nor U18643 (N_18643,N_11879,N_13006);
nand U18644 (N_18644,N_11201,N_10270);
nand U18645 (N_18645,N_14226,N_12731);
nor U18646 (N_18646,N_11521,N_12725);
xnor U18647 (N_18647,N_11365,N_10465);
xnor U18648 (N_18648,N_12435,N_10890);
or U18649 (N_18649,N_10520,N_10290);
and U18650 (N_18650,N_14141,N_13917);
nand U18651 (N_18651,N_10234,N_12335);
and U18652 (N_18652,N_11372,N_10182);
xnor U18653 (N_18653,N_14137,N_11432);
nand U18654 (N_18654,N_10125,N_10286);
and U18655 (N_18655,N_10673,N_13946);
and U18656 (N_18656,N_12513,N_11547);
nor U18657 (N_18657,N_10522,N_14646);
xor U18658 (N_18658,N_12458,N_12777);
nand U18659 (N_18659,N_12295,N_10002);
or U18660 (N_18660,N_13919,N_13057);
nor U18661 (N_18661,N_10324,N_10863);
or U18662 (N_18662,N_12800,N_12824);
or U18663 (N_18663,N_11575,N_13363);
or U18664 (N_18664,N_13415,N_11016);
nor U18665 (N_18665,N_12442,N_13864);
nor U18666 (N_18666,N_10529,N_12733);
and U18667 (N_18667,N_12868,N_12103);
or U18668 (N_18668,N_12045,N_10793);
or U18669 (N_18669,N_10779,N_10393);
nor U18670 (N_18670,N_11113,N_11598);
and U18671 (N_18671,N_11750,N_11117);
nand U18672 (N_18672,N_11542,N_12454);
xnor U18673 (N_18673,N_10788,N_14560);
nand U18674 (N_18674,N_12864,N_12823);
or U18675 (N_18675,N_12026,N_12815);
and U18676 (N_18676,N_11864,N_13003);
nand U18677 (N_18677,N_12499,N_13329);
or U18678 (N_18678,N_10185,N_10196);
nand U18679 (N_18679,N_12245,N_10128);
nor U18680 (N_18680,N_11593,N_14497);
or U18681 (N_18681,N_11729,N_13383);
xor U18682 (N_18682,N_13306,N_10390);
or U18683 (N_18683,N_14937,N_14136);
nor U18684 (N_18684,N_11878,N_12225);
nand U18685 (N_18685,N_12794,N_11285);
nor U18686 (N_18686,N_11440,N_14074);
nor U18687 (N_18687,N_14907,N_11262);
xnor U18688 (N_18688,N_12768,N_14309);
nand U18689 (N_18689,N_10800,N_11497);
nand U18690 (N_18690,N_13094,N_14518);
and U18691 (N_18691,N_13133,N_11721);
nor U18692 (N_18692,N_13751,N_14092);
nor U18693 (N_18693,N_11614,N_14268);
and U18694 (N_18694,N_10232,N_14998);
nor U18695 (N_18695,N_14955,N_13616);
and U18696 (N_18696,N_13019,N_11064);
nor U18697 (N_18697,N_13146,N_11935);
nor U18698 (N_18698,N_12590,N_11484);
and U18699 (N_18699,N_14653,N_13181);
and U18700 (N_18700,N_14511,N_13908);
and U18701 (N_18701,N_12131,N_13585);
nand U18702 (N_18702,N_14495,N_13256);
nor U18703 (N_18703,N_11512,N_13201);
nand U18704 (N_18704,N_12784,N_14716);
xnor U18705 (N_18705,N_12403,N_11225);
nand U18706 (N_18706,N_12816,N_13864);
nor U18707 (N_18707,N_11801,N_12080);
xnor U18708 (N_18708,N_11895,N_13020);
nor U18709 (N_18709,N_14790,N_10815);
nand U18710 (N_18710,N_13994,N_10152);
or U18711 (N_18711,N_12508,N_12841);
or U18712 (N_18712,N_14116,N_12049);
and U18713 (N_18713,N_12686,N_12880);
and U18714 (N_18714,N_11292,N_10207);
or U18715 (N_18715,N_13393,N_12628);
nand U18716 (N_18716,N_12981,N_14706);
nor U18717 (N_18717,N_11767,N_10766);
nand U18718 (N_18718,N_10939,N_14228);
nand U18719 (N_18719,N_12604,N_13379);
xnor U18720 (N_18720,N_13604,N_10304);
nor U18721 (N_18721,N_11360,N_13688);
nand U18722 (N_18722,N_12556,N_12325);
xnor U18723 (N_18723,N_12350,N_11647);
and U18724 (N_18724,N_10926,N_14920);
nand U18725 (N_18725,N_12118,N_13263);
and U18726 (N_18726,N_13940,N_12598);
or U18727 (N_18727,N_14314,N_10342);
nor U18728 (N_18728,N_11487,N_12067);
or U18729 (N_18729,N_12775,N_14465);
and U18730 (N_18730,N_14361,N_12898);
nand U18731 (N_18731,N_14281,N_11714);
nor U18732 (N_18732,N_12813,N_10063);
nor U18733 (N_18733,N_13416,N_10312);
and U18734 (N_18734,N_12592,N_11526);
or U18735 (N_18735,N_10694,N_13063);
nor U18736 (N_18736,N_13681,N_14532);
nand U18737 (N_18737,N_13139,N_14656);
or U18738 (N_18738,N_14022,N_11232);
nand U18739 (N_18739,N_12119,N_10176);
and U18740 (N_18740,N_12578,N_13528);
nor U18741 (N_18741,N_11281,N_12669);
nand U18742 (N_18742,N_13453,N_12331);
or U18743 (N_18743,N_10446,N_12336);
and U18744 (N_18744,N_13993,N_14894);
or U18745 (N_18745,N_13684,N_12309);
nor U18746 (N_18746,N_10962,N_14952);
nor U18747 (N_18747,N_11407,N_13304);
nand U18748 (N_18748,N_11665,N_10953);
nand U18749 (N_18749,N_11627,N_14636);
xnor U18750 (N_18750,N_13623,N_11818);
or U18751 (N_18751,N_10537,N_10827);
or U18752 (N_18752,N_13176,N_13511);
nand U18753 (N_18753,N_13796,N_10818);
and U18754 (N_18754,N_13302,N_11660);
nor U18755 (N_18755,N_13331,N_11395);
nor U18756 (N_18756,N_12478,N_13060);
or U18757 (N_18757,N_12193,N_13468);
nand U18758 (N_18758,N_11409,N_14847);
nor U18759 (N_18759,N_10963,N_10928);
and U18760 (N_18760,N_14909,N_11412);
or U18761 (N_18761,N_12272,N_12640);
or U18762 (N_18762,N_13720,N_11110);
and U18763 (N_18763,N_13149,N_11591);
nor U18764 (N_18764,N_11610,N_13341);
xor U18765 (N_18765,N_10279,N_14015);
or U18766 (N_18766,N_12326,N_10848);
xnor U18767 (N_18767,N_13787,N_13123);
xnor U18768 (N_18768,N_13936,N_11586);
and U18769 (N_18769,N_11642,N_11929);
or U18770 (N_18770,N_11695,N_12313);
and U18771 (N_18771,N_10335,N_13105);
and U18772 (N_18772,N_14523,N_13764);
nor U18773 (N_18773,N_12753,N_10080);
and U18774 (N_18774,N_13199,N_12618);
and U18775 (N_18775,N_10944,N_13380);
or U18776 (N_18776,N_14145,N_13610);
xor U18777 (N_18777,N_13142,N_12139);
nor U18778 (N_18778,N_13289,N_13547);
or U18779 (N_18779,N_10052,N_12781);
nor U18780 (N_18780,N_12272,N_10638);
and U18781 (N_18781,N_13556,N_12084);
nand U18782 (N_18782,N_13679,N_11125);
nor U18783 (N_18783,N_10334,N_10519);
and U18784 (N_18784,N_12838,N_10270);
or U18785 (N_18785,N_10173,N_12943);
or U18786 (N_18786,N_11954,N_12399);
or U18787 (N_18787,N_14259,N_14452);
nor U18788 (N_18788,N_11766,N_11035);
nand U18789 (N_18789,N_10009,N_14123);
nor U18790 (N_18790,N_12187,N_14278);
and U18791 (N_18791,N_14569,N_12517);
nor U18792 (N_18792,N_10272,N_12815);
or U18793 (N_18793,N_14495,N_10629);
and U18794 (N_18794,N_11204,N_12601);
nand U18795 (N_18795,N_14499,N_11587);
and U18796 (N_18796,N_14728,N_12368);
or U18797 (N_18797,N_10910,N_13615);
nand U18798 (N_18798,N_12549,N_10369);
nor U18799 (N_18799,N_10733,N_12384);
nand U18800 (N_18800,N_14935,N_11069);
nand U18801 (N_18801,N_12806,N_12101);
and U18802 (N_18802,N_12526,N_13412);
nand U18803 (N_18803,N_10915,N_14328);
nor U18804 (N_18804,N_10495,N_14096);
xor U18805 (N_18805,N_11666,N_12125);
nand U18806 (N_18806,N_10237,N_11434);
and U18807 (N_18807,N_12733,N_13399);
xnor U18808 (N_18808,N_11837,N_14023);
or U18809 (N_18809,N_10319,N_14009);
or U18810 (N_18810,N_11100,N_13251);
nor U18811 (N_18811,N_11454,N_10378);
or U18812 (N_18812,N_14498,N_14647);
xor U18813 (N_18813,N_11193,N_14694);
and U18814 (N_18814,N_11625,N_13305);
nand U18815 (N_18815,N_13029,N_13274);
nor U18816 (N_18816,N_13777,N_12888);
nand U18817 (N_18817,N_10975,N_13612);
xor U18818 (N_18818,N_14700,N_10607);
nand U18819 (N_18819,N_10962,N_14462);
or U18820 (N_18820,N_13538,N_11253);
and U18821 (N_18821,N_13468,N_13266);
xnor U18822 (N_18822,N_11482,N_14690);
or U18823 (N_18823,N_12673,N_12293);
nand U18824 (N_18824,N_14183,N_11450);
nor U18825 (N_18825,N_14402,N_14112);
nor U18826 (N_18826,N_10471,N_10067);
nor U18827 (N_18827,N_12400,N_10319);
or U18828 (N_18828,N_11070,N_10774);
xnor U18829 (N_18829,N_13931,N_13905);
nand U18830 (N_18830,N_12514,N_12405);
and U18831 (N_18831,N_12414,N_10766);
and U18832 (N_18832,N_11550,N_10244);
xnor U18833 (N_18833,N_12437,N_12201);
and U18834 (N_18834,N_10065,N_10809);
nand U18835 (N_18835,N_11044,N_11192);
nand U18836 (N_18836,N_12888,N_12628);
nor U18837 (N_18837,N_11881,N_12271);
and U18838 (N_18838,N_12353,N_10183);
nand U18839 (N_18839,N_10073,N_12602);
nor U18840 (N_18840,N_12416,N_12550);
nor U18841 (N_18841,N_10895,N_13354);
or U18842 (N_18842,N_10113,N_13882);
nor U18843 (N_18843,N_12248,N_10657);
or U18844 (N_18844,N_14046,N_12489);
and U18845 (N_18845,N_13582,N_14981);
nand U18846 (N_18846,N_11667,N_10828);
nor U18847 (N_18847,N_13634,N_14568);
nor U18848 (N_18848,N_12674,N_12696);
xor U18849 (N_18849,N_14374,N_13315);
or U18850 (N_18850,N_13779,N_14423);
nor U18851 (N_18851,N_11339,N_14102);
nor U18852 (N_18852,N_14740,N_11294);
nor U18853 (N_18853,N_11873,N_10124);
nand U18854 (N_18854,N_10297,N_11451);
or U18855 (N_18855,N_11981,N_13779);
nor U18856 (N_18856,N_10947,N_13645);
nor U18857 (N_18857,N_14549,N_13883);
nand U18858 (N_18858,N_12470,N_11371);
and U18859 (N_18859,N_10372,N_12856);
nand U18860 (N_18860,N_14587,N_12707);
nor U18861 (N_18861,N_13847,N_14886);
and U18862 (N_18862,N_10740,N_12331);
and U18863 (N_18863,N_13141,N_13943);
nand U18864 (N_18864,N_11916,N_14902);
or U18865 (N_18865,N_12179,N_12365);
nor U18866 (N_18866,N_14618,N_11278);
or U18867 (N_18867,N_11194,N_13325);
or U18868 (N_18868,N_10620,N_13664);
nor U18869 (N_18869,N_13416,N_12796);
nand U18870 (N_18870,N_10239,N_13940);
and U18871 (N_18871,N_10007,N_11016);
nor U18872 (N_18872,N_10035,N_13379);
and U18873 (N_18873,N_11414,N_14039);
or U18874 (N_18874,N_11463,N_11475);
nand U18875 (N_18875,N_13783,N_14616);
nor U18876 (N_18876,N_14523,N_10387);
nand U18877 (N_18877,N_14971,N_10632);
and U18878 (N_18878,N_13590,N_12593);
nor U18879 (N_18879,N_13455,N_14014);
nand U18880 (N_18880,N_10166,N_12803);
nand U18881 (N_18881,N_13767,N_14767);
nand U18882 (N_18882,N_10356,N_14973);
nor U18883 (N_18883,N_14668,N_13894);
and U18884 (N_18884,N_11334,N_10800);
or U18885 (N_18885,N_13818,N_12549);
and U18886 (N_18886,N_11068,N_13490);
and U18887 (N_18887,N_11803,N_10274);
nand U18888 (N_18888,N_11315,N_13466);
xor U18889 (N_18889,N_12410,N_14704);
or U18890 (N_18890,N_12465,N_14537);
and U18891 (N_18891,N_11013,N_11209);
nor U18892 (N_18892,N_12370,N_13266);
or U18893 (N_18893,N_11068,N_11786);
nand U18894 (N_18894,N_10304,N_11971);
nand U18895 (N_18895,N_14970,N_10958);
nor U18896 (N_18896,N_14762,N_11405);
nor U18897 (N_18897,N_13772,N_14901);
nor U18898 (N_18898,N_12747,N_12404);
and U18899 (N_18899,N_11927,N_10368);
and U18900 (N_18900,N_13193,N_10015);
nand U18901 (N_18901,N_13611,N_13078);
nor U18902 (N_18902,N_12674,N_10046);
xnor U18903 (N_18903,N_13647,N_11341);
and U18904 (N_18904,N_14047,N_13194);
and U18905 (N_18905,N_12092,N_10051);
nand U18906 (N_18906,N_12605,N_10795);
nand U18907 (N_18907,N_14702,N_14841);
nor U18908 (N_18908,N_11632,N_12651);
nor U18909 (N_18909,N_14527,N_12339);
nand U18910 (N_18910,N_10416,N_12472);
nor U18911 (N_18911,N_10581,N_12519);
and U18912 (N_18912,N_10980,N_14585);
nor U18913 (N_18913,N_13841,N_10079);
nor U18914 (N_18914,N_12648,N_14603);
and U18915 (N_18915,N_12578,N_10179);
nand U18916 (N_18916,N_12791,N_13834);
nor U18917 (N_18917,N_13079,N_13457);
or U18918 (N_18918,N_14525,N_10260);
nor U18919 (N_18919,N_13002,N_10153);
nand U18920 (N_18920,N_14393,N_12321);
and U18921 (N_18921,N_10552,N_12546);
and U18922 (N_18922,N_14480,N_12878);
or U18923 (N_18923,N_10356,N_10656);
and U18924 (N_18924,N_11672,N_11030);
xnor U18925 (N_18925,N_10155,N_12598);
nand U18926 (N_18926,N_11650,N_13726);
nor U18927 (N_18927,N_13249,N_12007);
xor U18928 (N_18928,N_12999,N_11221);
nand U18929 (N_18929,N_10849,N_11519);
xnor U18930 (N_18930,N_13377,N_10646);
or U18931 (N_18931,N_10051,N_13111);
and U18932 (N_18932,N_10328,N_13141);
nor U18933 (N_18933,N_12566,N_11065);
and U18934 (N_18934,N_10130,N_12336);
nand U18935 (N_18935,N_12422,N_12335);
and U18936 (N_18936,N_10982,N_11722);
nor U18937 (N_18937,N_10729,N_11733);
and U18938 (N_18938,N_14403,N_14757);
or U18939 (N_18939,N_12056,N_11836);
or U18940 (N_18940,N_13040,N_13280);
or U18941 (N_18941,N_13277,N_10982);
or U18942 (N_18942,N_12615,N_14178);
nand U18943 (N_18943,N_13766,N_11090);
nand U18944 (N_18944,N_13258,N_12888);
nor U18945 (N_18945,N_13663,N_12497);
and U18946 (N_18946,N_12866,N_14371);
and U18947 (N_18947,N_11312,N_12572);
nand U18948 (N_18948,N_10471,N_11738);
and U18949 (N_18949,N_11998,N_11009);
and U18950 (N_18950,N_10210,N_10538);
and U18951 (N_18951,N_14440,N_12939);
and U18952 (N_18952,N_12819,N_10368);
or U18953 (N_18953,N_10031,N_10809);
nor U18954 (N_18954,N_14625,N_10453);
nand U18955 (N_18955,N_14810,N_14385);
or U18956 (N_18956,N_12886,N_14710);
xnor U18957 (N_18957,N_14063,N_13645);
nor U18958 (N_18958,N_14977,N_12568);
or U18959 (N_18959,N_12890,N_14248);
nor U18960 (N_18960,N_10288,N_11919);
or U18961 (N_18961,N_12498,N_13954);
and U18962 (N_18962,N_10808,N_10538);
and U18963 (N_18963,N_14160,N_10868);
or U18964 (N_18964,N_10918,N_14629);
xnor U18965 (N_18965,N_11152,N_10018);
nand U18966 (N_18966,N_13816,N_10814);
nand U18967 (N_18967,N_11399,N_13440);
or U18968 (N_18968,N_12374,N_13805);
nand U18969 (N_18969,N_12864,N_12416);
or U18970 (N_18970,N_12308,N_14063);
xor U18971 (N_18971,N_12361,N_13766);
and U18972 (N_18972,N_11574,N_11678);
xnor U18973 (N_18973,N_12351,N_12507);
or U18974 (N_18974,N_10306,N_12921);
nand U18975 (N_18975,N_11923,N_11273);
nor U18976 (N_18976,N_13527,N_13555);
nand U18977 (N_18977,N_14957,N_13315);
nand U18978 (N_18978,N_12509,N_10357);
or U18979 (N_18979,N_13492,N_12530);
xnor U18980 (N_18980,N_10251,N_11742);
or U18981 (N_18981,N_14441,N_13844);
and U18982 (N_18982,N_10788,N_10511);
nand U18983 (N_18983,N_14468,N_11147);
xnor U18984 (N_18984,N_13017,N_14254);
or U18985 (N_18985,N_11078,N_14914);
and U18986 (N_18986,N_14284,N_10996);
and U18987 (N_18987,N_13463,N_10716);
nor U18988 (N_18988,N_11115,N_14225);
xnor U18989 (N_18989,N_11141,N_10323);
nand U18990 (N_18990,N_14992,N_13533);
and U18991 (N_18991,N_11166,N_12277);
and U18992 (N_18992,N_13957,N_14819);
or U18993 (N_18993,N_12348,N_13772);
and U18994 (N_18994,N_12730,N_12213);
or U18995 (N_18995,N_14580,N_12819);
and U18996 (N_18996,N_11166,N_10215);
or U18997 (N_18997,N_11188,N_11871);
nand U18998 (N_18998,N_13757,N_11673);
nand U18999 (N_18999,N_14904,N_12262);
nand U19000 (N_19000,N_14184,N_13893);
nor U19001 (N_19001,N_12608,N_11715);
nand U19002 (N_19002,N_12309,N_12850);
nor U19003 (N_19003,N_10113,N_10450);
nand U19004 (N_19004,N_13755,N_14896);
or U19005 (N_19005,N_13088,N_13401);
or U19006 (N_19006,N_12737,N_11113);
nand U19007 (N_19007,N_11858,N_14296);
nand U19008 (N_19008,N_12455,N_14583);
and U19009 (N_19009,N_12874,N_12675);
nand U19010 (N_19010,N_14372,N_11344);
and U19011 (N_19011,N_13569,N_14833);
and U19012 (N_19012,N_14477,N_14753);
and U19013 (N_19013,N_10851,N_11002);
or U19014 (N_19014,N_14563,N_11049);
nor U19015 (N_19015,N_14850,N_14705);
xor U19016 (N_19016,N_14385,N_11339);
or U19017 (N_19017,N_12893,N_13155);
nor U19018 (N_19018,N_13968,N_14764);
nor U19019 (N_19019,N_14076,N_14283);
or U19020 (N_19020,N_13747,N_10024);
nand U19021 (N_19021,N_12135,N_13857);
and U19022 (N_19022,N_12522,N_10330);
and U19023 (N_19023,N_14487,N_10412);
or U19024 (N_19024,N_12974,N_13115);
nand U19025 (N_19025,N_14114,N_10890);
xnor U19026 (N_19026,N_13716,N_14861);
and U19027 (N_19027,N_13067,N_13411);
nand U19028 (N_19028,N_10431,N_14965);
nand U19029 (N_19029,N_13041,N_13676);
and U19030 (N_19030,N_10192,N_11613);
nor U19031 (N_19031,N_10318,N_11423);
and U19032 (N_19032,N_11173,N_13267);
xor U19033 (N_19033,N_14578,N_14934);
nand U19034 (N_19034,N_13734,N_12232);
nand U19035 (N_19035,N_14519,N_11773);
or U19036 (N_19036,N_10209,N_12990);
or U19037 (N_19037,N_10039,N_12499);
nor U19038 (N_19038,N_10188,N_11640);
or U19039 (N_19039,N_11639,N_13599);
and U19040 (N_19040,N_10836,N_13392);
and U19041 (N_19041,N_13316,N_13378);
or U19042 (N_19042,N_10634,N_14484);
xor U19043 (N_19043,N_13414,N_11637);
xnor U19044 (N_19044,N_14391,N_11395);
and U19045 (N_19045,N_10301,N_12924);
or U19046 (N_19046,N_10557,N_10247);
and U19047 (N_19047,N_12609,N_13789);
nor U19048 (N_19048,N_10511,N_12251);
nor U19049 (N_19049,N_10368,N_14901);
nand U19050 (N_19050,N_14149,N_13897);
and U19051 (N_19051,N_12205,N_12281);
nand U19052 (N_19052,N_14850,N_14838);
or U19053 (N_19053,N_11337,N_11692);
xor U19054 (N_19054,N_13199,N_11424);
xor U19055 (N_19055,N_13753,N_12438);
and U19056 (N_19056,N_11454,N_14705);
nor U19057 (N_19057,N_10672,N_11105);
xor U19058 (N_19058,N_10933,N_10201);
and U19059 (N_19059,N_10956,N_10307);
and U19060 (N_19060,N_10567,N_12781);
xnor U19061 (N_19061,N_11225,N_13286);
xor U19062 (N_19062,N_11861,N_11966);
xnor U19063 (N_19063,N_10766,N_12465);
and U19064 (N_19064,N_13933,N_14565);
nor U19065 (N_19065,N_12031,N_11656);
nand U19066 (N_19066,N_14126,N_14170);
nor U19067 (N_19067,N_10608,N_12373);
or U19068 (N_19068,N_12786,N_10173);
nor U19069 (N_19069,N_12713,N_11648);
and U19070 (N_19070,N_11310,N_11238);
or U19071 (N_19071,N_12376,N_10310);
or U19072 (N_19072,N_13572,N_13537);
or U19073 (N_19073,N_10196,N_13193);
nand U19074 (N_19074,N_10263,N_13823);
xnor U19075 (N_19075,N_11329,N_10161);
and U19076 (N_19076,N_13594,N_11367);
and U19077 (N_19077,N_13360,N_10037);
nor U19078 (N_19078,N_13814,N_14571);
and U19079 (N_19079,N_13413,N_11549);
nor U19080 (N_19080,N_10277,N_13173);
nor U19081 (N_19081,N_12754,N_10947);
or U19082 (N_19082,N_11878,N_11682);
nor U19083 (N_19083,N_10800,N_13066);
xnor U19084 (N_19084,N_12534,N_10823);
nand U19085 (N_19085,N_12117,N_11666);
xnor U19086 (N_19086,N_11281,N_12610);
or U19087 (N_19087,N_14893,N_11716);
nand U19088 (N_19088,N_11597,N_14659);
or U19089 (N_19089,N_10759,N_10783);
xor U19090 (N_19090,N_14831,N_10298);
nand U19091 (N_19091,N_13671,N_10998);
nor U19092 (N_19092,N_14064,N_14369);
nand U19093 (N_19093,N_11013,N_11765);
nor U19094 (N_19094,N_11630,N_10628);
nand U19095 (N_19095,N_13170,N_12002);
nor U19096 (N_19096,N_10267,N_13484);
or U19097 (N_19097,N_11700,N_11342);
nor U19098 (N_19098,N_11847,N_12152);
nor U19099 (N_19099,N_14039,N_10500);
nor U19100 (N_19100,N_12381,N_11230);
xnor U19101 (N_19101,N_13563,N_14997);
nand U19102 (N_19102,N_13361,N_14070);
nand U19103 (N_19103,N_11279,N_13826);
xnor U19104 (N_19104,N_12052,N_11403);
nand U19105 (N_19105,N_10543,N_11120);
and U19106 (N_19106,N_10447,N_14830);
or U19107 (N_19107,N_13203,N_14322);
xnor U19108 (N_19108,N_12187,N_10080);
nor U19109 (N_19109,N_13031,N_12369);
or U19110 (N_19110,N_10171,N_12543);
xor U19111 (N_19111,N_10676,N_12124);
or U19112 (N_19112,N_12410,N_13353);
nand U19113 (N_19113,N_10898,N_14472);
xnor U19114 (N_19114,N_13884,N_10273);
or U19115 (N_19115,N_10404,N_12109);
and U19116 (N_19116,N_12408,N_12589);
or U19117 (N_19117,N_14011,N_10797);
nand U19118 (N_19118,N_11459,N_11213);
and U19119 (N_19119,N_12258,N_10579);
and U19120 (N_19120,N_14274,N_14442);
and U19121 (N_19121,N_12779,N_14518);
and U19122 (N_19122,N_11069,N_13341);
nor U19123 (N_19123,N_11259,N_12062);
or U19124 (N_19124,N_10590,N_13006);
and U19125 (N_19125,N_11704,N_10980);
and U19126 (N_19126,N_10765,N_10096);
nor U19127 (N_19127,N_12597,N_14333);
nor U19128 (N_19128,N_13141,N_13581);
nand U19129 (N_19129,N_12209,N_13829);
and U19130 (N_19130,N_11943,N_11617);
nor U19131 (N_19131,N_13296,N_13450);
or U19132 (N_19132,N_14832,N_13267);
xnor U19133 (N_19133,N_11062,N_12529);
and U19134 (N_19134,N_14255,N_12399);
nor U19135 (N_19135,N_11634,N_13194);
and U19136 (N_19136,N_11549,N_14206);
nand U19137 (N_19137,N_14520,N_11197);
nor U19138 (N_19138,N_10788,N_12488);
and U19139 (N_19139,N_12108,N_10969);
xnor U19140 (N_19140,N_13090,N_14474);
nor U19141 (N_19141,N_14055,N_13697);
or U19142 (N_19142,N_11187,N_13805);
or U19143 (N_19143,N_14941,N_13383);
nor U19144 (N_19144,N_14796,N_13452);
nor U19145 (N_19145,N_13505,N_14070);
and U19146 (N_19146,N_13898,N_13545);
nand U19147 (N_19147,N_14896,N_10967);
or U19148 (N_19148,N_13479,N_12843);
xnor U19149 (N_19149,N_12336,N_13495);
nor U19150 (N_19150,N_12229,N_11582);
nor U19151 (N_19151,N_10335,N_14860);
and U19152 (N_19152,N_11128,N_11733);
or U19153 (N_19153,N_11904,N_10263);
xor U19154 (N_19154,N_14677,N_12775);
and U19155 (N_19155,N_14181,N_12833);
nand U19156 (N_19156,N_11528,N_12236);
and U19157 (N_19157,N_13904,N_14009);
or U19158 (N_19158,N_13998,N_13988);
nor U19159 (N_19159,N_13002,N_13226);
or U19160 (N_19160,N_14319,N_10822);
nor U19161 (N_19161,N_11252,N_10524);
and U19162 (N_19162,N_10721,N_11140);
nand U19163 (N_19163,N_14235,N_14983);
nand U19164 (N_19164,N_14075,N_14509);
and U19165 (N_19165,N_14818,N_13016);
and U19166 (N_19166,N_10561,N_10364);
and U19167 (N_19167,N_12424,N_10908);
nand U19168 (N_19168,N_13125,N_10761);
nor U19169 (N_19169,N_13745,N_11679);
or U19170 (N_19170,N_11687,N_11501);
nand U19171 (N_19171,N_12967,N_12455);
nand U19172 (N_19172,N_12828,N_12226);
xnor U19173 (N_19173,N_10094,N_12312);
nand U19174 (N_19174,N_12541,N_13451);
nand U19175 (N_19175,N_12065,N_10367);
nand U19176 (N_19176,N_14667,N_11454);
nor U19177 (N_19177,N_13526,N_13429);
or U19178 (N_19178,N_11727,N_14979);
or U19179 (N_19179,N_10760,N_14266);
or U19180 (N_19180,N_10104,N_10599);
xnor U19181 (N_19181,N_12119,N_13986);
or U19182 (N_19182,N_13544,N_13219);
nand U19183 (N_19183,N_14194,N_10426);
and U19184 (N_19184,N_10868,N_13159);
nor U19185 (N_19185,N_13369,N_10403);
or U19186 (N_19186,N_11114,N_11283);
or U19187 (N_19187,N_14532,N_12329);
nand U19188 (N_19188,N_11429,N_13352);
and U19189 (N_19189,N_14773,N_12371);
nor U19190 (N_19190,N_10563,N_10305);
nand U19191 (N_19191,N_11050,N_14070);
or U19192 (N_19192,N_12007,N_10543);
or U19193 (N_19193,N_13512,N_11570);
or U19194 (N_19194,N_11524,N_13511);
or U19195 (N_19195,N_14549,N_11399);
nand U19196 (N_19196,N_10935,N_14558);
nor U19197 (N_19197,N_14804,N_10125);
nor U19198 (N_19198,N_14810,N_14615);
or U19199 (N_19199,N_14211,N_11508);
nor U19200 (N_19200,N_12831,N_10885);
nand U19201 (N_19201,N_14532,N_13645);
and U19202 (N_19202,N_11485,N_14120);
nor U19203 (N_19203,N_14721,N_10226);
xor U19204 (N_19204,N_14080,N_14631);
nand U19205 (N_19205,N_13557,N_13079);
xnor U19206 (N_19206,N_14013,N_10133);
and U19207 (N_19207,N_11549,N_12007);
or U19208 (N_19208,N_13920,N_10290);
nand U19209 (N_19209,N_11337,N_13709);
nor U19210 (N_19210,N_13568,N_14481);
and U19211 (N_19211,N_11715,N_10988);
nand U19212 (N_19212,N_11836,N_14062);
nand U19213 (N_19213,N_13795,N_11529);
and U19214 (N_19214,N_14357,N_13058);
or U19215 (N_19215,N_10730,N_12760);
or U19216 (N_19216,N_12171,N_13184);
nor U19217 (N_19217,N_11516,N_11490);
or U19218 (N_19218,N_13431,N_11586);
and U19219 (N_19219,N_10726,N_13860);
nand U19220 (N_19220,N_12247,N_13783);
nor U19221 (N_19221,N_11538,N_13642);
or U19222 (N_19222,N_10923,N_13223);
nand U19223 (N_19223,N_14493,N_11446);
nand U19224 (N_19224,N_14708,N_10423);
nor U19225 (N_19225,N_13955,N_11751);
nand U19226 (N_19226,N_11313,N_12165);
nor U19227 (N_19227,N_13995,N_11023);
nor U19228 (N_19228,N_13922,N_11756);
nor U19229 (N_19229,N_13650,N_11318);
and U19230 (N_19230,N_13576,N_12507);
or U19231 (N_19231,N_13765,N_13399);
or U19232 (N_19232,N_11381,N_11387);
nor U19233 (N_19233,N_12835,N_13614);
and U19234 (N_19234,N_10840,N_10844);
nor U19235 (N_19235,N_13867,N_12073);
or U19236 (N_19236,N_13463,N_14865);
nor U19237 (N_19237,N_12669,N_12384);
nor U19238 (N_19238,N_14888,N_11950);
or U19239 (N_19239,N_13956,N_12255);
or U19240 (N_19240,N_14661,N_11608);
and U19241 (N_19241,N_13699,N_14473);
and U19242 (N_19242,N_10858,N_11078);
nor U19243 (N_19243,N_11955,N_11276);
or U19244 (N_19244,N_10667,N_14106);
xnor U19245 (N_19245,N_12338,N_14524);
nor U19246 (N_19246,N_13714,N_10894);
or U19247 (N_19247,N_12518,N_14839);
nor U19248 (N_19248,N_14770,N_14152);
and U19249 (N_19249,N_10044,N_14216);
nand U19250 (N_19250,N_10450,N_14735);
nand U19251 (N_19251,N_11691,N_14446);
or U19252 (N_19252,N_12169,N_14349);
or U19253 (N_19253,N_10375,N_11246);
and U19254 (N_19254,N_11735,N_12722);
nor U19255 (N_19255,N_13550,N_12418);
nand U19256 (N_19256,N_12952,N_14512);
nor U19257 (N_19257,N_10591,N_12668);
nand U19258 (N_19258,N_12634,N_10261);
nor U19259 (N_19259,N_14984,N_13313);
xnor U19260 (N_19260,N_14700,N_14516);
and U19261 (N_19261,N_13469,N_10505);
or U19262 (N_19262,N_11240,N_11056);
and U19263 (N_19263,N_12846,N_14654);
nand U19264 (N_19264,N_14709,N_11055);
nor U19265 (N_19265,N_11904,N_10806);
nor U19266 (N_19266,N_10757,N_12386);
nor U19267 (N_19267,N_14701,N_10361);
nor U19268 (N_19268,N_10847,N_14459);
and U19269 (N_19269,N_14015,N_11439);
nor U19270 (N_19270,N_11483,N_14254);
nor U19271 (N_19271,N_10518,N_11003);
xnor U19272 (N_19272,N_10025,N_13618);
nand U19273 (N_19273,N_10382,N_13934);
and U19274 (N_19274,N_12485,N_10380);
nor U19275 (N_19275,N_13900,N_11197);
or U19276 (N_19276,N_14054,N_10145);
or U19277 (N_19277,N_10933,N_14608);
xor U19278 (N_19278,N_11805,N_10775);
and U19279 (N_19279,N_14971,N_14003);
xnor U19280 (N_19280,N_11539,N_12990);
nand U19281 (N_19281,N_12837,N_12332);
nor U19282 (N_19282,N_10571,N_10606);
nor U19283 (N_19283,N_13871,N_10804);
and U19284 (N_19284,N_11348,N_12006);
nor U19285 (N_19285,N_14829,N_11655);
or U19286 (N_19286,N_12309,N_12716);
and U19287 (N_19287,N_13954,N_13008);
and U19288 (N_19288,N_13014,N_12620);
and U19289 (N_19289,N_13694,N_10071);
or U19290 (N_19290,N_12949,N_11666);
or U19291 (N_19291,N_10752,N_11395);
nor U19292 (N_19292,N_10258,N_12065);
and U19293 (N_19293,N_14456,N_14497);
nand U19294 (N_19294,N_13540,N_13022);
xnor U19295 (N_19295,N_10247,N_11455);
nand U19296 (N_19296,N_14223,N_11997);
or U19297 (N_19297,N_14889,N_12566);
nand U19298 (N_19298,N_12378,N_13615);
nand U19299 (N_19299,N_14638,N_11446);
or U19300 (N_19300,N_10062,N_12112);
or U19301 (N_19301,N_14385,N_10655);
or U19302 (N_19302,N_12083,N_13677);
nand U19303 (N_19303,N_13720,N_11567);
and U19304 (N_19304,N_14436,N_13317);
nand U19305 (N_19305,N_13652,N_14934);
and U19306 (N_19306,N_14022,N_10861);
or U19307 (N_19307,N_12940,N_13884);
or U19308 (N_19308,N_14416,N_14403);
nor U19309 (N_19309,N_14102,N_10574);
and U19310 (N_19310,N_11302,N_11361);
xnor U19311 (N_19311,N_12167,N_14040);
nor U19312 (N_19312,N_14207,N_11936);
nand U19313 (N_19313,N_12655,N_13000);
nand U19314 (N_19314,N_12153,N_12960);
nor U19315 (N_19315,N_13081,N_13662);
or U19316 (N_19316,N_13855,N_10038);
nand U19317 (N_19317,N_10971,N_12561);
nand U19318 (N_19318,N_10573,N_14252);
nor U19319 (N_19319,N_13439,N_14222);
nand U19320 (N_19320,N_11427,N_12978);
and U19321 (N_19321,N_11970,N_14003);
nor U19322 (N_19322,N_10694,N_11912);
nor U19323 (N_19323,N_11332,N_10169);
xor U19324 (N_19324,N_10760,N_12229);
nand U19325 (N_19325,N_14233,N_12972);
nor U19326 (N_19326,N_13442,N_14367);
and U19327 (N_19327,N_11906,N_12172);
nor U19328 (N_19328,N_14030,N_14829);
nor U19329 (N_19329,N_13313,N_10925);
nor U19330 (N_19330,N_13040,N_13153);
and U19331 (N_19331,N_12108,N_12051);
or U19332 (N_19332,N_13340,N_13991);
nor U19333 (N_19333,N_11173,N_11833);
and U19334 (N_19334,N_12368,N_10238);
xor U19335 (N_19335,N_10706,N_10796);
nand U19336 (N_19336,N_10750,N_12527);
or U19337 (N_19337,N_11167,N_11030);
or U19338 (N_19338,N_10771,N_10941);
and U19339 (N_19339,N_12167,N_14058);
and U19340 (N_19340,N_10567,N_14425);
nor U19341 (N_19341,N_11718,N_10317);
nor U19342 (N_19342,N_12347,N_14888);
xnor U19343 (N_19343,N_13270,N_11725);
and U19344 (N_19344,N_10027,N_12514);
or U19345 (N_19345,N_14884,N_14090);
nand U19346 (N_19346,N_13234,N_12856);
nand U19347 (N_19347,N_12617,N_11455);
nor U19348 (N_19348,N_11394,N_13171);
or U19349 (N_19349,N_13156,N_10129);
or U19350 (N_19350,N_10360,N_14007);
nor U19351 (N_19351,N_11431,N_11375);
and U19352 (N_19352,N_11721,N_10443);
nand U19353 (N_19353,N_10464,N_14982);
and U19354 (N_19354,N_12559,N_11906);
and U19355 (N_19355,N_11740,N_12924);
and U19356 (N_19356,N_10057,N_13470);
nor U19357 (N_19357,N_10109,N_12646);
or U19358 (N_19358,N_10646,N_10261);
or U19359 (N_19359,N_13404,N_10684);
or U19360 (N_19360,N_13870,N_10333);
nor U19361 (N_19361,N_10772,N_12973);
nor U19362 (N_19362,N_12343,N_10307);
nor U19363 (N_19363,N_13464,N_14018);
nand U19364 (N_19364,N_11999,N_10099);
or U19365 (N_19365,N_12760,N_13480);
xnor U19366 (N_19366,N_11124,N_11209);
and U19367 (N_19367,N_14784,N_14830);
or U19368 (N_19368,N_13267,N_11288);
nand U19369 (N_19369,N_13888,N_12222);
and U19370 (N_19370,N_14778,N_12258);
or U19371 (N_19371,N_13711,N_10676);
and U19372 (N_19372,N_13189,N_11691);
nand U19373 (N_19373,N_12586,N_10037);
nor U19374 (N_19374,N_13407,N_10444);
or U19375 (N_19375,N_10114,N_10421);
nor U19376 (N_19376,N_10757,N_13487);
or U19377 (N_19377,N_14329,N_11449);
or U19378 (N_19378,N_14662,N_13350);
nor U19379 (N_19379,N_12979,N_13027);
or U19380 (N_19380,N_14184,N_13940);
or U19381 (N_19381,N_13820,N_11332);
nor U19382 (N_19382,N_10026,N_12666);
nand U19383 (N_19383,N_12741,N_14406);
xnor U19384 (N_19384,N_11074,N_10008);
nor U19385 (N_19385,N_12648,N_13531);
nor U19386 (N_19386,N_13796,N_10382);
and U19387 (N_19387,N_10061,N_10976);
nand U19388 (N_19388,N_14401,N_11675);
and U19389 (N_19389,N_14569,N_12566);
nand U19390 (N_19390,N_11369,N_10410);
nand U19391 (N_19391,N_10584,N_11157);
nand U19392 (N_19392,N_11894,N_10195);
xnor U19393 (N_19393,N_10297,N_13003);
or U19394 (N_19394,N_14018,N_13842);
nand U19395 (N_19395,N_14145,N_13772);
and U19396 (N_19396,N_10410,N_11882);
nor U19397 (N_19397,N_12605,N_12440);
nor U19398 (N_19398,N_12115,N_13101);
nor U19399 (N_19399,N_13744,N_14302);
xor U19400 (N_19400,N_10463,N_11322);
xnor U19401 (N_19401,N_11929,N_14012);
or U19402 (N_19402,N_14940,N_11447);
nor U19403 (N_19403,N_13392,N_10230);
xor U19404 (N_19404,N_11476,N_13878);
and U19405 (N_19405,N_10958,N_12760);
and U19406 (N_19406,N_10586,N_14636);
and U19407 (N_19407,N_14272,N_10398);
and U19408 (N_19408,N_11684,N_14808);
nand U19409 (N_19409,N_14590,N_11753);
xnor U19410 (N_19410,N_10998,N_11343);
nor U19411 (N_19411,N_12939,N_13936);
xnor U19412 (N_19412,N_14801,N_13836);
and U19413 (N_19413,N_12960,N_11520);
xor U19414 (N_19414,N_12470,N_14865);
nor U19415 (N_19415,N_10361,N_11964);
nand U19416 (N_19416,N_11256,N_13650);
or U19417 (N_19417,N_11932,N_13838);
or U19418 (N_19418,N_10266,N_11364);
or U19419 (N_19419,N_11720,N_14096);
nand U19420 (N_19420,N_13459,N_11805);
or U19421 (N_19421,N_12267,N_12401);
and U19422 (N_19422,N_14444,N_14440);
xor U19423 (N_19423,N_13688,N_13534);
nand U19424 (N_19424,N_12629,N_14632);
nand U19425 (N_19425,N_12337,N_10869);
xor U19426 (N_19426,N_12868,N_14620);
nand U19427 (N_19427,N_13665,N_14713);
nor U19428 (N_19428,N_12319,N_12276);
nor U19429 (N_19429,N_12268,N_12179);
xnor U19430 (N_19430,N_13177,N_12195);
nand U19431 (N_19431,N_13036,N_10570);
or U19432 (N_19432,N_11502,N_13581);
nand U19433 (N_19433,N_12066,N_12400);
or U19434 (N_19434,N_13123,N_11120);
or U19435 (N_19435,N_11531,N_13963);
xnor U19436 (N_19436,N_14029,N_13148);
and U19437 (N_19437,N_14353,N_14481);
and U19438 (N_19438,N_10319,N_14257);
and U19439 (N_19439,N_14032,N_10463);
and U19440 (N_19440,N_13704,N_14157);
nand U19441 (N_19441,N_10206,N_14016);
and U19442 (N_19442,N_11505,N_13622);
or U19443 (N_19443,N_12901,N_11508);
nand U19444 (N_19444,N_13584,N_14219);
nand U19445 (N_19445,N_10205,N_12454);
and U19446 (N_19446,N_14106,N_12773);
xor U19447 (N_19447,N_12205,N_10525);
or U19448 (N_19448,N_14485,N_11329);
or U19449 (N_19449,N_11372,N_11819);
nand U19450 (N_19450,N_10864,N_14722);
nand U19451 (N_19451,N_11558,N_10894);
nor U19452 (N_19452,N_11750,N_14950);
or U19453 (N_19453,N_12035,N_14281);
nand U19454 (N_19454,N_13616,N_12119);
and U19455 (N_19455,N_14775,N_11308);
nand U19456 (N_19456,N_12393,N_10563);
and U19457 (N_19457,N_10192,N_11936);
and U19458 (N_19458,N_12699,N_14026);
and U19459 (N_19459,N_13118,N_11286);
and U19460 (N_19460,N_12618,N_10289);
and U19461 (N_19461,N_14145,N_14745);
and U19462 (N_19462,N_10642,N_12997);
or U19463 (N_19463,N_10221,N_12143);
and U19464 (N_19464,N_12369,N_12943);
nand U19465 (N_19465,N_11362,N_12553);
nor U19466 (N_19466,N_10479,N_14286);
and U19467 (N_19467,N_10527,N_12062);
and U19468 (N_19468,N_14769,N_11136);
or U19469 (N_19469,N_14942,N_12109);
nand U19470 (N_19470,N_14219,N_14183);
xor U19471 (N_19471,N_14520,N_10590);
nor U19472 (N_19472,N_13863,N_13687);
nand U19473 (N_19473,N_10997,N_11414);
and U19474 (N_19474,N_11449,N_14275);
and U19475 (N_19475,N_13126,N_11802);
and U19476 (N_19476,N_11190,N_10874);
and U19477 (N_19477,N_14089,N_10440);
and U19478 (N_19478,N_11640,N_12708);
and U19479 (N_19479,N_10917,N_13794);
and U19480 (N_19480,N_13444,N_13917);
nor U19481 (N_19481,N_11090,N_12728);
nor U19482 (N_19482,N_10709,N_13200);
nor U19483 (N_19483,N_10109,N_14268);
xnor U19484 (N_19484,N_14949,N_12093);
and U19485 (N_19485,N_13248,N_14292);
or U19486 (N_19486,N_14717,N_12299);
xnor U19487 (N_19487,N_12837,N_13185);
xor U19488 (N_19488,N_10970,N_11680);
xor U19489 (N_19489,N_10720,N_13100);
or U19490 (N_19490,N_13245,N_12781);
and U19491 (N_19491,N_14455,N_10178);
nor U19492 (N_19492,N_10942,N_14909);
nand U19493 (N_19493,N_14841,N_12474);
or U19494 (N_19494,N_13584,N_11286);
nor U19495 (N_19495,N_11150,N_12233);
nor U19496 (N_19496,N_14687,N_14107);
or U19497 (N_19497,N_11654,N_14463);
nand U19498 (N_19498,N_12756,N_14618);
nor U19499 (N_19499,N_11071,N_12041);
nor U19500 (N_19500,N_12607,N_12225);
xor U19501 (N_19501,N_11195,N_14789);
or U19502 (N_19502,N_10652,N_14767);
nor U19503 (N_19503,N_11103,N_11574);
nor U19504 (N_19504,N_10967,N_12454);
xnor U19505 (N_19505,N_12810,N_13211);
and U19506 (N_19506,N_10539,N_13499);
or U19507 (N_19507,N_12816,N_12580);
nand U19508 (N_19508,N_14249,N_10378);
and U19509 (N_19509,N_11985,N_12192);
or U19510 (N_19510,N_10318,N_12780);
nand U19511 (N_19511,N_14569,N_14804);
or U19512 (N_19512,N_11456,N_12115);
xor U19513 (N_19513,N_11544,N_11180);
nand U19514 (N_19514,N_10316,N_11118);
or U19515 (N_19515,N_10685,N_11902);
and U19516 (N_19516,N_14501,N_14836);
nand U19517 (N_19517,N_11080,N_11122);
nand U19518 (N_19518,N_12395,N_12557);
or U19519 (N_19519,N_13310,N_10329);
and U19520 (N_19520,N_14442,N_13212);
nor U19521 (N_19521,N_10484,N_14680);
or U19522 (N_19522,N_11145,N_10458);
nand U19523 (N_19523,N_13102,N_14927);
or U19524 (N_19524,N_12637,N_13101);
nand U19525 (N_19525,N_12288,N_12348);
nand U19526 (N_19526,N_10248,N_13276);
nor U19527 (N_19527,N_13290,N_13201);
or U19528 (N_19528,N_13149,N_13588);
or U19529 (N_19529,N_10832,N_14362);
nand U19530 (N_19530,N_10079,N_12930);
xor U19531 (N_19531,N_13142,N_11819);
and U19532 (N_19532,N_13566,N_11570);
nand U19533 (N_19533,N_12660,N_13933);
or U19534 (N_19534,N_13960,N_12757);
and U19535 (N_19535,N_12312,N_10911);
xor U19536 (N_19536,N_10515,N_13988);
or U19537 (N_19537,N_13658,N_11260);
or U19538 (N_19538,N_10570,N_13739);
xnor U19539 (N_19539,N_11127,N_11697);
or U19540 (N_19540,N_14142,N_11590);
or U19541 (N_19541,N_12858,N_14448);
and U19542 (N_19542,N_12788,N_13060);
nand U19543 (N_19543,N_10343,N_13203);
nand U19544 (N_19544,N_14580,N_13397);
nand U19545 (N_19545,N_14218,N_13609);
nand U19546 (N_19546,N_14148,N_13962);
nor U19547 (N_19547,N_10459,N_10834);
and U19548 (N_19548,N_14713,N_13094);
or U19549 (N_19549,N_11885,N_13606);
xor U19550 (N_19550,N_11946,N_11150);
and U19551 (N_19551,N_12854,N_11954);
nor U19552 (N_19552,N_11781,N_11086);
xnor U19553 (N_19553,N_14176,N_14632);
or U19554 (N_19554,N_14698,N_13636);
nand U19555 (N_19555,N_12272,N_12087);
nor U19556 (N_19556,N_12404,N_12265);
and U19557 (N_19557,N_12740,N_10889);
and U19558 (N_19558,N_12869,N_12890);
or U19559 (N_19559,N_10265,N_11766);
nor U19560 (N_19560,N_11336,N_12113);
nor U19561 (N_19561,N_14086,N_10649);
nand U19562 (N_19562,N_12470,N_13307);
and U19563 (N_19563,N_11764,N_12295);
nand U19564 (N_19564,N_11122,N_10347);
and U19565 (N_19565,N_13235,N_11006);
nor U19566 (N_19566,N_12402,N_11703);
nor U19567 (N_19567,N_12484,N_13049);
and U19568 (N_19568,N_14360,N_12434);
or U19569 (N_19569,N_13292,N_10578);
and U19570 (N_19570,N_11885,N_10775);
or U19571 (N_19571,N_12563,N_10539);
nor U19572 (N_19572,N_12780,N_13754);
nand U19573 (N_19573,N_14700,N_12746);
nand U19574 (N_19574,N_12204,N_12334);
and U19575 (N_19575,N_14996,N_11601);
and U19576 (N_19576,N_13593,N_11504);
nand U19577 (N_19577,N_11826,N_14643);
or U19578 (N_19578,N_13024,N_10494);
and U19579 (N_19579,N_12688,N_12622);
nand U19580 (N_19580,N_10901,N_14284);
nand U19581 (N_19581,N_14628,N_14924);
nand U19582 (N_19582,N_13459,N_10378);
and U19583 (N_19583,N_10367,N_12663);
or U19584 (N_19584,N_11673,N_12003);
nand U19585 (N_19585,N_14900,N_12768);
xor U19586 (N_19586,N_12721,N_13507);
or U19587 (N_19587,N_13797,N_12871);
xnor U19588 (N_19588,N_14661,N_13107);
or U19589 (N_19589,N_14124,N_11117);
nand U19590 (N_19590,N_10238,N_10667);
nand U19591 (N_19591,N_13651,N_13112);
or U19592 (N_19592,N_10832,N_12300);
nor U19593 (N_19593,N_11802,N_14444);
and U19594 (N_19594,N_13275,N_13397);
nor U19595 (N_19595,N_14602,N_12698);
and U19596 (N_19596,N_12849,N_14921);
and U19597 (N_19597,N_10076,N_11429);
nand U19598 (N_19598,N_14001,N_13115);
and U19599 (N_19599,N_10871,N_10226);
nand U19600 (N_19600,N_13001,N_12281);
and U19601 (N_19601,N_14367,N_14349);
nand U19602 (N_19602,N_11779,N_10611);
or U19603 (N_19603,N_13833,N_14745);
or U19604 (N_19604,N_14015,N_12938);
and U19605 (N_19605,N_14903,N_12954);
nor U19606 (N_19606,N_14306,N_11120);
xor U19607 (N_19607,N_14899,N_10560);
and U19608 (N_19608,N_14782,N_10122);
nand U19609 (N_19609,N_11507,N_14537);
xor U19610 (N_19610,N_11418,N_10711);
xnor U19611 (N_19611,N_11196,N_13003);
nor U19612 (N_19612,N_10302,N_14059);
or U19613 (N_19613,N_11439,N_12759);
or U19614 (N_19614,N_12312,N_11920);
xnor U19615 (N_19615,N_12916,N_14452);
nand U19616 (N_19616,N_11451,N_11151);
nor U19617 (N_19617,N_12220,N_11597);
nor U19618 (N_19618,N_13744,N_12373);
nand U19619 (N_19619,N_13802,N_14413);
nor U19620 (N_19620,N_13773,N_12299);
nor U19621 (N_19621,N_14061,N_11732);
or U19622 (N_19622,N_11874,N_11846);
or U19623 (N_19623,N_11950,N_11733);
or U19624 (N_19624,N_11981,N_12432);
or U19625 (N_19625,N_14767,N_11381);
nand U19626 (N_19626,N_14779,N_13644);
nor U19627 (N_19627,N_14449,N_14482);
nor U19628 (N_19628,N_13106,N_11258);
nand U19629 (N_19629,N_11773,N_13367);
nor U19630 (N_19630,N_14464,N_13153);
xnor U19631 (N_19631,N_14846,N_14125);
xnor U19632 (N_19632,N_12323,N_14337);
nor U19633 (N_19633,N_14961,N_12532);
nor U19634 (N_19634,N_14608,N_13517);
and U19635 (N_19635,N_11544,N_10976);
and U19636 (N_19636,N_13321,N_10723);
xor U19637 (N_19637,N_13318,N_12963);
nand U19638 (N_19638,N_13890,N_11743);
or U19639 (N_19639,N_10243,N_14124);
nand U19640 (N_19640,N_12186,N_10944);
or U19641 (N_19641,N_13347,N_14005);
or U19642 (N_19642,N_12802,N_11267);
nand U19643 (N_19643,N_14568,N_11881);
nor U19644 (N_19644,N_14879,N_10421);
nand U19645 (N_19645,N_12599,N_10798);
or U19646 (N_19646,N_12132,N_13241);
nor U19647 (N_19647,N_14104,N_14909);
and U19648 (N_19648,N_10914,N_13655);
or U19649 (N_19649,N_13291,N_13785);
or U19650 (N_19650,N_12048,N_12386);
nor U19651 (N_19651,N_11510,N_12799);
and U19652 (N_19652,N_10662,N_12077);
and U19653 (N_19653,N_13218,N_13661);
or U19654 (N_19654,N_13233,N_12606);
nor U19655 (N_19655,N_14725,N_12631);
and U19656 (N_19656,N_14322,N_14812);
and U19657 (N_19657,N_13083,N_14622);
nand U19658 (N_19658,N_13308,N_13347);
nor U19659 (N_19659,N_14375,N_14684);
and U19660 (N_19660,N_14967,N_11379);
nand U19661 (N_19661,N_11010,N_12233);
or U19662 (N_19662,N_12153,N_13858);
nand U19663 (N_19663,N_12948,N_13634);
or U19664 (N_19664,N_10816,N_10297);
xor U19665 (N_19665,N_13581,N_10224);
nor U19666 (N_19666,N_13918,N_13923);
nor U19667 (N_19667,N_11455,N_10920);
nor U19668 (N_19668,N_10597,N_14767);
nor U19669 (N_19669,N_10451,N_11911);
nand U19670 (N_19670,N_11206,N_14545);
nor U19671 (N_19671,N_13179,N_13509);
or U19672 (N_19672,N_13418,N_11310);
nor U19673 (N_19673,N_10759,N_13266);
xnor U19674 (N_19674,N_13589,N_10420);
or U19675 (N_19675,N_10797,N_11322);
or U19676 (N_19676,N_13215,N_14597);
nor U19677 (N_19677,N_11429,N_10370);
or U19678 (N_19678,N_10458,N_11938);
and U19679 (N_19679,N_10232,N_13141);
or U19680 (N_19680,N_10323,N_11428);
or U19681 (N_19681,N_13063,N_11413);
xor U19682 (N_19682,N_11286,N_10016);
and U19683 (N_19683,N_14633,N_13297);
nor U19684 (N_19684,N_12279,N_13776);
nand U19685 (N_19685,N_14876,N_11649);
or U19686 (N_19686,N_13513,N_10047);
nand U19687 (N_19687,N_11726,N_14948);
nor U19688 (N_19688,N_10080,N_11452);
xor U19689 (N_19689,N_11416,N_13653);
xor U19690 (N_19690,N_10306,N_14450);
nor U19691 (N_19691,N_12332,N_12439);
and U19692 (N_19692,N_11445,N_13764);
nor U19693 (N_19693,N_11636,N_11719);
and U19694 (N_19694,N_14180,N_13484);
and U19695 (N_19695,N_14276,N_11535);
nand U19696 (N_19696,N_13515,N_14570);
nor U19697 (N_19697,N_11779,N_11262);
nor U19698 (N_19698,N_12941,N_10734);
nand U19699 (N_19699,N_14562,N_10399);
or U19700 (N_19700,N_13791,N_13731);
nand U19701 (N_19701,N_14162,N_11253);
xor U19702 (N_19702,N_11498,N_12845);
or U19703 (N_19703,N_12965,N_10328);
or U19704 (N_19704,N_11198,N_10471);
xnor U19705 (N_19705,N_10773,N_10944);
nand U19706 (N_19706,N_12903,N_12626);
and U19707 (N_19707,N_10885,N_11437);
or U19708 (N_19708,N_13988,N_13965);
and U19709 (N_19709,N_10032,N_12418);
nor U19710 (N_19710,N_13671,N_10739);
nor U19711 (N_19711,N_12649,N_11104);
xor U19712 (N_19712,N_13977,N_11502);
nor U19713 (N_19713,N_11010,N_13344);
and U19714 (N_19714,N_11264,N_14522);
nand U19715 (N_19715,N_14821,N_14536);
or U19716 (N_19716,N_10572,N_10817);
and U19717 (N_19717,N_14597,N_12862);
or U19718 (N_19718,N_13002,N_12744);
nor U19719 (N_19719,N_14724,N_12406);
and U19720 (N_19720,N_12481,N_10926);
nand U19721 (N_19721,N_11071,N_13651);
nor U19722 (N_19722,N_12214,N_14706);
nand U19723 (N_19723,N_13488,N_14936);
nor U19724 (N_19724,N_11806,N_12288);
nand U19725 (N_19725,N_11019,N_11227);
xnor U19726 (N_19726,N_13275,N_10965);
nand U19727 (N_19727,N_12450,N_12081);
nand U19728 (N_19728,N_13489,N_10447);
xnor U19729 (N_19729,N_14511,N_10291);
or U19730 (N_19730,N_13706,N_11493);
xor U19731 (N_19731,N_11590,N_14474);
or U19732 (N_19732,N_11305,N_13812);
or U19733 (N_19733,N_14855,N_11289);
nand U19734 (N_19734,N_14161,N_12462);
nand U19735 (N_19735,N_11187,N_13974);
and U19736 (N_19736,N_12474,N_13843);
and U19737 (N_19737,N_14404,N_12429);
nand U19738 (N_19738,N_10729,N_13349);
and U19739 (N_19739,N_14647,N_13250);
xor U19740 (N_19740,N_11015,N_13549);
xor U19741 (N_19741,N_13908,N_14874);
nand U19742 (N_19742,N_10528,N_12098);
and U19743 (N_19743,N_11650,N_14669);
nor U19744 (N_19744,N_10924,N_14105);
or U19745 (N_19745,N_13533,N_11722);
nand U19746 (N_19746,N_14954,N_10860);
and U19747 (N_19747,N_10068,N_12200);
or U19748 (N_19748,N_13506,N_10640);
nand U19749 (N_19749,N_13606,N_14692);
nand U19750 (N_19750,N_13265,N_13713);
nor U19751 (N_19751,N_11564,N_13898);
xnor U19752 (N_19752,N_11560,N_12580);
nand U19753 (N_19753,N_10427,N_11849);
and U19754 (N_19754,N_14502,N_14403);
and U19755 (N_19755,N_13888,N_10360);
and U19756 (N_19756,N_12446,N_14006);
xor U19757 (N_19757,N_12245,N_13445);
and U19758 (N_19758,N_10930,N_10059);
nand U19759 (N_19759,N_11418,N_13364);
xor U19760 (N_19760,N_11288,N_10101);
nand U19761 (N_19761,N_13044,N_12146);
nor U19762 (N_19762,N_14899,N_13403);
nor U19763 (N_19763,N_12257,N_13594);
nand U19764 (N_19764,N_12513,N_11383);
nor U19765 (N_19765,N_11171,N_11639);
nor U19766 (N_19766,N_11613,N_10704);
and U19767 (N_19767,N_12593,N_12317);
nor U19768 (N_19768,N_14830,N_14882);
and U19769 (N_19769,N_10583,N_12370);
and U19770 (N_19770,N_10429,N_14091);
and U19771 (N_19771,N_13825,N_11343);
nand U19772 (N_19772,N_11589,N_11687);
or U19773 (N_19773,N_12618,N_14425);
and U19774 (N_19774,N_14811,N_13331);
nand U19775 (N_19775,N_10595,N_12342);
and U19776 (N_19776,N_12731,N_11545);
nor U19777 (N_19777,N_13998,N_11731);
nand U19778 (N_19778,N_11333,N_10287);
nand U19779 (N_19779,N_13684,N_11940);
or U19780 (N_19780,N_12601,N_10680);
or U19781 (N_19781,N_12252,N_14705);
and U19782 (N_19782,N_11616,N_11527);
or U19783 (N_19783,N_11302,N_12652);
nor U19784 (N_19784,N_11332,N_13349);
or U19785 (N_19785,N_11392,N_14219);
nor U19786 (N_19786,N_13708,N_14009);
or U19787 (N_19787,N_12282,N_11683);
nand U19788 (N_19788,N_10322,N_11638);
and U19789 (N_19789,N_13101,N_10427);
nor U19790 (N_19790,N_11673,N_12038);
nand U19791 (N_19791,N_12071,N_12033);
nand U19792 (N_19792,N_10183,N_12165);
nand U19793 (N_19793,N_12131,N_11629);
or U19794 (N_19794,N_13836,N_12160);
nor U19795 (N_19795,N_11833,N_10028);
nor U19796 (N_19796,N_14291,N_13880);
nand U19797 (N_19797,N_12221,N_10948);
nor U19798 (N_19798,N_14766,N_10310);
nor U19799 (N_19799,N_14042,N_14455);
nand U19800 (N_19800,N_14526,N_12225);
or U19801 (N_19801,N_14855,N_13508);
nand U19802 (N_19802,N_12314,N_10452);
or U19803 (N_19803,N_11665,N_13756);
and U19804 (N_19804,N_13976,N_13034);
and U19805 (N_19805,N_12258,N_11594);
and U19806 (N_19806,N_10074,N_13253);
nor U19807 (N_19807,N_10228,N_14675);
or U19808 (N_19808,N_12562,N_11272);
nand U19809 (N_19809,N_12677,N_11474);
or U19810 (N_19810,N_13224,N_10404);
or U19811 (N_19811,N_13056,N_10953);
and U19812 (N_19812,N_13637,N_12984);
xor U19813 (N_19813,N_12094,N_14992);
nand U19814 (N_19814,N_14172,N_10357);
nor U19815 (N_19815,N_14233,N_13758);
and U19816 (N_19816,N_11146,N_12483);
or U19817 (N_19817,N_13988,N_14717);
nand U19818 (N_19818,N_12559,N_13113);
or U19819 (N_19819,N_13532,N_10010);
nor U19820 (N_19820,N_12516,N_12396);
or U19821 (N_19821,N_11620,N_12384);
and U19822 (N_19822,N_14622,N_14009);
and U19823 (N_19823,N_14572,N_13607);
or U19824 (N_19824,N_12297,N_12414);
nor U19825 (N_19825,N_14094,N_14868);
or U19826 (N_19826,N_13697,N_12211);
and U19827 (N_19827,N_12402,N_10189);
nor U19828 (N_19828,N_11684,N_13852);
nand U19829 (N_19829,N_11163,N_12935);
nor U19830 (N_19830,N_11315,N_14470);
nand U19831 (N_19831,N_12716,N_13062);
or U19832 (N_19832,N_13644,N_11424);
nor U19833 (N_19833,N_10704,N_13942);
or U19834 (N_19834,N_14218,N_12017);
nand U19835 (N_19835,N_13272,N_13707);
nand U19836 (N_19836,N_14888,N_14892);
or U19837 (N_19837,N_12967,N_14909);
nand U19838 (N_19838,N_14069,N_12287);
or U19839 (N_19839,N_13958,N_10471);
nand U19840 (N_19840,N_12816,N_12253);
nand U19841 (N_19841,N_11030,N_14195);
or U19842 (N_19842,N_10606,N_12961);
or U19843 (N_19843,N_11193,N_12175);
nor U19844 (N_19844,N_14371,N_12307);
nand U19845 (N_19845,N_14733,N_11369);
nor U19846 (N_19846,N_14111,N_13769);
or U19847 (N_19847,N_11843,N_13453);
nand U19848 (N_19848,N_12777,N_11137);
or U19849 (N_19849,N_13437,N_11087);
or U19850 (N_19850,N_10503,N_11305);
or U19851 (N_19851,N_12705,N_14028);
nor U19852 (N_19852,N_14829,N_14278);
nor U19853 (N_19853,N_14525,N_13970);
nor U19854 (N_19854,N_14701,N_13124);
nand U19855 (N_19855,N_14322,N_11813);
nand U19856 (N_19856,N_14194,N_14926);
xnor U19857 (N_19857,N_13367,N_10284);
or U19858 (N_19858,N_14199,N_14429);
nor U19859 (N_19859,N_12646,N_12415);
nor U19860 (N_19860,N_13253,N_12724);
nand U19861 (N_19861,N_10889,N_10028);
nor U19862 (N_19862,N_13122,N_12757);
nor U19863 (N_19863,N_14668,N_10456);
nor U19864 (N_19864,N_11258,N_12152);
nand U19865 (N_19865,N_11282,N_12520);
or U19866 (N_19866,N_11010,N_11251);
or U19867 (N_19867,N_11846,N_11736);
nor U19868 (N_19868,N_12883,N_13364);
or U19869 (N_19869,N_11914,N_10262);
nor U19870 (N_19870,N_14486,N_14764);
xor U19871 (N_19871,N_14166,N_11435);
or U19872 (N_19872,N_13239,N_12138);
nor U19873 (N_19873,N_10144,N_11835);
nand U19874 (N_19874,N_10584,N_12970);
xor U19875 (N_19875,N_11527,N_10793);
nor U19876 (N_19876,N_10089,N_13434);
or U19877 (N_19877,N_13540,N_12724);
or U19878 (N_19878,N_11726,N_14081);
nand U19879 (N_19879,N_11009,N_14859);
nor U19880 (N_19880,N_14003,N_13448);
xnor U19881 (N_19881,N_13065,N_14703);
and U19882 (N_19882,N_12233,N_11547);
nor U19883 (N_19883,N_13469,N_14320);
or U19884 (N_19884,N_14013,N_12094);
nand U19885 (N_19885,N_10953,N_12324);
and U19886 (N_19886,N_12199,N_13814);
nand U19887 (N_19887,N_10345,N_10870);
nand U19888 (N_19888,N_14080,N_12441);
and U19889 (N_19889,N_10623,N_13843);
nor U19890 (N_19890,N_11271,N_11970);
nor U19891 (N_19891,N_10242,N_12422);
or U19892 (N_19892,N_13607,N_11616);
or U19893 (N_19893,N_14379,N_13473);
nor U19894 (N_19894,N_13015,N_13837);
and U19895 (N_19895,N_10934,N_12779);
or U19896 (N_19896,N_12889,N_10678);
and U19897 (N_19897,N_12793,N_12211);
and U19898 (N_19898,N_14453,N_14298);
nor U19899 (N_19899,N_11186,N_13889);
and U19900 (N_19900,N_11453,N_12514);
nor U19901 (N_19901,N_14470,N_10626);
and U19902 (N_19902,N_12645,N_12241);
or U19903 (N_19903,N_11520,N_10918);
and U19904 (N_19904,N_14561,N_14001);
nand U19905 (N_19905,N_14828,N_13128);
nand U19906 (N_19906,N_10771,N_12192);
xnor U19907 (N_19907,N_11653,N_12029);
or U19908 (N_19908,N_13641,N_11904);
nor U19909 (N_19909,N_11799,N_13831);
nor U19910 (N_19910,N_12002,N_14684);
xor U19911 (N_19911,N_11232,N_11578);
or U19912 (N_19912,N_10948,N_12012);
and U19913 (N_19913,N_11071,N_10728);
xor U19914 (N_19914,N_12138,N_14050);
nand U19915 (N_19915,N_11487,N_13504);
xor U19916 (N_19916,N_13041,N_14130);
nor U19917 (N_19917,N_10565,N_12491);
nand U19918 (N_19918,N_10085,N_12031);
or U19919 (N_19919,N_11658,N_14528);
and U19920 (N_19920,N_10016,N_12913);
or U19921 (N_19921,N_11191,N_12130);
and U19922 (N_19922,N_14801,N_14348);
nor U19923 (N_19923,N_11349,N_13667);
or U19924 (N_19924,N_13664,N_14488);
nand U19925 (N_19925,N_13105,N_13146);
nand U19926 (N_19926,N_13836,N_14369);
or U19927 (N_19927,N_14578,N_11338);
and U19928 (N_19928,N_12064,N_14658);
or U19929 (N_19929,N_13934,N_12278);
nand U19930 (N_19930,N_14480,N_10007);
nand U19931 (N_19931,N_12274,N_10161);
xor U19932 (N_19932,N_14001,N_14828);
nand U19933 (N_19933,N_13125,N_13907);
and U19934 (N_19934,N_13458,N_12287);
or U19935 (N_19935,N_10181,N_11313);
or U19936 (N_19936,N_10655,N_12728);
nand U19937 (N_19937,N_10699,N_13517);
and U19938 (N_19938,N_12939,N_14935);
nand U19939 (N_19939,N_11633,N_13647);
nor U19940 (N_19940,N_10503,N_10791);
and U19941 (N_19941,N_13421,N_13458);
or U19942 (N_19942,N_12263,N_10128);
and U19943 (N_19943,N_12568,N_11162);
nor U19944 (N_19944,N_11801,N_12598);
or U19945 (N_19945,N_13280,N_11019);
nand U19946 (N_19946,N_13243,N_12616);
or U19947 (N_19947,N_11981,N_11200);
nor U19948 (N_19948,N_13509,N_14242);
and U19949 (N_19949,N_12596,N_12574);
nand U19950 (N_19950,N_10755,N_14514);
or U19951 (N_19951,N_12502,N_14756);
nand U19952 (N_19952,N_12570,N_12167);
nand U19953 (N_19953,N_13758,N_10436);
nand U19954 (N_19954,N_11782,N_14904);
nand U19955 (N_19955,N_10831,N_13076);
and U19956 (N_19956,N_12408,N_12915);
xor U19957 (N_19957,N_14880,N_10771);
and U19958 (N_19958,N_10146,N_13342);
and U19959 (N_19959,N_12576,N_12322);
nor U19960 (N_19960,N_14953,N_13511);
nand U19961 (N_19961,N_10132,N_14161);
xnor U19962 (N_19962,N_11104,N_11892);
or U19963 (N_19963,N_13107,N_11175);
nand U19964 (N_19964,N_10538,N_10292);
nor U19965 (N_19965,N_14572,N_13815);
and U19966 (N_19966,N_13651,N_14865);
nor U19967 (N_19967,N_13938,N_10845);
nor U19968 (N_19968,N_10293,N_14629);
nand U19969 (N_19969,N_14698,N_11951);
nand U19970 (N_19970,N_11309,N_14620);
nand U19971 (N_19971,N_13371,N_14614);
or U19972 (N_19972,N_11188,N_12476);
and U19973 (N_19973,N_13340,N_14879);
nand U19974 (N_19974,N_11421,N_12757);
and U19975 (N_19975,N_11459,N_11183);
nor U19976 (N_19976,N_11383,N_11514);
or U19977 (N_19977,N_11895,N_12399);
nor U19978 (N_19978,N_13970,N_12602);
nand U19979 (N_19979,N_10961,N_11174);
or U19980 (N_19980,N_10964,N_10859);
nand U19981 (N_19981,N_10876,N_14782);
and U19982 (N_19982,N_14511,N_13148);
nand U19983 (N_19983,N_12419,N_11855);
and U19984 (N_19984,N_12316,N_12875);
or U19985 (N_19985,N_14267,N_12642);
nor U19986 (N_19986,N_10416,N_10818);
or U19987 (N_19987,N_14921,N_11338);
or U19988 (N_19988,N_14868,N_12094);
nor U19989 (N_19989,N_13170,N_14592);
nand U19990 (N_19990,N_10290,N_13438);
or U19991 (N_19991,N_12170,N_13047);
xnor U19992 (N_19992,N_12437,N_14161);
nor U19993 (N_19993,N_10939,N_14926);
or U19994 (N_19994,N_13941,N_10407);
xor U19995 (N_19995,N_14482,N_12120);
or U19996 (N_19996,N_12911,N_12390);
xnor U19997 (N_19997,N_11894,N_13738);
nand U19998 (N_19998,N_12925,N_12847);
xor U19999 (N_19999,N_13824,N_14041);
nor UO_0 (O_0,N_18649,N_15007);
and UO_1 (O_1,N_17148,N_18761);
or UO_2 (O_2,N_17549,N_17505);
and UO_3 (O_3,N_18968,N_18438);
nand UO_4 (O_4,N_16670,N_19404);
nor UO_5 (O_5,N_17723,N_19847);
nand UO_6 (O_6,N_15107,N_17390);
or UO_7 (O_7,N_16472,N_18943);
and UO_8 (O_8,N_16057,N_18431);
nand UO_9 (O_9,N_19490,N_16060);
or UO_10 (O_10,N_15978,N_15172);
nand UO_11 (O_11,N_16582,N_17820);
nand UO_12 (O_12,N_16155,N_15158);
nor UO_13 (O_13,N_19809,N_19144);
nor UO_14 (O_14,N_17297,N_16065);
and UO_15 (O_15,N_19194,N_18753);
nor UO_16 (O_16,N_15842,N_17227);
nor UO_17 (O_17,N_16416,N_15723);
or UO_18 (O_18,N_16266,N_16506);
nor UO_19 (O_19,N_15064,N_19257);
nor UO_20 (O_20,N_15132,N_18688);
nor UO_21 (O_21,N_15315,N_19423);
or UO_22 (O_22,N_15281,N_18699);
and UO_23 (O_23,N_17407,N_18713);
and UO_24 (O_24,N_18567,N_16286);
or UO_25 (O_25,N_16733,N_16311);
or UO_26 (O_26,N_19470,N_18878);
nor UO_27 (O_27,N_15681,N_15276);
xnor UO_28 (O_28,N_19603,N_19259);
nand UO_29 (O_29,N_15628,N_17322);
and UO_30 (O_30,N_16487,N_19887);
or UO_31 (O_31,N_16227,N_16971);
or UO_32 (O_32,N_17886,N_16539);
and UO_33 (O_33,N_16666,N_19723);
and UO_34 (O_34,N_16097,N_19042);
and UO_35 (O_35,N_16943,N_17509);
nor UO_36 (O_36,N_17961,N_16451);
or UO_37 (O_37,N_19610,N_17191);
nand UO_38 (O_38,N_15316,N_18013);
nor UO_39 (O_39,N_15484,N_18091);
and UO_40 (O_40,N_19476,N_17526);
and UO_41 (O_41,N_18565,N_16455);
xnor UO_42 (O_42,N_16161,N_19577);
and UO_43 (O_43,N_18366,N_15971);
nand UO_44 (O_44,N_18802,N_18664);
and UO_45 (O_45,N_16383,N_18010);
xor UO_46 (O_46,N_16173,N_19881);
nand UO_47 (O_47,N_16657,N_16265);
nor UO_48 (O_48,N_19836,N_19837);
nor UO_49 (O_49,N_19653,N_18898);
nand UO_50 (O_50,N_16869,N_18864);
xor UO_51 (O_51,N_16120,N_16313);
xnor UO_52 (O_52,N_17144,N_16298);
and UO_53 (O_53,N_18238,N_18625);
xnor UO_54 (O_54,N_18750,N_18412);
and UO_55 (O_55,N_16805,N_18088);
and UO_56 (O_56,N_16691,N_16197);
nor UO_57 (O_57,N_16758,N_17474);
or UO_58 (O_58,N_15921,N_16151);
nor UO_59 (O_59,N_18103,N_19060);
or UO_60 (O_60,N_18200,N_19203);
nor UO_61 (O_61,N_19592,N_16415);
nand UO_62 (O_62,N_15037,N_16446);
xor UO_63 (O_63,N_18150,N_15476);
nor UO_64 (O_64,N_18665,N_19061);
or UO_65 (O_65,N_19954,N_16388);
nand UO_66 (O_66,N_17786,N_15433);
or UO_67 (O_67,N_16684,N_15072);
and UO_68 (O_68,N_16988,N_17596);
and UO_69 (O_69,N_19624,N_19889);
or UO_70 (O_70,N_16577,N_17317);
or UO_71 (O_71,N_16432,N_19830);
or UO_72 (O_72,N_15951,N_17442);
nand UO_73 (O_73,N_19396,N_16111);
nand UO_74 (O_74,N_19591,N_15332);
or UO_75 (O_75,N_18234,N_18759);
nand UO_76 (O_76,N_16548,N_16842);
nor UO_77 (O_77,N_16693,N_15954);
and UO_78 (O_78,N_15749,N_18166);
nand UO_79 (O_79,N_19411,N_19740);
nand UO_80 (O_80,N_16495,N_19466);
and UO_81 (O_81,N_18806,N_15306);
nor UO_82 (O_82,N_17612,N_17703);
and UO_83 (O_83,N_18354,N_15100);
and UO_84 (O_84,N_19155,N_15019);
nor UO_85 (O_85,N_16816,N_18810);
nand UO_86 (O_86,N_15732,N_16689);
or UO_87 (O_87,N_17041,N_19674);
or UO_88 (O_88,N_18774,N_15981);
nor UO_89 (O_89,N_15761,N_19448);
nor UO_90 (O_90,N_19397,N_16190);
nand UO_91 (O_91,N_16361,N_16747);
and UO_92 (O_92,N_16184,N_18380);
nor UO_93 (O_93,N_19403,N_18704);
or UO_94 (O_94,N_17221,N_16041);
nor UO_95 (O_95,N_16283,N_19364);
nor UO_96 (O_96,N_17768,N_16566);
xnor UO_97 (O_97,N_17887,N_17629);
nor UO_98 (O_98,N_15714,N_19020);
nor UO_99 (O_99,N_19129,N_19930);
nand UO_100 (O_100,N_17422,N_15730);
nor UO_101 (O_101,N_18573,N_18156);
and UO_102 (O_102,N_16037,N_15143);
nor UO_103 (O_103,N_16250,N_17534);
nand UO_104 (O_104,N_18757,N_16360);
and UO_105 (O_105,N_16384,N_18016);
xor UO_106 (O_106,N_16713,N_17999);
or UO_107 (O_107,N_17165,N_16620);
xor UO_108 (O_108,N_17329,N_17197);
nor UO_109 (O_109,N_19512,N_17980);
and UO_110 (O_110,N_18002,N_16522);
or UO_111 (O_111,N_16866,N_17518);
nor UO_112 (O_112,N_17065,N_16354);
and UO_113 (O_113,N_18106,N_17239);
and UO_114 (O_114,N_18832,N_18526);
nand UO_115 (O_115,N_17405,N_18468);
and UO_116 (O_116,N_18081,N_16434);
nand UO_117 (O_117,N_17118,N_16838);
nor UO_118 (O_118,N_18075,N_15376);
or UO_119 (O_119,N_17871,N_18187);
or UO_120 (O_120,N_19634,N_19128);
nand UO_121 (O_121,N_19119,N_15139);
xnor UO_122 (O_122,N_18805,N_18775);
or UO_123 (O_123,N_16230,N_16624);
nor UO_124 (O_124,N_17897,N_18529);
nand UO_125 (O_125,N_16382,N_15346);
nand UO_126 (O_126,N_15262,N_16952);
nand UO_127 (O_127,N_19359,N_15341);
nand UO_128 (O_128,N_19385,N_16160);
nand UO_129 (O_129,N_17040,N_18951);
nor UO_130 (O_130,N_16557,N_16514);
nor UO_131 (O_131,N_15534,N_17485);
nor UO_132 (O_132,N_17052,N_18610);
and UO_133 (O_133,N_16132,N_17155);
nand UO_134 (O_134,N_17465,N_18451);
or UO_135 (O_135,N_18432,N_17353);
nand UO_136 (O_136,N_17689,N_16223);
nor UO_137 (O_137,N_17778,N_15024);
or UO_138 (O_138,N_18278,N_19799);
xnor UO_139 (O_139,N_19538,N_16251);
nand UO_140 (O_140,N_15350,N_15848);
nand UO_141 (O_141,N_16245,N_19272);
and UO_142 (O_142,N_16853,N_19794);
or UO_143 (O_143,N_19525,N_18299);
xnor UO_144 (O_144,N_19695,N_15631);
nor UO_145 (O_145,N_15919,N_17210);
nand UO_146 (O_146,N_17904,N_15223);
nor UO_147 (O_147,N_15897,N_19140);
nor UO_148 (O_148,N_19635,N_18603);
or UO_149 (O_149,N_15725,N_18770);
and UO_150 (O_150,N_15349,N_18457);
or UO_151 (O_151,N_15685,N_19981);
or UO_152 (O_152,N_15912,N_16049);
and UO_153 (O_153,N_15461,N_19692);
nor UO_154 (O_154,N_15133,N_16088);
nor UO_155 (O_155,N_16902,N_18701);
and UO_156 (O_156,N_16603,N_18100);
or UO_157 (O_157,N_19824,N_18478);
and UO_158 (O_158,N_19783,N_17995);
or UO_159 (O_159,N_16810,N_17108);
nor UO_160 (O_160,N_19846,N_19668);
or UO_161 (O_161,N_18912,N_18913);
xor UO_162 (O_162,N_16204,N_18495);
or UO_163 (O_163,N_17630,N_17741);
or UO_164 (O_164,N_18054,N_15585);
or UO_165 (O_165,N_17050,N_19711);
xor UO_166 (O_166,N_15013,N_16452);
nand UO_167 (O_167,N_18522,N_18962);
nand UO_168 (O_168,N_15970,N_15129);
and UO_169 (O_169,N_16968,N_17624);
and UO_170 (O_170,N_18110,N_16370);
and UO_171 (O_171,N_19627,N_17367);
and UO_172 (O_172,N_15495,N_17023);
nor UO_173 (O_173,N_17319,N_19189);
nand UO_174 (O_174,N_15156,N_19518);
and UO_175 (O_175,N_17313,N_19308);
nand UO_176 (O_176,N_19307,N_16477);
nand UO_177 (O_177,N_18552,N_18575);
nor UO_178 (O_178,N_16653,N_18858);
or UO_179 (O_179,N_19870,N_17571);
nor UO_180 (O_180,N_19372,N_17361);
xor UO_181 (O_181,N_15200,N_17079);
nand UO_182 (O_182,N_17446,N_17996);
nor UO_183 (O_183,N_17062,N_17335);
or UO_184 (O_184,N_15151,N_16612);
nand UO_185 (O_185,N_16519,N_18637);
and UO_186 (O_186,N_15115,N_15014);
and UO_187 (O_187,N_16763,N_15320);
nor UO_188 (O_188,N_16987,N_17379);
nor UO_189 (O_189,N_19884,N_15003);
nor UO_190 (O_190,N_16659,N_17873);
nand UO_191 (O_191,N_15253,N_17014);
nand UO_192 (O_192,N_16321,N_17912);
nand UO_193 (O_193,N_17365,N_17676);
nor UO_194 (O_194,N_18697,N_18833);
and UO_195 (O_195,N_16780,N_17675);
or UO_196 (O_196,N_17966,N_19110);
or UO_197 (O_197,N_15773,N_15998);
nor UO_198 (O_198,N_15410,N_18952);
nor UO_199 (O_199,N_16078,N_16471);
nor UO_200 (O_200,N_19011,N_16211);
nand UO_201 (O_201,N_18190,N_15793);
or UO_202 (O_202,N_18974,N_15106);
or UO_203 (O_203,N_16328,N_19533);
and UO_204 (O_204,N_16880,N_16158);
or UO_205 (O_205,N_17487,N_18309);
xor UO_206 (O_206,N_15162,N_19242);
and UO_207 (O_207,N_19974,N_17910);
xor UO_208 (O_208,N_15250,N_15237);
nand UO_209 (O_209,N_19088,N_16808);
and UO_210 (O_210,N_16395,N_19588);
nand UO_211 (O_211,N_15302,N_18365);
or UO_212 (O_212,N_19206,N_17936);
or UO_213 (O_213,N_19178,N_19219);
or UO_214 (O_214,N_15458,N_18225);
nor UO_215 (O_215,N_17240,N_15050);
or UO_216 (O_216,N_15896,N_19728);
nand UO_217 (O_217,N_19299,N_19698);
nor UO_218 (O_218,N_17756,N_17266);
and UO_219 (O_219,N_19891,N_15508);
nor UO_220 (O_220,N_16007,N_15811);
nand UO_221 (O_221,N_17718,N_17145);
and UO_222 (O_222,N_15471,N_17383);
and UO_223 (O_223,N_19014,N_19945);
or UO_224 (O_224,N_17759,N_17073);
nor UO_225 (O_225,N_18071,N_18420);
or UO_226 (O_226,N_15418,N_18494);
nand UO_227 (O_227,N_16921,N_15591);
nor UO_228 (O_228,N_19217,N_19554);
xnor UO_229 (O_229,N_16473,N_17906);
nor UO_230 (O_230,N_16532,N_15383);
nand UO_231 (O_231,N_17994,N_18658);
or UO_232 (O_232,N_16903,N_18542);
nand UO_233 (O_233,N_17782,N_18941);
nand UO_234 (O_234,N_16925,N_15527);
nand UO_235 (O_235,N_18095,N_15928);
and UO_236 (O_236,N_15940,N_19682);
nand UO_237 (O_237,N_15385,N_16962);
or UO_238 (O_238,N_18749,N_16525);
nor UO_239 (O_239,N_16549,N_18674);
nand UO_240 (O_240,N_19116,N_18696);
nor UO_241 (O_241,N_19828,N_15096);
nand UO_242 (O_242,N_18053,N_18535);
and UO_243 (O_243,N_17781,N_16623);
xor UO_244 (O_244,N_16789,N_17628);
nand UO_245 (O_245,N_15199,N_19139);
or UO_246 (O_246,N_17730,N_16505);
xnor UO_247 (O_247,N_18728,N_17397);
and UO_248 (O_248,N_16708,N_15536);
or UO_249 (O_249,N_19233,N_16671);
nor UO_250 (O_250,N_16084,N_15803);
nand UO_251 (O_251,N_15326,N_15309);
and UO_252 (O_252,N_18406,N_15056);
and UO_253 (O_253,N_18639,N_18385);
nand UO_254 (O_254,N_17924,N_17593);
or UO_255 (O_255,N_16504,N_15000);
nor UO_256 (O_256,N_19036,N_18230);
and UO_257 (O_257,N_18007,N_15266);
nor UO_258 (O_258,N_16106,N_17874);
nand UO_259 (O_259,N_18690,N_19105);
or UO_260 (O_260,N_17229,N_17029);
or UO_261 (O_261,N_15179,N_15322);
or UO_262 (O_262,N_19795,N_19278);
and UO_263 (O_263,N_18397,N_15043);
xor UO_264 (O_264,N_16734,N_16819);
nand UO_265 (O_265,N_15916,N_15157);
nand UO_266 (O_266,N_17137,N_16464);
or UO_267 (O_267,N_19422,N_16494);
nor UO_268 (O_268,N_17671,N_19157);
nand UO_269 (O_269,N_16064,N_19399);
xnor UO_270 (O_270,N_18289,N_19328);
and UO_271 (O_271,N_17194,N_19851);
xor UO_272 (O_272,N_19633,N_15230);
nand UO_273 (O_273,N_15123,N_18598);
nor UO_274 (O_274,N_15573,N_18694);
or UO_275 (O_275,N_17708,N_16811);
nand UO_276 (O_276,N_16293,N_17214);
and UO_277 (O_277,N_17774,N_19387);
or UO_278 (O_278,N_17889,N_19125);
and UO_279 (O_279,N_19949,N_15756);
xor UO_280 (O_280,N_15336,N_15864);
nor UO_281 (O_281,N_19858,N_18956);
and UO_282 (O_282,N_17370,N_17440);
nand UO_283 (O_283,N_19748,N_15593);
xor UO_284 (O_284,N_16428,N_19504);
or UO_285 (O_285,N_15816,N_15218);
nor UO_286 (O_286,N_15128,N_18987);
and UO_287 (O_287,N_15190,N_16255);
nand UO_288 (O_288,N_18734,N_19860);
or UO_289 (O_289,N_18812,N_16741);
nor UO_290 (O_290,N_18467,N_17316);
and UO_291 (O_291,N_19195,N_19706);
nand UO_292 (O_292,N_18957,N_18989);
and UO_293 (O_293,N_17410,N_18825);
or UO_294 (O_294,N_19268,N_19790);
nor UO_295 (O_295,N_18969,N_18964);
nand UO_296 (O_296,N_19853,N_15985);
or UO_297 (O_297,N_17153,N_15224);
nor UO_298 (O_298,N_19408,N_16417);
nor UO_299 (O_299,N_15833,N_16220);
nand UO_300 (O_300,N_15070,N_15746);
nor UO_301 (O_301,N_17270,N_15615);
nand UO_302 (O_302,N_16716,N_17441);
and UO_303 (O_303,N_15255,N_17539);
or UO_304 (O_304,N_16222,N_15890);
nor UO_305 (O_305,N_17072,N_16901);
or UO_306 (O_306,N_16202,N_16583);
nand UO_307 (O_307,N_17501,N_17622);
and UO_308 (O_308,N_17706,N_15878);
and UO_309 (O_309,N_18312,N_15541);
or UO_310 (O_310,N_17085,N_19933);
nand UO_311 (O_311,N_19762,N_17687);
nor UO_312 (O_312,N_19305,N_16209);
xnor UO_313 (O_313,N_18151,N_15435);
or UO_314 (O_314,N_17794,N_15339);
and UO_315 (O_315,N_17445,N_17942);
or UO_316 (O_316,N_19644,N_15695);
xnor UO_317 (O_317,N_18814,N_19076);
and UO_318 (O_318,N_15022,N_18576);
or UO_319 (O_319,N_18772,N_17780);
xnor UO_320 (O_320,N_19663,N_16710);
nor UO_321 (O_321,N_19885,N_16697);
nand UO_322 (O_322,N_15930,N_19713);
and UO_323 (O_323,N_18816,N_17664);
and UO_324 (O_324,N_18656,N_15693);
and UO_325 (O_325,N_16721,N_16679);
nor UO_326 (O_326,N_18771,N_19226);
nor UO_327 (O_327,N_17056,N_15360);
nand UO_328 (O_328,N_17017,N_17638);
xnor UO_329 (O_329,N_16774,N_19587);
nor UO_330 (O_330,N_18521,N_15328);
nand UO_331 (O_331,N_15203,N_19877);
and UO_332 (O_332,N_19875,N_15727);
and UO_333 (O_333,N_15044,N_19551);
or UO_334 (O_334,N_19276,N_16674);
nor UO_335 (O_335,N_17089,N_18792);
nand UO_336 (O_336,N_16807,N_16114);
nor UO_337 (O_337,N_15668,N_15026);
or UO_338 (O_338,N_19555,N_16405);
nand UO_339 (O_339,N_19872,N_17574);
and UO_340 (O_340,N_15267,N_19031);
nand UO_341 (O_341,N_19501,N_16601);
and UO_342 (O_342,N_18676,N_18523);
nand UO_343 (O_343,N_17101,N_16840);
or UO_344 (O_344,N_16595,N_15915);
or UO_345 (O_345,N_16849,N_17607);
and UO_346 (O_346,N_16813,N_15491);
and UO_347 (O_347,N_19979,N_15983);
or UO_348 (O_348,N_16099,N_16180);
and UO_349 (O_349,N_15721,N_17340);
nand UO_350 (O_350,N_17952,N_19109);
and UO_351 (O_351,N_15895,N_15497);
nor UO_352 (O_352,N_15412,N_16662);
or UO_353 (O_353,N_19353,N_18837);
and UO_354 (O_354,N_17958,N_16731);
xnor UO_355 (O_355,N_17790,N_17369);
nand UO_356 (O_356,N_16996,N_19279);
nand UO_357 (O_357,N_16579,N_17251);
nand UO_358 (O_358,N_18907,N_16023);
nor UO_359 (O_359,N_18279,N_16890);
nor UO_360 (O_360,N_15119,N_16823);
or UO_361 (O_361,N_19833,N_18465);
or UO_362 (O_362,N_19960,N_15041);
or UO_363 (O_363,N_18601,N_19688);
and UO_364 (O_364,N_16559,N_19694);
nand UO_365 (O_365,N_15432,N_15662);
or UO_366 (O_366,N_18211,N_19322);
nand UO_367 (O_367,N_15015,N_15236);
or UO_368 (O_368,N_18390,N_18471);
and UO_369 (O_369,N_15280,N_17668);
and UO_370 (O_370,N_17005,N_15856);
nand UO_371 (O_371,N_19802,N_17296);
or UO_372 (O_372,N_17585,N_18396);
and UO_373 (O_373,N_18120,N_17838);
and UO_374 (O_374,N_17193,N_19229);
or UO_375 (O_375,N_17181,N_16711);
nand UO_376 (O_376,N_17081,N_18580);
and UO_377 (O_377,N_19499,N_19453);
xor UO_378 (O_378,N_19536,N_18698);
nand UO_379 (O_379,N_18970,N_15545);
nand UO_380 (O_380,N_17553,N_15321);
nand UO_381 (O_381,N_15138,N_17990);
nand UO_382 (O_382,N_17477,N_15170);
and UO_383 (O_383,N_18624,N_15171);
nand UO_384 (O_384,N_19942,N_15514);
or UO_385 (O_385,N_16225,N_18766);
and UO_386 (O_386,N_17196,N_16143);
and UO_387 (O_387,N_17180,N_16873);
nand UO_388 (O_388,N_17746,N_19906);
nor UO_389 (O_389,N_15987,N_18651);
and UO_390 (O_390,N_17413,N_19817);
nor UO_391 (O_391,N_18443,N_15305);
nor UO_392 (O_392,N_16034,N_16331);
or UO_393 (O_393,N_19452,N_15411);
xnor UO_394 (O_394,N_18003,N_15430);
nor UO_395 (O_395,N_19911,N_19106);
nor UO_396 (O_396,N_18283,N_19211);
or UO_397 (O_397,N_19888,N_15755);
and UO_398 (O_398,N_17154,N_15087);
or UO_399 (O_399,N_18561,N_15574);
nand UO_400 (O_400,N_18558,N_17821);
and UO_401 (O_401,N_19463,N_16993);
nand UO_402 (O_402,N_19366,N_17070);
xnor UO_403 (O_403,N_17479,N_15726);
and UO_404 (O_404,N_18615,N_16589);
xnor UO_405 (O_405,N_16492,N_16000);
nand UO_406 (O_406,N_17749,N_15215);
nor UO_407 (O_407,N_15269,N_16627);
and UO_408 (O_408,N_17614,N_19969);
nor UO_409 (O_409,N_16110,N_19134);
nand UO_410 (O_410,N_19440,N_16172);
nand UO_411 (O_411,N_18301,N_15283);
or UO_412 (O_412,N_17158,N_19045);
nor UO_413 (O_413,N_18963,N_19039);
and UO_414 (O_414,N_15790,N_17491);
nor UO_415 (O_415,N_16288,N_17719);
nor UO_416 (O_416,N_16994,N_18901);
or UO_417 (O_417,N_18873,N_18270);
xnor UO_418 (O_418,N_17374,N_17895);
nand UO_419 (O_419,N_16296,N_18714);
nand UO_420 (O_420,N_15565,N_17927);
nor UO_421 (O_421,N_15871,N_18203);
nand UO_422 (O_422,N_17293,N_16435);
nor UO_423 (O_423,N_15039,N_16010);
nor UO_424 (O_424,N_18219,N_16584);
nand UO_425 (O_425,N_19277,N_19444);
xnor UO_426 (O_426,N_17276,N_15994);
or UO_427 (O_427,N_19863,N_17439);
nand UO_428 (O_428,N_19773,N_19731);
and UO_429 (O_429,N_18796,N_18577);
and UO_430 (O_430,N_18992,N_16366);
or UO_431 (O_431,N_17829,N_16485);
or UO_432 (O_432,N_19642,N_19526);
xor UO_433 (O_433,N_16350,N_19368);
or UO_434 (O_434,N_15210,N_17617);
nand UO_435 (O_435,N_15563,N_19816);
or UO_436 (O_436,N_17716,N_15807);
nand UO_437 (O_437,N_18860,N_17496);
nor UO_438 (O_438,N_16934,N_19021);
nor UO_439 (O_439,N_17854,N_16013);
nor UO_440 (O_440,N_15991,N_15607);
and UO_441 (O_441,N_15325,N_16900);
nand UO_442 (O_442,N_15144,N_16746);
nand UO_443 (O_443,N_16597,N_19047);
nor UO_444 (O_444,N_15976,N_17604);
or UO_445 (O_445,N_16730,N_18514);
nand UO_446 (O_446,N_18326,N_17851);
nand UO_447 (O_447,N_15247,N_17970);
and UO_448 (O_448,N_17536,N_16437);
nor UO_449 (O_449,N_15380,N_15415);
and UO_450 (O_450,N_16919,N_17126);
nand UO_451 (O_451,N_19481,N_18090);
nor UO_452 (O_452,N_17212,N_18622);
nand UO_453 (O_453,N_17142,N_17391);
or UO_454 (O_454,N_19212,N_17171);
or UO_455 (O_455,N_15549,N_15677);
or UO_456 (O_456,N_18980,N_15823);
and UO_457 (O_457,N_15313,N_19114);
or UO_458 (O_458,N_16257,N_15038);
and UO_459 (O_459,N_17876,N_19344);
nand UO_460 (O_460,N_16308,N_19460);
and UO_461 (O_461,N_19205,N_19787);
nor UO_462 (O_462,N_15924,N_16163);
or UO_463 (O_463,N_16751,N_17803);
xnor UO_464 (O_464,N_16337,N_19651);
nor UO_465 (O_465,N_16409,N_15844);
and UO_466 (O_466,N_15486,N_19750);
nor UO_467 (O_467,N_19753,N_15675);
and UO_468 (O_468,N_18448,N_17688);
or UO_469 (O_469,N_17850,N_19376);
nand UO_470 (O_470,N_15487,N_18865);
nor UO_471 (O_471,N_16867,N_19213);
nor UO_472 (O_472,N_16563,N_19121);
nand UO_473 (O_473,N_17121,N_19473);
nand UO_474 (O_474,N_18178,N_15712);
nand UO_475 (O_475,N_17475,N_18925);
nand UO_476 (O_476,N_18466,N_18485);
nand UO_477 (O_477,N_15051,N_17058);
nor UO_478 (O_478,N_15225,N_19778);
xnor UO_479 (O_479,N_16486,N_18174);
and UO_480 (O_480,N_18971,N_17339);
and UO_481 (O_481,N_17324,N_15462);
nand UO_482 (O_482,N_19521,N_18729);
xnor UO_483 (O_483,N_19742,N_17564);
or UO_484 (O_484,N_15509,N_16241);
nand UO_485 (O_485,N_15455,N_19545);
nand UO_486 (O_486,N_17039,N_17457);
nand UO_487 (O_487,N_15165,N_16829);
nor UO_488 (O_488,N_18844,N_17993);
or UO_489 (O_489,N_16374,N_16134);
and UO_490 (O_490,N_19874,N_16775);
nand UO_491 (O_491,N_19931,N_16314);
and UO_492 (O_492,N_16668,N_19494);
and UO_493 (O_493,N_17368,N_19509);
nand UO_494 (O_494,N_15686,N_19446);
and UO_495 (O_495,N_15990,N_17366);
or UO_496 (O_496,N_15368,N_17576);
or UO_497 (O_497,N_17362,N_17054);
nor UO_498 (O_498,N_18984,N_16149);
or UO_499 (O_499,N_15758,N_19928);
and UO_500 (O_500,N_15475,N_19883);
nand UO_501 (O_501,N_18922,N_17386);
and UO_502 (O_502,N_16884,N_18257);
nand UO_503 (O_503,N_16246,N_17068);
nor UO_504 (O_504,N_15813,N_18997);
nor UO_505 (O_505,N_16358,N_15271);
nor UO_506 (O_506,N_15904,N_16407);
and UO_507 (O_507,N_17454,N_18492);
nor UO_508 (O_508,N_15760,N_16856);
nand UO_509 (O_509,N_18063,N_18846);
nor UO_510 (O_510,N_17423,N_16018);
and UO_511 (O_511,N_18756,N_15893);
or UO_512 (O_512,N_19892,N_15244);
nor UO_513 (O_513,N_18596,N_19621);
nor UO_514 (O_514,N_19656,N_19686);
or UO_515 (O_515,N_17772,N_19345);
nor UO_516 (O_516,N_16553,N_15818);
nor UO_517 (O_517,N_19222,N_19298);
nand UO_518 (O_518,N_19244,N_16044);
or UO_519 (O_519,N_16578,N_19821);
and UO_520 (O_520,N_19230,N_15010);
and UO_521 (O_521,N_19122,N_19434);
and UO_522 (O_522,N_18679,N_16944);
or UO_523 (O_523,N_15579,N_18029);
nand UO_524 (O_524,N_16187,N_17591);
or UO_525 (O_525,N_17681,N_19867);
nand UO_526 (O_526,N_15887,N_16947);
or UO_527 (O_527,N_19745,N_19113);
nand UO_528 (O_528,N_16586,N_19987);
and UO_529 (O_529,N_19161,N_15468);
or UO_530 (O_530,N_16826,N_16294);
or UO_531 (O_531,N_18206,N_18998);
and UO_532 (O_532,N_19604,N_15988);
nand UO_533 (O_533,N_16963,N_16636);
and UO_534 (O_534,N_15189,N_16784);
or UO_535 (O_535,N_15754,N_17930);
and UO_536 (O_536,N_18946,N_17665);
nor UO_537 (O_537,N_19339,N_17766);
nor UO_538 (O_538,N_19123,N_18249);
nor UO_539 (O_539,N_15304,N_17972);
or UO_540 (O_540,N_15530,N_16213);
nor UO_541 (O_541,N_16082,N_17395);
nand UO_542 (O_542,N_17736,N_15097);
nand UO_543 (O_543,N_15572,N_17810);
nor UO_544 (O_544,N_15620,N_15494);
nor UO_545 (O_545,N_19825,N_17831);
nand UO_546 (O_546,N_18189,N_18118);
and UO_547 (O_547,N_16936,N_16107);
nor UO_548 (O_548,N_17608,N_18079);
and UO_549 (O_549,N_19447,N_18000);
nand UO_550 (O_550,N_18733,N_19303);
nor UO_551 (O_551,N_16385,N_16369);
or UO_552 (O_552,N_17594,N_15092);
nand UO_553 (O_553,N_17863,N_19876);
nor UO_554 (O_554,N_15715,N_19561);
and UO_555 (O_555,N_17235,N_18209);
nor UO_556 (O_556,N_18194,N_18253);
nor UO_557 (O_557,N_15957,N_18708);
nand UO_558 (O_558,N_19670,N_19607);
nor UO_559 (O_559,N_16812,N_17466);
xnor UO_560 (O_560,N_18916,N_16027);
nor UO_561 (O_561,N_19534,N_15613);
or UO_562 (O_562,N_19182,N_17667);
nor UO_563 (O_563,N_19746,N_15057);
or UO_564 (O_564,N_15684,N_18107);
and UO_565 (O_565,N_15245,N_17320);
or UO_566 (O_566,N_17203,N_18269);
and UO_567 (O_567,N_16261,N_19486);
or UO_568 (O_568,N_15300,N_17414);
nand UO_569 (O_569,N_17643,N_17908);
and UO_570 (O_570,N_19160,N_15287);
nor UO_571 (O_571,N_17330,N_19370);
xnor UO_572 (O_572,N_19218,N_15927);
nand UO_573 (O_573,N_19975,N_19034);
and UO_574 (O_574,N_18499,N_18815);
or UO_575 (O_575,N_16463,N_18197);
and UO_576 (O_576,N_18486,N_16339);
or UO_577 (O_577,N_18069,N_15016);
or UO_578 (O_578,N_16749,N_19868);
nor UO_579 (O_579,N_16699,N_15002);
and UO_580 (O_580,N_16070,N_18232);
and UO_581 (O_581,N_17502,N_19179);
nor UO_582 (O_582,N_15903,N_17113);
xnor UO_583 (O_583,N_16568,N_16752);
and UO_584 (O_584,N_18272,N_18906);
nor UO_585 (O_585,N_16637,N_17818);
or UO_586 (O_586,N_19075,N_18294);
and UO_587 (O_587,N_16028,N_16871);
nand UO_588 (O_588,N_19840,N_15554);
and UO_589 (O_589,N_16176,N_18965);
nand UO_590 (O_590,N_19815,N_15664);
nand UO_591 (O_591,N_19003,N_19275);
or UO_592 (O_592,N_17537,N_18583);
nand UO_593 (O_593,N_17734,N_15974);
nand UO_594 (O_594,N_17544,N_18305);
xor UO_595 (O_595,N_19721,N_19620);
nand UO_596 (O_596,N_19565,N_19826);
and UO_597 (O_597,N_15053,N_15469);
nor UO_598 (O_598,N_19631,N_17130);
or UO_599 (O_599,N_18813,N_15969);
xor UO_600 (O_600,N_17650,N_16997);
nor UO_601 (O_601,N_16843,N_16864);
nand UO_602 (O_602,N_19207,N_15065);
xor UO_603 (O_603,N_19970,N_16528);
or UO_604 (O_604,N_15967,N_15489);
xnor UO_605 (O_605,N_17464,N_18462);
nor UO_606 (O_606,N_18045,N_16717);
or UO_607 (O_607,N_19660,N_19570);
xor UO_608 (O_608,N_18310,N_19562);
and UO_609 (O_609,N_15420,N_18460);
nor UO_610 (O_610,N_18038,N_15825);
nor UO_611 (O_611,N_18924,N_16551);
nor UO_612 (O_612,N_15744,N_18553);
nor UO_613 (O_613,N_15384,N_15343);
or UO_614 (O_614,N_16353,N_18152);
nor UO_615 (O_615,N_16897,N_16439);
and UO_616 (O_616,N_18236,N_15941);
nand UO_617 (O_617,N_18470,N_18322);
nor UO_618 (O_618,N_16558,N_19752);
or UO_619 (O_619,N_15279,N_16103);
or UO_620 (O_620,N_17714,N_19321);
and UO_621 (O_621,N_15590,N_15616);
and UO_622 (O_622,N_16252,N_19791);
nand UO_623 (O_623,N_17740,N_19373);
or UO_624 (O_624,N_18668,N_17484);
or UO_625 (O_625,N_18456,N_18760);
and UO_626 (O_626,N_18543,N_16404);
and UO_627 (O_627,N_15521,N_19349);
xnor UO_628 (O_628,N_18001,N_17738);
nand UO_629 (O_629,N_15586,N_17114);
and UO_630 (O_630,N_15876,N_18335);
nand UO_631 (O_631,N_19496,N_15704);
nor UO_632 (O_632,N_16429,N_16304);
or UO_633 (O_633,N_17760,N_18635);
and UO_634 (O_634,N_17898,N_19772);
and UO_635 (O_635,N_18154,N_17347);
nand UO_636 (O_636,N_18590,N_19082);
nor UO_637 (O_637,N_15787,N_17957);
or UO_638 (O_638,N_17449,N_17822);
nor UO_639 (O_639,N_19792,N_15979);
or UO_640 (O_640,N_17636,N_17525);
nor UO_641 (O_641,N_15373,N_17275);
or UO_642 (O_642,N_17905,N_18191);
nor UO_643 (O_643,N_18886,N_19556);
nand UO_644 (O_644,N_18928,N_16596);
nand UO_645 (O_645,N_18165,N_18762);
or UO_646 (O_646,N_18262,N_19506);
nand UO_647 (O_647,N_15382,N_15622);
and UO_648 (O_648,N_18508,N_17215);
nand UO_649 (O_649,N_16011,N_18387);
or UO_650 (O_650,N_16726,N_17499);
or UO_651 (O_651,N_19813,N_18363);
and UO_652 (O_652,N_15193,N_18513);
nor UO_653 (O_653,N_16116,N_17758);
nand UO_654 (O_654,N_19549,N_17879);
nand UO_655 (O_655,N_17209,N_19789);
nand UO_656 (O_656,N_19502,N_18560);
or UO_657 (O_657,N_17901,N_15962);
and UO_658 (O_658,N_18351,N_16125);
or UO_659 (O_659,N_15216,N_15260);
nand UO_660 (O_660,N_15397,N_17808);
and UO_661 (O_661,N_16215,N_16425);
or UO_662 (O_662,N_16408,N_17301);
nand UO_663 (O_663,N_19315,N_18383);
nand UO_664 (O_664,N_16145,N_19484);
nand UO_665 (O_665,N_16850,N_18422);
and UO_666 (O_666,N_17837,N_19197);
nand UO_667 (O_667,N_16402,N_17314);
or UO_668 (O_668,N_17865,N_15342);
and UO_669 (O_669,N_18005,N_18893);
or UO_670 (O_670,N_19751,N_17160);
xor UO_671 (O_671,N_17258,N_18130);
and UO_672 (O_672,N_18228,N_15734);
and UO_673 (O_673,N_18401,N_19083);
or UO_674 (O_674,N_15122,N_15802);
nor UO_675 (O_675,N_15299,N_19176);
and UO_676 (O_676,N_17864,N_15556);
nor UO_677 (O_677,N_15778,N_19839);
and UO_678 (O_678,N_19727,N_16965);
or UO_679 (O_679,N_15239,N_15676);
nor UO_680 (O_680,N_19167,N_16660);
or UO_681 (O_681,N_18082,N_16663);
nand UO_682 (O_682,N_18923,N_19464);
nor UO_683 (O_683,N_15795,N_17204);
nand UO_684 (O_684,N_17468,N_18687);
nand UO_685 (O_685,N_15030,N_17960);
or UO_686 (O_686,N_15699,N_15112);
and UO_687 (O_687,N_16095,N_15197);
or UO_688 (O_688,N_17247,N_17773);
or UO_689 (O_689,N_16009,N_17257);
nand UO_690 (O_690,N_17903,N_17046);
nor UO_691 (O_691,N_15735,N_17069);
nor UO_692 (O_692,N_17104,N_17610);
nand UO_693 (O_693,N_17406,N_15578);
nand UO_694 (O_694,N_15597,N_18483);
nor UO_695 (O_695,N_16980,N_19010);
and UO_696 (O_696,N_19412,N_17812);
nor UO_697 (O_697,N_15571,N_19142);
nor UO_698 (O_698,N_15931,N_19081);
nor UO_699 (O_699,N_18336,N_17157);
xor UO_700 (O_700,N_19690,N_18403);
and UO_701 (O_701,N_19678,N_19126);
and UO_702 (O_702,N_16373,N_16772);
and UO_703 (O_703,N_16393,N_19159);
nand UO_704 (O_704,N_15358,N_16561);
and UO_705 (O_705,N_19894,N_16830);
and UO_706 (O_706,N_16556,N_18859);
nor UO_707 (O_707,N_17115,N_15798);
nand UO_708 (O_708,N_18052,N_15551);
or UO_709 (O_709,N_19908,N_18669);
nand UO_710 (O_710,N_17834,N_18845);
and UO_711 (O_711,N_15198,N_19602);
and UO_712 (O_712,N_15542,N_16682);
nor UO_713 (O_713,N_19421,N_19586);
and UO_714 (O_714,N_16152,N_19051);
or UO_715 (O_715,N_16825,N_15398);
and UO_716 (O_716,N_16333,N_19707);
xor UO_717 (O_717,N_16680,N_15598);
xnor UO_718 (O_718,N_16712,N_19703);
or UO_719 (O_719,N_17077,N_16285);
nor UO_720 (O_720,N_15046,N_15526);
or UO_721 (O_721,N_16210,N_18484);
nand UO_722 (O_722,N_18167,N_18160);
nand UO_723 (O_723,N_16119,N_18650);
or UO_724 (O_724,N_19769,N_19726);
nand UO_725 (O_725,N_19169,N_18417);
and UO_726 (O_726,N_15757,N_19595);
nor UO_727 (O_727,N_17563,N_17860);
and UO_728 (O_728,N_18605,N_18654);
nand UO_729 (O_729,N_17682,N_15329);
or UO_730 (O_730,N_18357,N_19932);
nand UO_731 (O_731,N_17030,N_15846);
nand UO_732 (O_732,N_19483,N_16729);
nor UO_733 (O_733,N_15294,N_18824);
or UO_734 (O_734,N_19382,N_16759);
nand UO_735 (O_735,N_19956,N_15400);
and UO_736 (O_736,N_19019,N_15575);
and UO_737 (O_737,N_15869,N_17381);
nor UO_738 (O_738,N_15539,N_16835);
and UO_739 (O_739,N_15131,N_19316);
xor UO_740 (O_740,N_15679,N_19571);
or UO_741 (O_741,N_17015,N_15606);
nor UO_742 (O_742,N_19026,N_18817);
and UO_743 (O_743,N_18933,N_17044);
and UO_744 (O_744,N_18064,N_16198);
and UO_745 (O_745,N_19094,N_15792);
nor UO_746 (O_746,N_16083,N_18988);
nor UO_747 (O_747,N_16481,N_16984);
nor UO_748 (O_748,N_19280,N_16723);
xnor UO_749 (O_749,N_15389,N_19058);
nand UO_750 (O_750,N_18181,N_19346);
nand UO_751 (O_751,N_15018,N_19469);
or UO_752 (O_752,N_18012,N_15184);
nand UO_753 (O_753,N_16517,N_18442);
xor UO_754 (O_754,N_17712,N_19468);
nor UO_755 (O_755,N_15647,N_16592);
nand UO_756 (O_756,N_18659,N_15705);
nor UO_757 (O_757,N_17562,N_19360);
nand UO_758 (O_758,N_15703,N_18948);
nor UO_759 (O_759,N_16348,N_18306);
nor UO_760 (O_760,N_19768,N_15118);
nand UO_761 (O_761,N_16868,N_15035);
and UO_762 (O_762,N_17882,N_19164);
nand UO_763 (O_763,N_19563,N_18618);
nor UO_764 (O_764,N_15920,N_18578);
nand UO_765 (O_765,N_19231,N_17911);
nand UO_766 (O_766,N_18288,N_17348);
xor UO_767 (O_767,N_16920,N_18628);
and UO_768 (O_768,N_15331,N_15923);
or UO_769 (O_769,N_16979,N_16336);
nand UO_770 (O_770,N_18843,N_18680);
nor UO_771 (O_771,N_15449,N_17735);
nand UO_772 (O_772,N_15145,N_19569);
nand UO_773 (O_773,N_15289,N_16422);
nand UO_774 (O_774,N_18265,N_15812);
xor UO_775 (O_775,N_19177,N_18179);
nor UO_776 (O_776,N_17300,N_18501);
nor UO_777 (O_777,N_18936,N_17232);
nor UO_778 (O_778,N_19287,N_15088);
nor UO_779 (O_779,N_17452,N_15722);
or UO_780 (O_780,N_17447,N_15370);
nor UO_781 (O_781,N_18059,N_19878);
and UO_782 (O_782,N_19032,N_17694);
and UO_783 (O_783,N_17211,N_17064);
or UO_784 (O_784,N_15369,N_15399);
and UO_785 (O_785,N_18085,N_18518);
nor UO_786 (O_786,N_18260,N_19283);
and UO_787 (O_787,N_17739,N_16765);
and UO_788 (O_788,N_19990,N_19027);
nor UO_789 (O_789,N_18721,N_19462);
xnor UO_790 (O_790,N_19285,N_19171);
nand UO_791 (O_791,N_16511,N_17870);
nand UO_792 (O_792,N_18255,N_16303);
or UO_793 (O_793,N_15314,N_19953);
or UO_794 (O_794,N_15752,N_15080);
or UO_795 (O_795,N_18828,N_17680);
nor UO_796 (O_796,N_16542,N_19622);
and UO_797 (O_797,N_16948,N_16226);
and UO_798 (O_798,N_19215,N_19361);
nand UO_799 (O_799,N_16779,N_16076);
nand UO_800 (O_800,N_17093,N_18015);
or UO_801 (O_801,N_15503,N_19940);
nor UO_802 (O_802,N_15102,N_15619);
and UO_803 (O_803,N_16630,N_19038);
and UO_804 (O_804,N_16445,N_15029);
nand UO_805 (O_805,N_16909,N_15095);
nor UO_806 (O_806,N_16496,N_15640);
nand UO_807 (O_807,N_17249,N_18904);
nand UO_808 (O_808,N_18769,N_17926);
nor UO_809 (O_809,N_18453,N_15364);
and UO_810 (O_810,N_18132,N_17311);
nand UO_811 (O_811,N_19735,N_15739);
or UO_812 (O_812,N_16576,N_15537);
and UO_813 (O_813,N_15964,N_19059);
or UO_814 (O_814,N_19302,N_16295);
nand UO_815 (O_815,N_15716,N_15810);
and UO_816 (O_816,N_16686,N_15454);
and UO_817 (O_817,N_16547,N_17582);
nor UO_818 (O_818,N_17343,N_18426);
or UO_819 (O_819,N_15648,N_18205);
xnor UO_820 (O_820,N_18379,N_18527);
nand UO_821 (O_821,N_16170,N_17547);
nand UO_822 (O_822,N_18131,N_18633);
nand UO_823 (O_823,N_18515,N_15109);
nor UO_824 (O_824,N_18285,N_18113);
nor UO_825 (O_825,N_19724,N_16950);
nor UO_826 (O_826,N_17916,N_16195);
and UO_827 (O_827,N_18849,N_15910);
nand UO_828 (O_828,N_18227,N_19514);
nor UO_829 (O_829,N_18014,N_19699);
and UO_830 (O_830,N_18715,N_15894);
xnor UO_831 (O_831,N_17827,N_19293);
and UO_832 (O_832,N_19270,N_16841);
and UO_833 (O_833,N_17721,N_16368);
and UO_834 (O_834,N_18256,N_17707);
nand UO_835 (O_835,N_16916,N_15747);
and UO_836 (O_836,N_18787,N_16520);
nor UO_837 (O_837,N_18888,N_15689);
or UO_838 (O_838,N_18037,N_17341);
or UO_839 (O_839,N_16690,N_19898);
nand UO_840 (O_840,N_18510,N_17010);
nand UO_841 (O_841,N_16834,N_17880);
and UO_842 (O_842,N_19734,N_18337);
xor UO_843 (O_843,N_19016,N_18183);
and UO_844 (O_844,N_15634,N_16324);
and UO_845 (O_845,N_19406,N_18647);
nor UO_846 (O_846,N_15764,N_19333);
nand UO_847 (O_847,N_17111,N_19149);
nor UO_848 (O_848,N_16231,N_16162);
or UO_849 (O_849,N_18381,N_17226);
xnor UO_850 (O_850,N_15602,N_19427);
nand UO_851 (O_851,N_15609,N_19919);
nor UO_852 (O_852,N_17796,N_16063);
and UO_853 (O_853,N_19392,N_16908);
nor UO_854 (O_854,N_15820,N_16806);
xnor UO_855 (O_855,N_17045,N_17578);
nand UO_856 (O_856,N_15178,N_18180);
or UO_857 (O_857,N_18410,N_16802);
or UO_858 (O_858,N_16899,N_18990);
and UO_859 (O_859,N_17493,N_16735);
or UO_860 (O_860,N_16932,N_16012);
xnor UO_861 (O_861,N_15452,N_18937);
nor UO_862 (O_862,N_17698,N_19478);
nor UO_863 (O_863,N_19078,N_16881);
and UO_864 (O_864,N_15627,N_17644);
nand UO_865 (O_865,N_17861,N_15001);
nor UO_866 (O_866,N_16970,N_15135);
or UO_867 (O_867,N_19743,N_18604);
or UO_868 (O_868,N_16554,N_18842);
nand UO_869 (O_869,N_17290,N_16883);
nand UO_870 (O_870,N_17611,N_19952);
nor UO_871 (O_871,N_18999,N_15580);
nand UO_872 (O_872,N_18251,N_19617);
or UO_873 (O_873,N_15308,N_18271);
nand UO_874 (O_874,N_19921,N_18214);
nand UO_875 (O_875,N_19912,N_15443);
nor UO_876 (O_876,N_17151,N_15387);
or UO_877 (O_877,N_16574,N_16102);
or UO_878 (O_878,N_17653,N_15837);
nand UO_879 (O_879,N_18710,N_19202);
nor UO_880 (O_880,N_16696,N_16238);
nand UO_881 (O_881,N_15783,N_15815);
and UO_882 (O_882,N_17978,N_16817);
nor UO_883 (O_883,N_16203,N_15687);
and UO_884 (O_884,N_18070,N_15975);
nor UO_885 (O_885,N_19154,N_19429);
nand UO_886 (O_886,N_15791,N_19223);
and UO_887 (O_887,N_15205,N_16091);
and UO_888 (O_888,N_18653,N_16832);
or UO_889 (O_889,N_15540,N_18973);
nand UO_890 (O_890,N_18350,N_19882);
or UO_891 (O_891,N_16922,N_16706);
or UO_892 (O_892,N_19823,N_15167);
and UO_893 (O_893,N_19866,N_15702);
nand UO_894 (O_894,N_17025,N_16036);
nor UO_895 (O_895,N_16942,N_19098);
or UO_896 (O_896,N_18991,N_17967);
or UO_897 (O_897,N_19629,N_17584);
nor UO_898 (O_898,N_16221,N_16194);
and UO_899 (O_899,N_19220,N_16330);
or UO_900 (O_900,N_15535,N_18857);
nand UO_901 (O_901,N_18608,N_16536);
nor UO_902 (O_902,N_17750,N_18861);
xor UO_903 (O_903,N_18469,N_17839);
or UO_904 (O_904,N_16771,N_19834);
and UO_905 (O_905,N_15720,N_16315);
nand UO_906 (O_906,N_18732,N_16955);
nand UO_907 (O_907,N_18018,N_16676);
or UO_908 (O_908,N_16535,N_19063);
or UO_909 (O_909,N_19201,N_16567);
nand UO_910 (O_910,N_16862,N_15960);
nor UO_911 (O_911,N_19386,N_18616);
and UO_912 (O_912,N_18221,N_16133);
or UO_913 (O_913,N_18525,N_16797);
nor UO_914 (O_914,N_19615,N_19963);
nand UO_915 (O_915,N_16976,N_18114);
and UO_916 (O_916,N_17116,N_15959);
nand UO_917 (O_917,N_18048,N_15547);
or UO_918 (O_918,N_19676,N_18717);
xnor UO_919 (O_919,N_15074,N_16235);
nand UO_920 (O_920,N_16858,N_19012);
nand UO_921 (O_921,N_17988,N_15045);
nand UO_922 (O_922,N_15691,N_15076);
xor UO_923 (O_923,N_15180,N_17455);
nor UO_924 (O_924,N_17337,N_16267);
and UO_925 (O_925,N_19191,N_15751);
xnor UO_926 (O_926,N_19389,N_18581);
xor UO_927 (O_927,N_17119,N_19973);
nand UO_928 (O_928,N_15505,N_19696);
nor UO_929 (O_929,N_19236,N_16675);
nand UO_930 (O_930,N_15857,N_17642);
and UO_931 (O_931,N_16935,N_18324);
or UO_932 (O_932,N_19327,N_19465);
nor UO_933 (O_933,N_15220,N_17776);
and UO_934 (O_934,N_18055,N_17955);
or UO_935 (O_935,N_16891,N_16727);
nand UO_936 (O_936,N_18144,N_15713);
xnor UO_937 (O_937,N_18847,N_19265);
nand UO_938 (O_938,N_19013,N_18222);
and UO_939 (O_939,N_19934,N_19535);
and UO_940 (O_940,N_18275,N_19574);
and UO_941 (O_941,N_15159,N_16045);
nor UO_942 (O_942,N_18866,N_16725);
nor UO_943 (O_943,N_15450,N_17530);
nand UO_944 (O_944,N_17453,N_15496);
xor UO_945 (O_945,N_19002,N_17557);
or UO_946 (O_946,N_16704,N_18720);
and UO_947 (O_947,N_16888,N_15012);
and UO_948 (O_948,N_16989,N_16510);
and UO_949 (O_949,N_19077,N_18177);
nor UO_950 (O_950,N_15945,N_19606);
and UO_951 (O_951,N_16646,N_19965);
and UO_952 (O_952,N_16639,N_19946);
xor UO_953 (O_953,N_16544,N_16722);
or UO_954 (O_954,N_18334,N_16564);
nor UO_955 (O_955,N_18932,N_19767);
and UO_956 (O_956,N_19407,N_15161);
and UO_957 (O_957,N_16069,N_18237);
or UO_958 (O_958,N_17514,N_19352);
and UO_959 (O_959,N_15523,N_19029);
and UO_960 (O_960,N_15651,N_17599);
and UO_961 (O_961,N_16893,N_17224);
and UO_962 (O_962,N_18742,N_17495);
nand UO_963 (O_963,N_19680,N_17117);
and UO_964 (O_964,N_19820,N_17779);
or UO_965 (O_965,N_19761,N_17082);
nor UO_966 (O_966,N_15303,N_17817);
and UO_967 (O_967,N_16694,N_17883);
nand UO_968 (O_968,N_17959,N_16008);
and UO_969 (O_969,N_18136,N_18452);
nand UO_970 (O_970,N_15060,N_15845);
or UO_971 (O_971,N_17550,N_18536);
or UO_972 (O_972,N_18360,N_17346);
xor UO_973 (O_973,N_15972,N_15213);
nor UO_974 (O_974,N_17729,N_19788);
and UO_975 (O_975,N_19519,N_18557);
nand UO_976 (O_976,N_18129,N_17541);
and UO_977 (O_977,N_17372,N_17049);
xor UO_978 (O_978,N_19937,N_16527);
or UO_979 (O_979,N_15918,N_17619);
nand UO_980 (O_980,N_16081,N_19893);
and UO_981 (O_981,N_18433,N_15459);
nand UO_982 (O_982,N_17832,N_16118);
and UO_983 (O_983,N_18607,N_19033);
and UO_984 (O_984,N_16411,N_15868);
nor UO_985 (O_985,N_16509,N_19738);
or UO_986 (O_986,N_15879,N_17285);
or UO_987 (O_987,N_15374,N_18730);
or UO_988 (O_988,N_15767,N_15063);
nor UO_989 (O_989,N_17124,N_19290);
nand UO_990 (O_990,N_17208,N_17016);
xor UO_991 (O_991,N_16904,N_19237);
or UO_992 (O_992,N_16958,N_17245);
xor UO_993 (O_993,N_19964,N_19684);
and UO_994 (O_994,N_15337,N_17080);
and UO_995 (O_995,N_16327,N_17938);
and UO_996 (O_996,N_19901,N_16702);
nor UO_997 (O_997,N_18564,N_15555);
xnor UO_998 (O_998,N_19312,N_15865);
nor UO_999 (O_999,N_16999,N_18503);
nor UO_1000 (O_1000,N_19801,N_15641);
nand UO_1001 (O_1001,N_16608,N_17338);
nand UO_1002 (O_1002,N_17974,N_15408);
nand UO_1003 (O_1003,N_15117,N_15465);
and UO_1004 (O_1004,N_16764,N_19972);
nor UO_1005 (O_1005,N_15099,N_16467);
nand UO_1006 (O_1006,N_17053,N_16598);
nor UO_1007 (O_1007,N_16644,N_19297);
nand UO_1008 (O_1008,N_17219,N_19147);
nand UO_1009 (O_1009,N_16401,N_16137);
or UO_1010 (O_1010,N_15690,N_15866);
or UO_1011 (O_1011,N_17298,N_19438);
and UO_1012 (O_1012,N_15973,N_18892);
nor UO_1013 (O_1013,N_17336,N_16212);
and UO_1014 (O_1014,N_16396,N_18600);
and UO_1015 (O_1015,N_15036,N_17917);
and UO_1016 (O_1016,N_15083,N_16933);
nand UO_1017 (O_1017,N_17169,N_19273);
nand UO_1018 (O_1018,N_15243,N_16066);
nand UO_1019 (O_1019,N_18851,N_18146);
and UO_1020 (O_1020,N_19301,N_19797);
or UO_1021 (O_1021,N_18108,N_18153);
and UO_1022 (O_1022,N_15137,N_16135);
nand UO_1023 (O_1023,N_17754,N_19131);
nor UO_1024 (O_1024,N_18884,N_18021);
and UO_1025 (O_1025,N_18282,N_18487);
nor UO_1026 (O_1026,N_17849,N_18876);
nor UO_1027 (O_1027,N_17663,N_18881);
and UO_1028 (O_1028,N_16974,N_15771);
nand UO_1029 (O_1029,N_17060,N_18528);
or UO_1030 (O_1030,N_16130,N_16390);
and UO_1031 (O_1031,N_19861,N_15701);
xor UO_1032 (O_1032,N_19133,N_17328);
xnor UO_1033 (O_1033,N_19553,N_15168);
or UO_1034 (O_1034,N_17546,N_17743);
nor UO_1035 (O_1035,N_18848,N_17601);
and UO_1036 (O_1036,N_17968,N_18489);
and UO_1037 (O_1037,N_16157,N_19691);
nand UO_1038 (O_1038,N_19416,N_17545);
nor UO_1039 (O_1039,N_15552,N_19388);
xnor UO_1040 (O_1040,N_16108,N_19310);
xor UO_1041 (O_1041,N_16208,N_18955);
and UO_1042 (O_1042,N_15457,N_16159);
and UO_1043 (O_1043,N_15472,N_19198);
and UO_1044 (O_1044,N_15366,N_15839);
nand UO_1045 (O_1045,N_15093,N_19899);
nand UO_1046 (O_1046,N_18374,N_16821);
and UO_1047 (O_1047,N_16270,N_19812);
xnor UO_1048 (O_1048,N_16441,N_19228);
and UO_1049 (O_1049,N_16156,N_18830);
or UO_1050 (O_1050,N_17389,N_15901);
or UO_1051 (O_1051,N_17609,N_17388);
and UO_1052 (O_1052,N_18533,N_17842);
nand UO_1053 (O_1053,N_19330,N_17163);
nand UO_1054 (O_1054,N_17595,N_19759);
nand UO_1055 (O_1055,N_17515,N_17985);
nand UO_1056 (O_1056,N_19028,N_16625);
nand UO_1057 (O_1057,N_19493,N_19249);
or UO_1058 (O_1058,N_19363,N_19255);
nor UO_1059 (O_1059,N_19168,N_16475);
xnor UO_1060 (O_1060,N_18137,N_19733);
nand UO_1061 (O_1061,N_19777,N_16121);
nand UO_1062 (O_1062,N_16092,N_17078);
nand UO_1063 (O_1063,N_16200,N_15789);
nor UO_1064 (O_1064,N_18327,N_18193);
nand UO_1065 (O_1065,N_17508,N_15852);
nand UO_1066 (O_1066,N_17103,N_18078);
or UO_1067 (O_1067,N_16937,N_18502);
or UO_1068 (O_1068,N_15595,N_19136);
or UO_1069 (O_1069,N_15248,N_16844);
nand UO_1070 (O_1070,N_17432,N_15728);
or UO_1071 (O_1071,N_18303,N_16397);
xnor UO_1072 (O_1072,N_17254,N_18675);
nand UO_1073 (O_1073,N_19103,N_17350);
and UO_1074 (O_1074,N_17928,N_18073);
nor UO_1075 (O_1075,N_17556,N_19712);
and UO_1076 (O_1076,N_16191,N_18788);
nand UO_1077 (O_1077,N_15804,N_18168);
nor UO_1078 (O_1078,N_15396,N_19827);
xor UO_1079 (O_1079,N_17020,N_19055);
nor UO_1080 (O_1080,N_18158,N_15581);
or UO_1081 (O_1081,N_19537,N_19505);
nor UO_1082 (O_1082,N_15413,N_18570);
nand UO_1083 (O_1083,N_19319,N_19543);
nor UO_1084 (O_1084,N_15438,N_17217);
nand UO_1085 (O_1085,N_15782,N_16929);
or UO_1086 (O_1086,N_17267,N_18927);
nor UO_1087 (O_1087,N_15021,N_19367);
or UO_1088 (O_1088,N_17067,N_18124);
and UO_1089 (O_1089,N_18025,N_18885);
nor UO_1090 (O_1090,N_15160,N_15091);
xor UO_1091 (O_1091,N_16489,N_17991);
or UO_1092 (O_1092,N_15499,N_17867);
nor UO_1093 (O_1093,N_17963,N_17590);
nand UO_1094 (O_1094,N_19437,N_15605);
and UO_1095 (O_1095,N_16001,N_17357);
or UO_1096 (O_1096,N_16631,N_16498);
or UO_1097 (O_1097,N_16572,N_19643);
nand UO_1098 (O_1098,N_15624,N_17915);
nand UO_1099 (O_1099,N_16256,N_18549);
nand UO_1100 (O_1100,N_15882,N_19532);
and UO_1101 (O_1101,N_15474,N_16665);
and UO_1102 (O_1102,N_16466,N_16709);
nand UO_1103 (O_1103,N_18682,N_17947);
and UO_1104 (O_1104,N_18877,N_19980);
or UO_1105 (O_1105,N_18434,N_19626);
xor UO_1106 (O_1106,N_15819,N_18532);
and UO_1107 (O_1107,N_19048,N_15576);
nand UO_1108 (O_1108,N_16503,N_17315);
and UO_1109 (O_1109,N_19127,N_15427);
nor UO_1110 (O_1110,N_17787,N_17511);
xnor UO_1111 (O_1111,N_17188,N_15997);
xor UO_1112 (O_1112,N_19675,N_18958);
and UO_1113 (O_1113,N_17486,N_16634);
and UO_1114 (O_1114,N_15906,N_18049);
or UO_1115 (O_1115,N_17674,N_15729);
or UO_1116 (O_1116,N_19239,N_19523);
nor UO_1117 (O_1117,N_18157,N_19857);
and UO_1118 (O_1118,N_15377,N_17522);
xnor UO_1119 (O_1119,N_19648,N_18498);
nor UO_1120 (O_1120,N_19879,N_17123);
nor UO_1121 (O_1121,N_19754,N_18891);
nor UO_1122 (O_1122,N_15011,N_15794);
or UO_1123 (O_1123,N_19024,N_19845);
and UO_1124 (O_1124,N_18996,N_17327);
nor UO_1125 (O_1125,N_18488,N_15201);
nand UO_1126 (O_1126,N_16459,N_17331);
nor UO_1127 (O_1127,N_19025,N_18287);
nor UO_1128 (O_1128,N_19594,N_16524);
and UO_1129 (O_1129,N_15052,N_19107);
or UO_1130 (O_1130,N_15520,N_19234);
and UO_1131 (O_1131,N_19181,N_17132);
or UO_1132 (O_1132,N_19766,N_18566);
and UO_1133 (O_1133,N_15982,N_18746);
or UO_1134 (O_1134,N_17419,N_15860);
nor UO_1135 (O_1135,N_18854,N_19548);
nand UO_1136 (O_1136,N_16626,N_18917);
and UO_1137 (O_1137,N_19650,N_18463);
nor UO_1138 (O_1138,N_15914,N_18030);
xor UO_1139 (O_1139,N_16126,N_15867);
and UO_1140 (O_1140,N_19950,N_18872);
nand UO_1141 (O_1141,N_15694,N_19433);
and UO_1142 (O_1142,N_18979,N_17881);
nand UO_1143 (O_1143,N_19112,N_15362);
or UO_1144 (O_1144,N_18947,N_18273);
nand UO_1145 (O_1145,N_18388,N_17592);
and UO_1146 (O_1146,N_17294,N_15345);
and UO_1147 (O_1147,N_18202,N_15126);
xnor UO_1148 (O_1148,N_19683,N_16219);
nand UO_1149 (O_1149,N_16164,N_19842);
nand UO_1150 (O_1150,N_19269,N_19057);
or UO_1151 (O_1151,N_18455,N_15629);
xor UO_1152 (O_1152,N_15872,N_15946);
or UO_1153 (O_1153,N_16575,N_15781);
nor UO_1154 (O_1154,N_17618,N_15958);
and UO_1155 (O_1155,N_15445,N_19917);
and UO_1156 (O_1156,N_16724,N_19457);
nor UO_1157 (O_1157,N_17631,N_19757);
and UO_1158 (O_1158,N_15678,N_17686);
nor UO_1159 (O_1159,N_18011,N_17814);
or UO_1160 (O_1160,N_18229,N_15293);
nand UO_1161 (O_1161,N_15493,N_16673);
nor UO_1162 (O_1162,N_16375,N_18507);
or UO_1163 (O_1163,N_19150,N_19174);
or UO_1164 (O_1164,N_19704,N_16822);
or UO_1165 (O_1165,N_15463,N_16930);
or UO_1166 (O_1166,N_15635,N_18882);
nor UO_1167 (O_1167,N_16128,N_19677);
or UO_1168 (O_1168,N_16456,N_18297);
and UO_1169 (O_1169,N_18640,N_19336);
and UO_1170 (O_1170,N_15273,N_15477);
xor UO_1171 (O_1171,N_15291,N_17277);
or UO_1172 (O_1172,N_19041,N_18899);
and UO_1173 (O_1173,N_15492,N_19471);
xnor UO_1174 (O_1174,N_17635,N_16848);
xnor UO_1175 (O_1175,N_15683,N_19998);
nand UO_1176 (O_1176,N_19507,N_17979);
and UO_1177 (O_1177,N_15993,N_16113);
or UO_1178 (O_1178,N_16389,N_18919);
and UO_1179 (O_1179,N_17122,N_17529);
or UO_1180 (O_1180,N_17711,N_18737);
nor UO_1181 (O_1181,N_18261,N_19542);
and UO_1182 (O_1182,N_15584,N_15059);
or UO_1183 (O_1183,N_15980,N_16024);
nand UO_1184 (O_1184,N_18176,N_16089);
and UO_1185 (O_1185,N_18985,N_19613);
or UO_1186 (O_1186,N_16461,N_15738);
and UO_1187 (O_1187,N_16109,N_17084);
or UO_1188 (O_1188,N_16179,N_17767);
and UO_1189 (O_1189,N_19971,N_16148);
or UO_1190 (O_1190,N_17075,N_16541);
nor UO_1191 (O_1191,N_17731,N_16655);
or UO_1192 (O_1192,N_16284,N_16479);
and UO_1193 (O_1193,N_17434,N_17951);
xnor UO_1194 (O_1194,N_19771,N_15242);
or UO_1195 (O_1195,N_17771,N_18829);
nor UO_1196 (O_1196,N_18398,N_19304);
and UO_1197 (O_1197,N_19568,N_17809);
or UO_1198 (O_1198,N_19996,N_17633);
or UO_1199 (O_1199,N_18673,N_16609);
nand UO_1200 (O_1200,N_15570,N_17983);
and UO_1201 (O_1201,N_18841,N_15618);
nor UO_1202 (O_1202,N_19317,N_16300);
or UO_1203 (O_1203,N_15934,N_17236);
or UO_1204 (O_1204,N_17481,N_15992);
and UO_1205 (O_1205,N_18546,N_18332);
or UO_1206 (O_1206,N_17127,N_19546);
or UO_1207 (O_1207,N_16365,N_17352);
or UO_1208 (O_1208,N_16928,N_15352);
or UO_1209 (O_1209,N_18314,N_15361);
and UO_1210 (O_1210,N_17376,N_15632);
nor UO_1211 (O_1211,N_17325,N_15186);
and UO_1212 (O_1212,N_15841,N_17805);
and UO_1213 (O_1213,N_18242,N_17616);
nor UO_1214 (O_1214,N_17202,N_18855);
and UO_1215 (O_1215,N_18695,N_19657);
nor UO_1216 (O_1216,N_17387,N_19485);
nor UO_1217 (O_1217,N_18281,N_18461);
nand UO_1218 (O_1218,N_18953,N_18818);
and UO_1219 (O_1219,N_19095,N_17373);
and UO_1220 (O_1220,N_19609,N_16782);
nor UO_1221 (O_1221,N_17885,N_15371);
or UO_1222 (O_1222,N_15800,N_17382);
or UO_1223 (O_1223,N_16444,N_15665);
nand UO_1224 (O_1224,N_17106,N_15292);
nor UO_1225 (O_1225,N_18863,N_17032);
nand UO_1226 (O_1226,N_18940,N_18718);
and UO_1227 (O_1227,N_19068,N_15840);
or UO_1228 (O_1228,N_16906,N_17975);
or UO_1229 (O_1229,N_17807,N_16783);
or UO_1230 (O_1230,N_15386,N_19583);
or UO_1231 (O_1231,N_18938,N_17566);
nor UO_1232 (O_1232,N_18318,N_19737);
nand UO_1233 (O_1233,N_17066,N_17690);
xnor UO_1234 (O_1234,N_17094,N_16512);
nand UO_1235 (O_1235,N_15929,N_17533);
nor UO_1236 (O_1236,N_19567,N_15599);
or UO_1237 (O_1237,N_16206,N_17506);
nand UO_1238 (O_1238,N_16534,N_16292);
nor UO_1239 (O_1239,N_15933,N_17710);
and UO_1240 (O_1240,N_17517,N_16995);
or UO_1241 (O_1241,N_18439,N_19282);
nand UO_1242 (O_1242,N_15434,N_16860);
nor UO_1243 (O_1243,N_15078,N_18138);
xnor UO_1244 (O_1244,N_17651,N_17848);
nand UO_1245 (O_1245,N_19137,N_16692);
nor UO_1246 (O_1246,N_18982,N_18104);
or UO_1247 (O_1247,N_15922,N_18328);
nand UO_1248 (O_1248,N_16004,N_15393);
nor UO_1249 (O_1249,N_15564,N_17003);
nor UO_1250 (O_1250,N_16913,N_15217);
xor UO_1251 (O_1251,N_18677,N_16345);
or UO_1252 (O_1252,N_19186,N_19747);
or UO_1253 (O_1253,N_15639,N_17143);
and UO_1254 (O_1254,N_18252,N_19685);
or UO_1255 (O_1255,N_18084,N_19539);
nor UO_1256 (O_1256,N_17695,N_15356);
or UO_1257 (O_1257,N_16006,N_18046);
and UO_1258 (O_1258,N_19914,N_15405);
and UO_1259 (O_1259,N_16683,N_15282);
or UO_1260 (O_1260,N_16154,N_15513);
nor UO_1261 (O_1261,N_17172,N_18776);
and UO_1262 (O_1262,N_17195,N_18506);
xor UO_1263 (O_1263,N_16847,N_18791);
nor UO_1264 (O_1264,N_16490,N_17265);
and UO_1265 (O_1265,N_19982,N_17935);
and UO_1266 (O_1266,N_19993,N_17621);
nor UO_1267 (O_1267,N_15324,N_19904);
nand UO_1268 (O_1268,N_16938,N_15502);
or UO_1269 (O_1269,N_17047,N_16607);
xnor UO_1270 (O_1270,N_16237,N_19064);
and UO_1271 (O_1271,N_17176,N_19852);
or UO_1272 (O_1272,N_18819,N_18493);
xnor UO_1273 (O_1273,N_19153,N_19480);
nand UO_1274 (O_1274,N_17312,N_18475);
nor UO_1275 (O_1275,N_17724,N_18119);
xnor UO_1276 (O_1276,N_17220,N_15338);
and UO_1277 (O_1277,N_17131,N_19050);
or UO_1278 (O_1278,N_15256,N_15416);
nor UO_1279 (O_1279,N_19522,N_17852);
and UO_1280 (O_1280,N_15560,N_18135);
nand UO_1281 (O_1281,N_15284,N_16240);
nand UO_1282 (O_1282,N_16166,N_15334);
or UO_1283 (O_1283,N_15669,N_19296);
and UO_1284 (O_1284,N_18562,N_19920);
or UO_1285 (O_1285,N_15192,N_19248);
nor UO_1286 (O_1286,N_17945,N_16484);
or UO_1287 (O_1287,N_16071,N_16317);
nor UO_1288 (O_1288,N_19199,N_15378);
xor UO_1289 (O_1289,N_17789,N_17488);
nand UO_1290 (O_1290,N_15529,N_17027);
or UO_1291 (O_1291,N_18413,N_18072);
nand UO_1292 (O_1292,N_19288,N_16035);
and UO_1293 (O_1293,N_15196,N_17872);
and UO_1294 (O_1294,N_18155,N_18547);
nor UO_1295 (O_1295,N_18959,N_15525);
nand UO_1296 (O_1296,N_18449,N_16677);
or UO_1297 (O_1297,N_15421,N_17823);
nand UO_1298 (O_1298,N_17399,N_19647);
and UO_1299 (O_1299,N_15824,N_15173);
nor UO_1300 (O_1300,N_15796,N_17002);
and UO_1301 (O_1301,N_18182,N_19124);
or UO_1302 (O_1302,N_16055,N_17252);
xnor UO_1303 (O_1303,N_18544,N_16621);
or UO_1304 (O_1304,N_19774,N_15006);
or UO_1305 (O_1305,N_18172,N_18143);
nor UO_1306 (O_1306,N_19593,N_15422);
nor UO_1307 (O_1307,N_18722,N_17833);
nand UO_1308 (O_1308,N_16762,N_15770);
or UO_1309 (O_1309,N_19326,N_18820);
and UO_1310 (O_1310,N_19925,N_16282);
or UO_1311 (O_1311,N_18076,N_16242);
nand UO_1312 (O_1312,N_17869,N_15623);
or UO_1313 (O_1313,N_19281,N_16760);
and UO_1314 (O_1314,N_15071,N_18300);
xnor UO_1315 (O_1315,N_15381,N_16887);
nor UO_1316 (O_1316,N_16911,N_18921);
and UO_1317 (O_1317,N_15984,N_19432);
nand UO_1318 (O_1318,N_15152,N_15532);
and UO_1319 (O_1319,N_19814,N_18716);
or UO_1320 (O_1320,N_18724,N_15176);
xnor UO_1321 (O_1321,N_16552,N_17408);
nor UO_1322 (O_1322,N_17919,N_19730);
nand UO_1323 (O_1323,N_18799,N_19560);
or UO_1324 (O_1324,N_17168,N_18423);
nor UO_1325 (O_1325,N_16642,N_17190);
or UO_1326 (O_1326,N_17360,N_17139);
xnor UO_1327 (O_1327,N_17034,N_17662);
nor UO_1328 (O_1328,N_15401,N_17333);
nor UO_1329 (O_1329,N_15801,N_16488);
and UO_1330 (O_1330,N_17430,N_15114);
nor UO_1331 (O_1331,N_16643,N_16545);
or UO_1332 (O_1332,N_16508,N_16828);
nor UO_1333 (O_1333,N_15423,N_17540);
or UO_1334 (O_1334,N_15067,N_19384);
and UO_1335 (O_1335,N_17855,N_17281);
nor UO_1336 (O_1336,N_17483,N_17061);
and UO_1337 (O_1337,N_17813,N_16332);
nor UO_1338 (O_1338,N_19618,N_15711);
nand UO_1339 (O_1339,N_16061,N_15195);
or UO_1340 (O_1340,N_15008,N_16460);
nand UO_1341 (O_1341,N_17672,N_16483);
nand UO_1342 (O_1342,N_16002,N_17098);
or UO_1343 (O_1343,N_15777,N_15333);
nor UO_1344 (O_1344,N_15288,N_18995);
nor UO_1345 (O_1345,N_16142,N_16040);
or UO_1346 (O_1346,N_19101,N_15392);
nand UO_1347 (O_1347,N_16915,N_18784);
and UO_1348 (O_1348,N_19984,N_19661);
or UO_1349 (O_1349,N_18588,N_19451);
xor UO_1350 (O_1350,N_16129,N_19072);
nor UO_1351 (O_1351,N_17185,N_17001);
or UO_1352 (O_1352,N_16606,N_18464);
nand UO_1353 (O_1353,N_15663,N_18127);
and UO_1354 (O_1354,N_19992,N_16969);
nor UO_1355 (O_1355,N_18371,N_17450);
or UO_1356 (O_1356,N_19708,N_19679);
or UO_1357 (O_1357,N_16244,N_16743);
or UO_1358 (O_1358,N_18061,N_16038);
and UO_1359 (O_1359,N_16181,N_16687);
xnor UO_1360 (O_1360,N_18949,N_16604);
nand UO_1361 (O_1361,N_18538,N_16550);
and UO_1362 (O_1362,N_17949,N_18340);
nand UO_1363 (O_1363,N_17490,N_17791);
and UO_1364 (O_1364,N_16233,N_16507);
or UO_1365 (O_1365,N_16442,N_16565);
nor UO_1366 (O_1366,N_19413,N_18584);
nor UO_1367 (O_1367,N_16738,N_15367);
nand UO_1368 (O_1368,N_19628,N_17283);
nand UO_1369 (O_1369,N_19351,N_16861);
nor UO_1370 (O_1370,N_16372,N_19625);
nor UO_1371 (O_1371,N_18223,N_16043);
or UO_1372 (O_1372,N_17661,N_19672);
nand UO_1373 (O_1373,N_17378,N_18097);
nand UO_1374 (O_1374,N_15127,N_17223);
or UO_1375 (O_1375,N_15874,N_19941);
nor UO_1376 (O_1376,N_16318,N_15995);
and UO_1377 (O_1377,N_16413,N_17732);
and UO_1378 (O_1378,N_17868,N_16030);
nand UO_1379 (O_1379,N_18035,N_16791);
nand UO_1380 (O_1380,N_17412,N_16927);
nor UO_1381 (O_1381,N_19090,N_19175);
nand UO_1382 (O_1382,N_17377,N_19238);
and UO_1383 (O_1383,N_15859,N_19263);
nor UO_1384 (O_1384,N_15630,N_17894);
and UO_1385 (O_1385,N_19377,N_15451);
and UO_1386 (O_1386,N_18587,N_15444);
nand UO_1387 (O_1387,N_16248,N_18109);
nand UO_1388 (O_1388,N_15447,N_17028);
nor UO_1389 (O_1389,N_19331,N_17092);
nor UO_1390 (O_1390,N_15566,N_16239);
or UO_1391 (O_1391,N_19645,N_19720);
nand UO_1392 (O_1392,N_19632,N_16362);
and UO_1393 (O_1393,N_15049,N_17922);
and UO_1394 (O_1394,N_19776,N_18905);
and UO_1395 (O_1395,N_19117,N_15120);
nand UO_1396 (O_1396,N_18630,N_16046);
or UO_1397 (O_1397,N_15917,N_17657);
nand UO_1398 (O_1398,N_18516,N_18934);
xnor UO_1399 (O_1399,N_15111,N_16391);
nand UO_1400 (O_1400,N_15069,N_16638);
xnor UO_1401 (O_1401,N_17206,N_15164);
nand UO_1402 (O_1402,N_17884,N_15697);
and UO_1403 (O_1403,N_18626,N_16982);
or UO_1404 (O_1404,N_16855,N_18524);
or UO_1405 (O_1405,N_18051,N_19402);
nand UO_1406 (O_1406,N_18740,N_17087);
xnor UO_1407 (O_1407,N_15301,N_16610);
xor UO_1408 (O_1408,N_16319,N_15429);
nor UO_1409 (O_1409,N_16654,N_18427);
nor UO_1410 (O_1410,N_17437,N_19871);
and UO_1411 (O_1411,N_18731,N_19639);
and UO_1412 (O_1412,N_18198,N_16260);
nand UO_1413 (O_1413,N_18939,N_15084);
nor UO_1414 (O_1414,N_17568,N_19313);
or UO_1415 (O_1415,N_18117,N_18020);
or UO_1416 (O_1416,N_15577,N_18201);
nor UO_1417 (O_1417,N_19781,N_18856);
xor UO_1418 (O_1418,N_17931,N_16299);
and UO_1419 (O_1419,N_19986,N_17722);
or UO_1420 (O_1420,N_19655,N_18368);
or UO_1421 (O_1421,N_18042,N_16872);
and UO_1422 (O_1422,N_16312,N_17261);
nor UO_1423 (O_1423,N_19089,N_17356);
nor UO_1424 (O_1424,N_18391,N_15768);
nand UO_1425 (O_1425,N_17523,N_16588);
xnor UO_1426 (O_1426,N_19410,N_16876);
nor UO_1427 (O_1427,N_15261,N_16272);
or UO_1428 (O_1428,N_19841,N_17700);
and UO_1429 (O_1429,N_15558,N_18186);
nor UO_1430 (O_1430,N_15559,N_16491);
nand UO_1431 (O_1431,N_15272,N_18727);
nor UO_1432 (O_1432,N_17891,N_19378);
nor UO_1433 (O_1433,N_19916,N_15943);
or UO_1434 (O_1434,N_17292,N_18291);
and UO_1435 (O_1435,N_16818,N_19375);
nand UO_1436 (O_1436,N_15688,N_17401);
xor UO_1437 (O_1437,N_17021,N_15141);
nand UO_1438 (O_1438,N_15885,N_19260);
or UO_1439 (O_1439,N_19037,N_15479);
or UO_1440 (O_1440,N_19520,N_16581);
nor UO_1441 (O_1441,N_16048,N_18691);
nor UO_1442 (O_1442,N_17504,N_19258);
or UO_1443 (O_1443,N_15843,N_18376);
nand UO_1444 (O_1444,N_16297,N_15753);
or UO_1445 (O_1445,N_15403,N_16323);
xor UO_1446 (O_1446,N_18415,N_15913);
xor UO_1447 (O_1447,N_19939,N_19611);
nor UO_1448 (O_1448,N_17183,N_18121);
nand UO_1449 (O_1449,N_18369,N_19096);
nand UO_1450 (O_1450,N_19896,N_15740);
or UO_1451 (O_1451,N_18623,N_18632);
nor UO_1452 (O_1452,N_18531,N_17673);
or UO_1453 (O_1453,N_17755,N_16377);
and UO_1454 (O_1454,N_15395,N_16015);
nand UO_1455 (O_1455,N_15680,N_15467);
or UO_1456 (O_1456,N_17006,N_19152);
nand UO_1457 (O_1457,N_19764,N_17110);
nor UO_1458 (O_1458,N_18648,N_18474);
nor UO_1459 (O_1459,N_15548,N_17273);
or UO_1460 (O_1460,N_15612,N_17459);
or UO_1461 (O_1461,N_19356,N_17944);
and UO_1462 (O_1462,N_19803,N_15658);
or UO_1463 (O_1463,N_17189,N_17569);
or UO_1464 (O_1464,N_15296,N_17939);
and UO_1465 (O_1465,N_17583,N_15977);
xnor UO_1466 (O_1466,N_19455,N_18897);
and UO_1467 (O_1467,N_16628,N_19811);
nand UO_1468 (O_1468,N_15061,N_19585);
nand UO_1469 (O_1469,N_15009,N_18033);
or UO_1470 (O_1470,N_19271,N_17344);
xor UO_1471 (O_1471,N_18425,N_17570);
or UO_1472 (O_1472,N_19718,N_16546);
xor UO_1473 (O_1473,N_18192,N_18188);
or UO_1474 (O_1474,N_17182,N_16342);
nor UO_1475 (O_1475,N_16632,N_17835);
and UO_1476 (O_1476,N_15347,N_15937);
and UO_1477 (O_1477,N_18500,N_17645);
xnor UO_1478 (O_1478,N_17640,N_15480);
nor UO_1479 (O_1479,N_18122,N_15511);
nor UO_1480 (O_1480,N_19909,N_19441);
nor UO_1481 (O_1481,N_18149,N_16234);
nor UO_1482 (O_1482,N_17299,N_16750);
nand UO_1483 (O_1483,N_16975,N_19700);
and UO_1484 (O_1484,N_18115,N_18226);
nor UO_1485 (O_1485,N_19944,N_19151);
nand UO_1486 (O_1486,N_16414,N_17589);
nor UO_1487 (O_1487,N_19442,N_18370);
and UO_1488 (O_1488,N_18663,N_17830);
nand UO_1489 (O_1489,N_16978,N_16253);
or UO_1490 (O_1490,N_16325,N_19062);
and UO_1491 (O_1491,N_16316,N_19915);
and UO_1492 (O_1492,N_16427,N_15855);
or UO_1493 (O_1493,N_15965,N_17770);
nand UO_1494 (O_1494,N_18993,N_17543);
or UO_1495 (O_1495,N_17765,N_19337);
nor UO_1496 (O_1496,N_18217,N_19524);
nor UO_1497 (O_1497,N_18926,N_17000);
nand UO_1498 (O_1498,N_17801,N_15355);
nand UO_1499 (O_1499,N_15274,N_16594);
nor UO_1500 (O_1500,N_15437,N_17637);
and UO_1501 (O_1501,N_17199,N_15340);
nand UO_1502 (O_1502,N_16879,N_19143);
xor UO_1503 (O_1503,N_18418,N_15707);
or UO_1504 (O_1504,N_16966,N_16280);
or UO_1505 (O_1505,N_17769,N_19640);
nor UO_1506 (O_1506,N_17426,N_17921);
or UO_1507 (O_1507,N_18367,N_17482);
nand UO_1508 (O_1508,N_18634,N_17184);
or UO_1509 (O_1509,N_19365,N_16761);
and UO_1510 (O_1510,N_16787,N_16218);
nor UO_1511 (O_1511,N_17478,N_16016);
and UO_1512 (O_1512,N_15594,N_17448);
and UO_1513 (O_1513,N_15748,N_15048);
and UO_1514 (O_1514,N_17263,N_18779);
nand UO_1515 (O_1515,N_16236,N_15544);
or UO_1516 (O_1516,N_16905,N_16349);
nand UO_1517 (O_1517,N_19379,N_15175);
nor UO_1518 (O_1518,N_19449,N_19578);
and UO_1519 (O_1519,N_15311,N_15775);
nor UO_1520 (O_1520,N_17909,N_18808);
nand UO_1521 (O_1521,N_15645,N_15880);
nor UO_1522 (O_1522,N_18019,N_18867);
nand UO_1523 (O_1523,N_19510,N_16199);
or UO_1524 (O_1524,N_16815,N_16165);
nand UO_1525 (O_1525,N_17332,N_17304);
and UO_1526 (O_1526,N_18105,N_16617);
nand UO_1527 (O_1527,N_19500,N_16773);
and UO_1528 (O_1528,N_17551,N_19409);
nand UO_1529 (O_1529,N_16054,N_19873);
and UO_1530 (O_1530,N_16468,N_18349);
and UO_1531 (O_1531,N_16605,N_16973);
and UO_1532 (O_1532,N_17697,N_19436);
xnor UO_1533 (O_1533,N_19324,N_18161);
xnor UO_1534 (O_1534,N_18652,N_19390);
or UO_1535 (O_1535,N_17274,N_16305);
and UO_1536 (O_1536,N_18751,N_17234);
nand UO_1537 (O_1537,N_17334,N_15643);
and UO_1538 (O_1538,N_18644,N_18725);
nor UO_1539 (O_1539,N_15142,N_18280);
nor UO_1540 (O_1540,N_18642,N_18028);
or UO_1541 (O_1541,N_16436,N_16513);
xnor UO_1542 (O_1542,N_18047,N_18173);
nor UO_1543 (O_1543,N_17305,N_16355);
xnor UO_1544 (O_1544,N_19435,N_16249);
and UO_1545 (O_1545,N_19017,N_16521);
nor UO_1546 (O_1546,N_19332,N_17977);
and UO_1547 (O_1547,N_18404,N_16334);
nand UO_1548 (O_1548,N_16228,N_19689);
or UO_1549 (O_1549,N_15583,N_15966);
or UO_1550 (O_1550,N_17083,N_19666);
or UO_1551 (O_1551,N_19673,N_15750);
and UO_1552 (O_1552,N_17141,N_17976);
and UO_1553 (O_1553,N_18246,N_18706);
and UO_1554 (O_1554,N_16067,N_17174);
and UO_1555 (O_1555,N_15892,N_16310);
and UO_1556 (O_1556,N_16560,N_18429);
and UO_1557 (O_1557,N_19716,N_19204);
and UO_1558 (O_1558,N_17532,N_16359);
nor UO_1559 (O_1559,N_17684,N_17658);
xor UO_1560 (O_1560,N_16367,N_17271);
or UO_1561 (O_1561,N_19214,N_19978);
or UO_1562 (O_1562,N_18210,N_15899);
nand UO_1563 (O_1563,N_15512,N_15490);
nand UO_1564 (O_1564,N_19722,N_19461);
xnor UO_1565 (O_1565,N_17393,N_17272);
nor UO_1566 (O_1566,N_17097,N_17134);
nor UO_1567 (O_1567,N_17748,N_17857);
or UO_1568 (O_1568,N_15600,N_19232);
nand UO_1569 (O_1569,N_17278,N_16277);
or UO_1570 (O_1570,N_17811,N_15961);
xor UO_1571 (O_1571,N_18428,N_17828);
nor UO_1572 (O_1572,N_15672,N_16410);
xor UO_1573 (O_1573,N_16926,N_16100);
nor UO_1574 (O_1574,N_17146,N_18768);
nor UO_1575 (O_1575,N_17606,N_15174);
nor UO_1576 (O_1576,N_19957,N_16093);
and UO_1577 (O_1577,N_19115,N_17565);
and UO_1578 (O_1578,N_18534,N_16985);
nor UO_1579 (O_1579,N_15568,N_16430);
or UO_1580 (O_1580,N_19573,N_17166);
and UO_1581 (O_1581,N_15212,N_16629);
and UO_1582 (O_1582,N_18295,N_19544);
or UO_1583 (O_1583,N_17753,N_15406);
nand UO_1584 (O_1584,N_18408,N_15670);
and UO_1585 (O_1585,N_19601,N_18619);
nor UO_1586 (O_1586,N_15891,N_19111);
or UO_1587 (O_1587,N_18593,N_16188);
or UO_1588 (O_1588,N_17186,N_18184);
xnor UO_1589 (O_1589,N_16795,N_15849);
and UO_1590 (O_1590,N_15068,N_19216);
xnor UO_1591 (O_1591,N_19221,N_18785);
and UO_1592 (O_1592,N_18254,N_17013);
nor UO_1593 (O_1593,N_17404,N_18800);
nor UO_1594 (O_1594,N_15307,N_18744);
and UO_1595 (O_1595,N_18931,N_15470);
or UO_1596 (O_1596,N_16640,N_17602);
or UO_1597 (O_1597,N_18080,N_16122);
and UO_1598 (O_1598,N_18382,N_15938);
nand UO_1599 (O_1599,N_17677,N_18356);
nor UO_1600 (O_1600,N_18057,N_19369);
or UO_1601 (O_1601,N_17561,N_16247);
nor UO_1602 (O_1602,N_15440,N_15582);
and UO_1603 (O_1603,N_17262,N_15017);
nor UO_1604 (O_1604,N_17354,N_16104);
nand UO_1605 (O_1605,N_15297,N_15032);
or UO_1606 (O_1606,N_16516,N_19619);
xnor UO_1607 (O_1607,N_17364,N_18621);
or UO_1608 (O_1608,N_15696,N_19649);
nor UO_1609 (O_1609,N_19357,N_19576);
xor UO_1610 (O_1610,N_17011,N_17178);
or UO_1611 (O_1611,N_18372,N_16259);
and UO_1612 (O_1612,N_18479,N_19864);
nand UO_1613 (O_1613,N_18393,N_17679);
and UO_1614 (O_1614,N_17231,N_19779);
nor UO_1615 (O_1615,N_16371,N_17646);
and UO_1616 (O_1616,N_17965,N_16562);
xor UO_1617 (O_1617,N_16658,N_15905);
nand UO_1618 (O_1618,N_19697,N_17559);
nor UO_1619 (O_1619,N_16801,N_16615);
and UO_1620 (O_1620,N_17159,N_16171);
nor UO_1621 (O_1621,N_19458,N_15553);
xnor UO_1622 (O_1622,N_17950,N_18870);
or UO_1623 (O_1623,N_17701,N_18477);
nor UO_1624 (O_1624,N_19358,N_15290);
nand UO_1625 (O_1625,N_16224,N_19267);
or UO_1626 (O_1626,N_17268,N_15955);
xnor UO_1627 (O_1627,N_15140,N_17953);
xor UO_1628 (O_1628,N_19646,N_19531);
nand UO_1629 (O_1629,N_18355,N_17042);
nor UO_1630 (O_1630,N_19566,N_18207);
and UO_1631 (O_1631,N_16183,N_17498);
xor UO_1632 (O_1632,N_17948,N_16529);
or UO_1633 (O_1633,N_17836,N_19849);
or UO_1634 (O_1634,N_17349,N_15257);
nand UO_1635 (O_1635,N_19665,N_18599);
nor UO_1636 (O_1636,N_15772,N_19528);
nor UO_1637 (O_1637,N_15353,N_18409);
xnor UO_1638 (O_1638,N_15745,N_18850);
or UO_1639 (O_1639,N_18505,N_15614);
or UO_1640 (O_1640,N_18711,N_17579);
or UO_1641 (O_1641,N_18497,N_17914);
and UO_1642 (O_1642,N_19482,N_17656);
nand UO_1643 (O_1643,N_19431,N_18216);
nand UO_1644 (O_1644,N_18333,N_19854);
and UO_1645 (O_1645,N_18099,N_16961);
nand UO_1646 (O_1646,N_19922,N_17858);
nor UO_1647 (O_1647,N_19831,N_15098);
or UO_1648 (O_1648,N_17295,N_17287);
nor UO_1649 (O_1649,N_19924,N_16814);
and UO_1650 (O_1650,N_16656,N_17802);
or UO_1651 (O_1651,N_19517,N_19800);
nor UO_1652 (O_1652,N_16269,N_15344);
and UO_1653 (O_1653,N_15524,N_18726);
nor UO_1654 (O_1654,N_19513,N_15155);
xor UO_1655 (O_1655,N_18794,N_18798);
or UO_1656 (O_1656,N_17841,N_19044);
and UO_1657 (O_1657,N_18977,N_17720);
or UO_1658 (O_1658,N_15488,N_15737);
nand UO_1659 (O_1659,N_15219,N_17164);
or UO_1660 (O_1660,N_15105,N_19529);
nor UO_1661 (O_1661,N_17102,N_15226);
nor UO_1662 (O_1662,N_19638,N_16757);
or UO_1663 (O_1663,N_16570,N_17456);
and UO_1664 (O_1664,N_16480,N_17696);
nand UO_1665 (O_1665,N_18248,N_18667);
and UO_1666 (O_1666,N_16344,N_15166);
nand UO_1667 (O_1667,N_15424,N_17647);
nor UO_1668 (O_1668,N_18807,N_18994);
nor UO_1669 (O_1669,N_17480,N_18308);
xnor UO_1670 (O_1670,N_17900,N_17411);
nor UO_1671 (O_1671,N_16719,N_18102);
or UO_1672 (O_1672,N_18689,N_19630);
and UO_1673 (O_1673,N_19880,N_19770);
nor UO_1674 (O_1674,N_15562,N_18430);
or UO_1675 (O_1675,N_16232,N_16117);
or UO_1676 (O_1676,N_15146,N_18631);
or UO_1677 (O_1677,N_15557,N_17321);
and UO_1678 (O_1678,N_18321,N_15034);
or UO_1679 (O_1679,N_19118,N_19018);
nor UO_1680 (O_1680,N_19926,N_15925);
nand UO_1681 (O_1681,N_17008,N_19652);
nand UO_1682 (O_1682,N_17425,N_18853);
nand UO_1683 (O_1683,N_18629,N_15638);
and UO_1684 (O_1684,N_15656,N_15936);
xor UO_1685 (O_1685,N_16959,N_15124);
or UO_1686 (O_1686,N_15817,N_17913);
nor UO_1687 (O_1687,N_17973,N_18834);
or UO_1688 (O_1688,N_17394,N_16931);
xor UO_1689 (O_1689,N_17416,N_18763);
nor UO_1690 (O_1690,N_17443,N_16254);
nor UO_1691 (O_1691,N_17946,N_15148);
and UO_1692 (O_1692,N_18822,N_16264);
or UO_1693 (O_1693,N_16647,N_16229);
or UO_1694 (O_1694,N_18062,N_17510);
nand UO_1695 (O_1695,N_18224,N_19503);
xor UO_1696 (O_1696,N_15832,N_18267);
nor UO_1697 (O_1697,N_19439,N_17024);
xnor UO_1698 (O_1698,N_15150,N_17632);
or UO_1699 (O_1699,N_17286,N_16648);
nor UO_1700 (O_1700,N_19241,N_17552);
nand UO_1701 (O_1701,N_19425,N_17853);
xnor UO_1702 (O_1702,N_16870,N_17433);
and UO_1703 (O_1703,N_15953,N_17291);
xor UO_1704 (O_1704,N_18274,N_15323);
or UO_1705 (O_1705,N_16175,N_19245);
or UO_1706 (O_1706,N_18655,N_18681);
and UO_1707 (O_1707,N_19454,N_15863);
nor UO_1708 (O_1708,N_17733,N_17535);
nand UO_1709 (O_1709,N_18268,N_15177);
and UO_1710 (O_1710,N_19070,N_16493);
nor UO_1711 (O_1711,N_16141,N_18006);
xnor UO_1712 (O_1712,N_17899,N_16462);
nand UO_1713 (O_1713,N_19250,N_18700);
or UO_1714 (O_1714,N_16770,N_17620);
and UO_1715 (O_1715,N_15731,N_17558);
nand UO_1716 (O_1716,N_19637,N_19948);
nand UO_1717 (O_1717,N_17785,N_17004);
nor UO_1718 (O_1718,N_18094,N_16664);
and UO_1719 (O_1719,N_15086,N_19456);
or UO_1720 (O_1720,N_17469,N_16939);
nor UO_1721 (O_1721,N_16400,N_17984);
and UO_1722 (O_1722,N_17847,N_19938);
or UO_1723 (O_1723,N_18978,N_15611);
nand UO_1724 (O_1724,N_16877,N_17012);
nor UO_1725 (O_1725,N_19417,N_17704);
and UO_1726 (O_1726,N_18348,N_15233);
and UO_1727 (O_1727,N_19318,N_19196);
or UO_1728 (O_1728,N_19023,N_18313);
nor UO_1729 (O_1729,N_18147,N_15265);
or UO_1730 (O_1730,N_15407,N_19498);
and UO_1731 (O_1731,N_16449,N_19309);
nor UO_1732 (O_1732,N_15365,N_16885);
xor UO_1733 (O_1733,N_18666,N_19052);
xor UO_1734 (O_1734,N_15858,N_18133);
nand UO_1735 (O_1735,N_16458,N_19074);
nor UO_1736 (O_1736,N_18220,N_17091);
or UO_1737 (O_1737,N_16799,N_19641);
nand UO_1738 (O_1738,N_18871,N_16329);
nor UO_1739 (O_1739,N_16178,N_15453);
or UO_1740 (O_1740,N_18961,N_17147);
or UO_1741 (O_1741,N_15431,N_19994);
or UO_1742 (O_1742,N_19856,N_16912);
nor UO_1743 (O_1743,N_17438,N_19210);
or UO_1744 (O_1744,N_17048,N_17737);
or UO_1745 (O_1745,N_17424,N_16346);
nand UO_1746 (O_1746,N_18004,N_15351);
and UO_1747 (O_1747,N_17136,N_17161);
and UO_1748 (O_1748,N_18758,N_18068);
nand UO_1749 (O_1749,N_15831,N_18353);
nor UO_1750 (O_1750,N_15485,N_18259);
xor UO_1751 (O_1751,N_18386,N_18517);
nor UO_1752 (O_1752,N_17462,N_15134);
or UO_1753 (O_1753,N_17216,N_19192);
or UO_1754 (O_1754,N_18591,N_17542);
nor UO_1755 (O_1755,N_18446,N_15466);
nor UO_1756 (O_1756,N_18693,N_16476);
nor UO_1757 (O_1757,N_18142,N_16587);
and UO_1758 (O_1758,N_19508,N_17969);
nand UO_1759 (O_1759,N_19918,N_17243);
and UO_1760 (O_1760,N_17238,N_18389);
nor UO_1761 (O_1761,N_19658,N_15094);
and UO_1762 (O_1762,N_18169,N_16898);
nor UO_1763 (O_1763,N_17205,N_16649);
nand UO_1764 (O_1764,N_19739,N_15822);
or UO_1765 (O_1765,N_18879,N_16454);
nor UO_1766 (O_1766,N_18540,N_19927);
and UO_1767 (O_1767,N_16831,N_17877);
nor UO_1768 (O_1768,N_18231,N_19782);
or UO_1769 (O_1769,N_19066,N_18777);
nand UO_1770 (O_1770,N_16739,N_15372);
nand UO_1771 (O_1771,N_16744,N_19053);
or UO_1772 (O_1772,N_17888,N_19043);
nand UO_1773 (O_1773,N_15673,N_19848);
and UO_1774 (O_1774,N_15285,N_16804);
nand UO_1775 (O_1775,N_17225,N_17795);
nor UO_1776 (O_1776,N_17548,N_18950);
nor UO_1777 (O_1777,N_18767,N_17717);
and UO_1778 (O_1778,N_18661,N_15187);
or UO_1779 (O_1779,N_16748,N_19608);
xor UO_1780 (O_1780,N_17396,N_17902);
xor UO_1781 (O_1781,N_19756,N_17409);
nand UO_1782 (O_1782,N_18050,N_16399);
nand UO_1783 (O_1783,N_18935,N_17603);
nand UO_1784 (O_1784,N_15655,N_18307);
nand UO_1785 (O_1785,N_15227,N_17634);
xnor UO_1786 (O_1786,N_15989,N_18293);
nand UO_1787 (O_1787,N_16894,N_15330);
or UO_1788 (O_1788,N_18914,N_15949);
nand UO_1789 (O_1789,N_15436,N_18908);
or UO_1790 (O_1790,N_18685,N_15108);
nand UO_1791 (O_1791,N_17815,N_15646);
nand UO_1792 (O_1792,N_18929,N_15442);
nor UO_1793 (O_1793,N_19251,N_15950);
and UO_1794 (O_1794,N_19749,N_16940);
and UO_1795 (O_1795,N_19166,N_18862);
xor UO_1796 (O_1796,N_15700,N_18060);
or UO_1797 (O_1797,N_18378,N_18339);
nand UO_1798 (O_1798,N_15214,N_18739);
nand UO_1799 (O_1799,N_16056,N_17201);
nand UO_1800 (O_1800,N_16025,N_17989);
and UO_1801 (O_1801,N_16440,N_18678);
and UO_1802 (O_1802,N_15228,N_18606);
xnor UO_1803 (O_1803,N_19715,N_18185);
or UO_1804 (O_1804,N_15252,N_15785);
xnor UO_1805 (O_1805,N_16398,N_16177);
nor UO_1806 (O_1806,N_19477,N_18196);
nand UO_1807 (O_1807,N_17255,N_16123);
xnor UO_1808 (O_1808,N_17043,N_18245);
or UO_1809 (O_1809,N_18331,N_19495);
nor UO_1810 (O_1810,N_16085,N_15717);
nand UO_1811 (O_1811,N_16301,N_17678);
and UO_1812 (O_1812,N_17088,N_16701);
nand UO_1813 (O_1813,N_15875,N_19492);
nor UO_1814 (O_1814,N_16745,N_19475);
nand UO_1815 (O_1815,N_15653,N_17371);
nor UO_1816 (O_1816,N_18748,N_19314);
and UO_1817 (O_1817,N_17538,N_18852);
nor UO_1818 (O_1818,N_18900,N_18745);
nand UO_1819 (O_1819,N_16020,N_19988);
nand UO_1820 (O_1820,N_16019,N_17932);
and UO_1821 (O_1821,N_17472,N_19097);
nor UO_1822 (O_1822,N_15110,N_19132);
xnor UO_1823 (O_1823,N_18083,N_19580);
or UO_1824 (O_1824,N_15617,N_17318);
or UO_1825 (O_1825,N_19488,N_18384);
and UO_1826 (O_1826,N_18595,N_18159);
nor UO_1827 (O_1827,N_18782,N_18945);
and UO_1828 (O_1828,N_15661,N_18195);
nor UO_1829 (O_1829,N_15935,N_17162);
or UO_1830 (O_1830,N_17222,N_15531);
nand UO_1831 (O_1831,N_17890,N_18163);
nand UO_1832 (O_1832,N_18435,N_17669);
nor UO_1833 (O_1833,N_16910,N_19667);
xor UO_1834 (O_1834,N_18572,N_17308);
and UO_1835 (O_1835,N_15234,N_17648);
and UO_1836 (O_1836,N_19732,N_16050);
nor UO_1837 (O_1837,N_15710,N_16778);
nand UO_1838 (O_1838,N_18358,N_16923);
nand UO_1839 (O_1839,N_19008,N_18797);
nor UO_1840 (O_1840,N_15254,N_18747);
and UO_1841 (O_1841,N_17402,N_16079);
nor UO_1842 (O_1842,N_15546,N_17302);
nand UO_1843 (O_1843,N_17893,N_16379);
and UO_1844 (O_1844,N_19991,N_16953);
xor UO_1845 (O_1845,N_16167,N_19256);
or UO_1846 (O_1846,N_15589,N_18096);
or UO_1847 (O_1847,N_17964,N_19805);
nor UO_1848 (O_1848,N_19340,N_19599);
and UO_1849 (O_1849,N_19869,N_17520);
and UO_1850 (O_1850,N_18803,N_15163);
xor UO_1851 (O_1851,N_17380,N_15456);
nand UO_1852 (O_1852,N_17554,N_17342);
and UO_1853 (O_1853,N_16585,N_15357);
nor UO_1854 (O_1854,N_19170,N_16380);
or UO_1855 (O_1855,N_15838,N_16080);
nor UO_1856 (O_1856,N_18617,N_16146);
nand UO_1857 (O_1857,N_17435,N_19323);
xor UO_1858 (O_1858,N_16523,N_18592);
and UO_1859 (O_1859,N_16740,N_18125);
or UO_1860 (O_1860,N_18320,N_17288);
or UO_1861 (O_1861,N_15027,N_19741);
and UO_1862 (O_1862,N_19009,N_18645);
nor UO_1863 (O_1863,N_15592,N_15769);
or UO_1864 (O_1864,N_18032,N_19419);
xor UO_1865 (O_1865,N_17685,N_16854);
xnor UO_1866 (O_1866,N_17516,N_19362);
nor UO_1867 (O_1867,N_19347,N_19717);
or UO_1868 (O_1868,N_19246,N_15238);
nand UO_1869 (O_1869,N_17359,N_17099);
nand UO_1870 (O_1870,N_16193,N_16945);
nand UO_1871 (O_1871,N_17170,N_15881);
nand UO_1872 (O_1872,N_15986,N_16889);
nand UO_1873 (O_1873,N_17575,N_19835);
nand UO_1874 (O_1874,N_17256,N_17279);
and UO_1875 (O_1875,N_17705,N_19855);
nor UO_1876 (O_1876,N_16892,N_16753);
nand UO_1877 (O_1877,N_17655,N_16005);
and UO_1878 (O_1878,N_18067,N_16700);
xor UO_1879 (O_1879,N_17528,N_19616);
xor UO_1880 (O_1880,N_15543,N_16998);
and UO_1881 (O_1881,N_15473,N_15481);
and UO_1882 (O_1882,N_18098,N_19671);
nor UO_1883 (O_1883,N_16960,N_16448);
nand UO_1884 (O_1884,N_15085,N_17207);
nand UO_1885 (O_1885,N_17326,N_16074);
and UO_1886 (O_1886,N_19895,N_19744);
and UO_1887 (O_1887,N_16457,N_17956);
nor UO_1888 (O_1888,N_17715,N_19104);
nand UO_1889 (O_1889,N_17586,N_19714);
nor UO_1890 (O_1890,N_15853,N_18609);
and UO_1891 (O_1891,N_16788,N_16611);
or UO_1892 (O_1892,N_15674,N_15425);
and UO_1893 (O_1893,N_17775,N_16077);
nor UO_1894 (O_1894,N_18874,N_19636);
and UO_1895 (O_1895,N_18123,N_18736);
or UO_1896 (O_1896,N_16068,N_18009);
and UO_1897 (O_1897,N_15246,N_19084);
nor UO_1898 (O_1898,N_15417,N_16946);
nor UO_1899 (O_1899,N_17784,N_18795);
nor UO_1900 (O_1900,N_18594,N_15862);
nand UO_1901 (O_1901,N_19445,N_15101);
nand UO_1902 (O_1902,N_15319,N_19264);
or UO_1903 (O_1903,N_15908,N_17303);
and UO_1904 (O_1904,N_19614,N_15877);
and UO_1905 (O_1905,N_19763,N_18670);
nor UO_1906 (O_1906,N_17727,N_19240);
and UO_1907 (O_1907,N_18329,N_18044);
nor UO_1908 (O_1908,N_16695,N_16742);
or UO_1909 (O_1909,N_17398,N_19130);
or UO_1910 (O_1910,N_15208,N_16418);
and UO_1911 (O_1911,N_19935,N_18111);
nor UO_1912 (O_1912,N_17038,N_18910);
nand UO_1913 (O_1913,N_17138,N_19430);
xnor UO_1914 (O_1914,N_15149,N_15806);
nand UO_1915 (O_1915,N_18752,N_18702);
nand UO_1916 (O_1916,N_17149,N_17418);
nor UO_1917 (O_1917,N_15204,N_15025);
or UO_1918 (O_1918,N_15861,N_15359);
nor UO_1919 (O_1919,N_15850,N_15667);
and UO_1920 (O_1920,N_16924,N_15826);
and UO_1921 (O_1921,N_19208,N_19252);
nand UO_1922 (O_1922,N_18712,N_19995);
nor UO_1923 (O_1923,N_16518,N_16326);
nand UO_1924 (O_1924,N_19487,N_17804);
nor UO_1925 (O_1925,N_18586,N_16351);
nand UO_1926 (O_1926,N_15932,N_15258);
nand UO_1927 (O_1927,N_16756,N_15854);
nand UO_1928 (O_1928,N_19227,N_18571);
nor UO_1929 (O_1929,N_18330,N_19398);
or UO_1930 (O_1930,N_15999,N_16769);
nor UO_1931 (O_1931,N_17470,N_15633);
nor UO_1932 (O_1932,N_16273,N_18344);
nand UO_1933 (O_1933,N_16964,N_17660);
and UO_1934 (O_1934,N_18920,N_18662);
nand UO_1935 (O_1935,N_18139,N_18145);
nand UO_1936 (O_1936,N_18175,N_15033);
nor UO_1937 (O_1937,N_15441,N_18738);
or UO_1938 (O_1938,N_15005,N_16851);
and UO_1939 (O_1939,N_16641,N_19355);
and UO_1940 (O_1940,N_17692,N_18890);
or UO_1941 (O_1941,N_17998,N_17652);
nor UO_1942 (O_1942,N_18140,N_15169);
nand UO_1943 (O_1943,N_17489,N_18447);
nor UO_1944 (O_1944,N_15211,N_15528);
and UO_1945 (O_1945,N_15805,N_17747);
or UO_1946 (O_1946,N_15446,N_16423);
and UO_1947 (O_1947,N_16072,N_18315);
and UO_1948 (O_1948,N_16728,N_16652);
nor UO_1949 (O_1949,N_16447,N_16593);
and UO_1950 (O_1950,N_16499,N_19235);
nand UO_1951 (O_1951,N_18967,N_17129);
nand UO_1952 (O_1952,N_19428,N_18304);
nand UO_1953 (O_1953,N_15834,N_19557);
or UO_1954 (O_1954,N_19120,N_18944);
xnor UO_1955 (O_1955,N_15873,N_19348);
nand UO_1956 (O_1956,N_17463,N_17309);
nor UO_1957 (O_1957,N_16127,N_19818);
nand UO_1958 (O_1958,N_15394,N_16022);
nand UO_1959 (O_1959,N_17035,N_17866);
nand UO_1960 (O_1960,N_18126,N_15719);
nand UO_1961 (O_1961,N_15743,N_18692);
and UO_1962 (O_1962,N_16274,N_19654);
and UO_1963 (O_1963,N_18407,N_18058);
nor UO_1964 (O_1964,N_19547,N_17125);
xor UO_1965 (O_1965,N_15130,N_15809);
nor UO_1966 (O_1966,N_16412,N_15886);
nor UO_1967 (O_1967,N_19395,N_17793);
xor UO_1968 (O_1968,N_19977,N_18027);
nor UO_1969 (O_1969,N_16469,N_16021);
and UO_1970 (O_1970,N_16863,N_15264);
xor UO_1971 (O_1971,N_18574,N_16302);
and UO_1972 (O_1972,N_15055,N_16289);
nand UO_1973 (O_1973,N_17200,N_16139);
nand UO_1974 (O_1974,N_17403,N_18323);
nor UO_1975 (O_1975,N_17726,N_18875);
nor UO_1976 (O_1976,N_19850,N_18361);
nand UO_1977 (O_1977,N_18504,N_19474);
nand UO_1978 (O_1978,N_17788,N_17415);
nor UO_1979 (O_1979,N_17051,N_18395);
or UO_1980 (O_1980,N_15889,N_19472);
or UO_1981 (O_1981,N_15533,N_15682);
or UO_1982 (O_1982,N_19907,N_15671);
nand UO_1983 (O_1983,N_18826,N_15763);
nand UO_1984 (O_1984,N_19254,N_15081);
nor UO_1985 (O_1985,N_15506,N_19292);
or UO_1986 (O_1986,N_19807,N_16003);
or UO_1987 (O_1987,N_17037,N_18134);
or UO_1988 (O_1988,N_15235,N_15968);
or UO_1989 (O_1989,N_18568,N_17242);
nand UO_1990 (O_1990,N_18482,N_17246);
and UO_1991 (O_1991,N_18436,N_18087);
and UO_1992 (O_1992,N_15318,N_18375);
nand UO_1993 (O_1993,N_18887,N_19401);
nor UO_1994 (O_1994,N_15023,N_16737);
nor UO_1995 (O_1995,N_17355,N_15926);
or UO_1996 (O_1996,N_18346,N_18966);
and UO_1997 (O_1997,N_19079,N_15312);
and UO_1998 (O_1998,N_16186,N_19705);
and UO_1999 (O_1999,N_15601,N_15062);
and UO_2000 (O_2000,N_19796,N_17055);
xnor UO_2001 (O_2001,N_16715,N_15028);
nor UO_2002 (O_2002,N_18437,N_18065);
or UO_2003 (O_2003,N_19559,N_17152);
and UO_2004 (O_2004,N_19579,N_17460);
nor UO_2005 (O_2005,N_17587,N_15354);
and UO_2006 (O_2006,N_19393,N_17670);
nor UO_2007 (O_2007,N_17825,N_16363);
nor UO_2008 (O_2008,N_15996,N_16291);
nor UO_2009 (O_2009,N_17096,N_18783);
and UO_2010 (O_2010,N_17471,N_16058);
or UO_2011 (O_2011,N_17192,N_16357);
nand UO_2012 (O_2012,N_16767,N_15637);
and UO_2013 (O_2013,N_16150,N_16438);
nor UO_2014 (O_2014,N_15821,N_19415);
and UO_2015 (O_2015,N_15259,N_19274);
nand UO_2016 (O_2016,N_17140,N_19247);
xor UO_2017 (O_2017,N_19035,N_16785);
and UO_2018 (O_2018,N_18043,N_16263);
and UO_2019 (O_2019,N_18170,N_17237);
nor UO_2020 (O_2020,N_19808,N_16714);
or UO_2021 (O_2021,N_18657,N_19320);
and UO_2022 (O_2022,N_16530,N_19775);
and UO_2023 (O_2023,N_16859,N_19540);
and UO_2024 (O_2024,N_19575,N_16096);
nand UO_2025 (O_2025,N_18199,N_15814);
and UO_2026 (O_2026,N_17431,N_18641);
nand UO_2027 (O_2027,N_15625,N_15058);
nor UO_2028 (O_2028,N_16878,N_18723);
and UO_2029 (O_2029,N_17654,N_19765);
nor UO_2030 (O_2030,N_17095,N_15724);
or UO_2031 (O_2031,N_15515,N_16138);
and UO_2032 (O_2032,N_16322,N_16526);
or UO_2033 (O_2033,N_19162,N_15298);
and UO_2034 (O_2034,N_19108,N_17107);
and UO_2035 (O_2035,N_17156,N_18719);
or UO_2036 (O_2036,N_19829,N_16602);
and UO_2037 (O_2037,N_18008,N_18392);
nand UO_2038 (O_2038,N_18554,N_16571);
nand UO_2039 (O_2039,N_19702,N_17923);
and UO_2040 (O_2040,N_19966,N_19489);
nand UO_2041 (O_2041,N_16105,N_16306);
xor UO_2042 (O_2042,N_16431,N_18263);
and UO_2043 (O_2043,N_16718,N_16207);
or UO_2044 (O_2044,N_16101,N_17581);
and UO_2045 (O_2045,N_19844,N_17981);
nand UO_2046 (O_2046,N_19967,N_16991);
xnor UO_2047 (O_2047,N_15911,N_18056);
nor UO_2048 (O_2048,N_16651,N_15898);
or UO_2049 (O_2049,N_17792,N_16387);
xnor UO_2050 (O_2050,N_18302,N_16262);
or UO_2051 (O_2051,N_15125,N_16555);
or UO_2052 (O_2052,N_15780,N_15335);
xor UO_2053 (O_2053,N_19224,N_18290);
xor UO_2054 (O_2054,N_16090,N_16635);
nor UO_2055 (O_2055,N_18611,N_16075);
and UO_2056 (O_2056,N_17702,N_18773);
nand UO_2057 (O_2057,N_19725,N_19243);
xor UO_2058 (O_2058,N_17059,N_18258);
and UO_2059 (O_2059,N_18672,N_17500);
or UO_2060 (O_2060,N_18424,N_18491);
xor UO_2061 (O_2061,N_19450,N_18250);
nor UO_2062 (O_2062,N_17244,N_15278);
and UO_2063 (O_2063,N_18911,N_18377);
and UO_2064 (O_2064,N_17777,N_19086);
xnor UO_2065 (O_2065,N_19951,N_19188);
nand UO_2066 (O_2066,N_18074,N_16781);
nor UO_2067 (O_2067,N_19180,N_17918);
or UO_2068 (O_2068,N_19266,N_17289);
or UO_2069 (O_2069,N_17598,N_19284);
and UO_2070 (O_2070,N_17745,N_16754);
nor UO_2071 (O_2071,N_17943,N_15268);
nor UO_2072 (O_2072,N_16352,N_19793);
or UO_2073 (O_2073,N_17323,N_16335);
nand UO_2074 (O_2074,N_19190,N_17615);
or UO_2075 (O_2075,N_17007,N_16720);
or UO_2076 (O_2076,N_19822,N_18559);
or UO_2077 (O_2077,N_15501,N_18208);
and UO_2078 (O_2078,N_17177,N_16482);
and UO_2079 (O_2079,N_15569,N_15588);
nand UO_2080 (O_2080,N_18239,N_17987);
or UO_2081 (O_2081,N_15759,N_15708);
and UO_2082 (O_2082,N_16824,N_17627);
and UO_2083 (O_2083,N_17363,N_17250);
or UO_2084 (O_2084,N_17521,N_18790);
and UO_2085 (O_2085,N_19102,N_16052);
or UO_2086 (O_2086,N_19843,N_15090);
or UO_2087 (O_2087,N_19582,N_17253);
xor UO_2088 (O_2088,N_17639,N_17783);
nand UO_2089 (O_2089,N_15847,N_15136);
nand UO_2090 (O_2090,N_16678,N_19605);
and UO_2091 (O_2091,N_19798,N_18793);
xnor UO_2092 (O_2092,N_16667,N_19669);
and UO_2093 (O_2093,N_17797,N_15888);
or UO_2094 (O_2094,N_15516,N_18476);
nand UO_2095 (O_2095,N_19552,N_16650);
or UO_2096 (O_2096,N_15390,N_18112);
nand UO_2097 (O_2097,N_17497,N_16053);
and UO_2098 (O_2098,N_16433,N_17626);
or UO_2099 (O_2099,N_17929,N_19093);
or UO_2100 (O_2100,N_17691,N_15797);
nand UO_2101 (O_2101,N_15829,N_15621);
or UO_2102 (O_2102,N_16153,N_16792);
or UO_2103 (O_2103,N_17907,N_16378);
xor UO_2104 (O_2104,N_18754,N_16174);
nor UO_2105 (O_2105,N_19418,N_15827);
or UO_2106 (O_2106,N_16613,N_19564);
nor UO_2107 (O_2107,N_17920,N_17512);
nand UO_2108 (O_2108,N_18983,N_16992);
xor UO_2109 (O_2109,N_19286,N_17683);
xor UO_2110 (O_2110,N_18089,N_18296);
or UO_2111 (O_2111,N_18838,N_19709);
nand UO_2112 (O_2112,N_17233,N_18801);
xor UO_2113 (O_2113,N_17573,N_15698);
nor UO_2114 (O_2114,N_19516,N_16803);
nor UO_2115 (O_2115,N_15952,N_16707);
nand UO_2116 (O_2116,N_15121,N_15587);
nand UO_2117 (O_2117,N_19000,N_18894);
nand UO_2118 (O_2118,N_19073,N_19780);
or UO_2119 (O_2119,N_15089,N_18101);
nand UO_2120 (O_2120,N_16426,N_19976);
nand UO_2121 (O_2121,N_16836,N_15741);
and UO_2122 (O_2122,N_19343,N_15733);
or UO_2123 (O_2123,N_16633,N_16845);
nand UO_2124 (O_2124,N_19156,N_15550);
nand UO_2125 (O_2125,N_19736,N_15776);
and UO_2126 (O_2126,N_19838,N_16406);
or UO_2127 (O_2127,N_19080,N_19890);
and UO_2128 (O_2128,N_17997,N_16087);
or UO_2129 (O_2129,N_19291,N_18551);
nor UO_2130 (O_2130,N_19596,N_17307);
or UO_2131 (O_2131,N_17819,N_16833);
and UO_2132 (O_2132,N_15649,N_19091);
xor UO_2133 (O_2133,N_19354,N_15040);
or UO_2134 (O_2134,N_18545,N_18204);
nand UO_2135 (O_2135,N_19758,N_15603);
nand UO_2136 (O_2136,N_17623,N_18519);
and UO_2137 (O_2137,N_16026,N_15116);
or UO_2138 (O_2138,N_19497,N_16874);
nand UO_2139 (O_2139,N_17473,N_17666);
and UO_2140 (O_2140,N_18298,N_18530);
nand UO_2141 (O_2141,N_19558,N_18780);
nor UO_2142 (O_2142,N_19902,N_15181);
and UO_2143 (O_2143,N_15788,N_16705);
and UO_2144 (O_2144,N_17022,N_16537);
and UO_2145 (O_2145,N_16907,N_16798);
or UO_2146 (O_2146,N_18960,N_16364);
or UO_2147 (O_2147,N_18472,N_17467);
nand UO_2148 (O_2148,N_16258,N_17198);
nand UO_2149 (O_2149,N_17896,N_18164);
or UO_2150 (O_2150,N_18981,N_16029);
nand UO_2151 (O_2151,N_16214,N_18093);
nor UO_2152 (O_2152,N_18171,N_17071);
nor UO_2153 (O_2153,N_18705,N_16182);
nand UO_2154 (O_2154,N_19859,N_15404);
and UO_2155 (O_2155,N_16777,N_18022);
nor UO_2156 (O_2156,N_19584,N_17427);
and UO_2157 (O_2157,N_16192,N_18041);
or UO_2158 (O_2158,N_19662,N_18743);
xor UO_2159 (O_2159,N_19289,N_15185);
or UO_2160 (O_2160,N_15736,N_19681);
nand UO_2161 (O_2161,N_16875,N_18789);
nand UO_2162 (O_2162,N_17451,N_18496);
nand UO_2163 (O_2163,N_15799,N_19687);
xor UO_2164 (O_2164,N_18821,N_18373);
and UO_2165 (O_2165,N_15229,N_16419);
nor UO_2166 (O_2166,N_17844,N_18445);
nor UO_2167 (O_2167,N_19600,N_16918);
nor UO_2168 (O_2168,N_18589,N_17971);
nor UO_2169 (O_2169,N_15884,N_15830);
nor UO_2170 (O_2170,N_18286,N_18458);
and UO_2171 (O_2171,N_15498,N_17230);
nor UO_2172 (O_2172,N_17109,N_19085);
and UO_2173 (O_2173,N_16124,N_17962);
or UO_2174 (O_2174,N_15042,N_16776);
xnor UO_2175 (O_2175,N_16914,N_17625);
and UO_2176 (O_2176,N_15507,N_16047);
xor UO_2177 (O_2177,N_17228,N_18213);
or UO_2178 (O_2178,N_19804,N_15317);
nor UO_2179 (O_2179,N_19962,N_18023);
xnor UO_2180 (O_2180,N_16017,N_17744);
and UO_2181 (O_2181,N_19374,N_17764);
and UO_2182 (O_2182,N_18563,N_17659);
and UO_2183 (O_2183,N_15644,N_18266);
or UO_2184 (O_2184,N_17241,N_18024);
nor UO_2185 (O_2185,N_16394,N_16837);
nor UO_2186 (O_2186,N_17421,N_16661);
xor UO_2187 (O_2187,N_18086,N_17133);
nand UO_2188 (O_2188,N_19184,N_17458);
nand UO_2189 (O_2189,N_19572,N_19030);
xor UO_2190 (O_2190,N_17845,N_16309);
nand UO_2191 (O_2191,N_16443,N_15561);
or UO_2192 (O_2192,N_16538,N_18755);
and UO_2193 (O_2193,N_16381,N_17492);
or UO_2194 (O_2194,N_17358,N_16732);
and UO_2195 (O_2195,N_16972,N_15518);
or UO_2196 (O_2196,N_19329,N_19968);
or UO_2197 (O_2197,N_17649,N_18473);
and UO_2198 (O_2198,N_15883,N_16276);
nand UO_2199 (O_2199,N_18440,N_19959);
nor UO_2200 (O_2200,N_19100,N_16287);
xnor UO_2201 (O_2201,N_15947,N_19659);
nand UO_2202 (O_2202,N_19515,N_18454);
xor UO_2203 (O_2203,N_16347,N_17992);
nand UO_2204 (O_2204,N_17572,N_18359);
nor UO_2205 (O_2205,N_15448,N_19225);
and UO_2206 (O_2206,N_18880,N_16800);
and UO_2207 (O_2207,N_19173,N_18627);
nor UO_2208 (O_2208,N_16421,N_15402);
nor UO_2209 (O_2209,N_17513,N_19405);
and UO_2210 (O_2210,N_18233,N_17420);
or UO_2211 (O_2211,N_16941,N_15209);
nor UO_2212 (O_2212,N_18235,N_18247);
or UO_2213 (O_2213,N_16645,N_16216);
or UO_2214 (O_2214,N_19335,N_16217);
and UO_2215 (O_2215,N_15909,N_15948);
nor UO_2216 (O_2216,N_17120,N_19022);
nor UO_2217 (O_2217,N_18811,N_16275);
xor UO_2218 (O_2218,N_16600,N_15907);
xnor UO_2219 (O_2219,N_17800,N_17937);
or UO_2220 (O_2220,N_15500,N_16031);
or UO_2221 (O_2221,N_15221,N_16688);
nor UO_2222 (O_2222,N_18276,N_18537);
nor UO_2223 (O_2223,N_15939,N_19491);
and UO_2224 (O_2224,N_19049,N_18347);
nor UO_2225 (O_2225,N_18781,N_19172);
nand UO_2226 (O_2226,N_18416,N_17264);
and UO_2227 (O_2227,N_18831,N_19597);
xor UO_2228 (O_2228,N_15779,N_18316);
and UO_2229 (O_2229,N_16981,N_16669);
and UO_2230 (O_2230,N_18341,N_18889);
and UO_2231 (O_2231,N_17105,N_18128);
and UO_2232 (O_2232,N_16755,N_18582);
nand UO_2233 (O_2233,N_17806,N_16591);
and UO_2234 (O_2234,N_18548,N_17752);
nor UO_2235 (O_2235,N_17826,N_15596);
nor UO_2236 (O_2236,N_17986,N_17555);
and UO_2237 (O_2237,N_17954,N_17100);
and UO_2238 (O_2238,N_18036,N_16271);
nand UO_2239 (O_2239,N_18684,N_18244);
nor UO_2240 (O_2240,N_19936,N_16147);
nand UO_2241 (O_2241,N_18902,N_19071);
xor UO_2242 (O_2242,N_17519,N_18909);
or UO_2243 (O_2243,N_18836,N_17385);
nor UO_2244 (O_2244,N_15659,N_16515);
and UO_2245 (O_2245,N_19056,N_18240);
nor UO_2246 (O_2246,N_18414,N_15902);
xnor UO_2247 (O_2247,N_18918,N_19414);
nor UO_2248 (O_2248,N_18671,N_15956);
or UO_2249 (O_2249,N_15784,N_19865);
or UO_2250 (O_2250,N_17843,N_17494);
and UO_2251 (O_2251,N_15004,N_15183);
nand UO_2252 (O_2252,N_19459,N_17699);
xnor UO_2253 (O_2253,N_17567,N_16290);
nand UO_2254 (O_2254,N_15836,N_16590);
and UO_2255 (O_2255,N_17846,N_18976);
or UO_2256 (O_2256,N_17859,N_18511);
and UO_2257 (O_2257,N_18338,N_16796);
nand UO_2258 (O_2258,N_15762,N_16956);
nor UO_2259 (O_2259,N_18835,N_18869);
and UO_2260 (O_2260,N_16622,N_19383);
or UO_2261 (O_2261,N_16278,N_17282);
nor UO_2262 (O_2262,N_17179,N_19961);
nand UO_2263 (O_2263,N_17280,N_19099);
or UO_2264 (O_2264,N_16169,N_19183);
nor UO_2265 (O_2265,N_19381,N_16500);
nor UO_2266 (O_2266,N_18883,N_15104);
nor UO_2267 (O_2267,N_17090,N_15786);
nor UO_2268 (O_2268,N_15073,N_18555);
nand UO_2269 (O_2269,N_15075,N_16281);
or UO_2270 (O_2270,N_16736,N_15206);
xor UO_2271 (O_2271,N_19004,N_18823);
nor UO_2272 (O_2272,N_17531,N_18620);
or UO_2273 (O_2273,N_19001,N_18954);
nor UO_2274 (O_2274,N_16820,N_19819);
nand UO_2275 (O_2275,N_19785,N_19334);
and UO_2276 (O_2276,N_18400,N_16786);
nand UO_2277 (O_2277,N_15275,N_18569);
and UO_2278 (O_2278,N_17641,N_15478);
or UO_2279 (O_2279,N_17693,N_19295);
and UO_2280 (O_2280,N_15310,N_19999);
nand UO_2281 (O_2281,N_19985,N_17862);
nor UO_2282 (O_2282,N_18550,N_19165);
xor UO_2283 (O_2283,N_15348,N_16424);
and UO_2284 (O_2284,N_19443,N_17875);
or UO_2285 (O_2285,N_18930,N_16793);
nor UO_2286 (O_2286,N_19135,N_17934);
nand UO_2287 (O_2287,N_16531,N_17709);
or UO_2288 (O_2288,N_15522,N_19983);
or UO_2289 (O_2289,N_18735,N_16986);
or UO_2290 (O_2290,N_15295,N_15379);
xor UO_2291 (O_2291,N_17757,N_18707);
nor UO_2292 (O_2292,N_16540,N_16465);
and UO_2293 (O_2293,N_18311,N_15567);
xnor UO_2294 (O_2294,N_18039,N_19394);
and UO_2295 (O_2295,N_17074,N_18218);
or UO_2296 (O_2296,N_16703,N_15944);
or UO_2297 (O_2297,N_16392,N_18597);
nand UO_2298 (O_2298,N_15082,N_17213);
or UO_2299 (O_2299,N_19755,N_19200);
xnor UO_2300 (O_2300,N_15963,N_17940);
nand UO_2301 (O_2301,N_17150,N_16672);
or UO_2302 (O_2302,N_16839,N_19760);
and UO_2303 (O_2303,N_17816,N_15460);
or UO_2304 (O_2304,N_15870,N_19054);
or UO_2305 (O_2305,N_17135,N_19185);
and UO_2306 (O_2306,N_15504,N_15428);
or UO_2307 (O_2307,N_16619,N_19325);
or UO_2308 (O_2308,N_18614,N_17036);
or UO_2309 (O_2309,N_17086,N_17351);
or UO_2310 (O_2310,N_18362,N_16112);
or UO_2311 (O_2311,N_18660,N_16039);
xor UO_2312 (O_2312,N_16478,N_17269);
xor UO_2313 (O_2313,N_17260,N_17941);
nor UO_2314 (O_2314,N_15409,N_17982);
or UO_2315 (O_2315,N_15942,N_18903);
nand UO_2316 (O_2316,N_16403,N_15660);
or UO_2317 (O_2317,N_17063,N_15388);
or UO_2318 (O_2318,N_15636,N_18480);
nor UO_2319 (O_2319,N_16243,N_19550);
and UO_2320 (O_2320,N_18116,N_15153);
nand UO_2321 (O_2321,N_16032,N_15482);
nand UO_2322 (O_2322,N_19391,N_17713);
or UO_2323 (O_2323,N_15020,N_15113);
nand UO_2324 (O_2324,N_17306,N_17009);
or UO_2325 (O_2325,N_19342,N_18765);
xnor UO_2326 (O_2326,N_17428,N_18034);
nand UO_2327 (O_2327,N_16990,N_16059);
or UO_2328 (O_2328,N_16794,N_16115);
or UO_2329 (O_2329,N_17527,N_18827);
nand UO_2330 (O_2330,N_15263,N_19729);
nand UO_2331 (O_2331,N_15652,N_18215);
xor UO_2332 (O_2332,N_18512,N_18292);
and UO_2333 (O_2333,N_19193,N_18277);
nand UO_2334 (O_2334,N_15147,N_17524);
xor UO_2335 (O_2335,N_18636,N_18839);
and UO_2336 (O_2336,N_16543,N_18809);
xor UO_2337 (O_2337,N_17345,N_19138);
and UO_2338 (O_2338,N_19067,N_19947);
nor UO_2339 (O_2339,N_18683,N_17742);
nand UO_2340 (O_2340,N_19806,N_16896);
xor UO_2341 (O_2341,N_15610,N_17248);
nand UO_2342 (O_2342,N_15718,N_15608);
or UO_2343 (O_2343,N_18778,N_15419);
and UO_2344 (O_2344,N_18541,N_17173);
or UO_2345 (O_2345,N_19007,N_19380);
nand UO_2346 (O_2346,N_15517,N_19581);
nand UO_2347 (O_2347,N_15251,N_18212);
nor UO_2348 (O_2348,N_17112,N_16949);
nand UO_2349 (O_2349,N_19511,N_17580);
or UO_2350 (O_2350,N_16168,N_18638);
nand UO_2351 (O_2351,N_17026,N_17175);
nand UO_2352 (O_2352,N_19897,N_16886);
xor UO_2353 (O_2353,N_15414,N_15692);
xnor UO_2354 (O_2354,N_19612,N_18556);
or UO_2355 (O_2355,N_19905,N_18040);
and UO_2356 (O_2356,N_19300,N_16502);
or UO_2357 (O_2357,N_18325,N_18077);
and UO_2358 (O_2358,N_16042,N_16420);
or UO_2359 (O_2359,N_19253,N_15774);
and UO_2360 (O_2360,N_17033,N_16681);
nand UO_2361 (O_2361,N_18915,N_16501);
xnor UO_2362 (O_2362,N_15642,N_16917);
nand UO_2363 (O_2363,N_18481,N_16356);
nand UO_2364 (O_2364,N_17878,N_16614);
or UO_2365 (O_2365,N_19910,N_19311);
or UO_2366 (O_2366,N_15657,N_18148);
and UO_2367 (O_2367,N_15286,N_17751);
or UO_2368 (O_2368,N_19163,N_17417);
nor UO_2369 (O_2369,N_19701,N_17031);
and UO_2370 (O_2370,N_17762,N_15666);
nor UO_2371 (O_2371,N_15241,N_19158);
nor UO_2372 (O_2372,N_15828,N_19541);
nor UO_2373 (O_2373,N_17560,N_18319);
nor UO_2374 (O_2374,N_16185,N_18026);
and UO_2375 (O_2375,N_16768,N_16144);
and UO_2376 (O_2376,N_15765,N_15626);
xor UO_2377 (O_2377,N_19832,N_18017);
or UO_2378 (O_2378,N_18520,N_16954);
or UO_2379 (O_2379,N_16685,N_15077);
or UO_2380 (O_2380,N_19598,N_18942);
or UO_2381 (O_2381,N_19262,N_18643);
nand UO_2382 (O_2382,N_15709,N_16533);
or UO_2383 (O_2383,N_17259,N_18405);
nand UO_2384 (O_2384,N_15047,N_15277);
nand UO_2385 (O_2385,N_19146,N_16573);
nand UO_2386 (O_2386,N_16698,N_19784);
or UO_2387 (O_2387,N_19903,N_17763);
nor UO_2388 (O_2388,N_16967,N_16766);
nor UO_2389 (O_2389,N_19929,N_16977);
or UO_2390 (O_2390,N_18421,N_16268);
and UO_2391 (O_2391,N_18509,N_16827);
nand UO_2392 (O_2392,N_19710,N_15154);
and UO_2393 (O_2393,N_17167,N_19923);
and UO_2394 (O_2394,N_17461,N_19955);
nor UO_2395 (O_2395,N_19623,N_19400);
nand UO_2396 (O_2396,N_19664,N_17728);
or UO_2397 (O_2397,N_16338,N_16569);
nand UO_2398 (O_2398,N_17605,N_18840);
or UO_2399 (O_2399,N_16086,N_18345);
and UO_2400 (O_2400,N_18092,N_15851);
nor UO_2401 (O_2401,N_18646,N_17503);
nor UO_2402 (O_2402,N_19338,N_19141);
xor UO_2403 (O_2403,N_15207,N_16450);
nor UO_2404 (O_2404,N_19479,N_18804);
or UO_2405 (O_2405,N_19693,N_19997);
nand UO_2406 (O_2406,N_17128,N_18786);
xnor UO_2407 (O_2407,N_19040,N_19900);
xnor UO_2408 (O_2408,N_15079,N_18539);
and UO_2409 (O_2409,N_16882,N_15375);
and UO_2410 (O_2410,N_16279,N_15706);
xor UO_2411 (O_2411,N_17824,N_18364);
and UO_2412 (O_2412,N_19886,N_17798);
or UO_2413 (O_2413,N_16809,N_15835);
xnor UO_2414 (O_2414,N_17392,N_15240);
and UO_2415 (O_2415,N_18411,N_18394);
or UO_2416 (O_2416,N_16033,N_18764);
nand UO_2417 (O_2417,N_15650,N_16386);
and UO_2418 (O_2418,N_17613,N_15249);
nor UO_2419 (O_2419,N_18317,N_19786);
nand UO_2420 (O_2420,N_15808,N_16131);
and UO_2421 (O_2421,N_15054,N_16618);
nor UO_2422 (O_2422,N_15510,N_19092);
and UO_2423 (O_2423,N_16790,N_16599);
or UO_2424 (O_2424,N_15031,N_17057);
or UO_2425 (O_2425,N_16189,N_19341);
nor UO_2426 (O_2426,N_15363,N_15426);
or UO_2427 (O_2427,N_17933,N_19862);
and UO_2428 (O_2428,N_19590,N_17375);
and UO_2429 (O_2429,N_19810,N_18419);
xor UO_2430 (O_2430,N_17187,N_19065);
or UO_2431 (O_2431,N_15222,N_16497);
nand UO_2432 (O_2432,N_16580,N_18895);
and UO_2433 (O_2433,N_15766,N_15194);
or UO_2434 (O_2434,N_18342,N_18490);
nand UO_2435 (O_2435,N_18868,N_18444);
or UO_2436 (O_2436,N_15327,N_18284);
nand UO_2437 (O_2437,N_19420,N_18241);
nand UO_2438 (O_2438,N_16201,N_18975);
nand UO_2439 (O_2439,N_18066,N_15231);
and UO_2440 (O_2440,N_18141,N_15900);
or UO_2441 (O_2441,N_18402,N_17444);
and UO_2442 (O_2442,N_15483,N_17577);
and UO_2443 (O_2443,N_16852,N_16846);
and UO_2444 (O_2444,N_18352,N_15654);
nor UO_2445 (O_2445,N_16951,N_18741);
or UO_2446 (O_2446,N_17018,N_15519);
or UO_2447 (O_2447,N_19148,N_17799);
or UO_2448 (O_2448,N_16205,N_19306);
or UO_2449 (O_2449,N_16094,N_16014);
and UO_2450 (O_2450,N_16343,N_16140);
nor UO_2451 (O_2451,N_19530,N_17476);
nand UO_2452 (O_2452,N_17597,N_16098);
or UO_2453 (O_2453,N_18585,N_16320);
nor UO_2454 (O_2454,N_16857,N_16957);
nor UO_2455 (O_2455,N_18686,N_15538);
nor UO_2456 (O_2456,N_17310,N_17856);
xnor UO_2457 (O_2457,N_16983,N_18441);
nor UO_2458 (O_2458,N_16376,N_18264);
nand UO_2459 (O_2459,N_16196,N_17507);
xor UO_2460 (O_2460,N_16136,N_18343);
and UO_2461 (O_2461,N_17429,N_19719);
nand UO_2462 (O_2462,N_19958,N_18896);
and UO_2463 (O_2463,N_19006,N_15103);
nand UO_2464 (O_2464,N_16051,N_19294);
and UO_2465 (O_2465,N_19350,N_16453);
or UO_2466 (O_2466,N_15604,N_18243);
nor UO_2467 (O_2467,N_16073,N_19426);
xor UO_2468 (O_2468,N_19087,N_17925);
and UO_2469 (O_2469,N_15391,N_18972);
or UO_2470 (O_2470,N_17725,N_17076);
nor UO_2471 (O_2471,N_17284,N_17761);
nor UO_2472 (O_2472,N_19209,N_15188);
nor UO_2473 (O_2473,N_18450,N_19145);
nor UO_2474 (O_2474,N_18602,N_15464);
xnor UO_2475 (O_2475,N_19046,N_15066);
and UO_2476 (O_2476,N_15742,N_17588);
and UO_2477 (O_2477,N_18399,N_16474);
nand UO_2478 (O_2478,N_15439,N_19187);
or UO_2479 (O_2479,N_17400,N_19069);
nor UO_2480 (O_2480,N_15232,N_19527);
and UO_2481 (O_2481,N_18579,N_17218);
nand UO_2482 (O_2482,N_19015,N_15202);
nand UO_2483 (O_2483,N_16341,N_16470);
nor UO_2484 (O_2484,N_17600,N_16895);
or UO_2485 (O_2485,N_19261,N_18613);
nand UO_2486 (O_2486,N_19943,N_18986);
or UO_2487 (O_2487,N_19989,N_19467);
nand UO_2488 (O_2488,N_15182,N_16616);
nand UO_2489 (O_2489,N_19589,N_16340);
nor UO_2490 (O_2490,N_15191,N_19005);
or UO_2491 (O_2491,N_17840,N_17436);
nand UO_2492 (O_2492,N_19913,N_18709);
nand UO_2493 (O_2493,N_15270,N_18703);
or UO_2494 (O_2494,N_18459,N_17019);
nand UO_2495 (O_2495,N_18031,N_17892);
nor UO_2496 (O_2496,N_16307,N_19371);
or UO_2497 (O_2497,N_16062,N_19424);
or UO_2498 (O_2498,N_18612,N_16865);
nor UO_2499 (O_2499,N_17384,N_18162);
endmodule