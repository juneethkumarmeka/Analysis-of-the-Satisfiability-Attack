module basic_500_3000_500_6_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_154,In_134);
xor U1 (N_1,In_348,In_332);
nor U2 (N_2,In_319,In_226);
nor U3 (N_3,In_264,In_283);
nor U4 (N_4,In_446,In_150);
or U5 (N_5,In_377,In_478);
xnor U6 (N_6,In_441,In_102);
or U7 (N_7,In_144,In_479);
nand U8 (N_8,In_162,In_176);
xnor U9 (N_9,In_465,In_214);
nor U10 (N_10,In_422,In_300);
and U11 (N_11,In_367,In_216);
xor U12 (N_12,In_69,In_492);
xor U13 (N_13,In_420,In_288);
nor U14 (N_14,In_329,In_19);
or U15 (N_15,In_299,In_490);
nand U16 (N_16,In_67,In_29);
nand U17 (N_17,In_91,In_309);
nor U18 (N_18,In_239,In_237);
and U19 (N_19,In_499,In_114);
nand U20 (N_20,In_228,In_271);
or U21 (N_21,In_470,In_129);
nand U22 (N_22,In_388,In_54);
xor U23 (N_23,In_457,In_336);
nand U24 (N_24,In_431,In_368);
nor U25 (N_25,In_408,In_273);
nor U26 (N_26,In_2,In_27);
or U27 (N_27,In_168,In_217);
and U28 (N_28,In_241,In_170);
xnor U29 (N_29,In_439,In_254);
nor U30 (N_30,In_113,In_175);
nand U31 (N_31,In_22,In_167);
nor U32 (N_32,In_28,In_455);
xnor U33 (N_33,In_306,In_58);
nand U34 (N_34,In_375,In_249);
and U35 (N_35,In_342,In_235);
xnor U36 (N_36,In_65,In_157);
and U37 (N_37,In_253,In_463);
nor U38 (N_38,In_140,In_277);
nand U39 (N_39,In_469,In_234);
or U40 (N_40,In_247,In_250);
and U41 (N_41,In_355,In_89);
nor U42 (N_42,In_440,In_75);
and U43 (N_43,In_314,In_148);
and U44 (N_44,In_371,In_40);
and U45 (N_45,In_460,In_25);
nand U46 (N_46,In_409,In_96);
and U47 (N_47,In_7,In_396);
or U48 (N_48,In_407,In_198);
nand U49 (N_49,In_10,In_100);
xor U50 (N_50,In_321,In_328);
xor U51 (N_51,In_475,In_381);
nand U52 (N_52,In_77,In_155);
xnor U53 (N_53,In_401,In_106);
nor U54 (N_54,In_472,In_483);
and U55 (N_55,In_413,In_163);
or U56 (N_56,In_278,In_193);
xnor U57 (N_57,In_343,In_384);
or U58 (N_58,In_59,In_192);
and U59 (N_59,In_185,In_275);
nand U60 (N_60,In_191,In_379);
nand U61 (N_61,In_11,In_382);
or U62 (N_62,In_24,In_435);
and U63 (N_63,In_233,In_410);
or U64 (N_64,In_412,In_3);
xor U65 (N_65,In_444,In_145);
nor U66 (N_66,In_310,In_95);
or U67 (N_67,In_256,In_202);
xnor U68 (N_68,In_189,In_262);
nor U69 (N_69,In_52,In_138);
or U70 (N_70,In_484,In_279);
nand U71 (N_71,In_419,In_205);
and U72 (N_72,In_464,In_298);
xor U73 (N_73,In_60,In_203);
xnor U74 (N_74,In_4,In_426);
xnor U75 (N_75,In_97,In_304);
or U76 (N_76,In_130,In_20);
and U77 (N_77,In_180,In_161);
nor U78 (N_78,In_17,In_82);
xnor U79 (N_79,In_477,In_334);
xor U80 (N_80,In_125,In_90);
and U81 (N_81,In_160,In_195);
nor U82 (N_82,In_18,In_156);
or U83 (N_83,In_119,In_397);
nor U84 (N_84,In_317,In_196);
nand U85 (N_85,In_456,In_493);
nor U86 (N_86,In_392,In_146);
or U87 (N_87,In_378,In_281);
nor U88 (N_88,In_313,In_432);
nand U89 (N_89,In_93,In_56);
nor U90 (N_90,In_496,In_399);
and U91 (N_91,In_68,In_311);
xnor U92 (N_92,In_225,In_224);
nor U93 (N_93,In_221,In_359);
and U94 (N_94,In_26,In_108);
xnor U95 (N_95,In_395,In_248);
nor U96 (N_96,In_482,In_322);
or U97 (N_97,In_448,In_473);
nand U98 (N_98,In_172,In_383);
nand U99 (N_99,In_324,In_347);
xnor U100 (N_100,In_269,In_133);
nand U101 (N_101,In_474,In_428);
nor U102 (N_102,In_0,In_476);
nor U103 (N_103,In_284,In_462);
xor U104 (N_104,In_291,In_468);
nand U105 (N_105,In_165,In_307);
xnor U106 (N_106,In_453,In_323);
and U107 (N_107,In_230,In_268);
xnor U108 (N_108,In_101,In_66);
or U109 (N_109,In_8,In_201);
xor U110 (N_110,In_466,In_227);
nor U111 (N_111,In_364,In_238);
or U112 (N_112,In_6,In_489);
or U113 (N_113,In_84,In_416);
nor U114 (N_114,In_78,In_70);
nor U115 (N_115,In_480,In_151);
and U116 (N_116,In_251,In_427);
or U117 (N_117,In_210,In_337);
or U118 (N_118,In_481,In_71);
nand U119 (N_119,In_23,In_370);
or U120 (N_120,In_99,In_158);
or U121 (N_121,In_433,In_485);
nor U122 (N_122,In_385,In_13);
and U123 (N_123,In_153,In_449);
nor U124 (N_124,In_178,In_118);
xor U125 (N_125,In_37,In_1);
xnor U126 (N_126,In_445,In_361);
nor U127 (N_127,In_246,In_325);
nor U128 (N_128,In_139,In_423);
xnor U129 (N_129,In_120,In_83);
xnor U130 (N_130,In_169,In_174);
or U131 (N_131,In_286,In_41);
xor U132 (N_132,In_64,In_394);
and U133 (N_133,In_207,In_199);
and U134 (N_134,In_498,In_110);
and U135 (N_135,In_197,In_30);
and U136 (N_136,In_86,In_272);
nor U137 (N_137,In_187,In_265);
and U138 (N_138,In_81,In_400);
nand U139 (N_139,In_403,In_57);
and U140 (N_140,In_209,In_297);
and U141 (N_141,In_62,In_51);
and U142 (N_142,In_318,In_72);
and U143 (N_143,In_236,In_344);
nor U144 (N_144,In_424,In_380);
nor U145 (N_145,In_222,In_345);
nand U146 (N_146,In_231,In_471);
or U147 (N_147,In_141,In_351);
nor U148 (N_148,In_285,In_338);
nand U149 (N_149,In_16,In_31);
and U150 (N_150,In_142,In_458);
and U151 (N_151,In_147,In_346);
and U152 (N_152,In_88,In_121);
and U153 (N_153,In_208,In_443);
xor U154 (N_154,In_495,In_461);
nand U155 (N_155,In_46,In_244);
and U156 (N_156,In_255,In_166);
xnor U157 (N_157,In_267,In_74);
and U158 (N_158,In_402,In_429);
xnor U159 (N_159,In_190,In_127);
nor U160 (N_160,In_365,In_186);
xnor U161 (N_161,In_372,In_131);
nor U162 (N_162,In_450,In_117);
and U163 (N_163,In_15,In_260);
nand U164 (N_164,In_386,In_316);
or U165 (N_165,In_112,In_327);
or U166 (N_166,In_404,In_105);
or U167 (N_167,In_252,In_376);
and U168 (N_168,In_296,In_341);
nand U169 (N_169,In_358,In_94);
and U170 (N_170,In_135,In_21);
or U171 (N_171,In_352,In_497);
and U172 (N_172,In_47,In_418);
or U173 (N_173,In_92,In_374);
or U174 (N_174,In_486,In_350);
xor U175 (N_175,In_335,In_159);
nand U176 (N_176,In_390,In_293);
or U177 (N_177,In_290,In_173);
nor U178 (N_178,In_292,In_44);
nand U179 (N_179,In_398,In_276);
nand U180 (N_180,In_63,In_220);
xnor U181 (N_181,In_331,In_242);
and U182 (N_182,In_38,In_5);
nand U183 (N_183,In_451,In_48);
nor U184 (N_184,In_35,In_308);
or U185 (N_185,In_182,In_274);
or U186 (N_186,In_312,In_411);
xnor U187 (N_187,In_436,In_415);
and U188 (N_188,In_85,In_417);
nand U189 (N_189,In_393,In_76);
xnor U190 (N_190,In_266,In_188);
nor U191 (N_191,In_194,In_326);
nand U192 (N_192,In_315,In_289);
xor U193 (N_193,In_240,In_55);
or U194 (N_194,In_211,In_467);
xor U195 (N_195,In_164,In_137);
and U196 (N_196,In_184,In_109);
or U197 (N_197,In_103,In_366);
and U198 (N_198,In_282,In_179);
or U199 (N_199,In_49,In_183);
or U200 (N_200,In_333,In_421);
xnor U201 (N_201,In_123,In_434);
or U202 (N_202,In_305,In_438);
and U203 (N_203,In_301,In_212);
and U204 (N_204,In_124,In_107);
or U205 (N_205,In_330,In_181);
or U206 (N_206,In_459,In_295);
nand U207 (N_207,In_294,In_362);
xnor U208 (N_208,In_149,In_487);
and U209 (N_209,In_213,In_363);
nor U210 (N_210,In_302,In_339);
nor U211 (N_211,In_204,In_270);
xnor U212 (N_212,In_430,In_243);
nor U213 (N_213,In_61,In_9);
nand U214 (N_214,In_488,In_280);
and U215 (N_215,In_80,In_223);
and U216 (N_216,In_34,In_452);
xnor U217 (N_217,In_425,In_257);
or U218 (N_218,In_259,In_152);
xnor U219 (N_219,In_245,In_258);
nand U220 (N_220,In_360,In_387);
nor U221 (N_221,In_126,In_454);
or U222 (N_222,In_177,In_229);
xor U223 (N_223,In_215,In_132);
xnor U224 (N_224,In_219,In_45);
nand U225 (N_225,In_206,In_32);
or U226 (N_226,In_491,In_143);
xor U227 (N_227,In_122,In_53);
and U228 (N_228,In_14,In_115);
and U229 (N_229,In_87,In_303);
and U230 (N_230,In_414,In_12);
nand U231 (N_231,In_43,In_320);
nor U232 (N_232,In_354,In_50);
nor U233 (N_233,In_442,In_98);
and U234 (N_234,In_42,In_128);
or U235 (N_235,In_447,In_353);
or U236 (N_236,In_406,In_389);
nor U237 (N_237,In_79,In_494);
xnor U238 (N_238,In_104,In_232);
or U239 (N_239,In_261,In_39);
xor U240 (N_240,In_136,In_116);
or U241 (N_241,In_349,In_340);
nor U242 (N_242,In_391,In_437);
xnor U243 (N_243,In_373,In_200);
nor U244 (N_244,In_357,In_218);
nand U245 (N_245,In_356,In_73);
xnor U246 (N_246,In_263,In_287);
and U247 (N_247,In_33,In_36);
or U248 (N_248,In_111,In_369);
nor U249 (N_249,In_405,In_171);
nand U250 (N_250,In_119,In_88);
xnor U251 (N_251,In_282,In_311);
or U252 (N_252,In_73,In_42);
and U253 (N_253,In_465,In_318);
xor U254 (N_254,In_312,In_445);
nor U255 (N_255,In_42,In_396);
or U256 (N_256,In_268,In_254);
or U257 (N_257,In_472,In_216);
nand U258 (N_258,In_408,In_415);
nand U259 (N_259,In_133,In_293);
or U260 (N_260,In_386,In_224);
nor U261 (N_261,In_462,In_155);
and U262 (N_262,In_243,In_410);
and U263 (N_263,In_233,In_107);
nand U264 (N_264,In_351,In_117);
and U265 (N_265,In_489,In_280);
or U266 (N_266,In_84,In_19);
nand U267 (N_267,In_443,In_349);
nor U268 (N_268,In_460,In_448);
or U269 (N_269,In_226,In_211);
nand U270 (N_270,In_296,In_495);
xnor U271 (N_271,In_124,In_79);
nand U272 (N_272,In_213,In_368);
xor U273 (N_273,In_207,In_357);
nand U274 (N_274,In_78,In_281);
xnor U275 (N_275,In_495,In_71);
nor U276 (N_276,In_109,In_135);
xnor U277 (N_277,In_10,In_393);
and U278 (N_278,In_229,In_210);
xor U279 (N_279,In_256,In_401);
nor U280 (N_280,In_278,In_166);
nand U281 (N_281,In_471,In_305);
nand U282 (N_282,In_394,In_90);
nor U283 (N_283,In_483,In_128);
nand U284 (N_284,In_245,In_182);
and U285 (N_285,In_409,In_75);
nor U286 (N_286,In_96,In_370);
nor U287 (N_287,In_28,In_352);
nand U288 (N_288,In_297,In_94);
nand U289 (N_289,In_366,In_256);
nand U290 (N_290,In_315,In_400);
and U291 (N_291,In_474,In_264);
xor U292 (N_292,In_213,In_21);
or U293 (N_293,In_158,In_57);
nor U294 (N_294,In_445,In_11);
or U295 (N_295,In_390,In_477);
and U296 (N_296,In_360,In_263);
and U297 (N_297,In_253,In_492);
xor U298 (N_298,In_300,In_296);
and U299 (N_299,In_229,In_200);
nand U300 (N_300,In_433,In_488);
and U301 (N_301,In_132,In_462);
xor U302 (N_302,In_216,In_161);
nor U303 (N_303,In_326,In_137);
nor U304 (N_304,In_274,In_404);
or U305 (N_305,In_214,In_257);
and U306 (N_306,In_348,In_472);
xor U307 (N_307,In_359,In_30);
nand U308 (N_308,In_385,In_159);
nand U309 (N_309,In_233,In_405);
nand U310 (N_310,In_183,In_289);
nand U311 (N_311,In_321,In_215);
or U312 (N_312,In_367,In_364);
and U313 (N_313,In_388,In_187);
or U314 (N_314,In_50,In_70);
nand U315 (N_315,In_137,In_369);
nand U316 (N_316,In_30,In_489);
nor U317 (N_317,In_326,In_4);
nor U318 (N_318,In_111,In_385);
nor U319 (N_319,In_367,In_162);
nand U320 (N_320,In_46,In_317);
and U321 (N_321,In_259,In_8);
nand U322 (N_322,In_178,In_267);
nand U323 (N_323,In_192,In_155);
nand U324 (N_324,In_472,In_123);
nand U325 (N_325,In_315,In_407);
or U326 (N_326,In_459,In_178);
or U327 (N_327,In_300,In_340);
nor U328 (N_328,In_466,In_102);
nor U329 (N_329,In_113,In_432);
nand U330 (N_330,In_154,In_354);
and U331 (N_331,In_157,In_132);
nor U332 (N_332,In_143,In_371);
and U333 (N_333,In_226,In_483);
nor U334 (N_334,In_186,In_370);
and U335 (N_335,In_16,In_266);
nor U336 (N_336,In_430,In_464);
nand U337 (N_337,In_213,In_398);
xor U338 (N_338,In_69,In_409);
nor U339 (N_339,In_337,In_129);
xor U340 (N_340,In_66,In_51);
xnor U341 (N_341,In_156,In_416);
or U342 (N_342,In_398,In_417);
xor U343 (N_343,In_344,In_215);
nand U344 (N_344,In_17,In_142);
nor U345 (N_345,In_26,In_475);
nor U346 (N_346,In_26,In_77);
or U347 (N_347,In_496,In_103);
or U348 (N_348,In_298,In_428);
or U349 (N_349,In_477,In_412);
xnor U350 (N_350,In_142,In_272);
or U351 (N_351,In_390,In_488);
nor U352 (N_352,In_64,In_302);
nor U353 (N_353,In_206,In_252);
nand U354 (N_354,In_365,In_71);
or U355 (N_355,In_207,In_32);
or U356 (N_356,In_289,In_249);
or U357 (N_357,In_169,In_198);
nor U358 (N_358,In_250,In_31);
xnor U359 (N_359,In_320,In_56);
nand U360 (N_360,In_339,In_476);
and U361 (N_361,In_354,In_232);
nor U362 (N_362,In_125,In_353);
or U363 (N_363,In_34,In_357);
nor U364 (N_364,In_314,In_477);
xor U365 (N_365,In_219,In_294);
nor U366 (N_366,In_270,In_124);
and U367 (N_367,In_471,In_298);
nor U368 (N_368,In_125,In_189);
or U369 (N_369,In_179,In_206);
or U370 (N_370,In_41,In_428);
and U371 (N_371,In_213,In_169);
nor U372 (N_372,In_77,In_165);
xor U373 (N_373,In_424,In_415);
nand U374 (N_374,In_324,In_440);
nand U375 (N_375,In_488,In_338);
nand U376 (N_376,In_462,In_303);
xnor U377 (N_377,In_434,In_126);
and U378 (N_378,In_285,In_449);
nand U379 (N_379,In_261,In_275);
nand U380 (N_380,In_197,In_496);
nor U381 (N_381,In_31,In_124);
and U382 (N_382,In_407,In_242);
or U383 (N_383,In_185,In_351);
nor U384 (N_384,In_336,In_118);
xnor U385 (N_385,In_328,In_109);
and U386 (N_386,In_336,In_218);
and U387 (N_387,In_228,In_15);
xor U388 (N_388,In_3,In_401);
or U389 (N_389,In_246,In_110);
and U390 (N_390,In_127,In_476);
and U391 (N_391,In_9,In_171);
xnor U392 (N_392,In_198,In_385);
and U393 (N_393,In_125,In_208);
or U394 (N_394,In_64,In_122);
or U395 (N_395,In_279,In_143);
xor U396 (N_396,In_462,In_352);
nor U397 (N_397,In_174,In_151);
and U398 (N_398,In_59,In_287);
xor U399 (N_399,In_13,In_11);
or U400 (N_400,In_431,In_418);
or U401 (N_401,In_447,In_426);
xnor U402 (N_402,In_230,In_155);
nor U403 (N_403,In_185,In_236);
nor U404 (N_404,In_417,In_336);
and U405 (N_405,In_213,In_462);
or U406 (N_406,In_351,In_8);
xnor U407 (N_407,In_168,In_414);
xor U408 (N_408,In_304,In_157);
nor U409 (N_409,In_103,In_377);
nor U410 (N_410,In_73,In_441);
or U411 (N_411,In_480,In_97);
xnor U412 (N_412,In_192,In_330);
or U413 (N_413,In_50,In_39);
nand U414 (N_414,In_162,In_342);
and U415 (N_415,In_56,In_21);
nand U416 (N_416,In_203,In_442);
nor U417 (N_417,In_179,In_387);
and U418 (N_418,In_304,In_142);
and U419 (N_419,In_190,In_196);
xor U420 (N_420,In_273,In_472);
nand U421 (N_421,In_23,In_256);
nand U422 (N_422,In_460,In_225);
nor U423 (N_423,In_239,In_356);
and U424 (N_424,In_32,In_130);
nand U425 (N_425,In_440,In_245);
or U426 (N_426,In_413,In_329);
or U427 (N_427,In_263,In_60);
or U428 (N_428,In_309,In_76);
xnor U429 (N_429,In_122,In_447);
nor U430 (N_430,In_104,In_418);
nor U431 (N_431,In_366,In_245);
or U432 (N_432,In_476,In_110);
or U433 (N_433,In_141,In_489);
xor U434 (N_434,In_311,In_283);
and U435 (N_435,In_134,In_33);
and U436 (N_436,In_462,In_172);
xnor U437 (N_437,In_298,In_271);
or U438 (N_438,In_453,In_261);
and U439 (N_439,In_204,In_340);
nor U440 (N_440,In_22,In_148);
nand U441 (N_441,In_246,In_435);
nand U442 (N_442,In_471,In_42);
and U443 (N_443,In_276,In_345);
xor U444 (N_444,In_402,In_386);
nand U445 (N_445,In_347,In_353);
xnor U446 (N_446,In_429,In_473);
xor U447 (N_447,In_336,In_343);
xnor U448 (N_448,In_81,In_19);
xnor U449 (N_449,In_266,In_291);
xnor U450 (N_450,In_417,In_91);
or U451 (N_451,In_325,In_326);
xor U452 (N_452,In_486,In_347);
nand U453 (N_453,In_197,In_173);
nand U454 (N_454,In_210,In_355);
xor U455 (N_455,In_72,In_198);
or U456 (N_456,In_381,In_59);
nand U457 (N_457,In_321,In_310);
or U458 (N_458,In_411,In_125);
nor U459 (N_459,In_462,In_328);
nand U460 (N_460,In_232,In_483);
nor U461 (N_461,In_165,In_80);
nand U462 (N_462,In_372,In_476);
and U463 (N_463,In_203,In_130);
nand U464 (N_464,In_413,In_286);
and U465 (N_465,In_467,In_358);
xor U466 (N_466,In_284,In_137);
and U467 (N_467,In_164,In_191);
and U468 (N_468,In_179,In_38);
nor U469 (N_469,In_371,In_149);
and U470 (N_470,In_448,In_469);
xnor U471 (N_471,In_496,In_204);
or U472 (N_472,In_104,In_219);
nand U473 (N_473,In_96,In_328);
and U474 (N_474,In_419,In_432);
and U475 (N_475,In_39,In_190);
nand U476 (N_476,In_200,In_102);
or U477 (N_477,In_89,In_25);
and U478 (N_478,In_490,In_338);
xor U479 (N_479,In_133,In_186);
or U480 (N_480,In_446,In_23);
xnor U481 (N_481,In_498,In_279);
nand U482 (N_482,In_469,In_311);
nand U483 (N_483,In_455,In_356);
or U484 (N_484,In_157,In_22);
nand U485 (N_485,In_73,In_113);
xor U486 (N_486,In_462,In_483);
or U487 (N_487,In_316,In_297);
and U488 (N_488,In_138,In_107);
xnor U489 (N_489,In_275,In_245);
or U490 (N_490,In_415,In_491);
or U491 (N_491,In_177,In_198);
or U492 (N_492,In_361,In_271);
and U493 (N_493,In_303,In_387);
and U494 (N_494,In_208,In_428);
xor U495 (N_495,In_314,In_52);
and U496 (N_496,In_35,In_214);
nor U497 (N_497,In_144,In_38);
nand U498 (N_498,In_326,In_15);
nand U499 (N_499,In_364,In_223);
nor U500 (N_500,N_341,N_415);
or U501 (N_501,N_244,N_5);
nor U502 (N_502,N_405,N_272);
or U503 (N_503,N_306,N_419);
and U504 (N_504,N_39,N_497);
xor U505 (N_505,N_69,N_398);
and U506 (N_506,N_423,N_162);
or U507 (N_507,N_265,N_120);
xnor U508 (N_508,N_133,N_197);
xor U509 (N_509,N_414,N_212);
nor U510 (N_510,N_470,N_187);
nand U511 (N_511,N_79,N_492);
or U512 (N_512,N_125,N_234);
and U513 (N_513,N_377,N_61);
xnor U514 (N_514,N_2,N_116);
xnor U515 (N_515,N_150,N_432);
nor U516 (N_516,N_13,N_314);
xnor U517 (N_517,N_238,N_219);
nor U518 (N_518,N_413,N_337);
nor U519 (N_519,N_445,N_358);
and U520 (N_520,N_29,N_294);
or U521 (N_521,N_335,N_329);
or U522 (N_522,N_364,N_57);
xor U523 (N_523,N_453,N_394);
and U524 (N_524,N_190,N_17);
or U525 (N_525,N_312,N_87);
and U526 (N_526,N_449,N_235);
nor U527 (N_527,N_40,N_360);
nor U528 (N_528,N_399,N_457);
or U529 (N_529,N_9,N_33);
xor U530 (N_530,N_357,N_147);
nor U531 (N_531,N_459,N_195);
or U532 (N_532,N_319,N_223);
nor U533 (N_533,N_383,N_259);
nand U534 (N_534,N_436,N_417);
or U535 (N_535,N_282,N_151);
and U536 (N_536,N_22,N_11);
and U537 (N_537,N_28,N_209);
nand U538 (N_538,N_482,N_172);
or U539 (N_539,N_305,N_281);
nor U540 (N_540,N_455,N_88);
or U541 (N_541,N_300,N_160);
or U542 (N_542,N_480,N_134);
nand U543 (N_543,N_217,N_85);
nor U544 (N_544,N_117,N_372);
xor U545 (N_545,N_82,N_481);
nand U546 (N_546,N_468,N_443);
xnor U547 (N_547,N_205,N_166);
or U548 (N_548,N_58,N_253);
nand U549 (N_549,N_80,N_288);
and U550 (N_550,N_277,N_107);
nand U551 (N_551,N_71,N_437);
xor U552 (N_552,N_220,N_291);
and U553 (N_553,N_233,N_246);
or U554 (N_554,N_466,N_226);
and U555 (N_555,N_0,N_90);
nand U556 (N_556,N_189,N_10);
nand U557 (N_557,N_431,N_173);
or U558 (N_558,N_31,N_157);
and U559 (N_559,N_152,N_324);
nor U560 (N_560,N_274,N_193);
or U561 (N_561,N_355,N_68);
xnor U562 (N_562,N_370,N_304);
and U563 (N_563,N_179,N_106);
or U564 (N_564,N_263,N_483);
xnor U565 (N_565,N_137,N_261);
xnor U566 (N_566,N_180,N_119);
nor U567 (N_567,N_342,N_339);
and U568 (N_568,N_51,N_317);
nand U569 (N_569,N_178,N_241);
or U570 (N_570,N_269,N_429);
xnor U571 (N_571,N_391,N_138);
nor U572 (N_572,N_289,N_47);
or U573 (N_573,N_290,N_237);
or U574 (N_574,N_462,N_46);
xnor U575 (N_575,N_451,N_471);
nor U576 (N_576,N_174,N_73);
or U577 (N_577,N_34,N_109);
nor U578 (N_578,N_280,N_258);
nand U579 (N_579,N_296,N_77);
and U580 (N_580,N_322,N_21);
nand U581 (N_581,N_487,N_444);
and U582 (N_582,N_43,N_307);
nor U583 (N_583,N_385,N_256);
xor U584 (N_584,N_115,N_362);
nand U585 (N_585,N_126,N_93);
nor U586 (N_586,N_262,N_315);
and U587 (N_587,N_176,N_97);
nor U588 (N_588,N_32,N_194);
nor U589 (N_589,N_206,N_141);
or U590 (N_590,N_225,N_203);
nand U591 (N_591,N_59,N_389);
or U592 (N_592,N_363,N_128);
nor U593 (N_593,N_36,N_334);
nor U594 (N_594,N_236,N_214);
and U595 (N_595,N_245,N_308);
xnor U596 (N_596,N_316,N_440);
nand U597 (N_597,N_418,N_165);
xnor U598 (N_598,N_49,N_456);
xnor U599 (N_599,N_143,N_113);
or U600 (N_600,N_401,N_379);
and U601 (N_601,N_472,N_346);
or U602 (N_602,N_38,N_284);
or U603 (N_603,N_154,N_396);
or U604 (N_604,N_145,N_421);
and U605 (N_605,N_121,N_325);
nand U606 (N_606,N_331,N_359);
nor U607 (N_607,N_309,N_433);
xor U608 (N_608,N_376,N_386);
xor U609 (N_609,N_250,N_295);
or U610 (N_610,N_375,N_227);
nor U611 (N_611,N_146,N_55);
and U612 (N_612,N_397,N_321);
nand U613 (N_613,N_81,N_345);
or U614 (N_614,N_404,N_131);
or U615 (N_615,N_380,N_19);
xor U616 (N_616,N_279,N_495);
and U617 (N_617,N_177,N_169);
nor U618 (N_618,N_467,N_438);
nor U619 (N_619,N_100,N_124);
and U620 (N_620,N_276,N_76);
xnor U621 (N_621,N_350,N_153);
and U622 (N_622,N_243,N_488);
xnor U623 (N_623,N_491,N_102);
and U624 (N_624,N_273,N_249);
or U625 (N_625,N_287,N_349);
or U626 (N_626,N_252,N_328);
and U627 (N_627,N_8,N_84);
nand U628 (N_628,N_23,N_412);
xor U629 (N_629,N_320,N_27);
or U630 (N_630,N_452,N_353);
nand U631 (N_631,N_278,N_460);
xor U632 (N_632,N_30,N_94);
xor U633 (N_633,N_148,N_446);
or U634 (N_634,N_230,N_201);
xor U635 (N_635,N_298,N_101);
or U636 (N_636,N_275,N_213);
or U637 (N_637,N_499,N_479);
nor U638 (N_638,N_183,N_493);
or U639 (N_639,N_387,N_257);
nor U640 (N_640,N_163,N_50);
xor U641 (N_641,N_411,N_367);
nand U642 (N_642,N_198,N_292);
nand U643 (N_643,N_222,N_425);
or U644 (N_644,N_62,N_254);
nor U645 (N_645,N_476,N_208);
nand U646 (N_646,N_98,N_78);
xnor U647 (N_647,N_112,N_407);
xor U648 (N_648,N_229,N_477);
or U649 (N_649,N_310,N_142);
or U650 (N_650,N_330,N_108);
xor U651 (N_651,N_374,N_303);
or U652 (N_652,N_105,N_6);
nand U653 (N_653,N_323,N_168);
and U654 (N_654,N_104,N_53);
or U655 (N_655,N_442,N_25);
nand U656 (N_656,N_484,N_326);
or U657 (N_657,N_388,N_301);
or U658 (N_658,N_188,N_140);
or U659 (N_659,N_318,N_130);
nand U660 (N_660,N_454,N_224);
nor U661 (N_661,N_155,N_132);
and U662 (N_662,N_490,N_373);
xor U663 (N_663,N_75,N_378);
xor U664 (N_664,N_199,N_494);
nand U665 (N_665,N_416,N_381);
nor U666 (N_666,N_204,N_384);
or U667 (N_667,N_16,N_408);
or U668 (N_668,N_486,N_352);
and U669 (N_669,N_67,N_35);
nand U670 (N_670,N_65,N_103);
or U671 (N_671,N_285,N_450);
nor U672 (N_672,N_463,N_406);
or U673 (N_673,N_403,N_156);
and U674 (N_674,N_332,N_45);
nor U675 (N_675,N_458,N_158);
nand U676 (N_676,N_343,N_149);
nor U677 (N_677,N_207,N_283);
xnor U678 (N_678,N_336,N_186);
or U679 (N_679,N_139,N_302);
xnor U680 (N_680,N_369,N_420);
or U681 (N_681,N_351,N_422);
xor U682 (N_682,N_286,N_371);
and U683 (N_683,N_266,N_465);
and U684 (N_684,N_247,N_251);
nand U685 (N_685,N_340,N_441);
nand U686 (N_686,N_313,N_248);
or U687 (N_687,N_231,N_240);
nor U688 (N_688,N_135,N_70);
or U689 (N_689,N_184,N_327);
nor U690 (N_690,N_448,N_12);
or U691 (N_691,N_293,N_167);
nand U692 (N_692,N_232,N_159);
xnor U693 (N_693,N_26,N_48);
xnor U694 (N_694,N_56,N_3);
or U695 (N_695,N_42,N_427);
nor U696 (N_696,N_161,N_64);
xnor U697 (N_697,N_366,N_118);
xnor U698 (N_698,N_368,N_347);
nand U699 (N_699,N_338,N_164);
nand U700 (N_700,N_37,N_299);
nand U701 (N_701,N_297,N_83);
nand U702 (N_702,N_409,N_424);
nor U703 (N_703,N_72,N_410);
nor U704 (N_704,N_260,N_475);
nor U705 (N_705,N_171,N_99);
or U706 (N_706,N_15,N_255);
and U707 (N_707,N_18,N_434);
nor U708 (N_708,N_63,N_392);
or U709 (N_709,N_239,N_192);
nor U710 (N_710,N_464,N_181);
or U711 (N_711,N_91,N_54);
or U712 (N_712,N_202,N_430);
or U713 (N_713,N_344,N_439);
and U714 (N_714,N_182,N_210);
nor U715 (N_715,N_242,N_110);
or U716 (N_716,N_136,N_426);
or U717 (N_717,N_400,N_478);
nor U718 (N_718,N_127,N_74);
nand U719 (N_719,N_185,N_14);
and U720 (N_720,N_221,N_24);
nor U721 (N_721,N_41,N_218);
nand U722 (N_722,N_4,N_393);
nor U723 (N_723,N_60,N_111);
or U724 (N_724,N_485,N_365);
and U725 (N_725,N_216,N_489);
xnor U726 (N_726,N_96,N_271);
nor U727 (N_727,N_122,N_123);
nand U728 (N_728,N_356,N_170);
nor U729 (N_729,N_270,N_447);
nor U730 (N_730,N_348,N_311);
or U731 (N_731,N_435,N_228);
xnor U732 (N_732,N_1,N_200);
xnor U733 (N_733,N_395,N_402);
xnor U734 (N_734,N_333,N_382);
xor U735 (N_735,N_354,N_66);
and U736 (N_736,N_114,N_175);
and U737 (N_737,N_496,N_267);
and U738 (N_738,N_92,N_390);
and U739 (N_739,N_191,N_361);
nor U740 (N_740,N_469,N_428);
or U741 (N_741,N_461,N_215);
or U742 (N_742,N_474,N_86);
or U743 (N_743,N_264,N_7);
nor U744 (N_744,N_498,N_89);
or U745 (N_745,N_473,N_44);
or U746 (N_746,N_95,N_20);
nand U747 (N_747,N_144,N_52);
and U748 (N_748,N_129,N_211);
nand U749 (N_749,N_268,N_196);
nand U750 (N_750,N_1,N_475);
nor U751 (N_751,N_40,N_2);
nor U752 (N_752,N_51,N_494);
xor U753 (N_753,N_139,N_397);
nand U754 (N_754,N_152,N_140);
nand U755 (N_755,N_80,N_274);
nor U756 (N_756,N_254,N_391);
or U757 (N_757,N_96,N_492);
or U758 (N_758,N_364,N_427);
nor U759 (N_759,N_337,N_116);
or U760 (N_760,N_140,N_252);
or U761 (N_761,N_186,N_377);
or U762 (N_762,N_423,N_398);
nor U763 (N_763,N_181,N_437);
or U764 (N_764,N_418,N_178);
nand U765 (N_765,N_371,N_405);
nand U766 (N_766,N_317,N_288);
nand U767 (N_767,N_413,N_88);
xor U768 (N_768,N_477,N_192);
nand U769 (N_769,N_192,N_483);
xnor U770 (N_770,N_125,N_77);
nand U771 (N_771,N_231,N_333);
or U772 (N_772,N_212,N_331);
or U773 (N_773,N_129,N_374);
or U774 (N_774,N_100,N_193);
nor U775 (N_775,N_44,N_286);
and U776 (N_776,N_16,N_116);
or U777 (N_777,N_176,N_106);
xnor U778 (N_778,N_350,N_152);
nand U779 (N_779,N_318,N_362);
and U780 (N_780,N_360,N_211);
nand U781 (N_781,N_110,N_471);
and U782 (N_782,N_162,N_451);
or U783 (N_783,N_14,N_217);
nor U784 (N_784,N_151,N_448);
and U785 (N_785,N_471,N_372);
nor U786 (N_786,N_208,N_90);
and U787 (N_787,N_27,N_142);
xnor U788 (N_788,N_145,N_471);
or U789 (N_789,N_30,N_137);
xor U790 (N_790,N_0,N_191);
nand U791 (N_791,N_232,N_99);
nand U792 (N_792,N_410,N_152);
and U793 (N_793,N_98,N_55);
or U794 (N_794,N_7,N_10);
or U795 (N_795,N_308,N_410);
and U796 (N_796,N_121,N_317);
nor U797 (N_797,N_42,N_294);
or U798 (N_798,N_462,N_144);
and U799 (N_799,N_389,N_422);
and U800 (N_800,N_340,N_466);
nand U801 (N_801,N_197,N_336);
or U802 (N_802,N_243,N_224);
and U803 (N_803,N_141,N_446);
and U804 (N_804,N_46,N_345);
nand U805 (N_805,N_317,N_384);
or U806 (N_806,N_82,N_288);
xor U807 (N_807,N_50,N_460);
nand U808 (N_808,N_131,N_381);
and U809 (N_809,N_448,N_178);
nor U810 (N_810,N_384,N_402);
or U811 (N_811,N_420,N_251);
and U812 (N_812,N_14,N_295);
or U813 (N_813,N_283,N_477);
nor U814 (N_814,N_391,N_479);
nand U815 (N_815,N_473,N_113);
nand U816 (N_816,N_51,N_281);
nor U817 (N_817,N_255,N_498);
nor U818 (N_818,N_486,N_224);
xnor U819 (N_819,N_80,N_441);
xnor U820 (N_820,N_337,N_358);
or U821 (N_821,N_353,N_223);
and U822 (N_822,N_289,N_351);
nor U823 (N_823,N_251,N_54);
nand U824 (N_824,N_356,N_74);
and U825 (N_825,N_152,N_184);
nor U826 (N_826,N_133,N_388);
xnor U827 (N_827,N_344,N_186);
nor U828 (N_828,N_402,N_125);
nand U829 (N_829,N_381,N_151);
and U830 (N_830,N_429,N_295);
nor U831 (N_831,N_374,N_85);
and U832 (N_832,N_14,N_245);
nand U833 (N_833,N_194,N_449);
or U834 (N_834,N_225,N_108);
xnor U835 (N_835,N_477,N_27);
nand U836 (N_836,N_89,N_54);
nor U837 (N_837,N_369,N_340);
and U838 (N_838,N_150,N_489);
nor U839 (N_839,N_224,N_388);
and U840 (N_840,N_455,N_106);
xnor U841 (N_841,N_321,N_383);
nor U842 (N_842,N_240,N_196);
nand U843 (N_843,N_55,N_121);
nor U844 (N_844,N_366,N_159);
or U845 (N_845,N_428,N_59);
nand U846 (N_846,N_45,N_396);
nand U847 (N_847,N_498,N_48);
nand U848 (N_848,N_187,N_494);
xnor U849 (N_849,N_49,N_446);
nor U850 (N_850,N_267,N_464);
xnor U851 (N_851,N_179,N_34);
and U852 (N_852,N_126,N_433);
and U853 (N_853,N_499,N_370);
xnor U854 (N_854,N_89,N_35);
nand U855 (N_855,N_198,N_128);
xnor U856 (N_856,N_420,N_344);
nand U857 (N_857,N_189,N_413);
nand U858 (N_858,N_351,N_1);
or U859 (N_859,N_234,N_176);
nand U860 (N_860,N_337,N_138);
xnor U861 (N_861,N_88,N_248);
nor U862 (N_862,N_7,N_80);
xor U863 (N_863,N_475,N_257);
nor U864 (N_864,N_330,N_273);
xor U865 (N_865,N_387,N_144);
and U866 (N_866,N_253,N_454);
or U867 (N_867,N_101,N_435);
xnor U868 (N_868,N_125,N_294);
and U869 (N_869,N_266,N_297);
and U870 (N_870,N_342,N_208);
and U871 (N_871,N_457,N_198);
nand U872 (N_872,N_360,N_83);
nor U873 (N_873,N_268,N_475);
nand U874 (N_874,N_154,N_421);
and U875 (N_875,N_384,N_409);
and U876 (N_876,N_397,N_388);
and U877 (N_877,N_351,N_297);
nand U878 (N_878,N_82,N_491);
nor U879 (N_879,N_358,N_369);
nor U880 (N_880,N_231,N_338);
xor U881 (N_881,N_154,N_119);
and U882 (N_882,N_371,N_339);
xnor U883 (N_883,N_1,N_138);
xnor U884 (N_884,N_445,N_328);
xor U885 (N_885,N_187,N_343);
and U886 (N_886,N_442,N_87);
nand U887 (N_887,N_467,N_318);
and U888 (N_888,N_393,N_109);
nor U889 (N_889,N_67,N_375);
xor U890 (N_890,N_246,N_426);
xnor U891 (N_891,N_466,N_5);
and U892 (N_892,N_415,N_309);
or U893 (N_893,N_304,N_332);
and U894 (N_894,N_58,N_242);
and U895 (N_895,N_278,N_462);
nor U896 (N_896,N_419,N_185);
and U897 (N_897,N_270,N_318);
xnor U898 (N_898,N_56,N_270);
or U899 (N_899,N_167,N_349);
and U900 (N_900,N_364,N_497);
and U901 (N_901,N_0,N_203);
and U902 (N_902,N_457,N_119);
nor U903 (N_903,N_374,N_386);
nand U904 (N_904,N_219,N_156);
or U905 (N_905,N_329,N_141);
or U906 (N_906,N_42,N_219);
xnor U907 (N_907,N_126,N_171);
and U908 (N_908,N_125,N_348);
or U909 (N_909,N_263,N_89);
nand U910 (N_910,N_24,N_425);
nand U911 (N_911,N_449,N_23);
or U912 (N_912,N_167,N_392);
nor U913 (N_913,N_233,N_370);
xor U914 (N_914,N_476,N_457);
xor U915 (N_915,N_247,N_132);
xnor U916 (N_916,N_467,N_420);
xnor U917 (N_917,N_187,N_58);
and U918 (N_918,N_305,N_269);
nand U919 (N_919,N_218,N_476);
nor U920 (N_920,N_238,N_168);
nand U921 (N_921,N_203,N_324);
nand U922 (N_922,N_110,N_171);
xor U923 (N_923,N_312,N_305);
and U924 (N_924,N_225,N_236);
or U925 (N_925,N_214,N_241);
xor U926 (N_926,N_29,N_451);
nor U927 (N_927,N_125,N_23);
or U928 (N_928,N_177,N_379);
and U929 (N_929,N_422,N_234);
nor U930 (N_930,N_12,N_410);
or U931 (N_931,N_188,N_294);
and U932 (N_932,N_170,N_239);
and U933 (N_933,N_59,N_422);
xnor U934 (N_934,N_149,N_189);
nor U935 (N_935,N_475,N_493);
nand U936 (N_936,N_60,N_454);
xor U937 (N_937,N_250,N_205);
xnor U938 (N_938,N_90,N_244);
nor U939 (N_939,N_345,N_397);
nor U940 (N_940,N_182,N_310);
xor U941 (N_941,N_16,N_18);
xnor U942 (N_942,N_384,N_126);
and U943 (N_943,N_209,N_140);
xor U944 (N_944,N_409,N_174);
nor U945 (N_945,N_466,N_402);
or U946 (N_946,N_266,N_477);
or U947 (N_947,N_232,N_347);
or U948 (N_948,N_95,N_485);
nor U949 (N_949,N_322,N_189);
or U950 (N_950,N_94,N_296);
or U951 (N_951,N_24,N_443);
nor U952 (N_952,N_410,N_311);
and U953 (N_953,N_254,N_379);
or U954 (N_954,N_472,N_189);
nor U955 (N_955,N_478,N_301);
nor U956 (N_956,N_359,N_196);
and U957 (N_957,N_52,N_124);
nand U958 (N_958,N_497,N_295);
xnor U959 (N_959,N_264,N_184);
or U960 (N_960,N_113,N_138);
and U961 (N_961,N_278,N_480);
or U962 (N_962,N_488,N_468);
and U963 (N_963,N_324,N_130);
nor U964 (N_964,N_388,N_72);
nor U965 (N_965,N_21,N_361);
xnor U966 (N_966,N_256,N_250);
or U967 (N_967,N_368,N_221);
and U968 (N_968,N_253,N_265);
or U969 (N_969,N_477,N_321);
xnor U970 (N_970,N_329,N_343);
nor U971 (N_971,N_237,N_327);
and U972 (N_972,N_364,N_188);
nand U973 (N_973,N_380,N_182);
nand U974 (N_974,N_164,N_98);
and U975 (N_975,N_303,N_124);
or U976 (N_976,N_241,N_22);
and U977 (N_977,N_103,N_46);
xnor U978 (N_978,N_298,N_316);
xnor U979 (N_979,N_138,N_26);
and U980 (N_980,N_23,N_290);
nand U981 (N_981,N_388,N_452);
xnor U982 (N_982,N_163,N_128);
or U983 (N_983,N_233,N_373);
xnor U984 (N_984,N_166,N_270);
and U985 (N_985,N_398,N_327);
nand U986 (N_986,N_281,N_225);
or U987 (N_987,N_293,N_44);
xnor U988 (N_988,N_243,N_352);
nand U989 (N_989,N_102,N_62);
or U990 (N_990,N_454,N_357);
or U991 (N_991,N_322,N_57);
and U992 (N_992,N_379,N_430);
nor U993 (N_993,N_260,N_410);
or U994 (N_994,N_143,N_197);
and U995 (N_995,N_67,N_430);
nand U996 (N_996,N_138,N_41);
nor U997 (N_997,N_211,N_118);
nand U998 (N_998,N_214,N_32);
nand U999 (N_999,N_217,N_219);
and U1000 (N_1000,N_530,N_548);
nand U1001 (N_1001,N_696,N_925);
nand U1002 (N_1002,N_845,N_730);
or U1003 (N_1003,N_950,N_968);
and U1004 (N_1004,N_616,N_989);
and U1005 (N_1005,N_524,N_589);
nand U1006 (N_1006,N_573,N_533);
nor U1007 (N_1007,N_677,N_992);
and U1008 (N_1008,N_579,N_802);
nand U1009 (N_1009,N_654,N_863);
and U1010 (N_1010,N_706,N_617);
or U1011 (N_1011,N_581,N_927);
nor U1012 (N_1012,N_598,N_737);
xor U1013 (N_1013,N_745,N_621);
nand U1014 (N_1014,N_751,N_701);
or U1015 (N_1015,N_874,N_897);
nand U1016 (N_1016,N_661,N_886);
or U1017 (N_1017,N_994,N_972);
nand U1018 (N_1018,N_903,N_881);
nand U1019 (N_1019,N_712,N_645);
and U1020 (N_1020,N_791,N_952);
nor U1021 (N_1021,N_595,N_719);
nand U1022 (N_1022,N_642,N_918);
and U1023 (N_1023,N_669,N_640);
nor U1024 (N_1024,N_859,N_883);
and U1025 (N_1025,N_671,N_851);
xor U1026 (N_1026,N_867,N_539);
and U1027 (N_1027,N_762,N_838);
and U1028 (N_1028,N_656,N_861);
xor U1029 (N_1029,N_767,N_537);
or U1030 (N_1030,N_856,N_770);
and U1031 (N_1031,N_592,N_754);
xor U1032 (N_1032,N_603,N_519);
nand U1033 (N_1033,N_775,N_766);
nor U1034 (N_1034,N_890,N_674);
or U1035 (N_1035,N_700,N_778);
and U1036 (N_1036,N_790,N_545);
nor U1037 (N_1037,N_864,N_527);
nand U1038 (N_1038,N_878,N_833);
and U1039 (N_1039,N_752,N_765);
nor U1040 (N_1040,N_872,N_714);
or U1041 (N_1041,N_967,N_917);
nor U1042 (N_1042,N_792,N_964);
and U1043 (N_1043,N_943,N_866);
nor U1044 (N_1044,N_902,N_514);
and U1045 (N_1045,N_865,N_783);
and U1046 (N_1046,N_963,N_831);
nor U1047 (N_1047,N_815,N_882);
and U1048 (N_1048,N_977,N_538);
nand U1049 (N_1049,N_909,N_504);
nand U1050 (N_1050,N_522,N_687);
nor U1051 (N_1051,N_782,N_824);
or U1052 (N_1052,N_532,N_574);
xnor U1053 (N_1053,N_715,N_975);
or U1054 (N_1054,N_697,N_776);
or U1055 (N_1055,N_772,N_505);
xor U1056 (N_1056,N_500,N_551);
nand U1057 (N_1057,N_871,N_544);
or U1058 (N_1058,N_542,N_996);
or U1059 (N_1059,N_608,N_755);
or U1060 (N_1060,N_857,N_625);
nor U1061 (N_1061,N_836,N_686);
xor U1062 (N_1062,N_716,N_613);
nor U1063 (N_1063,N_921,N_508);
nor U1064 (N_1064,N_912,N_810);
xor U1065 (N_1065,N_502,N_931);
and U1066 (N_1066,N_757,N_868);
nand U1067 (N_1067,N_717,N_675);
and U1068 (N_1068,N_954,N_819);
nand U1069 (N_1069,N_988,N_799);
xor U1070 (N_1070,N_982,N_736);
nor U1071 (N_1071,N_667,N_713);
and U1072 (N_1072,N_584,N_554);
nor U1073 (N_1073,N_895,N_690);
nand U1074 (N_1074,N_536,N_681);
nor U1075 (N_1075,N_711,N_729);
or U1076 (N_1076,N_721,N_764);
nand U1077 (N_1077,N_528,N_743);
nand U1078 (N_1078,N_748,N_550);
nor U1079 (N_1079,N_614,N_699);
xnor U1080 (N_1080,N_834,N_797);
xor U1081 (N_1081,N_892,N_571);
nand U1082 (N_1082,N_884,N_920);
nand U1083 (N_1083,N_945,N_905);
nor U1084 (N_1084,N_855,N_786);
or U1085 (N_1085,N_956,N_801);
or U1086 (N_1086,N_893,N_606);
xor U1087 (N_1087,N_602,N_984);
nand U1088 (N_1088,N_873,N_683);
or U1089 (N_1089,N_807,N_814);
nor U1090 (N_1090,N_685,N_796);
xor U1091 (N_1091,N_900,N_568);
or U1092 (N_1092,N_846,N_987);
xor U1093 (N_1093,N_973,N_788);
nor U1094 (N_1094,N_942,N_941);
nor U1095 (N_1095,N_818,N_566);
xor U1096 (N_1096,N_590,N_709);
xor U1097 (N_1097,N_969,N_812);
and U1098 (N_1098,N_657,N_822);
nand U1099 (N_1099,N_580,N_634);
xnor U1100 (N_1100,N_756,N_933);
or U1101 (N_1101,N_628,N_887);
nand U1102 (N_1102,N_708,N_673);
nand U1103 (N_1103,N_948,N_885);
nand U1104 (N_1104,N_665,N_728);
nand U1105 (N_1105,N_844,N_959);
nand U1106 (N_1106,N_516,N_911);
or U1107 (N_1107,N_596,N_535);
and U1108 (N_1108,N_995,N_820);
or U1109 (N_1109,N_780,N_576);
or U1110 (N_1110,N_561,N_825);
nand U1111 (N_1111,N_841,N_908);
nor U1112 (N_1112,N_849,N_618);
nor U1113 (N_1113,N_720,N_759);
or U1114 (N_1114,N_922,N_585);
and U1115 (N_1115,N_693,N_901);
nor U1116 (N_1116,N_727,N_644);
xnor U1117 (N_1117,N_928,N_787);
and U1118 (N_1118,N_733,N_806);
and U1119 (N_1119,N_934,N_553);
and U1120 (N_1120,N_785,N_875);
nand U1121 (N_1121,N_541,N_501);
xor U1122 (N_1122,N_993,N_939);
nand U1123 (N_1123,N_774,N_682);
nand U1124 (N_1124,N_830,N_623);
or U1125 (N_1125,N_880,N_958);
and U1126 (N_1126,N_803,N_676);
or U1127 (N_1127,N_662,N_924);
xor U1128 (N_1128,N_643,N_735);
nor U1129 (N_1129,N_991,N_888);
and U1130 (N_1130,N_529,N_732);
nor U1131 (N_1131,N_929,N_965);
xnor U1132 (N_1132,N_672,N_947);
nor U1133 (N_1133,N_837,N_570);
nor U1134 (N_1134,N_930,N_639);
xor U1135 (N_1135,N_666,N_773);
nor U1136 (N_1136,N_702,N_913);
xnor U1137 (N_1137,N_688,N_558);
nand U1138 (N_1138,N_997,N_839);
nand U1139 (N_1139,N_694,N_670);
nand U1140 (N_1140,N_817,N_986);
nor U1141 (N_1141,N_649,N_562);
nand U1142 (N_1142,N_549,N_919);
and U1143 (N_1143,N_813,N_763);
nand U1144 (N_1144,N_646,N_635);
or U1145 (N_1145,N_559,N_705);
xnor U1146 (N_1146,N_509,N_985);
nand U1147 (N_1147,N_891,N_794);
and U1148 (N_1148,N_604,N_899);
nand U1149 (N_1149,N_840,N_843);
xor U1150 (N_1150,N_718,N_511);
nand U1151 (N_1151,N_594,N_605);
and U1152 (N_1152,N_907,N_915);
nor U1153 (N_1153,N_970,N_546);
nor U1154 (N_1154,N_842,N_703);
nor U1155 (N_1155,N_607,N_655);
xor U1156 (N_1156,N_599,N_565);
nor U1157 (N_1157,N_974,N_938);
or U1158 (N_1158,N_805,N_789);
nor U1159 (N_1159,N_629,N_591);
xnor U1160 (N_1160,N_521,N_914);
or U1161 (N_1161,N_771,N_575);
and U1162 (N_1162,N_684,N_932);
and U1163 (N_1163,N_534,N_858);
or U1164 (N_1164,N_650,N_531);
nor U1165 (N_1165,N_653,N_999);
nor U1166 (N_1166,N_626,N_513);
nor U1167 (N_1167,N_978,N_853);
nor U1168 (N_1168,N_746,N_567);
or U1169 (N_1169,N_707,N_946);
nor U1170 (N_1170,N_641,N_692);
nand U1171 (N_1171,N_647,N_648);
xnor U1172 (N_1172,N_808,N_829);
nand U1173 (N_1173,N_704,N_937);
xor U1174 (N_1174,N_523,N_557);
and U1175 (N_1175,N_747,N_510);
and U1176 (N_1176,N_652,N_633);
and U1177 (N_1177,N_503,N_753);
nor U1178 (N_1178,N_740,N_760);
or U1179 (N_1179,N_798,N_577);
or U1180 (N_1180,N_739,N_896);
nand U1181 (N_1181,N_777,N_940);
xor U1182 (N_1182,N_971,N_660);
nor U1183 (N_1183,N_800,N_862);
or U1184 (N_1184,N_586,N_722);
or U1185 (N_1185,N_741,N_935);
xor U1186 (N_1186,N_569,N_587);
nor U1187 (N_1187,N_651,N_520);
nor U1188 (N_1188,N_877,N_710);
nand U1189 (N_1189,N_638,N_744);
nand U1190 (N_1190,N_609,N_816);
and U1191 (N_1191,N_601,N_957);
nor U1192 (N_1192,N_979,N_784);
xnor U1193 (N_1193,N_560,N_906);
and U1194 (N_1194,N_506,N_734);
xnor U1195 (N_1195,N_981,N_870);
and U1196 (N_1196,N_889,N_552);
and U1197 (N_1197,N_582,N_852);
xnor U1198 (N_1198,N_564,N_679);
and U1199 (N_1199,N_526,N_726);
nand U1200 (N_1200,N_795,N_811);
and U1201 (N_1201,N_611,N_898);
xor U1202 (N_1202,N_738,N_749);
nor U1203 (N_1203,N_725,N_556);
or U1204 (N_1204,N_593,N_615);
xor U1205 (N_1205,N_678,N_949);
and U1206 (N_1206,N_953,N_876);
xnor U1207 (N_1207,N_691,N_622);
xnor U1208 (N_1208,N_944,N_632);
or U1209 (N_1209,N_512,N_804);
and U1210 (N_1210,N_631,N_624);
or U1211 (N_1211,N_998,N_976);
xor U1212 (N_1212,N_980,N_779);
and U1213 (N_1213,N_961,N_904);
nand U1214 (N_1214,N_809,N_854);
xor U1215 (N_1215,N_698,N_894);
nand U1216 (N_1216,N_731,N_983);
and U1217 (N_1217,N_630,N_723);
nor U1218 (N_1218,N_847,N_835);
xor U1219 (N_1219,N_768,N_627);
nand U1220 (N_1220,N_636,N_563);
xor U1221 (N_1221,N_695,N_724);
or U1222 (N_1222,N_664,N_600);
xnor U1223 (N_1223,N_781,N_823);
nand U1224 (N_1224,N_826,N_689);
xor U1225 (N_1225,N_518,N_620);
and U1226 (N_1226,N_850,N_821);
nand U1227 (N_1227,N_583,N_990);
nor U1228 (N_1228,N_610,N_793);
nand U1229 (N_1229,N_955,N_555);
xor U1230 (N_1230,N_543,N_619);
or U1231 (N_1231,N_879,N_926);
or U1232 (N_1232,N_750,N_525);
or U1233 (N_1233,N_761,N_916);
or U1234 (N_1234,N_860,N_517);
or U1235 (N_1235,N_578,N_848);
nor U1236 (N_1236,N_588,N_612);
nand U1237 (N_1237,N_663,N_966);
nand U1238 (N_1238,N_758,N_827);
or U1239 (N_1239,N_910,N_572);
and U1240 (N_1240,N_951,N_540);
nor U1241 (N_1241,N_828,N_507);
xor U1242 (N_1242,N_547,N_659);
nand U1243 (N_1243,N_832,N_668);
or U1244 (N_1244,N_637,N_923);
nand U1245 (N_1245,N_658,N_962);
xor U1246 (N_1246,N_960,N_769);
nor U1247 (N_1247,N_680,N_597);
nand U1248 (N_1248,N_742,N_869);
xnor U1249 (N_1249,N_515,N_936);
or U1250 (N_1250,N_778,N_853);
nor U1251 (N_1251,N_942,N_743);
nand U1252 (N_1252,N_532,N_997);
and U1253 (N_1253,N_757,N_690);
or U1254 (N_1254,N_695,N_889);
or U1255 (N_1255,N_532,N_979);
and U1256 (N_1256,N_580,N_584);
and U1257 (N_1257,N_888,N_900);
xor U1258 (N_1258,N_714,N_678);
or U1259 (N_1259,N_676,N_768);
and U1260 (N_1260,N_902,N_946);
or U1261 (N_1261,N_562,N_924);
and U1262 (N_1262,N_543,N_712);
or U1263 (N_1263,N_967,N_641);
xnor U1264 (N_1264,N_553,N_841);
nor U1265 (N_1265,N_628,N_764);
or U1266 (N_1266,N_744,N_551);
xor U1267 (N_1267,N_984,N_519);
nand U1268 (N_1268,N_645,N_976);
nor U1269 (N_1269,N_865,N_941);
nor U1270 (N_1270,N_513,N_551);
xnor U1271 (N_1271,N_731,N_840);
xnor U1272 (N_1272,N_552,N_996);
nor U1273 (N_1273,N_690,N_584);
xor U1274 (N_1274,N_834,N_558);
or U1275 (N_1275,N_877,N_533);
nand U1276 (N_1276,N_628,N_860);
or U1277 (N_1277,N_658,N_748);
xor U1278 (N_1278,N_664,N_687);
and U1279 (N_1279,N_947,N_744);
and U1280 (N_1280,N_723,N_825);
nand U1281 (N_1281,N_651,N_727);
nor U1282 (N_1282,N_788,N_852);
xnor U1283 (N_1283,N_723,N_942);
nor U1284 (N_1284,N_536,N_646);
and U1285 (N_1285,N_704,N_701);
nor U1286 (N_1286,N_744,N_505);
and U1287 (N_1287,N_636,N_788);
nand U1288 (N_1288,N_757,N_944);
xor U1289 (N_1289,N_983,N_882);
or U1290 (N_1290,N_722,N_682);
xor U1291 (N_1291,N_849,N_771);
nor U1292 (N_1292,N_774,N_712);
nor U1293 (N_1293,N_882,N_938);
and U1294 (N_1294,N_714,N_731);
and U1295 (N_1295,N_690,N_824);
xor U1296 (N_1296,N_843,N_656);
xor U1297 (N_1297,N_910,N_709);
and U1298 (N_1298,N_517,N_657);
and U1299 (N_1299,N_961,N_670);
and U1300 (N_1300,N_791,N_636);
nand U1301 (N_1301,N_535,N_735);
nand U1302 (N_1302,N_839,N_668);
and U1303 (N_1303,N_615,N_675);
nor U1304 (N_1304,N_998,N_872);
nor U1305 (N_1305,N_715,N_740);
nand U1306 (N_1306,N_856,N_854);
nand U1307 (N_1307,N_741,N_672);
or U1308 (N_1308,N_751,N_948);
nor U1309 (N_1309,N_930,N_705);
or U1310 (N_1310,N_509,N_726);
and U1311 (N_1311,N_621,N_855);
and U1312 (N_1312,N_952,N_593);
or U1313 (N_1313,N_951,N_564);
nor U1314 (N_1314,N_574,N_644);
xor U1315 (N_1315,N_726,N_691);
nor U1316 (N_1316,N_756,N_791);
and U1317 (N_1317,N_661,N_976);
xnor U1318 (N_1318,N_629,N_956);
xnor U1319 (N_1319,N_620,N_750);
or U1320 (N_1320,N_784,N_728);
nor U1321 (N_1321,N_971,N_828);
xor U1322 (N_1322,N_842,N_964);
xor U1323 (N_1323,N_696,N_547);
nand U1324 (N_1324,N_553,N_906);
and U1325 (N_1325,N_885,N_916);
or U1326 (N_1326,N_947,N_711);
nand U1327 (N_1327,N_895,N_539);
or U1328 (N_1328,N_892,N_550);
or U1329 (N_1329,N_517,N_922);
xor U1330 (N_1330,N_583,N_942);
or U1331 (N_1331,N_857,N_961);
or U1332 (N_1332,N_874,N_546);
nor U1333 (N_1333,N_601,N_708);
xor U1334 (N_1334,N_968,N_527);
nand U1335 (N_1335,N_744,N_565);
nor U1336 (N_1336,N_762,N_894);
nand U1337 (N_1337,N_860,N_721);
or U1338 (N_1338,N_880,N_777);
or U1339 (N_1339,N_611,N_897);
or U1340 (N_1340,N_800,N_861);
nand U1341 (N_1341,N_950,N_765);
nor U1342 (N_1342,N_550,N_953);
or U1343 (N_1343,N_832,N_780);
nand U1344 (N_1344,N_778,N_583);
nor U1345 (N_1345,N_734,N_738);
or U1346 (N_1346,N_775,N_680);
and U1347 (N_1347,N_564,N_578);
and U1348 (N_1348,N_967,N_527);
nor U1349 (N_1349,N_835,N_500);
and U1350 (N_1350,N_570,N_987);
xor U1351 (N_1351,N_537,N_502);
nor U1352 (N_1352,N_800,N_602);
and U1353 (N_1353,N_704,N_733);
nor U1354 (N_1354,N_662,N_896);
and U1355 (N_1355,N_840,N_556);
xnor U1356 (N_1356,N_888,N_802);
nor U1357 (N_1357,N_769,N_890);
nand U1358 (N_1358,N_913,N_557);
and U1359 (N_1359,N_915,N_787);
xor U1360 (N_1360,N_716,N_622);
and U1361 (N_1361,N_522,N_514);
nand U1362 (N_1362,N_593,N_873);
and U1363 (N_1363,N_634,N_775);
nand U1364 (N_1364,N_779,N_866);
and U1365 (N_1365,N_701,N_799);
xnor U1366 (N_1366,N_501,N_946);
xor U1367 (N_1367,N_632,N_879);
and U1368 (N_1368,N_709,N_637);
and U1369 (N_1369,N_901,N_649);
nor U1370 (N_1370,N_801,N_776);
and U1371 (N_1371,N_521,N_784);
and U1372 (N_1372,N_895,N_657);
or U1373 (N_1373,N_612,N_714);
nand U1374 (N_1374,N_525,N_677);
and U1375 (N_1375,N_735,N_768);
xnor U1376 (N_1376,N_687,N_549);
or U1377 (N_1377,N_584,N_605);
and U1378 (N_1378,N_701,N_516);
nand U1379 (N_1379,N_699,N_621);
nor U1380 (N_1380,N_512,N_850);
nor U1381 (N_1381,N_701,N_868);
or U1382 (N_1382,N_555,N_719);
nor U1383 (N_1383,N_623,N_705);
nor U1384 (N_1384,N_623,N_833);
xor U1385 (N_1385,N_556,N_573);
xnor U1386 (N_1386,N_876,N_539);
nor U1387 (N_1387,N_874,N_731);
nand U1388 (N_1388,N_622,N_719);
and U1389 (N_1389,N_695,N_893);
nor U1390 (N_1390,N_659,N_708);
xnor U1391 (N_1391,N_519,N_820);
and U1392 (N_1392,N_632,N_584);
nor U1393 (N_1393,N_558,N_943);
nor U1394 (N_1394,N_527,N_617);
xnor U1395 (N_1395,N_503,N_856);
nor U1396 (N_1396,N_942,N_719);
nand U1397 (N_1397,N_507,N_797);
and U1398 (N_1398,N_907,N_873);
xor U1399 (N_1399,N_501,N_956);
nor U1400 (N_1400,N_730,N_980);
nand U1401 (N_1401,N_787,N_897);
or U1402 (N_1402,N_725,N_731);
nand U1403 (N_1403,N_908,N_562);
and U1404 (N_1404,N_873,N_816);
or U1405 (N_1405,N_810,N_561);
and U1406 (N_1406,N_950,N_851);
nand U1407 (N_1407,N_873,N_766);
and U1408 (N_1408,N_960,N_870);
nor U1409 (N_1409,N_945,N_942);
nand U1410 (N_1410,N_517,N_618);
or U1411 (N_1411,N_858,N_922);
nor U1412 (N_1412,N_665,N_794);
and U1413 (N_1413,N_781,N_519);
or U1414 (N_1414,N_581,N_592);
and U1415 (N_1415,N_849,N_826);
xnor U1416 (N_1416,N_802,N_615);
or U1417 (N_1417,N_941,N_915);
or U1418 (N_1418,N_640,N_770);
xnor U1419 (N_1419,N_516,N_583);
nor U1420 (N_1420,N_580,N_651);
xor U1421 (N_1421,N_656,N_879);
and U1422 (N_1422,N_630,N_524);
nor U1423 (N_1423,N_742,N_876);
nor U1424 (N_1424,N_513,N_716);
or U1425 (N_1425,N_780,N_819);
and U1426 (N_1426,N_653,N_732);
and U1427 (N_1427,N_585,N_684);
and U1428 (N_1428,N_936,N_650);
xor U1429 (N_1429,N_936,N_573);
nor U1430 (N_1430,N_920,N_604);
or U1431 (N_1431,N_582,N_895);
nand U1432 (N_1432,N_885,N_546);
nor U1433 (N_1433,N_908,N_513);
xor U1434 (N_1434,N_794,N_874);
xor U1435 (N_1435,N_767,N_761);
nand U1436 (N_1436,N_676,N_550);
nand U1437 (N_1437,N_648,N_620);
xnor U1438 (N_1438,N_530,N_902);
xnor U1439 (N_1439,N_724,N_799);
or U1440 (N_1440,N_551,N_940);
and U1441 (N_1441,N_526,N_682);
or U1442 (N_1442,N_961,N_810);
or U1443 (N_1443,N_571,N_728);
nand U1444 (N_1444,N_651,N_775);
nor U1445 (N_1445,N_582,N_825);
nand U1446 (N_1446,N_895,N_824);
nor U1447 (N_1447,N_745,N_535);
or U1448 (N_1448,N_542,N_805);
nor U1449 (N_1449,N_628,N_790);
and U1450 (N_1450,N_806,N_504);
or U1451 (N_1451,N_572,N_521);
or U1452 (N_1452,N_976,N_518);
xnor U1453 (N_1453,N_510,N_645);
xor U1454 (N_1454,N_910,N_722);
xnor U1455 (N_1455,N_845,N_501);
or U1456 (N_1456,N_823,N_921);
nand U1457 (N_1457,N_638,N_856);
nor U1458 (N_1458,N_657,N_723);
nand U1459 (N_1459,N_562,N_756);
and U1460 (N_1460,N_690,N_883);
nand U1461 (N_1461,N_871,N_832);
xnor U1462 (N_1462,N_777,N_871);
nand U1463 (N_1463,N_838,N_540);
nor U1464 (N_1464,N_909,N_986);
xor U1465 (N_1465,N_933,N_710);
nand U1466 (N_1466,N_714,N_800);
xnor U1467 (N_1467,N_861,N_883);
or U1468 (N_1468,N_651,N_820);
or U1469 (N_1469,N_579,N_810);
or U1470 (N_1470,N_986,N_972);
nand U1471 (N_1471,N_735,N_879);
xnor U1472 (N_1472,N_689,N_853);
or U1473 (N_1473,N_672,N_612);
xor U1474 (N_1474,N_829,N_899);
and U1475 (N_1475,N_622,N_527);
nand U1476 (N_1476,N_538,N_881);
xor U1477 (N_1477,N_617,N_929);
nand U1478 (N_1478,N_963,N_683);
or U1479 (N_1479,N_826,N_754);
xnor U1480 (N_1480,N_878,N_611);
nand U1481 (N_1481,N_936,N_974);
or U1482 (N_1482,N_657,N_636);
nand U1483 (N_1483,N_991,N_923);
and U1484 (N_1484,N_523,N_889);
nand U1485 (N_1485,N_868,N_501);
nor U1486 (N_1486,N_747,N_682);
or U1487 (N_1487,N_662,N_760);
nand U1488 (N_1488,N_747,N_942);
and U1489 (N_1489,N_701,N_691);
nor U1490 (N_1490,N_884,N_892);
xor U1491 (N_1491,N_866,N_758);
and U1492 (N_1492,N_670,N_889);
and U1493 (N_1493,N_774,N_657);
and U1494 (N_1494,N_887,N_540);
and U1495 (N_1495,N_720,N_861);
nand U1496 (N_1496,N_863,N_742);
xor U1497 (N_1497,N_943,N_517);
and U1498 (N_1498,N_975,N_819);
nand U1499 (N_1499,N_942,N_880);
or U1500 (N_1500,N_1458,N_1471);
nor U1501 (N_1501,N_1440,N_1166);
nand U1502 (N_1502,N_1211,N_1455);
or U1503 (N_1503,N_1046,N_1138);
xnor U1504 (N_1504,N_1269,N_1282);
nand U1505 (N_1505,N_1145,N_1228);
xnor U1506 (N_1506,N_1447,N_1162);
xor U1507 (N_1507,N_1451,N_1490);
xnor U1508 (N_1508,N_1175,N_1273);
nor U1509 (N_1509,N_1395,N_1460);
xnor U1510 (N_1510,N_1141,N_1288);
or U1511 (N_1511,N_1310,N_1109);
or U1512 (N_1512,N_1427,N_1432);
nand U1513 (N_1513,N_1015,N_1087);
and U1514 (N_1514,N_1268,N_1384);
nand U1515 (N_1515,N_1097,N_1445);
or U1516 (N_1516,N_1420,N_1317);
nand U1517 (N_1517,N_1121,N_1105);
and U1518 (N_1518,N_1462,N_1203);
nor U1519 (N_1519,N_1345,N_1017);
or U1520 (N_1520,N_1235,N_1479);
and U1521 (N_1521,N_1204,N_1403);
nand U1522 (N_1522,N_1278,N_1494);
or U1523 (N_1523,N_1313,N_1208);
xnor U1524 (N_1524,N_1114,N_1311);
nor U1525 (N_1525,N_1116,N_1159);
nand U1526 (N_1526,N_1354,N_1298);
nand U1527 (N_1527,N_1104,N_1302);
and U1528 (N_1528,N_1429,N_1459);
or U1529 (N_1529,N_1349,N_1179);
nand U1530 (N_1530,N_1001,N_1233);
or U1531 (N_1531,N_1346,N_1169);
xor U1532 (N_1532,N_1035,N_1468);
nor U1533 (N_1533,N_1144,N_1358);
and U1534 (N_1534,N_1243,N_1068);
nor U1535 (N_1535,N_1315,N_1366);
nand U1536 (N_1536,N_1394,N_1393);
xnor U1537 (N_1537,N_1078,N_1423);
and U1538 (N_1538,N_1409,N_1096);
xnor U1539 (N_1539,N_1437,N_1333);
xnor U1540 (N_1540,N_1245,N_1338);
or U1541 (N_1541,N_1020,N_1289);
nand U1542 (N_1542,N_1405,N_1417);
nand U1543 (N_1543,N_1402,N_1454);
and U1544 (N_1544,N_1182,N_1491);
and U1545 (N_1545,N_1307,N_1083);
xnor U1546 (N_1546,N_1343,N_1122);
or U1547 (N_1547,N_1254,N_1305);
xor U1548 (N_1548,N_1091,N_1192);
or U1549 (N_1549,N_1465,N_1359);
or U1550 (N_1550,N_1266,N_1406);
nand U1551 (N_1551,N_1255,N_1498);
nor U1552 (N_1552,N_1456,N_1484);
nor U1553 (N_1553,N_1201,N_1388);
nor U1554 (N_1554,N_1251,N_1106);
or U1555 (N_1555,N_1347,N_1133);
and U1556 (N_1556,N_1416,N_1308);
xnor U1557 (N_1557,N_1030,N_1271);
nor U1558 (N_1558,N_1339,N_1265);
nor U1559 (N_1559,N_1022,N_1280);
and U1560 (N_1560,N_1323,N_1057);
xor U1561 (N_1561,N_1332,N_1139);
or U1562 (N_1562,N_1019,N_1263);
nor U1563 (N_1563,N_1277,N_1143);
or U1564 (N_1564,N_1051,N_1329);
nand U1565 (N_1565,N_1441,N_1295);
or U1566 (N_1566,N_1399,N_1063);
xor U1567 (N_1567,N_1130,N_1286);
xnor U1568 (N_1568,N_1348,N_1352);
nor U1569 (N_1569,N_1005,N_1188);
nand U1570 (N_1570,N_1336,N_1476);
or U1571 (N_1571,N_1331,N_1256);
nor U1572 (N_1572,N_1361,N_1061);
and U1573 (N_1573,N_1378,N_1442);
nor U1574 (N_1574,N_1043,N_1385);
nor U1575 (N_1575,N_1197,N_1418);
or U1576 (N_1576,N_1064,N_1422);
xnor U1577 (N_1577,N_1190,N_1241);
nor U1578 (N_1578,N_1391,N_1168);
or U1579 (N_1579,N_1004,N_1234);
and U1580 (N_1580,N_1200,N_1248);
nand U1581 (N_1581,N_1027,N_1085);
or U1582 (N_1582,N_1340,N_1038);
xor U1583 (N_1583,N_1226,N_1267);
and U1584 (N_1584,N_1443,N_1438);
nand U1585 (N_1585,N_1009,N_1062);
or U1586 (N_1586,N_1368,N_1189);
xnor U1587 (N_1587,N_1342,N_1316);
xor U1588 (N_1588,N_1360,N_1483);
xnor U1589 (N_1589,N_1127,N_1379);
nand U1590 (N_1590,N_1374,N_1079);
nor U1591 (N_1591,N_1052,N_1067);
nor U1592 (N_1592,N_1164,N_1060);
and U1593 (N_1593,N_1047,N_1018);
xnor U1594 (N_1594,N_1088,N_1082);
nor U1595 (N_1595,N_1152,N_1229);
or U1596 (N_1596,N_1353,N_1369);
nand U1597 (N_1597,N_1187,N_1253);
and U1598 (N_1598,N_1172,N_1031);
nor U1599 (N_1599,N_1177,N_1351);
and U1600 (N_1600,N_1246,N_1225);
and U1601 (N_1601,N_1236,N_1397);
xor U1602 (N_1602,N_1135,N_1012);
nor U1603 (N_1603,N_1016,N_1222);
or U1604 (N_1604,N_1325,N_1185);
nor U1605 (N_1605,N_1238,N_1173);
nor U1606 (N_1606,N_1037,N_1006);
and U1607 (N_1607,N_1421,N_1493);
nor U1608 (N_1608,N_1381,N_1089);
xnor U1609 (N_1609,N_1231,N_1430);
and U1610 (N_1610,N_1446,N_1297);
and U1611 (N_1611,N_1364,N_1119);
nor U1612 (N_1612,N_1489,N_1382);
xnor U1613 (N_1613,N_1485,N_1053);
xnor U1614 (N_1614,N_1193,N_1362);
and U1615 (N_1615,N_1470,N_1327);
and U1616 (N_1616,N_1099,N_1032);
xnor U1617 (N_1617,N_1337,N_1070);
or U1618 (N_1618,N_1448,N_1077);
or U1619 (N_1619,N_1370,N_1206);
nor U1620 (N_1620,N_1186,N_1080);
nor U1621 (N_1621,N_1147,N_1158);
nand U1622 (N_1622,N_1334,N_1326);
nand U1623 (N_1623,N_1244,N_1216);
xnor U1624 (N_1624,N_1452,N_1086);
xnor U1625 (N_1625,N_1492,N_1002);
or U1626 (N_1626,N_1058,N_1355);
xor U1627 (N_1627,N_1090,N_1098);
and U1628 (N_1628,N_1372,N_1010);
nand U1629 (N_1629,N_1034,N_1249);
xnor U1630 (N_1630,N_1367,N_1467);
nand U1631 (N_1631,N_1318,N_1174);
xnor U1632 (N_1632,N_1457,N_1259);
and U1633 (N_1633,N_1050,N_1044);
or U1634 (N_1634,N_1434,N_1300);
and U1635 (N_1635,N_1041,N_1167);
or U1636 (N_1636,N_1274,N_1309);
nor U1637 (N_1637,N_1040,N_1103);
nand U1638 (N_1638,N_1408,N_1163);
xor U1639 (N_1639,N_1217,N_1198);
nand U1640 (N_1640,N_1102,N_1486);
and U1641 (N_1641,N_1142,N_1180);
xor U1642 (N_1642,N_1081,N_1008);
xnor U1643 (N_1643,N_1312,N_1093);
nor U1644 (N_1644,N_1392,N_1299);
xnor U1645 (N_1645,N_1487,N_1373);
or U1646 (N_1646,N_1341,N_1330);
xnor U1647 (N_1647,N_1021,N_1048);
or U1648 (N_1648,N_1232,N_1252);
xor U1649 (N_1649,N_1357,N_1202);
or U1650 (N_1650,N_1075,N_1140);
nor U1651 (N_1651,N_1469,N_1480);
xor U1652 (N_1652,N_1137,N_1319);
or U1653 (N_1653,N_1224,N_1112);
xor U1654 (N_1654,N_1146,N_1281);
xnor U1655 (N_1655,N_1150,N_1261);
nor U1656 (N_1656,N_1320,N_1377);
and U1657 (N_1657,N_1328,N_1110);
nor U1658 (N_1658,N_1153,N_1400);
nand U1659 (N_1659,N_1161,N_1219);
nor U1660 (N_1660,N_1247,N_1107);
nor U1661 (N_1661,N_1404,N_1292);
nor U1662 (N_1662,N_1453,N_1213);
and U1663 (N_1663,N_1165,N_1149);
nand U1664 (N_1664,N_1113,N_1013);
nor U1665 (N_1665,N_1356,N_1157);
or U1666 (N_1666,N_1195,N_1258);
or U1667 (N_1667,N_1294,N_1184);
nand U1668 (N_1668,N_1321,N_1171);
xnor U1669 (N_1669,N_1024,N_1304);
or U1670 (N_1670,N_1444,N_1055);
or U1671 (N_1671,N_1215,N_1371);
or U1672 (N_1672,N_1426,N_1056);
nand U1673 (N_1673,N_1084,N_1324);
nand U1674 (N_1674,N_1071,N_1136);
and U1675 (N_1675,N_1218,N_1101);
or U1676 (N_1676,N_1496,N_1413);
nand U1677 (N_1677,N_1191,N_1431);
nand U1678 (N_1678,N_1449,N_1499);
nand U1679 (N_1679,N_1039,N_1412);
nand U1680 (N_1680,N_1131,N_1223);
and U1681 (N_1681,N_1205,N_1303);
nor U1682 (N_1682,N_1207,N_1495);
nand U1683 (N_1683,N_1293,N_1115);
or U1684 (N_1684,N_1296,N_1072);
nor U1685 (N_1685,N_1124,N_1466);
nand U1686 (N_1686,N_1125,N_1128);
nor U1687 (N_1687,N_1387,N_1196);
nor U1688 (N_1688,N_1066,N_1003);
nor U1689 (N_1689,N_1477,N_1335);
and U1690 (N_1690,N_1276,N_1497);
or U1691 (N_1691,N_1380,N_1474);
nand U1692 (N_1692,N_1132,N_1290);
nand U1693 (N_1693,N_1069,N_1283);
xor U1694 (N_1694,N_1410,N_1212);
and U1695 (N_1695,N_1419,N_1428);
nor U1696 (N_1696,N_1092,N_1117);
xor U1697 (N_1697,N_1054,N_1156);
and U1698 (N_1698,N_1436,N_1076);
or U1699 (N_1699,N_1414,N_1396);
nand U1700 (N_1700,N_1264,N_1194);
and U1701 (N_1701,N_1045,N_1023);
nand U1702 (N_1702,N_1134,N_1240);
and U1703 (N_1703,N_1221,N_1170);
xnor U1704 (N_1704,N_1450,N_1007);
and U1705 (N_1705,N_1183,N_1178);
or U1706 (N_1706,N_1478,N_1095);
nor U1707 (N_1707,N_1036,N_1433);
nor U1708 (N_1708,N_1209,N_1059);
and U1709 (N_1709,N_1074,N_1472);
nand U1710 (N_1710,N_1424,N_1464);
or U1711 (N_1711,N_1463,N_1287);
and U1712 (N_1712,N_1151,N_1482);
or U1713 (N_1713,N_1250,N_1401);
or U1714 (N_1714,N_1025,N_1389);
xnor U1715 (N_1715,N_1314,N_1411);
nand U1716 (N_1716,N_1257,N_1129);
nand U1717 (N_1717,N_1042,N_1108);
xor U1718 (N_1718,N_1285,N_1461);
xor U1719 (N_1719,N_1435,N_1383);
nand U1720 (N_1720,N_1210,N_1473);
and U1721 (N_1721,N_1155,N_1033);
nor U1722 (N_1722,N_1011,N_1301);
nor U1723 (N_1723,N_1398,N_1481);
or U1724 (N_1724,N_1123,N_1239);
or U1725 (N_1725,N_1230,N_1322);
or U1726 (N_1726,N_1407,N_1363);
xnor U1727 (N_1727,N_1390,N_1475);
nor U1728 (N_1728,N_1120,N_1237);
xnor U1729 (N_1729,N_1439,N_1260);
or U1730 (N_1730,N_1272,N_1014);
nor U1731 (N_1731,N_1181,N_1242);
xnor U1732 (N_1732,N_1065,N_1275);
and U1733 (N_1733,N_1029,N_1344);
nor U1734 (N_1734,N_1415,N_1376);
and U1735 (N_1735,N_1199,N_1148);
xnor U1736 (N_1736,N_1375,N_1220);
and U1737 (N_1737,N_1425,N_1049);
or U1738 (N_1738,N_1111,N_1488);
and U1739 (N_1739,N_1100,N_1227);
xnor U1740 (N_1740,N_1118,N_1154);
nand U1741 (N_1741,N_1291,N_1306);
and U1742 (N_1742,N_1284,N_1073);
xnor U1743 (N_1743,N_1126,N_1386);
xnor U1744 (N_1744,N_1262,N_1026);
xnor U1745 (N_1745,N_1094,N_1000);
and U1746 (N_1746,N_1350,N_1214);
xor U1747 (N_1747,N_1279,N_1270);
nor U1748 (N_1748,N_1028,N_1160);
nand U1749 (N_1749,N_1365,N_1176);
or U1750 (N_1750,N_1178,N_1050);
and U1751 (N_1751,N_1146,N_1210);
xnor U1752 (N_1752,N_1046,N_1475);
nor U1753 (N_1753,N_1305,N_1021);
or U1754 (N_1754,N_1308,N_1236);
xnor U1755 (N_1755,N_1206,N_1237);
nor U1756 (N_1756,N_1118,N_1021);
xnor U1757 (N_1757,N_1269,N_1250);
nand U1758 (N_1758,N_1277,N_1000);
nand U1759 (N_1759,N_1464,N_1337);
nor U1760 (N_1760,N_1040,N_1151);
nand U1761 (N_1761,N_1142,N_1341);
nor U1762 (N_1762,N_1484,N_1014);
xnor U1763 (N_1763,N_1117,N_1435);
xnor U1764 (N_1764,N_1036,N_1055);
nor U1765 (N_1765,N_1284,N_1198);
and U1766 (N_1766,N_1458,N_1281);
nand U1767 (N_1767,N_1030,N_1383);
or U1768 (N_1768,N_1344,N_1031);
nand U1769 (N_1769,N_1056,N_1212);
xnor U1770 (N_1770,N_1215,N_1128);
or U1771 (N_1771,N_1313,N_1202);
xnor U1772 (N_1772,N_1242,N_1021);
nand U1773 (N_1773,N_1175,N_1482);
nand U1774 (N_1774,N_1497,N_1082);
xor U1775 (N_1775,N_1005,N_1294);
nor U1776 (N_1776,N_1163,N_1319);
nand U1777 (N_1777,N_1131,N_1186);
or U1778 (N_1778,N_1204,N_1169);
nand U1779 (N_1779,N_1128,N_1296);
or U1780 (N_1780,N_1022,N_1094);
or U1781 (N_1781,N_1121,N_1196);
xor U1782 (N_1782,N_1113,N_1490);
and U1783 (N_1783,N_1251,N_1207);
or U1784 (N_1784,N_1402,N_1122);
nand U1785 (N_1785,N_1083,N_1141);
nor U1786 (N_1786,N_1005,N_1140);
and U1787 (N_1787,N_1217,N_1175);
or U1788 (N_1788,N_1241,N_1452);
and U1789 (N_1789,N_1495,N_1442);
nand U1790 (N_1790,N_1205,N_1085);
nor U1791 (N_1791,N_1287,N_1032);
nand U1792 (N_1792,N_1324,N_1411);
xnor U1793 (N_1793,N_1060,N_1481);
xor U1794 (N_1794,N_1364,N_1051);
nand U1795 (N_1795,N_1000,N_1212);
or U1796 (N_1796,N_1259,N_1347);
and U1797 (N_1797,N_1223,N_1197);
or U1798 (N_1798,N_1068,N_1408);
and U1799 (N_1799,N_1477,N_1210);
and U1800 (N_1800,N_1092,N_1047);
nand U1801 (N_1801,N_1030,N_1065);
xnor U1802 (N_1802,N_1140,N_1268);
or U1803 (N_1803,N_1300,N_1188);
and U1804 (N_1804,N_1061,N_1273);
or U1805 (N_1805,N_1180,N_1000);
xor U1806 (N_1806,N_1428,N_1306);
xnor U1807 (N_1807,N_1378,N_1069);
nor U1808 (N_1808,N_1152,N_1286);
nor U1809 (N_1809,N_1498,N_1197);
nand U1810 (N_1810,N_1284,N_1351);
nand U1811 (N_1811,N_1245,N_1472);
nand U1812 (N_1812,N_1177,N_1193);
and U1813 (N_1813,N_1032,N_1447);
and U1814 (N_1814,N_1336,N_1380);
and U1815 (N_1815,N_1275,N_1320);
and U1816 (N_1816,N_1223,N_1120);
or U1817 (N_1817,N_1167,N_1168);
nor U1818 (N_1818,N_1420,N_1132);
xnor U1819 (N_1819,N_1046,N_1274);
xnor U1820 (N_1820,N_1094,N_1220);
or U1821 (N_1821,N_1326,N_1033);
or U1822 (N_1822,N_1375,N_1183);
and U1823 (N_1823,N_1307,N_1106);
or U1824 (N_1824,N_1137,N_1353);
xor U1825 (N_1825,N_1457,N_1453);
or U1826 (N_1826,N_1085,N_1234);
nor U1827 (N_1827,N_1165,N_1492);
nor U1828 (N_1828,N_1095,N_1234);
or U1829 (N_1829,N_1215,N_1121);
nor U1830 (N_1830,N_1320,N_1302);
nor U1831 (N_1831,N_1399,N_1262);
xnor U1832 (N_1832,N_1415,N_1321);
nor U1833 (N_1833,N_1178,N_1340);
or U1834 (N_1834,N_1462,N_1286);
or U1835 (N_1835,N_1253,N_1256);
nand U1836 (N_1836,N_1246,N_1320);
nand U1837 (N_1837,N_1390,N_1426);
and U1838 (N_1838,N_1423,N_1451);
and U1839 (N_1839,N_1281,N_1282);
nand U1840 (N_1840,N_1051,N_1480);
nand U1841 (N_1841,N_1288,N_1226);
and U1842 (N_1842,N_1275,N_1395);
and U1843 (N_1843,N_1271,N_1092);
or U1844 (N_1844,N_1137,N_1415);
xor U1845 (N_1845,N_1372,N_1378);
nand U1846 (N_1846,N_1315,N_1115);
xnor U1847 (N_1847,N_1485,N_1341);
or U1848 (N_1848,N_1309,N_1460);
and U1849 (N_1849,N_1316,N_1042);
nor U1850 (N_1850,N_1310,N_1352);
nor U1851 (N_1851,N_1479,N_1376);
nor U1852 (N_1852,N_1237,N_1037);
nand U1853 (N_1853,N_1048,N_1175);
or U1854 (N_1854,N_1491,N_1405);
nor U1855 (N_1855,N_1170,N_1154);
nand U1856 (N_1856,N_1458,N_1236);
and U1857 (N_1857,N_1477,N_1013);
nand U1858 (N_1858,N_1288,N_1079);
and U1859 (N_1859,N_1384,N_1496);
and U1860 (N_1860,N_1475,N_1440);
and U1861 (N_1861,N_1361,N_1208);
and U1862 (N_1862,N_1081,N_1472);
and U1863 (N_1863,N_1286,N_1334);
or U1864 (N_1864,N_1473,N_1379);
xnor U1865 (N_1865,N_1234,N_1253);
and U1866 (N_1866,N_1305,N_1388);
xnor U1867 (N_1867,N_1222,N_1046);
or U1868 (N_1868,N_1454,N_1258);
or U1869 (N_1869,N_1238,N_1165);
or U1870 (N_1870,N_1311,N_1426);
nor U1871 (N_1871,N_1259,N_1218);
nand U1872 (N_1872,N_1447,N_1226);
xor U1873 (N_1873,N_1105,N_1039);
xor U1874 (N_1874,N_1334,N_1353);
xnor U1875 (N_1875,N_1003,N_1277);
or U1876 (N_1876,N_1092,N_1496);
and U1877 (N_1877,N_1207,N_1057);
xor U1878 (N_1878,N_1411,N_1091);
or U1879 (N_1879,N_1129,N_1392);
nand U1880 (N_1880,N_1354,N_1357);
nand U1881 (N_1881,N_1225,N_1266);
xnor U1882 (N_1882,N_1253,N_1293);
nand U1883 (N_1883,N_1115,N_1139);
nand U1884 (N_1884,N_1218,N_1366);
nand U1885 (N_1885,N_1282,N_1334);
and U1886 (N_1886,N_1409,N_1181);
nand U1887 (N_1887,N_1327,N_1352);
nor U1888 (N_1888,N_1031,N_1183);
nand U1889 (N_1889,N_1493,N_1382);
or U1890 (N_1890,N_1424,N_1317);
and U1891 (N_1891,N_1080,N_1159);
or U1892 (N_1892,N_1283,N_1334);
or U1893 (N_1893,N_1124,N_1345);
nor U1894 (N_1894,N_1243,N_1016);
and U1895 (N_1895,N_1435,N_1249);
or U1896 (N_1896,N_1342,N_1000);
nor U1897 (N_1897,N_1315,N_1111);
nor U1898 (N_1898,N_1291,N_1015);
xor U1899 (N_1899,N_1169,N_1483);
or U1900 (N_1900,N_1414,N_1340);
xor U1901 (N_1901,N_1262,N_1032);
nor U1902 (N_1902,N_1090,N_1144);
nand U1903 (N_1903,N_1421,N_1043);
or U1904 (N_1904,N_1008,N_1267);
and U1905 (N_1905,N_1452,N_1369);
nor U1906 (N_1906,N_1184,N_1322);
or U1907 (N_1907,N_1283,N_1029);
xnor U1908 (N_1908,N_1168,N_1261);
nand U1909 (N_1909,N_1171,N_1415);
nand U1910 (N_1910,N_1368,N_1355);
and U1911 (N_1911,N_1322,N_1052);
nand U1912 (N_1912,N_1078,N_1092);
or U1913 (N_1913,N_1003,N_1359);
or U1914 (N_1914,N_1436,N_1258);
xnor U1915 (N_1915,N_1465,N_1493);
nor U1916 (N_1916,N_1001,N_1015);
nand U1917 (N_1917,N_1214,N_1026);
and U1918 (N_1918,N_1290,N_1324);
xnor U1919 (N_1919,N_1471,N_1028);
and U1920 (N_1920,N_1320,N_1009);
nand U1921 (N_1921,N_1448,N_1401);
nor U1922 (N_1922,N_1432,N_1448);
and U1923 (N_1923,N_1272,N_1116);
nand U1924 (N_1924,N_1434,N_1313);
nor U1925 (N_1925,N_1378,N_1299);
xor U1926 (N_1926,N_1123,N_1189);
nor U1927 (N_1927,N_1061,N_1314);
or U1928 (N_1928,N_1316,N_1186);
xor U1929 (N_1929,N_1113,N_1284);
xor U1930 (N_1930,N_1133,N_1489);
nor U1931 (N_1931,N_1303,N_1445);
or U1932 (N_1932,N_1156,N_1197);
nor U1933 (N_1933,N_1207,N_1296);
and U1934 (N_1934,N_1206,N_1300);
nand U1935 (N_1935,N_1045,N_1394);
xor U1936 (N_1936,N_1418,N_1104);
and U1937 (N_1937,N_1000,N_1352);
nand U1938 (N_1938,N_1388,N_1351);
or U1939 (N_1939,N_1080,N_1116);
nand U1940 (N_1940,N_1250,N_1214);
xor U1941 (N_1941,N_1370,N_1235);
or U1942 (N_1942,N_1112,N_1482);
and U1943 (N_1943,N_1423,N_1260);
xor U1944 (N_1944,N_1017,N_1075);
xor U1945 (N_1945,N_1356,N_1360);
xnor U1946 (N_1946,N_1451,N_1186);
and U1947 (N_1947,N_1311,N_1450);
and U1948 (N_1948,N_1054,N_1037);
nor U1949 (N_1949,N_1439,N_1449);
or U1950 (N_1950,N_1207,N_1211);
nor U1951 (N_1951,N_1266,N_1125);
xnor U1952 (N_1952,N_1111,N_1229);
nand U1953 (N_1953,N_1259,N_1254);
and U1954 (N_1954,N_1103,N_1277);
nand U1955 (N_1955,N_1106,N_1354);
xor U1956 (N_1956,N_1132,N_1263);
and U1957 (N_1957,N_1169,N_1105);
or U1958 (N_1958,N_1177,N_1243);
xnor U1959 (N_1959,N_1386,N_1208);
nand U1960 (N_1960,N_1404,N_1060);
nor U1961 (N_1961,N_1338,N_1118);
xnor U1962 (N_1962,N_1031,N_1499);
nand U1963 (N_1963,N_1157,N_1053);
nor U1964 (N_1964,N_1440,N_1072);
nand U1965 (N_1965,N_1194,N_1394);
and U1966 (N_1966,N_1290,N_1323);
xor U1967 (N_1967,N_1278,N_1410);
or U1968 (N_1968,N_1097,N_1176);
nand U1969 (N_1969,N_1143,N_1159);
nand U1970 (N_1970,N_1400,N_1355);
or U1971 (N_1971,N_1415,N_1429);
or U1972 (N_1972,N_1178,N_1169);
and U1973 (N_1973,N_1392,N_1333);
nand U1974 (N_1974,N_1422,N_1238);
xor U1975 (N_1975,N_1135,N_1463);
or U1976 (N_1976,N_1082,N_1253);
xnor U1977 (N_1977,N_1421,N_1057);
xor U1978 (N_1978,N_1415,N_1244);
xor U1979 (N_1979,N_1284,N_1005);
or U1980 (N_1980,N_1027,N_1432);
or U1981 (N_1981,N_1461,N_1029);
or U1982 (N_1982,N_1474,N_1360);
xnor U1983 (N_1983,N_1296,N_1223);
xnor U1984 (N_1984,N_1226,N_1127);
or U1985 (N_1985,N_1446,N_1452);
and U1986 (N_1986,N_1472,N_1008);
nand U1987 (N_1987,N_1323,N_1340);
xnor U1988 (N_1988,N_1362,N_1259);
nand U1989 (N_1989,N_1074,N_1143);
xnor U1990 (N_1990,N_1449,N_1389);
nor U1991 (N_1991,N_1313,N_1308);
nor U1992 (N_1992,N_1200,N_1327);
and U1993 (N_1993,N_1489,N_1010);
nand U1994 (N_1994,N_1390,N_1379);
nor U1995 (N_1995,N_1197,N_1206);
and U1996 (N_1996,N_1021,N_1033);
nor U1997 (N_1997,N_1479,N_1062);
xor U1998 (N_1998,N_1455,N_1499);
or U1999 (N_1999,N_1301,N_1067);
or U2000 (N_2000,N_1579,N_1787);
nand U2001 (N_2001,N_1925,N_1941);
or U2002 (N_2002,N_1529,N_1693);
or U2003 (N_2003,N_1692,N_1739);
and U2004 (N_2004,N_1583,N_1895);
nor U2005 (N_2005,N_1537,N_1590);
nor U2006 (N_2006,N_1545,N_1868);
nor U2007 (N_2007,N_1942,N_1791);
nand U2008 (N_2008,N_1515,N_1632);
or U2009 (N_2009,N_1957,N_1792);
xnor U2010 (N_2010,N_1685,N_1520);
nand U2011 (N_2011,N_1843,N_1587);
or U2012 (N_2012,N_1778,N_1907);
or U2013 (N_2013,N_1997,N_1544);
xnor U2014 (N_2014,N_1728,N_1858);
xnor U2015 (N_2015,N_1839,N_1972);
or U2016 (N_2016,N_1795,N_1603);
xnor U2017 (N_2017,N_1646,N_1859);
and U2018 (N_2018,N_1666,N_1638);
and U2019 (N_2019,N_1541,N_1744);
and U2020 (N_2020,N_1500,N_1619);
xnor U2021 (N_2021,N_1917,N_1518);
and U2022 (N_2022,N_1840,N_1662);
nand U2023 (N_2023,N_1849,N_1650);
nor U2024 (N_2024,N_1533,N_1585);
xor U2025 (N_2025,N_1622,N_1887);
nor U2026 (N_2026,N_1749,N_1821);
or U2027 (N_2027,N_1834,N_1673);
or U2028 (N_2028,N_1540,N_1893);
xor U2029 (N_2029,N_1714,N_1885);
nor U2030 (N_2030,N_1629,N_1823);
nor U2031 (N_2031,N_1595,N_1551);
xnor U2032 (N_2032,N_1888,N_1920);
nand U2033 (N_2033,N_1855,N_1543);
or U2034 (N_2034,N_1562,N_1709);
xor U2035 (N_2035,N_1530,N_1674);
nor U2036 (N_2036,N_1794,N_1656);
nand U2037 (N_2037,N_1926,N_1737);
and U2038 (N_2038,N_1560,N_1642);
nor U2039 (N_2039,N_1940,N_1669);
and U2040 (N_2040,N_1526,N_1929);
nor U2041 (N_2041,N_1523,N_1575);
nand U2042 (N_2042,N_1862,N_1820);
or U2043 (N_2043,N_1557,N_1976);
nand U2044 (N_2044,N_1912,N_1829);
xnor U2045 (N_2045,N_1733,N_1747);
and U2046 (N_2046,N_1513,N_1886);
and U2047 (N_2047,N_1683,N_1775);
xor U2048 (N_2048,N_1731,N_1758);
xor U2049 (N_2049,N_1876,N_1814);
nand U2050 (N_2050,N_1591,N_1600);
and U2051 (N_2051,N_1548,N_1715);
nor U2052 (N_2052,N_1741,N_1952);
nand U2053 (N_2053,N_1784,N_1748);
nor U2054 (N_2054,N_1732,N_1863);
nand U2055 (N_2055,N_1798,N_1802);
or U2056 (N_2056,N_1527,N_1865);
nor U2057 (N_2057,N_1664,N_1634);
or U2058 (N_2058,N_1934,N_1670);
nand U2059 (N_2059,N_1780,N_1576);
nor U2060 (N_2060,N_1854,N_1652);
xor U2061 (N_2061,N_1531,N_1711);
xor U2062 (N_2062,N_1860,N_1809);
or U2063 (N_2063,N_1759,N_1723);
nand U2064 (N_2064,N_1751,N_1909);
or U2065 (N_2065,N_1774,N_1663);
or U2066 (N_2066,N_1640,N_1648);
or U2067 (N_2067,N_1736,N_1776);
and U2068 (N_2068,N_1954,N_1625);
xor U2069 (N_2069,N_1597,N_1695);
or U2070 (N_2070,N_1818,N_1610);
or U2071 (N_2071,N_1989,N_1686);
nor U2072 (N_2072,N_1841,N_1569);
or U2073 (N_2073,N_1913,N_1967);
or U2074 (N_2074,N_1788,N_1617);
nand U2075 (N_2075,N_1931,N_1914);
nor U2076 (N_2076,N_1897,N_1971);
xor U2077 (N_2077,N_1963,N_1742);
xor U2078 (N_2078,N_1980,N_1810);
nand U2079 (N_2079,N_1556,N_1719);
and U2080 (N_2080,N_1892,N_1826);
or U2081 (N_2081,N_1990,N_1985);
nor U2082 (N_2082,N_1573,N_1875);
xnor U2083 (N_2083,N_1512,N_1701);
or U2084 (N_2084,N_1800,N_1815);
nand U2085 (N_2085,N_1630,N_1570);
or U2086 (N_2086,N_1890,N_1994);
nand U2087 (N_2087,N_1961,N_1824);
xor U2088 (N_2088,N_1756,N_1785);
and U2089 (N_2089,N_1953,N_1986);
xor U2090 (N_2090,N_1832,N_1828);
or U2091 (N_2091,N_1665,N_1707);
nand U2092 (N_2092,N_1684,N_1535);
nor U2093 (N_2093,N_1555,N_1704);
nor U2094 (N_2094,N_1768,N_1996);
or U2095 (N_2095,N_1835,N_1697);
xor U2096 (N_2096,N_1633,N_1998);
nand U2097 (N_2097,N_1528,N_1611);
nor U2098 (N_2098,N_1702,N_1898);
nor U2099 (N_2099,N_1962,N_1613);
or U2100 (N_2100,N_1883,N_1869);
xor U2101 (N_2101,N_1593,N_1675);
or U2102 (N_2102,N_1988,N_1959);
and U2103 (N_2103,N_1750,N_1889);
xor U2104 (N_2104,N_1882,N_1866);
nor U2105 (N_2105,N_1752,N_1606);
nand U2106 (N_2106,N_1908,N_1844);
xor U2107 (N_2107,N_1667,N_1906);
xor U2108 (N_2108,N_1981,N_1838);
nor U2109 (N_2109,N_1745,N_1921);
and U2110 (N_2110,N_1760,N_1974);
nor U2111 (N_2111,N_1764,N_1729);
nor U2112 (N_2112,N_1822,N_1896);
xnor U2113 (N_2113,N_1509,N_1905);
xnor U2114 (N_2114,N_1574,N_1812);
xor U2115 (N_2115,N_1904,N_1726);
nand U2116 (N_2116,N_1973,N_1793);
and U2117 (N_2117,N_1644,N_1825);
and U2118 (N_2118,N_1521,N_1580);
nor U2119 (N_2119,N_1945,N_1502);
and U2120 (N_2120,N_1947,N_1511);
and U2121 (N_2121,N_1568,N_1903);
nand U2122 (N_2122,N_1561,N_1628);
or U2123 (N_2123,N_1660,N_1690);
nand U2124 (N_2124,N_1982,N_1682);
or U2125 (N_2125,N_1867,N_1979);
or U2126 (N_2126,N_1679,N_1517);
nor U2127 (N_2127,N_1939,N_1582);
xnor U2128 (N_2128,N_1938,N_1539);
or U2129 (N_2129,N_1577,N_1910);
nor U2130 (N_2130,N_1532,N_1836);
xnor U2131 (N_2131,N_1522,N_1703);
or U2132 (N_2132,N_1955,N_1857);
xor U2133 (N_2133,N_1618,N_1678);
xnor U2134 (N_2134,N_1668,N_1789);
nand U2135 (N_2135,N_1902,N_1722);
and U2136 (N_2136,N_1525,N_1738);
or U2137 (N_2137,N_1927,N_1688);
xor U2138 (N_2138,N_1861,N_1734);
and U2139 (N_2139,N_1599,N_1878);
nand U2140 (N_2140,N_1804,N_1969);
and U2141 (N_2141,N_1779,N_1873);
nor U2142 (N_2142,N_1833,N_1699);
nor U2143 (N_2143,N_1501,N_1853);
nand U2144 (N_2144,N_1566,N_1717);
or U2145 (N_2145,N_1647,N_1949);
nand U2146 (N_2146,N_1589,N_1880);
nor U2147 (N_2147,N_1546,N_1965);
or U2148 (N_2148,N_1598,N_1547);
nand U2149 (N_2149,N_1700,N_1643);
or U2150 (N_2150,N_1746,N_1870);
or U2151 (N_2151,N_1505,N_1725);
nor U2152 (N_2152,N_1637,N_1596);
nand U2153 (N_2153,N_1773,N_1559);
nor U2154 (N_2154,N_1842,N_1915);
xor U2155 (N_2155,N_1708,N_1616);
nand U2156 (N_2156,N_1783,N_1874);
or U2157 (N_2157,N_1992,N_1924);
or U2158 (N_2158,N_1901,N_1932);
nand U2159 (N_2159,N_1602,N_1594);
xnor U2160 (N_2160,N_1631,N_1916);
nor U2161 (N_2161,N_1645,N_1626);
nand U2162 (N_2162,N_1592,N_1805);
xnor U2163 (N_2163,N_1970,N_1718);
or U2164 (N_2164,N_1884,N_1609);
nand U2165 (N_2165,N_1837,N_1951);
or U2166 (N_2166,N_1654,N_1894);
nor U2167 (N_2167,N_1687,N_1659);
or U2168 (N_2168,N_1950,N_1935);
or U2169 (N_2169,N_1771,N_1510);
nor U2170 (N_2170,N_1677,N_1991);
xnor U2171 (N_2171,N_1584,N_1581);
nand U2172 (N_2172,N_1790,N_1724);
xor U2173 (N_2173,N_1588,N_1767);
nand U2174 (N_2174,N_1919,N_1524);
xnor U2175 (N_2175,N_1694,N_1765);
nor U2176 (N_2176,N_1864,N_1676);
and U2177 (N_2177,N_1655,N_1571);
xnor U2178 (N_2178,N_1946,N_1564);
xnor U2179 (N_2179,N_1827,N_1706);
nand U2180 (N_2180,N_1621,N_1984);
or U2181 (N_2181,N_1636,N_1830);
or U2182 (N_2182,N_1743,N_1993);
nor U2183 (N_2183,N_1504,N_1937);
xnor U2184 (N_2184,N_1769,N_1608);
or U2185 (N_2185,N_1691,N_1796);
and U2186 (N_2186,N_1657,N_1720);
xnor U2187 (N_2187,N_1772,N_1604);
xnor U2188 (N_2188,N_1508,N_1538);
and U2189 (N_2189,N_1923,N_1536);
and U2190 (N_2190,N_1730,N_1808);
xnor U2191 (N_2191,N_1936,N_1503);
and U2192 (N_2192,N_1554,N_1757);
or U2193 (N_2193,N_1671,N_1943);
and U2194 (N_2194,N_1506,N_1816);
or U2195 (N_2195,N_1968,N_1698);
nor U2196 (N_2196,N_1987,N_1807);
nor U2197 (N_2197,N_1845,N_1542);
xnor U2198 (N_2198,N_1507,N_1797);
nand U2199 (N_2199,N_1911,N_1766);
or U2200 (N_2200,N_1817,N_1627);
xor U2201 (N_2201,N_1620,N_1964);
nor U2202 (N_2202,N_1851,N_1977);
nand U2203 (N_2203,N_1705,N_1813);
nor U2204 (N_2204,N_1735,N_1777);
or U2205 (N_2205,N_1881,N_1534);
and U2206 (N_2206,N_1565,N_1516);
nand U2207 (N_2207,N_1801,N_1624);
and U2208 (N_2208,N_1721,N_1930);
nor U2209 (N_2209,N_1680,N_1614);
and U2210 (N_2210,N_1653,N_1761);
nand U2211 (N_2211,N_1672,N_1960);
nand U2212 (N_2212,N_1850,N_1763);
nor U2213 (N_2213,N_1607,N_1782);
nand U2214 (N_2214,N_1770,N_1786);
xnor U2215 (N_2215,N_1995,N_1944);
or U2216 (N_2216,N_1553,N_1716);
nand U2217 (N_2217,N_1948,N_1681);
nor U2218 (N_2218,N_1586,N_1856);
and U2219 (N_2219,N_1514,N_1572);
nor U2220 (N_2220,N_1848,N_1819);
or U2221 (N_2221,N_1891,N_1799);
xor U2222 (N_2222,N_1710,N_1900);
and U2223 (N_2223,N_1519,N_1605);
nor U2224 (N_2224,N_1740,N_1696);
xor U2225 (N_2225,N_1811,N_1754);
xor U2226 (N_2226,N_1975,N_1549);
and U2227 (N_2227,N_1831,N_1978);
and U2228 (N_2228,N_1933,N_1552);
xor U2229 (N_2229,N_1871,N_1899);
and U2230 (N_2230,N_1649,N_1966);
xnor U2231 (N_2231,N_1550,N_1658);
or U2232 (N_2232,N_1612,N_1641);
nor U2233 (N_2233,N_1872,N_1578);
xnor U2234 (N_2234,N_1601,N_1661);
nand U2235 (N_2235,N_1928,N_1803);
xor U2236 (N_2236,N_1918,N_1806);
nand U2237 (N_2237,N_1958,N_1689);
or U2238 (N_2238,N_1846,N_1639);
xnor U2239 (N_2239,N_1999,N_1852);
and U2240 (N_2240,N_1563,N_1558);
nand U2241 (N_2241,N_1879,N_1877);
nor U2242 (N_2242,N_1713,N_1755);
or U2243 (N_2243,N_1781,N_1615);
xor U2244 (N_2244,N_1983,N_1956);
or U2245 (N_2245,N_1623,N_1712);
and U2246 (N_2246,N_1922,N_1567);
nand U2247 (N_2247,N_1727,N_1847);
and U2248 (N_2248,N_1635,N_1651);
or U2249 (N_2249,N_1753,N_1762);
xnor U2250 (N_2250,N_1708,N_1649);
and U2251 (N_2251,N_1550,N_1597);
nor U2252 (N_2252,N_1821,N_1844);
or U2253 (N_2253,N_1819,N_1960);
or U2254 (N_2254,N_1529,N_1816);
xor U2255 (N_2255,N_1564,N_1574);
or U2256 (N_2256,N_1736,N_1728);
nor U2257 (N_2257,N_1736,N_1504);
nor U2258 (N_2258,N_1908,N_1879);
xnor U2259 (N_2259,N_1868,N_1840);
nand U2260 (N_2260,N_1817,N_1866);
or U2261 (N_2261,N_1601,N_1633);
or U2262 (N_2262,N_1590,N_1943);
or U2263 (N_2263,N_1989,N_1979);
nor U2264 (N_2264,N_1531,N_1710);
nand U2265 (N_2265,N_1533,N_1964);
nand U2266 (N_2266,N_1628,N_1995);
or U2267 (N_2267,N_1615,N_1859);
or U2268 (N_2268,N_1613,N_1593);
xor U2269 (N_2269,N_1996,N_1872);
nand U2270 (N_2270,N_1874,N_1748);
nor U2271 (N_2271,N_1546,N_1696);
and U2272 (N_2272,N_1888,N_1666);
nand U2273 (N_2273,N_1759,N_1584);
or U2274 (N_2274,N_1682,N_1811);
xor U2275 (N_2275,N_1657,N_1779);
xor U2276 (N_2276,N_1622,N_1505);
or U2277 (N_2277,N_1973,N_1775);
or U2278 (N_2278,N_1708,N_1998);
nand U2279 (N_2279,N_1538,N_1764);
and U2280 (N_2280,N_1622,N_1625);
nor U2281 (N_2281,N_1788,N_1710);
nor U2282 (N_2282,N_1960,N_1916);
and U2283 (N_2283,N_1689,N_1789);
nand U2284 (N_2284,N_1595,N_1591);
nand U2285 (N_2285,N_1783,N_1697);
and U2286 (N_2286,N_1971,N_1801);
nor U2287 (N_2287,N_1542,N_1884);
and U2288 (N_2288,N_1776,N_1534);
nand U2289 (N_2289,N_1506,N_1629);
nand U2290 (N_2290,N_1529,N_1704);
nor U2291 (N_2291,N_1608,N_1768);
nand U2292 (N_2292,N_1521,N_1789);
nand U2293 (N_2293,N_1724,N_1846);
nand U2294 (N_2294,N_1551,N_1665);
nand U2295 (N_2295,N_1698,N_1576);
nor U2296 (N_2296,N_1759,N_1951);
nor U2297 (N_2297,N_1850,N_1581);
and U2298 (N_2298,N_1643,N_1592);
nand U2299 (N_2299,N_1975,N_1719);
nor U2300 (N_2300,N_1724,N_1999);
xnor U2301 (N_2301,N_1536,N_1697);
xnor U2302 (N_2302,N_1605,N_1851);
nand U2303 (N_2303,N_1752,N_1647);
nand U2304 (N_2304,N_1757,N_1599);
or U2305 (N_2305,N_1690,N_1586);
nor U2306 (N_2306,N_1892,N_1992);
and U2307 (N_2307,N_1841,N_1675);
xor U2308 (N_2308,N_1539,N_1545);
nor U2309 (N_2309,N_1783,N_1939);
and U2310 (N_2310,N_1602,N_1567);
nand U2311 (N_2311,N_1610,N_1718);
and U2312 (N_2312,N_1817,N_1907);
or U2313 (N_2313,N_1709,N_1592);
xor U2314 (N_2314,N_1894,N_1534);
and U2315 (N_2315,N_1768,N_1616);
xor U2316 (N_2316,N_1819,N_1727);
or U2317 (N_2317,N_1822,N_1977);
or U2318 (N_2318,N_1598,N_1694);
nand U2319 (N_2319,N_1813,N_1682);
nor U2320 (N_2320,N_1840,N_1668);
xor U2321 (N_2321,N_1785,N_1924);
and U2322 (N_2322,N_1544,N_1564);
nor U2323 (N_2323,N_1841,N_1747);
or U2324 (N_2324,N_1699,N_1963);
and U2325 (N_2325,N_1578,N_1631);
nor U2326 (N_2326,N_1871,N_1867);
and U2327 (N_2327,N_1687,N_1749);
nand U2328 (N_2328,N_1941,N_1754);
nand U2329 (N_2329,N_1890,N_1760);
xor U2330 (N_2330,N_1610,N_1681);
xnor U2331 (N_2331,N_1809,N_1659);
xnor U2332 (N_2332,N_1868,N_1659);
or U2333 (N_2333,N_1727,N_1985);
nor U2334 (N_2334,N_1603,N_1686);
nor U2335 (N_2335,N_1685,N_1738);
nor U2336 (N_2336,N_1648,N_1858);
and U2337 (N_2337,N_1878,N_1877);
nand U2338 (N_2338,N_1931,N_1998);
and U2339 (N_2339,N_1879,N_1510);
xnor U2340 (N_2340,N_1745,N_1684);
nor U2341 (N_2341,N_1757,N_1935);
or U2342 (N_2342,N_1683,N_1928);
nand U2343 (N_2343,N_1505,N_1710);
and U2344 (N_2344,N_1561,N_1855);
nand U2345 (N_2345,N_1907,N_1770);
or U2346 (N_2346,N_1878,N_1672);
and U2347 (N_2347,N_1557,N_1885);
or U2348 (N_2348,N_1536,N_1552);
and U2349 (N_2349,N_1982,N_1791);
and U2350 (N_2350,N_1618,N_1946);
nor U2351 (N_2351,N_1936,N_1511);
nand U2352 (N_2352,N_1912,N_1629);
nor U2353 (N_2353,N_1881,N_1578);
nand U2354 (N_2354,N_1767,N_1676);
or U2355 (N_2355,N_1507,N_1834);
nand U2356 (N_2356,N_1523,N_1938);
nand U2357 (N_2357,N_1911,N_1560);
xnor U2358 (N_2358,N_1581,N_1823);
or U2359 (N_2359,N_1910,N_1558);
xor U2360 (N_2360,N_1647,N_1867);
or U2361 (N_2361,N_1500,N_1982);
and U2362 (N_2362,N_1585,N_1794);
nor U2363 (N_2363,N_1656,N_1904);
or U2364 (N_2364,N_1528,N_1842);
nor U2365 (N_2365,N_1805,N_1910);
or U2366 (N_2366,N_1628,N_1509);
nand U2367 (N_2367,N_1687,N_1955);
nor U2368 (N_2368,N_1585,N_1830);
xnor U2369 (N_2369,N_1680,N_1814);
nor U2370 (N_2370,N_1512,N_1705);
or U2371 (N_2371,N_1800,N_1796);
or U2372 (N_2372,N_1896,N_1655);
xor U2373 (N_2373,N_1820,N_1954);
or U2374 (N_2374,N_1766,N_1860);
nand U2375 (N_2375,N_1590,N_1921);
and U2376 (N_2376,N_1676,N_1621);
or U2377 (N_2377,N_1754,N_1869);
or U2378 (N_2378,N_1787,N_1840);
and U2379 (N_2379,N_1601,N_1698);
and U2380 (N_2380,N_1935,N_1771);
or U2381 (N_2381,N_1522,N_1608);
xor U2382 (N_2382,N_1884,N_1721);
or U2383 (N_2383,N_1673,N_1810);
or U2384 (N_2384,N_1573,N_1874);
xor U2385 (N_2385,N_1541,N_1778);
xnor U2386 (N_2386,N_1945,N_1589);
or U2387 (N_2387,N_1544,N_1790);
or U2388 (N_2388,N_1938,N_1969);
xnor U2389 (N_2389,N_1649,N_1696);
or U2390 (N_2390,N_1636,N_1529);
xnor U2391 (N_2391,N_1707,N_1530);
nor U2392 (N_2392,N_1899,N_1863);
nand U2393 (N_2393,N_1733,N_1984);
and U2394 (N_2394,N_1673,N_1696);
nor U2395 (N_2395,N_1829,N_1608);
and U2396 (N_2396,N_1738,N_1924);
or U2397 (N_2397,N_1912,N_1874);
xnor U2398 (N_2398,N_1815,N_1924);
and U2399 (N_2399,N_1773,N_1505);
nor U2400 (N_2400,N_1809,N_1848);
nor U2401 (N_2401,N_1767,N_1967);
or U2402 (N_2402,N_1736,N_1877);
or U2403 (N_2403,N_1817,N_1550);
nor U2404 (N_2404,N_1822,N_1763);
and U2405 (N_2405,N_1586,N_1678);
and U2406 (N_2406,N_1857,N_1508);
and U2407 (N_2407,N_1874,N_1839);
or U2408 (N_2408,N_1722,N_1555);
nor U2409 (N_2409,N_1988,N_1835);
or U2410 (N_2410,N_1942,N_1523);
nand U2411 (N_2411,N_1739,N_1843);
xor U2412 (N_2412,N_1583,N_1773);
nor U2413 (N_2413,N_1611,N_1833);
or U2414 (N_2414,N_1623,N_1607);
nand U2415 (N_2415,N_1631,N_1759);
xor U2416 (N_2416,N_1999,N_1625);
xor U2417 (N_2417,N_1710,N_1577);
xnor U2418 (N_2418,N_1692,N_1756);
nor U2419 (N_2419,N_1573,N_1886);
nand U2420 (N_2420,N_1747,N_1640);
and U2421 (N_2421,N_1660,N_1894);
xnor U2422 (N_2422,N_1783,N_1992);
and U2423 (N_2423,N_1866,N_1760);
or U2424 (N_2424,N_1824,N_1601);
or U2425 (N_2425,N_1950,N_1505);
nor U2426 (N_2426,N_1584,N_1603);
nor U2427 (N_2427,N_1803,N_1692);
xor U2428 (N_2428,N_1880,N_1540);
nand U2429 (N_2429,N_1786,N_1560);
nor U2430 (N_2430,N_1807,N_1936);
nor U2431 (N_2431,N_1710,N_1672);
and U2432 (N_2432,N_1926,N_1623);
or U2433 (N_2433,N_1652,N_1721);
or U2434 (N_2434,N_1610,N_1647);
and U2435 (N_2435,N_1902,N_1542);
and U2436 (N_2436,N_1821,N_1702);
and U2437 (N_2437,N_1554,N_1742);
or U2438 (N_2438,N_1993,N_1843);
nand U2439 (N_2439,N_1518,N_1552);
and U2440 (N_2440,N_1986,N_1651);
and U2441 (N_2441,N_1851,N_1664);
nand U2442 (N_2442,N_1920,N_1991);
and U2443 (N_2443,N_1599,N_1921);
nor U2444 (N_2444,N_1595,N_1628);
or U2445 (N_2445,N_1962,N_1569);
xnor U2446 (N_2446,N_1959,N_1574);
or U2447 (N_2447,N_1879,N_1944);
nand U2448 (N_2448,N_1579,N_1589);
xnor U2449 (N_2449,N_1822,N_1816);
nand U2450 (N_2450,N_1594,N_1743);
nor U2451 (N_2451,N_1697,N_1513);
nand U2452 (N_2452,N_1849,N_1653);
and U2453 (N_2453,N_1674,N_1780);
and U2454 (N_2454,N_1579,N_1927);
xor U2455 (N_2455,N_1853,N_1564);
xnor U2456 (N_2456,N_1937,N_1532);
or U2457 (N_2457,N_1840,N_1553);
nand U2458 (N_2458,N_1634,N_1808);
xor U2459 (N_2459,N_1521,N_1616);
and U2460 (N_2460,N_1728,N_1757);
or U2461 (N_2461,N_1560,N_1664);
nor U2462 (N_2462,N_1511,N_1540);
and U2463 (N_2463,N_1888,N_1767);
xor U2464 (N_2464,N_1783,N_1520);
xor U2465 (N_2465,N_1569,N_1577);
and U2466 (N_2466,N_1846,N_1810);
and U2467 (N_2467,N_1598,N_1918);
nand U2468 (N_2468,N_1894,N_1773);
or U2469 (N_2469,N_1821,N_1835);
nand U2470 (N_2470,N_1578,N_1541);
and U2471 (N_2471,N_1761,N_1609);
and U2472 (N_2472,N_1680,N_1641);
and U2473 (N_2473,N_1621,N_1957);
xnor U2474 (N_2474,N_1640,N_1568);
and U2475 (N_2475,N_1895,N_1818);
nand U2476 (N_2476,N_1880,N_1879);
and U2477 (N_2477,N_1859,N_1525);
nor U2478 (N_2478,N_1745,N_1533);
or U2479 (N_2479,N_1810,N_1850);
nand U2480 (N_2480,N_1693,N_1922);
and U2481 (N_2481,N_1653,N_1660);
nor U2482 (N_2482,N_1931,N_1992);
or U2483 (N_2483,N_1631,N_1704);
xnor U2484 (N_2484,N_1707,N_1569);
nand U2485 (N_2485,N_1569,N_1969);
and U2486 (N_2486,N_1894,N_1512);
nor U2487 (N_2487,N_1947,N_1604);
and U2488 (N_2488,N_1683,N_1728);
or U2489 (N_2489,N_1725,N_1666);
nor U2490 (N_2490,N_1502,N_1541);
nor U2491 (N_2491,N_1562,N_1902);
xor U2492 (N_2492,N_1790,N_1810);
xor U2493 (N_2493,N_1669,N_1909);
xnor U2494 (N_2494,N_1529,N_1777);
xnor U2495 (N_2495,N_1756,N_1640);
nor U2496 (N_2496,N_1933,N_1687);
and U2497 (N_2497,N_1894,N_1752);
nand U2498 (N_2498,N_1942,N_1987);
xnor U2499 (N_2499,N_1892,N_1971);
or U2500 (N_2500,N_2150,N_2236);
or U2501 (N_2501,N_2258,N_2168);
or U2502 (N_2502,N_2260,N_2494);
xor U2503 (N_2503,N_2390,N_2272);
and U2504 (N_2504,N_2283,N_2454);
or U2505 (N_2505,N_2297,N_2185);
nor U2506 (N_2506,N_2391,N_2405);
xnor U2507 (N_2507,N_2189,N_2426);
nand U2508 (N_2508,N_2292,N_2221);
and U2509 (N_2509,N_2481,N_2413);
nor U2510 (N_2510,N_2455,N_2135);
nand U2511 (N_2511,N_2395,N_2007);
or U2512 (N_2512,N_2015,N_2242);
nand U2513 (N_2513,N_2480,N_2336);
or U2514 (N_2514,N_2274,N_2371);
or U2515 (N_2515,N_2042,N_2203);
and U2516 (N_2516,N_2459,N_2347);
xor U2517 (N_2517,N_2416,N_2079);
nand U2518 (N_2518,N_2190,N_2499);
xnor U2519 (N_2519,N_2381,N_2198);
nand U2520 (N_2520,N_2224,N_2364);
nand U2521 (N_2521,N_2139,N_2112);
xor U2522 (N_2522,N_2180,N_2345);
or U2523 (N_2523,N_2490,N_2386);
nand U2524 (N_2524,N_2448,N_2475);
nor U2525 (N_2525,N_2473,N_2451);
and U2526 (N_2526,N_2360,N_2136);
nand U2527 (N_2527,N_2389,N_2038);
nor U2528 (N_2528,N_2172,N_2484);
or U2529 (N_2529,N_2308,N_2328);
xor U2530 (N_2530,N_2127,N_2465);
and U2531 (N_2531,N_2085,N_2115);
or U2532 (N_2532,N_2187,N_2338);
nor U2533 (N_2533,N_2287,N_2429);
xnor U2534 (N_2534,N_2011,N_2425);
xor U2535 (N_2535,N_2119,N_2398);
and U2536 (N_2536,N_2132,N_2331);
nor U2537 (N_2537,N_2109,N_2472);
nor U2538 (N_2538,N_2106,N_2232);
xnor U2539 (N_2539,N_2211,N_2148);
or U2540 (N_2540,N_2333,N_2262);
xor U2541 (N_2541,N_2419,N_2169);
or U2542 (N_2542,N_2313,N_2051);
nand U2543 (N_2543,N_2470,N_2254);
nand U2544 (N_2544,N_2036,N_2237);
nand U2545 (N_2545,N_2202,N_2267);
and U2546 (N_2546,N_2299,N_2259);
or U2547 (N_2547,N_2018,N_2305);
nand U2548 (N_2548,N_2463,N_2175);
nor U2549 (N_2549,N_2016,N_2197);
xnor U2550 (N_2550,N_2485,N_2279);
or U2551 (N_2551,N_2376,N_2466);
nor U2552 (N_2552,N_2092,N_2452);
nand U2553 (N_2553,N_2444,N_2143);
xor U2554 (N_2554,N_2446,N_2210);
nor U2555 (N_2555,N_2012,N_2076);
or U2556 (N_2556,N_2462,N_2072);
or U2557 (N_2557,N_2369,N_2029);
nor U2558 (N_2558,N_2204,N_2094);
nand U2559 (N_2559,N_2154,N_2177);
nand U2560 (N_2560,N_2370,N_2165);
xor U2561 (N_2561,N_2327,N_2002);
nor U2562 (N_2562,N_2403,N_2030);
nor U2563 (N_2563,N_2288,N_2492);
xnor U2564 (N_2564,N_2225,N_2184);
nand U2565 (N_2565,N_2301,N_2495);
nor U2566 (N_2566,N_2013,N_2447);
nand U2567 (N_2567,N_2006,N_2230);
or U2568 (N_2568,N_2393,N_2399);
nor U2569 (N_2569,N_2257,N_2087);
and U2570 (N_2570,N_2041,N_2003);
or U2571 (N_2571,N_2304,N_2082);
and U2572 (N_2572,N_2020,N_2129);
and U2573 (N_2573,N_2050,N_2430);
xnor U2574 (N_2574,N_2427,N_2032);
nand U2575 (N_2575,N_2471,N_2479);
nand U2576 (N_2576,N_2159,N_2397);
xnor U2577 (N_2577,N_2238,N_2021);
nor U2578 (N_2578,N_2083,N_2066);
xor U2579 (N_2579,N_2207,N_2432);
nor U2580 (N_2580,N_2057,N_2251);
xor U2581 (N_2581,N_2332,N_2483);
nor U2582 (N_2582,N_2081,N_2205);
or U2583 (N_2583,N_2061,N_2149);
nor U2584 (N_2584,N_2114,N_2497);
xor U2585 (N_2585,N_2354,N_2467);
nor U2586 (N_2586,N_2401,N_2163);
nand U2587 (N_2587,N_2035,N_2117);
or U2588 (N_2588,N_2124,N_2049);
nor U2589 (N_2589,N_2162,N_2241);
nor U2590 (N_2590,N_2441,N_2167);
nor U2591 (N_2591,N_2487,N_2385);
or U2592 (N_2592,N_2256,N_2340);
nand U2593 (N_2593,N_2017,N_2488);
and U2594 (N_2594,N_2378,N_2222);
nor U2595 (N_2595,N_2157,N_2145);
nand U2596 (N_2596,N_2218,N_2456);
or U2597 (N_2597,N_2152,N_2045);
or U2598 (N_2598,N_2265,N_2196);
nor U2599 (N_2599,N_2068,N_2384);
or U2600 (N_2600,N_2069,N_2247);
nand U2601 (N_2601,N_2239,N_2146);
and U2602 (N_2602,N_2240,N_2275);
and U2603 (N_2603,N_2276,N_2025);
nor U2604 (N_2604,N_2337,N_2439);
and U2605 (N_2605,N_2243,N_2442);
nor U2606 (N_2606,N_2043,N_2191);
nor U2607 (N_2607,N_2010,N_2449);
or U2608 (N_2608,N_2486,N_2101);
nand U2609 (N_2609,N_2402,N_2103);
nor U2610 (N_2610,N_2155,N_2080);
nand U2611 (N_2611,N_2458,N_2130);
and U2612 (N_2612,N_2248,N_2273);
nand U2613 (N_2613,N_2478,N_2496);
nand U2614 (N_2614,N_2435,N_2408);
nor U2615 (N_2615,N_2111,N_2353);
and U2616 (N_2616,N_2100,N_2414);
xnor U2617 (N_2617,N_2476,N_2291);
nor U2618 (N_2618,N_2176,N_2261);
nor U2619 (N_2619,N_2394,N_2412);
and U2620 (N_2620,N_2296,N_2290);
or U2621 (N_2621,N_2144,N_2311);
xnor U2622 (N_2622,N_2178,N_2437);
nor U2623 (N_2623,N_2110,N_2329);
nand U2624 (N_2624,N_2344,N_2063);
nor U2625 (N_2625,N_2026,N_2316);
and U2626 (N_2626,N_2253,N_2024);
nor U2627 (N_2627,N_2477,N_2460);
and U2628 (N_2628,N_2420,N_2491);
and U2629 (N_2629,N_2014,N_2269);
nor U2630 (N_2630,N_2365,N_2160);
nand U2631 (N_2631,N_2095,N_2493);
and U2632 (N_2632,N_2421,N_2088);
xnor U2633 (N_2633,N_2392,N_2411);
or U2634 (N_2634,N_2341,N_2450);
nor U2635 (N_2635,N_2404,N_2436);
or U2636 (N_2636,N_2352,N_2089);
nand U2637 (N_2637,N_2125,N_2141);
and U2638 (N_2638,N_2188,N_2334);
and U2639 (N_2639,N_2245,N_2443);
or U2640 (N_2640,N_2244,N_2346);
or U2641 (N_2641,N_2368,N_2406);
nor U2642 (N_2642,N_2031,N_2303);
and U2643 (N_2643,N_2415,N_2022);
and U2644 (N_2644,N_2396,N_2461);
or U2645 (N_2645,N_2161,N_2231);
or U2646 (N_2646,N_2055,N_2065);
and U2647 (N_2647,N_2064,N_2498);
nor U2648 (N_2648,N_2053,N_2326);
nand U2649 (N_2649,N_2116,N_2005);
nand U2650 (N_2650,N_2034,N_2489);
nand U2651 (N_2651,N_2009,N_2086);
xor U2652 (N_2652,N_2208,N_2004);
nor U2653 (N_2653,N_2330,N_2044);
and U2654 (N_2654,N_2315,N_2325);
nand U2655 (N_2655,N_2362,N_2090);
and U2656 (N_2656,N_2054,N_2246);
and U2657 (N_2657,N_2212,N_2128);
and U2658 (N_2658,N_2234,N_2037);
and U2659 (N_2659,N_2310,N_2373);
or U2660 (N_2660,N_2000,N_2309);
or U2661 (N_2661,N_2366,N_2343);
and U2662 (N_2662,N_2300,N_2118);
nor U2663 (N_2663,N_2201,N_2379);
nor U2664 (N_2664,N_2361,N_2131);
and U2665 (N_2665,N_2056,N_2335);
or U2666 (N_2666,N_2348,N_2046);
xor U2667 (N_2667,N_2209,N_2424);
nor U2668 (N_2668,N_2084,N_2445);
xnor U2669 (N_2669,N_2440,N_2280);
nand U2670 (N_2670,N_2339,N_2363);
and U2671 (N_2671,N_2105,N_2174);
or U2672 (N_2672,N_2070,N_2268);
or U2673 (N_2673,N_2423,N_2108);
nand U2674 (N_2674,N_2200,N_2133);
nand U2675 (N_2675,N_2284,N_2271);
or U2676 (N_2676,N_2324,N_2147);
nand U2677 (N_2677,N_2252,N_2302);
and U2678 (N_2678,N_2278,N_2097);
xnor U2679 (N_2679,N_2058,N_2048);
nor U2680 (N_2680,N_2377,N_2074);
and U2681 (N_2681,N_2409,N_2418);
nor U2682 (N_2682,N_2374,N_2121);
nand U2683 (N_2683,N_2314,N_2215);
xor U2684 (N_2684,N_2104,N_2289);
and U2685 (N_2685,N_2192,N_2220);
nand U2686 (N_2686,N_2073,N_2306);
and U2687 (N_2687,N_2319,N_2227);
xnor U2688 (N_2688,N_2216,N_2431);
and U2689 (N_2689,N_2033,N_2438);
nand U2690 (N_2690,N_2138,N_2023);
xnor U2691 (N_2691,N_2098,N_2170);
xor U2692 (N_2692,N_2342,N_2142);
xor U2693 (N_2693,N_2266,N_2349);
and U2694 (N_2694,N_2099,N_2482);
xor U2695 (N_2695,N_2350,N_2285);
nand U2696 (N_2696,N_2277,N_2195);
and U2697 (N_2697,N_2059,N_2270);
nand U2698 (N_2698,N_2213,N_2294);
nand U2699 (N_2699,N_2317,N_2356);
or U2700 (N_2700,N_2067,N_2249);
nor U2701 (N_2701,N_2153,N_2199);
nor U2702 (N_2702,N_2107,N_2250);
nand U2703 (N_2703,N_2226,N_2323);
and U2704 (N_2704,N_2214,N_2120);
nand U2705 (N_2705,N_2194,N_2134);
nand U2706 (N_2706,N_2286,N_2469);
or U2707 (N_2707,N_2182,N_2001);
and U2708 (N_2708,N_2183,N_2229);
nor U2709 (N_2709,N_2355,N_2040);
nor U2710 (N_2710,N_2282,N_2171);
nor U2711 (N_2711,N_2295,N_2400);
or U2712 (N_2712,N_2052,N_2358);
or U2713 (N_2713,N_2474,N_2410);
and U2714 (N_2714,N_2217,N_2096);
or U2715 (N_2715,N_2351,N_2235);
or U2716 (N_2716,N_2307,N_2428);
xnor U2717 (N_2717,N_2071,N_2164);
and U2718 (N_2718,N_2464,N_2359);
and U2719 (N_2719,N_2264,N_2047);
nor U2720 (N_2720,N_2422,N_2140);
xor U2721 (N_2721,N_2113,N_2223);
nor U2722 (N_2722,N_2102,N_2078);
nand U2723 (N_2723,N_2375,N_2434);
and U2724 (N_2724,N_2028,N_2219);
nor U2725 (N_2725,N_2060,N_2179);
xor U2726 (N_2726,N_2158,N_2263);
xnor U2727 (N_2727,N_2137,N_2321);
xnor U2728 (N_2728,N_2388,N_2453);
nor U2729 (N_2729,N_2298,N_2156);
and U2730 (N_2730,N_2312,N_2233);
or U2731 (N_2731,N_2322,N_2186);
and U2732 (N_2732,N_2091,N_2166);
or U2733 (N_2733,N_2126,N_2062);
or U2734 (N_2734,N_2019,N_2383);
nor U2735 (N_2735,N_2417,N_2193);
xnor U2736 (N_2736,N_2093,N_2433);
nor U2737 (N_2737,N_2255,N_2027);
xnor U2738 (N_2738,N_2382,N_2320);
xor U2739 (N_2739,N_2457,N_2077);
nand U2740 (N_2740,N_2075,N_2008);
xnor U2741 (N_2741,N_2293,N_2387);
xnor U2742 (N_2742,N_2039,N_2357);
nor U2743 (N_2743,N_2372,N_2367);
or U2744 (N_2744,N_2181,N_2123);
nor U2745 (N_2745,N_2281,N_2407);
nor U2746 (N_2746,N_2122,N_2151);
nand U2747 (N_2747,N_2173,N_2318);
nor U2748 (N_2748,N_2468,N_2380);
nor U2749 (N_2749,N_2228,N_2206);
or U2750 (N_2750,N_2445,N_2093);
nor U2751 (N_2751,N_2247,N_2261);
and U2752 (N_2752,N_2346,N_2428);
nor U2753 (N_2753,N_2140,N_2090);
nor U2754 (N_2754,N_2415,N_2081);
or U2755 (N_2755,N_2194,N_2286);
xor U2756 (N_2756,N_2294,N_2031);
nand U2757 (N_2757,N_2136,N_2327);
nand U2758 (N_2758,N_2462,N_2075);
and U2759 (N_2759,N_2125,N_2348);
or U2760 (N_2760,N_2179,N_2462);
and U2761 (N_2761,N_2492,N_2060);
nor U2762 (N_2762,N_2251,N_2052);
or U2763 (N_2763,N_2226,N_2138);
nand U2764 (N_2764,N_2350,N_2333);
and U2765 (N_2765,N_2294,N_2445);
xnor U2766 (N_2766,N_2475,N_2324);
nor U2767 (N_2767,N_2495,N_2393);
nand U2768 (N_2768,N_2242,N_2161);
nand U2769 (N_2769,N_2360,N_2444);
xor U2770 (N_2770,N_2493,N_2197);
nor U2771 (N_2771,N_2263,N_2470);
nand U2772 (N_2772,N_2203,N_2208);
and U2773 (N_2773,N_2295,N_2296);
and U2774 (N_2774,N_2349,N_2434);
or U2775 (N_2775,N_2372,N_2239);
and U2776 (N_2776,N_2364,N_2160);
nand U2777 (N_2777,N_2490,N_2414);
or U2778 (N_2778,N_2414,N_2319);
xnor U2779 (N_2779,N_2389,N_2360);
or U2780 (N_2780,N_2369,N_2014);
nand U2781 (N_2781,N_2170,N_2149);
nor U2782 (N_2782,N_2399,N_2036);
nand U2783 (N_2783,N_2060,N_2303);
or U2784 (N_2784,N_2173,N_2472);
nand U2785 (N_2785,N_2426,N_2382);
or U2786 (N_2786,N_2296,N_2483);
nor U2787 (N_2787,N_2294,N_2420);
xnor U2788 (N_2788,N_2353,N_2403);
nor U2789 (N_2789,N_2046,N_2448);
nor U2790 (N_2790,N_2489,N_2242);
xor U2791 (N_2791,N_2070,N_2165);
or U2792 (N_2792,N_2386,N_2304);
or U2793 (N_2793,N_2395,N_2180);
or U2794 (N_2794,N_2176,N_2111);
xnor U2795 (N_2795,N_2138,N_2063);
nor U2796 (N_2796,N_2395,N_2465);
or U2797 (N_2797,N_2272,N_2426);
xnor U2798 (N_2798,N_2102,N_2088);
xor U2799 (N_2799,N_2376,N_2178);
or U2800 (N_2800,N_2426,N_2352);
and U2801 (N_2801,N_2351,N_2047);
xor U2802 (N_2802,N_2030,N_2103);
nand U2803 (N_2803,N_2143,N_2016);
and U2804 (N_2804,N_2316,N_2169);
xnor U2805 (N_2805,N_2055,N_2233);
or U2806 (N_2806,N_2324,N_2262);
nor U2807 (N_2807,N_2395,N_2038);
nor U2808 (N_2808,N_2274,N_2072);
or U2809 (N_2809,N_2315,N_2390);
or U2810 (N_2810,N_2047,N_2169);
xnor U2811 (N_2811,N_2034,N_2198);
and U2812 (N_2812,N_2245,N_2165);
and U2813 (N_2813,N_2416,N_2259);
or U2814 (N_2814,N_2353,N_2317);
and U2815 (N_2815,N_2128,N_2152);
nand U2816 (N_2816,N_2422,N_2000);
or U2817 (N_2817,N_2029,N_2251);
nand U2818 (N_2818,N_2123,N_2047);
nor U2819 (N_2819,N_2481,N_2132);
xnor U2820 (N_2820,N_2407,N_2317);
nand U2821 (N_2821,N_2406,N_2077);
nor U2822 (N_2822,N_2424,N_2033);
nand U2823 (N_2823,N_2207,N_2192);
nand U2824 (N_2824,N_2392,N_2127);
nor U2825 (N_2825,N_2013,N_2282);
nand U2826 (N_2826,N_2065,N_2118);
and U2827 (N_2827,N_2403,N_2357);
nand U2828 (N_2828,N_2412,N_2427);
xnor U2829 (N_2829,N_2068,N_2391);
xnor U2830 (N_2830,N_2023,N_2409);
nor U2831 (N_2831,N_2320,N_2124);
or U2832 (N_2832,N_2090,N_2109);
and U2833 (N_2833,N_2209,N_2283);
and U2834 (N_2834,N_2070,N_2482);
and U2835 (N_2835,N_2009,N_2136);
or U2836 (N_2836,N_2247,N_2338);
xor U2837 (N_2837,N_2355,N_2228);
nand U2838 (N_2838,N_2401,N_2031);
nand U2839 (N_2839,N_2406,N_2476);
nand U2840 (N_2840,N_2420,N_2006);
nand U2841 (N_2841,N_2177,N_2359);
and U2842 (N_2842,N_2321,N_2205);
xnor U2843 (N_2843,N_2340,N_2071);
nor U2844 (N_2844,N_2058,N_2434);
xnor U2845 (N_2845,N_2157,N_2480);
nand U2846 (N_2846,N_2221,N_2416);
nor U2847 (N_2847,N_2073,N_2107);
or U2848 (N_2848,N_2402,N_2474);
nand U2849 (N_2849,N_2096,N_2059);
and U2850 (N_2850,N_2127,N_2171);
nor U2851 (N_2851,N_2042,N_2006);
or U2852 (N_2852,N_2343,N_2347);
nand U2853 (N_2853,N_2028,N_2488);
nand U2854 (N_2854,N_2275,N_2494);
nor U2855 (N_2855,N_2407,N_2243);
xor U2856 (N_2856,N_2097,N_2289);
or U2857 (N_2857,N_2492,N_2052);
xnor U2858 (N_2858,N_2245,N_2239);
xor U2859 (N_2859,N_2293,N_2452);
or U2860 (N_2860,N_2068,N_2458);
nor U2861 (N_2861,N_2423,N_2166);
nand U2862 (N_2862,N_2442,N_2330);
nand U2863 (N_2863,N_2374,N_2352);
and U2864 (N_2864,N_2357,N_2375);
nor U2865 (N_2865,N_2485,N_2272);
and U2866 (N_2866,N_2284,N_2406);
and U2867 (N_2867,N_2392,N_2135);
nand U2868 (N_2868,N_2065,N_2432);
and U2869 (N_2869,N_2250,N_2445);
and U2870 (N_2870,N_2062,N_2054);
and U2871 (N_2871,N_2308,N_2421);
xor U2872 (N_2872,N_2053,N_2394);
nand U2873 (N_2873,N_2209,N_2397);
or U2874 (N_2874,N_2087,N_2028);
nand U2875 (N_2875,N_2472,N_2386);
nand U2876 (N_2876,N_2248,N_2315);
nand U2877 (N_2877,N_2058,N_2310);
xor U2878 (N_2878,N_2306,N_2380);
xor U2879 (N_2879,N_2427,N_2083);
nor U2880 (N_2880,N_2450,N_2016);
nor U2881 (N_2881,N_2384,N_2438);
and U2882 (N_2882,N_2268,N_2116);
xor U2883 (N_2883,N_2482,N_2297);
or U2884 (N_2884,N_2233,N_2198);
nor U2885 (N_2885,N_2005,N_2099);
or U2886 (N_2886,N_2331,N_2409);
xnor U2887 (N_2887,N_2166,N_2451);
nor U2888 (N_2888,N_2214,N_2497);
xor U2889 (N_2889,N_2118,N_2015);
or U2890 (N_2890,N_2493,N_2085);
or U2891 (N_2891,N_2262,N_2359);
xnor U2892 (N_2892,N_2224,N_2043);
xnor U2893 (N_2893,N_2336,N_2088);
nor U2894 (N_2894,N_2122,N_2331);
nor U2895 (N_2895,N_2256,N_2180);
or U2896 (N_2896,N_2412,N_2402);
xnor U2897 (N_2897,N_2239,N_2288);
and U2898 (N_2898,N_2360,N_2271);
nor U2899 (N_2899,N_2087,N_2282);
nand U2900 (N_2900,N_2354,N_2458);
xnor U2901 (N_2901,N_2431,N_2333);
xor U2902 (N_2902,N_2194,N_2284);
or U2903 (N_2903,N_2475,N_2468);
xor U2904 (N_2904,N_2172,N_2299);
xor U2905 (N_2905,N_2313,N_2008);
nand U2906 (N_2906,N_2333,N_2120);
nor U2907 (N_2907,N_2337,N_2072);
or U2908 (N_2908,N_2091,N_2193);
or U2909 (N_2909,N_2284,N_2332);
or U2910 (N_2910,N_2133,N_2300);
nor U2911 (N_2911,N_2016,N_2279);
xor U2912 (N_2912,N_2451,N_2268);
nand U2913 (N_2913,N_2447,N_2304);
xnor U2914 (N_2914,N_2035,N_2127);
or U2915 (N_2915,N_2405,N_2189);
nor U2916 (N_2916,N_2056,N_2452);
xnor U2917 (N_2917,N_2125,N_2049);
or U2918 (N_2918,N_2316,N_2269);
and U2919 (N_2919,N_2173,N_2054);
and U2920 (N_2920,N_2104,N_2252);
xnor U2921 (N_2921,N_2229,N_2304);
and U2922 (N_2922,N_2304,N_2117);
nor U2923 (N_2923,N_2499,N_2329);
xor U2924 (N_2924,N_2481,N_2211);
nand U2925 (N_2925,N_2116,N_2436);
or U2926 (N_2926,N_2092,N_2182);
xor U2927 (N_2927,N_2420,N_2186);
nor U2928 (N_2928,N_2456,N_2415);
nor U2929 (N_2929,N_2154,N_2331);
xor U2930 (N_2930,N_2206,N_2334);
nand U2931 (N_2931,N_2378,N_2149);
xnor U2932 (N_2932,N_2013,N_2418);
xnor U2933 (N_2933,N_2288,N_2041);
xor U2934 (N_2934,N_2215,N_2037);
or U2935 (N_2935,N_2447,N_2248);
nand U2936 (N_2936,N_2330,N_2147);
xor U2937 (N_2937,N_2186,N_2363);
or U2938 (N_2938,N_2352,N_2363);
and U2939 (N_2939,N_2270,N_2296);
or U2940 (N_2940,N_2382,N_2197);
xor U2941 (N_2941,N_2125,N_2351);
and U2942 (N_2942,N_2004,N_2290);
and U2943 (N_2943,N_2479,N_2327);
nor U2944 (N_2944,N_2219,N_2349);
nor U2945 (N_2945,N_2235,N_2496);
nand U2946 (N_2946,N_2332,N_2203);
or U2947 (N_2947,N_2404,N_2439);
nand U2948 (N_2948,N_2087,N_2185);
and U2949 (N_2949,N_2446,N_2022);
or U2950 (N_2950,N_2244,N_2389);
or U2951 (N_2951,N_2076,N_2158);
nor U2952 (N_2952,N_2045,N_2206);
and U2953 (N_2953,N_2401,N_2297);
xor U2954 (N_2954,N_2108,N_2012);
xnor U2955 (N_2955,N_2326,N_2451);
or U2956 (N_2956,N_2222,N_2371);
nand U2957 (N_2957,N_2337,N_2441);
or U2958 (N_2958,N_2082,N_2291);
or U2959 (N_2959,N_2498,N_2339);
or U2960 (N_2960,N_2177,N_2021);
nand U2961 (N_2961,N_2344,N_2385);
xor U2962 (N_2962,N_2057,N_2462);
nand U2963 (N_2963,N_2236,N_2115);
nor U2964 (N_2964,N_2047,N_2052);
nand U2965 (N_2965,N_2196,N_2262);
xor U2966 (N_2966,N_2325,N_2064);
or U2967 (N_2967,N_2312,N_2405);
nor U2968 (N_2968,N_2045,N_2125);
and U2969 (N_2969,N_2129,N_2097);
nor U2970 (N_2970,N_2040,N_2124);
xor U2971 (N_2971,N_2319,N_2274);
nor U2972 (N_2972,N_2043,N_2063);
xor U2973 (N_2973,N_2111,N_2103);
nand U2974 (N_2974,N_2138,N_2215);
and U2975 (N_2975,N_2100,N_2205);
xnor U2976 (N_2976,N_2459,N_2041);
nor U2977 (N_2977,N_2479,N_2030);
or U2978 (N_2978,N_2410,N_2213);
or U2979 (N_2979,N_2379,N_2036);
and U2980 (N_2980,N_2108,N_2057);
and U2981 (N_2981,N_2062,N_2323);
or U2982 (N_2982,N_2432,N_2048);
or U2983 (N_2983,N_2164,N_2231);
and U2984 (N_2984,N_2323,N_2361);
nor U2985 (N_2985,N_2352,N_2493);
or U2986 (N_2986,N_2422,N_2056);
nor U2987 (N_2987,N_2122,N_2303);
nor U2988 (N_2988,N_2358,N_2369);
or U2989 (N_2989,N_2007,N_2286);
nand U2990 (N_2990,N_2461,N_2418);
xnor U2991 (N_2991,N_2371,N_2003);
and U2992 (N_2992,N_2399,N_2090);
nor U2993 (N_2993,N_2268,N_2343);
nand U2994 (N_2994,N_2294,N_2435);
nor U2995 (N_2995,N_2205,N_2168);
or U2996 (N_2996,N_2445,N_2402);
or U2997 (N_2997,N_2449,N_2107);
nand U2998 (N_2998,N_2217,N_2484);
xnor U2999 (N_2999,N_2415,N_2102);
nor UO_0 (O_0,N_2882,N_2886);
and UO_1 (O_1,N_2787,N_2977);
and UO_2 (O_2,N_2654,N_2723);
nor UO_3 (O_3,N_2692,N_2592);
xor UO_4 (O_4,N_2552,N_2546);
xnor UO_5 (O_5,N_2567,N_2668);
xor UO_6 (O_6,N_2768,N_2855);
or UO_7 (O_7,N_2843,N_2842);
nand UO_8 (O_8,N_2603,N_2973);
nor UO_9 (O_9,N_2719,N_2921);
and UO_10 (O_10,N_2744,N_2745);
or UO_11 (O_11,N_2816,N_2953);
and UO_12 (O_12,N_2697,N_2534);
nand UO_13 (O_13,N_2937,N_2758);
and UO_14 (O_14,N_2608,N_2877);
nor UO_15 (O_15,N_2941,N_2845);
and UO_16 (O_16,N_2818,N_2984);
and UO_17 (O_17,N_2897,N_2677);
or UO_18 (O_18,N_2620,N_2743);
nor UO_19 (O_19,N_2910,N_2658);
xor UO_20 (O_20,N_2811,N_2720);
or UO_21 (O_21,N_2789,N_2601);
and UO_22 (O_22,N_2988,N_2721);
or UO_23 (O_23,N_2571,N_2894);
nor UO_24 (O_24,N_2929,N_2577);
nand UO_25 (O_25,N_2597,N_2547);
or UO_26 (O_26,N_2793,N_2559);
nor UO_27 (O_27,N_2610,N_2670);
nand UO_28 (O_28,N_2504,N_2702);
or UO_29 (O_29,N_2801,N_2932);
xnor UO_30 (O_30,N_2591,N_2565);
nor UO_31 (O_31,N_2675,N_2931);
xnor UO_32 (O_32,N_2917,N_2604);
nor UO_33 (O_33,N_2649,N_2735);
xnor UO_34 (O_34,N_2911,N_2706);
or UO_35 (O_35,N_2667,N_2684);
xor UO_36 (O_36,N_2536,N_2933);
xor UO_37 (O_37,N_2802,N_2583);
xor UO_38 (O_38,N_2934,N_2893);
nor UO_39 (O_39,N_2832,N_2656);
or UO_40 (O_40,N_2874,N_2650);
nand UO_41 (O_41,N_2781,N_2724);
nor UO_42 (O_42,N_2713,N_2967);
and UO_43 (O_43,N_2507,N_2896);
or UO_44 (O_44,N_2772,N_2646);
and UO_45 (O_45,N_2541,N_2555);
nand UO_46 (O_46,N_2639,N_2944);
or UO_47 (O_47,N_2727,N_2776);
xor UO_48 (O_48,N_2873,N_2867);
nand UO_49 (O_49,N_2965,N_2773);
xnor UO_50 (O_50,N_2746,N_2834);
or UO_51 (O_51,N_2605,N_2569);
and UO_52 (O_52,N_2810,N_2957);
or UO_53 (O_53,N_2598,N_2714);
nand UO_54 (O_54,N_2815,N_2794);
or UO_55 (O_55,N_2521,N_2846);
nand UO_56 (O_56,N_2553,N_2586);
xnor UO_57 (O_57,N_2587,N_2860);
nand UO_58 (O_58,N_2892,N_2596);
or UO_59 (O_59,N_2737,N_2628);
or UO_60 (O_60,N_2759,N_2859);
and UO_61 (O_61,N_2829,N_2606);
nor UO_62 (O_62,N_2854,N_2875);
and UO_63 (O_63,N_2537,N_2819);
nor UO_64 (O_64,N_2919,N_2958);
nor UO_65 (O_65,N_2607,N_2907);
or UO_66 (O_66,N_2991,N_2618);
or UO_67 (O_67,N_2733,N_2865);
nand UO_68 (O_68,N_2916,N_2522);
and UO_69 (O_69,N_2696,N_2614);
nand UO_70 (O_70,N_2764,N_2835);
and UO_71 (O_71,N_2572,N_2978);
nor UO_72 (O_72,N_2732,N_2870);
xnor UO_73 (O_73,N_2661,N_2568);
xnor UO_74 (O_74,N_2699,N_2518);
nand UO_75 (O_75,N_2756,N_2726);
xor UO_76 (O_76,N_2852,N_2543);
nor UO_77 (O_77,N_2716,N_2970);
nand UO_78 (O_78,N_2891,N_2955);
xnor UO_79 (O_79,N_2695,N_2969);
and UO_80 (O_80,N_2950,N_2729);
nor UO_81 (O_81,N_2906,N_2943);
xnor UO_82 (O_82,N_2954,N_2889);
xnor UO_83 (O_83,N_2674,N_2980);
nand UO_84 (O_84,N_2752,N_2928);
nor UO_85 (O_85,N_2836,N_2786);
xor UO_86 (O_86,N_2902,N_2655);
nand UO_87 (O_87,N_2579,N_2806);
and UO_88 (O_88,N_2853,N_2997);
or UO_89 (O_89,N_2866,N_2775);
or UO_90 (O_90,N_2848,N_2833);
and UO_91 (O_91,N_2709,N_2666);
nand UO_92 (O_92,N_2679,N_2993);
nor UO_93 (O_93,N_2613,N_2558);
xnor UO_94 (O_94,N_2599,N_2619);
xnor UO_95 (O_95,N_2615,N_2523);
xnor UO_96 (O_96,N_2871,N_2839);
or UO_97 (O_97,N_2557,N_2827);
xor UO_98 (O_98,N_2771,N_2672);
nand UO_99 (O_99,N_2517,N_2511);
xnor UO_100 (O_100,N_2918,N_2982);
and UO_101 (O_101,N_2840,N_2738);
or UO_102 (O_102,N_2938,N_2635);
nand UO_103 (O_103,N_2509,N_2798);
nor UO_104 (O_104,N_2638,N_2705);
nor UO_105 (O_105,N_2817,N_2535);
nand UO_106 (O_106,N_2778,N_2609);
nor UO_107 (O_107,N_2685,N_2627);
xor UO_108 (O_108,N_2964,N_2570);
and UO_109 (O_109,N_2593,N_2660);
xnor UO_110 (O_110,N_2711,N_2508);
and UO_111 (O_111,N_2942,N_2981);
or UO_112 (O_112,N_2945,N_2566);
and UO_113 (O_113,N_2971,N_2883);
nor UO_114 (O_114,N_2922,N_2899);
nand UO_115 (O_115,N_2576,N_2750);
or UO_116 (O_116,N_2755,N_2687);
xnor UO_117 (O_117,N_2512,N_2653);
and UO_118 (O_118,N_2799,N_2616);
and UO_119 (O_119,N_2779,N_2968);
or UO_120 (O_120,N_2531,N_2515);
nand UO_121 (O_121,N_2588,N_2795);
nand UO_122 (O_122,N_2636,N_2584);
nor UO_123 (O_123,N_2644,N_2528);
and UO_124 (O_124,N_2760,N_2510);
or UO_125 (O_125,N_2533,N_2939);
nand UO_126 (O_126,N_2920,N_2946);
and UO_127 (O_127,N_2514,N_2662);
nand UO_128 (O_128,N_2647,N_2952);
nor UO_129 (O_129,N_2851,N_2573);
nand UO_130 (O_130,N_2757,N_2673);
and UO_131 (O_131,N_2739,N_2863);
or UO_132 (O_132,N_2602,N_2904);
nand UO_133 (O_133,N_2700,N_2751);
and UO_134 (O_134,N_2761,N_2783);
xor UO_135 (O_135,N_2722,N_2825);
or UO_136 (O_136,N_2671,N_2689);
nor UO_137 (O_137,N_2502,N_2809);
nand UO_138 (O_138,N_2903,N_2681);
or UO_139 (O_139,N_2625,N_2540);
nand UO_140 (O_140,N_2949,N_2680);
nand UO_141 (O_141,N_2525,N_2763);
nor UO_142 (O_142,N_2748,N_2561);
nor UO_143 (O_143,N_2999,N_2847);
xnor UO_144 (O_144,N_2913,N_2935);
nor UO_145 (O_145,N_2730,N_2741);
or UO_146 (O_146,N_2753,N_2693);
xnor UO_147 (O_147,N_2669,N_2790);
nor UO_148 (O_148,N_2611,N_2595);
nor UO_149 (O_149,N_2962,N_2849);
nor UO_150 (O_150,N_2526,N_2823);
xnor UO_151 (O_151,N_2972,N_2959);
nor UO_152 (O_152,N_2563,N_2814);
and UO_153 (O_153,N_2506,N_2538);
nand UO_154 (O_154,N_2881,N_2983);
nor UO_155 (O_155,N_2879,N_2861);
nand UO_156 (O_156,N_2960,N_2664);
or UO_157 (O_157,N_2864,N_2912);
nand UO_158 (O_158,N_2782,N_2698);
or UO_159 (O_159,N_2905,N_2624);
xnor UO_160 (O_160,N_2927,N_2898);
and UO_161 (O_161,N_2678,N_2947);
nand UO_162 (O_162,N_2986,N_2956);
nand UO_163 (O_163,N_2708,N_2803);
xnor UO_164 (O_164,N_2651,N_2976);
nand UO_165 (O_165,N_2989,N_2712);
or UO_166 (O_166,N_2808,N_2725);
or UO_167 (O_167,N_2856,N_2837);
or UO_168 (O_168,N_2631,N_2715);
nand UO_169 (O_169,N_2564,N_2749);
xnor UO_170 (O_170,N_2996,N_2686);
xor UO_171 (O_171,N_2747,N_2582);
nor UO_172 (O_172,N_2915,N_2626);
nor UO_173 (O_173,N_2797,N_2994);
xnor UO_174 (O_174,N_2767,N_2629);
and UO_175 (O_175,N_2831,N_2728);
nor UO_176 (O_176,N_2926,N_2807);
and UO_177 (O_177,N_2858,N_2520);
and UO_178 (O_178,N_2643,N_2844);
xnor UO_179 (O_179,N_2961,N_2805);
and UO_180 (O_180,N_2812,N_2914);
or UO_181 (O_181,N_2524,N_2513);
and UO_182 (O_182,N_2788,N_2551);
xor UO_183 (O_183,N_2880,N_2769);
and UO_184 (O_184,N_2500,N_2731);
and UO_185 (O_185,N_2574,N_2545);
nor UO_186 (O_186,N_2501,N_2539);
or UO_187 (O_187,N_2633,N_2777);
and UO_188 (O_188,N_2657,N_2532);
nand UO_189 (O_189,N_2641,N_2703);
or UO_190 (O_190,N_2663,N_2718);
nand UO_191 (O_191,N_2659,N_2742);
and UO_192 (O_192,N_2857,N_2530);
nor UO_193 (O_193,N_2908,N_2979);
nor UO_194 (O_194,N_2734,N_2717);
and UO_195 (O_195,N_2707,N_2640);
xnor UO_196 (O_196,N_2974,N_2796);
nand UO_197 (O_197,N_2765,N_2888);
nand UO_198 (O_198,N_2923,N_2940);
or UO_199 (O_199,N_2998,N_2648);
xor UO_200 (O_200,N_2838,N_2556);
and UO_201 (O_201,N_2590,N_2694);
nor UO_202 (O_202,N_2822,N_2930);
xnor UO_203 (O_203,N_2754,N_2527);
or UO_204 (O_204,N_2529,N_2951);
or UO_205 (O_205,N_2623,N_2544);
and UO_206 (O_206,N_2887,N_2548);
or UO_207 (O_207,N_2676,N_2876);
and UO_208 (O_208,N_2804,N_2740);
nand UO_209 (O_209,N_2762,N_2701);
xnor UO_210 (O_210,N_2990,N_2542);
xor UO_211 (O_211,N_2813,N_2683);
and UO_212 (O_212,N_2630,N_2652);
and UO_213 (O_213,N_2909,N_2868);
nand UO_214 (O_214,N_2987,N_2828);
nor UO_215 (O_215,N_2503,N_2780);
nand UO_216 (O_216,N_2617,N_2560);
nor UO_217 (O_217,N_2800,N_2600);
and UO_218 (O_218,N_2900,N_2637);
and UO_219 (O_219,N_2691,N_2594);
nand UO_220 (O_220,N_2784,N_2690);
nand UO_221 (O_221,N_2885,N_2821);
and UO_222 (O_222,N_2792,N_2995);
and UO_223 (O_223,N_2830,N_2710);
xor UO_224 (O_224,N_2966,N_2901);
or UO_225 (O_225,N_2622,N_2575);
nor UO_226 (O_226,N_2585,N_2766);
or UO_227 (O_227,N_2704,N_2890);
nand UO_228 (O_228,N_2554,N_2872);
nor UO_229 (O_229,N_2820,N_2884);
or UO_230 (O_230,N_2634,N_2862);
or UO_231 (O_231,N_2774,N_2785);
nand UO_232 (O_232,N_2841,N_2824);
nand UO_233 (O_233,N_2642,N_2682);
nor UO_234 (O_234,N_2975,N_2621);
nor UO_235 (O_235,N_2632,N_2519);
nor UO_236 (O_236,N_2581,N_2578);
xnor UO_237 (O_237,N_2770,N_2791);
nand UO_238 (O_238,N_2612,N_2869);
or UO_239 (O_239,N_2826,N_2924);
xor UO_240 (O_240,N_2562,N_2985);
and UO_241 (O_241,N_2665,N_2936);
xnor UO_242 (O_242,N_2850,N_2992);
xor UO_243 (O_243,N_2736,N_2505);
or UO_244 (O_244,N_2925,N_2963);
nor UO_245 (O_245,N_2645,N_2895);
or UO_246 (O_246,N_2550,N_2878);
and UO_247 (O_247,N_2580,N_2516);
and UO_248 (O_248,N_2948,N_2589);
or UO_249 (O_249,N_2549,N_2688);
and UO_250 (O_250,N_2579,N_2618);
nor UO_251 (O_251,N_2753,N_2825);
nor UO_252 (O_252,N_2811,N_2852);
nor UO_253 (O_253,N_2729,N_2814);
or UO_254 (O_254,N_2782,N_2743);
and UO_255 (O_255,N_2517,N_2687);
nor UO_256 (O_256,N_2804,N_2618);
or UO_257 (O_257,N_2507,N_2611);
xor UO_258 (O_258,N_2794,N_2698);
nor UO_259 (O_259,N_2988,N_2777);
xnor UO_260 (O_260,N_2818,N_2663);
and UO_261 (O_261,N_2860,N_2599);
nand UO_262 (O_262,N_2503,N_2863);
nor UO_263 (O_263,N_2781,N_2597);
and UO_264 (O_264,N_2926,N_2673);
nor UO_265 (O_265,N_2841,N_2811);
or UO_266 (O_266,N_2927,N_2925);
or UO_267 (O_267,N_2818,N_2960);
and UO_268 (O_268,N_2619,N_2715);
xor UO_269 (O_269,N_2645,N_2925);
and UO_270 (O_270,N_2549,N_2647);
nor UO_271 (O_271,N_2852,N_2941);
xnor UO_272 (O_272,N_2515,N_2925);
xnor UO_273 (O_273,N_2789,N_2584);
nor UO_274 (O_274,N_2867,N_2632);
or UO_275 (O_275,N_2692,N_2694);
and UO_276 (O_276,N_2529,N_2722);
nand UO_277 (O_277,N_2700,N_2915);
nor UO_278 (O_278,N_2731,N_2849);
nand UO_279 (O_279,N_2553,N_2618);
and UO_280 (O_280,N_2993,N_2911);
or UO_281 (O_281,N_2574,N_2859);
or UO_282 (O_282,N_2943,N_2968);
or UO_283 (O_283,N_2586,N_2845);
nor UO_284 (O_284,N_2683,N_2558);
xor UO_285 (O_285,N_2833,N_2757);
nand UO_286 (O_286,N_2740,N_2974);
nand UO_287 (O_287,N_2656,N_2755);
and UO_288 (O_288,N_2973,N_2894);
and UO_289 (O_289,N_2688,N_2682);
and UO_290 (O_290,N_2990,N_2597);
nor UO_291 (O_291,N_2729,N_2794);
and UO_292 (O_292,N_2692,N_2626);
and UO_293 (O_293,N_2863,N_2605);
nor UO_294 (O_294,N_2738,N_2980);
and UO_295 (O_295,N_2582,N_2556);
xor UO_296 (O_296,N_2682,N_2887);
xor UO_297 (O_297,N_2595,N_2505);
nand UO_298 (O_298,N_2803,N_2939);
or UO_299 (O_299,N_2863,N_2829);
nor UO_300 (O_300,N_2987,N_2981);
xor UO_301 (O_301,N_2904,N_2883);
and UO_302 (O_302,N_2742,N_2876);
xnor UO_303 (O_303,N_2528,N_2547);
and UO_304 (O_304,N_2946,N_2980);
nor UO_305 (O_305,N_2831,N_2810);
and UO_306 (O_306,N_2849,N_2787);
or UO_307 (O_307,N_2573,N_2959);
nand UO_308 (O_308,N_2556,N_2607);
or UO_309 (O_309,N_2977,N_2668);
nand UO_310 (O_310,N_2614,N_2649);
nand UO_311 (O_311,N_2510,N_2984);
and UO_312 (O_312,N_2975,N_2750);
xnor UO_313 (O_313,N_2706,N_2762);
xor UO_314 (O_314,N_2904,N_2738);
and UO_315 (O_315,N_2683,N_2852);
nor UO_316 (O_316,N_2710,N_2645);
xor UO_317 (O_317,N_2537,N_2916);
xnor UO_318 (O_318,N_2513,N_2924);
xor UO_319 (O_319,N_2678,N_2714);
nand UO_320 (O_320,N_2896,N_2570);
xnor UO_321 (O_321,N_2718,N_2986);
nand UO_322 (O_322,N_2773,N_2920);
or UO_323 (O_323,N_2759,N_2765);
or UO_324 (O_324,N_2559,N_2730);
nor UO_325 (O_325,N_2838,N_2821);
or UO_326 (O_326,N_2776,N_2996);
and UO_327 (O_327,N_2704,N_2655);
and UO_328 (O_328,N_2566,N_2624);
and UO_329 (O_329,N_2576,N_2717);
nor UO_330 (O_330,N_2817,N_2760);
nand UO_331 (O_331,N_2858,N_2919);
xor UO_332 (O_332,N_2934,N_2605);
or UO_333 (O_333,N_2910,N_2706);
nand UO_334 (O_334,N_2665,N_2627);
xor UO_335 (O_335,N_2661,N_2768);
or UO_336 (O_336,N_2662,N_2614);
or UO_337 (O_337,N_2635,N_2516);
nor UO_338 (O_338,N_2652,N_2588);
nand UO_339 (O_339,N_2725,N_2694);
or UO_340 (O_340,N_2880,N_2639);
xnor UO_341 (O_341,N_2792,N_2969);
and UO_342 (O_342,N_2999,N_2519);
and UO_343 (O_343,N_2837,N_2698);
xnor UO_344 (O_344,N_2847,N_2831);
and UO_345 (O_345,N_2810,N_2500);
and UO_346 (O_346,N_2831,N_2504);
xor UO_347 (O_347,N_2821,N_2708);
and UO_348 (O_348,N_2843,N_2923);
xnor UO_349 (O_349,N_2825,N_2828);
and UO_350 (O_350,N_2978,N_2536);
or UO_351 (O_351,N_2645,N_2518);
nand UO_352 (O_352,N_2749,N_2584);
or UO_353 (O_353,N_2547,N_2841);
xnor UO_354 (O_354,N_2629,N_2545);
nand UO_355 (O_355,N_2791,N_2754);
or UO_356 (O_356,N_2858,N_2762);
nor UO_357 (O_357,N_2712,N_2825);
and UO_358 (O_358,N_2585,N_2873);
nor UO_359 (O_359,N_2541,N_2895);
or UO_360 (O_360,N_2989,N_2893);
nand UO_361 (O_361,N_2629,N_2719);
xor UO_362 (O_362,N_2693,N_2509);
nor UO_363 (O_363,N_2597,N_2929);
xor UO_364 (O_364,N_2530,N_2930);
nand UO_365 (O_365,N_2504,N_2687);
xnor UO_366 (O_366,N_2517,N_2888);
nor UO_367 (O_367,N_2610,N_2976);
or UO_368 (O_368,N_2646,N_2706);
xor UO_369 (O_369,N_2749,N_2545);
nand UO_370 (O_370,N_2852,N_2685);
nand UO_371 (O_371,N_2918,N_2998);
nor UO_372 (O_372,N_2737,N_2939);
and UO_373 (O_373,N_2596,N_2823);
or UO_374 (O_374,N_2790,N_2981);
nand UO_375 (O_375,N_2561,N_2744);
or UO_376 (O_376,N_2821,N_2510);
xnor UO_377 (O_377,N_2753,N_2821);
nand UO_378 (O_378,N_2725,N_2749);
and UO_379 (O_379,N_2786,N_2919);
or UO_380 (O_380,N_2778,N_2588);
xor UO_381 (O_381,N_2523,N_2555);
and UO_382 (O_382,N_2553,N_2508);
nand UO_383 (O_383,N_2880,N_2515);
or UO_384 (O_384,N_2760,N_2845);
nand UO_385 (O_385,N_2871,N_2867);
and UO_386 (O_386,N_2947,N_2781);
or UO_387 (O_387,N_2883,N_2939);
xnor UO_388 (O_388,N_2581,N_2846);
and UO_389 (O_389,N_2550,N_2650);
xor UO_390 (O_390,N_2599,N_2815);
and UO_391 (O_391,N_2576,N_2651);
nand UO_392 (O_392,N_2671,N_2976);
xor UO_393 (O_393,N_2656,N_2520);
nor UO_394 (O_394,N_2727,N_2720);
or UO_395 (O_395,N_2529,N_2825);
xnor UO_396 (O_396,N_2716,N_2961);
nand UO_397 (O_397,N_2960,N_2925);
xnor UO_398 (O_398,N_2970,N_2976);
nand UO_399 (O_399,N_2545,N_2993);
xor UO_400 (O_400,N_2841,N_2599);
or UO_401 (O_401,N_2601,N_2687);
nand UO_402 (O_402,N_2982,N_2718);
and UO_403 (O_403,N_2780,N_2880);
and UO_404 (O_404,N_2584,N_2953);
and UO_405 (O_405,N_2753,N_2873);
nand UO_406 (O_406,N_2834,N_2802);
nor UO_407 (O_407,N_2836,N_2862);
and UO_408 (O_408,N_2520,N_2657);
nand UO_409 (O_409,N_2704,N_2592);
and UO_410 (O_410,N_2970,N_2663);
nor UO_411 (O_411,N_2735,N_2951);
nand UO_412 (O_412,N_2990,N_2929);
or UO_413 (O_413,N_2676,N_2578);
or UO_414 (O_414,N_2922,N_2750);
or UO_415 (O_415,N_2564,N_2774);
nor UO_416 (O_416,N_2986,N_2996);
and UO_417 (O_417,N_2908,N_2651);
and UO_418 (O_418,N_2679,N_2590);
nand UO_419 (O_419,N_2665,N_2843);
or UO_420 (O_420,N_2787,N_2682);
xnor UO_421 (O_421,N_2936,N_2776);
or UO_422 (O_422,N_2531,N_2622);
nor UO_423 (O_423,N_2570,N_2657);
or UO_424 (O_424,N_2571,N_2850);
or UO_425 (O_425,N_2670,N_2817);
nand UO_426 (O_426,N_2504,N_2778);
or UO_427 (O_427,N_2663,N_2834);
and UO_428 (O_428,N_2856,N_2540);
nor UO_429 (O_429,N_2872,N_2635);
xnor UO_430 (O_430,N_2635,N_2775);
nor UO_431 (O_431,N_2592,N_2701);
and UO_432 (O_432,N_2715,N_2625);
and UO_433 (O_433,N_2852,N_2550);
or UO_434 (O_434,N_2674,N_2519);
and UO_435 (O_435,N_2870,N_2711);
xor UO_436 (O_436,N_2666,N_2930);
and UO_437 (O_437,N_2842,N_2582);
or UO_438 (O_438,N_2781,N_2614);
or UO_439 (O_439,N_2609,N_2654);
and UO_440 (O_440,N_2702,N_2567);
nor UO_441 (O_441,N_2593,N_2923);
nor UO_442 (O_442,N_2610,N_2762);
nor UO_443 (O_443,N_2898,N_2911);
nand UO_444 (O_444,N_2500,N_2975);
nand UO_445 (O_445,N_2642,N_2742);
nor UO_446 (O_446,N_2957,N_2782);
or UO_447 (O_447,N_2713,N_2753);
or UO_448 (O_448,N_2668,N_2987);
or UO_449 (O_449,N_2911,N_2528);
nand UO_450 (O_450,N_2631,N_2914);
and UO_451 (O_451,N_2539,N_2875);
or UO_452 (O_452,N_2904,N_2501);
or UO_453 (O_453,N_2692,N_2799);
or UO_454 (O_454,N_2611,N_2628);
xnor UO_455 (O_455,N_2589,N_2634);
xor UO_456 (O_456,N_2678,N_2554);
xnor UO_457 (O_457,N_2518,N_2678);
xnor UO_458 (O_458,N_2741,N_2857);
nor UO_459 (O_459,N_2649,N_2753);
or UO_460 (O_460,N_2518,N_2738);
xnor UO_461 (O_461,N_2923,N_2636);
nor UO_462 (O_462,N_2842,N_2841);
xnor UO_463 (O_463,N_2661,N_2623);
xor UO_464 (O_464,N_2524,N_2964);
nand UO_465 (O_465,N_2937,N_2840);
and UO_466 (O_466,N_2653,N_2712);
or UO_467 (O_467,N_2916,N_2799);
xor UO_468 (O_468,N_2851,N_2753);
nor UO_469 (O_469,N_2786,N_2772);
xor UO_470 (O_470,N_2860,N_2585);
nand UO_471 (O_471,N_2646,N_2849);
or UO_472 (O_472,N_2514,N_2864);
nor UO_473 (O_473,N_2854,N_2743);
nor UO_474 (O_474,N_2897,N_2767);
or UO_475 (O_475,N_2640,N_2991);
nand UO_476 (O_476,N_2906,N_2545);
xor UO_477 (O_477,N_2901,N_2962);
nand UO_478 (O_478,N_2845,N_2642);
nand UO_479 (O_479,N_2638,N_2873);
nand UO_480 (O_480,N_2856,N_2505);
xnor UO_481 (O_481,N_2636,N_2823);
nand UO_482 (O_482,N_2858,N_2794);
nand UO_483 (O_483,N_2939,N_2766);
nand UO_484 (O_484,N_2870,N_2888);
nor UO_485 (O_485,N_2721,N_2607);
xor UO_486 (O_486,N_2775,N_2731);
nor UO_487 (O_487,N_2544,N_2731);
nand UO_488 (O_488,N_2749,N_2505);
nand UO_489 (O_489,N_2813,N_2852);
or UO_490 (O_490,N_2538,N_2853);
nor UO_491 (O_491,N_2627,N_2805);
nor UO_492 (O_492,N_2859,N_2767);
and UO_493 (O_493,N_2586,N_2853);
nand UO_494 (O_494,N_2729,N_2631);
nor UO_495 (O_495,N_2899,N_2513);
nor UO_496 (O_496,N_2765,N_2938);
xor UO_497 (O_497,N_2631,N_2627);
xor UO_498 (O_498,N_2965,N_2539);
and UO_499 (O_499,N_2599,N_2770);
endmodule