module basic_500_3000_500_5_levels_1xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_154,In_207);
or U1 (N_1,In_283,In_230);
and U2 (N_2,In_61,In_18);
and U3 (N_3,In_82,In_340);
or U4 (N_4,In_29,In_9);
nor U5 (N_5,In_68,In_429);
or U6 (N_6,In_351,In_231);
or U7 (N_7,In_146,In_31);
and U8 (N_8,In_265,In_364);
or U9 (N_9,In_424,In_41);
nor U10 (N_10,In_363,In_456);
nor U11 (N_11,In_347,In_143);
nand U12 (N_12,In_305,In_357);
nand U13 (N_13,In_219,In_448);
nand U14 (N_14,In_324,In_235);
or U15 (N_15,In_76,In_38);
or U16 (N_16,In_260,In_455);
nand U17 (N_17,In_332,In_229);
and U18 (N_18,In_7,In_482);
or U19 (N_19,In_169,In_220);
nand U20 (N_20,In_433,In_385);
or U21 (N_21,In_126,In_3);
and U22 (N_22,In_187,In_97);
or U23 (N_23,In_227,In_107);
or U24 (N_24,In_270,In_390);
nand U25 (N_25,In_284,In_37);
or U26 (N_26,In_333,In_313);
or U27 (N_27,In_413,In_155);
and U28 (N_28,In_202,In_464);
nand U29 (N_29,In_262,In_228);
nor U30 (N_30,In_2,In_81);
nor U31 (N_31,In_257,In_392);
and U32 (N_32,In_271,In_497);
and U33 (N_33,In_254,In_291);
nor U34 (N_34,In_449,In_240);
nor U35 (N_35,In_58,In_200);
and U36 (N_36,In_495,In_386);
or U37 (N_37,In_21,In_216);
nand U38 (N_38,In_312,In_241);
nor U39 (N_39,In_277,In_408);
nor U40 (N_40,In_105,In_179);
nand U41 (N_41,In_272,In_173);
or U42 (N_42,In_388,In_276);
and U43 (N_43,In_17,In_188);
and U44 (N_44,In_310,In_157);
and U45 (N_45,In_63,In_415);
and U46 (N_46,In_70,In_314);
and U47 (N_47,In_86,In_181);
or U48 (N_48,In_339,In_439);
nor U49 (N_49,In_129,In_441);
nor U50 (N_50,In_204,In_25);
and U51 (N_51,In_160,In_472);
or U52 (N_52,In_474,In_62);
nor U53 (N_53,In_156,In_328);
or U54 (N_54,In_110,In_35);
nand U55 (N_55,In_373,In_432);
and U56 (N_56,In_483,In_402);
nor U57 (N_57,In_345,In_24);
or U58 (N_58,In_72,In_89);
nor U59 (N_59,In_434,In_123);
nand U60 (N_60,In_191,In_412);
nor U61 (N_61,In_486,In_327);
and U62 (N_62,In_114,In_201);
nand U63 (N_63,In_33,In_193);
or U64 (N_64,In_221,In_350);
nor U65 (N_65,In_478,In_22);
and U66 (N_66,In_67,In_421);
and U67 (N_67,In_95,In_263);
or U68 (N_68,In_279,In_69);
and U69 (N_69,In_379,In_302);
and U70 (N_70,In_316,In_300);
nand U71 (N_71,In_246,In_491);
and U72 (N_72,In_44,In_335);
nor U73 (N_73,In_459,In_295);
and U74 (N_74,In_376,In_12);
or U75 (N_75,In_147,In_223);
or U76 (N_76,In_1,In_59);
nor U77 (N_77,In_118,In_83);
nor U78 (N_78,In_419,In_293);
or U79 (N_79,In_286,In_494);
nand U80 (N_80,In_406,In_281);
nor U81 (N_81,In_39,In_233);
and U82 (N_82,In_131,In_132);
nand U83 (N_83,In_268,In_150);
and U84 (N_84,In_489,In_329);
nor U85 (N_85,In_488,In_396);
nor U86 (N_86,In_435,In_426);
and U87 (N_87,In_93,In_299);
nand U88 (N_88,In_322,In_389);
and U89 (N_89,In_30,In_440);
or U90 (N_90,In_369,In_487);
or U91 (N_91,In_91,In_102);
nor U92 (N_92,In_217,In_192);
and U93 (N_93,In_337,In_404);
nand U94 (N_94,In_346,In_292);
or U95 (N_95,In_323,In_248);
nand U96 (N_96,In_334,In_403);
or U97 (N_97,In_460,In_318);
and U98 (N_98,In_99,In_165);
nor U99 (N_99,In_422,In_480);
and U100 (N_100,In_280,In_282);
or U101 (N_101,In_238,In_0);
and U102 (N_102,In_236,In_414);
and U103 (N_103,In_8,In_368);
nor U104 (N_104,In_142,In_119);
and U105 (N_105,In_367,In_13);
or U106 (N_106,In_380,In_210);
nand U107 (N_107,In_384,In_101);
or U108 (N_108,In_109,In_247);
nand U109 (N_109,In_46,In_250);
or U110 (N_110,In_139,In_375);
and U111 (N_111,In_80,In_269);
and U112 (N_112,In_461,In_354);
nand U113 (N_113,In_261,In_103);
or U114 (N_114,In_196,In_43);
or U115 (N_115,In_203,In_251);
and U116 (N_116,In_387,In_409);
nand U117 (N_117,In_355,In_208);
nand U118 (N_118,In_471,In_467);
xor U119 (N_119,In_36,In_294);
and U120 (N_120,In_53,In_317);
and U121 (N_121,In_258,In_111);
and U122 (N_122,In_85,In_447);
nand U123 (N_123,In_431,In_135);
and U124 (N_124,In_397,In_49);
nand U125 (N_125,In_242,In_115);
nor U126 (N_126,In_430,In_226);
or U127 (N_127,In_57,In_395);
or U128 (N_128,In_326,In_436);
nor U129 (N_129,In_342,In_381);
and U130 (N_130,In_209,In_442);
and U131 (N_131,In_234,In_133);
and U132 (N_132,In_417,In_353);
nor U133 (N_133,In_453,In_4);
nor U134 (N_134,In_5,In_232);
nor U135 (N_135,In_125,In_56);
nor U136 (N_136,In_171,In_266);
nor U137 (N_137,In_359,In_370);
nand U138 (N_138,In_166,In_194);
or U139 (N_139,In_116,In_446);
nand U140 (N_140,In_152,In_399);
nand U141 (N_141,In_79,In_20);
and U142 (N_142,In_325,In_457);
nand U143 (N_143,In_176,In_259);
nand U144 (N_144,In_273,In_98);
xnor U145 (N_145,In_66,In_214);
nand U146 (N_146,In_71,In_55);
and U147 (N_147,In_361,In_290);
or U148 (N_148,In_34,In_26);
or U149 (N_149,In_438,In_470);
or U150 (N_150,In_215,In_104);
xor U151 (N_151,In_393,In_64);
nand U152 (N_152,In_149,In_23);
nor U153 (N_153,In_443,In_122);
and U154 (N_154,In_479,In_485);
or U155 (N_155,In_19,In_225);
and U156 (N_156,In_127,In_330);
nor U157 (N_157,In_65,In_428);
or U158 (N_158,In_42,In_183);
and U159 (N_159,In_121,In_498);
or U160 (N_160,In_47,In_163);
nand U161 (N_161,In_331,In_213);
or U162 (N_162,In_212,In_45);
and U163 (N_163,In_374,In_75);
and U164 (N_164,In_245,In_100);
or U165 (N_165,In_382,In_469);
and U166 (N_166,In_444,In_137);
and U167 (N_167,In_174,In_252);
and U168 (N_168,In_303,In_407);
nor U169 (N_169,In_378,In_128);
or U170 (N_170,In_50,In_400);
and U171 (N_171,In_141,In_159);
nand U172 (N_172,In_343,In_356);
and U173 (N_173,In_224,In_306);
and U174 (N_174,In_197,In_211);
or U175 (N_175,In_320,In_420);
or U176 (N_176,In_167,In_198);
or U177 (N_177,In_336,In_278);
or U178 (N_178,In_427,In_362);
nand U179 (N_179,In_140,In_6);
nor U180 (N_180,In_338,In_410);
nor U181 (N_181,In_452,In_73);
nand U182 (N_182,In_120,In_264);
nand U183 (N_183,In_170,In_78);
xnor U184 (N_184,In_398,In_138);
nor U185 (N_185,In_425,In_130);
nor U186 (N_186,In_124,In_383);
nand U187 (N_187,In_321,In_256);
nand U188 (N_188,In_274,In_285);
nor U189 (N_189,In_249,In_496);
nor U190 (N_190,In_177,In_161);
or U191 (N_191,In_365,In_11);
or U192 (N_192,In_401,In_451);
nand U193 (N_193,In_96,In_108);
nor U194 (N_194,In_366,In_90);
nor U195 (N_195,In_15,In_309);
nor U196 (N_196,In_40,In_344);
and U197 (N_197,In_311,In_186);
nand U198 (N_198,In_287,In_391);
nand U199 (N_199,In_32,In_136);
nand U200 (N_200,In_275,In_298);
nand U201 (N_201,In_463,In_190);
and U202 (N_202,In_168,In_199);
and U203 (N_203,In_466,In_189);
nand U204 (N_204,In_148,In_319);
nand U205 (N_205,In_54,In_493);
or U206 (N_206,In_255,In_106);
nor U207 (N_207,In_468,In_16);
and U208 (N_208,In_301,In_296);
nand U209 (N_209,In_492,In_243);
nor U210 (N_210,In_88,In_477);
and U211 (N_211,In_454,In_341);
nor U212 (N_212,In_352,In_92);
nand U213 (N_213,In_372,In_237);
nand U214 (N_214,In_172,In_308);
nand U215 (N_215,In_315,In_476);
nand U216 (N_216,In_411,In_117);
xor U217 (N_217,In_52,In_267);
nor U218 (N_218,In_462,In_112);
nor U219 (N_219,In_289,In_60);
and U220 (N_220,In_297,In_206);
nor U221 (N_221,In_244,In_158);
nand U222 (N_222,In_164,In_371);
nand U223 (N_223,In_84,In_222);
or U224 (N_224,In_304,In_445);
nand U225 (N_225,In_151,In_180);
and U226 (N_226,In_153,In_113);
or U227 (N_227,In_94,In_218);
or U228 (N_228,In_475,In_349);
or U229 (N_229,In_437,In_465);
nor U230 (N_230,In_28,In_162);
nand U231 (N_231,In_288,In_178);
nor U232 (N_232,In_184,In_27);
and U233 (N_233,In_394,In_195);
and U234 (N_234,In_253,In_144);
or U235 (N_235,In_481,In_348);
nand U236 (N_236,In_473,In_185);
nor U237 (N_237,In_405,In_450);
nand U238 (N_238,In_239,In_418);
and U239 (N_239,In_360,In_10);
nor U240 (N_240,In_48,In_307);
or U241 (N_241,In_74,In_423);
or U242 (N_242,In_484,In_358);
or U243 (N_243,In_77,In_175);
and U244 (N_244,In_205,In_87);
nand U245 (N_245,In_377,In_51);
nand U246 (N_246,In_416,In_490);
nor U247 (N_247,In_182,In_134);
or U248 (N_248,In_458,In_145);
nor U249 (N_249,In_14,In_499);
nor U250 (N_250,In_78,In_276);
nand U251 (N_251,In_475,In_263);
nor U252 (N_252,In_340,In_39);
nand U253 (N_253,In_94,In_347);
nor U254 (N_254,In_38,In_154);
nand U255 (N_255,In_181,In_264);
nand U256 (N_256,In_96,In_88);
nand U257 (N_257,In_49,In_135);
nand U258 (N_258,In_127,In_208);
nor U259 (N_259,In_184,In_146);
nor U260 (N_260,In_35,In_94);
and U261 (N_261,In_236,In_257);
nand U262 (N_262,In_411,In_420);
or U263 (N_263,In_292,In_149);
and U264 (N_264,In_86,In_445);
nand U265 (N_265,In_192,In_109);
and U266 (N_266,In_485,In_133);
and U267 (N_267,In_101,In_442);
and U268 (N_268,In_400,In_423);
or U269 (N_269,In_324,In_162);
and U270 (N_270,In_387,In_403);
nand U271 (N_271,In_417,In_308);
nor U272 (N_272,In_40,In_229);
nor U273 (N_273,In_413,In_438);
or U274 (N_274,In_200,In_470);
and U275 (N_275,In_143,In_148);
or U276 (N_276,In_373,In_9);
and U277 (N_277,In_135,In_134);
nor U278 (N_278,In_401,In_218);
or U279 (N_279,In_225,In_316);
nor U280 (N_280,In_493,In_449);
and U281 (N_281,In_140,In_295);
or U282 (N_282,In_184,In_33);
nand U283 (N_283,In_200,In_496);
nand U284 (N_284,In_330,In_462);
and U285 (N_285,In_481,In_120);
or U286 (N_286,In_384,In_452);
or U287 (N_287,In_129,In_69);
and U288 (N_288,In_257,In_457);
xor U289 (N_289,In_115,In_403);
nand U290 (N_290,In_421,In_373);
and U291 (N_291,In_191,In_462);
or U292 (N_292,In_60,In_348);
nor U293 (N_293,In_205,In_257);
and U294 (N_294,In_260,In_10);
nand U295 (N_295,In_262,In_203);
and U296 (N_296,In_488,In_175);
or U297 (N_297,In_28,In_158);
nand U298 (N_298,In_281,In_336);
and U299 (N_299,In_325,In_27);
nor U300 (N_300,In_115,In_404);
nor U301 (N_301,In_491,In_216);
nor U302 (N_302,In_112,In_108);
xnor U303 (N_303,In_281,In_215);
and U304 (N_304,In_442,In_57);
and U305 (N_305,In_372,In_105);
nor U306 (N_306,In_187,In_419);
and U307 (N_307,In_480,In_103);
nand U308 (N_308,In_267,In_129);
or U309 (N_309,In_254,In_133);
nor U310 (N_310,In_187,In_341);
and U311 (N_311,In_46,In_238);
or U312 (N_312,In_30,In_260);
and U313 (N_313,In_415,In_206);
and U314 (N_314,In_345,In_240);
nor U315 (N_315,In_175,In_378);
or U316 (N_316,In_100,In_365);
nor U317 (N_317,In_171,In_77);
nor U318 (N_318,In_44,In_154);
nand U319 (N_319,In_115,In_130);
nand U320 (N_320,In_416,In_161);
or U321 (N_321,In_183,In_129);
nor U322 (N_322,In_372,In_303);
nand U323 (N_323,In_182,In_200);
nor U324 (N_324,In_495,In_235);
or U325 (N_325,In_337,In_31);
and U326 (N_326,In_492,In_306);
nor U327 (N_327,In_32,In_11);
nor U328 (N_328,In_69,In_381);
or U329 (N_329,In_217,In_65);
or U330 (N_330,In_427,In_62);
or U331 (N_331,In_90,In_295);
nor U332 (N_332,In_114,In_179);
nand U333 (N_333,In_221,In_300);
nand U334 (N_334,In_433,In_282);
nand U335 (N_335,In_412,In_391);
or U336 (N_336,In_60,In_332);
or U337 (N_337,In_106,In_373);
and U338 (N_338,In_432,In_45);
or U339 (N_339,In_141,In_167);
and U340 (N_340,In_139,In_449);
nand U341 (N_341,In_216,In_371);
nand U342 (N_342,In_117,In_179);
or U343 (N_343,In_106,In_442);
nor U344 (N_344,In_335,In_328);
or U345 (N_345,In_200,In_138);
nor U346 (N_346,In_150,In_87);
and U347 (N_347,In_114,In_11);
nand U348 (N_348,In_375,In_98);
xor U349 (N_349,In_215,In_277);
or U350 (N_350,In_62,In_133);
and U351 (N_351,In_152,In_438);
nand U352 (N_352,In_402,In_155);
nand U353 (N_353,In_469,In_296);
and U354 (N_354,In_62,In_104);
nand U355 (N_355,In_415,In_248);
or U356 (N_356,In_183,In_134);
and U357 (N_357,In_204,In_74);
and U358 (N_358,In_108,In_240);
nand U359 (N_359,In_354,In_53);
nand U360 (N_360,In_189,In_251);
nand U361 (N_361,In_176,In_355);
nor U362 (N_362,In_210,In_331);
nor U363 (N_363,In_32,In_307);
and U364 (N_364,In_239,In_452);
and U365 (N_365,In_202,In_494);
nor U366 (N_366,In_258,In_282);
nand U367 (N_367,In_375,In_1);
nor U368 (N_368,In_84,In_493);
and U369 (N_369,In_190,In_280);
nor U370 (N_370,In_91,In_40);
nor U371 (N_371,In_81,In_96);
nor U372 (N_372,In_431,In_444);
or U373 (N_373,In_292,In_70);
nor U374 (N_374,In_428,In_293);
nand U375 (N_375,In_79,In_204);
nand U376 (N_376,In_292,In_301);
and U377 (N_377,In_331,In_189);
nand U378 (N_378,In_335,In_262);
xnor U379 (N_379,In_61,In_106);
and U380 (N_380,In_464,In_148);
nand U381 (N_381,In_128,In_213);
nor U382 (N_382,In_450,In_195);
and U383 (N_383,In_41,In_47);
nor U384 (N_384,In_18,In_268);
and U385 (N_385,In_132,In_241);
or U386 (N_386,In_199,In_227);
nor U387 (N_387,In_18,In_228);
nand U388 (N_388,In_392,In_353);
nand U389 (N_389,In_392,In_355);
and U390 (N_390,In_270,In_59);
or U391 (N_391,In_85,In_327);
nand U392 (N_392,In_102,In_187);
or U393 (N_393,In_316,In_322);
and U394 (N_394,In_393,In_412);
nand U395 (N_395,In_1,In_463);
nand U396 (N_396,In_264,In_495);
and U397 (N_397,In_206,In_408);
nor U398 (N_398,In_382,In_38);
and U399 (N_399,In_287,In_437);
or U400 (N_400,In_169,In_111);
and U401 (N_401,In_54,In_65);
nand U402 (N_402,In_293,In_281);
or U403 (N_403,In_166,In_13);
nand U404 (N_404,In_32,In_194);
nor U405 (N_405,In_191,In_456);
or U406 (N_406,In_59,In_333);
nor U407 (N_407,In_227,In_308);
nand U408 (N_408,In_200,In_485);
nor U409 (N_409,In_166,In_497);
nand U410 (N_410,In_126,In_453);
or U411 (N_411,In_125,In_264);
nor U412 (N_412,In_274,In_426);
or U413 (N_413,In_7,In_386);
or U414 (N_414,In_290,In_475);
and U415 (N_415,In_459,In_376);
nor U416 (N_416,In_314,In_12);
or U417 (N_417,In_139,In_133);
and U418 (N_418,In_122,In_86);
nor U419 (N_419,In_347,In_430);
nor U420 (N_420,In_437,In_316);
and U421 (N_421,In_319,In_273);
nor U422 (N_422,In_483,In_372);
or U423 (N_423,In_209,In_386);
and U424 (N_424,In_147,In_163);
nor U425 (N_425,In_495,In_314);
nor U426 (N_426,In_485,In_156);
or U427 (N_427,In_349,In_452);
or U428 (N_428,In_59,In_466);
xor U429 (N_429,In_220,In_19);
or U430 (N_430,In_360,In_190);
or U431 (N_431,In_220,In_435);
or U432 (N_432,In_69,In_123);
or U433 (N_433,In_405,In_495);
nor U434 (N_434,In_136,In_404);
nor U435 (N_435,In_484,In_63);
nor U436 (N_436,In_128,In_346);
nor U437 (N_437,In_244,In_59);
or U438 (N_438,In_463,In_489);
nand U439 (N_439,In_454,In_88);
and U440 (N_440,In_16,In_241);
nor U441 (N_441,In_1,In_94);
or U442 (N_442,In_275,In_161);
nand U443 (N_443,In_387,In_234);
or U444 (N_444,In_304,In_28);
or U445 (N_445,In_298,In_491);
nand U446 (N_446,In_228,In_321);
and U447 (N_447,In_273,In_390);
or U448 (N_448,In_426,In_407);
nor U449 (N_449,In_442,In_198);
nor U450 (N_450,In_225,In_426);
nand U451 (N_451,In_82,In_335);
or U452 (N_452,In_185,In_280);
nand U453 (N_453,In_209,In_387);
nand U454 (N_454,In_125,In_25);
nor U455 (N_455,In_372,In_215);
or U456 (N_456,In_165,In_263);
nand U457 (N_457,In_12,In_125);
or U458 (N_458,In_483,In_26);
or U459 (N_459,In_264,In_345);
and U460 (N_460,In_294,In_295);
nor U461 (N_461,In_19,In_45);
xnor U462 (N_462,In_6,In_273);
or U463 (N_463,In_166,In_368);
nor U464 (N_464,In_194,In_158);
and U465 (N_465,In_254,In_175);
and U466 (N_466,In_439,In_95);
xnor U467 (N_467,In_247,In_439);
or U468 (N_468,In_231,In_477);
and U469 (N_469,In_297,In_23);
nand U470 (N_470,In_278,In_338);
and U471 (N_471,In_292,In_86);
or U472 (N_472,In_483,In_422);
nor U473 (N_473,In_286,In_144);
nor U474 (N_474,In_87,In_353);
nor U475 (N_475,In_78,In_360);
nand U476 (N_476,In_202,In_71);
and U477 (N_477,In_193,In_172);
or U478 (N_478,In_312,In_276);
nor U479 (N_479,In_202,In_331);
or U480 (N_480,In_439,In_342);
nor U481 (N_481,In_268,In_121);
nor U482 (N_482,In_177,In_493);
and U483 (N_483,In_9,In_0);
or U484 (N_484,In_117,In_71);
or U485 (N_485,In_128,In_166);
nand U486 (N_486,In_410,In_411);
nand U487 (N_487,In_11,In_179);
or U488 (N_488,In_130,In_249);
or U489 (N_489,In_452,In_227);
nor U490 (N_490,In_97,In_55);
nor U491 (N_491,In_5,In_196);
nand U492 (N_492,In_76,In_276);
and U493 (N_493,In_46,In_312);
or U494 (N_494,In_26,In_99);
or U495 (N_495,In_206,In_220);
nor U496 (N_496,In_399,In_337);
or U497 (N_497,In_74,In_160);
or U498 (N_498,In_19,In_146);
xor U499 (N_499,In_52,In_219);
nand U500 (N_500,In_212,In_230);
and U501 (N_501,In_180,In_221);
or U502 (N_502,In_465,In_332);
or U503 (N_503,In_11,In_358);
or U504 (N_504,In_497,In_401);
and U505 (N_505,In_498,In_360);
nand U506 (N_506,In_371,In_66);
nor U507 (N_507,In_168,In_240);
nor U508 (N_508,In_5,In_303);
nor U509 (N_509,In_464,In_168);
nand U510 (N_510,In_378,In_124);
or U511 (N_511,In_389,In_379);
nand U512 (N_512,In_470,In_117);
nand U513 (N_513,In_394,In_317);
xnor U514 (N_514,In_242,In_7);
nor U515 (N_515,In_374,In_305);
nor U516 (N_516,In_458,In_348);
nor U517 (N_517,In_132,In_494);
and U518 (N_518,In_28,In_271);
nor U519 (N_519,In_236,In_302);
or U520 (N_520,In_255,In_180);
nand U521 (N_521,In_142,In_336);
or U522 (N_522,In_129,In_75);
nor U523 (N_523,In_335,In_270);
and U524 (N_524,In_138,In_238);
or U525 (N_525,In_169,In_245);
and U526 (N_526,In_163,In_220);
and U527 (N_527,In_86,In_359);
nor U528 (N_528,In_207,In_389);
nor U529 (N_529,In_149,In_466);
or U530 (N_530,In_145,In_91);
nand U531 (N_531,In_143,In_32);
or U532 (N_532,In_4,In_450);
nand U533 (N_533,In_337,In_298);
nand U534 (N_534,In_163,In_285);
nand U535 (N_535,In_290,In_484);
nand U536 (N_536,In_250,In_329);
nor U537 (N_537,In_321,In_8);
or U538 (N_538,In_488,In_446);
nand U539 (N_539,In_159,In_7);
nor U540 (N_540,In_372,In_264);
and U541 (N_541,In_145,In_57);
and U542 (N_542,In_395,In_269);
nor U543 (N_543,In_86,In_4);
nand U544 (N_544,In_477,In_484);
and U545 (N_545,In_326,In_366);
or U546 (N_546,In_228,In_106);
and U547 (N_547,In_457,In_306);
nand U548 (N_548,In_280,In_249);
or U549 (N_549,In_201,In_348);
and U550 (N_550,In_213,In_101);
and U551 (N_551,In_128,In_361);
nor U552 (N_552,In_202,In_378);
and U553 (N_553,In_32,In_485);
nor U554 (N_554,In_373,In_23);
or U555 (N_555,In_279,In_489);
or U556 (N_556,In_439,In_26);
nor U557 (N_557,In_359,In_136);
and U558 (N_558,In_278,In_311);
or U559 (N_559,In_68,In_219);
or U560 (N_560,In_202,In_430);
nand U561 (N_561,In_381,In_201);
and U562 (N_562,In_376,In_108);
or U563 (N_563,In_206,In_161);
nand U564 (N_564,In_56,In_5);
nand U565 (N_565,In_348,In_98);
and U566 (N_566,In_195,In_417);
nand U567 (N_567,In_443,In_175);
nor U568 (N_568,In_423,In_494);
and U569 (N_569,In_371,In_410);
or U570 (N_570,In_295,In_419);
and U571 (N_571,In_257,In_228);
nor U572 (N_572,In_357,In_203);
and U573 (N_573,In_18,In_120);
nor U574 (N_574,In_139,In_3);
and U575 (N_575,In_104,In_111);
nand U576 (N_576,In_217,In_205);
nand U577 (N_577,In_346,In_360);
nor U578 (N_578,In_31,In_95);
or U579 (N_579,In_72,In_3);
nor U580 (N_580,In_374,In_295);
or U581 (N_581,In_163,In_269);
nor U582 (N_582,In_237,In_300);
nor U583 (N_583,In_418,In_421);
or U584 (N_584,In_358,In_380);
or U585 (N_585,In_226,In_29);
nand U586 (N_586,In_388,In_329);
or U587 (N_587,In_483,In_400);
and U588 (N_588,In_230,In_191);
or U589 (N_589,In_239,In_408);
nor U590 (N_590,In_229,In_282);
and U591 (N_591,In_468,In_420);
nor U592 (N_592,In_229,In_118);
nor U593 (N_593,In_482,In_190);
nor U594 (N_594,In_184,In_88);
nand U595 (N_595,In_255,In_492);
nand U596 (N_596,In_489,In_415);
nor U597 (N_597,In_369,In_232);
or U598 (N_598,In_208,In_41);
nor U599 (N_599,In_105,In_199);
and U600 (N_600,N_510,N_166);
or U601 (N_601,N_263,N_556);
xnor U602 (N_602,N_597,N_137);
or U603 (N_603,N_204,N_460);
and U604 (N_604,N_524,N_282);
nand U605 (N_605,N_598,N_242);
nand U606 (N_606,N_373,N_341);
and U607 (N_607,N_56,N_287);
and U608 (N_608,N_225,N_291);
xnor U609 (N_609,N_335,N_69);
and U610 (N_610,N_60,N_207);
nand U611 (N_611,N_477,N_299);
nand U612 (N_612,N_508,N_509);
and U613 (N_613,N_439,N_237);
or U614 (N_614,N_275,N_231);
nor U615 (N_615,N_549,N_127);
or U616 (N_616,N_221,N_454);
nor U617 (N_617,N_300,N_90);
nor U618 (N_618,N_314,N_548);
nand U619 (N_619,N_243,N_408);
or U620 (N_620,N_72,N_61);
nand U621 (N_621,N_293,N_353);
or U622 (N_622,N_47,N_591);
or U623 (N_623,N_20,N_119);
or U624 (N_624,N_414,N_134);
or U625 (N_625,N_308,N_145);
or U626 (N_626,N_585,N_226);
nor U627 (N_627,N_148,N_389);
and U628 (N_628,N_379,N_109);
nand U629 (N_629,N_248,N_192);
or U630 (N_630,N_499,N_284);
nand U631 (N_631,N_165,N_64);
or U632 (N_632,N_254,N_594);
or U633 (N_633,N_513,N_334);
and U634 (N_634,N_575,N_582);
or U635 (N_635,N_0,N_512);
nor U636 (N_636,N_362,N_95);
nor U637 (N_637,N_465,N_62);
and U638 (N_638,N_208,N_235);
xnor U639 (N_639,N_444,N_289);
and U640 (N_640,N_484,N_23);
or U641 (N_641,N_218,N_211);
or U642 (N_642,N_177,N_401);
and U643 (N_643,N_160,N_34);
nor U644 (N_644,N_312,N_365);
or U645 (N_645,N_330,N_132);
or U646 (N_646,N_419,N_281);
or U647 (N_647,N_9,N_453);
and U648 (N_648,N_294,N_249);
or U649 (N_649,N_112,N_1);
nand U650 (N_650,N_339,N_506);
nand U651 (N_651,N_313,N_345);
or U652 (N_652,N_178,N_50);
or U653 (N_653,N_283,N_121);
nand U654 (N_654,N_104,N_153);
nor U655 (N_655,N_187,N_11);
or U656 (N_656,N_396,N_21);
nor U657 (N_657,N_496,N_167);
and U658 (N_658,N_435,N_410);
nand U659 (N_659,N_361,N_318);
or U660 (N_660,N_52,N_151);
and U661 (N_661,N_196,N_459);
xnor U662 (N_662,N_443,N_413);
and U663 (N_663,N_333,N_271);
xnor U664 (N_664,N_246,N_307);
or U665 (N_665,N_245,N_98);
or U666 (N_666,N_257,N_468);
or U667 (N_667,N_189,N_403);
nand U668 (N_668,N_467,N_126);
or U669 (N_669,N_523,N_532);
nor U670 (N_670,N_309,N_324);
or U671 (N_671,N_431,N_206);
or U672 (N_672,N_327,N_570);
nand U673 (N_673,N_28,N_219);
and U674 (N_674,N_531,N_550);
xor U675 (N_675,N_40,N_3);
nand U676 (N_676,N_150,N_27);
nor U677 (N_677,N_65,N_86);
and U678 (N_678,N_240,N_123);
and U679 (N_679,N_344,N_168);
and U680 (N_680,N_7,N_436);
and U681 (N_681,N_441,N_547);
or U682 (N_682,N_393,N_424);
or U683 (N_683,N_392,N_210);
nand U684 (N_684,N_409,N_212);
nand U685 (N_685,N_171,N_337);
or U686 (N_686,N_162,N_110);
nand U687 (N_687,N_558,N_175);
and U688 (N_688,N_437,N_446);
nor U689 (N_689,N_486,N_473);
nor U690 (N_690,N_449,N_423);
nand U691 (N_691,N_458,N_233);
nand U692 (N_692,N_286,N_131);
and U693 (N_693,N_82,N_536);
and U694 (N_694,N_336,N_452);
nor U695 (N_695,N_525,N_39);
or U696 (N_696,N_228,N_426);
nand U697 (N_697,N_35,N_319);
and U698 (N_698,N_561,N_43);
nor U699 (N_699,N_588,N_227);
nor U700 (N_700,N_518,N_348);
or U701 (N_701,N_391,N_93);
and U702 (N_702,N_377,N_76);
nor U703 (N_703,N_285,N_37);
nand U704 (N_704,N_495,N_77);
nor U705 (N_705,N_343,N_573);
nand U706 (N_706,N_315,N_417);
or U707 (N_707,N_464,N_522);
nand U708 (N_708,N_328,N_280);
nand U709 (N_709,N_136,N_567);
nor U710 (N_710,N_310,N_476);
nand U711 (N_711,N_164,N_253);
nor U712 (N_712,N_38,N_277);
nor U713 (N_713,N_388,N_407);
nand U714 (N_714,N_36,N_321);
nor U715 (N_715,N_596,N_295);
nor U716 (N_716,N_492,N_478);
and U717 (N_717,N_350,N_138);
nand U718 (N_718,N_128,N_360);
nand U719 (N_719,N_519,N_516);
or U720 (N_720,N_250,N_583);
or U721 (N_721,N_102,N_63);
nand U722 (N_722,N_576,N_256);
nor U723 (N_723,N_180,N_397);
and U724 (N_724,N_264,N_412);
and U725 (N_725,N_186,N_179);
nand U726 (N_726,N_113,N_357);
nand U727 (N_727,N_170,N_51);
nand U728 (N_728,N_526,N_197);
nor U729 (N_729,N_562,N_381);
nand U730 (N_730,N_529,N_411);
nand U731 (N_731,N_566,N_191);
or U732 (N_732,N_45,N_267);
or U733 (N_733,N_149,N_405);
nand U734 (N_734,N_528,N_111);
nor U735 (N_735,N_258,N_58);
and U736 (N_736,N_470,N_74);
nor U737 (N_737,N_555,N_442);
nand U738 (N_738,N_84,N_209);
and U739 (N_739,N_400,N_83);
or U740 (N_740,N_428,N_322);
nand U741 (N_741,N_195,N_354);
or U742 (N_742,N_406,N_457);
nand U743 (N_743,N_367,N_346);
and U744 (N_744,N_143,N_376);
nand U745 (N_745,N_122,N_87);
nand U746 (N_746,N_41,N_317);
nor U747 (N_747,N_92,N_586);
or U748 (N_748,N_542,N_97);
or U749 (N_749,N_469,N_323);
or U750 (N_750,N_366,N_572);
nor U751 (N_751,N_497,N_13);
nor U752 (N_752,N_269,N_584);
nor U753 (N_753,N_6,N_296);
nor U754 (N_754,N_265,N_577);
nand U755 (N_755,N_370,N_22);
nor U756 (N_756,N_565,N_91);
and U757 (N_757,N_368,N_68);
or U758 (N_758,N_130,N_432);
nor U759 (N_759,N_182,N_599);
or U760 (N_760,N_504,N_456);
or U761 (N_761,N_181,N_185);
or U762 (N_762,N_463,N_232);
and U763 (N_763,N_216,N_12);
nor U764 (N_764,N_455,N_450);
or U765 (N_765,N_503,N_199);
or U766 (N_766,N_57,N_502);
and U767 (N_767,N_445,N_255);
nor U768 (N_768,N_223,N_487);
and U769 (N_769,N_416,N_96);
and U770 (N_770,N_16,N_188);
and U771 (N_771,N_500,N_303);
and U772 (N_772,N_351,N_18);
nand U773 (N_773,N_349,N_215);
nor U774 (N_774,N_129,N_114);
nand U775 (N_775,N_142,N_4);
nand U776 (N_776,N_118,N_480);
and U777 (N_777,N_268,N_539);
nand U778 (N_778,N_404,N_479);
and U779 (N_779,N_371,N_147);
nand U780 (N_780,N_107,N_169);
or U781 (N_781,N_290,N_135);
nand U782 (N_782,N_387,N_320);
and U783 (N_783,N_311,N_244);
nor U784 (N_784,N_8,N_238);
nand U785 (N_785,N_203,N_152);
nor U786 (N_786,N_262,N_194);
and U787 (N_787,N_106,N_5);
nand U788 (N_788,N_386,N_305);
nand U789 (N_789,N_176,N_578);
nor U790 (N_790,N_260,N_448);
and U791 (N_791,N_491,N_358);
nand U792 (N_792,N_494,N_521);
nand U793 (N_793,N_85,N_474);
nand U794 (N_794,N_217,N_274);
and U795 (N_795,N_580,N_54);
nor U796 (N_796,N_251,N_272);
and U797 (N_797,N_259,N_292);
or U798 (N_798,N_438,N_372);
nor U799 (N_799,N_155,N_571);
or U800 (N_800,N_141,N_306);
nor U801 (N_801,N_482,N_421);
and U802 (N_802,N_230,N_301);
or U803 (N_803,N_198,N_190);
nor U804 (N_804,N_116,N_515);
nor U805 (N_805,N_342,N_139);
nand U806 (N_806,N_507,N_46);
and U807 (N_807,N_587,N_325);
and U808 (N_808,N_384,N_73);
and U809 (N_809,N_471,N_78);
nor U810 (N_810,N_159,N_278);
nand U811 (N_811,N_17,N_234);
or U812 (N_812,N_184,N_67);
and U813 (N_813,N_541,N_273);
xnor U814 (N_814,N_19,N_581);
xnor U815 (N_815,N_538,N_356);
and U816 (N_816,N_363,N_557);
or U817 (N_817,N_589,N_553);
nor U818 (N_818,N_53,N_425);
and U819 (N_819,N_537,N_288);
and U820 (N_820,N_560,N_544);
and U821 (N_821,N_239,N_229);
or U822 (N_822,N_462,N_201);
nor U823 (N_823,N_574,N_472);
or U824 (N_824,N_563,N_214);
nor U825 (N_825,N_385,N_200);
nor U826 (N_826,N_202,N_174);
and U827 (N_827,N_355,N_340);
or U828 (N_828,N_304,N_375);
and U829 (N_829,N_434,N_42);
nor U830 (N_830,N_220,N_501);
or U831 (N_831,N_552,N_48);
nand U832 (N_832,N_402,N_533);
nand U833 (N_833,N_489,N_390);
or U834 (N_834,N_579,N_103);
or U835 (N_835,N_88,N_125);
and U836 (N_836,N_44,N_205);
or U837 (N_837,N_415,N_24);
nor U838 (N_838,N_158,N_475);
and U839 (N_839,N_514,N_483);
nor U840 (N_840,N_568,N_451);
or U841 (N_841,N_173,N_593);
nand U842 (N_842,N_261,N_422);
nand U843 (N_843,N_157,N_352);
or U844 (N_844,N_29,N_543);
nor U845 (N_845,N_347,N_163);
nor U846 (N_846,N_156,N_331);
nand U847 (N_847,N_124,N_546);
nand U848 (N_848,N_493,N_332);
nand U849 (N_849,N_590,N_535);
nand U850 (N_850,N_420,N_276);
nand U851 (N_851,N_183,N_55);
nor U852 (N_852,N_2,N_418);
nand U853 (N_853,N_302,N_15);
or U854 (N_854,N_146,N_33);
and U855 (N_855,N_485,N_133);
or U856 (N_856,N_359,N_447);
or U857 (N_857,N_490,N_383);
nor U858 (N_858,N_117,N_193);
or U859 (N_859,N_247,N_338);
nand U860 (N_860,N_236,N_105);
or U861 (N_861,N_75,N_461);
or U862 (N_862,N_140,N_364);
nor U863 (N_863,N_569,N_564);
and U864 (N_864,N_380,N_270);
nor U865 (N_865,N_25,N_241);
nand U866 (N_866,N_14,N_530);
and U867 (N_867,N_595,N_433);
nor U868 (N_868,N_224,N_329);
nor U869 (N_869,N_498,N_81);
nand U870 (N_870,N_279,N_213);
or U871 (N_871,N_59,N_79);
and U872 (N_872,N_66,N_298);
nand U873 (N_873,N_488,N_551);
or U874 (N_874,N_89,N_554);
and U875 (N_875,N_481,N_430);
and U876 (N_876,N_100,N_222);
and U877 (N_877,N_505,N_517);
and U878 (N_878,N_71,N_26);
and U879 (N_879,N_399,N_10);
and U880 (N_880,N_520,N_378);
and U881 (N_881,N_120,N_94);
nor U882 (N_882,N_369,N_511);
nand U883 (N_883,N_427,N_154);
and U884 (N_884,N_440,N_161);
nor U885 (N_885,N_429,N_101);
or U886 (N_886,N_32,N_30);
nand U887 (N_887,N_398,N_592);
nor U888 (N_888,N_99,N_540);
or U889 (N_889,N_316,N_70);
nand U890 (N_890,N_297,N_394);
nor U891 (N_891,N_108,N_252);
nand U892 (N_892,N_466,N_31);
and U893 (N_893,N_395,N_80);
nor U894 (N_894,N_559,N_374);
nand U895 (N_895,N_144,N_534);
and U896 (N_896,N_115,N_527);
or U897 (N_897,N_326,N_266);
nor U898 (N_898,N_49,N_382);
and U899 (N_899,N_545,N_172);
nor U900 (N_900,N_162,N_216);
or U901 (N_901,N_449,N_18);
nor U902 (N_902,N_329,N_355);
nand U903 (N_903,N_258,N_207);
and U904 (N_904,N_450,N_284);
nor U905 (N_905,N_369,N_565);
and U906 (N_906,N_32,N_442);
nand U907 (N_907,N_193,N_90);
nor U908 (N_908,N_469,N_372);
or U909 (N_909,N_410,N_180);
and U910 (N_910,N_2,N_109);
nor U911 (N_911,N_560,N_190);
nand U912 (N_912,N_185,N_438);
or U913 (N_913,N_328,N_289);
nor U914 (N_914,N_379,N_186);
and U915 (N_915,N_173,N_334);
nand U916 (N_916,N_463,N_26);
nand U917 (N_917,N_387,N_365);
or U918 (N_918,N_424,N_122);
or U919 (N_919,N_86,N_117);
nor U920 (N_920,N_216,N_572);
or U921 (N_921,N_586,N_140);
nor U922 (N_922,N_17,N_357);
nor U923 (N_923,N_175,N_387);
nand U924 (N_924,N_12,N_140);
nand U925 (N_925,N_4,N_371);
and U926 (N_926,N_551,N_422);
and U927 (N_927,N_107,N_51);
and U928 (N_928,N_218,N_111);
nor U929 (N_929,N_412,N_53);
nor U930 (N_930,N_350,N_590);
nor U931 (N_931,N_547,N_533);
and U932 (N_932,N_79,N_118);
nor U933 (N_933,N_228,N_402);
nor U934 (N_934,N_70,N_84);
and U935 (N_935,N_192,N_364);
or U936 (N_936,N_460,N_577);
nor U937 (N_937,N_522,N_214);
and U938 (N_938,N_372,N_21);
nor U939 (N_939,N_40,N_326);
or U940 (N_940,N_551,N_260);
or U941 (N_941,N_393,N_354);
nor U942 (N_942,N_46,N_76);
or U943 (N_943,N_421,N_549);
or U944 (N_944,N_461,N_568);
and U945 (N_945,N_265,N_160);
nor U946 (N_946,N_79,N_278);
nor U947 (N_947,N_211,N_13);
or U948 (N_948,N_133,N_548);
nor U949 (N_949,N_476,N_488);
nand U950 (N_950,N_301,N_17);
and U951 (N_951,N_376,N_341);
nand U952 (N_952,N_516,N_328);
xnor U953 (N_953,N_496,N_230);
or U954 (N_954,N_25,N_572);
and U955 (N_955,N_86,N_155);
and U956 (N_956,N_292,N_251);
nand U957 (N_957,N_507,N_101);
nand U958 (N_958,N_395,N_467);
nor U959 (N_959,N_365,N_543);
nor U960 (N_960,N_139,N_185);
or U961 (N_961,N_506,N_349);
nand U962 (N_962,N_22,N_347);
nor U963 (N_963,N_260,N_354);
and U964 (N_964,N_470,N_26);
nand U965 (N_965,N_245,N_512);
nand U966 (N_966,N_480,N_135);
nor U967 (N_967,N_294,N_87);
nor U968 (N_968,N_324,N_243);
and U969 (N_969,N_187,N_112);
nor U970 (N_970,N_190,N_338);
nor U971 (N_971,N_377,N_444);
and U972 (N_972,N_108,N_380);
nor U973 (N_973,N_215,N_242);
nand U974 (N_974,N_260,N_117);
nor U975 (N_975,N_448,N_117);
nor U976 (N_976,N_402,N_152);
nand U977 (N_977,N_361,N_197);
or U978 (N_978,N_439,N_387);
and U979 (N_979,N_271,N_141);
or U980 (N_980,N_542,N_497);
and U981 (N_981,N_189,N_64);
nor U982 (N_982,N_322,N_378);
nand U983 (N_983,N_376,N_322);
nand U984 (N_984,N_134,N_213);
nor U985 (N_985,N_341,N_124);
or U986 (N_986,N_338,N_241);
and U987 (N_987,N_399,N_107);
nand U988 (N_988,N_244,N_364);
or U989 (N_989,N_440,N_57);
nand U990 (N_990,N_316,N_246);
nand U991 (N_991,N_29,N_469);
or U992 (N_992,N_463,N_597);
nand U993 (N_993,N_199,N_583);
nand U994 (N_994,N_572,N_329);
or U995 (N_995,N_286,N_15);
or U996 (N_996,N_384,N_528);
nand U997 (N_997,N_499,N_386);
nand U998 (N_998,N_54,N_80);
nor U999 (N_999,N_458,N_50);
nand U1000 (N_1000,N_93,N_54);
nand U1001 (N_1001,N_360,N_408);
nand U1002 (N_1002,N_470,N_436);
nand U1003 (N_1003,N_535,N_228);
and U1004 (N_1004,N_196,N_56);
nor U1005 (N_1005,N_44,N_589);
or U1006 (N_1006,N_435,N_204);
nor U1007 (N_1007,N_370,N_528);
nand U1008 (N_1008,N_449,N_321);
nand U1009 (N_1009,N_257,N_574);
and U1010 (N_1010,N_27,N_43);
nand U1011 (N_1011,N_438,N_558);
nor U1012 (N_1012,N_319,N_373);
nor U1013 (N_1013,N_45,N_88);
or U1014 (N_1014,N_117,N_325);
nand U1015 (N_1015,N_486,N_414);
and U1016 (N_1016,N_128,N_40);
nor U1017 (N_1017,N_563,N_432);
nor U1018 (N_1018,N_27,N_100);
nand U1019 (N_1019,N_65,N_243);
and U1020 (N_1020,N_239,N_167);
or U1021 (N_1021,N_491,N_312);
and U1022 (N_1022,N_184,N_375);
and U1023 (N_1023,N_568,N_491);
nand U1024 (N_1024,N_93,N_247);
nor U1025 (N_1025,N_358,N_199);
and U1026 (N_1026,N_450,N_579);
and U1027 (N_1027,N_144,N_234);
and U1028 (N_1028,N_574,N_268);
nand U1029 (N_1029,N_11,N_486);
or U1030 (N_1030,N_174,N_143);
nand U1031 (N_1031,N_263,N_418);
nand U1032 (N_1032,N_262,N_448);
nor U1033 (N_1033,N_153,N_295);
nor U1034 (N_1034,N_41,N_480);
and U1035 (N_1035,N_41,N_138);
and U1036 (N_1036,N_531,N_167);
nor U1037 (N_1037,N_68,N_443);
nand U1038 (N_1038,N_507,N_77);
and U1039 (N_1039,N_228,N_392);
nor U1040 (N_1040,N_320,N_214);
nand U1041 (N_1041,N_584,N_404);
and U1042 (N_1042,N_4,N_271);
nand U1043 (N_1043,N_372,N_163);
and U1044 (N_1044,N_94,N_356);
or U1045 (N_1045,N_221,N_520);
nor U1046 (N_1046,N_195,N_591);
nor U1047 (N_1047,N_73,N_174);
nor U1048 (N_1048,N_552,N_491);
and U1049 (N_1049,N_22,N_291);
nand U1050 (N_1050,N_433,N_237);
nand U1051 (N_1051,N_264,N_209);
nand U1052 (N_1052,N_9,N_25);
nor U1053 (N_1053,N_436,N_583);
and U1054 (N_1054,N_518,N_168);
and U1055 (N_1055,N_41,N_248);
nand U1056 (N_1056,N_275,N_284);
nand U1057 (N_1057,N_404,N_451);
nand U1058 (N_1058,N_116,N_110);
nand U1059 (N_1059,N_194,N_443);
or U1060 (N_1060,N_152,N_220);
or U1061 (N_1061,N_8,N_35);
or U1062 (N_1062,N_476,N_299);
or U1063 (N_1063,N_42,N_559);
and U1064 (N_1064,N_470,N_395);
and U1065 (N_1065,N_495,N_289);
nand U1066 (N_1066,N_457,N_416);
and U1067 (N_1067,N_487,N_562);
nand U1068 (N_1068,N_537,N_500);
nor U1069 (N_1069,N_492,N_494);
nor U1070 (N_1070,N_117,N_276);
nor U1071 (N_1071,N_403,N_493);
or U1072 (N_1072,N_105,N_172);
nand U1073 (N_1073,N_100,N_57);
or U1074 (N_1074,N_543,N_301);
nand U1075 (N_1075,N_202,N_383);
or U1076 (N_1076,N_143,N_200);
or U1077 (N_1077,N_30,N_535);
nand U1078 (N_1078,N_52,N_284);
xnor U1079 (N_1079,N_551,N_511);
or U1080 (N_1080,N_334,N_401);
or U1081 (N_1081,N_493,N_256);
nor U1082 (N_1082,N_358,N_108);
nand U1083 (N_1083,N_21,N_476);
nand U1084 (N_1084,N_541,N_230);
nor U1085 (N_1085,N_523,N_544);
and U1086 (N_1086,N_380,N_293);
or U1087 (N_1087,N_530,N_231);
nor U1088 (N_1088,N_290,N_151);
nor U1089 (N_1089,N_474,N_234);
nor U1090 (N_1090,N_451,N_75);
nor U1091 (N_1091,N_121,N_330);
or U1092 (N_1092,N_206,N_102);
nor U1093 (N_1093,N_523,N_111);
or U1094 (N_1094,N_158,N_453);
and U1095 (N_1095,N_391,N_478);
nand U1096 (N_1096,N_361,N_186);
or U1097 (N_1097,N_303,N_474);
and U1098 (N_1098,N_207,N_251);
and U1099 (N_1099,N_239,N_135);
nor U1100 (N_1100,N_35,N_272);
nor U1101 (N_1101,N_257,N_170);
nand U1102 (N_1102,N_519,N_344);
nand U1103 (N_1103,N_77,N_188);
and U1104 (N_1104,N_452,N_481);
nand U1105 (N_1105,N_402,N_366);
nand U1106 (N_1106,N_165,N_271);
nor U1107 (N_1107,N_60,N_90);
nand U1108 (N_1108,N_187,N_107);
and U1109 (N_1109,N_487,N_440);
or U1110 (N_1110,N_156,N_35);
and U1111 (N_1111,N_50,N_333);
or U1112 (N_1112,N_134,N_401);
nand U1113 (N_1113,N_412,N_246);
nand U1114 (N_1114,N_182,N_300);
nand U1115 (N_1115,N_404,N_286);
nor U1116 (N_1116,N_269,N_380);
and U1117 (N_1117,N_6,N_572);
nor U1118 (N_1118,N_469,N_105);
nand U1119 (N_1119,N_120,N_382);
and U1120 (N_1120,N_89,N_81);
nor U1121 (N_1121,N_417,N_100);
and U1122 (N_1122,N_524,N_2);
nand U1123 (N_1123,N_382,N_542);
and U1124 (N_1124,N_512,N_32);
nor U1125 (N_1125,N_545,N_207);
nand U1126 (N_1126,N_571,N_198);
nand U1127 (N_1127,N_407,N_286);
and U1128 (N_1128,N_519,N_456);
or U1129 (N_1129,N_594,N_491);
nor U1130 (N_1130,N_362,N_406);
nor U1131 (N_1131,N_372,N_428);
nand U1132 (N_1132,N_217,N_322);
nor U1133 (N_1133,N_358,N_322);
nand U1134 (N_1134,N_432,N_75);
and U1135 (N_1135,N_477,N_428);
or U1136 (N_1136,N_348,N_203);
nand U1137 (N_1137,N_328,N_100);
or U1138 (N_1138,N_297,N_594);
nor U1139 (N_1139,N_284,N_30);
and U1140 (N_1140,N_420,N_271);
xnor U1141 (N_1141,N_502,N_158);
or U1142 (N_1142,N_154,N_389);
nand U1143 (N_1143,N_136,N_95);
or U1144 (N_1144,N_147,N_9);
nand U1145 (N_1145,N_414,N_89);
nor U1146 (N_1146,N_522,N_255);
or U1147 (N_1147,N_65,N_339);
xnor U1148 (N_1148,N_38,N_526);
and U1149 (N_1149,N_150,N_180);
or U1150 (N_1150,N_125,N_298);
and U1151 (N_1151,N_412,N_284);
nand U1152 (N_1152,N_108,N_221);
and U1153 (N_1153,N_311,N_567);
or U1154 (N_1154,N_228,N_206);
nand U1155 (N_1155,N_231,N_10);
nor U1156 (N_1156,N_175,N_538);
or U1157 (N_1157,N_332,N_513);
nor U1158 (N_1158,N_429,N_248);
and U1159 (N_1159,N_198,N_109);
and U1160 (N_1160,N_279,N_115);
or U1161 (N_1161,N_263,N_444);
nor U1162 (N_1162,N_143,N_47);
nor U1163 (N_1163,N_263,N_431);
or U1164 (N_1164,N_589,N_404);
or U1165 (N_1165,N_526,N_372);
and U1166 (N_1166,N_162,N_176);
nor U1167 (N_1167,N_389,N_598);
nand U1168 (N_1168,N_313,N_321);
or U1169 (N_1169,N_123,N_563);
or U1170 (N_1170,N_453,N_216);
nor U1171 (N_1171,N_385,N_279);
nand U1172 (N_1172,N_349,N_569);
nor U1173 (N_1173,N_219,N_192);
nor U1174 (N_1174,N_36,N_598);
or U1175 (N_1175,N_186,N_203);
or U1176 (N_1176,N_250,N_529);
and U1177 (N_1177,N_465,N_430);
nand U1178 (N_1178,N_387,N_53);
nand U1179 (N_1179,N_481,N_489);
and U1180 (N_1180,N_40,N_247);
and U1181 (N_1181,N_573,N_264);
and U1182 (N_1182,N_338,N_124);
or U1183 (N_1183,N_247,N_486);
or U1184 (N_1184,N_354,N_374);
or U1185 (N_1185,N_327,N_49);
and U1186 (N_1186,N_43,N_479);
nor U1187 (N_1187,N_380,N_285);
or U1188 (N_1188,N_313,N_589);
and U1189 (N_1189,N_536,N_585);
and U1190 (N_1190,N_13,N_500);
or U1191 (N_1191,N_449,N_497);
nand U1192 (N_1192,N_186,N_426);
nand U1193 (N_1193,N_42,N_250);
nor U1194 (N_1194,N_1,N_574);
nor U1195 (N_1195,N_292,N_149);
or U1196 (N_1196,N_571,N_132);
nand U1197 (N_1197,N_1,N_387);
and U1198 (N_1198,N_211,N_174);
and U1199 (N_1199,N_328,N_365);
and U1200 (N_1200,N_635,N_613);
nor U1201 (N_1201,N_1012,N_1038);
nand U1202 (N_1202,N_937,N_1010);
or U1203 (N_1203,N_1145,N_944);
nor U1204 (N_1204,N_802,N_1146);
nor U1205 (N_1205,N_1026,N_1082);
nand U1206 (N_1206,N_861,N_789);
or U1207 (N_1207,N_706,N_822);
nand U1208 (N_1208,N_946,N_963);
and U1209 (N_1209,N_731,N_759);
nor U1210 (N_1210,N_1060,N_1075);
and U1211 (N_1211,N_1053,N_719);
nand U1212 (N_1212,N_1137,N_602);
nor U1213 (N_1213,N_751,N_1159);
or U1214 (N_1214,N_1059,N_661);
nor U1215 (N_1215,N_859,N_903);
or U1216 (N_1216,N_630,N_1179);
or U1217 (N_1217,N_942,N_729);
nor U1218 (N_1218,N_806,N_987);
nor U1219 (N_1219,N_614,N_703);
nor U1220 (N_1220,N_1002,N_670);
and U1221 (N_1221,N_1017,N_619);
nand U1222 (N_1222,N_1167,N_1153);
or U1223 (N_1223,N_960,N_989);
nand U1224 (N_1224,N_967,N_1125);
or U1225 (N_1225,N_1093,N_810);
or U1226 (N_1226,N_880,N_608);
or U1227 (N_1227,N_625,N_780);
and U1228 (N_1228,N_1191,N_823);
nor U1229 (N_1229,N_951,N_632);
and U1230 (N_1230,N_1165,N_844);
nor U1231 (N_1231,N_919,N_607);
nor U1232 (N_1232,N_1094,N_674);
or U1233 (N_1233,N_1158,N_935);
nand U1234 (N_1234,N_1003,N_1031);
nor U1235 (N_1235,N_1047,N_933);
nand U1236 (N_1236,N_883,N_926);
and U1237 (N_1237,N_768,N_742);
or U1238 (N_1238,N_882,N_1154);
nor U1239 (N_1239,N_1149,N_988);
and U1240 (N_1240,N_626,N_1120);
nand U1241 (N_1241,N_778,N_1008);
nor U1242 (N_1242,N_1086,N_835);
and U1243 (N_1243,N_1077,N_1076);
nor U1244 (N_1244,N_1113,N_836);
nand U1245 (N_1245,N_773,N_1068);
or U1246 (N_1246,N_743,N_1126);
or U1247 (N_1247,N_1161,N_715);
nand U1248 (N_1248,N_720,N_783);
nor U1249 (N_1249,N_985,N_1065);
nand U1250 (N_1250,N_1078,N_744);
nor U1251 (N_1251,N_764,N_870);
or U1252 (N_1252,N_872,N_1180);
nand U1253 (N_1253,N_1186,N_840);
and U1254 (N_1254,N_1122,N_722);
nor U1255 (N_1255,N_955,N_1178);
and U1256 (N_1256,N_665,N_622);
nand U1257 (N_1257,N_1133,N_811);
or U1258 (N_1258,N_957,N_925);
and U1259 (N_1259,N_677,N_1193);
and U1260 (N_1260,N_659,N_890);
or U1261 (N_1261,N_634,N_1172);
nor U1262 (N_1262,N_1173,N_908);
and U1263 (N_1263,N_996,N_650);
nor U1264 (N_1264,N_915,N_612);
nor U1265 (N_1265,N_749,N_754);
nand U1266 (N_1266,N_816,N_833);
and U1267 (N_1267,N_1088,N_879);
and U1268 (N_1268,N_777,N_938);
nand U1269 (N_1269,N_927,N_799);
nand U1270 (N_1270,N_1147,N_920);
or U1271 (N_1271,N_637,N_668);
nand U1272 (N_1272,N_1168,N_1030);
or U1273 (N_1273,N_714,N_683);
or U1274 (N_1274,N_1058,N_784);
nand U1275 (N_1275,N_748,N_1170);
nor U1276 (N_1276,N_1091,N_818);
nand U1277 (N_1277,N_948,N_643);
nand U1278 (N_1278,N_769,N_853);
nand U1279 (N_1279,N_1101,N_984);
and U1280 (N_1280,N_889,N_793);
nor U1281 (N_1281,N_1032,N_997);
nor U1282 (N_1282,N_841,N_1092);
nand U1283 (N_1283,N_1039,N_953);
or U1284 (N_1284,N_1070,N_660);
nor U1285 (N_1285,N_724,N_1176);
nand U1286 (N_1286,N_991,N_687);
nand U1287 (N_1287,N_707,N_856);
nand U1288 (N_1288,N_1081,N_1062);
or U1289 (N_1289,N_717,N_819);
and U1290 (N_1290,N_797,N_849);
nand U1291 (N_1291,N_1066,N_847);
nor U1292 (N_1292,N_747,N_852);
or U1293 (N_1293,N_1162,N_1118);
or U1294 (N_1294,N_831,N_671);
nor U1295 (N_1295,N_1006,N_974);
nor U1296 (N_1296,N_615,N_1020);
or U1297 (N_1297,N_961,N_979);
or U1298 (N_1298,N_1109,N_860);
nor U1299 (N_1299,N_1019,N_804);
nand U1300 (N_1300,N_788,N_1014);
and U1301 (N_1301,N_854,N_845);
nand U1302 (N_1302,N_969,N_970);
nor U1303 (N_1303,N_959,N_1029);
nand U1304 (N_1304,N_1067,N_672);
xnor U1305 (N_1305,N_881,N_857);
nor U1306 (N_1306,N_1073,N_994);
and U1307 (N_1307,N_894,N_1181);
and U1308 (N_1308,N_805,N_1187);
or U1309 (N_1309,N_791,N_1139);
nand U1310 (N_1310,N_776,N_990);
and U1311 (N_1311,N_851,N_976);
or U1312 (N_1312,N_617,N_1069);
and U1313 (N_1313,N_1027,N_691);
nand U1314 (N_1314,N_718,N_1198);
or U1315 (N_1315,N_873,N_897);
nor U1316 (N_1316,N_1185,N_954);
nor U1317 (N_1317,N_971,N_1143);
nor U1318 (N_1318,N_763,N_843);
nand U1319 (N_1319,N_821,N_792);
nor U1320 (N_1320,N_832,N_815);
nand U1321 (N_1321,N_1123,N_877);
nor U1322 (N_1322,N_709,N_760);
nand U1323 (N_1323,N_995,N_1061);
nand U1324 (N_1324,N_1104,N_1130);
nand U1325 (N_1325,N_980,N_1097);
nor U1326 (N_1326,N_912,N_886);
nand U1327 (N_1327,N_1131,N_610);
nor U1328 (N_1328,N_605,N_1046);
nand U1329 (N_1329,N_1024,N_770);
nor U1330 (N_1330,N_733,N_1085);
and U1331 (N_1331,N_694,N_962);
nand U1332 (N_1332,N_892,N_936);
nor U1333 (N_1333,N_726,N_1051);
and U1334 (N_1334,N_848,N_1044);
and U1335 (N_1335,N_716,N_855);
and U1336 (N_1336,N_1112,N_1140);
nand U1337 (N_1337,N_1037,N_940);
or U1338 (N_1338,N_690,N_1119);
and U1339 (N_1339,N_898,N_956);
nand U1340 (N_1340,N_738,N_647);
nor U1341 (N_1341,N_675,N_633);
or U1342 (N_1342,N_1188,N_623);
nor U1343 (N_1343,N_928,N_1174);
and U1344 (N_1344,N_711,N_875);
or U1345 (N_1345,N_1064,N_1111);
nor U1346 (N_1346,N_922,N_1045);
nand U1347 (N_1347,N_1115,N_1013);
and U1348 (N_1348,N_1128,N_850);
and U1349 (N_1349,N_1169,N_1175);
nand U1350 (N_1350,N_752,N_905);
nand U1351 (N_1351,N_829,N_1184);
and U1352 (N_1352,N_758,N_775);
nor U1353 (N_1353,N_900,N_1098);
nor U1354 (N_1354,N_1035,N_745);
nor U1355 (N_1355,N_917,N_1054);
and U1356 (N_1356,N_712,N_1132);
nand U1357 (N_1357,N_1144,N_1056);
nand U1358 (N_1358,N_680,N_621);
nand U1359 (N_1359,N_930,N_1049);
nor U1360 (N_1360,N_771,N_986);
or U1361 (N_1361,N_878,N_772);
nand U1362 (N_1362,N_869,N_998);
nand U1363 (N_1363,N_866,N_713);
or U1364 (N_1364,N_787,N_658);
nand U1365 (N_1365,N_732,N_601);
and U1366 (N_1366,N_1087,N_1004);
nand U1367 (N_1367,N_803,N_884);
nand U1368 (N_1368,N_1021,N_685);
nand U1369 (N_1369,N_973,N_641);
and U1370 (N_1370,N_1141,N_727);
or U1371 (N_1371,N_828,N_1142);
or U1372 (N_1372,N_846,N_891);
or U1373 (N_1373,N_1116,N_746);
nand U1374 (N_1374,N_876,N_1164);
nand U1375 (N_1375,N_666,N_686);
or U1376 (N_1376,N_708,N_1057);
and U1377 (N_1377,N_669,N_636);
nand U1378 (N_1378,N_688,N_1136);
nand U1379 (N_1379,N_1190,N_1157);
nand U1380 (N_1380,N_826,N_741);
or U1381 (N_1381,N_858,N_1022);
or U1382 (N_1382,N_790,N_862);
nand U1383 (N_1383,N_887,N_1033);
and U1384 (N_1384,N_618,N_1007);
nor U1385 (N_1385,N_649,N_983);
or U1386 (N_1386,N_624,N_616);
and U1387 (N_1387,N_904,N_604);
or U1388 (N_1388,N_739,N_918);
and U1389 (N_1389,N_1106,N_939);
and U1390 (N_1390,N_721,N_934);
and U1391 (N_1391,N_653,N_921);
nand U1392 (N_1392,N_824,N_992);
nor U1393 (N_1393,N_838,N_639);
nand U1394 (N_1394,N_631,N_1196);
and U1395 (N_1395,N_1127,N_627);
or U1396 (N_1396,N_1199,N_1018);
and U1397 (N_1397,N_950,N_662);
nor U1398 (N_1398,N_1100,N_696);
nand U1399 (N_1399,N_1011,N_981);
and U1400 (N_1400,N_902,N_867);
or U1401 (N_1401,N_914,N_684);
nor U1402 (N_1402,N_931,N_1192);
nand U1403 (N_1403,N_1000,N_896);
or U1404 (N_1404,N_678,N_728);
nand U1405 (N_1405,N_699,N_1028);
nor U1406 (N_1406,N_1083,N_972);
and U1407 (N_1407,N_893,N_885);
nand U1408 (N_1408,N_1023,N_664);
or U1409 (N_1409,N_1121,N_767);
and U1410 (N_1410,N_999,N_638);
nand U1411 (N_1411,N_642,N_975);
or U1412 (N_1412,N_700,N_945);
nand U1413 (N_1413,N_663,N_646);
or U1414 (N_1414,N_913,N_1084);
nor U1415 (N_1415,N_730,N_817);
or U1416 (N_1416,N_895,N_1005);
nor U1417 (N_1417,N_1009,N_786);
and U1418 (N_1418,N_1050,N_809);
nand U1419 (N_1419,N_785,N_1197);
nor U1420 (N_1420,N_907,N_736);
and U1421 (N_1421,N_798,N_628);
nand U1422 (N_1422,N_1063,N_1195);
nor U1423 (N_1423,N_1079,N_606);
nor U1424 (N_1424,N_1052,N_1041);
and U1425 (N_1425,N_657,N_943);
nand U1426 (N_1426,N_1089,N_864);
nand U1427 (N_1427,N_651,N_734);
nand U1428 (N_1428,N_737,N_1124);
and U1429 (N_1429,N_1182,N_1074);
and U1430 (N_1430,N_1090,N_949);
or U1431 (N_1431,N_1025,N_725);
or U1432 (N_1432,N_766,N_756);
nand U1433 (N_1433,N_689,N_1148);
nand U1434 (N_1434,N_757,N_656);
nor U1435 (N_1435,N_947,N_1040);
nor U1436 (N_1436,N_808,N_1156);
nand U1437 (N_1437,N_702,N_909);
nand U1438 (N_1438,N_1099,N_812);
or U1439 (N_1439,N_901,N_1110);
nand U1440 (N_1440,N_1135,N_1107);
and U1441 (N_1441,N_993,N_1150);
or U1442 (N_1442,N_761,N_735);
and U1443 (N_1443,N_1152,N_871);
or U1444 (N_1444,N_781,N_1042);
nor U1445 (N_1445,N_753,N_977);
nor U1446 (N_1446,N_1095,N_1134);
nand U1447 (N_1447,N_842,N_652);
nand U1448 (N_1448,N_1105,N_982);
or U1449 (N_1449,N_1102,N_1177);
and U1450 (N_1450,N_800,N_704);
nor U1451 (N_1451,N_705,N_1015);
nor U1452 (N_1452,N_1080,N_762);
or U1453 (N_1453,N_1151,N_827);
and U1454 (N_1454,N_1016,N_1163);
or U1455 (N_1455,N_911,N_1189);
or U1456 (N_1456,N_1138,N_1171);
nand U1457 (N_1457,N_1166,N_1034);
and U1458 (N_1458,N_807,N_654);
and U1459 (N_1459,N_837,N_600);
and U1460 (N_1460,N_888,N_774);
and U1461 (N_1461,N_865,N_1043);
xor U1462 (N_1462,N_863,N_782);
and U1463 (N_1463,N_740,N_899);
nand U1464 (N_1464,N_924,N_701);
nand U1465 (N_1465,N_603,N_1129);
or U1466 (N_1466,N_679,N_673);
nor U1467 (N_1467,N_620,N_910);
or U1468 (N_1468,N_964,N_1072);
nand U1469 (N_1469,N_923,N_874);
nand U1470 (N_1470,N_813,N_645);
nand U1471 (N_1471,N_814,N_1117);
nand U1472 (N_1472,N_952,N_695);
nor U1473 (N_1473,N_825,N_1048);
and U1474 (N_1474,N_1160,N_839);
nand U1475 (N_1475,N_1103,N_609);
or U1476 (N_1476,N_929,N_978);
xor U1477 (N_1477,N_648,N_906);
nor U1478 (N_1478,N_834,N_1096);
or U1479 (N_1479,N_966,N_801);
or U1480 (N_1480,N_697,N_1183);
nor U1481 (N_1481,N_667,N_916);
nor U1482 (N_1482,N_941,N_693);
or U1483 (N_1483,N_968,N_965);
and U1484 (N_1484,N_1001,N_682);
and U1485 (N_1485,N_640,N_1108);
and U1486 (N_1486,N_765,N_1036);
nor U1487 (N_1487,N_676,N_796);
nand U1488 (N_1488,N_830,N_1194);
or U1489 (N_1489,N_655,N_692);
or U1490 (N_1490,N_755,N_1155);
nor U1491 (N_1491,N_820,N_681);
nand U1492 (N_1492,N_794,N_723);
nor U1493 (N_1493,N_629,N_795);
and U1494 (N_1494,N_644,N_1114);
and U1495 (N_1495,N_698,N_868);
or U1496 (N_1496,N_611,N_1055);
nor U1497 (N_1497,N_750,N_779);
and U1498 (N_1498,N_932,N_710);
nand U1499 (N_1499,N_1071,N_958);
and U1500 (N_1500,N_746,N_792);
and U1501 (N_1501,N_874,N_843);
nor U1502 (N_1502,N_1146,N_931);
nand U1503 (N_1503,N_1099,N_870);
and U1504 (N_1504,N_1163,N_1188);
nand U1505 (N_1505,N_736,N_901);
nand U1506 (N_1506,N_1086,N_631);
or U1507 (N_1507,N_878,N_1102);
and U1508 (N_1508,N_1046,N_674);
and U1509 (N_1509,N_1003,N_781);
nand U1510 (N_1510,N_865,N_837);
or U1511 (N_1511,N_970,N_783);
and U1512 (N_1512,N_750,N_1124);
nand U1513 (N_1513,N_830,N_1146);
nor U1514 (N_1514,N_682,N_730);
and U1515 (N_1515,N_647,N_747);
and U1516 (N_1516,N_975,N_861);
nand U1517 (N_1517,N_1089,N_1156);
and U1518 (N_1518,N_642,N_813);
and U1519 (N_1519,N_1125,N_942);
or U1520 (N_1520,N_675,N_1035);
nand U1521 (N_1521,N_1075,N_813);
or U1522 (N_1522,N_844,N_782);
and U1523 (N_1523,N_828,N_1154);
and U1524 (N_1524,N_799,N_1180);
and U1525 (N_1525,N_1073,N_1031);
and U1526 (N_1526,N_695,N_1042);
nor U1527 (N_1527,N_1086,N_980);
nor U1528 (N_1528,N_1060,N_960);
nor U1529 (N_1529,N_624,N_1181);
or U1530 (N_1530,N_1082,N_1060);
nand U1531 (N_1531,N_850,N_1090);
and U1532 (N_1532,N_773,N_849);
nor U1533 (N_1533,N_656,N_1087);
nand U1534 (N_1534,N_974,N_939);
and U1535 (N_1535,N_767,N_1197);
nor U1536 (N_1536,N_716,N_1081);
nand U1537 (N_1537,N_960,N_999);
or U1538 (N_1538,N_1154,N_845);
nor U1539 (N_1539,N_1025,N_1018);
nor U1540 (N_1540,N_1122,N_897);
or U1541 (N_1541,N_1015,N_872);
nor U1542 (N_1542,N_795,N_1095);
nor U1543 (N_1543,N_1070,N_650);
nand U1544 (N_1544,N_640,N_768);
and U1545 (N_1545,N_765,N_1136);
and U1546 (N_1546,N_850,N_699);
nand U1547 (N_1547,N_780,N_893);
or U1548 (N_1548,N_857,N_957);
and U1549 (N_1549,N_660,N_814);
nor U1550 (N_1550,N_889,N_833);
and U1551 (N_1551,N_953,N_1103);
and U1552 (N_1552,N_973,N_797);
nand U1553 (N_1553,N_666,N_1170);
nand U1554 (N_1554,N_973,N_778);
nor U1555 (N_1555,N_782,N_1092);
nor U1556 (N_1556,N_761,N_743);
nor U1557 (N_1557,N_807,N_673);
nor U1558 (N_1558,N_850,N_984);
and U1559 (N_1559,N_1051,N_1056);
nor U1560 (N_1560,N_601,N_605);
nor U1561 (N_1561,N_661,N_873);
nand U1562 (N_1562,N_1147,N_766);
and U1563 (N_1563,N_615,N_1095);
nor U1564 (N_1564,N_845,N_739);
and U1565 (N_1565,N_977,N_915);
nand U1566 (N_1566,N_618,N_716);
or U1567 (N_1567,N_666,N_1183);
or U1568 (N_1568,N_673,N_832);
nor U1569 (N_1569,N_629,N_1087);
and U1570 (N_1570,N_944,N_1124);
or U1571 (N_1571,N_1076,N_744);
or U1572 (N_1572,N_737,N_968);
nand U1573 (N_1573,N_780,N_736);
nand U1574 (N_1574,N_619,N_1039);
nand U1575 (N_1575,N_1044,N_896);
nor U1576 (N_1576,N_1051,N_859);
or U1577 (N_1577,N_794,N_864);
or U1578 (N_1578,N_722,N_816);
nor U1579 (N_1579,N_979,N_879);
and U1580 (N_1580,N_722,N_931);
nor U1581 (N_1581,N_606,N_848);
or U1582 (N_1582,N_1126,N_752);
nand U1583 (N_1583,N_831,N_948);
nand U1584 (N_1584,N_629,N_1148);
or U1585 (N_1585,N_961,N_1144);
or U1586 (N_1586,N_829,N_735);
nor U1587 (N_1587,N_903,N_711);
nand U1588 (N_1588,N_685,N_654);
nand U1589 (N_1589,N_926,N_1136);
nand U1590 (N_1590,N_886,N_960);
and U1591 (N_1591,N_1062,N_1072);
nand U1592 (N_1592,N_646,N_696);
and U1593 (N_1593,N_1074,N_888);
nor U1594 (N_1594,N_874,N_692);
or U1595 (N_1595,N_1118,N_1032);
or U1596 (N_1596,N_715,N_898);
nor U1597 (N_1597,N_792,N_737);
nand U1598 (N_1598,N_1155,N_765);
or U1599 (N_1599,N_923,N_604);
nor U1600 (N_1600,N_1054,N_867);
or U1601 (N_1601,N_630,N_993);
nand U1602 (N_1602,N_638,N_1089);
and U1603 (N_1603,N_1063,N_877);
or U1604 (N_1604,N_1003,N_1024);
nand U1605 (N_1605,N_1097,N_897);
and U1606 (N_1606,N_886,N_1102);
nor U1607 (N_1607,N_1063,N_853);
nand U1608 (N_1608,N_1126,N_618);
and U1609 (N_1609,N_1147,N_611);
and U1610 (N_1610,N_1150,N_1164);
nand U1611 (N_1611,N_800,N_678);
xor U1612 (N_1612,N_906,N_1119);
nand U1613 (N_1613,N_787,N_862);
and U1614 (N_1614,N_988,N_662);
nor U1615 (N_1615,N_969,N_1194);
nand U1616 (N_1616,N_894,N_984);
nor U1617 (N_1617,N_1017,N_959);
and U1618 (N_1618,N_1093,N_1055);
nor U1619 (N_1619,N_991,N_910);
or U1620 (N_1620,N_660,N_1061);
or U1621 (N_1621,N_707,N_943);
nor U1622 (N_1622,N_600,N_1139);
nor U1623 (N_1623,N_650,N_677);
nand U1624 (N_1624,N_1126,N_1027);
nand U1625 (N_1625,N_606,N_835);
and U1626 (N_1626,N_932,N_918);
and U1627 (N_1627,N_922,N_679);
and U1628 (N_1628,N_1176,N_742);
nor U1629 (N_1629,N_823,N_1105);
and U1630 (N_1630,N_1041,N_914);
or U1631 (N_1631,N_903,N_959);
nand U1632 (N_1632,N_771,N_758);
nand U1633 (N_1633,N_911,N_925);
nor U1634 (N_1634,N_923,N_1161);
and U1635 (N_1635,N_778,N_791);
or U1636 (N_1636,N_675,N_816);
nor U1637 (N_1637,N_1089,N_835);
nand U1638 (N_1638,N_775,N_1097);
nor U1639 (N_1639,N_1103,N_606);
and U1640 (N_1640,N_961,N_880);
or U1641 (N_1641,N_973,N_1000);
and U1642 (N_1642,N_943,N_1105);
or U1643 (N_1643,N_860,N_955);
or U1644 (N_1644,N_934,N_720);
nor U1645 (N_1645,N_1134,N_769);
nand U1646 (N_1646,N_758,N_859);
and U1647 (N_1647,N_990,N_912);
or U1648 (N_1648,N_1181,N_635);
nor U1649 (N_1649,N_604,N_818);
nor U1650 (N_1650,N_1185,N_964);
and U1651 (N_1651,N_866,N_928);
nand U1652 (N_1652,N_735,N_1116);
nand U1653 (N_1653,N_1022,N_740);
nor U1654 (N_1654,N_977,N_1085);
nand U1655 (N_1655,N_931,N_935);
nand U1656 (N_1656,N_809,N_1122);
nand U1657 (N_1657,N_1012,N_1044);
and U1658 (N_1658,N_1156,N_635);
nor U1659 (N_1659,N_683,N_868);
nor U1660 (N_1660,N_1168,N_1102);
nand U1661 (N_1661,N_1072,N_757);
nor U1662 (N_1662,N_1089,N_1044);
nor U1663 (N_1663,N_1024,N_1172);
or U1664 (N_1664,N_844,N_1164);
nor U1665 (N_1665,N_801,N_887);
and U1666 (N_1666,N_1033,N_1015);
and U1667 (N_1667,N_674,N_881);
nand U1668 (N_1668,N_1094,N_654);
nand U1669 (N_1669,N_839,N_945);
or U1670 (N_1670,N_873,N_1142);
nor U1671 (N_1671,N_1043,N_1059);
or U1672 (N_1672,N_1119,N_951);
nand U1673 (N_1673,N_680,N_913);
or U1674 (N_1674,N_847,N_715);
or U1675 (N_1675,N_999,N_996);
and U1676 (N_1676,N_836,N_1114);
nand U1677 (N_1677,N_879,N_956);
nand U1678 (N_1678,N_1145,N_769);
and U1679 (N_1679,N_1071,N_615);
nor U1680 (N_1680,N_835,N_1047);
nand U1681 (N_1681,N_717,N_1123);
xor U1682 (N_1682,N_965,N_957);
or U1683 (N_1683,N_691,N_892);
nand U1684 (N_1684,N_1068,N_1146);
nand U1685 (N_1685,N_1017,N_814);
nand U1686 (N_1686,N_977,N_1037);
nand U1687 (N_1687,N_616,N_630);
and U1688 (N_1688,N_968,N_1148);
and U1689 (N_1689,N_613,N_1015);
nand U1690 (N_1690,N_1163,N_1031);
or U1691 (N_1691,N_762,N_898);
or U1692 (N_1692,N_639,N_1075);
nand U1693 (N_1693,N_1030,N_870);
or U1694 (N_1694,N_947,N_662);
and U1695 (N_1695,N_1192,N_1131);
nand U1696 (N_1696,N_604,N_723);
or U1697 (N_1697,N_807,N_1073);
and U1698 (N_1698,N_795,N_668);
and U1699 (N_1699,N_1021,N_765);
nand U1700 (N_1700,N_983,N_729);
or U1701 (N_1701,N_949,N_804);
nand U1702 (N_1702,N_1073,N_822);
or U1703 (N_1703,N_1153,N_1004);
nor U1704 (N_1704,N_960,N_1107);
and U1705 (N_1705,N_1014,N_623);
and U1706 (N_1706,N_927,N_970);
nand U1707 (N_1707,N_860,N_639);
and U1708 (N_1708,N_1183,N_871);
or U1709 (N_1709,N_913,N_1064);
or U1710 (N_1710,N_966,N_1069);
nor U1711 (N_1711,N_806,N_1101);
nand U1712 (N_1712,N_689,N_1169);
nor U1713 (N_1713,N_996,N_776);
nor U1714 (N_1714,N_713,N_925);
and U1715 (N_1715,N_609,N_929);
nor U1716 (N_1716,N_1011,N_660);
nor U1717 (N_1717,N_875,N_1154);
or U1718 (N_1718,N_633,N_1090);
nor U1719 (N_1719,N_1023,N_608);
and U1720 (N_1720,N_1088,N_624);
and U1721 (N_1721,N_871,N_988);
nand U1722 (N_1722,N_991,N_946);
or U1723 (N_1723,N_895,N_1034);
and U1724 (N_1724,N_851,N_634);
nor U1725 (N_1725,N_1019,N_778);
or U1726 (N_1726,N_1136,N_733);
or U1727 (N_1727,N_606,N_893);
and U1728 (N_1728,N_858,N_848);
nor U1729 (N_1729,N_940,N_789);
nand U1730 (N_1730,N_951,N_1179);
or U1731 (N_1731,N_1004,N_1159);
nand U1732 (N_1732,N_946,N_624);
nor U1733 (N_1733,N_1040,N_1072);
nor U1734 (N_1734,N_873,N_903);
nand U1735 (N_1735,N_948,N_1194);
and U1736 (N_1736,N_679,N_822);
nand U1737 (N_1737,N_783,N_900);
and U1738 (N_1738,N_682,N_741);
nand U1739 (N_1739,N_764,N_1135);
nand U1740 (N_1740,N_837,N_1032);
and U1741 (N_1741,N_960,N_926);
or U1742 (N_1742,N_990,N_987);
or U1743 (N_1743,N_1098,N_601);
or U1744 (N_1744,N_697,N_1114);
or U1745 (N_1745,N_683,N_712);
and U1746 (N_1746,N_1091,N_1141);
or U1747 (N_1747,N_939,N_1072);
nand U1748 (N_1748,N_1037,N_742);
nand U1749 (N_1749,N_738,N_620);
and U1750 (N_1750,N_829,N_883);
nor U1751 (N_1751,N_637,N_988);
nand U1752 (N_1752,N_1077,N_1074);
or U1753 (N_1753,N_1156,N_846);
and U1754 (N_1754,N_948,N_762);
nor U1755 (N_1755,N_607,N_923);
or U1756 (N_1756,N_1154,N_1024);
or U1757 (N_1757,N_809,N_1077);
or U1758 (N_1758,N_725,N_1197);
or U1759 (N_1759,N_712,N_909);
nand U1760 (N_1760,N_847,N_1008);
nor U1761 (N_1761,N_1186,N_695);
nor U1762 (N_1762,N_1188,N_770);
nor U1763 (N_1763,N_635,N_814);
or U1764 (N_1764,N_1187,N_846);
nor U1765 (N_1765,N_1040,N_962);
nand U1766 (N_1766,N_833,N_840);
and U1767 (N_1767,N_880,N_840);
or U1768 (N_1768,N_1133,N_1036);
nand U1769 (N_1769,N_955,N_929);
nor U1770 (N_1770,N_1069,N_801);
nor U1771 (N_1771,N_1116,N_825);
nand U1772 (N_1772,N_1103,N_809);
and U1773 (N_1773,N_691,N_1101);
nand U1774 (N_1774,N_1039,N_985);
nor U1775 (N_1775,N_888,N_713);
nand U1776 (N_1776,N_700,N_1148);
and U1777 (N_1777,N_659,N_1084);
and U1778 (N_1778,N_1041,N_865);
or U1779 (N_1779,N_749,N_882);
nor U1780 (N_1780,N_966,N_1012);
xnor U1781 (N_1781,N_745,N_1005);
or U1782 (N_1782,N_973,N_857);
or U1783 (N_1783,N_687,N_864);
nor U1784 (N_1784,N_750,N_782);
and U1785 (N_1785,N_946,N_868);
nand U1786 (N_1786,N_815,N_1149);
nand U1787 (N_1787,N_838,N_637);
or U1788 (N_1788,N_772,N_746);
nand U1789 (N_1789,N_801,N_725);
or U1790 (N_1790,N_770,N_1161);
or U1791 (N_1791,N_1077,N_834);
xnor U1792 (N_1792,N_704,N_807);
nor U1793 (N_1793,N_761,N_732);
nand U1794 (N_1794,N_1060,N_1107);
or U1795 (N_1795,N_704,N_918);
nor U1796 (N_1796,N_939,N_907);
or U1797 (N_1797,N_737,N_808);
and U1798 (N_1798,N_895,N_812);
nand U1799 (N_1799,N_873,N_882);
and U1800 (N_1800,N_1522,N_1301);
nand U1801 (N_1801,N_1450,N_1518);
nand U1802 (N_1802,N_1405,N_1656);
or U1803 (N_1803,N_1508,N_1299);
nor U1804 (N_1804,N_1429,N_1676);
nor U1805 (N_1805,N_1385,N_1602);
and U1806 (N_1806,N_1487,N_1747);
or U1807 (N_1807,N_1681,N_1729);
or U1808 (N_1808,N_1368,N_1332);
nor U1809 (N_1809,N_1463,N_1734);
and U1810 (N_1810,N_1361,N_1346);
nor U1811 (N_1811,N_1239,N_1709);
nand U1812 (N_1812,N_1467,N_1349);
or U1813 (N_1813,N_1704,N_1410);
and U1814 (N_1814,N_1271,N_1644);
nand U1815 (N_1815,N_1531,N_1351);
nand U1816 (N_1816,N_1678,N_1295);
nand U1817 (N_1817,N_1314,N_1481);
nor U1818 (N_1818,N_1534,N_1521);
nand U1819 (N_1819,N_1697,N_1698);
nand U1820 (N_1820,N_1752,N_1660);
nor U1821 (N_1821,N_1461,N_1366);
nand U1822 (N_1822,N_1473,N_1695);
and U1823 (N_1823,N_1782,N_1613);
nand U1824 (N_1824,N_1370,N_1603);
nand U1825 (N_1825,N_1633,N_1503);
nand U1826 (N_1826,N_1340,N_1722);
nor U1827 (N_1827,N_1587,N_1251);
and U1828 (N_1828,N_1737,N_1680);
nand U1829 (N_1829,N_1427,N_1624);
or U1830 (N_1830,N_1262,N_1650);
nor U1831 (N_1831,N_1542,N_1514);
nor U1832 (N_1832,N_1399,N_1341);
nor U1833 (N_1833,N_1753,N_1780);
and U1834 (N_1834,N_1581,N_1327);
nand U1835 (N_1835,N_1770,N_1592);
nor U1836 (N_1836,N_1528,N_1312);
and U1837 (N_1837,N_1758,N_1474);
nand U1838 (N_1838,N_1347,N_1649);
or U1839 (N_1839,N_1754,N_1721);
or U1840 (N_1840,N_1775,N_1537);
nor U1841 (N_1841,N_1478,N_1710);
xnor U1842 (N_1842,N_1339,N_1438);
nor U1843 (N_1843,N_1549,N_1557);
or U1844 (N_1844,N_1502,N_1672);
or U1845 (N_1845,N_1477,N_1310);
and U1846 (N_1846,N_1714,N_1456);
nor U1847 (N_1847,N_1589,N_1673);
or U1848 (N_1848,N_1416,N_1631);
nor U1849 (N_1849,N_1716,N_1488);
or U1850 (N_1850,N_1317,N_1376);
or U1851 (N_1851,N_1509,N_1543);
or U1852 (N_1852,N_1216,N_1261);
nor U1853 (N_1853,N_1516,N_1595);
or U1854 (N_1854,N_1789,N_1621);
nor U1855 (N_1855,N_1367,N_1764);
or U1856 (N_1856,N_1428,N_1215);
or U1857 (N_1857,N_1316,N_1238);
nand U1858 (N_1858,N_1523,N_1558);
and U1859 (N_1859,N_1415,N_1241);
and U1860 (N_1860,N_1344,N_1419);
nor U1861 (N_1861,N_1425,N_1568);
and U1862 (N_1862,N_1496,N_1283);
or U1863 (N_1863,N_1433,N_1690);
or U1864 (N_1864,N_1622,N_1607);
nor U1865 (N_1865,N_1653,N_1320);
nand U1866 (N_1866,N_1363,N_1772);
and U1867 (N_1867,N_1640,N_1281);
or U1868 (N_1868,N_1655,N_1381);
nor U1869 (N_1869,N_1489,N_1548);
or U1870 (N_1870,N_1658,N_1342);
nand U1871 (N_1871,N_1634,N_1535);
xnor U1872 (N_1872,N_1675,N_1407);
nor U1873 (N_1873,N_1297,N_1619);
and U1874 (N_1874,N_1554,N_1318);
nor U1875 (N_1875,N_1530,N_1757);
nand U1876 (N_1876,N_1616,N_1377);
and U1877 (N_1877,N_1545,N_1499);
or U1878 (N_1878,N_1232,N_1420);
or U1879 (N_1879,N_1769,N_1552);
nor U1880 (N_1880,N_1766,N_1401);
nor U1881 (N_1881,N_1491,N_1765);
and U1882 (N_1882,N_1541,N_1567);
nor U1883 (N_1883,N_1390,N_1533);
xor U1884 (N_1884,N_1564,N_1276);
nor U1885 (N_1885,N_1486,N_1388);
nand U1886 (N_1886,N_1739,N_1268);
and U1887 (N_1887,N_1696,N_1771);
nand U1888 (N_1888,N_1451,N_1750);
or U1889 (N_1889,N_1468,N_1479);
nor U1890 (N_1890,N_1609,N_1735);
or U1891 (N_1891,N_1235,N_1392);
or U1892 (N_1892,N_1434,N_1665);
nor U1893 (N_1893,N_1718,N_1453);
or U1894 (N_1894,N_1610,N_1788);
nand U1895 (N_1895,N_1406,N_1569);
nor U1896 (N_1896,N_1457,N_1555);
nor U1897 (N_1897,N_1620,N_1638);
nor U1898 (N_1898,N_1266,N_1500);
or U1899 (N_1899,N_1454,N_1286);
nand U1900 (N_1900,N_1231,N_1490);
and U1901 (N_1901,N_1439,N_1713);
nand U1902 (N_1902,N_1412,N_1730);
or U1903 (N_1903,N_1354,N_1424);
or U1904 (N_1904,N_1413,N_1661);
nand U1905 (N_1905,N_1662,N_1596);
nor U1906 (N_1906,N_1645,N_1411);
and U1907 (N_1907,N_1220,N_1515);
and U1908 (N_1908,N_1498,N_1207);
and U1909 (N_1909,N_1641,N_1458);
nand U1910 (N_1910,N_1594,N_1601);
nor U1911 (N_1911,N_1396,N_1611);
or U1912 (N_1912,N_1728,N_1374);
or U1913 (N_1913,N_1355,N_1623);
nand U1914 (N_1914,N_1677,N_1513);
and U1915 (N_1915,N_1493,N_1325);
and U1916 (N_1916,N_1761,N_1781);
nand U1917 (N_1917,N_1570,N_1201);
or U1918 (N_1918,N_1315,N_1553);
nor U1919 (N_1919,N_1445,N_1257);
and U1920 (N_1920,N_1466,N_1391);
and U1921 (N_1921,N_1475,N_1352);
nand U1922 (N_1922,N_1205,N_1504);
or U1923 (N_1923,N_1336,N_1637);
nor U1924 (N_1924,N_1560,N_1359);
xor U1925 (N_1925,N_1308,N_1218);
nor U1926 (N_1926,N_1208,N_1236);
and U1927 (N_1927,N_1703,N_1795);
and U1928 (N_1928,N_1269,N_1706);
or U1929 (N_1929,N_1329,N_1459);
and U1930 (N_1930,N_1485,N_1224);
nand U1931 (N_1931,N_1615,N_1234);
and U1932 (N_1932,N_1628,N_1209);
nand U1933 (N_1933,N_1582,N_1304);
xor U1934 (N_1934,N_1626,N_1330);
nand U1935 (N_1935,N_1666,N_1360);
and U1936 (N_1936,N_1506,N_1501);
nor U1937 (N_1937,N_1432,N_1785);
nand U1938 (N_1938,N_1402,N_1512);
nand U1939 (N_1939,N_1260,N_1277);
nand U1940 (N_1940,N_1264,N_1408);
nand U1941 (N_1941,N_1300,N_1776);
nor U1942 (N_1942,N_1797,N_1612);
nand U1943 (N_1943,N_1302,N_1298);
and U1944 (N_1944,N_1394,N_1258);
nand U1945 (N_1945,N_1667,N_1751);
nor U1946 (N_1946,N_1383,N_1632);
nor U1947 (N_1947,N_1460,N_1723);
nand U1948 (N_1948,N_1293,N_1480);
nand U1949 (N_1949,N_1333,N_1326);
nand U1950 (N_1950,N_1719,N_1743);
nor U1951 (N_1951,N_1756,N_1223);
and U1952 (N_1952,N_1646,N_1384);
nor U1953 (N_1953,N_1296,N_1436);
or U1954 (N_1954,N_1538,N_1540);
nand U1955 (N_1955,N_1755,N_1219);
nand U1956 (N_1956,N_1294,N_1688);
nand U1957 (N_1957,N_1636,N_1353);
nor U1958 (N_1958,N_1767,N_1256);
and U1959 (N_1959,N_1430,N_1712);
nand U1960 (N_1960,N_1726,N_1711);
nand U1961 (N_1961,N_1448,N_1437);
or U1962 (N_1962,N_1275,N_1563);
nor U1963 (N_1963,N_1787,N_1572);
nand U1964 (N_1964,N_1455,N_1248);
nand U1965 (N_1965,N_1689,N_1606);
or U1966 (N_1966,N_1322,N_1762);
and U1967 (N_1967,N_1246,N_1778);
nand U1968 (N_1968,N_1544,N_1345);
and U1969 (N_1969,N_1497,N_1211);
or U1970 (N_1970,N_1417,N_1627);
and U1971 (N_1971,N_1289,N_1240);
and U1972 (N_1972,N_1337,N_1768);
nor U1973 (N_1973,N_1243,N_1259);
nor U1974 (N_1974,N_1715,N_1784);
and U1975 (N_1975,N_1674,N_1311);
nor U1976 (N_1976,N_1288,N_1278);
nand U1977 (N_1977,N_1447,N_1387);
nor U1978 (N_1978,N_1790,N_1323);
or U1979 (N_1979,N_1306,N_1604);
or U1980 (N_1980,N_1397,N_1577);
nor U1981 (N_1981,N_1287,N_1382);
nand U1982 (N_1982,N_1335,N_1559);
nand U1983 (N_1983,N_1204,N_1731);
xor U1984 (N_1984,N_1643,N_1793);
or U1985 (N_1985,N_1669,N_1692);
nand U1986 (N_1986,N_1472,N_1443);
or U1987 (N_1987,N_1575,N_1593);
nand U1988 (N_1988,N_1214,N_1249);
and U1989 (N_1989,N_1303,N_1629);
and U1990 (N_1990,N_1510,N_1244);
nor U1991 (N_1991,N_1449,N_1608);
nand U1992 (N_1992,N_1635,N_1422);
and U1993 (N_1993,N_1682,N_1319);
nand U1994 (N_1994,N_1727,N_1444);
xnor U1995 (N_1995,N_1328,N_1561);
and U1996 (N_1996,N_1740,N_1324);
or U1997 (N_1997,N_1597,N_1685);
nor U1998 (N_1998,N_1380,N_1442);
nor U1999 (N_1999,N_1483,N_1520);
or U2000 (N_2000,N_1639,N_1741);
nand U2001 (N_2001,N_1600,N_1441);
nand U2002 (N_2002,N_1663,N_1230);
and U2003 (N_2003,N_1724,N_1431);
xor U2004 (N_2004,N_1228,N_1398);
nor U2005 (N_2005,N_1524,N_1254);
or U2006 (N_2006,N_1505,N_1371);
and U2007 (N_2007,N_1423,N_1736);
nand U2008 (N_2008,N_1556,N_1253);
or U2009 (N_2009,N_1657,N_1748);
and U2010 (N_2010,N_1414,N_1774);
nor U2011 (N_2011,N_1378,N_1732);
nand U2012 (N_2012,N_1580,N_1792);
nor U2013 (N_2013,N_1791,N_1763);
and U2014 (N_2014,N_1562,N_1693);
or U2015 (N_2015,N_1309,N_1679);
or U2016 (N_2016,N_1700,N_1334);
or U2017 (N_2017,N_1794,N_1440);
xor U2018 (N_2018,N_1579,N_1465);
and U2019 (N_2019,N_1708,N_1694);
nand U2020 (N_2020,N_1511,N_1786);
or U2021 (N_2021,N_1527,N_1305);
and U2022 (N_2022,N_1222,N_1746);
and U2023 (N_2023,N_1773,N_1206);
nand U2024 (N_2024,N_1707,N_1494);
nand U2025 (N_2025,N_1670,N_1536);
nand U2026 (N_2026,N_1307,N_1242);
nand U2027 (N_2027,N_1725,N_1701);
nor U2028 (N_2028,N_1369,N_1446);
and U2029 (N_2029,N_1476,N_1282);
or U2030 (N_2030,N_1798,N_1668);
nor U2031 (N_2031,N_1280,N_1760);
nand U2032 (N_2032,N_1212,N_1225);
nor U2033 (N_2033,N_1226,N_1284);
nor U2034 (N_2034,N_1285,N_1270);
or U2035 (N_2035,N_1343,N_1364);
nor U2036 (N_2036,N_1221,N_1777);
nand U2037 (N_2037,N_1372,N_1614);
nor U2038 (N_2038,N_1588,N_1591);
or U2039 (N_2039,N_1686,N_1358);
or U2040 (N_2040,N_1691,N_1274);
nor U2041 (N_2041,N_1252,N_1452);
nand U2042 (N_2042,N_1617,N_1482);
nand U2043 (N_2043,N_1630,N_1373);
nor U2044 (N_2044,N_1571,N_1237);
or U2045 (N_2045,N_1495,N_1565);
and U2046 (N_2046,N_1599,N_1583);
nand U2047 (N_2047,N_1625,N_1550);
nor U2048 (N_2048,N_1464,N_1586);
nor U2049 (N_2049,N_1799,N_1210);
and U2050 (N_2050,N_1400,N_1338);
and U2051 (N_2051,N_1426,N_1203);
nand U2052 (N_2052,N_1759,N_1733);
xnor U2053 (N_2053,N_1532,N_1331);
or U2054 (N_2054,N_1738,N_1507);
nor U2055 (N_2055,N_1313,N_1539);
xor U2056 (N_2056,N_1403,N_1742);
nor U2057 (N_2057,N_1356,N_1365);
or U2058 (N_2058,N_1783,N_1267);
nor U2059 (N_2059,N_1265,N_1291);
or U2060 (N_2060,N_1749,N_1517);
or U2061 (N_2061,N_1470,N_1379);
or U2062 (N_2062,N_1664,N_1418);
nor U2063 (N_2063,N_1651,N_1605);
nand U2064 (N_2064,N_1566,N_1547);
nor U2065 (N_2065,N_1471,N_1350);
and U2066 (N_2066,N_1389,N_1551);
and U2067 (N_2067,N_1393,N_1717);
and U2068 (N_2068,N_1574,N_1654);
and U2069 (N_2069,N_1578,N_1421);
nand U2070 (N_2070,N_1386,N_1526);
and U2071 (N_2071,N_1642,N_1671);
nand U2072 (N_2072,N_1683,N_1321);
nand U2073 (N_2073,N_1279,N_1357);
or U2074 (N_2074,N_1529,N_1202);
and U2075 (N_2075,N_1705,N_1213);
or U2076 (N_2076,N_1229,N_1546);
or U2077 (N_2077,N_1598,N_1484);
and U2078 (N_2078,N_1492,N_1409);
or U2079 (N_2079,N_1779,N_1573);
nand U2080 (N_2080,N_1217,N_1745);
and U2081 (N_2081,N_1796,N_1584);
or U2082 (N_2082,N_1250,N_1348);
or U2083 (N_2083,N_1702,N_1469);
and U2084 (N_2084,N_1247,N_1618);
nor U2085 (N_2085,N_1263,N_1585);
nand U2086 (N_2086,N_1290,N_1375);
or U2087 (N_2087,N_1659,N_1233);
nand U2088 (N_2088,N_1647,N_1576);
nand U2089 (N_2089,N_1462,N_1687);
and U2090 (N_2090,N_1435,N_1404);
nand U2091 (N_2091,N_1684,N_1200);
or U2092 (N_2092,N_1255,N_1362);
nor U2093 (N_2093,N_1519,N_1652);
and U2094 (N_2094,N_1744,N_1525);
nor U2095 (N_2095,N_1273,N_1395);
nand U2096 (N_2096,N_1590,N_1648);
nand U2097 (N_2097,N_1245,N_1272);
nor U2098 (N_2098,N_1720,N_1292);
or U2099 (N_2099,N_1227,N_1699);
and U2100 (N_2100,N_1353,N_1646);
or U2101 (N_2101,N_1209,N_1313);
or U2102 (N_2102,N_1530,N_1344);
nor U2103 (N_2103,N_1522,N_1428);
nand U2104 (N_2104,N_1320,N_1448);
or U2105 (N_2105,N_1388,N_1499);
nor U2106 (N_2106,N_1450,N_1537);
nor U2107 (N_2107,N_1549,N_1648);
nor U2108 (N_2108,N_1685,N_1346);
nor U2109 (N_2109,N_1604,N_1768);
and U2110 (N_2110,N_1574,N_1345);
nand U2111 (N_2111,N_1729,N_1662);
nor U2112 (N_2112,N_1757,N_1289);
nand U2113 (N_2113,N_1243,N_1231);
or U2114 (N_2114,N_1577,N_1718);
or U2115 (N_2115,N_1631,N_1762);
nand U2116 (N_2116,N_1735,N_1627);
and U2117 (N_2117,N_1576,N_1776);
nand U2118 (N_2118,N_1366,N_1249);
xnor U2119 (N_2119,N_1530,N_1552);
nor U2120 (N_2120,N_1741,N_1346);
nand U2121 (N_2121,N_1336,N_1370);
or U2122 (N_2122,N_1309,N_1427);
nor U2123 (N_2123,N_1684,N_1673);
or U2124 (N_2124,N_1452,N_1732);
or U2125 (N_2125,N_1291,N_1594);
nand U2126 (N_2126,N_1221,N_1772);
and U2127 (N_2127,N_1432,N_1627);
nand U2128 (N_2128,N_1314,N_1442);
nor U2129 (N_2129,N_1609,N_1405);
nor U2130 (N_2130,N_1402,N_1682);
and U2131 (N_2131,N_1668,N_1649);
nand U2132 (N_2132,N_1718,N_1434);
and U2133 (N_2133,N_1592,N_1304);
nor U2134 (N_2134,N_1361,N_1271);
nand U2135 (N_2135,N_1750,N_1318);
or U2136 (N_2136,N_1537,N_1490);
and U2137 (N_2137,N_1481,N_1710);
or U2138 (N_2138,N_1286,N_1538);
or U2139 (N_2139,N_1522,N_1433);
or U2140 (N_2140,N_1575,N_1774);
or U2141 (N_2141,N_1516,N_1662);
and U2142 (N_2142,N_1652,N_1403);
or U2143 (N_2143,N_1380,N_1560);
nand U2144 (N_2144,N_1701,N_1411);
nand U2145 (N_2145,N_1387,N_1378);
and U2146 (N_2146,N_1245,N_1269);
or U2147 (N_2147,N_1406,N_1756);
nand U2148 (N_2148,N_1312,N_1748);
or U2149 (N_2149,N_1375,N_1349);
and U2150 (N_2150,N_1345,N_1760);
or U2151 (N_2151,N_1776,N_1588);
nor U2152 (N_2152,N_1586,N_1691);
and U2153 (N_2153,N_1650,N_1492);
or U2154 (N_2154,N_1559,N_1280);
and U2155 (N_2155,N_1703,N_1636);
or U2156 (N_2156,N_1611,N_1624);
and U2157 (N_2157,N_1667,N_1560);
and U2158 (N_2158,N_1269,N_1379);
or U2159 (N_2159,N_1514,N_1742);
nand U2160 (N_2160,N_1778,N_1646);
nand U2161 (N_2161,N_1342,N_1512);
nand U2162 (N_2162,N_1546,N_1612);
or U2163 (N_2163,N_1322,N_1585);
nor U2164 (N_2164,N_1735,N_1491);
and U2165 (N_2165,N_1413,N_1706);
and U2166 (N_2166,N_1776,N_1323);
and U2167 (N_2167,N_1439,N_1605);
and U2168 (N_2168,N_1610,N_1584);
nor U2169 (N_2169,N_1544,N_1573);
or U2170 (N_2170,N_1204,N_1229);
and U2171 (N_2171,N_1294,N_1521);
and U2172 (N_2172,N_1339,N_1291);
nor U2173 (N_2173,N_1476,N_1687);
and U2174 (N_2174,N_1451,N_1466);
or U2175 (N_2175,N_1236,N_1639);
or U2176 (N_2176,N_1525,N_1576);
and U2177 (N_2177,N_1426,N_1245);
nor U2178 (N_2178,N_1384,N_1661);
or U2179 (N_2179,N_1691,N_1480);
nand U2180 (N_2180,N_1785,N_1258);
nor U2181 (N_2181,N_1369,N_1551);
or U2182 (N_2182,N_1474,N_1239);
or U2183 (N_2183,N_1659,N_1627);
nand U2184 (N_2184,N_1446,N_1501);
and U2185 (N_2185,N_1517,N_1268);
and U2186 (N_2186,N_1507,N_1753);
nor U2187 (N_2187,N_1774,N_1374);
or U2188 (N_2188,N_1363,N_1634);
nor U2189 (N_2189,N_1477,N_1569);
nor U2190 (N_2190,N_1790,N_1346);
and U2191 (N_2191,N_1417,N_1280);
or U2192 (N_2192,N_1706,N_1450);
nor U2193 (N_2193,N_1672,N_1445);
nand U2194 (N_2194,N_1746,N_1724);
and U2195 (N_2195,N_1583,N_1470);
or U2196 (N_2196,N_1444,N_1539);
and U2197 (N_2197,N_1775,N_1345);
nand U2198 (N_2198,N_1231,N_1669);
nor U2199 (N_2199,N_1465,N_1708);
or U2200 (N_2200,N_1266,N_1666);
and U2201 (N_2201,N_1776,N_1689);
nand U2202 (N_2202,N_1699,N_1476);
nand U2203 (N_2203,N_1689,N_1653);
and U2204 (N_2204,N_1479,N_1228);
and U2205 (N_2205,N_1754,N_1542);
nor U2206 (N_2206,N_1641,N_1356);
nor U2207 (N_2207,N_1695,N_1419);
nor U2208 (N_2208,N_1611,N_1447);
nor U2209 (N_2209,N_1469,N_1367);
and U2210 (N_2210,N_1254,N_1544);
and U2211 (N_2211,N_1323,N_1205);
and U2212 (N_2212,N_1621,N_1319);
and U2213 (N_2213,N_1514,N_1690);
and U2214 (N_2214,N_1264,N_1213);
nor U2215 (N_2215,N_1442,N_1282);
and U2216 (N_2216,N_1277,N_1411);
nor U2217 (N_2217,N_1696,N_1399);
nand U2218 (N_2218,N_1580,N_1349);
nor U2219 (N_2219,N_1368,N_1260);
nand U2220 (N_2220,N_1430,N_1234);
nand U2221 (N_2221,N_1381,N_1365);
nor U2222 (N_2222,N_1484,N_1653);
or U2223 (N_2223,N_1547,N_1767);
and U2224 (N_2224,N_1248,N_1659);
and U2225 (N_2225,N_1455,N_1608);
or U2226 (N_2226,N_1695,N_1403);
or U2227 (N_2227,N_1297,N_1309);
and U2228 (N_2228,N_1782,N_1250);
nand U2229 (N_2229,N_1566,N_1470);
nor U2230 (N_2230,N_1675,N_1544);
and U2231 (N_2231,N_1672,N_1302);
and U2232 (N_2232,N_1727,N_1249);
or U2233 (N_2233,N_1645,N_1472);
nor U2234 (N_2234,N_1310,N_1737);
nor U2235 (N_2235,N_1443,N_1418);
nand U2236 (N_2236,N_1762,N_1317);
and U2237 (N_2237,N_1618,N_1289);
nand U2238 (N_2238,N_1450,N_1204);
nand U2239 (N_2239,N_1427,N_1391);
and U2240 (N_2240,N_1672,N_1612);
nor U2241 (N_2241,N_1761,N_1687);
nor U2242 (N_2242,N_1426,N_1635);
nor U2243 (N_2243,N_1529,N_1314);
or U2244 (N_2244,N_1224,N_1394);
nor U2245 (N_2245,N_1473,N_1234);
and U2246 (N_2246,N_1421,N_1283);
nand U2247 (N_2247,N_1710,N_1575);
nand U2248 (N_2248,N_1697,N_1355);
nor U2249 (N_2249,N_1320,N_1559);
nand U2250 (N_2250,N_1364,N_1200);
or U2251 (N_2251,N_1747,N_1472);
or U2252 (N_2252,N_1691,N_1551);
and U2253 (N_2253,N_1392,N_1304);
or U2254 (N_2254,N_1619,N_1655);
nand U2255 (N_2255,N_1307,N_1273);
and U2256 (N_2256,N_1587,N_1351);
and U2257 (N_2257,N_1694,N_1752);
nor U2258 (N_2258,N_1486,N_1577);
or U2259 (N_2259,N_1438,N_1242);
nor U2260 (N_2260,N_1265,N_1245);
and U2261 (N_2261,N_1269,N_1538);
nor U2262 (N_2262,N_1564,N_1782);
nand U2263 (N_2263,N_1543,N_1366);
and U2264 (N_2264,N_1243,N_1629);
or U2265 (N_2265,N_1595,N_1757);
nor U2266 (N_2266,N_1219,N_1205);
nor U2267 (N_2267,N_1495,N_1641);
xnor U2268 (N_2268,N_1578,N_1754);
nor U2269 (N_2269,N_1280,N_1322);
nor U2270 (N_2270,N_1525,N_1530);
nand U2271 (N_2271,N_1301,N_1396);
nor U2272 (N_2272,N_1376,N_1654);
nor U2273 (N_2273,N_1508,N_1245);
or U2274 (N_2274,N_1515,N_1766);
nor U2275 (N_2275,N_1552,N_1437);
xor U2276 (N_2276,N_1341,N_1321);
xnor U2277 (N_2277,N_1312,N_1433);
or U2278 (N_2278,N_1663,N_1324);
and U2279 (N_2279,N_1285,N_1433);
and U2280 (N_2280,N_1383,N_1747);
xnor U2281 (N_2281,N_1666,N_1558);
and U2282 (N_2282,N_1561,N_1579);
nand U2283 (N_2283,N_1799,N_1596);
nand U2284 (N_2284,N_1326,N_1643);
nor U2285 (N_2285,N_1578,N_1701);
nand U2286 (N_2286,N_1373,N_1272);
nor U2287 (N_2287,N_1581,N_1329);
and U2288 (N_2288,N_1601,N_1237);
and U2289 (N_2289,N_1687,N_1359);
or U2290 (N_2290,N_1507,N_1535);
and U2291 (N_2291,N_1403,N_1447);
nand U2292 (N_2292,N_1558,N_1537);
nand U2293 (N_2293,N_1544,N_1319);
or U2294 (N_2294,N_1306,N_1577);
nand U2295 (N_2295,N_1488,N_1612);
or U2296 (N_2296,N_1527,N_1690);
nand U2297 (N_2297,N_1704,N_1615);
nand U2298 (N_2298,N_1721,N_1246);
or U2299 (N_2299,N_1322,N_1370);
xor U2300 (N_2300,N_1240,N_1228);
nor U2301 (N_2301,N_1263,N_1222);
or U2302 (N_2302,N_1540,N_1329);
nand U2303 (N_2303,N_1726,N_1688);
nand U2304 (N_2304,N_1673,N_1399);
nor U2305 (N_2305,N_1744,N_1634);
or U2306 (N_2306,N_1223,N_1683);
or U2307 (N_2307,N_1202,N_1781);
nand U2308 (N_2308,N_1247,N_1373);
or U2309 (N_2309,N_1257,N_1628);
nand U2310 (N_2310,N_1638,N_1324);
or U2311 (N_2311,N_1521,N_1685);
and U2312 (N_2312,N_1629,N_1617);
or U2313 (N_2313,N_1362,N_1224);
nor U2314 (N_2314,N_1492,N_1571);
nor U2315 (N_2315,N_1741,N_1705);
or U2316 (N_2316,N_1397,N_1759);
nand U2317 (N_2317,N_1453,N_1226);
nand U2318 (N_2318,N_1332,N_1375);
nor U2319 (N_2319,N_1736,N_1313);
nor U2320 (N_2320,N_1742,N_1573);
nor U2321 (N_2321,N_1388,N_1769);
and U2322 (N_2322,N_1275,N_1289);
and U2323 (N_2323,N_1460,N_1475);
and U2324 (N_2324,N_1212,N_1299);
nor U2325 (N_2325,N_1571,N_1494);
or U2326 (N_2326,N_1409,N_1224);
nor U2327 (N_2327,N_1425,N_1628);
or U2328 (N_2328,N_1252,N_1341);
and U2329 (N_2329,N_1396,N_1626);
or U2330 (N_2330,N_1286,N_1209);
nand U2331 (N_2331,N_1484,N_1604);
xnor U2332 (N_2332,N_1750,N_1535);
nand U2333 (N_2333,N_1325,N_1680);
nor U2334 (N_2334,N_1431,N_1565);
or U2335 (N_2335,N_1777,N_1232);
xor U2336 (N_2336,N_1518,N_1555);
and U2337 (N_2337,N_1369,N_1212);
nor U2338 (N_2338,N_1765,N_1223);
and U2339 (N_2339,N_1362,N_1760);
xnor U2340 (N_2340,N_1381,N_1691);
nand U2341 (N_2341,N_1462,N_1485);
or U2342 (N_2342,N_1506,N_1328);
or U2343 (N_2343,N_1524,N_1339);
nor U2344 (N_2344,N_1303,N_1529);
or U2345 (N_2345,N_1743,N_1489);
nand U2346 (N_2346,N_1293,N_1462);
and U2347 (N_2347,N_1648,N_1681);
or U2348 (N_2348,N_1683,N_1609);
nand U2349 (N_2349,N_1242,N_1734);
nand U2350 (N_2350,N_1738,N_1276);
nor U2351 (N_2351,N_1719,N_1730);
nand U2352 (N_2352,N_1791,N_1695);
and U2353 (N_2353,N_1607,N_1430);
or U2354 (N_2354,N_1345,N_1464);
xor U2355 (N_2355,N_1365,N_1278);
and U2356 (N_2356,N_1497,N_1709);
or U2357 (N_2357,N_1701,N_1251);
nor U2358 (N_2358,N_1687,N_1631);
and U2359 (N_2359,N_1236,N_1729);
or U2360 (N_2360,N_1761,N_1629);
nand U2361 (N_2361,N_1716,N_1634);
or U2362 (N_2362,N_1364,N_1234);
nor U2363 (N_2363,N_1713,N_1645);
and U2364 (N_2364,N_1306,N_1603);
nand U2365 (N_2365,N_1570,N_1661);
and U2366 (N_2366,N_1250,N_1642);
nor U2367 (N_2367,N_1317,N_1383);
nand U2368 (N_2368,N_1299,N_1709);
nor U2369 (N_2369,N_1578,N_1739);
nor U2370 (N_2370,N_1417,N_1290);
and U2371 (N_2371,N_1372,N_1557);
and U2372 (N_2372,N_1285,N_1403);
or U2373 (N_2373,N_1437,N_1256);
or U2374 (N_2374,N_1486,N_1776);
and U2375 (N_2375,N_1202,N_1795);
nor U2376 (N_2376,N_1333,N_1253);
and U2377 (N_2377,N_1287,N_1649);
or U2378 (N_2378,N_1340,N_1516);
nand U2379 (N_2379,N_1227,N_1226);
or U2380 (N_2380,N_1385,N_1329);
and U2381 (N_2381,N_1675,N_1606);
and U2382 (N_2382,N_1306,N_1656);
nor U2383 (N_2383,N_1245,N_1336);
nor U2384 (N_2384,N_1777,N_1748);
nand U2385 (N_2385,N_1283,N_1631);
nand U2386 (N_2386,N_1529,N_1331);
nor U2387 (N_2387,N_1692,N_1707);
nand U2388 (N_2388,N_1302,N_1204);
nand U2389 (N_2389,N_1640,N_1677);
xor U2390 (N_2390,N_1561,N_1751);
or U2391 (N_2391,N_1624,N_1335);
and U2392 (N_2392,N_1793,N_1596);
and U2393 (N_2393,N_1569,N_1724);
nor U2394 (N_2394,N_1587,N_1652);
nor U2395 (N_2395,N_1749,N_1232);
and U2396 (N_2396,N_1372,N_1514);
nor U2397 (N_2397,N_1345,N_1237);
nor U2398 (N_2398,N_1319,N_1418);
and U2399 (N_2399,N_1367,N_1289);
and U2400 (N_2400,N_2356,N_2352);
or U2401 (N_2401,N_1949,N_1864);
xor U2402 (N_2402,N_1927,N_2378);
or U2403 (N_2403,N_1867,N_1852);
and U2404 (N_2404,N_2266,N_2288);
or U2405 (N_2405,N_2177,N_2327);
nor U2406 (N_2406,N_2300,N_1945);
nor U2407 (N_2407,N_2121,N_2070);
and U2408 (N_2408,N_2253,N_2375);
or U2409 (N_2409,N_2149,N_2062);
and U2410 (N_2410,N_2211,N_2204);
nand U2411 (N_2411,N_1907,N_1912);
nand U2412 (N_2412,N_2275,N_2210);
or U2413 (N_2413,N_2243,N_1800);
nand U2414 (N_2414,N_2087,N_2305);
and U2415 (N_2415,N_2311,N_2080);
and U2416 (N_2416,N_1895,N_2372);
nor U2417 (N_2417,N_2027,N_1847);
nand U2418 (N_2418,N_2169,N_2245);
nand U2419 (N_2419,N_2045,N_2010);
nor U2420 (N_2420,N_2161,N_2174);
and U2421 (N_2421,N_2159,N_2178);
or U2422 (N_2422,N_1801,N_2004);
nand U2423 (N_2423,N_1804,N_2384);
and U2424 (N_2424,N_1996,N_1951);
or U2425 (N_2425,N_2152,N_2168);
nand U2426 (N_2426,N_2196,N_1834);
and U2427 (N_2427,N_1859,N_2312);
nand U2428 (N_2428,N_2213,N_2217);
nand U2429 (N_2429,N_1906,N_2342);
and U2430 (N_2430,N_2392,N_2255);
or U2431 (N_2431,N_1981,N_2291);
or U2432 (N_2432,N_2272,N_2101);
or U2433 (N_2433,N_2322,N_2258);
and U2434 (N_2434,N_1937,N_2123);
or U2435 (N_2435,N_2247,N_2280);
nand U2436 (N_2436,N_1944,N_2308);
nor U2437 (N_2437,N_2382,N_2130);
and U2438 (N_2438,N_2381,N_2285);
nor U2439 (N_2439,N_1989,N_2398);
and U2440 (N_2440,N_2369,N_2002);
nand U2441 (N_2441,N_2205,N_2119);
nor U2442 (N_2442,N_2012,N_1980);
nor U2443 (N_2443,N_2359,N_2059);
or U2444 (N_2444,N_2343,N_1971);
and U2445 (N_2445,N_2218,N_2099);
and U2446 (N_2446,N_1810,N_2220);
or U2447 (N_2447,N_2313,N_2246);
nor U2448 (N_2448,N_1934,N_2297);
nor U2449 (N_2449,N_2110,N_2183);
nor U2450 (N_2450,N_1894,N_2223);
nand U2451 (N_2451,N_1836,N_1974);
or U2452 (N_2452,N_1809,N_2031);
nand U2453 (N_2453,N_2024,N_1930);
or U2454 (N_2454,N_2175,N_2107);
nor U2455 (N_2455,N_1883,N_2187);
nor U2456 (N_2456,N_2339,N_1808);
nand U2457 (N_2457,N_2271,N_2036);
nor U2458 (N_2458,N_1956,N_1873);
and U2459 (N_2459,N_2257,N_2154);
xor U2460 (N_2460,N_2042,N_1817);
and U2461 (N_2461,N_2287,N_2254);
and U2462 (N_2462,N_2180,N_1922);
nor U2463 (N_2463,N_2063,N_1822);
nand U2464 (N_2464,N_2048,N_2108);
nand U2465 (N_2465,N_2338,N_2188);
nor U2466 (N_2466,N_1990,N_2032);
nand U2467 (N_2467,N_2078,N_2345);
nand U2468 (N_2468,N_1841,N_1831);
nor U2469 (N_2469,N_1964,N_1874);
or U2470 (N_2470,N_2232,N_2006);
or U2471 (N_2471,N_2324,N_1878);
nand U2472 (N_2472,N_1875,N_2018);
and U2473 (N_2473,N_2035,N_2301);
nand U2474 (N_2474,N_1839,N_2349);
nand U2475 (N_2475,N_2017,N_2334);
or U2476 (N_2476,N_2380,N_2057);
nor U2477 (N_2477,N_1879,N_1943);
or U2478 (N_2478,N_2049,N_2316);
nand U2479 (N_2479,N_1925,N_2094);
nand U2480 (N_2480,N_2216,N_1899);
nand U2481 (N_2481,N_1967,N_2296);
or U2482 (N_2482,N_2114,N_1940);
nor U2483 (N_2483,N_2028,N_2084);
and U2484 (N_2484,N_2391,N_2228);
xnor U2485 (N_2485,N_2157,N_2292);
and U2486 (N_2486,N_2377,N_2109);
or U2487 (N_2487,N_1898,N_2170);
or U2488 (N_2488,N_2267,N_2111);
nand U2489 (N_2489,N_2022,N_2052);
or U2490 (N_2490,N_2385,N_1850);
or U2491 (N_2491,N_2276,N_2047);
or U2492 (N_2492,N_1938,N_2182);
and U2493 (N_2493,N_2357,N_2132);
or U2494 (N_2494,N_2089,N_2390);
and U2495 (N_2495,N_1903,N_1993);
nor U2496 (N_2496,N_1815,N_2368);
and U2497 (N_2497,N_1885,N_1916);
or U2498 (N_2498,N_2241,N_2076);
xnor U2499 (N_2499,N_1845,N_1914);
or U2500 (N_2500,N_2127,N_1881);
and U2501 (N_2501,N_1892,N_1900);
nor U2502 (N_2502,N_2172,N_1803);
or U2503 (N_2503,N_1868,N_2014);
and U2504 (N_2504,N_1921,N_1819);
xnor U2505 (N_2505,N_2103,N_2242);
nor U2506 (N_2506,N_2310,N_2184);
nand U2507 (N_2507,N_1987,N_2374);
and U2508 (N_2508,N_2299,N_2209);
nand U2509 (N_2509,N_2038,N_1977);
nor U2510 (N_2510,N_2140,N_1968);
nand U2511 (N_2511,N_2064,N_1848);
and U2512 (N_2512,N_1860,N_2284);
or U2513 (N_2513,N_2278,N_1904);
nor U2514 (N_2514,N_1941,N_2263);
and U2515 (N_2515,N_1837,N_1954);
nor U2516 (N_2516,N_1915,N_1833);
or U2517 (N_2517,N_2333,N_2155);
nand U2518 (N_2518,N_2056,N_2293);
and U2519 (N_2519,N_2237,N_1973);
nor U2520 (N_2520,N_2189,N_2354);
or U2521 (N_2521,N_1835,N_2050);
and U2522 (N_2522,N_1985,N_1863);
and U2523 (N_2523,N_2396,N_2171);
and U2524 (N_2524,N_2201,N_2091);
nor U2525 (N_2525,N_2234,N_2197);
nor U2526 (N_2526,N_1880,N_1959);
or U2527 (N_2527,N_2207,N_1812);
nand U2528 (N_2528,N_2095,N_2315);
nand U2529 (N_2529,N_2088,N_2348);
nor U2530 (N_2530,N_2306,N_2222);
nand U2531 (N_2531,N_1887,N_2071);
nand U2532 (N_2532,N_2259,N_1826);
nand U2533 (N_2533,N_2083,N_2145);
xor U2534 (N_2534,N_1935,N_1929);
nor U2535 (N_2535,N_2147,N_2033);
nor U2536 (N_2536,N_2105,N_2008);
nor U2537 (N_2537,N_2151,N_1849);
and U2538 (N_2538,N_1856,N_2126);
nor U2539 (N_2539,N_2365,N_2138);
nand U2540 (N_2540,N_1893,N_1979);
nor U2541 (N_2541,N_2336,N_2156);
nor U2542 (N_2542,N_2388,N_2116);
nand U2543 (N_2543,N_1924,N_2117);
and U2544 (N_2544,N_1830,N_2023);
and U2545 (N_2545,N_2016,N_2097);
nor U2546 (N_2546,N_1986,N_2096);
nand U2547 (N_2547,N_2055,N_1952);
or U2548 (N_2548,N_2112,N_1861);
or U2549 (N_2549,N_2081,N_2163);
or U2550 (N_2550,N_2331,N_2141);
nor U2551 (N_2551,N_2072,N_2394);
or U2552 (N_2552,N_2104,N_2212);
nor U2553 (N_2553,N_2393,N_2219);
nor U2554 (N_2554,N_2043,N_2206);
and U2555 (N_2555,N_2001,N_2137);
nor U2556 (N_2556,N_1983,N_1997);
or U2557 (N_2557,N_1872,N_1953);
nor U2558 (N_2558,N_2021,N_2165);
nand U2559 (N_2559,N_2011,N_2283);
nor U2560 (N_2560,N_2034,N_2185);
and U2561 (N_2561,N_2009,N_2135);
or U2562 (N_2562,N_2239,N_2249);
nand U2563 (N_2563,N_2061,N_2133);
or U2564 (N_2564,N_2166,N_2355);
nor U2565 (N_2565,N_1853,N_2226);
xor U2566 (N_2566,N_1939,N_1802);
nand U2567 (N_2567,N_2093,N_1829);
or U2568 (N_2568,N_2120,N_1910);
nor U2569 (N_2569,N_2317,N_2373);
nor U2570 (N_2570,N_2214,N_2221);
or U2571 (N_2571,N_1871,N_1902);
nand U2572 (N_2572,N_2361,N_2128);
nand U2573 (N_2573,N_2265,N_2250);
nor U2574 (N_2574,N_2026,N_2383);
nand U2575 (N_2575,N_1958,N_1955);
and U2576 (N_2576,N_2227,N_2321);
and U2577 (N_2577,N_1988,N_1926);
and U2578 (N_2578,N_2173,N_1960);
xnor U2579 (N_2579,N_2181,N_1840);
nand U2580 (N_2580,N_1825,N_2100);
or U2581 (N_2581,N_2019,N_2325);
or U2582 (N_2582,N_2146,N_2347);
nand U2583 (N_2583,N_2198,N_1814);
nand U2584 (N_2584,N_1947,N_2215);
nand U2585 (N_2585,N_1969,N_2134);
or U2586 (N_2586,N_2225,N_2389);
nand U2587 (N_2587,N_2039,N_2307);
nor U2588 (N_2588,N_2003,N_2252);
nor U2589 (N_2589,N_2238,N_1890);
nand U2590 (N_2590,N_1919,N_1870);
and U2591 (N_2591,N_2125,N_1909);
and U2592 (N_2592,N_2158,N_1946);
nand U2593 (N_2593,N_2203,N_2379);
xnor U2594 (N_2594,N_1984,N_2186);
nor U2595 (N_2595,N_2286,N_1928);
or U2596 (N_2596,N_2264,N_2054);
nand U2597 (N_2597,N_2060,N_2304);
xor U2598 (N_2598,N_2294,N_2085);
or U2599 (N_2599,N_1975,N_2044);
nand U2600 (N_2600,N_2150,N_1931);
nand U2601 (N_2601,N_2268,N_2199);
nor U2602 (N_2602,N_1882,N_2233);
or U2603 (N_2603,N_1972,N_1832);
nor U2604 (N_2604,N_2353,N_1978);
nand U2605 (N_2605,N_2086,N_2037);
or U2606 (N_2606,N_2191,N_1994);
or U2607 (N_2607,N_2330,N_2364);
nor U2608 (N_2608,N_2320,N_1932);
or U2609 (N_2609,N_1888,N_2256);
or U2610 (N_2610,N_1999,N_2144);
and U2611 (N_2611,N_2376,N_1820);
nor U2612 (N_2612,N_1824,N_1908);
nand U2613 (N_2613,N_2277,N_2162);
and U2614 (N_2614,N_1811,N_2013);
or U2615 (N_2615,N_1998,N_1970);
nand U2616 (N_2616,N_2098,N_2068);
nor U2617 (N_2617,N_2399,N_1862);
or U2618 (N_2618,N_2153,N_1913);
nand U2619 (N_2619,N_2073,N_2340);
nand U2620 (N_2620,N_2040,N_2350);
nand U2621 (N_2621,N_1995,N_1876);
nand U2622 (N_2622,N_2041,N_1807);
and U2623 (N_2623,N_2229,N_2351);
or U2624 (N_2624,N_2367,N_1877);
nor U2625 (N_2625,N_1851,N_1855);
nand U2626 (N_2626,N_2335,N_1948);
nor U2627 (N_2627,N_2397,N_2289);
xnor U2628 (N_2628,N_2142,N_1858);
or U2629 (N_2629,N_2136,N_2236);
or U2630 (N_2630,N_2323,N_2332);
nand U2631 (N_2631,N_2290,N_1838);
nand U2632 (N_2632,N_2069,N_2122);
nor U2633 (N_2633,N_1961,N_2139);
and U2634 (N_2634,N_2200,N_2074);
or U2635 (N_2635,N_1842,N_2118);
nand U2636 (N_2636,N_2190,N_2279);
nand U2637 (N_2637,N_2058,N_1854);
and U2638 (N_2638,N_1911,N_2160);
and U2639 (N_2639,N_2371,N_2148);
and U2640 (N_2640,N_1806,N_2230);
and U2641 (N_2641,N_2262,N_1869);
and U2642 (N_2642,N_2370,N_1966);
nand U2643 (N_2643,N_1920,N_1886);
and U2644 (N_2644,N_2176,N_1923);
nand U2645 (N_2645,N_2179,N_2143);
nand U2646 (N_2646,N_2395,N_2224);
and U2647 (N_2647,N_2235,N_2106);
and U2648 (N_2648,N_2303,N_2053);
xor U2649 (N_2649,N_2067,N_1816);
nor U2650 (N_2650,N_1897,N_2309);
or U2651 (N_2651,N_2090,N_2326);
nor U2652 (N_2652,N_2007,N_2387);
and U2653 (N_2653,N_2092,N_1992);
or U2654 (N_2654,N_2131,N_2193);
or U2655 (N_2655,N_2113,N_2281);
nor U2656 (N_2656,N_2260,N_2363);
nor U2657 (N_2657,N_2386,N_2020);
or U2658 (N_2658,N_1813,N_1818);
and U2659 (N_2659,N_2029,N_2248);
nor U2660 (N_2660,N_2282,N_1982);
or U2661 (N_2661,N_1857,N_1991);
nor U2662 (N_2662,N_2000,N_2195);
nor U2663 (N_2663,N_2251,N_2362);
nor U2664 (N_2664,N_2079,N_2025);
or U2665 (N_2665,N_2075,N_2102);
nor U2666 (N_2666,N_1821,N_2329);
and U2667 (N_2667,N_2261,N_1942);
and U2668 (N_2668,N_2366,N_1866);
nand U2669 (N_2669,N_2346,N_2065);
nor U2670 (N_2670,N_2129,N_2030);
or U2671 (N_2671,N_1933,N_2269);
nand U2672 (N_2672,N_1950,N_1884);
and U2673 (N_2673,N_2344,N_2202);
or U2674 (N_2674,N_2318,N_1962);
or U2675 (N_2675,N_2046,N_2231);
and U2676 (N_2676,N_2015,N_2124);
and U2677 (N_2677,N_1865,N_2314);
nor U2678 (N_2678,N_1889,N_1828);
or U2679 (N_2679,N_2192,N_1918);
nand U2680 (N_2680,N_1965,N_2270);
or U2681 (N_2681,N_1976,N_2358);
or U2682 (N_2682,N_2208,N_2360);
nor U2683 (N_2683,N_1843,N_2066);
nand U2684 (N_2684,N_2273,N_2295);
and U2685 (N_2685,N_1936,N_2341);
nand U2686 (N_2686,N_1891,N_1901);
or U2687 (N_2687,N_1805,N_2167);
or U2688 (N_2688,N_2115,N_2328);
nand U2689 (N_2689,N_2302,N_1905);
or U2690 (N_2690,N_2319,N_2298);
nor U2691 (N_2691,N_1957,N_2244);
and U2692 (N_2692,N_2164,N_2194);
and U2693 (N_2693,N_1963,N_2077);
nor U2694 (N_2694,N_1844,N_1846);
nand U2695 (N_2695,N_1823,N_2082);
nor U2696 (N_2696,N_2051,N_1827);
nand U2697 (N_2697,N_2274,N_2240);
or U2698 (N_2698,N_2337,N_1896);
or U2699 (N_2699,N_1917,N_2005);
or U2700 (N_2700,N_1835,N_2011);
nor U2701 (N_2701,N_1952,N_2084);
nand U2702 (N_2702,N_2126,N_2349);
or U2703 (N_2703,N_1931,N_2383);
nand U2704 (N_2704,N_1952,N_1977);
nand U2705 (N_2705,N_2324,N_2399);
or U2706 (N_2706,N_1866,N_1840);
nand U2707 (N_2707,N_1975,N_2180);
nand U2708 (N_2708,N_2029,N_2214);
and U2709 (N_2709,N_1894,N_2187);
nand U2710 (N_2710,N_2067,N_2066);
or U2711 (N_2711,N_1895,N_2363);
and U2712 (N_2712,N_1894,N_2100);
nor U2713 (N_2713,N_2123,N_2245);
nand U2714 (N_2714,N_2024,N_2122);
and U2715 (N_2715,N_1811,N_1903);
nand U2716 (N_2716,N_2282,N_2233);
nand U2717 (N_2717,N_2109,N_2153);
or U2718 (N_2718,N_1843,N_2109);
or U2719 (N_2719,N_2014,N_1916);
or U2720 (N_2720,N_2179,N_2195);
and U2721 (N_2721,N_2030,N_2062);
and U2722 (N_2722,N_1905,N_1834);
nand U2723 (N_2723,N_1883,N_1963);
nor U2724 (N_2724,N_2292,N_2135);
and U2725 (N_2725,N_1860,N_2299);
or U2726 (N_2726,N_2228,N_2393);
and U2727 (N_2727,N_1834,N_2152);
or U2728 (N_2728,N_2399,N_2172);
and U2729 (N_2729,N_1957,N_2093);
nand U2730 (N_2730,N_1911,N_2338);
and U2731 (N_2731,N_2003,N_2036);
and U2732 (N_2732,N_1933,N_2345);
and U2733 (N_2733,N_2075,N_2323);
nor U2734 (N_2734,N_1946,N_2122);
or U2735 (N_2735,N_2140,N_2172);
or U2736 (N_2736,N_1852,N_2366);
nand U2737 (N_2737,N_1920,N_1822);
and U2738 (N_2738,N_1825,N_2247);
and U2739 (N_2739,N_1859,N_2156);
and U2740 (N_2740,N_1890,N_2350);
nand U2741 (N_2741,N_2316,N_2270);
or U2742 (N_2742,N_2265,N_2114);
or U2743 (N_2743,N_1835,N_2236);
or U2744 (N_2744,N_2256,N_2208);
nand U2745 (N_2745,N_2343,N_1894);
and U2746 (N_2746,N_2137,N_2203);
nor U2747 (N_2747,N_1815,N_2209);
or U2748 (N_2748,N_2391,N_2100);
or U2749 (N_2749,N_2289,N_2312);
nor U2750 (N_2750,N_2209,N_2213);
nand U2751 (N_2751,N_2157,N_2193);
nor U2752 (N_2752,N_2050,N_1801);
or U2753 (N_2753,N_2127,N_2184);
nor U2754 (N_2754,N_2088,N_2041);
nor U2755 (N_2755,N_2033,N_2107);
nor U2756 (N_2756,N_1945,N_2268);
nand U2757 (N_2757,N_1808,N_2309);
or U2758 (N_2758,N_1909,N_2369);
or U2759 (N_2759,N_1944,N_2343);
nor U2760 (N_2760,N_1959,N_2065);
or U2761 (N_2761,N_2355,N_2159);
and U2762 (N_2762,N_1935,N_2289);
and U2763 (N_2763,N_2036,N_2287);
and U2764 (N_2764,N_2325,N_1851);
or U2765 (N_2765,N_2001,N_1952);
nand U2766 (N_2766,N_2123,N_1984);
nor U2767 (N_2767,N_2075,N_1921);
and U2768 (N_2768,N_2020,N_2011);
and U2769 (N_2769,N_2376,N_2378);
and U2770 (N_2770,N_1989,N_1956);
nor U2771 (N_2771,N_2020,N_1981);
nor U2772 (N_2772,N_2307,N_2214);
nand U2773 (N_2773,N_2050,N_2131);
nand U2774 (N_2774,N_2200,N_1814);
and U2775 (N_2775,N_2037,N_2116);
or U2776 (N_2776,N_1980,N_1957);
nand U2777 (N_2777,N_1948,N_2179);
nor U2778 (N_2778,N_2200,N_1829);
nand U2779 (N_2779,N_1858,N_2349);
and U2780 (N_2780,N_2370,N_2071);
and U2781 (N_2781,N_2329,N_2300);
and U2782 (N_2782,N_2243,N_2043);
and U2783 (N_2783,N_2353,N_2228);
nand U2784 (N_2784,N_2021,N_2115);
nor U2785 (N_2785,N_2159,N_2020);
nor U2786 (N_2786,N_2012,N_2139);
nor U2787 (N_2787,N_1954,N_1850);
or U2788 (N_2788,N_2339,N_2317);
nand U2789 (N_2789,N_2296,N_2219);
nand U2790 (N_2790,N_2094,N_2064);
nor U2791 (N_2791,N_2182,N_2307);
nand U2792 (N_2792,N_2361,N_1958);
and U2793 (N_2793,N_1950,N_2373);
and U2794 (N_2794,N_2258,N_2164);
nor U2795 (N_2795,N_1965,N_2239);
or U2796 (N_2796,N_1884,N_2145);
or U2797 (N_2797,N_1934,N_2249);
or U2798 (N_2798,N_2070,N_2375);
and U2799 (N_2799,N_1981,N_1966);
nand U2800 (N_2800,N_2279,N_1920);
nand U2801 (N_2801,N_1859,N_2287);
and U2802 (N_2802,N_1847,N_1963);
and U2803 (N_2803,N_1950,N_2016);
and U2804 (N_2804,N_1863,N_2068);
nand U2805 (N_2805,N_2105,N_2127);
and U2806 (N_2806,N_2087,N_1951);
nand U2807 (N_2807,N_2353,N_1878);
or U2808 (N_2808,N_2008,N_2261);
and U2809 (N_2809,N_2360,N_1877);
nand U2810 (N_2810,N_1982,N_2288);
nand U2811 (N_2811,N_2011,N_2062);
nor U2812 (N_2812,N_1958,N_1904);
nor U2813 (N_2813,N_1837,N_1986);
or U2814 (N_2814,N_2329,N_2084);
or U2815 (N_2815,N_2327,N_1892);
and U2816 (N_2816,N_2056,N_2127);
or U2817 (N_2817,N_2247,N_2009);
and U2818 (N_2818,N_2040,N_2076);
or U2819 (N_2819,N_2388,N_2143);
and U2820 (N_2820,N_1953,N_2254);
nor U2821 (N_2821,N_2276,N_2091);
or U2822 (N_2822,N_1947,N_2173);
and U2823 (N_2823,N_2241,N_2087);
or U2824 (N_2824,N_1990,N_2006);
nand U2825 (N_2825,N_2231,N_2286);
nand U2826 (N_2826,N_2016,N_2078);
nand U2827 (N_2827,N_2017,N_2108);
or U2828 (N_2828,N_2124,N_2086);
or U2829 (N_2829,N_2054,N_1840);
and U2830 (N_2830,N_2196,N_2358);
nor U2831 (N_2831,N_2244,N_2317);
or U2832 (N_2832,N_1855,N_2009);
nand U2833 (N_2833,N_1860,N_1824);
or U2834 (N_2834,N_2095,N_2237);
or U2835 (N_2835,N_1963,N_2273);
and U2836 (N_2836,N_2393,N_1835);
or U2837 (N_2837,N_2363,N_1992);
and U2838 (N_2838,N_2176,N_2133);
nor U2839 (N_2839,N_2304,N_2170);
nor U2840 (N_2840,N_1877,N_1953);
or U2841 (N_2841,N_2333,N_1958);
and U2842 (N_2842,N_2033,N_2358);
or U2843 (N_2843,N_1937,N_2128);
or U2844 (N_2844,N_2383,N_2170);
and U2845 (N_2845,N_2084,N_1892);
nor U2846 (N_2846,N_2101,N_2169);
or U2847 (N_2847,N_2115,N_2045);
and U2848 (N_2848,N_1997,N_2306);
nand U2849 (N_2849,N_1805,N_2158);
nor U2850 (N_2850,N_2226,N_1997);
or U2851 (N_2851,N_2365,N_1989);
or U2852 (N_2852,N_2245,N_2281);
nand U2853 (N_2853,N_2192,N_2375);
and U2854 (N_2854,N_2353,N_1895);
and U2855 (N_2855,N_2101,N_1863);
nor U2856 (N_2856,N_1955,N_2045);
or U2857 (N_2857,N_2255,N_2316);
or U2858 (N_2858,N_2025,N_2333);
nand U2859 (N_2859,N_2394,N_2052);
nor U2860 (N_2860,N_2082,N_2392);
nand U2861 (N_2861,N_2194,N_2199);
nand U2862 (N_2862,N_1956,N_2155);
nor U2863 (N_2863,N_2081,N_1949);
and U2864 (N_2864,N_2187,N_2292);
nand U2865 (N_2865,N_2120,N_2070);
or U2866 (N_2866,N_2238,N_1937);
and U2867 (N_2867,N_1996,N_2149);
nand U2868 (N_2868,N_2064,N_2136);
or U2869 (N_2869,N_2312,N_1876);
nor U2870 (N_2870,N_1899,N_2313);
nand U2871 (N_2871,N_1890,N_2305);
nor U2872 (N_2872,N_2170,N_2025);
nor U2873 (N_2873,N_1999,N_1836);
nor U2874 (N_2874,N_2081,N_2230);
or U2875 (N_2875,N_2034,N_2387);
nand U2876 (N_2876,N_2339,N_2358);
nand U2877 (N_2877,N_2241,N_2385);
nor U2878 (N_2878,N_2246,N_1909);
or U2879 (N_2879,N_2056,N_2388);
nand U2880 (N_2880,N_2097,N_1803);
nand U2881 (N_2881,N_2117,N_2048);
nor U2882 (N_2882,N_2018,N_2056);
or U2883 (N_2883,N_2093,N_2309);
or U2884 (N_2884,N_1967,N_2152);
or U2885 (N_2885,N_1813,N_2064);
or U2886 (N_2886,N_1970,N_2205);
and U2887 (N_2887,N_2156,N_2057);
and U2888 (N_2888,N_2177,N_2266);
and U2889 (N_2889,N_2053,N_1825);
or U2890 (N_2890,N_2294,N_2195);
and U2891 (N_2891,N_1914,N_2021);
and U2892 (N_2892,N_2371,N_1866);
nor U2893 (N_2893,N_2240,N_2173);
and U2894 (N_2894,N_2034,N_1822);
or U2895 (N_2895,N_2173,N_1948);
nor U2896 (N_2896,N_2071,N_1989);
nand U2897 (N_2897,N_1833,N_2222);
and U2898 (N_2898,N_1937,N_1819);
nor U2899 (N_2899,N_1977,N_2200);
and U2900 (N_2900,N_2195,N_2219);
or U2901 (N_2901,N_2369,N_1836);
or U2902 (N_2902,N_2166,N_2249);
or U2903 (N_2903,N_2158,N_2266);
nand U2904 (N_2904,N_2190,N_2040);
nand U2905 (N_2905,N_1892,N_2367);
or U2906 (N_2906,N_2107,N_2212);
and U2907 (N_2907,N_2027,N_2053);
nor U2908 (N_2908,N_1956,N_2018);
xor U2909 (N_2909,N_2061,N_2335);
nand U2910 (N_2910,N_1840,N_2358);
nand U2911 (N_2911,N_2292,N_2195);
or U2912 (N_2912,N_1950,N_2238);
nand U2913 (N_2913,N_1842,N_2373);
and U2914 (N_2914,N_1811,N_1831);
nor U2915 (N_2915,N_2196,N_2017);
or U2916 (N_2916,N_1840,N_2210);
nor U2917 (N_2917,N_2342,N_2310);
nor U2918 (N_2918,N_1853,N_2275);
nand U2919 (N_2919,N_2059,N_1955);
and U2920 (N_2920,N_1806,N_1944);
or U2921 (N_2921,N_2192,N_2143);
nand U2922 (N_2922,N_1828,N_2202);
and U2923 (N_2923,N_1845,N_1953);
and U2924 (N_2924,N_2037,N_1903);
and U2925 (N_2925,N_2265,N_2008);
or U2926 (N_2926,N_1877,N_2063);
and U2927 (N_2927,N_2285,N_2292);
or U2928 (N_2928,N_2190,N_2338);
xnor U2929 (N_2929,N_2147,N_2286);
nand U2930 (N_2930,N_1923,N_2208);
and U2931 (N_2931,N_2292,N_1811);
and U2932 (N_2932,N_2014,N_2287);
xor U2933 (N_2933,N_1930,N_1852);
and U2934 (N_2934,N_1802,N_2169);
and U2935 (N_2935,N_2178,N_1830);
nor U2936 (N_2936,N_2038,N_2215);
or U2937 (N_2937,N_1874,N_2307);
or U2938 (N_2938,N_1968,N_2206);
and U2939 (N_2939,N_2134,N_1832);
nand U2940 (N_2940,N_2049,N_2152);
nand U2941 (N_2941,N_1976,N_1831);
nor U2942 (N_2942,N_1913,N_2397);
or U2943 (N_2943,N_2104,N_2174);
and U2944 (N_2944,N_1980,N_2060);
nor U2945 (N_2945,N_2271,N_2045);
nand U2946 (N_2946,N_2118,N_2205);
nand U2947 (N_2947,N_2091,N_2373);
and U2948 (N_2948,N_1853,N_2162);
or U2949 (N_2949,N_2044,N_1885);
or U2950 (N_2950,N_2212,N_1827);
nor U2951 (N_2951,N_2048,N_1819);
or U2952 (N_2952,N_1801,N_2120);
or U2953 (N_2953,N_1996,N_1857);
xor U2954 (N_2954,N_1910,N_2301);
and U2955 (N_2955,N_2225,N_1930);
and U2956 (N_2956,N_1915,N_1878);
and U2957 (N_2957,N_2089,N_2001);
or U2958 (N_2958,N_2158,N_2108);
or U2959 (N_2959,N_1961,N_2016);
or U2960 (N_2960,N_2065,N_2319);
nand U2961 (N_2961,N_1884,N_1963);
or U2962 (N_2962,N_2032,N_2102);
xnor U2963 (N_2963,N_2391,N_2106);
and U2964 (N_2964,N_1848,N_2216);
nand U2965 (N_2965,N_2088,N_2134);
or U2966 (N_2966,N_2250,N_1814);
nand U2967 (N_2967,N_1856,N_2029);
nand U2968 (N_2968,N_2316,N_1932);
nor U2969 (N_2969,N_1899,N_2137);
nand U2970 (N_2970,N_1892,N_2054);
and U2971 (N_2971,N_2052,N_2209);
nor U2972 (N_2972,N_2018,N_2204);
or U2973 (N_2973,N_1830,N_1852);
or U2974 (N_2974,N_1935,N_2002);
and U2975 (N_2975,N_1939,N_2098);
nand U2976 (N_2976,N_2227,N_2026);
nand U2977 (N_2977,N_2140,N_1958);
and U2978 (N_2978,N_1941,N_1905);
nand U2979 (N_2979,N_2240,N_2151);
or U2980 (N_2980,N_2018,N_2038);
and U2981 (N_2981,N_2338,N_2315);
and U2982 (N_2982,N_2303,N_1838);
nor U2983 (N_2983,N_2248,N_2136);
nand U2984 (N_2984,N_1954,N_2007);
and U2985 (N_2985,N_1983,N_2080);
nor U2986 (N_2986,N_1867,N_1897);
and U2987 (N_2987,N_1996,N_1807);
and U2988 (N_2988,N_1855,N_2108);
or U2989 (N_2989,N_2251,N_2215);
or U2990 (N_2990,N_2292,N_2339);
or U2991 (N_2991,N_1812,N_1838);
nand U2992 (N_2992,N_1973,N_2279);
and U2993 (N_2993,N_2313,N_1902);
nand U2994 (N_2994,N_1878,N_2043);
and U2995 (N_2995,N_2126,N_1848);
or U2996 (N_2996,N_2083,N_2334);
nand U2997 (N_2997,N_2394,N_1905);
or U2998 (N_2998,N_1839,N_1908);
or U2999 (N_2999,N_2078,N_1917);
or UO_0 (O_0,N_2953,N_2504);
nand UO_1 (O_1,N_2692,N_2988);
nor UO_2 (O_2,N_2539,N_2864);
and UO_3 (O_3,N_2746,N_2830);
nor UO_4 (O_4,N_2532,N_2652);
or UO_5 (O_5,N_2724,N_2419);
or UO_6 (O_6,N_2883,N_2612);
or UO_7 (O_7,N_2929,N_2514);
nor UO_8 (O_8,N_2491,N_2770);
and UO_9 (O_9,N_2975,N_2817);
and UO_10 (O_10,N_2457,N_2408);
nand UO_11 (O_11,N_2730,N_2905);
nand UO_12 (O_12,N_2498,N_2586);
nand UO_13 (O_13,N_2446,N_2956);
nand UO_14 (O_14,N_2952,N_2632);
nor UO_15 (O_15,N_2540,N_2793);
nand UO_16 (O_16,N_2554,N_2927);
and UO_17 (O_17,N_2462,N_2958);
nand UO_18 (O_18,N_2932,N_2976);
nand UO_19 (O_19,N_2937,N_2996);
nand UO_20 (O_20,N_2897,N_2798);
or UO_21 (O_21,N_2574,N_2659);
and UO_22 (O_22,N_2892,N_2890);
nand UO_23 (O_23,N_2541,N_2781);
and UO_24 (O_24,N_2807,N_2486);
nand UO_25 (O_25,N_2997,N_2577);
nand UO_26 (O_26,N_2722,N_2465);
nand UO_27 (O_27,N_2573,N_2678);
nor UO_28 (O_28,N_2492,N_2410);
nor UO_29 (O_29,N_2720,N_2570);
nand UO_30 (O_30,N_2422,N_2756);
xor UO_31 (O_31,N_2585,N_2912);
nand UO_32 (O_32,N_2881,N_2971);
nor UO_33 (O_33,N_2863,N_2458);
or UO_34 (O_34,N_2903,N_2911);
nand UO_35 (O_35,N_2417,N_2780);
or UO_36 (O_36,N_2551,N_2944);
and UO_37 (O_37,N_2593,N_2868);
nand UO_38 (O_38,N_2943,N_2758);
and UO_39 (O_39,N_2950,N_2870);
and UO_40 (O_40,N_2493,N_2699);
nand UO_41 (O_41,N_2442,N_2655);
and UO_42 (O_42,N_2649,N_2978);
and UO_43 (O_43,N_2472,N_2445);
nor UO_44 (O_44,N_2487,N_2945);
nand UO_45 (O_45,N_2751,N_2764);
or UO_46 (O_46,N_2799,N_2528);
and UO_47 (O_47,N_2850,N_2977);
or UO_48 (O_48,N_2569,N_2832);
or UO_49 (O_49,N_2467,N_2902);
nand UO_50 (O_50,N_2672,N_2979);
and UO_51 (O_51,N_2477,N_2584);
and UO_52 (O_52,N_2617,N_2796);
nor UO_53 (O_53,N_2974,N_2494);
and UO_54 (O_54,N_2572,N_2925);
or UO_55 (O_55,N_2928,N_2402);
or UO_56 (O_56,N_2833,N_2682);
nor UO_57 (O_57,N_2827,N_2683);
or UO_58 (O_58,N_2431,N_2463);
or UO_59 (O_59,N_2866,N_2851);
and UO_60 (O_60,N_2450,N_2860);
and UO_61 (O_61,N_2765,N_2676);
nor UO_62 (O_62,N_2602,N_2856);
nand UO_63 (O_63,N_2846,N_2638);
and UO_64 (O_64,N_2518,N_2600);
and UO_65 (O_65,N_2835,N_2715);
nor UO_66 (O_66,N_2984,N_2665);
and UO_67 (O_67,N_2790,N_2961);
or UO_68 (O_68,N_2575,N_2875);
nor UO_69 (O_69,N_2964,N_2441);
nand UO_70 (O_70,N_2747,N_2544);
nor UO_71 (O_71,N_2814,N_2667);
nor UO_72 (O_72,N_2762,N_2871);
nand UO_73 (O_73,N_2533,N_2861);
or UO_74 (O_74,N_2635,N_2565);
and UO_75 (O_75,N_2898,N_2853);
nand UO_76 (O_76,N_2436,N_2841);
and UO_77 (O_77,N_2411,N_2429);
nor UO_78 (O_78,N_2967,N_2695);
or UO_79 (O_79,N_2962,N_2657);
and UO_80 (O_80,N_2865,N_2522);
nor UO_81 (O_81,N_2645,N_2688);
and UO_82 (O_82,N_2689,N_2412);
nor UO_83 (O_83,N_2938,N_2786);
nor UO_84 (O_84,N_2718,N_2480);
nor UO_85 (O_85,N_2433,N_2736);
nand UO_86 (O_86,N_2475,N_2435);
or UO_87 (O_87,N_2805,N_2908);
nor UO_88 (O_88,N_2685,N_2628);
and UO_89 (O_89,N_2656,N_2428);
nand UO_90 (O_90,N_2500,N_2918);
nand UO_91 (O_91,N_2413,N_2773);
and UO_92 (O_92,N_2503,N_2869);
nand UO_93 (O_93,N_2924,N_2693);
nor UO_94 (O_94,N_2557,N_2766);
and UO_95 (O_95,N_2716,N_2947);
nor UO_96 (O_96,N_2543,N_2536);
nor UO_97 (O_97,N_2739,N_2591);
or UO_98 (O_98,N_2820,N_2456);
nor UO_99 (O_99,N_2468,N_2794);
nand UO_100 (O_100,N_2440,N_2742);
nor UO_101 (O_101,N_2749,N_2893);
and UO_102 (O_102,N_2791,N_2954);
nand UO_103 (O_103,N_2671,N_2753);
and UO_104 (O_104,N_2867,N_2712);
nand UO_105 (O_105,N_2713,N_2508);
or UO_106 (O_106,N_2873,N_2401);
or UO_107 (O_107,N_2862,N_2596);
and UO_108 (O_108,N_2727,N_2914);
nand UO_109 (O_109,N_2737,N_2788);
nor UO_110 (O_110,N_2845,N_2717);
and UO_111 (O_111,N_2858,N_2641);
or UO_112 (O_112,N_2555,N_2459);
and UO_113 (O_113,N_2679,N_2530);
or UO_114 (O_114,N_2496,N_2432);
nor UO_115 (O_115,N_2831,N_2825);
nor UO_116 (O_116,N_2627,N_2703);
nor UO_117 (O_117,N_2711,N_2763);
nand UO_118 (O_118,N_2843,N_2453);
and UO_119 (O_119,N_2587,N_2815);
or UO_120 (O_120,N_2804,N_2529);
nand UO_121 (O_121,N_2681,N_2725);
and UO_122 (O_122,N_2728,N_2455);
or UO_123 (O_123,N_2647,N_2696);
or UO_124 (O_124,N_2707,N_2666);
or UO_125 (O_125,N_2754,N_2704);
or UO_126 (O_126,N_2499,N_2818);
and UO_127 (O_127,N_2660,N_2631);
or UO_128 (O_128,N_2545,N_2708);
and UO_129 (O_129,N_2603,N_2779);
or UO_130 (O_130,N_2661,N_2620);
and UO_131 (O_131,N_2792,N_2917);
nor UO_132 (O_132,N_2438,N_2669);
nand UO_133 (O_133,N_2848,N_2731);
nor UO_134 (O_134,N_2537,N_2829);
or UO_135 (O_135,N_2633,N_2414);
nor UO_136 (O_136,N_2980,N_2973);
nand UO_137 (O_137,N_2824,N_2416);
nand UO_138 (O_138,N_2723,N_2625);
nor UO_139 (O_139,N_2469,N_2624);
or UO_140 (O_140,N_2760,N_2963);
nand UO_141 (O_141,N_2513,N_2721);
or UO_142 (O_142,N_2889,N_2534);
nand UO_143 (O_143,N_2481,N_2690);
nor UO_144 (O_144,N_2615,N_2705);
nor UO_145 (O_145,N_2710,N_2839);
and UO_146 (O_146,N_2616,N_2470);
or UO_147 (O_147,N_2430,N_2443);
and UO_148 (O_148,N_2771,N_2916);
nor UO_149 (O_149,N_2854,N_2418);
and UO_150 (O_150,N_2546,N_2564);
nand UO_151 (O_151,N_2409,N_2608);
or UO_152 (O_152,N_2733,N_2806);
and UO_153 (O_153,N_2592,N_2684);
nand UO_154 (O_154,N_2582,N_2535);
nand UO_155 (O_155,N_2872,N_2994);
nor UO_156 (O_156,N_2935,N_2662);
and UO_157 (O_157,N_2567,N_2939);
nand UO_158 (O_158,N_2990,N_2901);
nand UO_159 (O_159,N_2523,N_2729);
and UO_160 (O_160,N_2895,N_2425);
or UO_161 (O_161,N_2599,N_2538);
nand UO_162 (O_162,N_2913,N_2750);
and UO_163 (O_163,N_2951,N_2969);
or UO_164 (O_164,N_2836,N_2816);
or UO_165 (O_165,N_2885,N_2650);
nand UO_166 (O_166,N_2821,N_2478);
and UO_167 (O_167,N_2857,N_2775);
or UO_168 (O_168,N_2941,N_2420);
nand UO_169 (O_169,N_2842,N_2787);
nor UO_170 (O_170,N_2965,N_2454);
nand UO_171 (O_171,N_2719,N_2489);
or UO_172 (O_172,N_2777,N_2697);
and UO_173 (O_173,N_2512,N_2561);
or UO_174 (O_174,N_2621,N_2614);
nand UO_175 (O_175,N_2785,N_2899);
or UO_176 (O_176,N_2946,N_2651);
and UO_177 (O_177,N_2542,N_2642);
nand UO_178 (O_178,N_2502,N_2910);
nand UO_179 (O_179,N_2847,N_2664);
or UO_180 (O_180,N_2801,N_2619);
nor UO_181 (O_181,N_2476,N_2844);
nor UO_182 (O_182,N_2884,N_2802);
and UO_183 (O_183,N_2516,N_2876);
nor UO_184 (O_184,N_2415,N_2404);
nand UO_185 (O_185,N_2549,N_2560);
and UO_186 (O_186,N_2734,N_2859);
nor UO_187 (O_187,N_2837,N_2485);
nand UO_188 (O_188,N_2479,N_2406);
and UO_189 (O_189,N_2982,N_2957);
and UO_190 (O_190,N_2968,N_2427);
nand UO_191 (O_191,N_2448,N_2646);
or UO_192 (O_192,N_2654,N_2797);
or UO_193 (O_193,N_2687,N_2548);
nand UO_194 (O_194,N_2515,N_2778);
and UO_195 (O_195,N_2808,N_2840);
nand UO_196 (O_196,N_2686,N_2940);
or UO_197 (O_197,N_2623,N_2767);
and UO_198 (O_198,N_2519,N_2501);
nor UO_199 (O_199,N_2789,N_2639);
and UO_200 (O_200,N_2673,N_2812);
nand UO_201 (O_201,N_2887,N_2547);
nor UO_202 (O_202,N_2464,N_2474);
nand UO_203 (O_203,N_2904,N_2849);
or UO_204 (O_204,N_2588,N_2991);
and UO_205 (O_205,N_2579,N_2714);
nor UO_206 (O_206,N_2670,N_2421);
nor UO_207 (O_207,N_2505,N_2526);
or UO_208 (O_208,N_2640,N_2674);
and UO_209 (O_209,N_2795,N_2999);
and UO_210 (O_210,N_2447,N_2838);
nand UO_211 (O_211,N_2981,N_2668);
nand UO_212 (O_212,N_2774,N_2966);
and UO_213 (O_213,N_2581,N_2611);
or UO_214 (O_214,N_2698,N_2637);
nand UO_215 (O_215,N_2738,N_2888);
or UO_216 (O_216,N_2769,N_2826);
and UO_217 (O_217,N_2878,N_2740);
nand UO_218 (O_218,N_2566,N_2748);
nor UO_219 (O_219,N_2896,N_2922);
nand UO_220 (O_220,N_2813,N_2828);
nor UO_221 (O_221,N_2834,N_2658);
and UO_222 (O_222,N_2784,N_2553);
nand UO_223 (O_223,N_2403,N_2488);
nor UO_224 (O_224,N_2634,N_2583);
or UO_225 (O_225,N_2460,N_2653);
nand UO_226 (O_226,N_2755,N_2589);
and UO_227 (O_227,N_2590,N_2506);
nor UO_228 (O_228,N_2563,N_2983);
or UO_229 (O_229,N_2772,N_2955);
nand UO_230 (O_230,N_2407,N_2992);
nand UO_231 (O_231,N_2926,N_2618);
and UO_232 (O_232,N_2644,N_2426);
nand UO_233 (O_233,N_2580,N_2894);
nand UO_234 (O_234,N_2610,N_2520);
or UO_235 (O_235,N_2909,N_2819);
nand UO_236 (O_236,N_2702,N_2521);
or UO_237 (O_237,N_2607,N_2986);
or UO_238 (O_238,N_2907,N_2597);
and UO_239 (O_239,N_2972,N_2741);
nor UO_240 (O_240,N_2768,N_2595);
or UO_241 (O_241,N_2700,N_2490);
nand UO_242 (O_242,N_2613,N_2761);
nor UO_243 (O_243,N_2510,N_2726);
nand UO_244 (O_244,N_2752,N_2423);
nand UO_245 (O_245,N_2874,N_2757);
nand UO_246 (O_246,N_2879,N_2648);
nor UO_247 (O_247,N_2483,N_2745);
or UO_248 (O_248,N_2424,N_2629);
nor UO_249 (O_249,N_2743,N_2782);
or UO_250 (O_250,N_2601,N_2552);
and UO_251 (O_251,N_2452,N_2550);
or UO_252 (O_252,N_2675,N_2562);
and UO_253 (O_253,N_2882,N_2449);
and UO_254 (O_254,N_2527,N_2594);
nor UO_255 (O_255,N_2604,N_2571);
nor UO_256 (O_256,N_2473,N_2511);
nand UO_257 (O_257,N_2663,N_2461);
nor UO_258 (O_258,N_2891,N_2437);
or UO_259 (O_259,N_2886,N_2811);
nand UO_260 (O_260,N_2985,N_2880);
or UO_261 (O_261,N_2568,N_2484);
nand UO_262 (O_262,N_2934,N_2949);
and UO_263 (O_263,N_2482,N_2556);
nand UO_264 (O_264,N_2525,N_2919);
or UO_265 (O_265,N_2524,N_2942);
or UO_266 (O_266,N_2507,N_2852);
xnor UO_267 (O_267,N_2993,N_2630);
nand UO_268 (O_268,N_2906,N_2609);
nand UO_269 (O_269,N_2987,N_2931);
or UO_270 (O_270,N_2989,N_2809);
xor UO_271 (O_271,N_2559,N_2576);
and UO_272 (O_272,N_2732,N_2694);
and UO_273 (O_273,N_2400,N_2517);
nor UO_274 (O_274,N_2677,N_2691);
nor UO_275 (O_275,N_2759,N_2606);
and UO_276 (O_276,N_2923,N_2598);
or UO_277 (O_277,N_2643,N_2405);
or UO_278 (O_278,N_2471,N_2970);
or UO_279 (O_279,N_2509,N_2466);
nand UO_280 (O_280,N_2803,N_2451);
or UO_281 (O_281,N_2776,N_2626);
or UO_282 (O_282,N_2495,N_2995);
or UO_283 (O_283,N_2915,N_2998);
and UO_284 (O_284,N_2877,N_2622);
nand UO_285 (O_285,N_2735,N_2636);
nand UO_286 (O_286,N_2709,N_2855);
and UO_287 (O_287,N_2706,N_2936);
and UO_288 (O_288,N_2822,N_2948);
or UO_289 (O_289,N_2800,N_2900);
nand UO_290 (O_290,N_2920,N_2783);
or UO_291 (O_291,N_2531,N_2744);
nor UO_292 (O_292,N_2434,N_2680);
nor UO_293 (O_293,N_2823,N_2444);
nor UO_294 (O_294,N_2578,N_2921);
or UO_295 (O_295,N_2810,N_2497);
nor UO_296 (O_296,N_2959,N_2960);
nor UO_297 (O_297,N_2439,N_2558);
or UO_298 (O_298,N_2930,N_2605);
and UO_299 (O_299,N_2701,N_2933);
nor UO_300 (O_300,N_2919,N_2713);
or UO_301 (O_301,N_2954,N_2458);
nand UO_302 (O_302,N_2757,N_2888);
nor UO_303 (O_303,N_2447,N_2953);
or UO_304 (O_304,N_2756,N_2942);
nor UO_305 (O_305,N_2919,N_2540);
or UO_306 (O_306,N_2613,N_2470);
nand UO_307 (O_307,N_2867,N_2750);
nand UO_308 (O_308,N_2508,N_2650);
nor UO_309 (O_309,N_2674,N_2993);
and UO_310 (O_310,N_2621,N_2527);
nor UO_311 (O_311,N_2725,N_2533);
nand UO_312 (O_312,N_2478,N_2481);
nand UO_313 (O_313,N_2661,N_2598);
nor UO_314 (O_314,N_2568,N_2675);
and UO_315 (O_315,N_2882,N_2677);
nand UO_316 (O_316,N_2591,N_2561);
and UO_317 (O_317,N_2844,N_2493);
nand UO_318 (O_318,N_2494,N_2920);
and UO_319 (O_319,N_2517,N_2553);
or UO_320 (O_320,N_2688,N_2834);
nand UO_321 (O_321,N_2544,N_2681);
and UO_322 (O_322,N_2872,N_2603);
nor UO_323 (O_323,N_2636,N_2519);
or UO_324 (O_324,N_2633,N_2962);
or UO_325 (O_325,N_2787,N_2873);
and UO_326 (O_326,N_2853,N_2525);
nand UO_327 (O_327,N_2567,N_2821);
and UO_328 (O_328,N_2811,N_2578);
and UO_329 (O_329,N_2753,N_2522);
nor UO_330 (O_330,N_2833,N_2903);
nand UO_331 (O_331,N_2889,N_2537);
or UO_332 (O_332,N_2500,N_2921);
and UO_333 (O_333,N_2643,N_2611);
nand UO_334 (O_334,N_2716,N_2619);
nor UO_335 (O_335,N_2813,N_2442);
or UO_336 (O_336,N_2748,N_2404);
or UO_337 (O_337,N_2997,N_2816);
and UO_338 (O_338,N_2744,N_2524);
nand UO_339 (O_339,N_2630,N_2804);
nand UO_340 (O_340,N_2776,N_2849);
and UO_341 (O_341,N_2769,N_2956);
or UO_342 (O_342,N_2717,N_2676);
and UO_343 (O_343,N_2550,N_2830);
nor UO_344 (O_344,N_2446,N_2966);
nand UO_345 (O_345,N_2546,N_2792);
nand UO_346 (O_346,N_2748,N_2926);
nand UO_347 (O_347,N_2746,N_2939);
and UO_348 (O_348,N_2442,N_2542);
nand UO_349 (O_349,N_2744,N_2532);
or UO_350 (O_350,N_2559,N_2650);
nor UO_351 (O_351,N_2583,N_2822);
and UO_352 (O_352,N_2796,N_2625);
nor UO_353 (O_353,N_2458,N_2627);
nand UO_354 (O_354,N_2718,N_2662);
nor UO_355 (O_355,N_2614,N_2583);
or UO_356 (O_356,N_2986,N_2911);
and UO_357 (O_357,N_2613,N_2592);
and UO_358 (O_358,N_2856,N_2885);
nand UO_359 (O_359,N_2715,N_2981);
or UO_360 (O_360,N_2408,N_2634);
nand UO_361 (O_361,N_2770,N_2737);
nand UO_362 (O_362,N_2903,N_2561);
or UO_363 (O_363,N_2481,N_2651);
or UO_364 (O_364,N_2679,N_2883);
and UO_365 (O_365,N_2563,N_2453);
nor UO_366 (O_366,N_2842,N_2638);
nand UO_367 (O_367,N_2953,N_2508);
or UO_368 (O_368,N_2877,N_2715);
and UO_369 (O_369,N_2550,N_2519);
or UO_370 (O_370,N_2679,N_2657);
and UO_371 (O_371,N_2489,N_2873);
nand UO_372 (O_372,N_2419,N_2856);
nor UO_373 (O_373,N_2467,N_2424);
nor UO_374 (O_374,N_2806,N_2542);
nor UO_375 (O_375,N_2504,N_2768);
nor UO_376 (O_376,N_2536,N_2528);
nand UO_377 (O_377,N_2748,N_2570);
or UO_378 (O_378,N_2404,N_2484);
and UO_379 (O_379,N_2893,N_2723);
and UO_380 (O_380,N_2427,N_2929);
nand UO_381 (O_381,N_2950,N_2660);
and UO_382 (O_382,N_2926,N_2455);
or UO_383 (O_383,N_2902,N_2918);
nor UO_384 (O_384,N_2926,N_2443);
and UO_385 (O_385,N_2720,N_2487);
or UO_386 (O_386,N_2691,N_2926);
nand UO_387 (O_387,N_2776,N_2586);
nand UO_388 (O_388,N_2595,N_2624);
xnor UO_389 (O_389,N_2980,N_2916);
and UO_390 (O_390,N_2498,N_2853);
nor UO_391 (O_391,N_2814,N_2883);
nor UO_392 (O_392,N_2850,N_2788);
nor UO_393 (O_393,N_2523,N_2935);
and UO_394 (O_394,N_2488,N_2978);
nand UO_395 (O_395,N_2576,N_2427);
or UO_396 (O_396,N_2506,N_2482);
nor UO_397 (O_397,N_2769,N_2861);
or UO_398 (O_398,N_2616,N_2678);
nor UO_399 (O_399,N_2994,N_2814);
and UO_400 (O_400,N_2747,N_2871);
nand UO_401 (O_401,N_2459,N_2674);
nand UO_402 (O_402,N_2779,N_2800);
nor UO_403 (O_403,N_2839,N_2891);
nor UO_404 (O_404,N_2650,N_2791);
nand UO_405 (O_405,N_2982,N_2689);
nand UO_406 (O_406,N_2672,N_2429);
and UO_407 (O_407,N_2810,N_2812);
or UO_408 (O_408,N_2682,N_2884);
or UO_409 (O_409,N_2987,N_2688);
or UO_410 (O_410,N_2723,N_2726);
and UO_411 (O_411,N_2755,N_2638);
nor UO_412 (O_412,N_2931,N_2502);
or UO_413 (O_413,N_2823,N_2578);
and UO_414 (O_414,N_2407,N_2820);
nor UO_415 (O_415,N_2898,N_2774);
nand UO_416 (O_416,N_2448,N_2850);
or UO_417 (O_417,N_2728,N_2893);
nor UO_418 (O_418,N_2763,N_2690);
or UO_419 (O_419,N_2514,N_2528);
nor UO_420 (O_420,N_2490,N_2540);
or UO_421 (O_421,N_2953,N_2720);
nand UO_422 (O_422,N_2644,N_2985);
nor UO_423 (O_423,N_2852,N_2465);
and UO_424 (O_424,N_2634,N_2543);
nand UO_425 (O_425,N_2927,N_2792);
and UO_426 (O_426,N_2811,N_2436);
nor UO_427 (O_427,N_2419,N_2483);
or UO_428 (O_428,N_2448,N_2956);
nand UO_429 (O_429,N_2850,N_2564);
or UO_430 (O_430,N_2421,N_2486);
nand UO_431 (O_431,N_2988,N_2843);
nand UO_432 (O_432,N_2630,N_2881);
and UO_433 (O_433,N_2760,N_2762);
and UO_434 (O_434,N_2463,N_2885);
nor UO_435 (O_435,N_2566,N_2809);
or UO_436 (O_436,N_2760,N_2502);
and UO_437 (O_437,N_2407,N_2807);
or UO_438 (O_438,N_2933,N_2586);
or UO_439 (O_439,N_2684,N_2737);
xnor UO_440 (O_440,N_2927,N_2873);
nand UO_441 (O_441,N_2496,N_2695);
and UO_442 (O_442,N_2838,N_2843);
and UO_443 (O_443,N_2493,N_2426);
nor UO_444 (O_444,N_2630,N_2667);
or UO_445 (O_445,N_2706,N_2546);
nand UO_446 (O_446,N_2706,N_2511);
or UO_447 (O_447,N_2975,N_2566);
nor UO_448 (O_448,N_2934,N_2601);
and UO_449 (O_449,N_2812,N_2626);
nor UO_450 (O_450,N_2503,N_2951);
and UO_451 (O_451,N_2471,N_2819);
and UO_452 (O_452,N_2720,N_2669);
nand UO_453 (O_453,N_2657,N_2676);
or UO_454 (O_454,N_2440,N_2567);
or UO_455 (O_455,N_2558,N_2507);
or UO_456 (O_456,N_2561,N_2692);
nor UO_457 (O_457,N_2988,N_2471);
nand UO_458 (O_458,N_2901,N_2997);
or UO_459 (O_459,N_2960,N_2837);
nand UO_460 (O_460,N_2692,N_2820);
or UO_461 (O_461,N_2439,N_2516);
and UO_462 (O_462,N_2993,N_2955);
nand UO_463 (O_463,N_2809,N_2760);
or UO_464 (O_464,N_2990,N_2648);
nor UO_465 (O_465,N_2633,N_2954);
nor UO_466 (O_466,N_2429,N_2577);
nor UO_467 (O_467,N_2528,N_2997);
or UO_468 (O_468,N_2853,N_2597);
nor UO_469 (O_469,N_2740,N_2889);
and UO_470 (O_470,N_2430,N_2425);
nor UO_471 (O_471,N_2436,N_2417);
and UO_472 (O_472,N_2457,N_2412);
nand UO_473 (O_473,N_2810,N_2965);
nand UO_474 (O_474,N_2792,N_2607);
nor UO_475 (O_475,N_2658,N_2902);
or UO_476 (O_476,N_2659,N_2423);
or UO_477 (O_477,N_2488,N_2983);
and UO_478 (O_478,N_2510,N_2807);
nand UO_479 (O_479,N_2911,N_2927);
nor UO_480 (O_480,N_2626,N_2831);
and UO_481 (O_481,N_2538,N_2764);
nand UO_482 (O_482,N_2960,N_2516);
nor UO_483 (O_483,N_2650,N_2997);
or UO_484 (O_484,N_2916,N_2524);
or UO_485 (O_485,N_2415,N_2523);
nand UO_486 (O_486,N_2411,N_2658);
nor UO_487 (O_487,N_2784,N_2548);
or UO_488 (O_488,N_2473,N_2407);
or UO_489 (O_489,N_2819,N_2720);
and UO_490 (O_490,N_2803,N_2873);
nand UO_491 (O_491,N_2821,N_2825);
and UO_492 (O_492,N_2447,N_2639);
nand UO_493 (O_493,N_2676,N_2504);
or UO_494 (O_494,N_2943,N_2542);
or UO_495 (O_495,N_2630,N_2618);
or UO_496 (O_496,N_2753,N_2625);
or UO_497 (O_497,N_2918,N_2640);
nor UO_498 (O_498,N_2731,N_2929);
and UO_499 (O_499,N_2820,N_2505);
endmodule