module basic_1500_15000_2000_15_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
or U0 (N_0,In_63,In_109);
xor U1 (N_1,In_274,In_332);
xor U2 (N_2,In_728,In_1005);
xnor U3 (N_3,In_1006,In_1036);
and U4 (N_4,In_1233,In_1290);
and U5 (N_5,In_471,In_199);
and U6 (N_6,In_758,In_921);
and U7 (N_7,In_222,In_1240);
nand U8 (N_8,In_731,In_278);
xnor U9 (N_9,In_1160,In_312);
and U10 (N_10,In_263,In_957);
xor U11 (N_11,In_407,In_719);
nand U12 (N_12,In_563,In_265);
or U13 (N_13,In_118,In_1028);
nor U14 (N_14,In_445,In_532);
nor U15 (N_15,In_754,In_1312);
or U16 (N_16,In_1490,In_1482);
or U17 (N_17,In_33,In_889);
and U18 (N_18,In_1321,In_353);
and U19 (N_19,In_865,In_805);
nand U20 (N_20,In_1298,In_1425);
and U21 (N_21,In_588,In_166);
and U22 (N_22,In_1161,In_656);
or U23 (N_23,In_469,In_1463);
nand U24 (N_24,In_857,In_1385);
xnor U25 (N_25,In_1038,In_210);
nand U26 (N_26,In_768,In_248);
nand U27 (N_27,In_365,In_846);
and U28 (N_28,In_447,In_714);
nand U29 (N_29,In_1143,In_432);
nand U30 (N_30,In_1384,In_1471);
and U31 (N_31,In_257,In_1042);
nor U32 (N_32,In_57,In_1352);
and U33 (N_33,In_1022,In_872);
nor U34 (N_34,In_1051,In_43);
and U35 (N_35,In_894,In_305);
nand U36 (N_36,In_297,In_510);
xor U37 (N_37,In_1162,In_851);
xor U38 (N_38,In_621,In_387);
xor U39 (N_39,In_1158,In_925);
xor U40 (N_40,In_80,In_249);
nand U41 (N_41,In_195,In_1242);
or U42 (N_42,In_1415,In_1202);
and U43 (N_43,In_1236,In_196);
nor U44 (N_44,In_1098,In_735);
or U45 (N_45,In_558,In_1099);
and U46 (N_46,In_1235,In_835);
xnor U47 (N_47,In_900,In_111);
and U48 (N_48,In_766,In_74);
or U49 (N_49,In_785,In_811);
xor U50 (N_50,In_726,In_1103);
nand U51 (N_51,In_647,In_600);
xor U52 (N_52,In_551,In_137);
and U53 (N_53,In_255,In_369);
or U54 (N_54,In_84,In_706);
nand U55 (N_55,In_285,In_1068);
nand U56 (N_56,In_1192,In_1000);
nor U57 (N_57,In_670,In_983);
and U58 (N_58,In_1040,In_179);
nor U59 (N_59,In_1134,In_973);
nor U60 (N_60,In_465,In_1094);
nor U61 (N_61,In_636,In_205);
or U62 (N_62,In_49,In_717);
nand U63 (N_63,In_560,In_1150);
xor U64 (N_64,In_93,In_293);
nor U65 (N_65,In_7,In_523);
xnor U66 (N_66,In_227,In_709);
xor U67 (N_67,In_832,In_1483);
xnor U68 (N_68,In_262,In_695);
or U69 (N_69,In_108,In_1306);
xor U70 (N_70,In_1464,In_1095);
xnor U71 (N_71,In_713,In_1194);
nand U72 (N_72,In_246,In_85);
nor U73 (N_73,In_1414,In_494);
and U74 (N_74,In_1374,In_1174);
or U75 (N_75,In_635,In_932);
xnor U76 (N_76,In_400,In_1112);
and U77 (N_77,In_940,In_1113);
xnor U78 (N_78,In_1353,In_742);
nor U79 (N_79,In_596,In_1327);
and U80 (N_80,In_951,In_966);
xor U81 (N_81,In_1149,In_1115);
or U82 (N_82,In_193,In_1082);
xor U83 (N_83,In_1391,In_1289);
nand U84 (N_84,In_530,In_923);
and U85 (N_85,In_73,In_421);
nand U86 (N_86,In_684,In_994);
xor U87 (N_87,In_1397,In_1087);
or U88 (N_88,In_859,In_724);
and U89 (N_89,In_1039,In_1248);
xnor U90 (N_90,In_1007,In_1027);
nand U91 (N_91,In_1424,In_1246);
nor U92 (N_92,In_942,In_5);
nor U93 (N_93,In_303,In_534);
and U94 (N_94,In_663,In_545);
nand U95 (N_95,In_94,In_1480);
nor U96 (N_96,In_504,In_393);
and U97 (N_97,In_1309,In_397);
xor U98 (N_98,In_1043,In_787);
nand U99 (N_99,In_1485,In_963);
nor U100 (N_100,In_1459,In_611);
or U101 (N_101,In_1338,In_1436);
xnor U102 (N_102,In_223,In_1423);
nand U103 (N_103,In_550,In_2);
and U104 (N_104,In_1468,In_1360);
nor U105 (N_105,In_1421,In_829);
and U106 (N_106,In_786,In_134);
or U107 (N_107,In_554,In_1448);
and U108 (N_108,In_1266,In_1379);
or U109 (N_109,In_1120,In_37);
or U110 (N_110,In_1343,In_420);
and U111 (N_111,In_398,In_653);
nand U112 (N_112,In_1227,In_949);
xnor U113 (N_113,In_1177,In_186);
or U114 (N_114,In_1016,In_759);
and U115 (N_115,In_67,In_1487);
or U116 (N_116,In_182,In_242);
xnor U117 (N_117,In_929,In_329);
or U118 (N_118,In_1450,In_893);
or U119 (N_119,In_732,In_649);
nand U120 (N_120,In_440,In_299);
xor U121 (N_121,In_956,In_816);
and U122 (N_122,In_70,In_637);
nor U123 (N_123,In_292,In_391);
nor U124 (N_124,In_273,In_1388);
nand U125 (N_125,In_56,In_824);
nor U126 (N_126,In_338,In_375);
and U127 (N_127,In_307,In_1315);
and U128 (N_128,In_1069,In_562);
or U129 (N_129,In_650,In_845);
nand U130 (N_130,In_1406,In_595);
nand U131 (N_131,In_664,In_858);
xnor U132 (N_132,In_382,In_499);
or U133 (N_133,In_773,In_22);
xor U134 (N_134,In_798,In_891);
nor U135 (N_135,In_394,In_493);
xor U136 (N_136,In_698,In_388);
xor U137 (N_137,In_568,In_623);
xnor U138 (N_138,In_95,In_1473);
nand U139 (N_139,In_1444,In_174);
or U140 (N_140,In_266,In_593);
xnor U141 (N_141,In_1109,In_642);
xor U142 (N_142,In_1294,In_789);
nand U143 (N_143,In_868,In_1079);
and U144 (N_144,In_830,In_333);
nand U145 (N_145,In_997,In_103);
nand U146 (N_146,In_537,In_898);
xnor U147 (N_147,In_996,In_1469);
xnor U148 (N_148,In_740,In_1254);
nand U149 (N_149,In_1131,In_225);
or U150 (N_150,In_372,In_213);
and U151 (N_151,In_1055,In_20);
and U152 (N_152,In_247,In_476);
and U153 (N_153,In_200,In_46);
xnor U154 (N_154,In_395,In_971);
or U155 (N_155,In_902,In_1299);
xnor U156 (N_156,In_1080,In_1142);
nand U157 (N_157,In_1489,In_498);
xor U158 (N_158,In_123,In_1437);
nand U159 (N_159,In_1071,In_122);
nand U160 (N_160,In_959,In_1435);
and U161 (N_161,In_970,In_401);
or U162 (N_162,In_426,In_1328);
nor U163 (N_163,In_437,In_771);
nand U164 (N_164,In_290,In_968);
and U165 (N_165,In_1457,In_120);
xor U166 (N_166,In_967,In_987);
nor U167 (N_167,In_1361,In_539);
or U168 (N_168,In_26,In_264);
or U169 (N_169,In_301,In_747);
nor U170 (N_170,In_1096,In_191);
or U171 (N_171,In_54,In_1214);
nand U172 (N_172,In_681,In_1191);
nor U173 (N_173,In_1408,In_442);
or U174 (N_174,In_1476,In_371);
xnor U175 (N_175,In_1456,In_1398);
nor U176 (N_176,In_876,In_1176);
nand U177 (N_177,In_567,In_89);
nand U178 (N_178,In_295,In_1380);
nor U179 (N_179,In_575,In_91);
xnor U180 (N_180,In_842,In_379);
or U181 (N_181,In_1400,In_1445);
nand U182 (N_182,In_870,In_1118);
nand U183 (N_183,In_1116,In_1337);
nand U184 (N_184,In_909,In_634);
or U185 (N_185,In_1495,In_838);
nand U186 (N_186,In_1228,In_906);
nor U187 (N_187,In_1372,In_1188);
nor U188 (N_188,In_1128,In_573);
nor U189 (N_189,In_1245,In_916);
and U190 (N_190,In_308,In_528);
or U191 (N_191,In_462,In_1264);
nor U192 (N_192,In_1198,In_1389);
nand U193 (N_193,In_1260,In_704);
nor U194 (N_194,In_507,In_1124);
nand U195 (N_195,In_1147,In_1129);
xnor U196 (N_196,In_1332,In_1104);
nand U197 (N_197,In_1063,In_1373);
or U198 (N_198,In_460,In_1224);
or U199 (N_199,In_1195,In_458);
and U200 (N_200,In_319,In_124);
xor U201 (N_201,In_1204,In_1308);
nor U202 (N_202,In_1076,In_946);
xor U203 (N_203,In_1132,In_599);
or U204 (N_204,In_705,In_677);
nor U205 (N_205,In_416,In_580);
or U206 (N_206,In_322,In_339);
xor U207 (N_207,In_1386,In_1029);
nor U208 (N_208,In_638,In_947);
or U209 (N_209,In_777,In_1170);
or U210 (N_210,In_1291,In_927);
and U211 (N_211,In_612,In_1247);
or U212 (N_212,In_513,In_1370);
nor U213 (N_213,In_406,In_418);
xnor U214 (N_214,In_1278,In_886);
and U215 (N_215,In_461,In_1037);
xnor U216 (N_216,In_151,In_1368);
nand U217 (N_217,In_161,In_1154);
and U218 (N_218,In_866,In_1359);
or U219 (N_219,In_208,In_574);
nor U220 (N_220,In_616,In_203);
nand U221 (N_221,In_904,In_107);
and U222 (N_222,In_630,In_1272);
nand U223 (N_223,In_632,In_1117);
or U224 (N_224,In_1196,In_1135);
and U225 (N_225,In_217,In_609);
nand U226 (N_226,In_473,In_302);
and U227 (N_227,In_526,In_455);
nor U228 (N_228,In_837,In_608);
nor U229 (N_229,In_129,In_1077);
nand U230 (N_230,In_1108,In_1238);
xnor U231 (N_231,In_14,In_757);
and U232 (N_232,In_597,In_1271);
or U233 (N_233,In_683,In_1419);
or U234 (N_234,In_45,In_1475);
nor U235 (N_235,In_689,In_723);
nor U236 (N_236,In_1172,In_502);
xnor U237 (N_237,In_806,In_1014);
nor U238 (N_238,In_1169,In_1255);
nand U239 (N_239,In_1031,In_390);
and U240 (N_240,In_587,In_559);
nor U241 (N_241,In_1393,In_351);
and U242 (N_242,In_1089,In_366);
xnor U243 (N_243,In_711,In_1369);
nand U244 (N_244,In_472,In_1009);
or U245 (N_245,In_581,In_481);
nor U246 (N_246,In_701,In_602);
xor U247 (N_247,In_86,In_1122);
xor U248 (N_248,In_88,In_911);
nand U249 (N_249,In_412,In_235);
nand U250 (N_250,In_75,In_189);
nor U251 (N_251,In_1025,In_1032);
or U252 (N_252,In_470,In_1030);
or U253 (N_253,In_669,In_508);
or U254 (N_254,In_306,In_665);
or U255 (N_255,In_542,In_1411);
nor U256 (N_256,In_32,In_1243);
and U257 (N_257,In_183,In_707);
or U258 (N_258,In_209,In_962);
and U259 (N_259,In_1454,In_452);
nor U260 (N_260,In_1097,In_1320);
and U261 (N_261,In_564,In_298);
and U262 (N_262,In_549,In_819);
nand U263 (N_263,In_8,In_730);
xnor U264 (N_264,In_907,In_799);
and U265 (N_265,In_19,In_1394);
or U266 (N_266,In_1253,In_121);
nand U267 (N_267,In_69,In_328);
and U268 (N_268,In_887,In_168);
nor U269 (N_269,In_782,In_1270);
and U270 (N_270,In_779,In_438);
nor U271 (N_271,In_281,In_38);
and U272 (N_272,In_590,In_1241);
or U273 (N_273,In_466,In_879);
and U274 (N_274,In_619,In_141);
nand U275 (N_275,In_501,In_1267);
nor U276 (N_276,In_659,In_566);
xor U277 (N_277,In_463,In_39);
nor U278 (N_278,In_1348,In_1447);
and U279 (N_279,In_796,In_569);
xnor U280 (N_280,In_443,In_555);
and U281 (N_281,In_678,In_1035);
or U282 (N_282,In_516,In_428);
nand U283 (N_283,In_1313,In_256);
nand U284 (N_284,In_96,In_1011);
nand U285 (N_285,In_459,In_1216);
nand U286 (N_286,In_607,In_521);
xnor U287 (N_287,In_1070,In_687);
and U288 (N_288,In_583,In_1078);
or U289 (N_289,In_1229,In_1365);
xnor U290 (N_290,In_617,In_435);
and U291 (N_291,In_601,In_354);
and U292 (N_292,In_181,In_1330);
and U293 (N_293,In_628,In_1404);
xnor U294 (N_294,In_9,In_253);
nor U295 (N_295,In_950,In_1288);
nand U296 (N_296,In_1334,In_148);
and U297 (N_297,In_1081,In_1057);
nor U298 (N_298,In_60,In_984);
and U299 (N_299,In_110,In_769);
and U300 (N_300,In_1034,In_287);
nor U301 (N_301,In_1146,In_1212);
nand U302 (N_302,In_1184,In_877);
and U303 (N_303,In_775,In_739);
or U304 (N_304,In_640,In_436);
nand U305 (N_305,In_1086,In_1206);
nor U306 (N_306,In_652,In_218);
xnor U307 (N_307,In_1467,In_1390);
nor U308 (N_308,In_980,In_972);
and U309 (N_309,In_1329,In_511);
xor U310 (N_310,In_453,In_854);
nor U311 (N_311,In_703,In_856);
nor U312 (N_312,In_874,In_82);
xor U313 (N_313,In_928,In_65);
xnor U314 (N_314,In_1497,In_1075);
and U315 (N_315,In_1017,In_645);
xor U316 (N_316,In_4,In_556);
nand U317 (N_317,In_674,In_1276);
xnor U318 (N_318,In_1127,In_198);
nor U319 (N_319,In_425,In_774);
nor U320 (N_320,In_1023,In_1366);
and U321 (N_321,In_1152,In_673);
nand U322 (N_322,In_643,In_417);
nor U323 (N_323,In_1341,In_943);
nor U324 (N_324,In_809,In_16);
and U325 (N_325,In_1455,In_1265);
and U326 (N_326,In_324,In_1324);
or U327 (N_327,In_250,In_519);
or U328 (N_328,In_871,In_87);
and U329 (N_329,In_1383,In_1351);
or U330 (N_330,In_1156,In_841);
nor U331 (N_331,In_1056,In_776);
nand U332 (N_332,In_651,In_439);
and U333 (N_333,In_176,In_1367);
nor U334 (N_334,In_800,In_988);
and U335 (N_335,In_1479,In_860);
or U336 (N_336,In_955,In_803);
or U337 (N_337,In_744,In_727);
or U338 (N_338,In_855,In_802);
xnor U339 (N_339,In_657,In_41);
and U340 (N_340,In_1470,In_1249);
nand U341 (N_341,In_982,In_1085);
nor U342 (N_342,In_1484,In_0);
and U343 (N_343,In_47,In_48);
nor U344 (N_344,In_514,In_331);
and U345 (N_345,In_78,In_990);
nand U346 (N_346,In_389,In_919);
nand U347 (N_347,In_1207,In_232);
nand U348 (N_348,In_641,In_1449);
xnor U349 (N_349,In_862,In_1439);
nor U350 (N_350,In_1049,In_500);
nor U351 (N_351,In_1432,In_1319);
xnor U352 (N_352,In_1015,In_688);
or U353 (N_353,In_127,In_505);
nor U354 (N_354,In_1178,In_1251);
nand U355 (N_355,In_304,In_679);
or U356 (N_356,In_145,In_772);
or U357 (N_357,In_102,In_1208);
and U358 (N_358,In_277,In_756);
or U359 (N_359,In_454,In_1252);
and U360 (N_360,In_146,In_781);
nor U361 (N_361,In_861,In_524);
or U362 (N_362,In_167,In_1434);
or U363 (N_363,In_1059,In_214);
nor U364 (N_364,In_363,In_1244);
nand U365 (N_365,In_487,In_1314);
nand U366 (N_366,In_912,In_1004);
nor U367 (N_367,In_880,In_90);
nor U368 (N_368,In_1125,In_1067);
nor U369 (N_369,In_844,In_964);
nor U370 (N_370,In_1494,In_1141);
xor U371 (N_371,In_527,In_553);
nor U372 (N_372,In_831,In_1024);
xor U373 (N_373,In_999,In_360);
xnor U374 (N_374,In_370,In_221);
xnor U375 (N_375,In_478,In_10);
nand U376 (N_376,In_1066,In_468);
nand U377 (N_377,In_535,In_892);
and U378 (N_378,In_1430,In_101);
nand U379 (N_379,In_267,In_503);
nor U380 (N_380,In_258,In_356);
xor U381 (N_381,In_883,In_961);
and U382 (N_382,In_488,In_1323);
xor U383 (N_383,In_344,In_840);
nand U384 (N_384,In_976,In_937);
xnor U385 (N_385,In_1452,In_1218);
nor U386 (N_386,In_197,In_444);
or U387 (N_387,In_422,In_318);
and U388 (N_388,In_1460,In_1199);
nor U389 (N_389,In_890,In_42);
nand U390 (N_390,In_310,In_910);
xor U391 (N_391,In_380,In_908);
and U392 (N_392,In_138,In_1442);
or U393 (N_393,In_169,In_1165);
or U394 (N_394,In_565,In_1402);
nor U395 (N_395,In_409,In_467);
nand U396 (N_396,In_125,In_931);
xnor U397 (N_397,In_1438,In_40);
and U398 (N_398,In_780,In_1041);
and U399 (N_399,In_1133,In_700);
xor U400 (N_400,In_483,In_449);
nor U401 (N_401,In_1416,In_130);
or U402 (N_402,In_1336,In_177);
and U403 (N_403,In_1105,In_827);
or U404 (N_404,In_606,In_1310);
xor U405 (N_405,In_1164,In_1033);
nand U406 (N_406,In_658,In_741);
xnor U407 (N_407,In_1209,In_68);
and U408 (N_408,In_92,In_315);
and U409 (N_409,In_431,In_541);
and U410 (N_410,In_598,In_251);
nand U411 (N_411,In_944,In_357);
nor U412 (N_412,In_1428,In_18);
nand U413 (N_413,In_577,In_1297);
nor U414 (N_414,In_77,In_1045);
xor U415 (N_415,In_896,In_1062);
nor U416 (N_416,In_784,In_1396);
xnor U417 (N_417,In_1285,In_475);
nor U418 (N_418,In_410,In_464);
xnor U419 (N_419,In_313,In_1155);
xnor U420 (N_420,In_1190,In_284);
and U421 (N_421,In_1481,In_810);
nor U422 (N_422,In_79,In_269);
nand U423 (N_423,In_571,In_62);
nor U424 (N_424,In_325,In_788);
or U425 (N_425,In_6,In_1325);
xor U426 (N_426,In_386,In_725);
and U427 (N_427,In_484,In_808);
and U428 (N_428,In_1026,In_254);
or U429 (N_429,In_676,In_1064);
nand U430 (N_430,In_903,In_969);
nor U431 (N_431,In_543,In_974);
and U432 (N_432,In_901,In_133);
and U433 (N_433,In_424,In_28);
nand U434 (N_434,In_1060,In_31);
xor U435 (N_435,In_506,In_381);
or U436 (N_436,In_34,In_639);
and U437 (N_437,In_343,In_812);
or U438 (N_438,In_1136,In_286);
or U439 (N_439,In_823,In_1493);
or U440 (N_440,In_104,In_114);
or U441 (N_441,In_1151,In_160);
and U442 (N_442,In_1179,In_185);
and U443 (N_443,In_456,In_1286);
xor U444 (N_444,In_1020,In_1201);
nand U445 (N_445,In_531,In_309);
nand U446 (N_446,In_522,In_288);
and U447 (N_447,In_836,In_1401);
xnor U448 (N_448,In_1111,In_586);
nor U449 (N_449,In_975,In_922);
nand U450 (N_450,In_1318,In_1061);
xor U451 (N_451,In_17,In_648);
and U452 (N_452,In_1311,In_100);
or U453 (N_453,In_515,In_1472);
nor U454 (N_454,In_1258,In_13);
nor U455 (N_455,In_1058,In_1382);
nor U456 (N_456,In_404,In_157);
nor U457 (N_457,In_825,In_59);
nor U458 (N_458,In_1292,In_1441);
and U459 (N_459,In_760,In_1403);
or U460 (N_460,In_154,In_98);
xor U461 (N_461,In_1084,In_362);
nor U462 (N_462,In_228,In_1263);
nand U463 (N_463,In_1410,In_761);
xnor U464 (N_464,In_1417,In_1126);
nand U465 (N_465,In_1200,In_405);
nand U466 (N_466,In_509,In_282);
xor U467 (N_467,In_1280,In_1203);
nor U468 (N_468,In_275,In_172);
or U469 (N_469,In_1317,In_413);
nor U470 (N_470,In_241,In_1231);
xor U471 (N_471,In_383,In_790);
nor U472 (N_472,In_938,In_396);
nand U473 (N_473,In_367,In_1250);
and U474 (N_474,In_1322,In_1102);
xnor U475 (N_475,In_584,In_132);
nor U476 (N_476,In_105,In_1210);
and U477 (N_477,In_1275,In_1364);
xnor U478 (N_478,In_589,In_1375);
nor U479 (N_479,In_536,In_765);
xor U480 (N_480,In_849,In_646);
and U481 (N_481,In_1072,In_699);
xor U482 (N_482,In_952,In_1205);
or U483 (N_483,In_668,In_520);
or U484 (N_484,In_1326,In_839);
nand U485 (N_485,In_279,In_44);
and U486 (N_486,In_149,In_119);
and U487 (N_487,In_1220,In_495);
and U488 (N_488,In_1305,In_1130);
nor U489 (N_489,In_833,In_935);
nand U490 (N_490,In_340,In_311);
xor U491 (N_491,In_1381,In_604);
nand U492 (N_492,In_797,In_863);
xnor U493 (N_493,In_231,In_491);
and U494 (N_494,In_548,In_128);
or U495 (N_495,In_1407,In_716);
or U496 (N_496,In_27,In_1046);
xnor U497 (N_497,In_660,In_1137);
and U498 (N_498,In_655,In_97);
nor U499 (N_499,In_30,In_140);
xor U500 (N_500,In_1018,In_419);
nand U501 (N_501,In_211,In_112);
and U502 (N_502,In_252,In_1239);
nor U503 (N_503,In_1427,In_1222);
nor U504 (N_504,In_159,In_675);
or U505 (N_505,In_215,In_1496);
nor U506 (N_506,In_1499,In_457);
nor U507 (N_507,In_336,In_147);
nand U508 (N_508,In_1287,In_429);
and U509 (N_509,In_995,In_1054);
or U510 (N_510,In_822,In_820);
nor U511 (N_511,In_53,In_1073);
or U512 (N_512,In_276,In_1);
nor U513 (N_513,In_546,In_1230);
nand U514 (N_514,In_913,In_1012);
xor U515 (N_515,In_807,In_1226);
and U516 (N_516,In_1123,In_1168);
nand U517 (N_517,In_627,In_733);
nor U518 (N_518,In_66,In_989);
nor U519 (N_519,In_155,In_489);
or U520 (N_520,In_1100,In_1167);
and U521 (N_521,In_355,In_55);
and U522 (N_522,In_289,In_346);
and U523 (N_523,In_1013,In_1387);
or U524 (N_524,In_72,In_603);
or U525 (N_525,In_512,In_585);
xor U526 (N_526,In_373,In_490);
nand U527 (N_527,In_605,In_486);
nand U528 (N_528,In_592,In_337);
or U529 (N_529,In_1088,In_259);
xnor U530 (N_530,In_187,In_582);
and U531 (N_531,In_126,In_1277);
xor U532 (N_532,In_618,In_933);
nor U533 (N_533,In_1295,In_818);
nor U534 (N_534,In_152,In_207);
nand U535 (N_535,In_1371,In_1092);
nand U536 (N_536,In_939,In_434);
nor U537 (N_537,In_986,In_347);
or U538 (N_538,In_117,In_992);
nand U539 (N_539,In_143,In_1217);
nor U540 (N_540,In_821,In_978);
nor U541 (N_541,In_682,In_1052);
nand U542 (N_542,In_358,In_377);
nor U543 (N_543,In_1355,In_35);
nand U544 (N_544,In_1010,In_1362);
nor U545 (N_545,In_941,In_1193);
nor U546 (N_546,In_25,In_615);
nand U547 (N_547,In_11,In_361);
or U548 (N_548,In_878,In_485);
nor U549 (N_549,In_1268,In_61);
nand U550 (N_550,In_1331,In_1185);
nor U551 (N_551,In_446,In_1296);
xor U552 (N_552,In_194,In_920);
nor U553 (N_553,In_135,In_1189);
nand U554 (N_554,In_899,In_712);
nand U555 (N_555,In_352,In_136);
xnor U556 (N_556,In_686,In_884);
nand U557 (N_557,In_1148,In_991);
nor U558 (N_558,In_778,In_690);
nand U559 (N_559,In_1157,In_1183);
xor U560 (N_560,In_864,In_1093);
or U561 (N_561,In_1140,In_794);
and U562 (N_562,In_572,In_954);
nor U563 (N_563,In_834,In_236);
nand U564 (N_564,In_1300,In_384);
nor U565 (N_565,In_153,In_321);
xor U566 (N_566,In_738,In_1376);
xor U567 (N_567,In_1458,In_1302);
or U568 (N_568,In_1350,In_58);
and U569 (N_569,In_1283,In_1259);
nand U570 (N_570,In_610,In_702);
and U571 (N_571,In_3,In_1451);
nand U572 (N_572,In_1426,In_492);
and U573 (N_573,In_271,In_694);
xnor U574 (N_574,In_317,In_1492);
xor U575 (N_575,In_629,In_561);
nor U576 (N_576,In_245,In_1119);
nor U577 (N_577,In_1465,In_1433);
and U578 (N_578,In_1139,In_239);
xnor U579 (N_579,In_1232,In_948);
and U580 (N_580,In_737,In_547);
nor U581 (N_581,In_721,In_960);
nor U582 (N_582,In_1145,In_296);
or U583 (N_583,In_764,In_1187);
nand U584 (N_584,In_106,In_165);
xor U585 (N_585,In_1443,In_1461);
xor U586 (N_586,In_631,In_654);
or U587 (N_587,In_917,In_693);
nor U588 (N_588,In_374,In_661);
nor U589 (N_589,In_238,In_848);
and U590 (N_590,In_206,In_1008);
or U591 (N_591,In_1197,In_897);
and U592 (N_592,In_692,In_614);
xnor U593 (N_593,In_753,In_1110);
and U594 (N_594,In_791,In_233);
and U595 (N_595,In_1486,In_666);
nand U596 (N_596,In_1478,In_229);
and U597 (N_597,In_544,In_83);
nor U598 (N_598,In_1159,In_1175);
nand U599 (N_599,In_345,In_1378);
and U600 (N_600,In_734,In_722);
nand U601 (N_601,In_326,In_1392);
and U602 (N_602,In_1186,In_378);
nor U603 (N_603,In_188,In_411);
nand U604 (N_604,In_552,In_915);
nand U605 (N_605,In_1262,In_482);
nor U606 (N_606,In_763,In_736);
nor U607 (N_607,In_349,In_1153);
xor U608 (N_608,In_1180,In_323);
nor U609 (N_609,In_710,In_875);
nor U610 (N_610,In_930,In_1002);
xor U611 (N_611,In_51,In_1121);
and U612 (N_612,In_570,In_1395);
nor U613 (N_613,In_691,In_1215);
or U614 (N_614,In_451,In_1412);
or U615 (N_615,In_15,In_662);
xnor U616 (N_616,In_624,In_450);
and U617 (N_617,In_219,In_767);
nand U618 (N_618,In_936,In_142);
xor U619 (N_619,In_1274,In_671);
or U620 (N_620,In_1405,In_1003);
nor U621 (N_621,In_50,In_625);
or U622 (N_622,In_116,In_1171);
or U623 (N_623,In_924,In_762);
nand U624 (N_624,In_1281,In_1347);
nand U625 (N_625,In_320,In_163);
or U626 (N_626,In_1420,In_525);
nor U627 (N_627,In_873,In_399);
nor U628 (N_628,In_1340,In_847);
and U629 (N_629,In_745,In_99);
or U630 (N_630,In_1101,In_672);
xnor U631 (N_631,In_815,In_1429);
nand U632 (N_632,In_620,In_385);
or U633 (N_633,In_1440,In_1413);
xnor U634 (N_634,In_1377,In_517);
xnor U635 (N_635,In_408,In_477);
nor U636 (N_636,In_888,In_1333);
xor U637 (N_637,In_272,In_1409);
or U638 (N_638,In_718,In_270);
nor U639 (N_639,In_12,In_1050);
xnor U640 (N_640,In_843,In_792);
or U641 (N_641,In_260,In_1474);
and U642 (N_642,In_538,In_192);
xnor U643 (N_643,In_291,In_1219);
nand U644 (N_644,In_1256,In_294);
or U645 (N_645,In_697,In_748);
and U646 (N_646,In_867,In_144);
and U647 (N_647,In_190,In_402);
nor U648 (N_648,In_918,In_1357);
and U649 (N_649,In_1431,In_178);
nor U650 (N_650,In_81,In_335);
xor U651 (N_651,In_743,In_230);
or U652 (N_652,In_204,In_1114);
or U653 (N_653,In_1106,In_885);
and U654 (N_654,In_1083,In_1363);
nand U655 (N_655,In_1303,In_1453);
nand U656 (N_656,In_23,In_364);
or U657 (N_657,In_1346,In_348);
xor U658 (N_658,In_578,In_180);
nor U659 (N_659,In_448,In_1462);
and U660 (N_660,In_430,In_21);
nand U661 (N_661,In_914,In_1354);
nor U662 (N_662,In_685,In_1349);
nor U663 (N_663,In_985,In_202);
xnor U664 (N_664,In_853,In_474);
or U665 (N_665,In_1044,In_156);
nand U666 (N_666,In_633,In_234);
or U667 (N_667,In_591,In_801);
and U668 (N_668,In_557,In_350);
or U669 (N_669,In_115,In_1399);
nor U670 (N_670,In_977,In_300);
xnor U671 (N_671,In_1021,In_1418);
nand U672 (N_672,In_175,In_814);
and U673 (N_673,In_131,In_220);
or U674 (N_674,In_330,In_403);
nand U675 (N_675,In_533,In_1335);
and U676 (N_676,In_1342,In_427);
and U677 (N_677,In_750,In_341);
nor U678 (N_678,In_1488,In_1065);
or U679 (N_679,In_993,In_644);
or U680 (N_680,In_1182,In_622);
or U681 (N_681,In_71,In_1316);
and U682 (N_682,In_1282,In_953);
nand U683 (N_683,In_905,In_24);
or U684 (N_684,In_795,In_1053);
and U685 (N_685,In_376,In_479);
and U686 (N_686,In_576,In_184);
nand U687 (N_687,In_1047,In_626);
xor U688 (N_688,In_496,In_1293);
xnor U689 (N_689,In_162,In_1358);
xor U690 (N_690,In_1498,In_334);
and U691 (N_691,In_158,In_1269);
nand U692 (N_692,In_1163,In_1138);
or U693 (N_693,In_433,In_139);
nand U694 (N_694,In_755,In_752);
and U695 (N_695,In_1339,In_613);
xnor U696 (N_696,In_1237,In_280);
nor U697 (N_697,In_881,In_783);
or U698 (N_698,In_170,In_680);
nand U699 (N_699,In_1090,In_76);
or U700 (N_700,In_850,In_1446);
xor U701 (N_701,In_1166,In_415);
and U702 (N_702,In_1344,In_1211);
and U703 (N_703,In_64,In_594);
xnor U704 (N_704,In_164,In_1307);
and U705 (N_705,In_979,In_52);
xnor U706 (N_706,In_667,In_1257);
and U707 (N_707,In_171,In_240);
and U708 (N_708,In_1304,In_715);
and U709 (N_709,In_708,In_1356);
nor U710 (N_710,In_243,In_1019);
xor U711 (N_711,In_1345,In_29);
xnor U712 (N_712,In_1466,In_1223);
nand U713 (N_713,In_958,In_212);
xor U714 (N_714,In_414,In_244);
nor U715 (N_715,In_869,In_368);
xnor U716 (N_716,In_423,In_316);
nand U717 (N_717,In_998,In_314);
nand U718 (N_718,In_1181,In_261);
and U719 (N_719,In_540,In_237);
nand U720 (N_720,In_1261,In_1284);
nand U721 (N_721,In_729,In_579);
or U722 (N_722,In_852,In_926);
nor U723 (N_723,In_1234,In_518);
nor U724 (N_724,In_173,In_746);
and U725 (N_725,In_342,In_720);
and U726 (N_726,In_224,In_770);
and U727 (N_727,In_1107,In_749);
nand U728 (N_728,In_1091,In_1001);
nor U729 (N_729,In_1273,In_201);
or U730 (N_730,In_150,In_793);
or U731 (N_731,In_1422,In_36);
or U732 (N_732,In_817,In_226);
or U733 (N_733,In_392,In_268);
xor U734 (N_734,In_1221,In_981);
and U735 (N_735,In_359,In_1491);
or U736 (N_736,In_945,In_480);
or U737 (N_737,In_804,In_1477);
or U738 (N_738,In_895,In_965);
or U739 (N_739,In_1074,In_934);
or U740 (N_740,In_327,In_813);
nand U741 (N_741,In_751,In_1213);
nor U742 (N_742,In_1279,In_1301);
xnor U743 (N_743,In_529,In_1048);
nor U744 (N_744,In_216,In_882);
or U745 (N_745,In_283,In_441);
nand U746 (N_746,In_1173,In_828);
or U747 (N_747,In_113,In_1225);
xnor U748 (N_748,In_497,In_696);
nor U749 (N_749,In_826,In_1144);
or U750 (N_750,In_769,In_594);
and U751 (N_751,In_349,In_201);
or U752 (N_752,In_7,In_55);
nand U753 (N_753,In_623,In_120);
and U754 (N_754,In_227,In_1227);
xnor U755 (N_755,In_812,In_1273);
or U756 (N_756,In_1225,In_151);
nor U757 (N_757,In_695,In_864);
nor U758 (N_758,In_1350,In_469);
xnor U759 (N_759,In_785,In_856);
nand U760 (N_760,In_281,In_957);
and U761 (N_761,In_211,In_4);
nand U762 (N_762,In_735,In_1020);
xnor U763 (N_763,In_1156,In_1352);
or U764 (N_764,In_1057,In_926);
nor U765 (N_765,In_251,In_89);
and U766 (N_766,In_1298,In_646);
xor U767 (N_767,In_1490,In_234);
nor U768 (N_768,In_1320,In_526);
or U769 (N_769,In_1091,In_1213);
or U770 (N_770,In_2,In_432);
nor U771 (N_771,In_97,In_905);
xor U772 (N_772,In_959,In_1064);
or U773 (N_773,In_1123,In_1472);
or U774 (N_774,In_87,In_1493);
xnor U775 (N_775,In_1043,In_488);
nand U776 (N_776,In_1493,In_286);
or U777 (N_777,In_638,In_756);
or U778 (N_778,In_967,In_1);
nor U779 (N_779,In_877,In_645);
nand U780 (N_780,In_565,In_1063);
or U781 (N_781,In_74,In_92);
and U782 (N_782,In_376,In_1136);
nor U783 (N_783,In_1193,In_982);
nand U784 (N_784,In_66,In_249);
or U785 (N_785,In_72,In_2);
and U786 (N_786,In_1125,In_997);
or U787 (N_787,In_1025,In_218);
xnor U788 (N_788,In_1045,In_1037);
xor U789 (N_789,In_621,In_911);
or U790 (N_790,In_929,In_412);
nor U791 (N_791,In_1032,In_747);
and U792 (N_792,In_1060,In_977);
xor U793 (N_793,In_1062,In_1271);
nand U794 (N_794,In_421,In_881);
and U795 (N_795,In_1004,In_389);
or U796 (N_796,In_1472,In_1420);
and U797 (N_797,In_840,In_1272);
or U798 (N_798,In_858,In_398);
and U799 (N_799,In_1159,In_623);
and U800 (N_800,In_1354,In_1364);
nand U801 (N_801,In_851,In_872);
nor U802 (N_802,In_1056,In_996);
nand U803 (N_803,In_399,In_1347);
nand U804 (N_804,In_1038,In_371);
nand U805 (N_805,In_952,In_815);
nor U806 (N_806,In_536,In_771);
nand U807 (N_807,In_183,In_1202);
nor U808 (N_808,In_218,In_585);
nand U809 (N_809,In_1344,In_1052);
nor U810 (N_810,In_921,In_886);
nand U811 (N_811,In_342,In_1296);
and U812 (N_812,In_966,In_865);
nand U813 (N_813,In_466,In_957);
and U814 (N_814,In_1048,In_752);
or U815 (N_815,In_147,In_1113);
and U816 (N_816,In_760,In_840);
or U817 (N_817,In_494,In_690);
nand U818 (N_818,In_1376,In_818);
xor U819 (N_819,In_370,In_482);
xor U820 (N_820,In_15,In_1190);
nor U821 (N_821,In_14,In_561);
xor U822 (N_822,In_249,In_827);
and U823 (N_823,In_642,In_818);
and U824 (N_824,In_375,In_1115);
xnor U825 (N_825,In_680,In_964);
nor U826 (N_826,In_1020,In_646);
xor U827 (N_827,In_767,In_691);
nor U828 (N_828,In_1021,In_742);
and U829 (N_829,In_654,In_357);
and U830 (N_830,In_1443,In_911);
nor U831 (N_831,In_1008,In_1027);
nand U832 (N_832,In_943,In_1448);
and U833 (N_833,In_878,In_562);
or U834 (N_834,In_1051,In_904);
nor U835 (N_835,In_384,In_301);
nand U836 (N_836,In_590,In_1410);
nor U837 (N_837,In_1426,In_454);
nor U838 (N_838,In_1317,In_348);
nand U839 (N_839,In_1020,In_1371);
or U840 (N_840,In_673,In_854);
nand U841 (N_841,In_1415,In_500);
or U842 (N_842,In_710,In_691);
nand U843 (N_843,In_508,In_359);
nand U844 (N_844,In_163,In_646);
and U845 (N_845,In_993,In_1498);
or U846 (N_846,In_359,In_1400);
nand U847 (N_847,In_750,In_134);
nor U848 (N_848,In_1253,In_1321);
nor U849 (N_849,In_799,In_283);
nor U850 (N_850,In_1112,In_940);
xnor U851 (N_851,In_778,In_1439);
xor U852 (N_852,In_1436,In_1134);
or U853 (N_853,In_1424,In_14);
nor U854 (N_854,In_1436,In_383);
nor U855 (N_855,In_891,In_1020);
nor U856 (N_856,In_867,In_515);
and U857 (N_857,In_779,In_487);
nand U858 (N_858,In_1310,In_1090);
nand U859 (N_859,In_1012,In_267);
nand U860 (N_860,In_997,In_1472);
xnor U861 (N_861,In_792,In_21);
nand U862 (N_862,In_1353,In_190);
and U863 (N_863,In_135,In_627);
or U864 (N_864,In_1022,In_616);
nor U865 (N_865,In_1432,In_778);
nand U866 (N_866,In_371,In_1118);
xor U867 (N_867,In_992,In_1049);
nand U868 (N_868,In_737,In_1259);
nor U869 (N_869,In_920,In_666);
nor U870 (N_870,In_1080,In_376);
xor U871 (N_871,In_902,In_1498);
nand U872 (N_872,In_342,In_832);
or U873 (N_873,In_110,In_1365);
and U874 (N_874,In_590,In_495);
nand U875 (N_875,In_841,In_910);
and U876 (N_876,In_1161,In_305);
and U877 (N_877,In_1140,In_251);
and U878 (N_878,In_1146,In_319);
nor U879 (N_879,In_651,In_1042);
xor U880 (N_880,In_307,In_781);
or U881 (N_881,In_1499,In_464);
xnor U882 (N_882,In_778,In_1489);
nand U883 (N_883,In_1339,In_424);
xnor U884 (N_884,In_629,In_1499);
xor U885 (N_885,In_627,In_1189);
nor U886 (N_886,In_160,In_613);
nand U887 (N_887,In_424,In_955);
xnor U888 (N_888,In_21,In_1491);
xnor U889 (N_889,In_1236,In_1226);
nand U890 (N_890,In_1304,In_1156);
nand U891 (N_891,In_1235,In_987);
nor U892 (N_892,In_474,In_248);
or U893 (N_893,In_628,In_1116);
xor U894 (N_894,In_787,In_603);
and U895 (N_895,In_1484,In_883);
or U896 (N_896,In_449,In_902);
nand U897 (N_897,In_498,In_10);
xnor U898 (N_898,In_987,In_702);
nand U899 (N_899,In_157,In_1072);
nor U900 (N_900,In_108,In_1017);
and U901 (N_901,In_308,In_1289);
nand U902 (N_902,In_104,In_1045);
or U903 (N_903,In_1051,In_778);
nand U904 (N_904,In_676,In_440);
and U905 (N_905,In_344,In_823);
and U906 (N_906,In_728,In_246);
xnor U907 (N_907,In_562,In_474);
and U908 (N_908,In_1492,In_780);
xnor U909 (N_909,In_61,In_1287);
or U910 (N_910,In_114,In_7);
nand U911 (N_911,In_1255,In_92);
and U912 (N_912,In_1074,In_154);
or U913 (N_913,In_1296,In_29);
and U914 (N_914,In_270,In_103);
nand U915 (N_915,In_513,In_175);
and U916 (N_916,In_2,In_88);
xnor U917 (N_917,In_1234,In_708);
and U918 (N_918,In_68,In_902);
or U919 (N_919,In_1105,In_580);
and U920 (N_920,In_877,In_459);
nand U921 (N_921,In_41,In_446);
and U922 (N_922,In_167,In_1487);
nor U923 (N_923,In_333,In_1071);
and U924 (N_924,In_1306,In_896);
xor U925 (N_925,In_1235,In_75);
nor U926 (N_926,In_262,In_728);
or U927 (N_927,In_1205,In_766);
nand U928 (N_928,In_832,In_628);
or U929 (N_929,In_201,In_1374);
nor U930 (N_930,In_372,In_1020);
or U931 (N_931,In_458,In_984);
nor U932 (N_932,In_69,In_803);
and U933 (N_933,In_674,In_1297);
xnor U934 (N_934,In_1161,In_436);
nand U935 (N_935,In_1161,In_52);
and U936 (N_936,In_938,In_238);
and U937 (N_937,In_457,In_1190);
or U938 (N_938,In_1246,In_243);
or U939 (N_939,In_240,In_255);
and U940 (N_940,In_1022,In_116);
nor U941 (N_941,In_679,In_31);
or U942 (N_942,In_941,In_1191);
xor U943 (N_943,In_318,In_1130);
and U944 (N_944,In_162,In_85);
xnor U945 (N_945,In_1351,In_425);
nand U946 (N_946,In_141,In_1442);
nor U947 (N_947,In_201,In_247);
or U948 (N_948,In_44,In_632);
nand U949 (N_949,In_114,In_472);
nor U950 (N_950,In_993,In_104);
or U951 (N_951,In_949,In_60);
xnor U952 (N_952,In_642,In_9);
nand U953 (N_953,In_605,In_69);
xnor U954 (N_954,In_1047,In_706);
and U955 (N_955,In_1215,In_1375);
or U956 (N_956,In_1345,In_1341);
nor U957 (N_957,In_611,In_541);
xnor U958 (N_958,In_68,In_1252);
or U959 (N_959,In_167,In_41);
and U960 (N_960,In_1234,In_1078);
nand U961 (N_961,In_1336,In_330);
and U962 (N_962,In_54,In_494);
and U963 (N_963,In_633,In_807);
nor U964 (N_964,In_759,In_177);
and U965 (N_965,In_199,In_409);
and U966 (N_966,In_246,In_173);
xnor U967 (N_967,In_1196,In_1458);
and U968 (N_968,In_408,In_1003);
or U969 (N_969,In_311,In_1035);
nand U970 (N_970,In_495,In_1197);
nor U971 (N_971,In_600,In_1181);
nor U972 (N_972,In_229,In_435);
and U973 (N_973,In_1320,In_206);
xnor U974 (N_974,In_643,In_1414);
or U975 (N_975,In_1484,In_884);
xnor U976 (N_976,In_357,In_64);
xnor U977 (N_977,In_171,In_1163);
nor U978 (N_978,In_580,In_1089);
nand U979 (N_979,In_709,In_796);
or U980 (N_980,In_169,In_1429);
xor U981 (N_981,In_1407,In_973);
xnor U982 (N_982,In_1476,In_201);
nand U983 (N_983,In_1286,In_62);
xor U984 (N_984,In_545,In_595);
or U985 (N_985,In_1465,In_936);
nor U986 (N_986,In_401,In_428);
and U987 (N_987,In_668,In_626);
xnor U988 (N_988,In_1223,In_1296);
nor U989 (N_989,In_945,In_1242);
nand U990 (N_990,In_109,In_169);
nand U991 (N_991,In_637,In_1175);
nor U992 (N_992,In_421,In_1211);
nand U993 (N_993,In_937,In_1487);
or U994 (N_994,In_531,In_1115);
xnor U995 (N_995,In_817,In_544);
nand U996 (N_996,In_754,In_1083);
or U997 (N_997,In_1121,In_219);
and U998 (N_998,In_665,In_780);
nor U999 (N_999,In_1318,In_184);
or U1000 (N_1000,N_86,N_67);
and U1001 (N_1001,N_817,N_509);
and U1002 (N_1002,N_870,N_107);
and U1003 (N_1003,N_0,N_816);
xnor U1004 (N_1004,N_951,N_595);
nor U1005 (N_1005,N_197,N_258);
nor U1006 (N_1006,N_678,N_871);
and U1007 (N_1007,N_770,N_479);
nand U1008 (N_1008,N_291,N_662);
nand U1009 (N_1009,N_126,N_933);
and U1010 (N_1010,N_369,N_720);
nand U1011 (N_1011,N_744,N_234);
or U1012 (N_1012,N_121,N_285);
or U1013 (N_1013,N_572,N_322);
xor U1014 (N_1014,N_526,N_819);
xnor U1015 (N_1015,N_616,N_801);
and U1016 (N_1016,N_552,N_294);
nand U1017 (N_1017,N_134,N_431);
or U1018 (N_1018,N_229,N_594);
and U1019 (N_1019,N_331,N_200);
nand U1020 (N_1020,N_206,N_838);
nand U1021 (N_1021,N_149,N_854);
nand U1022 (N_1022,N_123,N_209);
xor U1023 (N_1023,N_246,N_940);
nor U1024 (N_1024,N_73,N_239);
and U1025 (N_1025,N_860,N_87);
or U1026 (N_1026,N_943,N_268);
xnor U1027 (N_1027,N_625,N_670);
and U1028 (N_1028,N_58,N_252);
nor U1029 (N_1029,N_373,N_729);
nand U1030 (N_1030,N_383,N_357);
xnor U1031 (N_1031,N_936,N_654);
xnor U1032 (N_1032,N_208,N_789);
xor U1033 (N_1033,N_668,N_592);
or U1034 (N_1034,N_634,N_549);
nor U1035 (N_1035,N_599,N_261);
nor U1036 (N_1036,N_397,N_809);
or U1037 (N_1037,N_645,N_972);
nor U1038 (N_1038,N_227,N_122);
or U1039 (N_1039,N_846,N_604);
nand U1040 (N_1040,N_800,N_637);
xnor U1041 (N_1041,N_336,N_866);
nand U1042 (N_1042,N_257,N_248);
or U1043 (N_1043,N_8,N_955);
or U1044 (N_1044,N_6,N_308);
or U1045 (N_1045,N_105,N_942);
nand U1046 (N_1046,N_284,N_146);
or U1047 (N_1047,N_803,N_400);
nand U1048 (N_1048,N_694,N_213);
or U1049 (N_1049,N_57,N_938);
nor U1050 (N_1050,N_243,N_773);
xor U1051 (N_1051,N_27,N_748);
and U1052 (N_1052,N_799,N_84);
nand U1053 (N_1053,N_71,N_689);
nand U1054 (N_1054,N_108,N_33);
or U1055 (N_1055,N_872,N_858);
nand U1056 (N_1056,N_436,N_775);
nor U1057 (N_1057,N_602,N_349);
and U1058 (N_1058,N_862,N_539);
or U1059 (N_1059,N_484,N_715);
and U1060 (N_1060,N_347,N_88);
and U1061 (N_1061,N_100,N_304);
nor U1062 (N_1062,N_598,N_899);
nor U1063 (N_1063,N_719,N_51);
xor U1064 (N_1064,N_147,N_774);
and U1065 (N_1065,N_432,N_632);
or U1066 (N_1066,N_867,N_458);
xor U1067 (N_1067,N_853,N_771);
nand U1068 (N_1068,N_732,N_254);
and U1069 (N_1069,N_647,N_957);
nor U1070 (N_1070,N_89,N_808);
nor U1071 (N_1071,N_441,N_181);
xnor U1072 (N_1072,N_507,N_739);
nor U1073 (N_1073,N_319,N_993);
xor U1074 (N_1074,N_106,N_559);
nand U1075 (N_1075,N_93,N_362);
and U1076 (N_1076,N_512,N_873);
nor U1077 (N_1077,N_535,N_570);
xor U1078 (N_1078,N_198,N_511);
and U1079 (N_1079,N_671,N_672);
or U1080 (N_1080,N_863,N_387);
or U1081 (N_1081,N_528,N_309);
xnor U1082 (N_1082,N_48,N_939);
nand U1083 (N_1083,N_180,N_641);
nor U1084 (N_1084,N_714,N_405);
xnor U1085 (N_1085,N_425,N_326);
and U1086 (N_1086,N_544,N_17);
or U1087 (N_1087,N_618,N_573);
and U1088 (N_1088,N_201,N_850);
and U1089 (N_1089,N_840,N_682);
nand U1090 (N_1090,N_734,N_736);
nor U1091 (N_1091,N_302,N_231);
and U1092 (N_1092,N_138,N_548);
nand U1093 (N_1093,N_56,N_300);
xnor U1094 (N_1094,N_408,N_342);
xor U1095 (N_1095,N_669,N_474);
or U1096 (N_1096,N_157,N_905);
or U1097 (N_1097,N_576,N_313);
nand U1098 (N_1098,N_412,N_651);
or U1099 (N_1099,N_949,N_25);
or U1100 (N_1100,N_170,N_579);
or U1101 (N_1101,N_790,N_700);
nand U1102 (N_1102,N_167,N_464);
nor U1103 (N_1103,N_96,N_470);
and U1104 (N_1104,N_880,N_364);
nor U1105 (N_1105,N_50,N_990);
nand U1106 (N_1106,N_203,N_150);
nor U1107 (N_1107,N_148,N_883);
nor U1108 (N_1108,N_821,N_179);
nor U1109 (N_1109,N_416,N_31);
nand U1110 (N_1110,N_53,N_115);
or U1111 (N_1111,N_385,N_659);
nor U1112 (N_1112,N_447,N_786);
xnor U1113 (N_1113,N_414,N_434);
or U1114 (N_1114,N_966,N_660);
or U1115 (N_1115,N_60,N_19);
nor U1116 (N_1116,N_785,N_494);
and U1117 (N_1117,N_463,N_462);
nor U1118 (N_1118,N_588,N_529);
and U1119 (N_1119,N_542,N_473);
and U1120 (N_1120,N_295,N_63);
or U1121 (N_1121,N_376,N_3);
and U1122 (N_1122,N_155,N_151);
nand U1123 (N_1123,N_45,N_532);
nand U1124 (N_1124,N_15,N_610);
nand U1125 (N_1125,N_379,N_389);
nor U1126 (N_1126,N_363,N_12);
or U1127 (N_1127,N_190,N_965);
xnor U1128 (N_1128,N_834,N_657);
nor U1129 (N_1129,N_489,N_236);
or U1130 (N_1130,N_292,N_563);
nor U1131 (N_1131,N_941,N_353);
xor U1132 (N_1132,N_102,N_128);
nor U1133 (N_1133,N_574,N_249);
xnor U1134 (N_1134,N_903,N_611);
or U1135 (N_1135,N_718,N_601);
nand U1136 (N_1136,N_454,N_184);
or U1137 (N_1137,N_293,N_169);
or U1138 (N_1138,N_445,N_350);
nand U1139 (N_1139,N_520,N_37);
xor U1140 (N_1140,N_455,N_320);
nor U1141 (N_1141,N_346,N_724);
nand U1142 (N_1142,N_956,N_478);
nand U1143 (N_1143,N_869,N_255);
nand U1144 (N_1144,N_130,N_538);
or U1145 (N_1145,N_891,N_504);
or U1146 (N_1146,N_806,N_653);
or U1147 (N_1147,N_335,N_501);
xor U1148 (N_1148,N_828,N_44);
or U1149 (N_1149,N_496,N_558);
nor U1150 (N_1150,N_276,N_66);
nor U1151 (N_1151,N_42,N_182);
nor U1152 (N_1152,N_219,N_564);
nor U1153 (N_1153,N_525,N_856);
nor U1154 (N_1154,N_352,N_900);
nand U1155 (N_1155,N_833,N_339);
xnor U1156 (N_1156,N_843,N_764);
and U1157 (N_1157,N_704,N_418);
and U1158 (N_1158,N_986,N_907);
or U1159 (N_1159,N_829,N_673);
xnor U1160 (N_1160,N_827,N_620);
and U1161 (N_1161,N_995,N_597);
nor U1162 (N_1162,N_204,N_792);
nor U1163 (N_1163,N_983,N_580);
xor U1164 (N_1164,N_288,N_70);
xor U1165 (N_1165,N_554,N_581);
and U1166 (N_1166,N_269,N_119);
nor U1167 (N_1167,N_699,N_712);
nor U1168 (N_1168,N_368,N_530);
nor U1169 (N_1169,N_422,N_609);
and U1170 (N_1170,N_240,N_237);
nand U1171 (N_1171,N_807,N_59);
or U1172 (N_1172,N_10,N_902);
nor U1173 (N_1173,N_894,N_475);
and U1174 (N_1174,N_482,N_571);
or U1175 (N_1175,N_901,N_186);
nand U1176 (N_1176,N_329,N_868);
or U1177 (N_1177,N_981,N_575);
nand U1178 (N_1178,N_21,N_438);
or U1179 (N_1179,N_35,N_7);
nand U1180 (N_1180,N_685,N_747);
nor U1181 (N_1181,N_547,N_264);
xnor U1182 (N_1182,N_18,N_259);
or U1183 (N_1183,N_781,N_131);
and U1184 (N_1184,N_517,N_429);
and U1185 (N_1185,N_915,N_946);
nand U1186 (N_1186,N_354,N_160);
nand U1187 (N_1187,N_413,N_677);
nand U1188 (N_1188,N_199,N_793);
nor U1189 (N_1189,N_844,N_521);
xnor U1190 (N_1190,N_24,N_876);
or U1191 (N_1191,N_428,N_218);
or U1192 (N_1192,N_553,N_804);
nand U1193 (N_1193,N_629,N_881);
xnor U1194 (N_1194,N_557,N_693);
xnor U1195 (N_1195,N_82,N_877);
or U1196 (N_1196,N_394,N_228);
and U1197 (N_1197,N_984,N_443);
nand U1198 (N_1198,N_191,N_896);
nand U1199 (N_1199,N_381,N_759);
nand U1200 (N_1200,N_226,N_371);
nand U1201 (N_1201,N_265,N_608);
nor U1202 (N_1202,N_29,N_433);
nor U1203 (N_1203,N_77,N_934);
nand U1204 (N_1204,N_664,N_442);
and U1205 (N_1205,N_382,N_527);
nand U1206 (N_1206,N_717,N_196);
nand U1207 (N_1207,N_307,N_540);
and U1208 (N_1208,N_918,N_534);
nand U1209 (N_1209,N_481,N_613);
xnor U1210 (N_1210,N_120,N_224);
xor U1211 (N_1211,N_762,N_892);
nor U1212 (N_1212,N_585,N_314);
nor U1213 (N_1213,N_374,N_317);
xnor U1214 (N_1214,N_702,N_423);
nand U1215 (N_1215,N_855,N_923);
nand U1216 (N_1216,N_235,N_193);
nor U1217 (N_1217,N_378,N_992);
and U1218 (N_1218,N_913,N_999);
or U1219 (N_1219,N_603,N_779);
nor U1220 (N_1220,N_953,N_878);
and U1221 (N_1221,N_419,N_95);
nand U1222 (N_1222,N_639,N_908);
and U1223 (N_1223,N_4,N_777);
xor U1224 (N_1224,N_667,N_20);
nor U1225 (N_1225,N_46,N_695);
nand U1226 (N_1226,N_958,N_546);
and U1227 (N_1227,N_752,N_755);
nor U1228 (N_1228,N_968,N_109);
nand U1229 (N_1229,N_256,N_973);
or U1230 (N_1230,N_403,N_780);
nor U1231 (N_1231,N_158,N_471);
nor U1232 (N_1232,N_679,N_343);
or U1233 (N_1233,N_805,N_731);
nand U1234 (N_1234,N_410,N_830);
or U1235 (N_1235,N_175,N_340);
and U1236 (N_1236,N_624,N_137);
and U1237 (N_1237,N_117,N_426);
nor U1238 (N_1238,N_141,N_277);
nor U1239 (N_1239,N_404,N_101);
or U1240 (N_1240,N_366,N_430);
xnor U1241 (N_1241,N_143,N_22);
and U1242 (N_1242,N_345,N_728);
and U1243 (N_1243,N_997,N_696);
nand U1244 (N_1244,N_152,N_519);
xnor U1245 (N_1245,N_708,N_270);
xnor U1246 (N_1246,N_756,N_114);
and U1247 (N_1247,N_132,N_959);
or U1248 (N_1248,N_851,N_566);
and U1249 (N_1249,N_306,N_393);
or U1250 (N_1250,N_524,N_650);
nand U1251 (N_1251,N_578,N_245);
xnor U1252 (N_1252,N_145,N_503);
and U1253 (N_1253,N_43,N_283);
or U1254 (N_1254,N_163,N_716);
xor U1255 (N_1255,N_112,N_605);
and U1256 (N_1256,N_638,N_927);
or U1257 (N_1257,N_621,N_859);
nand U1258 (N_1258,N_411,N_750);
xor U1259 (N_1259,N_788,N_187);
nor U1260 (N_1260,N_861,N_351);
xnor U1261 (N_1261,N_543,N_92);
and U1262 (N_1262,N_13,N_505);
xor U1263 (N_1263,N_2,N_769);
xnor U1264 (N_1264,N_926,N_882);
nand U1265 (N_1265,N_982,N_826);
and U1266 (N_1266,N_241,N_476);
or U1267 (N_1267,N_697,N_701);
xnor U1268 (N_1268,N_726,N_440);
xnor U1269 (N_1269,N_401,N_221);
nand U1270 (N_1270,N_640,N_344);
nand U1271 (N_1271,N_166,N_684);
xor U1272 (N_1272,N_78,N_280);
nand U1273 (N_1273,N_407,N_811);
or U1274 (N_1274,N_970,N_483);
xor U1275 (N_1275,N_439,N_296);
nor U1276 (N_1276,N_636,N_94);
nand U1277 (N_1277,N_301,N_386);
and U1278 (N_1278,N_656,N_189);
nor U1279 (N_1279,N_622,N_133);
nor U1280 (N_1280,N_948,N_852);
nand U1281 (N_1281,N_874,N_745);
nand U1282 (N_1282,N_207,N_361);
xor U1283 (N_1283,N_490,N_848);
nor U1284 (N_1284,N_266,N_456);
nor U1285 (N_1285,N_633,N_692);
xnor U1286 (N_1286,N_758,N_584);
or U1287 (N_1287,N_560,N_623);
xor U1288 (N_1288,N_398,N_614);
nor U1289 (N_1289,N_791,N_960);
or U1290 (N_1290,N_568,N_772);
nand U1291 (N_1291,N_453,N_355);
or U1292 (N_1292,N_583,N_74);
nand U1293 (N_1293,N_250,N_707);
nor U1294 (N_1294,N_127,N_330);
or U1295 (N_1295,N_281,N_154);
xor U1296 (N_1296,N_205,N_705);
or U1297 (N_1297,N_783,N_740);
nor U1298 (N_1298,N_837,N_34);
and U1299 (N_1299,N_904,N_690);
xor U1300 (N_1300,N_761,N_922);
nor U1301 (N_1301,N_536,N_81);
nor U1302 (N_1302,N_402,N_920);
xnor U1303 (N_1303,N_537,N_487);
and U1304 (N_1304,N_615,N_49);
and U1305 (N_1305,N_924,N_606);
nor U1306 (N_1306,N_845,N_5);
and U1307 (N_1307,N_810,N_502);
nand U1308 (N_1308,N_327,N_681);
xnor U1309 (N_1309,N_287,N_332);
nor U1310 (N_1310,N_988,N_865);
nor U1311 (N_1311,N_38,N_969);
and U1312 (N_1312,N_778,N_192);
nor U1313 (N_1313,N_477,N_749);
and U1314 (N_1314,N_514,N_299);
nor U1315 (N_1315,N_162,N_721);
and U1316 (N_1316,N_360,N_271);
nand U1317 (N_1317,N_887,N_643);
xor U1318 (N_1318,N_153,N_935);
or U1319 (N_1319,N_90,N_399);
xnor U1320 (N_1320,N_97,N_743);
xor U1321 (N_1321,N_674,N_80);
nor U1322 (N_1322,N_273,N_663);
xnor U1323 (N_1323,N_488,N_75);
xnor U1324 (N_1324,N_565,N_760);
xnor U1325 (N_1325,N_784,N_52);
or U1326 (N_1326,N_897,N_522);
and U1327 (N_1327,N_472,N_99);
and U1328 (N_1328,N_825,N_135);
or U1329 (N_1329,N_310,N_164);
nor U1330 (N_1330,N_321,N_680);
xnor U1331 (N_1331,N_14,N_54);
and U1332 (N_1332,N_289,N_55);
and U1333 (N_1333,N_358,N_303);
and U1334 (N_1334,N_28,N_977);
or U1335 (N_1335,N_195,N_136);
nand U1336 (N_1336,N_395,N_311);
nor U1337 (N_1337,N_885,N_921);
nand U1338 (N_1338,N_61,N_964);
or U1339 (N_1339,N_686,N_963);
or U1340 (N_1340,N_824,N_884);
nor U1341 (N_1341,N_916,N_427);
and U1342 (N_1342,N_589,N_417);
nand U1343 (N_1343,N_409,N_593);
and U1344 (N_1344,N_766,N_518);
xnor U1345 (N_1345,N_646,N_836);
nor U1346 (N_1346,N_129,N_485);
xnor U1347 (N_1347,N_550,N_415);
nand U1348 (N_1348,N_79,N_142);
nand U1349 (N_1349,N_642,N_178);
and U1350 (N_1350,N_962,N_971);
xnor U1351 (N_1351,N_676,N_356);
or U1352 (N_1352,N_709,N_323);
or U1353 (N_1353,N_183,N_710);
or U1354 (N_1354,N_467,N_776);
and U1355 (N_1355,N_11,N_286);
nand U1356 (N_1356,N_723,N_556);
nand U1357 (N_1357,N_895,N_380);
or U1358 (N_1358,N_104,N_391);
nor U1359 (N_1359,N_813,N_569);
and U1360 (N_1360,N_909,N_174);
nor U1361 (N_1361,N_247,N_794);
nor U1362 (N_1362,N_531,N_435);
nor U1363 (N_1363,N_334,N_365);
nor U1364 (N_1364,N_220,N_797);
and U1365 (N_1365,N_480,N_279);
nand U1366 (N_1366,N_666,N_91);
and U1367 (N_1367,N_64,N_274);
nor U1368 (N_1368,N_98,N_493);
nor U1369 (N_1369,N_630,N_945);
or U1370 (N_1370,N_26,N_110);
and U1371 (N_1371,N_460,N_815);
xor U1372 (N_1372,N_161,N_928);
nor U1373 (N_1373,N_424,N_910);
and U1374 (N_1374,N_139,N_980);
xor U1375 (N_1375,N_188,N_486);
xnor U1376 (N_1376,N_113,N_492);
and U1377 (N_1377,N_388,N_911);
or U1378 (N_1378,N_39,N_567);
and U1379 (N_1379,N_944,N_545);
or U1380 (N_1380,N_312,N_782);
nand U1381 (N_1381,N_491,N_727);
nand U1382 (N_1382,N_16,N_738);
nor U1383 (N_1383,N_998,N_751);
nor U1384 (N_1384,N_683,N_979);
nand U1385 (N_1385,N_889,N_994);
or U1386 (N_1386,N_577,N_172);
and U1387 (N_1387,N_437,N_847);
nand U1388 (N_1388,N_406,N_802);
and U1389 (N_1389,N_555,N_763);
or U1390 (N_1390,N_318,N_886);
xnor U1391 (N_1391,N_30,N_967);
nor U1392 (N_1392,N_420,N_253);
nand U1393 (N_1393,N_814,N_341);
or U1394 (N_1394,N_665,N_996);
nor U1395 (N_1395,N_823,N_40);
or U1396 (N_1396,N_165,N_297);
or U1397 (N_1397,N_703,N_144);
and U1398 (N_1398,N_32,N_421);
nor U1399 (N_1399,N_839,N_465);
nand U1400 (N_1400,N_298,N_932);
and U1401 (N_1401,N_925,N_251);
xor U1402 (N_1402,N_211,N_742);
nand U1403 (N_1403,N_469,N_590);
xor U1404 (N_1404,N_324,N_171);
or U1405 (N_1405,N_831,N_607);
or U1406 (N_1406,N_372,N_735);
and U1407 (N_1407,N_582,N_515);
xnor U1408 (N_1408,N_290,N_978);
nand U1409 (N_1409,N_62,N_591);
xnor U1410 (N_1410,N_85,N_516);
or U1411 (N_1411,N_818,N_627);
nand U1412 (N_1412,N_628,N_626);
nor U1413 (N_1413,N_23,N_631);
and U1414 (N_1414,N_111,N_466);
and U1415 (N_1415,N_975,N_675);
and U1416 (N_1416,N_72,N_232);
nand U1417 (N_1417,N_370,N_41);
xor U1418 (N_1418,N_698,N_533);
xor U1419 (N_1419,N_244,N_338);
nand U1420 (N_1420,N_730,N_711);
nor U1421 (N_1421,N_337,N_468);
and U1422 (N_1422,N_961,N_500);
nor U1423 (N_1423,N_929,N_596);
nor U1424 (N_1424,N_210,N_262);
and U1425 (N_1425,N_587,N_194);
nand U1426 (N_1426,N_217,N_156);
and U1427 (N_1427,N_691,N_68);
xor U1428 (N_1428,N_315,N_612);
nand U1429 (N_1429,N_448,N_375);
or U1430 (N_1430,N_185,N_450);
nor U1431 (N_1431,N_176,N_333);
and U1432 (N_1432,N_523,N_931);
nand U1433 (N_1433,N_498,N_222);
or U1434 (N_1434,N_457,N_214);
or U1435 (N_1435,N_648,N_275);
nand U1436 (N_1436,N_919,N_842);
and U1437 (N_1437,N_746,N_733);
nand U1438 (N_1438,N_917,N_173);
nor U1439 (N_1439,N_974,N_688);
and U1440 (N_1440,N_83,N_952);
xnor U1441 (N_1441,N_849,N_223);
xnor U1442 (N_1442,N_649,N_449);
xor U1443 (N_1443,N_989,N_741);
and U1444 (N_1444,N_890,N_812);
or U1445 (N_1445,N_652,N_562);
or U1446 (N_1446,N_822,N_272);
nand U1447 (N_1447,N_754,N_864);
nand U1448 (N_1448,N_737,N_1);
xnor U1449 (N_1449,N_875,N_658);
and U1450 (N_1450,N_795,N_392);
and U1451 (N_1451,N_377,N_768);
xnor U1452 (N_1452,N_36,N_459);
or U1453 (N_1453,N_359,N_497);
nand U1454 (N_1454,N_820,N_233);
nand U1455 (N_1455,N_396,N_225);
or U1456 (N_1456,N_499,N_796);
nor U1457 (N_1457,N_987,N_367);
xor U1458 (N_1458,N_937,N_260);
and U1459 (N_1459,N_140,N_888);
nor U1460 (N_1460,N_976,N_510);
nor U1461 (N_1461,N_947,N_103);
xnor U1462 (N_1462,N_841,N_898);
nand U1463 (N_1463,N_159,N_787);
and U1464 (N_1464,N_390,N_446);
and U1465 (N_1465,N_316,N_586);
nand U1466 (N_1466,N_541,N_461);
and U1467 (N_1467,N_384,N_212);
xnor U1468 (N_1468,N_69,N_617);
or U1469 (N_1469,N_267,N_495);
nor U1470 (N_1470,N_985,N_906);
and U1471 (N_1471,N_561,N_857);
and U1472 (N_1472,N_991,N_238);
xor U1473 (N_1473,N_215,N_444);
xor U1474 (N_1474,N_168,N_65);
xnor U1475 (N_1475,N_798,N_655);
and U1476 (N_1476,N_644,N_305);
nand U1477 (N_1477,N_177,N_76);
or U1478 (N_1478,N_47,N_706);
and U1479 (N_1479,N_767,N_832);
nand U1480 (N_1480,N_619,N_600);
nor U1481 (N_1481,N_954,N_879);
xnor U1482 (N_1482,N_635,N_116);
or U1483 (N_1483,N_930,N_202);
nor U1484 (N_1484,N_508,N_325);
xor U1485 (N_1485,N_506,N_513);
or U1486 (N_1486,N_950,N_661);
nor U1487 (N_1487,N_282,N_753);
xor U1488 (N_1488,N_278,N_722);
and U1489 (N_1489,N_118,N_328);
nor U1490 (N_1490,N_230,N_835);
xor U1491 (N_1491,N_124,N_893);
nor U1492 (N_1492,N_765,N_263);
nor U1493 (N_1493,N_242,N_9);
and U1494 (N_1494,N_452,N_713);
nor U1495 (N_1495,N_451,N_914);
xor U1496 (N_1496,N_216,N_757);
and U1497 (N_1497,N_551,N_912);
nor U1498 (N_1498,N_725,N_125);
or U1499 (N_1499,N_348,N_687);
nor U1500 (N_1500,N_910,N_146);
or U1501 (N_1501,N_289,N_360);
nor U1502 (N_1502,N_28,N_688);
and U1503 (N_1503,N_927,N_757);
xor U1504 (N_1504,N_767,N_626);
or U1505 (N_1505,N_880,N_960);
and U1506 (N_1506,N_341,N_308);
and U1507 (N_1507,N_142,N_869);
or U1508 (N_1508,N_212,N_469);
nor U1509 (N_1509,N_618,N_166);
nand U1510 (N_1510,N_903,N_930);
or U1511 (N_1511,N_824,N_586);
and U1512 (N_1512,N_737,N_17);
and U1513 (N_1513,N_975,N_234);
or U1514 (N_1514,N_937,N_901);
xor U1515 (N_1515,N_521,N_100);
nand U1516 (N_1516,N_233,N_746);
nand U1517 (N_1517,N_713,N_351);
xor U1518 (N_1518,N_134,N_591);
xor U1519 (N_1519,N_280,N_605);
nand U1520 (N_1520,N_359,N_695);
nor U1521 (N_1521,N_253,N_779);
nand U1522 (N_1522,N_507,N_75);
and U1523 (N_1523,N_534,N_179);
xor U1524 (N_1524,N_657,N_120);
nand U1525 (N_1525,N_329,N_800);
nor U1526 (N_1526,N_647,N_152);
xor U1527 (N_1527,N_382,N_994);
nand U1528 (N_1528,N_3,N_418);
nand U1529 (N_1529,N_978,N_678);
nor U1530 (N_1530,N_736,N_194);
xnor U1531 (N_1531,N_264,N_383);
and U1532 (N_1532,N_974,N_851);
nand U1533 (N_1533,N_470,N_975);
nor U1534 (N_1534,N_808,N_142);
and U1535 (N_1535,N_29,N_714);
nor U1536 (N_1536,N_514,N_172);
nor U1537 (N_1537,N_443,N_629);
xnor U1538 (N_1538,N_79,N_191);
and U1539 (N_1539,N_226,N_964);
nor U1540 (N_1540,N_644,N_268);
nor U1541 (N_1541,N_590,N_351);
nor U1542 (N_1542,N_120,N_372);
nor U1543 (N_1543,N_540,N_502);
or U1544 (N_1544,N_936,N_784);
xor U1545 (N_1545,N_312,N_329);
nand U1546 (N_1546,N_574,N_506);
nor U1547 (N_1547,N_434,N_181);
nand U1548 (N_1548,N_143,N_752);
nand U1549 (N_1549,N_881,N_749);
or U1550 (N_1550,N_956,N_542);
and U1551 (N_1551,N_238,N_397);
xnor U1552 (N_1552,N_0,N_403);
or U1553 (N_1553,N_413,N_833);
xnor U1554 (N_1554,N_509,N_51);
nand U1555 (N_1555,N_178,N_271);
xor U1556 (N_1556,N_38,N_481);
nand U1557 (N_1557,N_780,N_119);
and U1558 (N_1558,N_507,N_539);
xor U1559 (N_1559,N_896,N_509);
and U1560 (N_1560,N_7,N_181);
nand U1561 (N_1561,N_568,N_443);
and U1562 (N_1562,N_247,N_54);
or U1563 (N_1563,N_326,N_632);
or U1564 (N_1564,N_105,N_123);
xor U1565 (N_1565,N_730,N_874);
and U1566 (N_1566,N_568,N_407);
nand U1567 (N_1567,N_898,N_470);
nand U1568 (N_1568,N_366,N_496);
and U1569 (N_1569,N_951,N_992);
nor U1570 (N_1570,N_683,N_971);
nor U1571 (N_1571,N_154,N_583);
xor U1572 (N_1572,N_102,N_645);
and U1573 (N_1573,N_371,N_728);
nand U1574 (N_1574,N_668,N_439);
and U1575 (N_1575,N_376,N_560);
xnor U1576 (N_1576,N_87,N_661);
nand U1577 (N_1577,N_67,N_127);
nand U1578 (N_1578,N_763,N_332);
or U1579 (N_1579,N_494,N_378);
nand U1580 (N_1580,N_608,N_482);
or U1581 (N_1581,N_306,N_338);
xor U1582 (N_1582,N_882,N_460);
nor U1583 (N_1583,N_149,N_572);
xor U1584 (N_1584,N_593,N_229);
nand U1585 (N_1585,N_202,N_864);
xor U1586 (N_1586,N_45,N_345);
or U1587 (N_1587,N_978,N_437);
or U1588 (N_1588,N_145,N_791);
nor U1589 (N_1589,N_489,N_633);
nand U1590 (N_1590,N_736,N_720);
xor U1591 (N_1591,N_379,N_174);
nand U1592 (N_1592,N_15,N_463);
nand U1593 (N_1593,N_67,N_588);
xor U1594 (N_1594,N_548,N_505);
nand U1595 (N_1595,N_433,N_855);
and U1596 (N_1596,N_467,N_791);
or U1597 (N_1597,N_434,N_492);
and U1598 (N_1598,N_600,N_503);
and U1599 (N_1599,N_504,N_614);
and U1600 (N_1600,N_77,N_605);
or U1601 (N_1601,N_249,N_961);
and U1602 (N_1602,N_891,N_778);
nor U1603 (N_1603,N_148,N_776);
nand U1604 (N_1604,N_668,N_249);
xnor U1605 (N_1605,N_797,N_976);
nand U1606 (N_1606,N_644,N_8);
nor U1607 (N_1607,N_330,N_415);
nor U1608 (N_1608,N_420,N_150);
xnor U1609 (N_1609,N_241,N_610);
and U1610 (N_1610,N_941,N_439);
xor U1611 (N_1611,N_834,N_310);
nor U1612 (N_1612,N_225,N_782);
nand U1613 (N_1613,N_542,N_237);
nor U1614 (N_1614,N_530,N_234);
or U1615 (N_1615,N_549,N_317);
nor U1616 (N_1616,N_22,N_257);
nor U1617 (N_1617,N_497,N_20);
nor U1618 (N_1618,N_544,N_26);
nand U1619 (N_1619,N_35,N_597);
or U1620 (N_1620,N_834,N_708);
and U1621 (N_1621,N_735,N_863);
and U1622 (N_1622,N_948,N_271);
or U1623 (N_1623,N_971,N_412);
nand U1624 (N_1624,N_181,N_71);
nand U1625 (N_1625,N_132,N_600);
and U1626 (N_1626,N_559,N_562);
or U1627 (N_1627,N_516,N_605);
and U1628 (N_1628,N_243,N_301);
xnor U1629 (N_1629,N_772,N_363);
nor U1630 (N_1630,N_164,N_765);
xnor U1631 (N_1631,N_954,N_767);
or U1632 (N_1632,N_785,N_908);
nor U1633 (N_1633,N_804,N_830);
and U1634 (N_1634,N_987,N_46);
nand U1635 (N_1635,N_886,N_307);
xor U1636 (N_1636,N_385,N_103);
nor U1637 (N_1637,N_268,N_417);
nand U1638 (N_1638,N_533,N_173);
nand U1639 (N_1639,N_725,N_993);
and U1640 (N_1640,N_799,N_299);
nand U1641 (N_1641,N_981,N_273);
nand U1642 (N_1642,N_447,N_45);
nand U1643 (N_1643,N_765,N_334);
or U1644 (N_1644,N_168,N_413);
and U1645 (N_1645,N_21,N_104);
and U1646 (N_1646,N_859,N_778);
and U1647 (N_1647,N_459,N_387);
or U1648 (N_1648,N_38,N_63);
nand U1649 (N_1649,N_907,N_820);
nor U1650 (N_1650,N_759,N_690);
nand U1651 (N_1651,N_813,N_631);
or U1652 (N_1652,N_115,N_300);
and U1653 (N_1653,N_370,N_217);
xnor U1654 (N_1654,N_288,N_308);
and U1655 (N_1655,N_208,N_305);
nor U1656 (N_1656,N_150,N_381);
xor U1657 (N_1657,N_324,N_152);
nor U1658 (N_1658,N_115,N_525);
nand U1659 (N_1659,N_796,N_622);
or U1660 (N_1660,N_912,N_678);
xor U1661 (N_1661,N_639,N_47);
or U1662 (N_1662,N_159,N_36);
and U1663 (N_1663,N_992,N_610);
nor U1664 (N_1664,N_841,N_918);
or U1665 (N_1665,N_64,N_422);
xor U1666 (N_1666,N_822,N_184);
and U1667 (N_1667,N_371,N_432);
and U1668 (N_1668,N_450,N_253);
nand U1669 (N_1669,N_249,N_628);
nor U1670 (N_1670,N_14,N_727);
and U1671 (N_1671,N_749,N_531);
xnor U1672 (N_1672,N_222,N_513);
or U1673 (N_1673,N_104,N_686);
xnor U1674 (N_1674,N_927,N_545);
nor U1675 (N_1675,N_109,N_612);
nand U1676 (N_1676,N_385,N_405);
nor U1677 (N_1677,N_265,N_956);
nand U1678 (N_1678,N_882,N_886);
nand U1679 (N_1679,N_110,N_553);
or U1680 (N_1680,N_870,N_566);
nand U1681 (N_1681,N_997,N_338);
nor U1682 (N_1682,N_309,N_852);
nand U1683 (N_1683,N_125,N_279);
nand U1684 (N_1684,N_88,N_400);
or U1685 (N_1685,N_29,N_939);
nand U1686 (N_1686,N_865,N_593);
nor U1687 (N_1687,N_363,N_642);
nand U1688 (N_1688,N_828,N_938);
and U1689 (N_1689,N_876,N_133);
nand U1690 (N_1690,N_683,N_957);
nand U1691 (N_1691,N_737,N_846);
nor U1692 (N_1692,N_457,N_158);
nand U1693 (N_1693,N_166,N_101);
nor U1694 (N_1694,N_16,N_660);
and U1695 (N_1695,N_985,N_819);
nor U1696 (N_1696,N_334,N_129);
xnor U1697 (N_1697,N_792,N_73);
nand U1698 (N_1698,N_439,N_385);
nor U1699 (N_1699,N_450,N_998);
nand U1700 (N_1700,N_519,N_17);
nor U1701 (N_1701,N_197,N_489);
nor U1702 (N_1702,N_414,N_741);
xnor U1703 (N_1703,N_757,N_694);
nor U1704 (N_1704,N_107,N_280);
xnor U1705 (N_1705,N_702,N_154);
or U1706 (N_1706,N_970,N_571);
xor U1707 (N_1707,N_765,N_688);
and U1708 (N_1708,N_731,N_324);
nor U1709 (N_1709,N_800,N_546);
nand U1710 (N_1710,N_101,N_716);
nor U1711 (N_1711,N_719,N_544);
xor U1712 (N_1712,N_251,N_865);
or U1713 (N_1713,N_947,N_686);
or U1714 (N_1714,N_942,N_138);
or U1715 (N_1715,N_851,N_595);
or U1716 (N_1716,N_181,N_463);
nor U1717 (N_1717,N_318,N_687);
nand U1718 (N_1718,N_868,N_123);
nand U1719 (N_1719,N_641,N_247);
nand U1720 (N_1720,N_254,N_406);
and U1721 (N_1721,N_491,N_391);
and U1722 (N_1722,N_815,N_905);
xnor U1723 (N_1723,N_777,N_303);
and U1724 (N_1724,N_637,N_382);
nand U1725 (N_1725,N_152,N_275);
nor U1726 (N_1726,N_468,N_465);
or U1727 (N_1727,N_487,N_708);
and U1728 (N_1728,N_75,N_32);
and U1729 (N_1729,N_898,N_876);
or U1730 (N_1730,N_123,N_568);
nand U1731 (N_1731,N_547,N_473);
or U1732 (N_1732,N_740,N_180);
and U1733 (N_1733,N_719,N_867);
or U1734 (N_1734,N_503,N_335);
and U1735 (N_1735,N_713,N_531);
nor U1736 (N_1736,N_925,N_771);
and U1737 (N_1737,N_347,N_931);
xnor U1738 (N_1738,N_289,N_804);
nand U1739 (N_1739,N_287,N_199);
xor U1740 (N_1740,N_611,N_129);
nand U1741 (N_1741,N_494,N_224);
and U1742 (N_1742,N_280,N_877);
nor U1743 (N_1743,N_562,N_669);
xnor U1744 (N_1744,N_940,N_855);
and U1745 (N_1745,N_948,N_771);
nor U1746 (N_1746,N_711,N_685);
nor U1747 (N_1747,N_272,N_152);
and U1748 (N_1748,N_46,N_379);
and U1749 (N_1749,N_380,N_891);
or U1750 (N_1750,N_895,N_654);
xor U1751 (N_1751,N_268,N_942);
nand U1752 (N_1752,N_940,N_291);
and U1753 (N_1753,N_190,N_424);
nand U1754 (N_1754,N_530,N_408);
nor U1755 (N_1755,N_106,N_373);
xnor U1756 (N_1756,N_357,N_671);
and U1757 (N_1757,N_774,N_572);
nand U1758 (N_1758,N_52,N_710);
and U1759 (N_1759,N_69,N_754);
xnor U1760 (N_1760,N_600,N_555);
nand U1761 (N_1761,N_848,N_123);
and U1762 (N_1762,N_314,N_803);
and U1763 (N_1763,N_82,N_463);
and U1764 (N_1764,N_121,N_816);
or U1765 (N_1765,N_170,N_48);
xor U1766 (N_1766,N_632,N_476);
or U1767 (N_1767,N_646,N_356);
nor U1768 (N_1768,N_602,N_122);
xnor U1769 (N_1769,N_665,N_675);
nor U1770 (N_1770,N_236,N_147);
and U1771 (N_1771,N_847,N_561);
nor U1772 (N_1772,N_972,N_713);
nor U1773 (N_1773,N_176,N_709);
or U1774 (N_1774,N_784,N_117);
or U1775 (N_1775,N_257,N_594);
or U1776 (N_1776,N_796,N_865);
nand U1777 (N_1777,N_361,N_614);
or U1778 (N_1778,N_433,N_458);
nand U1779 (N_1779,N_94,N_806);
nand U1780 (N_1780,N_230,N_264);
and U1781 (N_1781,N_683,N_832);
or U1782 (N_1782,N_691,N_264);
nor U1783 (N_1783,N_980,N_544);
nand U1784 (N_1784,N_544,N_302);
and U1785 (N_1785,N_553,N_891);
xor U1786 (N_1786,N_862,N_753);
or U1787 (N_1787,N_605,N_885);
nand U1788 (N_1788,N_461,N_30);
nor U1789 (N_1789,N_22,N_727);
or U1790 (N_1790,N_906,N_686);
xnor U1791 (N_1791,N_475,N_287);
xnor U1792 (N_1792,N_55,N_939);
and U1793 (N_1793,N_818,N_881);
and U1794 (N_1794,N_351,N_401);
nor U1795 (N_1795,N_111,N_657);
and U1796 (N_1796,N_888,N_715);
xnor U1797 (N_1797,N_612,N_609);
nor U1798 (N_1798,N_102,N_931);
or U1799 (N_1799,N_263,N_128);
xnor U1800 (N_1800,N_824,N_259);
nor U1801 (N_1801,N_202,N_791);
nor U1802 (N_1802,N_105,N_531);
and U1803 (N_1803,N_267,N_953);
nand U1804 (N_1804,N_951,N_719);
or U1805 (N_1805,N_422,N_66);
xnor U1806 (N_1806,N_363,N_491);
nand U1807 (N_1807,N_940,N_220);
xnor U1808 (N_1808,N_856,N_420);
nor U1809 (N_1809,N_229,N_141);
or U1810 (N_1810,N_189,N_317);
nor U1811 (N_1811,N_8,N_800);
and U1812 (N_1812,N_989,N_501);
or U1813 (N_1813,N_127,N_232);
or U1814 (N_1814,N_681,N_692);
and U1815 (N_1815,N_516,N_190);
or U1816 (N_1816,N_469,N_138);
nor U1817 (N_1817,N_234,N_314);
and U1818 (N_1818,N_523,N_919);
xor U1819 (N_1819,N_639,N_970);
nand U1820 (N_1820,N_904,N_881);
xnor U1821 (N_1821,N_743,N_5);
and U1822 (N_1822,N_817,N_768);
and U1823 (N_1823,N_410,N_581);
xor U1824 (N_1824,N_933,N_109);
nand U1825 (N_1825,N_456,N_527);
and U1826 (N_1826,N_580,N_489);
nand U1827 (N_1827,N_220,N_925);
and U1828 (N_1828,N_883,N_964);
and U1829 (N_1829,N_562,N_3);
nand U1830 (N_1830,N_697,N_451);
nor U1831 (N_1831,N_268,N_993);
nand U1832 (N_1832,N_731,N_79);
xor U1833 (N_1833,N_517,N_524);
nand U1834 (N_1834,N_634,N_611);
nor U1835 (N_1835,N_529,N_602);
nand U1836 (N_1836,N_167,N_626);
or U1837 (N_1837,N_695,N_23);
and U1838 (N_1838,N_886,N_623);
nor U1839 (N_1839,N_479,N_344);
and U1840 (N_1840,N_113,N_605);
nor U1841 (N_1841,N_408,N_373);
or U1842 (N_1842,N_741,N_958);
and U1843 (N_1843,N_232,N_624);
nor U1844 (N_1844,N_573,N_312);
and U1845 (N_1845,N_220,N_439);
or U1846 (N_1846,N_537,N_82);
nor U1847 (N_1847,N_972,N_238);
nor U1848 (N_1848,N_398,N_712);
nand U1849 (N_1849,N_217,N_443);
and U1850 (N_1850,N_574,N_740);
xor U1851 (N_1851,N_554,N_894);
nor U1852 (N_1852,N_111,N_973);
and U1853 (N_1853,N_759,N_178);
and U1854 (N_1854,N_541,N_466);
or U1855 (N_1855,N_604,N_539);
xor U1856 (N_1856,N_981,N_754);
and U1857 (N_1857,N_68,N_871);
nor U1858 (N_1858,N_874,N_866);
nand U1859 (N_1859,N_171,N_533);
nor U1860 (N_1860,N_391,N_442);
nor U1861 (N_1861,N_669,N_542);
and U1862 (N_1862,N_187,N_742);
xnor U1863 (N_1863,N_262,N_163);
xor U1864 (N_1864,N_431,N_53);
nor U1865 (N_1865,N_918,N_995);
nor U1866 (N_1866,N_839,N_801);
nand U1867 (N_1867,N_168,N_776);
nor U1868 (N_1868,N_568,N_666);
xnor U1869 (N_1869,N_563,N_283);
nor U1870 (N_1870,N_404,N_593);
nand U1871 (N_1871,N_984,N_671);
xnor U1872 (N_1872,N_705,N_418);
nor U1873 (N_1873,N_621,N_758);
and U1874 (N_1874,N_212,N_770);
or U1875 (N_1875,N_434,N_425);
nand U1876 (N_1876,N_266,N_203);
nand U1877 (N_1877,N_261,N_813);
nor U1878 (N_1878,N_898,N_727);
nor U1879 (N_1879,N_963,N_43);
xor U1880 (N_1880,N_950,N_218);
nand U1881 (N_1881,N_41,N_873);
xnor U1882 (N_1882,N_553,N_870);
and U1883 (N_1883,N_539,N_400);
nand U1884 (N_1884,N_173,N_714);
and U1885 (N_1885,N_588,N_282);
nand U1886 (N_1886,N_792,N_506);
nor U1887 (N_1887,N_756,N_174);
nor U1888 (N_1888,N_216,N_381);
nor U1889 (N_1889,N_973,N_859);
or U1890 (N_1890,N_705,N_903);
xnor U1891 (N_1891,N_4,N_337);
xor U1892 (N_1892,N_703,N_120);
xnor U1893 (N_1893,N_526,N_99);
or U1894 (N_1894,N_943,N_507);
xor U1895 (N_1895,N_652,N_800);
nand U1896 (N_1896,N_876,N_834);
nor U1897 (N_1897,N_923,N_224);
and U1898 (N_1898,N_599,N_480);
and U1899 (N_1899,N_680,N_141);
xnor U1900 (N_1900,N_234,N_436);
xor U1901 (N_1901,N_453,N_163);
nor U1902 (N_1902,N_312,N_686);
nand U1903 (N_1903,N_276,N_315);
or U1904 (N_1904,N_196,N_293);
or U1905 (N_1905,N_689,N_457);
xnor U1906 (N_1906,N_673,N_186);
nand U1907 (N_1907,N_37,N_457);
xor U1908 (N_1908,N_409,N_986);
nand U1909 (N_1909,N_722,N_340);
nor U1910 (N_1910,N_766,N_921);
xor U1911 (N_1911,N_528,N_864);
and U1912 (N_1912,N_591,N_829);
nor U1913 (N_1913,N_998,N_899);
nand U1914 (N_1914,N_264,N_108);
nor U1915 (N_1915,N_2,N_63);
or U1916 (N_1916,N_438,N_66);
nor U1917 (N_1917,N_824,N_456);
and U1918 (N_1918,N_171,N_746);
nor U1919 (N_1919,N_34,N_581);
xor U1920 (N_1920,N_177,N_84);
and U1921 (N_1921,N_341,N_919);
or U1922 (N_1922,N_233,N_647);
nand U1923 (N_1923,N_362,N_861);
and U1924 (N_1924,N_583,N_692);
xor U1925 (N_1925,N_726,N_882);
nand U1926 (N_1926,N_87,N_592);
or U1927 (N_1927,N_80,N_661);
xor U1928 (N_1928,N_957,N_272);
xnor U1929 (N_1929,N_802,N_157);
and U1930 (N_1930,N_643,N_704);
xor U1931 (N_1931,N_533,N_256);
nor U1932 (N_1932,N_230,N_253);
nor U1933 (N_1933,N_21,N_782);
xnor U1934 (N_1934,N_946,N_56);
or U1935 (N_1935,N_637,N_113);
xor U1936 (N_1936,N_919,N_712);
nand U1937 (N_1937,N_34,N_808);
nor U1938 (N_1938,N_370,N_363);
nor U1939 (N_1939,N_608,N_974);
or U1940 (N_1940,N_387,N_118);
and U1941 (N_1941,N_417,N_988);
nor U1942 (N_1942,N_428,N_676);
nand U1943 (N_1943,N_53,N_306);
or U1944 (N_1944,N_336,N_697);
nand U1945 (N_1945,N_384,N_985);
nor U1946 (N_1946,N_948,N_93);
or U1947 (N_1947,N_144,N_518);
or U1948 (N_1948,N_964,N_49);
nor U1949 (N_1949,N_429,N_267);
xnor U1950 (N_1950,N_459,N_468);
nor U1951 (N_1951,N_956,N_157);
xor U1952 (N_1952,N_361,N_69);
nand U1953 (N_1953,N_341,N_789);
and U1954 (N_1954,N_965,N_403);
and U1955 (N_1955,N_203,N_702);
xnor U1956 (N_1956,N_84,N_943);
xor U1957 (N_1957,N_722,N_923);
nand U1958 (N_1958,N_641,N_230);
nand U1959 (N_1959,N_422,N_723);
and U1960 (N_1960,N_202,N_577);
nand U1961 (N_1961,N_314,N_627);
nor U1962 (N_1962,N_723,N_416);
or U1963 (N_1963,N_238,N_221);
and U1964 (N_1964,N_319,N_415);
and U1965 (N_1965,N_33,N_174);
nand U1966 (N_1966,N_294,N_570);
xnor U1967 (N_1967,N_621,N_353);
nand U1968 (N_1968,N_749,N_919);
xnor U1969 (N_1969,N_239,N_191);
nor U1970 (N_1970,N_383,N_784);
xor U1971 (N_1971,N_718,N_482);
and U1972 (N_1972,N_880,N_514);
or U1973 (N_1973,N_750,N_314);
nor U1974 (N_1974,N_98,N_209);
xnor U1975 (N_1975,N_468,N_838);
nor U1976 (N_1976,N_961,N_699);
nand U1977 (N_1977,N_980,N_255);
nand U1978 (N_1978,N_759,N_105);
nor U1979 (N_1979,N_833,N_144);
nand U1980 (N_1980,N_570,N_431);
nor U1981 (N_1981,N_834,N_63);
and U1982 (N_1982,N_262,N_474);
and U1983 (N_1983,N_13,N_338);
or U1984 (N_1984,N_618,N_262);
and U1985 (N_1985,N_378,N_134);
and U1986 (N_1986,N_332,N_764);
nand U1987 (N_1987,N_147,N_713);
nand U1988 (N_1988,N_617,N_271);
or U1989 (N_1989,N_990,N_683);
and U1990 (N_1990,N_780,N_298);
xor U1991 (N_1991,N_349,N_387);
or U1992 (N_1992,N_693,N_5);
nand U1993 (N_1993,N_889,N_51);
xnor U1994 (N_1994,N_709,N_455);
and U1995 (N_1995,N_833,N_28);
nor U1996 (N_1996,N_173,N_601);
nor U1997 (N_1997,N_175,N_142);
xor U1998 (N_1998,N_541,N_539);
xnor U1999 (N_1999,N_65,N_220);
nor U2000 (N_2000,N_1448,N_1591);
nor U2001 (N_2001,N_1502,N_1018);
and U2002 (N_2002,N_1428,N_1839);
and U2003 (N_2003,N_1741,N_1935);
or U2004 (N_2004,N_1518,N_1889);
and U2005 (N_2005,N_1348,N_1961);
nor U2006 (N_2006,N_1792,N_1442);
and U2007 (N_2007,N_1795,N_1415);
or U2008 (N_2008,N_1864,N_1747);
nand U2009 (N_2009,N_1579,N_1109);
xor U2010 (N_2010,N_1509,N_1954);
or U2011 (N_2011,N_1708,N_1359);
or U2012 (N_2012,N_1270,N_1944);
and U2013 (N_2013,N_1079,N_1520);
or U2014 (N_2014,N_1312,N_1044);
nor U2015 (N_2015,N_1342,N_1580);
nor U2016 (N_2016,N_1821,N_1832);
nor U2017 (N_2017,N_1854,N_1843);
or U2018 (N_2018,N_1040,N_1240);
xor U2019 (N_2019,N_1534,N_1541);
nand U2020 (N_2020,N_1715,N_1464);
or U2021 (N_2021,N_1337,N_1141);
or U2022 (N_2022,N_1144,N_1016);
or U2023 (N_2023,N_1196,N_1288);
or U2024 (N_2024,N_1530,N_1666);
xor U2025 (N_2025,N_1164,N_1896);
xnor U2026 (N_2026,N_1368,N_1411);
or U2027 (N_2027,N_1631,N_1965);
or U2028 (N_2028,N_1149,N_1172);
nand U2029 (N_2029,N_1835,N_1135);
or U2030 (N_2030,N_1734,N_1540);
and U2031 (N_2031,N_1081,N_1251);
xnor U2032 (N_2032,N_1638,N_1655);
nand U2033 (N_2033,N_1093,N_1515);
or U2034 (N_2034,N_1231,N_1074);
and U2035 (N_2035,N_1301,N_1077);
nand U2036 (N_2036,N_1254,N_1159);
and U2037 (N_2037,N_1067,N_1269);
xnor U2038 (N_2038,N_1879,N_1942);
or U2039 (N_2039,N_1460,N_1228);
nand U2040 (N_2040,N_1725,N_1105);
xor U2041 (N_2041,N_1969,N_1165);
nor U2042 (N_2042,N_1786,N_1177);
or U2043 (N_2043,N_1863,N_1952);
or U2044 (N_2044,N_1053,N_1717);
and U2045 (N_2045,N_1204,N_1116);
nor U2046 (N_2046,N_1552,N_1769);
nand U2047 (N_2047,N_1709,N_1878);
or U2048 (N_2048,N_1227,N_1134);
xor U2049 (N_2049,N_1259,N_1533);
xnor U2050 (N_2050,N_1023,N_1922);
or U2051 (N_2051,N_1635,N_1788);
or U2052 (N_2052,N_1924,N_1179);
or U2053 (N_2053,N_1380,N_1298);
xor U2054 (N_2054,N_1086,N_1388);
nand U2055 (N_2055,N_1949,N_1997);
and U2056 (N_2056,N_1966,N_1963);
nand U2057 (N_2057,N_1687,N_1557);
nor U2058 (N_2058,N_1375,N_1885);
and U2059 (N_2059,N_1385,N_1307);
or U2060 (N_2060,N_1595,N_1890);
nor U2061 (N_2061,N_1948,N_1094);
or U2062 (N_2062,N_1527,N_1775);
nand U2063 (N_2063,N_1265,N_1562);
or U2064 (N_2064,N_1893,N_1493);
and U2065 (N_2065,N_1229,N_1103);
nor U2066 (N_2066,N_1106,N_1536);
nor U2067 (N_2067,N_1294,N_1667);
and U2068 (N_2068,N_1358,N_1313);
nand U2069 (N_2069,N_1669,N_1009);
and U2070 (N_2070,N_1439,N_1146);
or U2071 (N_2071,N_1791,N_1903);
xnor U2072 (N_2072,N_1226,N_1455);
or U2073 (N_2073,N_1473,N_1751);
and U2074 (N_2074,N_1857,N_1977);
xor U2075 (N_2075,N_1783,N_1213);
and U2076 (N_2076,N_1360,N_1349);
xnor U2077 (N_2077,N_1812,N_1277);
nand U2078 (N_2078,N_1249,N_1987);
nand U2079 (N_2079,N_1431,N_1412);
and U2080 (N_2080,N_1723,N_1034);
nand U2081 (N_2081,N_1891,N_1160);
nand U2082 (N_2082,N_1133,N_1266);
or U2083 (N_2083,N_1754,N_1823);
or U2084 (N_2084,N_1874,N_1806);
or U2085 (N_2085,N_1553,N_1290);
nand U2086 (N_2086,N_1576,N_1753);
nand U2087 (N_2087,N_1653,N_1171);
xnor U2088 (N_2088,N_1524,N_1611);
nand U2089 (N_2089,N_1316,N_1841);
nand U2090 (N_2090,N_1237,N_1814);
xnor U2091 (N_2091,N_1472,N_1773);
and U2092 (N_2092,N_1690,N_1583);
or U2093 (N_2093,N_1733,N_1990);
and U2094 (N_2094,N_1590,N_1068);
nor U2095 (N_2095,N_1726,N_1789);
nor U2096 (N_2096,N_1759,N_1039);
or U2097 (N_2097,N_1427,N_1100);
nand U2098 (N_2098,N_1847,N_1858);
and U2099 (N_2099,N_1192,N_1742);
nor U2100 (N_2100,N_1189,N_1292);
nor U2101 (N_2101,N_1679,N_1441);
or U2102 (N_2102,N_1529,N_1008);
nand U2103 (N_2103,N_1853,N_1232);
nand U2104 (N_2104,N_1466,N_1550);
or U2105 (N_2105,N_1596,N_1822);
nand U2106 (N_2106,N_1933,N_1060);
nor U2107 (N_2107,N_1664,N_1461);
nor U2108 (N_2108,N_1410,N_1408);
or U2109 (N_2109,N_1284,N_1908);
xor U2110 (N_2110,N_1300,N_1767);
nand U2111 (N_2111,N_1481,N_1967);
and U2112 (N_2112,N_1123,N_1581);
nor U2113 (N_2113,N_1193,N_1303);
or U2114 (N_2114,N_1622,N_1125);
nand U2115 (N_2115,N_1030,N_1923);
nor U2116 (N_2116,N_1684,N_1994);
nand U2117 (N_2117,N_1444,N_1061);
xnor U2118 (N_2118,N_1201,N_1128);
nand U2119 (N_2119,N_1613,N_1402);
nor U2120 (N_2120,N_1906,N_1980);
nor U2121 (N_2121,N_1956,N_1943);
nor U2122 (N_2122,N_1918,N_1072);
or U2123 (N_2123,N_1744,N_1138);
nand U2124 (N_2124,N_1712,N_1048);
and U2125 (N_2125,N_1830,N_1117);
nor U2126 (N_2126,N_1677,N_1334);
xor U2127 (N_2127,N_1208,N_1505);
xnor U2128 (N_2128,N_1357,N_1275);
nor U2129 (N_2129,N_1434,N_1567);
xnor U2130 (N_2130,N_1148,N_1339);
nand U2131 (N_2131,N_1362,N_1291);
or U2132 (N_2132,N_1849,N_1364);
xnor U2133 (N_2133,N_1497,N_1834);
xnor U2134 (N_2134,N_1486,N_1819);
or U2135 (N_2135,N_1480,N_1031);
nor U2136 (N_2136,N_1054,N_1750);
and U2137 (N_2137,N_1500,N_1028);
nor U2138 (N_2138,N_1025,N_1003);
or U2139 (N_2139,N_1673,N_1572);
nand U2140 (N_2140,N_1945,N_1575);
and U2141 (N_2141,N_1245,N_1899);
nand U2142 (N_2142,N_1979,N_1671);
xnor U2143 (N_2143,N_1365,N_1212);
or U2144 (N_2144,N_1131,N_1153);
and U2145 (N_2145,N_1507,N_1716);
nor U2146 (N_2146,N_1384,N_1218);
or U2147 (N_2147,N_1454,N_1996);
nand U2148 (N_2148,N_1652,N_1701);
or U2149 (N_2149,N_1198,N_1356);
xor U2150 (N_2150,N_1501,N_1381);
and U2151 (N_2151,N_1665,N_1696);
nand U2152 (N_2152,N_1453,N_1563);
or U2153 (N_2153,N_1264,N_1901);
and U2154 (N_2154,N_1881,N_1186);
or U2155 (N_2155,N_1598,N_1098);
xor U2156 (N_2156,N_1621,N_1037);
nor U2157 (N_2157,N_1816,N_1970);
nor U2158 (N_2158,N_1634,N_1156);
or U2159 (N_2159,N_1763,N_1260);
xnor U2160 (N_2160,N_1605,N_1920);
nand U2161 (N_2161,N_1194,N_1147);
and U2162 (N_2162,N_1719,N_1538);
xor U2163 (N_2163,N_1882,N_1535);
xor U2164 (N_2164,N_1808,N_1555);
or U2165 (N_2165,N_1805,N_1941);
or U2166 (N_2166,N_1045,N_1324);
and U2167 (N_2167,N_1617,N_1962);
nand U2168 (N_2168,N_1309,N_1223);
and U2169 (N_2169,N_1958,N_1776);
nand U2170 (N_2170,N_1661,N_1482);
or U2171 (N_2171,N_1953,N_1981);
or U2172 (N_2172,N_1803,N_1021);
or U2173 (N_2173,N_1510,N_1475);
xnor U2174 (N_2174,N_1503,N_1571);
nor U2175 (N_2175,N_1258,N_1246);
and U2176 (N_2176,N_1235,N_1276);
nor U2177 (N_2177,N_1939,N_1624);
or U2178 (N_2178,N_1318,N_1799);
or U2179 (N_2179,N_1674,N_1247);
and U2180 (N_2180,N_1871,N_1568);
or U2181 (N_2181,N_1785,N_1478);
nand U2182 (N_2182,N_1930,N_1971);
or U2183 (N_2183,N_1096,N_1488);
xnor U2184 (N_2184,N_1985,N_1202);
nand U2185 (N_2185,N_1739,N_1066);
nor U2186 (N_2186,N_1566,N_1209);
and U2187 (N_2187,N_1872,N_1813);
nand U2188 (N_2188,N_1422,N_1090);
and U2189 (N_2189,N_1297,N_1038);
and U2190 (N_2190,N_1526,N_1451);
xor U2191 (N_2191,N_1333,N_1217);
or U2192 (N_2192,N_1440,N_1588);
and U2193 (N_2193,N_1487,N_1593);
or U2194 (N_2194,N_1817,N_1974);
or U2195 (N_2195,N_1836,N_1724);
and U2196 (N_2196,N_1564,N_1367);
xor U2197 (N_2197,N_1554,N_1975);
or U2198 (N_2198,N_1917,N_1216);
xnor U2199 (N_2199,N_1798,N_1938);
nor U2200 (N_2200,N_1335,N_1043);
nand U2201 (N_2201,N_1435,N_1080);
nor U2202 (N_2202,N_1386,N_1542);
and U2203 (N_2203,N_1946,N_1927);
nor U2204 (N_2204,N_1599,N_1433);
xnor U2205 (N_2205,N_1886,N_1104);
and U2206 (N_2206,N_1569,N_1406);
nand U2207 (N_2207,N_1326,N_1797);
or U2208 (N_2208,N_1910,N_1490);
or U2209 (N_2209,N_1657,N_1662);
or U2210 (N_2210,N_1166,N_1921);
nand U2211 (N_2211,N_1175,N_1085);
or U2212 (N_2212,N_1012,N_1728);
or U2213 (N_2213,N_1796,N_1089);
nor U2214 (N_2214,N_1187,N_1110);
nand U2215 (N_2215,N_1136,N_1860);
or U2216 (N_2216,N_1668,N_1594);
nor U2217 (N_2217,N_1115,N_1646);
xnor U2218 (N_2218,N_1285,N_1261);
and U2219 (N_2219,N_1727,N_1928);
nor U2220 (N_2220,N_1907,N_1852);
or U2221 (N_2221,N_1268,N_1810);
xnor U2222 (N_2222,N_1035,N_1888);
xnor U2223 (N_2223,N_1702,N_1140);
nor U2224 (N_2224,N_1831,N_1467);
nor U2225 (N_2225,N_1625,N_1984);
xor U2226 (N_2226,N_1376,N_1760);
and U2227 (N_2227,N_1102,N_1416);
nor U2228 (N_2228,N_1282,N_1620);
and U2229 (N_2229,N_1456,N_1614);
nor U2230 (N_2230,N_1001,N_1736);
nor U2231 (N_2231,N_1829,N_1310);
xor U2232 (N_2232,N_1837,N_1462);
nand U2233 (N_2233,N_1130,N_1710);
or U2234 (N_2234,N_1393,N_1644);
nand U2235 (N_2235,N_1573,N_1417);
and U2236 (N_2236,N_1523,N_1374);
or U2237 (N_2237,N_1982,N_1793);
nor U2238 (N_2238,N_1919,N_1256);
and U2239 (N_2239,N_1252,N_1663);
nor U2240 (N_2240,N_1768,N_1787);
nor U2241 (N_2241,N_1735,N_1900);
nor U2242 (N_2242,N_1940,N_1244);
or U2243 (N_2243,N_1629,N_1512);
nand U2244 (N_2244,N_1587,N_1586);
nor U2245 (N_2245,N_1051,N_1113);
nor U2246 (N_2246,N_1112,N_1851);
or U2247 (N_2247,N_1369,N_1828);
nand U2248 (N_2248,N_1957,N_1468);
xnor U2249 (N_2249,N_1818,N_1637);
and U2250 (N_2250,N_1731,N_1407);
or U2251 (N_2251,N_1092,N_1707);
nand U2252 (N_2252,N_1354,N_1761);
nor U2253 (N_2253,N_1366,N_1041);
and U2254 (N_2254,N_1405,N_1219);
and U2255 (N_2255,N_1641,N_1762);
nand U2256 (N_2256,N_1397,N_1479);
nand U2257 (N_2257,N_1145,N_1859);
xnor U2258 (N_2258,N_1685,N_1695);
nor U2259 (N_2259,N_1531,N_1826);
or U2260 (N_2260,N_1004,N_1332);
nor U2261 (N_2261,N_1833,N_1352);
nand U2262 (N_2262,N_1325,N_1314);
or U2263 (N_2263,N_1999,N_1027);
and U2264 (N_2264,N_1781,N_1511);
and U2265 (N_2265,N_1032,N_1937);
xor U2266 (N_2266,N_1181,N_1976);
and U2267 (N_2267,N_1111,N_1010);
or U2268 (N_2268,N_1532,N_1489);
xnor U2269 (N_2269,N_1525,N_1749);
nor U2270 (N_2270,N_1350,N_1336);
or U2271 (N_2271,N_1737,N_1764);
or U2272 (N_2272,N_1867,N_1912);
nor U2273 (N_2273,N_1271,N_1597);
or U2274 (N_2274,N_1191,N_1029);
or U2275 (N_2275,N_1391,N_1222);
nor U2276 (N_2276,N_1495,N_1255);
nand U2277 (N_2277,N_1328,N_1423);
xnor U2278 (N_2278,N_1049,N_1215);
xor U2279 (N_2279,N_1185,N_1378);
nor U2280 (N_2280,N_1399,N_1457);
xnor U2281 (N_2281,N_1017,N_1643);
nand U2282 (N_2282,N_1766,N_1295);
or U2283 (N_2283,N_1107,N_1862);
nand U2284 (N_2284,N_1913,N_1647);
or U2285 (N_2285,N_1331,N_1861);
and U2286 (N_2286,N_1800,N_1400);
xnor U2287 (N_2287,N_1689,N_1302);
and U2288 (N_2288,N_1551,N_1752);
xor U2289 (N_2289,N_1516,N_1404);
nor U2290 (N_2290,N_1437,N_1305);
nand U2291 (N_2291,N_1024,N_1273);
and U2292 (N_2292,N_1195,N_1603);
nand U2293 (N_2293,N_1755,N_1429);
nor U2294 (N_2294,N_1120,N_1340);
and U2295 (N_2295,N_1238,N_1746);
xnor U2296 (N_2296,N_1281,N_1809);
xor U2297 (N_2297,N_1320,N_1697);
nor U2298 (N_2298,N_1802,N_1543);
xnor U2299 (N_2299,N_1883,N_1866);
nand U2300 (N_2300,N_1811,N_1983);
nand U2301 (N_2301,N_1558,N_1430);
and U2302 (N_2302,N_1064,N_1827);
xor U2303 (N_2303,N_1248,N_1322);
nand U2304 (N_2304,N_1151,N_1925);
or U2305 (N_2305,N_1703,N_1680);
and U2306 (N_2306,N_1855,N_1865);
xnor U2307 (N_2307,N_1387,N_1779);
xnor U2308 (N_2308,N_1278,N_1065);
nand U2309 (N_2309,N_1355,N_1628);
nand U2310 (N_2310,N_1496,N_1063);
and U2311 (N_2311,N_1623,N_1126);
xor U2312 (N_2312,N_1926,N_1272);
and U2313 (N_2313,N_1197,N_1498);
xor U2314 (N_2314,N_1132,N_1492);
nor U2315 (N_2315,N_1820,N_1539);
xnor U2316 (N_2316,N_1678,N_1311);
xor U2317 (N_2317,N_1162,N_1119);
or U2318 (N_2318,N_1200,N_1875);
xor U2319 (N_2319,N_1506,N_1911);
xor U2320 (N_2320,N_1420,N_1998);
nand U2321 (N_2321,N_1155,N_1168);
xnor U2322 (N_2322,N_1091,N_1304);
nor U2323 (N_2323,N_1438,N_1377);
or U2324 (N_2324,N_1777,N_1729);
and U2325 (N_2325,N_1650,N_1955);
xnor U2326 (N_2326,N_1884,N_1286);
or U2327 (N_2327,N_1545,N_1528);
and U2328 (N_2328,N_1609,N_1289);
nand U2329 (N_2329,N_1398,N_1280);
xor U2330 (N_2330,N_1242,N_1183);
nand U2331 (N_2331,N_1452,N_1071);
or U2332 (N_2332,N_1721,N_1718);
or U2333 (N_2333,N_1392,N_1892);
xor U2334 (N_2334,N_1182,N_1559);
nor U2335 (N_2335,N_1902,N_1459);
and U2336 (N_2336,N_1062,N_1139);
and U2337 (N_2337,N_1790,N_1915);
nor U2338 (N_2338,N_1394,N_1263);
xor U2339 (N_2339,N_1672,N_1083);
nor U2340 (N_2340,N_1262,N_1167);
and U2341 (N_2341,N_1600,N_1042);
nor U2342 (N_2342,N_1383,N_1108);
or U2343 (N_2343,N_1005,N_1670);
xnor U2344 (N_2344,N_1341,N_1758);
nor U2345 (N_2345,N_1838,N_1073);
nor U2346 (N_2346,N_1577,N_1210);
or U2347 (N_2347,N_1711,N_1158);
or U2348 (N_2348,N_1287,N_1992);
nor U2349 (N_2349,N_1152,N_1693);
nor U2350 (N_2350,N_1801,N_1691);
xnor U2351 (N_2351,N_1639,N_1403);
xnor U2352 (N_2352,N_1253,N_1705);
nor U2353 (N_2353,N_1170,N_1959);
and U2354 (N_2354,N_1471,N_1330);
xnor U2355 (N_2355,N_1076,N_1447);
nor U2356 (N_2356,N_1909,N_1698);
and U2357 (N_2357,N_1589,N_1057);
xnor U2358 (N_2358,N_1163,N_1722);
nand U2359 (N_2359,N_1157,N_1544);
nor U2360 (N_2360,N_1418,N_1494);
nor U2361 (N_2361,N_1211,N_1905);
xnor U2362 (N_2362,N_1986,N_1056);
nor U2363 (N_2363,N_1425,N_1887);
nand U2364 (N_2364,N_1602,N_1221);
nand U2365 (N_2365,N_1648,N_1007);
xor U2366 (N_2366,N_1426,N_1880);
xor U2367 (N_2367,N_1842,N_1205);
and U2368 (N_2368,N_1476,N_1154);
and U2369 (N_2369,N_1960,N_1612);
nand U2370 (N_2370,N_1675,N_1561);
nand U2371 (N_2371,N_1804,N_1371);
nand U2372 (N_2372,N_1306,N_1274);
xnor U2373 (N_2373,N_1973,N_1346);
and U2374 (N_2374,N_1607,N_1379);
xnor U2375 (N_2375,N_1869,N_1772);
and U2376 (N_2376,N_1636,N_1345);
or U2377 (N_2377,N_1225,N_1700);
xnor U2378 (N_2378,N_1548,N_1449);
nand U2379 (N_2379,N_1848,N_1504);
or U2380 (N_2380,N_1771,N_1582);
nand U2381 (N_2381,N_1450,N_1950);
xnor U2382 (N_2382,N_1323,N_1180);
nor U2383 (N_2383,N_1936,N_1026);
nor U2384 (N_2384,N_1084,N_1432);
or U2385 (N_2385,N_1315,N_1730);
nor U2386 (N_2386,N_1382,N_1267);
nor U2387 (N_2387,N_1560,N_1161);
nand U2388 (N_2388,N_1220,N_1929);
and U2389 (N_2389,N_1150,N_1047);
and U2390 (N_2390,N_1932,N_1069);
and U2391 (N_2391,N_1856,N_1458);
or U2392 (N_2392,N_1142,N_1485);
nand U2393 (N_2393,N_1713,N_1389);
xnor U2394 (N_2394,N_1143,N_1978);
nand U2395 (N_2395,N_1088,N_1988);
nor U2396 (N_2396,N_1414,N_1070);
nand U2397 (N_2397,N_1514,N_1327);
nand U2398 (N_2398,N_1465,N_1995);
and U2399 (N_2399,N_1230,N_1549);
nand U2400 (N_2400,N_1840,N_1214);
nand U2401 (N_2401,N_1916,N_1784);
nand U2402 (N_2402,N_1206,N_1203);
nor U2403 (N_2403,N_1870,N_1199);
nor U2404 (N_2404,N_1250,N_1825);
or U2405 (N_2405,N_1129,N_1014);
xor U2406 (N_2406,N_1424,N_1319);
xor U2407 (N_2407,N_1483,N_1877);
or U2408 (N_2408,N_1618,N_1022);
nor U2409 (N_2409,N_1770,N_1344);
or U2410 (N_2410,N_1642,N_1293);
nand U2411 (N_2411,N_1658,N_1178);
and U2412 (N_2412,N_1714,N_1006);
and U2413 (N_2413,N_1876,N_1565);
or U2414 (N_2414,N_1615,N_1522);
and U2415 (N_2415,N_1015,N_1519);
nand U2416 (N_2416,N_1169,N_1633);
or U2417 (N_2417,N_1904,N_1127);
nor U2418 (N_2418,N_1396,N_1989);
nand U2419 (N_2419,N_1121,N_1207);
nor U2420 (N_2420,N_1075,N_1748);
xor U2421 (N_2421,N_1627,N_1363);
and U2422 (N_2422,N_1968,N_1436);
xnor U2423 (N_2423,N_1972,N_1329);
or U2424 (N_2424,N_1898,N_1894);
xnor U2425 (N_2425,N_1547,N_1055);
nand U2426 (N_2426,N_1610,N_1868);
nand U2427 (N_2427,N_1421,N_1188);
xnor U2428 (N_2428,N_1413,N_1844);
or U2429 (N_2429,N_1570,N_1019);
or U2430 (N_2430,N_1390,N_1176);
or U2431 (N_2431,N_1095,N_1521);
or U2432 (N_2432,N_1082,N_1608);
or U2433 (N_2433,N_1738,N_1616);
and U2434 (N_2434,N_1630,N_1078);
nand U2435 (N_2435,N_1353,N_1991);
xnor U2436 (N_2436,N_1578,N_1619);
and U2437 (N_2437,N_1470,N_1036);
nand U2438 (N_2438,N_1740,N_1584);
xnor U2439 (N_2439,N_1101,N_1592);
or U2440 (N_2440,N_1299,N_1745);
or U2441 (N_2441,N_1059,N_1824);
nor U2442 (N_2442,N_1118,N_1640);
xnor U2443 (N_2443,N_1321,N_1681);
nand U2444 (N_2444,N_1020,N_1914);
xor U2445 (N_2445,N_1477,N_1651);
or U2446 (N_2446,N_1243,N_1343);
and U2447 (N_2447,N_1757,N_1688);
xor U2448 (N_2448,N_1845,N_1947);
and U2449 (N_2449,N_1011,N_1308);
and U2450 (N_2450,N_1692,N_1013);
or U2451 (N_2451,N_1370,N_1720);
xor U2452 (N_2452,N_1234,N_1951);
nand U2453 (N_2453,N_1174,N_1469);
xor U2454 (N_2454,N_1517,N_1683);
xor U2455 (N_2455,N_1283,N_1445);
and U2456 (N_2456,N_1756,N_1137);
and U2457 (N_2457,N_1699,N_1484);
and U2458 (N_2458,N_1654,N_1704);
or U2459 (N_2459,N_1513,N_1537);
and U2460 (N_2460,N_1087,N_1765);
or U2461 (N_2461,N_1224,N_1897);
xnor U2462 (N_2462,N_1964,N_1052);
xor U2463 (N_2463,N_1317,N_1508);
nor U2464 (N_2464,N_1000,N_1645);
and U2465 (N_2465,N_1463,N_1419);
xnor U2466 (N_2466,N_1807,N_1491);
and U2467 (N_2467,N_1993,N_1184);
nand U2468 (N_2468,N_1122,N_1686);
nor U2469 (N_2469,N_1649,N_1190);
xor U2470 (N_2470,N_1794,N_1934);
nand U2471 (N_2471,N_1443,N_1173);
nand U2472 (N_2472,N_1401,N_1409);
nand U2473 (N_2473,N_1780,N_1743);
and U2474 (N_2474,N_1850,N_1395);
nor U2475 (N_2475,N_1233,N_1546);
nor U2476 (N_2476,N_1446,N_1556);
xor U2477 (N_2477,N_1241,N_1931);
and U2478 (N_2478,N_1676,N_1050);
xnor U2479 (N_2479,N_1296,N_1632);
nor U2480 (N_2480,N_1585,N_1499);
nand U2481 (N_2481,N_1474,N_1778);
nand U2482 (N_2482,N_1706,N_1046);
nor U2483 (N_2483,N_1604,N_1279);
nor U2484 (N_2484,N_1257,N_1774);
or U2485 (N_2485,N_1347,N_1372);
nand U2486 (N_2486,N_1002,N_1732);
or U2487 (N_2487,N_1815,N_1626);
xor U2488 (N_2488,N_1659,N_1682);
xnor U2489 (N_2489,N_1873,N_1236);
or U2490 (N_2490,N_1351,N_1373);
nor U2491 (N_2491,N_1239,N_1338);
or U2492 (N_2492,N_1694,N_1606);
or U2493 (N_2493,N_1058,N_1574);
xor U2494 (N_2494,N_1033,N_1846);
nor U2495 (N_2495,N_1099,N_1114);
or U2496 (N_2496,N_1124,N_1601);
or U2497 (N_2497,N_1361,N_1660);
and U2498 (N_2498,N_1097,N_1782);
nand U2499 (N_2499,N_1656,N_1895);
nor U2500 (N_2500,N_1426,N_1877);
nor U2501 (N_2501,N_1544,N_1177);
and U2502 (N_2502,N_1088,N_1275);
nand U2503 (N_2503,N_1645,N_1489);
or U2504 (N_2504,N_1363,N_1607);
and U2505 (N_2505,N_1792,N_1540);
nand U2506 (N_2506,N_1615,N_1410);
nor U2507 (N_2507,N_1647,N_1848);
or U2508 (N_2508,N_1334,N_1195);
nand U2509 (N_2509,N_1369,N_1922);
and U2510 (N_2510,N_1042,N_1668);
xnor U2511 (N_2511,N_1661,N_1513);
or U2512 (N_2512,N_1092,N_1199);
and U2513 (N_2513,N_1631,N_1717);
nand U2514 (N_2514,N_1665,N_1393);
nand U2515 (N_2515,N_1673,N_1609);
and U2516 (N_2516,N_1183,N_1268);
nor U2517 (N_2517,N_1240,N_1458);
and U2518 (N_2518,N_1660,N_1424);
xor U2519 (N_2519,N_1746,N_1408);
nor U2520 (N_2520,N_1280,N_1040);
nand U2521 (N_2521,N_1724,N_1995);
xor U2522 (N_2522,N_1359,N_1083);
or U2523 (N_2523,N_1424,N_1171);
and U2524 (N_2524,N_1409,N_1633);
or U2525 (N_2525,N_1918,N_1775);
nor U2526 (N_2526,N_1703,N_1926);
xor U2527 (N_2527,N_1408,N_1569);
nor U2528 (N_2528,N_1935,N_1236);
nand U2529 (N_2529,N_1748,N_1076);
nor U2530 (N_2530,N_1324,N_1724);
xnor U2531 (N_2531,N_1969,N_1817);
or U2532 (N_2532,N_1568,N_1630);
or U2533 (N_2533,N_1806,N_1426);
xnor U2534 (N_2534,N_1764,N_1623);
nand U2535 (N_2535,N_1208,N_1817);
or U2536 (N_2536,N_1167,N_1614);
and U2537 (N_2537,N_1013,N_1962);
nand U2538 (N_2538,N_1663,N_1476);
or U2539 (N_2539,N_1754,N_1627);
or U2540 (N_2540,N_1261,N_1842);
or U2541 (N_2541,N_1884,N_1791);
nand U2542 (N_2542,N_1275,N_1958);
nor U2543 (N_2543,N_1573,N_1702);
and U2544 (N_2544,N_1925,N_1623);
nor U2545 (N_2545,N_1041,N_1088);
nor U2546 (N_2546,N_1694,N_1003);
or U2547 (N_2547,N_1111,N_1874);
nand U2548 (N_2548,N_1013,N_1753);
and U2549 (N_2549,N_1802,N_1120);
or U2550 (N_2550,N_1657,N_1548);
or U2551 (N_2551,N_1924,N_1414);
and U2552 (N_2552,N_1903,N_1135);
and U2553 (N_2553,N_1035,N_1714);
nand U2554 (N_2554,N_1782,N_1278);
and U2555 (N_2555,N_1684,N_1751);
nand U2556 (N_2556,N_1152,N_1012);
and U2557 (N_2557,N_1821,N_1401);
nor U2558 (N_2558,N_1769,N_1996);
and U2559 (N_2559,N_1174,N_1239);
or U2560 (N_2560,N_1290,N_1746);
and U2561 (N_2561,N_1145,N_1246);
and U2562 (N_2562,N_1772,N_1913);
or U2563 (N_2563,N_1468,N_1612);
nand U2564 (N_2564,N_1316,N_1398);
and U2565 (N_2565,N_1978,N_1695);
and U2566 (N_2566,N_1250,N_1831);
nand U2567 (N_2567,N_1973,N_1371);
nand U2568 (N_2568,N_1433,N_1973);
nand U2569 (N_2569,N_1440,N_1142);
nand U2570 (N_2570,N_1234,N_1522);
xnor U2571 (N_2571,N_1761,N_1183);
xor U2572 (N_2572,N_1474,N_1812);
nor U2573 (N_2573,N_1772,N_1474);
nor U2574 (N_2574,N_1687,N_1857);
xor U2575 (N_2575,N_1309,N_1333);
and U2576 (N_2576,N_1378,N_1958);
and U2577 (N_2577,N_1473,N_1765);
nor U2578 (N_2578,N_1751,N_1390);
nor U2579 (N_2579,N_1513,N_1498);
or U2580 (N_2580,N_1932,N_1758);
nand U2581 (N_2581,N_1021,N_1495);
nand U2582 (N_2582,N_1209,N_1193);
nor U2583 (N_2583,N_1314,N_1047);
and U2584 (N_2584,N_1697,N_1137);
nor U2585 (N_2585,N_1494,N_1139);
or U2586 (N_2586,N_1294,N_1253);
and U2587 (N_2587,N_1064,N_1657);
nor U2588 (N_2588,N_1610,N_1479);
nand U2589 (N_2589,N_1899,N_1846);
xor U2590 (N_2590,N_1035,N_1431);
and U2591 (N_2591,N_1981,N_1669);
nand U2592 (N_2592,N_1332,N_1254);
and U2593 (N_2593,N_1235,N_1346);
xnor U2594 (N_2594,N_1629,N_1814);
nor U2595 (N_2595,N_1627,N_1902);
and U2596 (N_2596,N_1750,N_1210);
xor U2597 (N_2597,N_1880,N_1852);
nand U2598 (N_2598,N_1000,N_1761);
and U2599 (N_2599,N_1314,N_1840);
xnor U2600 (N_2600,N_1479,N_1525);
nand U2601 (N_2601,N_1371,N_1604);
or U2602 (N_2602,N_1408,N_1869);
and U2603 (N_2603,N_1993,N_1466);
nand U2604 (N_2604,N_1879,N_1290);
xnor U2605 (N_2605,N_1986,N_1231);
and U2606 (N_2606,N_1828,N_1835);
xor U2607 (N_2607,N_1742,N_1259);
and U2608 (N_2608,N_1380,N_1317);
xnor U2609 (N_2609,N_1979,N_1378);
xor U2610 (N_2610,N_1476,N_1078);
nand U2611 (N_2611,N_1766,N_1847);
or U2612 (N_2612,N_1488,N_1644);
nand U2613 (N_2613,N_1977,N_1424);
or U2614 (N_2614,N_1907,N_1685);
nor U2615 (N_2615,N_1330,N_1765);
xor U2616 (N_2616,N_1831,N_1459);
and U2617 (N_2617,N_1381,N_1950);
nor U2618 (N_2618,N_1342,N_1964);
nor U2619 (N_2619,N_1633,N_1236);
xnor U2620 (N_2620,N_1977,N_1213);
xnor U2621 (N_2621,N_1673,N_1307);
or U2622 (N_2622,N_1549,N_1353);
and U2623 (N_2623,N_1857,N_1359);
nand U2624 (N_2624,N_1517,N_1518);
nor U2625 (N_2625,N_1212,N_1481);
and U2626 (N_2626,N_1421,N_1744);
or U2627 (N_2627,N_1981,N_1282);
or U2628 (N_2628,N_1189,N_1246);
or U2629 (N_2629,N_1542,N_1170);
and U2630 (N_2630,N_1297,N_1880);
nor U2631 (N_2631,N_1713,N_1138);
nand U2632 (N_2632,N_1001,N_1007);
nand U2633 (N_2633,N_1613,N_1985);
nor U2634 (N_2634,N_1907,N_1774);
and U2635 (N_2635,N_1873,N_1123);
nor U2636 (N_2636,N_1369,N_1447);
nand U2637 (N_2637,N_1764,N_1805);
and U2638 (N_2638,N_1431,N_1894);
or U2639 (N_2639,N_1000,N_1321);
xor U2640 (N_2640,N_1964,N_1079);
and U2641 (N_2641,N_1639,N_1804);
and U2642 (N_2642,N_1003,N_1021);
or U2643 (N_2643,N_1854,N_1969);
xor U2644 (N_2644,N_1236,N_1338);
nand U2645 (N_2645,N_1119,N_1305);
nor U2646 (N_2646,N_1685,N_1939);
and U2647 (N_2647,N_1840,N_1279);
xor U2648 (N_2648,N_1645,N_1524);
xor U2649 (N_2649,N_1727,N_1934);
xor U2650 (N_2650,N_1880,N_1709);
nor U2651 (N_2651,N_1592,N_1790);
xnor U2652 (N_2652,N_1326,N_1743);
xor U2653 (N_2653,N_1340,N_1798);
xnor U2654 (N_2654,N_1271,N_1500);
nor U2655 (N_2655,N_1916,N_1151);
or U2656 (N_2656,N_1510,N_1132);
nand U2657 (N_2657,N_1663,N_1948);
or U2658 (N_2658,N_1423,N_1291);
or U2659 (N_2659,N_1484,N_1553);
or U2660 (N_2660,N_1185,N_1812);
nor U2661 (N_2661,N_1506,N_1532);
or U2662 (N_2662,N_1020,N_1281);
and U2663 (N_2663,N_1873,N_1903);
nand U2664 (N_2664,N_1584,N_1468);
or U2665 (N_2665,N_1286,N_1913);
and U2666 (N_2666,N_1974,N_1070);
xor U2667 (N_2667,N_1655,N_1555);
and U2668 (N_2668,N_1096,N_1711);
xor U2669 (N_2669,N_1896,N_1725);
and U2670 (N_2670,N_1342,N_1230);
or U2671 (N_2671,N_1910,N_1132);
nand U2672 (N_2672,N_1075,N_1373);
nand U2673 (N_2673,N_1050,N_1562);
and U2674 (N_2674,N_1534,N_1411);
xnor U2675 (N_2675,N_1174,N_1938);
and U2676 (N_2676,N_1031,N_1408);
nor U2677 (N_2677,N_1486,N_1658);
nand U2678 (N_2678,N_1327,N_1267);
xnor U2679 (N_2679,N_1587,N_1847);
nand U2680 (N_2680,N_1674,N_1910);
nand U2681 (N_2681,N_1149,N_1005);
and U2682 (N_2682,N_1177,N_1676);
or U2683 (N_2683,N_1415,N_1731);
xor U2684 (N_2684,N_1272,N_1736);
nor U2685 (N_2685,N_1718,N_1373);
and U2686 (N_2686,N_1050,N_1819);
or U2687 (N_2687,N_1726,N_1098);
xnor U2688 (N_2688,N_1259,N_1077);
xnor U2689 (N_2689,N_1789,N_1599);
or U2690 (N_2690,N_1968,N_1190);
or U2691 (N_2691,N_1005,N_1651);
or U2692 (N_2692,N_1716,N_1079);
nor U2693 (N_2693,N_1464,N_1302);
or U2694 (N_2694,N_1164,N_1159);
xor U2695 (N_2695,N_1530,N_1070);
and U2696 (N_2696,N_1925,N_1297);
and U2697 (N_2697,N_1764,N_1351);
nand U2698 (N_2698,N_1126,N_1491);
xnor U2699 (N_2699,N_1638,N_1478);
nand U2700 (N_2700,N_1123,N_1239);
nor U2701 (N_2701,N_1966,N_1313);
and U2702 (N_2702,N_1327,N_1713);
xor U2703 (N_2703,N_1390,N_1248);
or U2704 (N_2704,N_1703,N_1163);
xnor U2705 (N_2705,N_1187,N_1292);
xnor U2706 (N_2706,N_1757,N_1050);
xnor U2707 (N_2707,N_1266,N_1078);
nand U2708 (N_2708,N_1348,N_1843);
and U2709 (N_2709,N_1983,N_1846);
nor U2710 (N_2710,N_1236,N_1486);
xor U2711 (N_2711,N_1397,N_1630);
nor U2712 (N_2712,N_1039,N_1955);
or U2713 (N_2713,N_1370,N_1280);
and U2714 (N_2714,N_1692,N_1471);
or U2715 (N_2715,N_1825,N_1242);
xnor U2716 (N_2716,N_1123,N_1606);
nor U2717 (N_2717,N_1748,N_1381);
xor U2718 (N_2718,N_1410,N_1661);
or U2719 (N_2719,N_1253,N_1439);
nor U2720 (N_2720,N_1704,N_1447);
nand U2721 (N_2721,N_1551,N_1819);
and U2722 (N_2722,N_1483,N_1099);
and U2723 (N_2723,N_1223,N_1578);
xnor U2724 (N_2724,N_1792,N_1968);
and U2725 (N_2725,N_1187,N_1499);
nand U2726 (N_2726,N_1977,N_1933);
and U2727 (N_2727,N_1559,N_1336);
and U2728 (N_2728,N_1517,N_1275);
xor U2729 (N_2729,N_1819,N_1141);
nor U2730 (N_2730,N_1709,N_1270);
or U2731 (N_2731,N_1395,N_1889);
and U2732 (N_2732,N_1528,N_1898);
and U2733 (N_2733,N_1214,N_1926);
or U2734 (N_2734,N_1676,N_1229);
xor U2735 (N_2735,N_1796,N_1205);
xnor U2736 (N_2736,N_1139,N_1527);
nor U2737 (N_2737,N_1347,N_1152);
nand U2738 (N_2738,N_1904,N_1866);
xor U2739 (N_2739,N_1206,N_1673);
xor U2740 (N_2740,N_1357,N_1366);
xnor U2741 (N_2741,N_1603,N_1563);
nand U2742 (N_2742,N_1082,N_1567);
or U2743 (N_2743,N_1656,N_1155);
and U2744 (N_2744,N_1060,N_1028);
and U2745 (N_2745,N_1042,N_1943);
xor U2746 (N_2746,N_1835,N_1938);
xnor U2747 (N_2747,N_1238,N_1454);
and U2748 (N_2748,N_1684,N_1253);
nand U2749 (N_2749,N_1351,N_1804);
nand U2750 (N_2750,N_1533,N_1272);
nor U2751 (N_2751,N_1109,N_1454);
nor U2752 (N_2752,N_1525,N_1576);
or U2753 (N_2753,N_1721,N_1216);
or U2754 (N_2754,N_1072,N_1698);
nand U2755 (N_2755,N_1141,N_1463);
nor U2756 (N_2756,N_1104,N_1443);
nor U2757 (N_2757,N_1431,N_1812);
xor U2758 (N_2758,N_1150,N_1428);
nor U2759 (N_2759,N_1250,N_1614);
and U2760 (N_2760,N_1908,N_1330);
nor U2761 (N_2761,N_1356,N_1026);
or U2762 (N_2762,N_1064,N_1055);
xnor U2763 (N_2763,N_1050,N_1904);
nor U2764 (N_2764,N_1783,N_1497);
and U2765 (N_2765,N_1025,N_1918);
or U2766 (N_2766,N_1665,N_1843);
nor U2767 (N_2767,N_1905,N_1338);
nor U2768 (N_2768,N_1272,N_1232);
or U2769 (N_2769,N_1560,N_1863);
and U2770 (N_2770,N_1608,N_1162);
nor U2771 (N_2771,N_1639,N_1909);
xor U2772 (N_2772,N_1806,N_1610);
or U2773 (N_2773,N_1344,N_1252);
nand U2774 (N_2774,N_1979,N_1200);
or U2775 (N_2775,N_1940,N_1025);
xnor U2776 (N_2776,N_1711,N_1383);
nor U2777 (N_2777,N_1572,N_1468);
nor U2778 (N_2778,N_1629,N_1747);
nand U2779 (N_2779,N_1353,N_1803);
nand U2780 (N_2780,N_1837,N_1151);
or U2781 (N_2781,N_1931,N_1180);
or U2782 (N_2782,N_1022,N_1818);
xnor U2783 (N_2783,N_1583,N_1662);
or U2784 (N_2784,N_1939,N_1696);
xnor U2785 (N_2785,N_1260,N_1949);
xor U2786 (N_2786,N_1339,N_1253);
or U2787 (N_2787,N_1336,N_1995);
nor U2788 (N_2788,N_1098,N_1214);
and U2789 (N_2789,N_1188,N_1557);
xnor U2790 (N_2790,N_1892,N_1058);
or U2791 (N_2791,N_1487,N_1560);
or U2792 (N_2792,N_1972,N_1411);
nand U2793 (N_2793,N_1276,N_1462);
nor U2794 (N_2794,N_1860,N_1974);
xor U2795 (N_2795,N_1215,N_1068);
nand U2796 (N_2796,N_1249,N_1492);
and U2797 (N_2797,N_1331,N_1444);
xnor U2798 (N_2798,N_1560,N_1519);
or U2799 (N_2799,N_1370,N_1001);
or U2800 (N_2800,N_1648,N_1894);
or U2801 (N_2801,N_1473,N_1343);
nor U2802 (N_2802,N_1303,N_1437);
xnor U2803 (N_2803,N_1713,N_1271);
and U2804 (N_2804,N_1115,N_1730);
or U2805 (N_2805,N_1001,N_1596);
nor U2806 (N_2806,N_1807,N_1253);
and U2807 (N_2807,N_1130,N_1980);
nor U2808 (N_2808,N_1520,N_1429);
xor U2809 (N_2809,N_1018,N_1141);
xnor U2810 (N_2810,N_1222,N_1242);
nor U2811 (N_2811,N_1445,N_1535);
xor U2812 (N_2812,N_1036,N_1963);
and U2813 (N_2813,N_1862,N_1789);
and U2814 (N_2814,N_1605,N_1461);
or U2815 (N_2815,N_1538,N_1517);
nand U2816 (N_2816,N_1313,N_1488);
xor U2817 (N_2817,N_1594,N_1788);
xnor U2818 (N_2818,N_1903,N_1225);
and U2819 (N_2819,N_1367,N_1916);
nand U2820 (N_2820,N_1452,N_1499);
and U2821 (N_2821,N_1722,N_1502);
or U2822 (N_2822,N_1423,N_1307);
xnor U2823 (N_2823,N_1060,N_1209);
nor U2824 (N_2824,N_1255,N_1243);
nor U2825 (N_2825,N_1950,N_1915);
and U2826 (N_2826,N_1926,N_1280);
and U2827 (N_2827,N_1348,N_1987);
or U2828 (N_2828,N_1555,N_1048);
nor U2829 (N_2829,N_1909,N_1779);
nor U2830 (N_2830,N_1231,N_1243);
xor U2831 (N_2831,N_1963,N_1116);
or U2832 (N_2832,N_1768,N_1542);
nor U2833 (N_2833,N_1484,N_1545);
xnor U2834 (N_2834,N_1325,N_1483);
nor U2835 (N_2835,N_1340,N_1992);
xnor U2836 (N_2836,N_1712,N_1725);
and U2837 (N_2837,N_1454,N_1934);
and U2838 (N_2838,N_1484,N_1939);
nand U2839 (N_2839,N_1720,N_1677);
xor U2840 (N_2840,N_1050,N_1037);
nor U2841 (N_2841,N_1054,N_1434);
nand U2842 (N_2842,N_1480,N_1571);
xor U2843 (N_2843,N_1529,N_1198);
nor U2844 (N_2844,N_1335,N_1538);
nand U2845 (N_2845,N_1997,N_1523);
nor U2846 (N_2846,N_1177,N_1223);
and U2847 (N_2847,N_1009,N_1122);
nand U2848 (N_2848,N_1688,N_1502);
or U2849 (N_2849,N_1922,N_1580);
nand U2850 (N_2850,N_1745,N_1356);
nand U2851 (N_2851,N_1983,N_1061);
xor U2852 (N_2852,N_1941,N_1997);
xnor U2853 (N_2853,N_1016,N_1897);
nor U2854 (N_2854,N_1958,N_1507);
or U2855 (N_2855,N_1102,N_1613);
nor U2856 (N_2856,N_1377,N_1826);
nor U2857 (N_2857,N_1738,N_1668);
or U2858 (N_2858,N_1010,N_1050);
or U2859 (N_2859,N_1977,N_1169);
nor U2860 (N_2860,N_1935,N_1770);
nand U2861 (N_2861,N_1304,N_1383);
nand U2862 (N_2862,N_1245,N_1261);
and U2863 (N_2863,N_1639,N_1689);
xnor U2864 (N_2864,N_1053,N_1152);
nand U2865 (N_2865,N_1098,N_1901);
or U2866 (N_2866,N_1018,N_1973);
nand U2867 (N_2867,N_1079,N_1975);
xnor U2868 (N_2868,N_1483,N_1342);
xor U2869 (N_2869,N_1263,N_1342);
nor U2870 (N_2870,N_1019,N_1503);
or U2871 (N_2871,N_1535,N_1192);
nor U2872 (N_2872,N_1388,N_1405);
nor U2873 (N_2873,N_1783,N_1084);
nor U2874 (N_2874,N_1130,N_1777);
and U2875 (N_2875,N_1450,N_1084);
nor U2876 (N_2876,N_1712,N_1471);
nor U2877 (N_2877,N_1799,N_1638);
xnor U2878 (N_2878,N_1958,N_1021);
xor U2879 (N_2879,N_1536,N_1575);
or U2880 (N_2880,N_1325,N_1598);
nand U2881 (N_2881,N_1061,N_1286);
and U2882 (N_2882,N_1303,N_1268);
nor U2883 (N_2883,N_1636,N_1316);
or U2884 (N_2884,N_1124,N_1778);
and U2885 (N_2885,N_1492,N_1446);
nor U2886 (N_2886,N_1187,N_1775);
or U2887 (N_2887,N_1240,N_1454);
xor U2888 (N_2888,N_1109,N_1844);
nor U2889 (N_2889,N_1985,N_1670);
or U2890 (N_2890,N_1578,N_1229);
xnor U2891 (N_2891,N_1700,N_1758);
and U2892 (N_2892,N_1660,N_1713);
or U2893 (N_2893,N_1769,N_1016);
and U2894 (N_2894,N_1896,N_1127);
or U2895 (N_2895,N_1536,N_1223);
or U2896 (N_2896,N_1717,N_1040);
nand U2897 (N_2897,N_1610,N_1529);
nand U2898 (N_2898,N_1455,N_1246);
nand U2899 (N_2899,N_1612,N_1530);
nand U2900 (N_2900,N_1048,N_1372);
xnor U2901 (N_2901,N_1153,N_1637);
and U2902 (N_2902,N_1281,N_1693);
nor U2903 (N_2903,N_1164,N_1068);
xnor U2904 (N_2904,N_1467,N_1402);
and U2905 (N_2905,N_1205,N_1643);
and U2906 (N_2906,N_1870,N_1352);
nand U2907 (N_2907,N_1280,N_1681);
and U2908 (N_2908,N_1399,N_1986);
xor U2909 (N_2909,N_1312,N_1302);
or U2910 (N_2910,N_1979,N_1491);
nor U2911 (N_2911,N_1592,N_1886);
xor U2912 (N_2912,N_1452,N_1703);
nand U2913 (N_2913,N_1016,N_1762);
nor U2914 (N_2914,N_1285,N_1042);
and U2915 (N_2915,N_1077,N_1992);
and U2916 (N_2916,N_1668,N_1077);
nand U2917 (N_2917,N_1101,N_1037);
or U2918 (N_2918,N_1965,N_1610);
nand U2919 (N_2919,N_1189,N_1118);
nand U2920 (N_2920,N_1585,N_1038);
and U2921 (N_2921,N_1801,N_1351);
and U2922 (N_2922,N_1137,N_1046);
or U2923 (N_2923,N_1528,N_1872);
or U2924 (N_2924,N_1757,N_1919);
and U2925 (N_2925,N_1047,N_1044);
nor U2926 (N_2926,N_1158,N_1236);
or U2927 (N_2927,N_1190,N_1400);
xnor U2928 (N_2928,N_1058,N_1021);
or U2929 (N_2929,N_1210,N_1076);
xnor U2930 (N_2930,N_1070,N_1858);
and U2931 (N_2931,N_1949,N_1894);
xnor U2932 (N_2932,N_1140,N_1667);
xor U2933 (N_2933,N_1718,N_1632);
xnor U2934 (N_2934,N_1677,N_1704);
or U2935 (N_2935,N_1429,N_1644);
nor U2936 (N_2936,N_1237,N_1964);
and U2937 (N_2937,N_1724,N_1990);
nand U2938 (N_2938,N_1474,N_1426);
nor U2939 (N_2939,N_1627,N_1037);
or U2940 (N_2940,N_1733,N_1194);
nor U2941 (N_2941,N_1933,N_1369);
or U2942 (N_2942,N_1211,N_1185);
and U2943 (N_2943,N_1707,N_1779);
or U2944 (N_2944,N_1051,N_1786);
nand U2945 (N_2945,N_1505,N_1813);
or U2946 (N_2946,N_1837,N_1091);
xnor U2947 (N_2947,N_1298,N_1424);
or U2948 (N_2948,N_1124,N_1063);
and U2949 (N_2949,N_1985,N_1388);
nor U2950 (N_2950,N_1472,N_1662);
or U2951 (N_2951,N_1898,N_1768);
nor U2952 (N_2952,N_1603,N_1437);
and U2953 (N_2953,N_1102,N_1323);
and U2954 (N_2954,N_1293,N_1230);
nand U2955 (N_2955,N_1610,N_1981);
nor U2956 (N_2956,N_1002,N_1565);
xnor U2957 (N_2957,N_1659,N_1853);
nand U2958 (N_2958,N_1788,N_1006);
and U2959 (N_2959,N_1730,N_1488);
and U2960 (N_2960,N_1739,N_1118);
nand U2961 (N_2961,N_1545,N_1006);
xor U2962 (N_2962,N_1522,N_1867);
nor U2963 (N_2963,N_1271,N_1715);
nand U2964 (N_2964,N_1375,N_1107);
or U2965 (N_2965,N_1216,N_1667);
nor U2966 (N_2966,N_1925,N_1545);
nand U2967 (N_2967,N_1623,N_1193);
nand U2968 (N_2968,N_1386,N_1366);
nor U2969 (N_2969,N_1817,N_1391);
nand U2970 (N_2970,N_1263,N_1215);
and U2971 (N_2971,N_1536,N_1892);
xnor U2972 (N_2972,N_1551,N_1441);
and U2973 (N_2973,N_1902,N_1806);
or U2974 (N_2974,N_1489,N_1178);
nor U2975 (N_2975,N_1734,N_1055);
or U2976 (N_2976,N_1223,N_1923);
and U2977 (N_2977,N_1992,N_1893);
nor U2978 (N_2978,N_1711,N_1946);
or U2979 (N_2979,N_1287,N_1705);
or U2980 (N_2980,N_1553,N_1162);
xnor U2981 (N_2981,N_1078,N_1669);
nor U2982 (N_2982,N_1422,N_1156);
nand U2983 (N_2983,N_1980,N_1878);
or U2984 (N_2984,N_1988,N_1340);
nor U2985 (N_2985,N_1342,N_1382);
and U2986 (N_2986,N_1157,N_1464);
nor U2987 (N_2987,N_1507,N_1633);
nor U2988 (N_2988,N_1179,N_1685);
nand U2989 (N_2989,N_1349,N_1814);
and U2990 (N_2990,N_1867,N_1306);
or U2991 (N_2991,N_1086,N_1792);
nand U2992 (N_2992,N_1171,N_1974);
and U2993 (N_2993,N_1307,N_1118);
xnor U2994 (N_2994,N_1503,N_1938);
and U2995 (N_2995,N_1799,N_1278);
xor U2996 (N_2996,N_1218,N_1758);
and U2997 (N_2997,N_1738,N_1148);
or U2998 (N_2998,N_1289,N_1984);
nand U2999 (N_2999,N_1975,N_1339);
nand U3000 (N_3000,N_2690,N_2194);
nand U3001 (N_3001,N_2622,N_2003);
and U3002 (N_3002,N_2243,N_2180);
and U3003 (N_3003,N_2697,N_2551);
or U3004 (N_3004,N_2525,N_2860);
and U3005 (N_3005,N_2558,N_2193);
nand U3006 (N_3006,N_2612,N_2272);
xnor U3007 (N_3007,N_2893,N_2935);
nor U3008 (N_3008,N_2317,N_2997);
and U3009 (N_3009,N_2133,N_2228);
and U3010 (N_3010,N_2237,N_2462);
nand U3011 (N_3011,N_2419,N_2465);
xor U3012 (N_3012,N_2031,N_2235);
nand U3013 (N_3013,N_2751,N_2501);
xor U3014 (N_3014,N_2882,N_2738);
and U3015 (N_3015,N_2218,N_2667);
and U3016 (N_3016,N_2873,N_2124);
or U3017 (N_3017,N_2377,N_2684);
nand U3018 (N_3018,N_2066,N_2915);
and U3019 (N_3019,N_2740,N_2723);
nor U3020 (N_3020,N_2685,N_2715);
or U3021 (N_3021,N_2301,N_2632);
nand U3022 (N_3022,N_2264,N_2028);
nor U3023 (N_3023,N_2601,N_2646);
or U3024 (N_3024,N_2511,N_2993);
or U3025 (N_3025,N_2334,N_2947);
xor U3026 (N_3026,N_2345,N_2555);
and U3027 (N_3027,N_2466,N_2870);
nor U3028 (N_3028,N_2394,N_2504);
and U3029 (N_3029,N_2531,N_2025);
and U3030 (N_3030,N_2890,N_2857);
xor U3031 (N_3031,N_2621,N_2382);
xor U3032 (N_3032,N_2770,N_2091);
nand U3033 (N_3033,N_2204,N_2426);
nor U3034 (N_3034,N_2339,N_2244);
nand U3035 (N_3035,N_2479,N_2527);
and U3036 (N_3036,N_2246,N_2005);
nor U3037 (N_3037,N_2533,N_2414);
nor U3038 (N_3038,N_2855,N_2196);
and U3039 (N_3039,N_2842,N_2027);
nor U3040 (N_3040,N_2640,N_2637);
xnor U3041 (N_3041,N_2731,N_2909);
xnor U3042 (N_3042,N_2059,N_2790);
nand U3043 (N_3043,N_2013,N_2375);
and U3044 (N_3044,N_2987,N_2129);
nand U3045 (N_3045,N_2048,N_2507);
nor U3046 (N_3046,N_2582,N_2451);
and U3047 (N_3047,N_2960,N_2432);
nand U3048 (N_3048,N_2232,N_2598);
nand U3049 (N_3049,N_2876,N_2524);
xor U3050 (N_3050,N_2696,N_2177);
nand U3051 (N_3051,N_2625,N_2729);
xnor U3052 (N_3052,N_2104,N_2087);
nand U3053 (N_3053,N_2674,N_2134);
xor U3054 (N_3054,N_2055,N_2452);
xor U3055 (N_3055,N_2403,N_2164);
xor U3056 (N_3056,N_2138,N_2242);
nand U3057 (N_3057,N_2212,N_2223);
nor U3058 (N_3058,N_2221,N_2792);
nor U3059 (N_3059,N_2672,N_2686);
or U3060 (N_3060,N_2881,N_2121);
and U3061 (N_3061,N_2398,N_2406);
xnor U3062 (N_3062,N_2768,N_2747);
nand U3063 (N_3063,N_2061,N_2284);
and U3064 (N_3064,N_2162,N_2103);
and U3065 (N_3065,N_2833,N_2594);
nor U3066 (N_3066,N_2869,N_2712);
or U3067 (N_3067,N_2024,N_2644);
or U3068 (N_3068,N_2156,N_2270);
xor U3069 (N_3069,N_2880,N_2053);
and U3070 (N_3070,N_2142,N_2757);
or U3071 (N_3071,N_2057,N_2786);
nor U3072 (N_3072,N_2919,N_2328);
nand U3073 (N_3073,N_2476,N_2969);
nor U3074 (N_3074,N_2442,N_2772);
and U3075 (N_3075,N_2811,N_2549);
nor U3076 (N_3076,N_2937,N_2559);
or U3077 (N_3077,N_2166,N_2393);
and U3078 (N_3078,N_2649,N_2175);
or U3079 (N_3079,N_2940,N_2139);
or U3080 (N_3080,N_2459,N_2314);
nand U3081 (N_3081,N_2495,N_2670);
or U3082 (N_3082,N_2972,N_2127);
nor U3083 (N_3083,N_2516,N_2930);
and U3084 (N_3084,N_2288,N_2276);
nand U3085 (N_3085,N_2841,N_2383);
and U3086 (N_3086,N_2296,N_2736);
nor U3087 (N_3087,N_2325,N_2226);
nand U3088 (N_3088,N_2349,N_2404);
or U3089 (N_3089,N_2022,N_2396);
nor U3090 (N_3090,N_2160,N_2385);
or U3091 (N_3091,N_2399,N_2407);
xor U3092 (N_3092,N_2814,N_2205);
nor U3093 (N_3093,N_2846,N_2054);
or U3094 (N_3094,N_2150,N_2081);
nand U3095 (N_3095,N_2979,N_2100);
or U3096 (N_3096,N_2645,N_2034);
nor U3097 (N_3097,N_2826,N_2460);
nor U3098 (N_3098,N_2508,N_2981);
nor U3099 (N_3099,N_2484,N_2641);
or U3100 (N_3100,N_2077,N_2974);
and U3101 (N_3101,N_2942,N_2101);
xor U3102 (N_3102,N_2793,N_2256);
nand U3103 (N_3103,N_2209,N_2887);
nand U3104 (N_3104,N_2932,N_2183);
nand U3105 (N_3105,N_2102,N_2923);
or U3106 (N_3106,N_2457,N_2105);
nand U3107 (N_3107,N_2413,N_2862);
or U3108 (N_3108,N_2963,N_2629);
nand U3109 (N_3109,N_2410,N_2119);
or U3110 (N_3110,N_2132,N_2506);
nand U3111 (N_3111,N_2176,N_2648);
xor U3112 (N_3112,N_2809,N_2191);
or U3113 (N_3113,N_2557,N_2735);
and U3114 (N_3114,N_2656,N_2560);
xor U3115 (N_3115,N_2095,N_2941);
nor U3116 (N_3116,N_2018,N_2630);
xnor U3117 (N_3117,N_2788,N_2761);
or U3118 (N_3118,N_2954,N_2838);
nand U3119 (N_3119,N_2023,N_2872);
xor U3120 (N_3120,N_2660,N_2096);
xnor U3121 (N_3121,N_2618,N_2360);
or U3122 (N_3122,N_2454,N_2519);
or U3123 (N_3123,N_2851,N_2695);
and U3124 (N_3124,N_2145,N_2707);
and U3125 (N_3125,N_2720,N_2899);
nor U3126 (N_3126,N_2845,N_2536);
or U3127 (N_3127,N_2810,N_2082);
nor U3128 (N_3128,N_2709,N_2445);
and U3129 (N_3129,N_2908,N_2900);
and U3130 (N_3130,N_2830,N_2046);
nand U3131 (N_3131,N_2812,N_2889);
or U3132 (N_3132,N_2578,N_2153);
nand U3133 (N_3133,N_2680,N_2664);
nor U3134 (N_3134,N_2203,N_2975);
and U3135 (N_3135,N_2068,N_2021);
nand U3136 (N_3136,N_2781,N_2263);
or U3137 (N_3137,N_2600,N_2198);
and U3138 (N_3138,N_2951,N_2668);
or U3139 (N_3139,N_2389,N_2688);
nor U3140 (N_3140,N_2610,N_2813);
and U3141 (N_3141,N_2624,N_2719);
and U3142 (N_3142,N_2806,N_2920);
xnor U3143 (N_3143,N_2514,N_2001);
nand U3144 (N_3144,N_2450,N_2586);
or U3145 (N_3145,N_2895,N_2224);
xnor U3146 (N_3146,N_2148,N_2269);
or U3147 (N_3147,N_2787,N_2673);
xor U3148 (N_3148,N_2936,N_2388);
xnor U3149 (N_3149,N_2173,N_2321);
nand U3150 (N_3150,N_2229,N_2602);
and U3151 (N_3151,N_2038,N_2113);
nand U3152 (N_3152,N_2779,N_2892);
and U3153 (N_3153,N_2593,N_2829);
xnor U3154 (N_3154,N_2746,N_2886);
nor U3155 (N_3155,N_2297,N_2577);
nand U3156 (N_3156,N_2480,N_2315);
nand U3157 (N_3157,N_2964,N_2361);
nand U3158 (N_3158,N_2412,N_2366);
xnor U3159 (N_3159,N_2289,N_2849);
or U3160 (N_3160,N_2550,N_2905);
nand U3161 (N_3161,N_2633,N_2710);
nor U3162 (N_3162,N_2376,N_2004);
nand U3163 (N_3163,N_2433,N_2052);
or U3164 (N_3164,N_2765,N_2523);
and U3165 (N_3165,N_2789,N_2657);
and U3166 (N_3166,N_2040,N_2293);
and U3167 (N_3167,N_2058,N_2711);
nand U3168 (N_3168,N_2647,N_2784);
nand U3169 (N_3169,N_2397,N_2340);
nor U3170 (N_3170,N_2912,N_2754);
xnor U3171 (N_3171,N_2390,N_2878);
or U3172 (N_3172,N_2918,N_2934);
or U3173 (N_3173,N_2636,N_2141);
or U3174 (N_3174,N_2090,N_2921);
xor U3175 (N_3175,N_2554,N_2439);
nor U3176 (N_3176,N_2801,N_2745);
nand U3177 (N_3177,N_2891,N_2714);
and U3178 (N_3178,N_2159,N_2853);
or U3179 (N_3179,N_2543,N_2913);
nand U3180 (N_3180,N_2035,N_2216);
nor U3181 (N_3181,N_2357,N_2009);
and U3182 (N_3182,N_2295,N_2627);
xnor U3183 (N_3183,N_2443,N_2561);
or U3184 (N_3184,N_2326,N_2883);
nand U3185 (N_3185,N_2036,N_2369);
xnor U3186 (N_3186,N_2977,N_2362);
nand U3187 (N_3187,N_2758,N_2168);
or U3188 (N_3188,N_2251,N_2780);
nor U3189 (N_3189,N_2548,N_2888);
or U3190 (N_3190,N_2755,N_2576);
nor U3191 (N_3191,N_2373,N_2992);
and U3192 (N_3192,N_2140,N_2444);
nor U3193 (N_3193,N_2497,N_2238);
nor U3194 (N_3194,N_2584,N_2236);
nand U3195 (N_3195,N_2662,N_2333);
nor U3196 (N_3196,N_2944,N_2653);
and U3197 (N_3197,N_2438,N_2347);
and U3198 (N_3198,N_2078,N_2161);
xor U3199 (N_3199,N_2303,N_2721);
or U3200 (N_3200,N_2118,N_2885);
and U3201 (N_3201,N_2737,N_2098);
and U3202 (N_3202,N_2871,N_2917);
or U3203 (N_3203,N_2374,N_2861);
xnor U3204 (N_3204,N_2771,N_2286);
nand U3205 (N_3205,N_2725,N_2202);
and U3206 (N_3206,N_2300,N_2517);
or U3207 (N_3207,N_2774,N_2565);
xor U3208 (N_3208,N_2535,N_2566);
and U3209 (N_3209,N_2130,N_2722);
and U3210 (N_3210,N_2279,N_2717);
and U3211 (N_3211,N_2453,N_2691);
nor U3212 (N_3212,N_2184,N_2512);
nand U3213 (N_3213,N_2475,N_2877);
or U3214 (N_3214,N_2687,N_2590);
xnor U3215 (N_3215,N_2967,N_2982);
nor U3216 (N_3216,N_2795,N_2778);
nor U3217 (N_3217,N_2615,N_2835);
or U3218 (N_3218,N_2631,N_2060);
nand U3219 (N_3219,N_2174,N_2227);
xor U3220 (N_3220,N_2544,N_2863);
xnor U3221 (N_3221,N_2999,N_2949);
nand U3222 (N_3222,N_2607,N_2189);
nor U3223 (N_3223,N_2694,N_2456);
nand U3224 (N_3224,N_2197,N_2014);
and U3225 (N_3225,N_2182,N_2073);
and U3226 (N_3226,N_2015,N_2430);
and U3227 (N_3227,N_2207,N_2355);
or U3228 (N_3228,N_2047,N_2989);
or U3229 (N_3229,N_2294,N_2701);
nor U3230 (N_3230,N_2875,N_2639);
or U3231 (N_3231,N_2961,N_2939);
nor U3232 (N_3232,N_2994,N_2677);
nor U3233 (N_3233,N_2225,N_2461);
or U3234 (N_3234,N_2526,N_2782);
or U3235 (N_3235,N_2856,N_2545);
and U3236 (N_3236,N_2502,N_2117);
and U3237 (N_3237,N_2492,N_2776);
xnor U3238 (N_3238,N_2663,N_2816);
nor U3239 (N_3239,N_2032,N_2946);
xnor U3240 (N_3240,N_2931,N_2352);
nor U3241 (N_3241,N_2110,N_2431);
and U3242 (N_3242,N_2386,N_2671);
nand U3243 (N_3243,N_2617,N_2332);
xnor U3244 (N_3244,N_2666,N_2580);
xnor U3245 (N_3245,N_2020,N_2570);
nor U3246 (N_3246,N_2342,N_2151);
nor U3247 (N_3247,N_2844,N_2732);
and U3248 (N_3248,N_2287,N_2706);
or U3249 (N_3249,N_2505,N_2785);
xor U3250 (N_3250,N_2429,N_2274);
xor U3251 (N_3251,N_2734,N_2319);
nand U3252 (N_3252,N_2730,N_2894);
and U3253 (N_3253,N_2820,N_2298);
nor U3254 (N_3254,N_2742,N_2115);
nand U3255 (N_3255,N_2702,N_2528);
xnor U3256 (N_3256,N_2240,N_2112);
and U3257 (N_3257,N_2190,N_2083);
or U3258 (N_3258,N_2948,N_2316);
or U3259 (N_3259,N_2773,N_2750);
xnor U3260 (N_3260,N_2356,N_2897);
xor U3261 (N_3261,N_2259,N_2655);
or U3262 (N_3262,N_2017,N_2499);
or U3263 (N_3263,N_2471,N_2614);
nor U3264 (N_3264,N_2470,N_2029);
xor U3265 (N_3265,N_2985,N_2044);
nor U3266 (N_3266,N_2000,N_2943);
nor U3267 (N_3267,N_2292,N_2998);
and U3268 (N_3268,N_2125,N_2094);
nand U3269 (N_3269,N_2039,N_2070);
nand U3270 (N_3270,N_2596,N_2135);
nand U3271 (N_3271,N_2563,N_2748);
nand U3272 (N_3272,N_2699,N_2477);
and U3273 (N_3273,N_2401,N_2111);
xor U3274 (N_3274,N_2491,N_2042);
xnor U3275 (N_3275,N_2472,N_2214);
and U3276 (N_3276,N_2831,N_2815);
nand U3277 (N_3277,N_2268,N_2489);
and U3278 (N_3278,N_2973,N_2336);
nand U3279 (N_3279,N_2344,N_2929);
nor U3280 (N_3280,N_2562,N_2458);
xor U3281 (N_3281,N_2310,N_2126);
xnor U3282 (N_3282,N_2455,N_2306);
or U3283 (N_3283,N_2217,N_2192);
nand U3284 (N_3284,N_2661,N_2143);
xnor U3285 (N_3285,N_2144,N_2309);
or U3286 (N_3286,N_2320,N_2278);
nor U3287 (N_3287,N_2916,N_2595);
and U3288 (N_3288,N_2764,N_2072);
or U3289 (N_3289,N_2265,N_2490);
nor U3290 (N_3290,N_2063,N_2966);
nor U3291 (N_3291,N_2253,N_2836);
nor U3292 (N_3292,N_2354,N_2515);
and U3293 (N_3293,N_2819,N_2800);
nor U3294 (N_3294,N_2503,N_2798);
nand U3295 (N_3295,N_2064,N_2155);
xor U3296 (N_3296,N_2137,N_2775);
nor U3297 (N_3297,N_2983,N_2417);
nand U3298 (N_3298,N_2085,N_2323);
or U3299 (N_3299,N_2409,N_2304);
nor U3300 (N_3300,N_2075,N_2724);
or U3301 (N_3301,N_2002,N_2322);
and U3302 (N_3302,N_2832,N_2449);
nor U3303 (N_3303,N_2152,N_2726);
nand U3304 (N_3304,N_2359,N_2769);
or U3305 (N_3305,N_2041,N_2107);
or U3306 (N_3306,N_2675,N_2493);
nor U3307 (N_3307,N_2950,N_2222);
and U3308 (N_3308,N_2275,N_2283);
or U3309 (N_3309,N_2006,N_2330);
and U3310 (N_3310,N_2088,N_2635);
and U3311 (N_3311,N_2827,N_2247);
nand U3312 (N_3312,N_2858,N_2791);
xor U3313 (N_3313,N_2254,N_2652);
and U3314 (N_3314,N_2571,N_2626);
and U3315 (N_3315,N_2539,N_2447);
and U3316 (N_3316,N_2441,N_2821);
or U3317 (N_3317,N_2828,N_2220);
and U3318 (N_3318,N_2307,N_2199);
nand U3319 (N_3319,N_2086,N_2329);
nand U3320 (N_3320,N_2252,N_2379);
nand U3321 (N_3321,N_2537,N_2392);
and U3322 (N_3322,N_2261,N_2708);
nor U3323 (N_3323,N_2556,N_2968);
xor U3324 (N_3324,N_2420,N_2384);
nand U3325 (N_3325,N_2604,N_2766);
nor U3326 (N_3326,N_2169,N_2370);
and U3327 (N_3327,N_2305,N_2154);
nand U3328 (N_3328,N_2171,N_2416);
xor U3329 (N_3329,N_2381,N_2350);
nand U3330 (N_3330,N_2865,N_2924);
nor U3331 (N_3331,N_2703,N_2608);
and U3332 (N_3332,N_2727,N_2464);
and U3333 (N_3333,N_2324,N_2867);
or U3334 (N_3334,N_2007,N_2638);
xor U3335 (N_3335,N_2854,N_2158);
and U3336 (N_3336,N_2693,N_2011);
nand U3337 (N_3337,N_2541,N_2233);
and U3338 (N_3338,N_2933,N_2327);
xor U3339 (N_3339,N_2898,N_2089);
or U3340 (N_3340,N_2368,N_2187);
xnor U3341 (N_3341,N_2308,N_2290);
and U3342 (N_3342,N_2230,N_2147);
nand U3343 (N_3343,N_2518,N_2213);
nand U3344 (N_3344,N_2049,N_2522);
nand U3345 (N_3345,N_2093,N_2839);
and U3346 (N_3346,N_2682,N_2753);
or U3347 (N_3347,N_2817,N_2553);
nand U3348 (N_3348,N_2658,N_2965);
nor U3349 (N_3349,N_2803,N_2030);
nand U3350 (N_3350,N_2266,N_2606);
nor U3351 (N_3351,N_2874,N_2904);
or U3352 (N_3352,N_2884,N_2683);
or U3353 (N_3353,N_2076,N_2823);
or U3354 (N_3354,N_2763,N_2642);
nand U3355 (N_3355,N_2045,N_2245);
nand U3356 (N_3356,N_2425,N_2258);
xnor U3357 (N_3357,N_2108,N_2991);
and U3358 (N_3358,N_2170,N_2911);
nor U3359 (N_3359,N_2436,N_2868);
nor U3360 (N_3360,N_2538,N_2380);
nand U3361 (N_3361,N_2760,N_2201);
nor U3362 (N_3362,N_2446,N_2372);
xnor U3363 (N_3363,N_2583,N_2603);
and U3364 (N_3364,N_2084,N_2418);
xor U3365 (N_3365,N_2713,N_2804);
and U3366 (N_3366,N_2267,N_2273);
or U3367 (N_3367,N_2097,N_2605);
xnor U3368 (N_3368,N_2976,N_2415);
and U3369 (N_3369,N_2676,N_2071);
nand U3370 (N_3370,N_2837,N_2469);
nand U3371 (N_3371,N_2338,N_2131);
and U3372 (N_3372,N_2679,N_2260);
nand U3373 (N_3373,N_2692,N_2037);
xnor U3374 (N_3374,N_2611,N_2959);
or U3375 (N_3375,N_2206,N_2179);
xor U3376 (N_3376,N_2474,N_2952);
or U3377 (N_3377,N_2850,N_2498);
and U3378 (N_3378,N_2282,N_2521);
nand U3379 (N_3379,N_2530,N_2210);
or U3380 (N_3380,N_2487,N_2423);
and U3381 (N_3381,N_2435,N_2540);
nor U3382 (N_3382,N_2579,N_2534);
xor U3383 (N_3383,N_2271,N_2542);
and U3384 (N_3384,N_2619,N_2473);
nand U3385 (N_3385,N_2185,N_2799);
nor U3386 (N_3386,N_2681,N_2689);
xnor U3387 (N_3387,N_2654,N_2777);
and U3388 (N_3388,N_2970,N_2318);
xnor U3389 (N_3389,N_2588,N_2572);
or U3390 (N_3390,N_2739,N_2313);
xor U3391 (N_3391,N_2391,N_2520);
nand U3392 (N_3392,N_2906,N_2365);
or U3393 (N_3393,N_2343,N_2552);
or U3394 (N_3394,N_2925,N_2008);
and U3395 (N_3395,N_2106,N_2592);
nor U3396 (N_3396,N_2597,N_2996);
xnor U3397 (N_3397,N_2802,N_2958);
and U3398 (N_3398,N_2099,N_2587);
xnor U3399 (N_3399,N_2822,N_2752);
or U3400 (N_3400,N_2051,N_2564);
or U3401 (N_3401,N_2080,N_2926);
or U3402 (N_3402,N_2026,N_2331);
nand U3403 (N_3403,N_2114,N_2704);
nand U3404 (N_3404,N_2749,N_2248);
xor U3405 (N_3405,N_2255,N_2585);
or U3406 (N_3406,N_2262,N_2927);
nor U3407 (N_3407,N_2718,N_2574);
nor U3408 (N_3408,N_2234,N_2762);
nor U3409 (N_3409,N_2067,N_2613);
xor U3410 (N_3410,N_2211,N_2928);
xor U3411 (N_3411,N_2043,N_2405);
or U3412 (N_3412,N_2783,N_2402);
nor U3413 (N_3413,N_2195,N_2348);
or U3414 (N_3414,N_2743,N_2852);
xnor U3415 (N_3415,N_2428,N_2529);
nor U3416 (N_3416,N_2698,N_2651);
and U3417 (N_3417,N_2866,N_2285);
nand U3418 (N_3418,N_2079,N_2033);
and U3419 (N_3419,N_2988,N_2807);
or U3420 (N_3420,N_2478,N_2488);
nor U3421 (N_3421,N_2805,N_2486);
xor U3422 (N_3422,N_2312,N_2219);
nor U3423 (N_3423,N_2280,N_2136);
nor U3424 (N_3424,N_2367,N_2157);
nand U3425 (N_3425,N_2346,N_2896);
and U3426 (N_3426,N_2188,N_2879);
nor U3427 (N_3427,N_2728,N_2840);
and U3428 (N_3428,N_2400,N_2120);
nor U3429 (N_3429,N_2434,N_2109);
or U3430 (N_3430,N_2358,N_2744);
xor U3431 (N_3431,N_2065,N_2796);
or U3432 (N_3432,N_2794,N_2953);
xnor U3433 (N_3433,N_2463,N_2149);
nor U3434 (N_3434,N_2705,N_2716);
nand U3435 (N_3435,N_2074,N_2990);
or U3436 (N_3436,N_2971,N_2957);
xnor U3437 (N_3437,N_2546,N_2902);
xor U3438 (N_3438,N_2302,N_2843);
xnor U3439 (N_3439,N_2010,N_2669);
nor U3440 (N_3440,N_2231,N_2208);
xnor U3441 (N_3441,N_2568,N_2163);
or U3442 (N_3442,N_2364,N_2468);
xor U3443 (N_3443,N_2241,N_2165);
xor U3444 (N_3444,N_2181,N_2569);
or U3445 (N_3445,N_2440,N_2547);
xnor U3446 (N_3446,N_2422,N_2494);
or U3447 (N_3447,N_2859,N_2019);
and U3448 (N_3448,N_2509,N_2995);
nand U3449 (N_3449,N_2513,N_2984);
and U3450 (N_3450,N_2250,N_2864);
nor U3451 (N_3451,N_2659,N_2277);
nand U3452 (N_3452,N_2901,N_2200);
nand U3453 (N_3453,N_2483,N_2848);
or U3454 (N_3454,N_2408,N_2467);
nor U3455 (N_3455,N_2448,N_2986);
or U3456 (N_3456,N_2481,N_2834);
nor U3457 (N_3457,N_2825,N_2589);
xnor U3458 (N_3458,N_2581,N_2922);
nor U3459 (N_3459,N_2620,N_2186);
nand U3460 (N_3460,N_2062,N_2299);
and U3461 (N_3461,N_2824,N_2411);
xor U3462 (N_3462,N_2116,N_2281);
nor U3463 (N_3463,N_2907,N_2616);
and U3464 (N_3464,N_2741,N_2634);
xnor U3465 (N_3465,N_2978,N_2938);
xor U3466 (N_3466,N_2249,N_2609);
and U3467 (N_3467,N_2575,N_2239);
or U3468 (N_3468,N_2482,N_2650);
xnor U3469 (N_3469,N_2387,N_2643);
and U3470 (N_3470,N_2337,N_2500);
and U3471 (N_3471,N_2421,N_2215);
nor U3472 (N_3472,N_2123,N_2351);
or U3473 (N_3473,N_2756,N_2122);
xnor U3474 (N_3474,N_2903,N_2311);
or U3475 (N_3475,N_2371,N_2678);
and U3476 (N_3476,N_2980,N_2573);
nand U3477 (N_3477,N_2395,N_2172);
xor U3478 (N_3478,N_2759,N_2353);
or U3479 (N_3479,N_2808,N_2146);
nand U3480 (N_3480,N_2910,N_2914);
nor U3481 (N_3481,N_2128,N_2733);
nand U3482 (N_3482,N_2178,N_2496);
xnor U3483 (N_3483,N_2167,N_2092);
xor U3484 (N_3484,N_2363,N_2012);
xnor U3485 (N_3485,N_2665,N_2378);
nand U3486 (N_3486,N_2955,N_2532);
and U3487 (N_3487,N_2510,N_2427);
or U3488 (N_3488,N_2291,N_2700);
and U3489 (N_3489,N_2567,N_2797);
nand U3490 (N_3490,N_2962,N_2628);
nor U3491 (N_3491,N_2050,N_2847);
xor U3492 (N_3492,N_2056,N_2945);
nor U3493 (N_3493,N_2424,N_2591);
or U3494 (N_3494,N_2956,N_2016);
or U3495 (N_3495,N_2257,N_2623);
nor U3496 (N_3496,N_2818,N_2485);
and U3497 (N_3497,N_2599,N_2335);
xor U3498 (N_3498,N_2437,N_2341);
or U3499 (N_3499,N_2767,N_2069);
and U3500 (N_3500,N_2503,N_2700);
nor U3501 (N_3501,N_2155,N_2689);
and U3502 (N_3502,N_2199,N_2915);
xor U3503 (N_3503,N_2355,N_2787);
nor U3504 (N_3504,N_2429,N_2513);
or U3505 (N_3505,N_2658,N_2373);
nor U3506 (N_3506,N_2643,N_2562);
or U3507 (N_3507,N_2686,N_2119);
xor U3508 (N_3508,N_2583,N_2585);
xnor U3509 (N_3509,N_2782,N_2522);
or U3510 (N_3510,N_2223,N_2235);
nor U3511 (N_3511,N_2723,N_2360);
nor U3512 (N_3512,N_2030,N_2197);
xor U3513 (N_3513,N_2622,N_2378);
nand U3514 (N_3514,N_2226,N_2266);
xor U3515 (N_3515,N_2876,N_2409);
xnor U3516 (N_3516,N_2567,N_2009);
xor U3517 (N_3517,N_2373,N_2393);
and U3518 (N_3518,N_2078,N_2526);
nor U3519 (N_3519,N_2807,N_2617);
or U3520 (N_3520,N_2692,N_2963);
or U3521 (N_3521,N_2780,N_2283);
nor U3522 (N_3522,N_2689,N_2781);
nor U3523 (N_3523,N_2607,N_2337);
and U3524 (N_3524,N_2531,N_2627);
and U3525 (N_3525,N_2011,N_2360);
xor U3526 (N_3526,N_2670,N_2256);
xor U3527 (N_3527,N_2850,N_2630);
nand U3528 (N_3528,N_2578,N_2479);
and U3529 (N_3529,N_2995,N_2399);
or U3530 (N_3530,N_2647,N_2318);
nor U3531 (N_3531,N_2876,N_2110);
nand U3532 (N_3532,N_2417,N_2877);
xor U3533 (N_3533,N_2928,N_2837);
nor U3534 (N_3534,N_2339,N_2252);
nor U3535 (N_3535,N_2674,N_2525);
and U3536 (N_3536,N_2334,N_2432);
nand U3537 (N_3537,N_2132,N_2509);
xnor U3538 (N_3538,N_2413,N_2965);
nor U3539 (N_3539,N_2489,N_2128);
xor U3540 (N_3540,N_2663,N_2128);
nand U3541 (N_3541,N_2353,N_2836);
nor U3542 (N_3542,N_2746,N_2765);
nor U3543 (N_3543,N_2899,N_2925);
and U3544 (N_3544,N_2099,N_2885);
nand U3545 (N_3545,N_2813,N_2283);
xor U3546 (N_3546,N_2191,N_2987);
nor U3547 (N_3547,N_2507,N_2913);
nand U3548 (N_3548,N_2039,N_2233);
nor U3549 (N_3549,N_2034,N_2387);
nor U3550 (N_3550,N_2369,N_2583);
nand U3551 (N_3551,N_2936,N_2544);
xor U3552 (N_3552,N_2816,N_2932);
xnor U3553 (N_3553,N_2924,N_2647);
or U3554 (N_3554,N_2151,N_2111);
xnor U3555 (N_3555,N_2857,N_2833);
or U3556 (N_3556,N_2323,N_2653);
nor U3557 (N_3557,N_2670,N_2037);
or U3558 (N_3558,N_2721,N_2350);
and U3559 (N_3559,N_2480,N_2851);
nand U3560 (N_3560,N_2586,N_2140);
and U3561 (N_3561,N_2146,N_2716);
xnor U3562 (N_3562,N_2749,N_2658);
xnor U3563 (N_3563,N_2009,N_2577);
nand U3564 (N_3564,N_2820,N_2745);
and U3565 (N_3565,N_2028,N_2301);
and U3566 (N_3566,N_2368,N_2810);
xnor U3567 (N_3567,N_2179,N_2134);
and U3568 (N_3568,N_2117,N_2449);
or U3569 (N_3569,N_2328,N_2872);
nor U3570 (N_3570,N_2318,N_2437);
and U3571 (N_3571,N_2861,N_2179);
nand U3572 (N_3572,N_2547,N_2243);
and U3573 (N_3573,N_2357,N_2339);
nor U3574 (N_3574,N_2673,N_2470);
nor U3575 (N_3575,N_2032,N_2237);
xnor U3576 (N_3576,N_2346,N_2348);
nand U3577 (N_3577,N_2796,N_2321);
or U3578 (N_3578,N_2561,N_2932);
and U3579 (N_3579,N_2750,N_2925);
xnor U3580 (N_3580,N_2538,N_2993);
or U3581 (N_3581,N_2051,N_2420);
or U3582 (N_3582,N_2768,N_2721);
and U3583 (N_3583,N_2997,N_2824);
and U3584 (N_3584,N_2026,N_2978);
and U3585 (N_3585,N_2134,N_2182);
nor U3586 (N_3586,N_2463,N_2751);
xnor U3587 (N_3587,N_2358,N_2181);
nor U3588 (N_3588,N_2485,N_2347);
or U3589 (N_3589,N_2395,N_2613);
and U3590 (N_3590,N_2196,N_2146);
nand U3591 (N_3591,N_2658,N_2351);
nor U3592 (N_3592,N_2948,N_2689);
nor U3593 (N_3593,N_2190,N_2173);
nor U3594 (N_3594,N_2288,N_2767);
or U3595 (N_3595,N_2185,N_2642);
nor U3596 (N_3596,N_2103,N_2697);
or U3597 (N_3597,N_2606,N_2859);
nor U3598 (N_3598,N_2057,N_2674);
nor U3599 (N_3599,N_2254,N_2331);
nand U3600 (N_3600,N_2020,N_2525);
nand U3601 (N_3601,N_2700,N_2835);
and U3602 (N_3602,N_2270,N_2157);
xnor U3603 (N_3603,N_2825,N_2033);
nor U3604 (N_3604,N_2228,N_2619);
nor U3605 (N_3605,N_2635,N_2349);
xnor U3606 (N_3606,N_2767,N_2286);
nand U3607 (N_3607,N_2894,N_2911);
nor U3608 (N_3608,N_2176,N_2841);
and U3609 (N_3609,N_2884,N_2857);
nand U3610 (N_3610,N_2804,N_2625);
or U3611 (N_3611,N_2522,N_2374);
xor U3612 (N_3612,N_2934,N_2728);
or U3613 (N_3613,N_2452,N_2161);
nand U3614 (N_3614,N_2475,N_2262);
or U3615 (N_3615,N_2044,N_2470);
xor U3616 (N_3616,N_2929,N_2410);
nor U3617 (N_3617,N_2955,N_2570);
or U3618 (N_3618,N_2241,N_2718);
and U3619 (N_3619,N_2416,N_2502);
xnor U3620 (N_3620,N_2740,N_2665);
xor U3621 (N_3621,N_2949,N_2386);
and U3622 (N_3622,N_2539,N_2544);
nor U3623 (N_3623,N_2656,N_2429);
nor U3624 (N_3624,N_2649,N_2730);
or U3625 (N_3625,N_2324,N_2912);
nand U3626 (N_3626,N_2529,N_2064);
xor U3627 (N_3627,N_2265,N_2013);
and U3628 (N_3628,N_2380,N_2880);
nor U3629 (N_3629,N_2022,N_2563);
or U3630 (N_3630,N_2066,N_2071);
xor U3631 (N_3631,N_2027,N_2924);
and U3632 (N_3632,N_2671,N_2049);
nand U3633 (N_3633,N_2879,N_2642);
xor U3634 (N_3634,N_2505,N_2313);
nand U3635 (N_3635,N_2636,N_2605);
nor U3636 (N_3636,N_2625,N_2169);
nand U3637 (N_3637,N_2326,N_2065);
nand U3638 (N_3638,N_2728,N_2686);
or U3639 (N_3639,N_2646,N_2369);
nand U3640 (N_3640,N_2789,N_2480);
and U3641 (N_3641,N_2491,N_2282);
or U3642 (N_3642,N_2543,N_2220);
or U3643 (N_3643,N_2976,N_2529);
nor U3644 (N_3644,N_2986,N_2690);
and U3645 (N_3645,N_2713,N_2696);
or U3646 (N_3646,N_2167,N_2628);
or U3647 (N_3647,N_2364,N_2464);
nor U3648 (N_3648,N_2391,N_2281);
nor U3649 (N_3649,N_2857,N_2024);
and U3650 (N_3650,N_2317,N_2636);
or U3651 (N_3651,N_2072,N_2627);
nand U3652 (N_3652,N_2390,N_2058);
nand U3653 (N_3653,N_2092,N_2073);
xnor U3654 (N_3654,N_2768,N_2389);
xnor U3655 (N_3655,N_2156,N_2337);
nor U3656 (N_3656,N_2741,N_2832);
and U3657 (N_3657,N_2876,N_2379);
xor U3658 (N_3658,N_2202,N_2976);
nor U3659 (N_3659,N_2316,N_2352);
and U3660 (N_3660,N_2626,N_2763);
xor U3661 (N_3661,N_2504,N_2293);
or U3662 (N_3662,N_2036,N_2038);
and U3663 (N_3663,N_2720,N_2965);
nand U3664 (N_3664,N_2347,N_2648);
or U3665 (N_3665,N_2419,N_2642);
xor U3666 (N_3666,N_2063,N_2843);
xnor U3667 (N_3667,N_2765,N_2445);
nor U3668 (N_3668,N_2743,N_2808);
nand U3669 (N_3669,N_2826,N_2027);
and U3670 (N_3670,N_2946,N_2996);
nand U3671 (N_3671,N_2318,N_2377);
or U3672 (N_3672,N_2233,N_2072);
or U3673 (N_3673,N_2435,N_2202);
nand U3674 (N_3674,N_2772,N_2122);
and U3675 (N_3675,N_2700,N_2255);
nand U3676 (N_3676,N_2536,N_2126);
nor U3677 (N_3677,N_2681,N_2531);
nand U3678 (N_3678,N_2689,N_2300);
and U3679 (N_3679,N_2321,N_2880);
and U3680 (N_3680,N_2910,N_2532);
xnor U3681 (N_3681,N_2039,N_2177);
xnor U3682 (N_3682,N_2950,N_2960);
and U3683 (N_3683,N_2339,N_2152);
and U3684 (N_3684,N_2400,N_2074);
xor U3685 (N_3685,N_2780,N_2923);
xor U3686 (N_3686,N_2880,N_2147);
nand U3687 (N_3687,N_2950,N_2123);
or U3688 (N_3688,N_2980,N_2516);
xor U3689 (N_3689,N_2807,N_2202);
or U3690 (N_3690,N_2948,N_2772);
nor U3691 (N_3691,N_2072,N_2790);
nor U3692 (N_3692,N_2899,N_2454);
nand U3693 (N_3693,N_2046,N_2858);
xor U3694 (N_3694,N_2177,N_2434);
and U3695 (N_3695,N_2322,N_2359);
nor U3696 (N_3696,N_2115,N_2285);
and U3697 (N_3697,N_2112,N_2472);
and U3698 (N_3698,N_2740,N_2994);
or U3699 (N_3699,N_2150,N_2471);
xor U3700 (N_3700,N_2722,N_2562);
and U3701 (N_3701,N_2547,N_2062);
xor U3702 (N_3702,N_2618,N_2167);
xor U3703 (N_3703,N_2866,N_2225);
nand U3704 (N_3704,N_2848,N_2861);
nand U3705 (N_3705,N_2766,N_2683);
or U3706 (N_3706,N_2646,N_2293);
xnor U3707 (N_3707,N_2208,N_2915);
or U3708 (N_3708,N_2300,N_2112);
or U3709 (N_3709,N_2075,N_2255);
or U3710 (N_3710,N_2120,N_2983);
or U3711 (N_3711,N_2703,N_2656);
xnor U3712 (N_3712,N_2176,N_2853);
xnor U3713 (N_3713,N_2341,N_2703);
nor U3714 (N_3714,N_2150,N_2817);
nand U3715 (N_3715,N_2066,N_2841);
xor U3716 (N_3716,N_2386,N_2216);
or U3717 (N_3717,N_2555,N_2869);
nor U3718 (N_3718,N_2932,N_2291);
and U3719 (N_3719,N_2382,N_2001);
and U3720 (N_3720,N_2455,N_2503);
nor U3721 (N_3721,N_2737,N_2902);
and U3722 (N_3722,N_2483,N_2205);
nand U3723 (N_3723,N_2233,N_2809);
xnor U3724 (N_3724,N_2514,N_2521);
nor U3725 (N_3725,N_2569,N_2502);
nor U3726 (N_3726,N_2481,N_2371);
or U3727 (N_3727,N_2707,N_2228);
xor U3728 (N_3728,N_2137,N_2501);
nor U3729 (N_3729,N_2671,N_2871);
nor U3730 (N_3730,N_2029,N_2161);
nor U3731 (N_3731,N_2838,N_2302);
and U3732 (N_3732,N_2605,N_2973);
or U3733 (N_3733,N_2002,N_2487);
nor U3734 (N_3734,N_2569,N_2735);
xnor U3735 (N_3735,N_2842,N_2246);
nand U3736 (N_3736,N_2982,N_2979);
and U3737 (N_3737,N_2688,N_2523);
or U3738 (N_3738,N_2047,N_2019);
nor U3739 (N_3739,N_2082,N_2517);
and U3740 (N_3740,N_2055,N_2564);
or U3741 (N_3741,N_2519,N_2916);
xnor U3742 (N_3742,N_2440,N_2073);
and U3743 (N_3743,N_2609,N_2723);
or U3744 (N_3744,N_2567,N_2433);
xnor U3745 (N_3745,N_2976,N_2768);
or U3746 (N_3746,N_2317,N_2702);
xor U3747 (N_3747,N_2574,N_2497);
nor U3748 (N_3748,N_2262,N_2345);
nor U3749 (N_3749,N_2744,N_2150);
and U3750 (N_3750,N_2245,N_2588);
nand U3751 (N_3751,N_2909,N_2642);
or U3752 (N_3752,N_2872,N_2821);
or U3753 (N_3753,N_2238,N_2471);
nand U3754 (N_3754,N_2167,N_2360);
or U3755 (N_3755,N_2566,N_2933);
nand U3756 (N_3756,N_2750,N_2318);
or U3757 (N_3757,N_2918,N_2336);
nand U3758 (N_3758,N_2082,N_2265);
xor U3759 (N_3759,N_2116,N_2235);
nor U3760 (N_3760,N_2279,N_2086);
xor U3761 (N_3761,N_2878,N_2958);
nor U3762 (N_3762,N_2067,N_2701);
nor U3763 (N_3763,N_2760,N_2510);
nand U3764 (N_3764,N_2079,N_2559);
nand U3765 (N_3765,N_2083,N_2650);
and U3766 (N_3766,N_2853,N_2278);
nand U3767 (N_3767,N_2088,N_2249);
and U3768 (N_3768,N_2008,N_2705);
nor U3769 (N_3769,N_2916,N_2447);
and U3770 (N_3770,N_2567,N_2168);
or U3771 (N_3771,N_2810,N_2755);
and U3772 (N_3772,N_2486,N_2686);
nor U3773 (N_3773,N_2278,N_2471);
nor U3774 (N_3774,N_2208,N_2014);
nor U3775 (N_3775,N_2131,N_2947);
or U3776 (N_3776,N_2447,N_2050);
nor U3777 (N_3777,N_2099,N_2780);
and U3778 (N_3778,N_2519,N_2194);
or U3779 (N_3779,N_2692,N_2544);
xnor U3780 (N_3780,N_2092,N_2910);
and U3781 (N_3781,N_2778,N_2123);
nor U3782 (N_3782,N_2029,N_2109);
nor U3783 (N_3783,N_2169,N_2039);
or U3784 (N_3784,N_2318,N_2348);
xnor U3785 (N_3785,N_2012,N_2836);
or U3786 (N_3786,N_2811,N_2469);
xnor U3787 (N_3787,N_2088,N_2143);
xor U3788 (N_3788,N_2037,N_2880);
nand U3789 (N_3789,N_2578,N_2133);
nand U3790 (N_3790,N_2158,N_2738);
nor U3791 (N_3791,N_2771,N_2135);
xnor U3792 (N_3792,N_2833,N_2558);
and U3793 (N_3793,N_2007,N_2285);
xnor U3794 (N_3794,N_2402,N_2077);
and U3795 (N_3795,N_2056,N_2055);
or U3796 (N_3796,N_2486,N_2085);
xnor U3797 (N_3797,N_2765,N_2766);
and U3798 (N_3798,N_2463,N_2690);
and U3799 (N_3799,N_2980,N_2723);
nand U3800 (N_3800,N_2154,N_2031);
and U3801 (N_3801,N_2481,N_2465);
xor U3802 (N_3802,N_2017,N_2794);
and U3803 (N_3803,N_2576,N_2081);
nand U3804 (N_3804,N_2253,N_2869);
and U3805 (N_3805,N_2867,N_2406);
nor U3806 (N_3806,N_2080,N_2697);
or U3807 (N_3807,N_2251,N_2924);
nand U3808 (N_3808,N_2479,N_2220);
nand U3809 (N_3809,N_2244,N_2209);
xnor U3810 (N_3810,N_2127,N_2070);
nand U3811 (N_3811,N_2619,N_2359);
xnor U3812 (N_3812,N_2367,N_2046);
or U3813 (N_3813,N_2506,N_2597);
or U3814 (N_3814,N_2722,N_2040);
nand U3815 (N_3815,N_2922,N_2324);
or U3816 (N_3816,N_2714,N_2894);
nand U3817 (N_3817,N_2992,N_2310);
xor U3818 (N_3818,N_2843,N_2653);
and U3819 (N_3819,N_2584,N_2047);
and U3820 (N_3820,N_2854,N_2172);
nand U3821 (N_3821,N_2741,N_2334);
xor U3822 (N_3822,N_2267,N_2182);
xor U3823 (N_3823,N_2991,N_2950);
and U3824 (N_3824,N_2486,N_2723);
xnor U3825 (N_3825,N_2496,N_2713);
or U3826 (N_3826,N_2208,N_2517);
nand U3827 (N_3827,N_2579,N_2256);
xor U3828 (N_3828,N_2959,N_2239);
or U3829 (N_3829,N_2489,N_2870);
xnor U3830 (N_3830,N_2367,N_2114);
or U3831 (N_3831,N_2140,N_2323);
or U3832 (N_3832,N_2876,N_2950);
xor U3833 (N_3833,N_2171,N_2075);
and U3834 (N_3834,N_2352,N_2456);
and U3835 (N_3835,N_2802,N_2050);
or U3836 (N_3836,N_2078,N_2624);
or U3837 (N_3837,N_2759,N_2950);
nor U3838 (N_3838,N_2113,N_2747);
xor U3839 (N_3839,N_2286,N_2053);
or U3840 (N_3840,N_2019,N_2856);
nor U3841 (N_3841,N_2848,N_2462);
and U3842 (N_3842,N_2671,N_2024);
and U3843 (N_3843,N_2270,N_2563);
nor U3844 (N_3844,N_2445,N_2760);
or U3845 (N_3845,N_2902,N_2246);
nand U3846 (N_3846,N_2162,N_2762);
nor U3847 (N_3847,N_2403,N_2161);
xnor U3848 (N_3848,N_2927,N_2184);
or U3849 (N_3849,N_2647,N_2482);
nor U3850 (N_3850,N_2450,N_2621);
and U3851 (N_3851,N_2272,N_2114);
or U3852 (N_3852,N_2805,N_2748);
or U3853 (N_3853,N_2223,N_2038);
nor U3854 (N_3854,N_2650,N_2548);
or U3855 (N_3855,N_2192,N_2302);
and U3856 (N_3856,N_2600,N_2055);
nor U3857 (N_3857,N_2464,N_2002);
xnor U3858 (N_3858,N_2932,N_2463);
xnor U3859 (N_3859,N_2006,N_2069);
nor U3860 (N_3860,N_2419,N_2254);
nand U3861 (N_3861,N_2957,N_2183);
xor U3862 (N_3862,N_2963,N_2550);
and U3863 (N_3863,N_2760,N_2948);
and U3864 (N_3864,N_2699,N_2934);
xor U3865 (N_3865,N_2572,N_2072);
or U3866 (N_3866,N_2990,N_2161);
nor U3867 (N_3867,N_2807,N_2307);
or U3868 (N_3868,N_2256,N_2545);
nor U3869 (N_3869,N_2495,N_2790);
nor U3870 (N_3870,N_2837,N_2069);
xnor U3871 (N_3871,N_2932,N_2811);
nand U3872 (N_3872,N_2014,N_2251);
and U3873 (N_3873,N_2748,N_2927);
nor U3874 (N_3874,N_2257,N_2139);
nand U3875 (N_3875,N_2938,N_2264);
xor U3876 (N_3876,N_2963,N_2395);
or U3877 (N_3877,N_2160,N_2581);
or U3878 (N_3878,N_2030,N_2817);
nor U3879 (N_3879,N_2205,N_2610);
and U3880 (N_3880,N_2433,N_2978);
nand U3881 (N_3881,N_2994,N_2597);
and U3882 (N_3882,N_2956,N_2950);
and U3883 (N_3883,N_2185,N_2177);
and U3884 (N_3884,N_2916,N_2749);
or U3885 (N_3885,N_2050,N_2249);
and U3886 (N_3886,N_2121,N_2317);
nand U3887 (N_3887,N_2013,N_2505);
and U3888 (N_3888,N_2998,N_2393);
nor U3889 (N_3889,N_2635,N_2373);
nor U3890 (N_3890,N_2404,N_2908);
xor U3891 (N_3891,N_2086,N_2526);
nand U3892 (N_3892,N_2977,N_2031);
nor U3893 (N_3893,N_2175,N_2849);
and U3894 (N_3894,N_2983,N_2121);
xor U3895 (N_3895,N_2439,N_2770);
or U3896 (N_3896,N_2237,N_2047);
and U3897 (N_3897,N_2120,N_2748);
xor U3898 (N_3898,N_2661,N_2663);
nand U3899 (N_3899,N_2558,N_2128);
or U3900 (N_3900,N_2502,N_2619);
xnor U3901 (N_3901,N_2381,N_2642);
nor U3902 (N_3902,N_2119,N_2931);
and U3903 (N_3903,N_2848,N_2922);
and U3904 (N_3904,N_2775,N_2766);
xnor U3905 (N_3905,N_2036,N_2785);
xor U3906 (N_3906,N_2012,N_2760);
and U3907 (N_3907,N_2936,N_2693);
xnor U3908 (N_3908,N_2594,N_2232);
xnor U3909 (N_3909,N_2748,N_2152);
xnor U3910 (N_3910,N_2467,N_2907);
nor U3911 (N_3911,N_2433,N_2130);
nor U3912 (N_3912,N_2765,N_2692);
or U3913 (N_3913,N_2923,N_2476);
nor U3914 (N_3914,N_2684,N_2418);
nand U3915 (N_3915,N_2814,N_2176);
xor U3916 (N_3916,N_2665,N_2844);
and U3917 (N_3917,N_2725,N_2360);
and U3918 (N_3918,N_2676,N_2274);
xnor U3919 (N_3919,N_2869,N_2050);
or U3920 (N_3920,N_2854,N_2247);
xnor U3921 (N_3921,N_2520,N_2599);
or U3922 (N_3922,N_2750,N_2147);
nor U3923 (N_3923,N_2724,N_2212);
and U3924 (N_3924,N_2599,N_2112);
nor U3925 (N_3925,N_2845,N_2759);
xor U3926 (N_3926,N_2174,N_2581);
and U3927 (N_3927,N_2791,N_2333);
nand U3928 (N_3928,N_2949,N_2212);
xor U3929 (N_3929,N_2329,N_2308);
nand U3930 (N_3930,N_2759,N_2750);
or U3931 (N_3931,N_2515,N_2940);
nand U3932 (N_3932,N_2981,N_2827);
nor U3933 (N_3933,N_2290,N_2667);
or U3934 (N_3934,N_2867,N_2475);
and U3935 (N_3935,N_2494,N_2217);
and U3936 (N_3936,N_2125,N_2017);
and U3937 (N_3937,N_2196,N_2780);
nand U3938 (N_3938,N_2507,N_2859);
and U3939 (N_3939,N_2847,N_2205);
nor U3940 (N_3940,N_2560,N_2473);
nor U3941 (N_3941,N_2712,N_2299);
nand U3942 (N_3942,N_2607,N_2673);
nand U3943 (N_3943,N_2277,N_2801);
and U3944 (N_3944,N_2495,N_2822);
xnor U3945 (N_3945,N_2606,N_2279);
or U3946 (N_3946,N_2711,N_2429);
nor U3947 (N_3947,N_2845,N_2473);
nand U3948 (N_3948,N_2755,N_2811);
nand U3949 (N_3949,N_2351,N_2920);
nand U3950 (N_3950,N_2041,N_2584);
nand U3951 (N_3951,N_2158,N_2270);
and U3952 (N_3952,N_2808,N_2584);
and U3953 (N_3953,N_2581,N_2950);
or U3954 (N_3954,N_2867,N_2167);
nand U3955 (N_3955,N_2979,N_2909);
xor U3956 (N_3956,N_2412,N_2788);
or U3957 (N_3957,N_2350,N_2704);
and U3958 (N_3958,N_2058,N_2054);
xor U3959 (N_3959,N_2947,N_2151);
xor U3960 (N_3960,N_2771,N_2952);
and U3961 (N_3961,N_2095,N_2675);
nand U3962 (N_3962,N_2625,N_2548);
or U3963 (N_3963,N_2108,N_2871);
or U3964 (N_3964,N_2529,N_2128);
nor U3965 (N_3965,N_2909,N_2934);
xor U3966 (N_3966,N_2024,N_2974);
nand U3967 (N_3967,N_2515,N_2134);
xor U3968 (N_3968,N_2862,N_2089);
xnor U3969 (N_3969,N_2699,N_2408);
and U3970 (N_3970,N_2721,N_2059);
nand U3971 (N_3971,N_2765,N_2912);
xnor U3972 (N_3972,N_2543,N_2556);
or U3973 (N_3973,N_2239,N_2359);
nor U3974 (N_3974,N_2219,N_2721);
and U3975 (N_3975,N_2295,N_2434);
or U3976 (N_3976,N_2357,N_2140);
nor U3977 (N_3977,N_2707,N_2954);
and U3978 (N_3978,N_2479,N_2004);
nor U3979 (N_3979,N_2014,N_2455);
nor U3980 (N_3980,N_2903,N_2076);
xor U3981 (N_3981,N_2941,N_2228);
and U3982 (N_3982,N_2154,N_2472);
and U3983 (N_3983,N_2362,N_2689);
xnor U3984 (N_3984,N_2555,N_2482);
xnor U3985 (N_3985,N_2336,N_2798);
and U3986 (N_3986,N_2593,N_2626);
nand U3987 (N_3987,N_2412,N_2336);
and U3988 (N_3988,N_2896,N_2398);
nor U3989 (N_3989,N_2841,N_2537);
nand U3990 (N_3990,N_2057,N_2384);
and U3991 (N_3991,N_2516,N_2330);
nand U3992 (N_3992,N_2778,N_2931);
and U3993 (N_3993,N_2368,N_2597);
and U3994 (N_3994,N_2883,N_2716);
nand U3995 (N_3995,N_2584,N_2335);
xor U3996 (N_3996,N_2824,N_2505);
and U3997 (N_3997,N_2309,N_2414);
and U3998 (N_3998,N_2688,N_2500);
nor U3999 (N_3999,N_2279,N_2553);
nand U4000 (N_4000,N_3210,N_3844);
xor U4001 (N_4001,N_3868,N_3055);
nand U4002 (N_4002,N_3684,N_3119);
and U4003 (N_4003,N_3607,N_3577);
nand U4004 (N_4004,N_3826,N_3947);
or U4005 (N_4005,N_3489,N_3647);
nor U4006 (N_4006,N_3340,N_3061);
xor U4007 (N_4007,N_3729,N_3120);
xor U4008 (N_4008,N_3566,N_3394);
or U4009 (N_4009,N_3455,N_3905);
or U4010 (N_4010,N_3057,N_3374);
or U4011 (N_4011,N_3078,N_3346);
nor U4012 (N_4012,N_3580,N_3322);
and U4013 (N_4013,N_3658,N_3679);
nand U4014 (N_4014,N_3353,N_3629);
xnor U4015 (N_4015,N_3081,N_3895);
xnor U4016 (N_4016,N_3595,N_3156);
nor U4017 (N_4017,N_3635,N_3225);
nor U4018 (N_4018,N_3857,N_3750);
nand U4019 (N_4019,N_3508,N_3253);
nor U4020 (N_4020,N_3759,N_3646);
nor U4021 (N_4021,N_3415,N_3421);
nor U4022 (N_4022,N_3591,N_3468);
nor U4023 (N_4023,N_3674,N_3029);
and U4024 (N_4024,N_3632,N_3609);
nor U4025 (N_4025,N_3644,N_3515);
and U4026 (N_4026,N_3960,N_3027);
xor U4027 (N_4027,N_3981,N_3720);
nor U4028 (N_4028,N_3323,N_3086);
xnor U4029 (N_4029,N_3689,N_3973);
and U4030 (N_4030,N_3196,N_3224);
xnor U4031 (N_4031,N_3446,N_3083);
nand U4032 (N_4032,N_3882,N_3276);
or U4033 (N_4033,N_3259,N_3856);
xor U4034 (N_4034,N_3706,N_3915);
and U4035 (N_4035,N_3971,N_3033);
or U4036 (N_4036,N_3069,N_3418);
or U4037 (N_4037,N_3718,N_3157);
and U4038 (N_4038,N_3830,N_3552);
nor U4039 (N_4039,N_3479,N_3834);
and U4040 (N_4040,N_3953,N_3603);
or U4041 (N_4041,N_3496,N_3265);
nor U4042 (N_4042,N_3889,N_3139);
or U4043 (N_4043,N_3713,N_3954);
or U4044 (N_4044,N_3885,N_3306);
xnor U4045 (N_4045,N_3672,N_3762);
or U4046 (N_4046,N_3972,N_3929);
nand U4047 (N_4047,N_3664,N_3575);
or U4048 (N_4048,N_3443,N_3964);
and U4049 (N_4049,N_3336,N_3803);
or U4050 (N_4050,N_3622,N_3187);
or U4051 (N_4051,N_3652,N_3748);
and U4052 (N_4052,N_3553,N_3533);
nor U4053 (N_4053,N_3425,N_3153);
xor U4054 (N_4054,N_3653,N_3104);
and U4055 (N_4055,N_3420,N_3484);
and U4056 (N_4056,N_3760,N_3270);
nor U4057 (N_4057,N_3526,N_3648);
and U4058 (N_4058,N_3736,N_3463);
nand U4059 (N_4059,N_3093,N_3459);
nor U4060 (N_4060,N_3813,N_3890);
nor U4061 (N_4061,N_3843,N_3944);
nor U4062 (N_4062,N_3475,N_3962);
or U4063 (N_4063,N_3114,N_3606);
nor U4064 (N_4064,N_3507,N_3053);
nand U4065 (N_4065,N_3631,N_3516);
or U4066 (N_4066,N_3481,N_3619);
xor U4067 (N_4067,N_3556,N_3778);
nor U4068 (N_4068,N_3918,N_3182);
nor U4069 (N_4069,N_3339,N_3867);
nand U4070 (N_4070,N_3151,N_3669);
or U4071 (N_4071,N_3390,N_3135);
and U4072 (N_4072,N_3872,N_3583);
xor U4073 (N_4073,N_3103,N_3744);
xor U4074 (N_4074,N_3492,N_3290);
or U4075 (N_4075,N_3095,N_3261);
nor U4076 (N_4076,N_3520,N_3164);
nor U4077 (N_4077,N_3593,N_3561);
xnor U4078 (N_4078,N_3535,N_3544);
or U4079 (N_4079,N_3710,N_3796);
or U4080 (N_4080,N_3232,N_3304);
nor U4081 (N_4081,N_3839,N_3454);
or U4082 (N_4082,N_3649,N_3949);
nor U4083 (N_4083,N_3248,N_3350);
xnor U4084 (N_4084,N_3916,N_3431);
and U4085 (N_4085,N_3138,N_3023);
or U4086 (N_4086,N_3274,N_3866);
nand U4087 (N_4087,N_3026,N_3783);
nor U4088 (N_4088,N_3123,N_3959);
or U4089 (N_4089,N_3324,N_3747);
and U4090 (N_4090,N_3943,N_3117);
nor U4091 (N_4091,N_3140,N_3766);
nor U4092 (N_4092,N_3465,N_3541);
nor U4093 (N_4093,N_3392,N_3931);
nand U4094 (N_4094,N_3467,N_3560);
xnor U4095 (N_4095,N_3036,N_3227);
nand U4096 (N_4096,N_3342,N_3220);
xor U4097 (N_4097,N_3293,N_3850);
nor U4098 (N_4098,N_3877,N_3006);
or U4099 (N_4099,N_3297,N_3189);
and U4100 (N_4100,N_3945,N_3537);
nor U4101 (N_4101,N_3016,N_3773);
nand U4102 (N_4102,N_3230,N_3473);
and U4103 (N_4103,N_3772,N_3690);
nand U4104 (N_4104,N_3205,N_3510);
or U4105 (N_4105,N_3474,N_3377);
nand U4106 (N_4106,N_3173,N_3574);
xor U4107 (N_4107,N_3133,N_3318);
or U4108 (N_4108,N_3371,N_3438);
nor U4109 (N_4109,N_3605,N_3070);
nand U4110 (N_4110,N_3709,N_3416);
or U4111 (N_4111,N_3052,N_3291);
nand U4112 (N_4112,N_3343,N_3321);
nor U4113 (N_4113,N_3651,N_3495);
and U4114 (N_4114,N_3875,N_3251);
or U4115 (N_4115,N_3208,N_3222);
xnor U4116 (N_4116,N_3327,N_3207);
nor U4117 (N_4117,N_3673,N_3243);
nand U4118 (N_4118,N_3845,N_3968);
nand U4119 (N_4119,N_3922,N_3848);
nand U4120 (N_4120,N_3693,N_3668);
nand U4121 (N_4121,N_3966,N_3511);
or U4122 (N_4122,N_3010,N_3751);
nor U4123 (N_4123,N_3166,N_3235);
nand U4124 (N_4124,N_3776,N_3501);
nand U4125 (N_4125,N_3578,N_3121);
nor U4126 (N_4126,N_3469,N_3218);
nand U4127 (N_4127,N_3989,N_3988);
and U4128 (N_4128,N_3787,N_3209);
nand U4129 (N_4129,N_3798,N_3302);
xor U4130 (N_4130,N_3847,N_3381);
xor U4131 (N_4131,N_3045,N_3999);
nand U4132 (N_4132,N_3099,N_3247);
and U4133 (N_4133,N_3047,N_3723);
nand U4134 (N_4134,N_3129,N_3433);
nand U4135 (N_4135,N_3005,N_3965);
nor U4136 (N_4136,N_3414,N_3997);
xnor U4137 (N_4137,N_3044,N_3543);
nand U4138 (N_4138,N_3170,N_3429);
or U4139 (N_4139,N_3190,N_3660);
xor U4140 (N_4140,N_3065,N_3816);
or U4141 (N_4141,N_3345,N_3733);
or U4142 (N_4142,N_3017,N_3466);
nand U4143 (N_4143,N_3800,N_3172);
xnor U4144 (N_4144,N_3058,N_3912);
or U4145 (N_4145,N_3464,N_3852);
and U4146 (N_4146,N_3478,N_3775);
or U4147 (N_4147,N_3849,N_3814);
xor U4148 (N_4148,N_3871,N_3528);
nor U4149 (N_4149,N_3162,N_3077);
or U4150 (N_4150,N_3941,N_3946);
xnor U4151 (N_4151,N_3623,N_3639);
nor U4152 (N_4152,N_3366,N_3245);
xnor U4153 (N_4153,N_3558,N_3899);
xnor U4154 (N_4154,N_3785,N_3487);
nand U4155 (N_4155,N_3236,N_3211);
nand U4156 (N_4156,N_3493,N_3665);
nand U4157 (N_4157,N_3832,N_3254);
and U4158 (N_4158,N_3793,N_3289);
xnor U4159 (N_4159,N_3958,N_3328);
and U4160 (N_4160,N_3881,N_3432);
nor U4161 (N_4161,N_3280,N_3488);
and U4162 (N_4162,N_3483,N_3695);
nor U4163 (N_4163,N_3035,N_3676);
nand U4164 (N_4164,N_3296,N_3707);
or U4165 (N_4165,N_3716,N_3627);
nand U4166 (N_4166,N_3268,N_3934);
or U4167 (N_4167,N_3400,N_3616);
and U4168 (N_4168,N_3378,N_3801);
xor U4169 (N_4169,N_3907,N_3952);
nand U4170 (N_4170,N_3891,N_3364);
nand U4171 (N_4171,N_3184,N_3592);
and U4172 (N_4172,N_3539,N_3192);
nor U4173 (N_4173,N_3150,N_3191);
and U4174 (N_4174,N_3898,N_3092);
xor U4175 (N_4175,N_3074,N_3795);
nor U4176 (N_4176,N_3011,N_3283);
nand U4177 (N_4177,N_3549,N_3115);
or U4178 (N_4178,N_3435,N_3909);
xor U4179 (N_4179,N_3084,N_3441);
and U4180 (N_4180,N_3870,N_3292);
and U4181 (N_4181,N_3611,N_3951);
nor U4182 (N_4182,N_3079,N_3360);
xor U4183 (N_4183,N_3049,N_3688);
and U4184 (N_4184,N_3050,N_3383);
and U4185 (N_4185,N_3538,N_3835);
and U4186 (N_4186,N_3348,N_3329);
nor U4187 (N_4187,N_3264,N_3417);
and U4188 (N_4188,N_3199,N_3223);
nand U4189 (N_4189,N_3137,N_3066);
xnor U4190 (N_4190,N_3085,N_3376);
nor U4191 (N_4191,N_3731,N_3317);
and U4192 (N_4192,N_3942,N_3682);
or U4193 (N_4193,N_3337,N_3820);
xor U4194 (N_4194,N_3708,N_3503);
nand U4195 (N_4195,N_3012,N_3613);
and U4196 (N_4196,N_3691,N_3216);
xnor U4197 (N_4197,N_3320,N_3094);
nor U4198 (N_4198,N_3308,N_3048);
or U4199 (N_4199,N_3132,N_3221);
or U4200 (N_4200,N_3054,N_3822);
nor U4201 (N_4201,N_3449,N_3779);
xnor U4202 (N_4202,N_3836,N_3699);
xor U4203 (N_4203,N_3249,N_3740);
xor U4204 (N_4204,N_3703,N_3263);
nand U4205 (N_4205,N_3453,N_3357);
xor U4206 (N_4206,N_3039,N_3018);
xor U4207 (N_4207,N_3024,N_3457);
or U4208 (N_4208,N_3542,N_3145);
nand U4209 (N_4209,N_3349,N_3331);
xor U4210 (N_4210,N_3124,N_3257);
and U4211 (N_4211,N_3309,N_3600);
and U4212 (N_4212,N_3734,N_3098);
and U4213 (N_4213,N_3112,N_3358);
or U4214 (N_4214,N_3677,N_3313);
and U4215 (N_4215,N_3799,N_3565);
or U4216 (N_4216,N_3266,N_3788);
xnor U4217 (N_4217,N_3697,N_3101);
or U4218 (N_4218,N_3728,N_3186);
nor U4219 (N_4219,N_3823,N_3064);
and U4220 (N_4220,N_3448,N_3683);
or U4221 (N_4221,N_3303,N_3957);
and U4222 (N_4222,N_3940,N_3534);
or U4223 (N_4223,N_3754,N_3900);
nand U4224 (N_4224,N_3926,N_3105);
xor U4225 (N_4225,N_3332,N_3874);
and U4226 (N_4226,N_3752,N_3144);
nor U4227 (N_4227,N_3702,N_3923);
nor U4228 (N_4228,N_3128,N_3146);
nand U4229 (N_4229,N_3147,N_3051);
and U4230 (N_4230,N_3524,N_3768);
and U4231 (N_4231,N_3424,N_3601);
nor U4232 (N_4232,N_3821,N_3531);
xor U4233 (N_4233,N_3833,N_3919);
or U4234 (N_4234,N_3384,N_3726);
or U4235 (N_4235,N_3599,N_3628);
or U4236 (N_4236,N_3618,N_3073);
xor U4237 (N_4237,N_3271,N_3305);
xnor U4238 (N_4238,N_3131,N_3260);
xor U4239 (N_4239,N_3091,N_3163);
nor U4240 (N_4240,N_3670,N_3884);
nor U4241 (N_4241,N_3278,N_3551);
nand U4242 (N_4242,N_3897,N_3914);
nor U4243 (N_4243,N_3666,N_3168);
and U4244 (N_4244,N_3370,N_3594);
and U4245 (N_4245,N_3831,N_3853);
nand U4246 (N_4246,N_3442,N_3359);
and U4247 (N_4247,N_3995,N_3529);
and U4248 (N_4248,N_3491,N_3979);
nand U4249 (N_4249,N_3810,N_3930);
nor U4250 (N_4250,N_3267,N_3996);
nor U4251 (N_4251,N_3506,N_3749);
nand U4252 (N_4252,N_3298,N_3287);
xor U4253 (N_4253,N_3687,N_3518);
nand U4254 (N_4254,N_3521,N_3312);
and U4255 (N_4255,N_3859,N_3982);
and U4256 (N_4256,N_3395,N_3177);
or U4257 (N_4257,N_3936,N_3590);
nor U4258 (N_4258,N_3214,N_3269);
nor U4259 (N_4259,N_3143,N_3841);
nand U4260 (N_4260,N_3719,N_3771);
nand U4261 (N_4261,N_3967,N_3686);
nor U4262 (N_4262,N_3273,N_3925);
xor U4263 (N_4263,N_3201,N_3586);
xnor U4264 (N_4264,N_3241,N_3715);
nor U4265 (N_4265,N_3540,N_3258);
xor U4266 (N_4266,N_3880,N_3068);
nand U4267 (N_4267,N_3855,N_3587);
nand U4268 (N_4268,N_3774,N_3238);
nor U4269 (N_4269,N_3840,N_3125);
and U4270 (N_4270,N_3502,N_3908);
and U4271 (N_4271,N_3555,N_3917);
nand U4272 (N_4272,N_3512,N_3584);
nor U4273 (N_4273,N_3545,N_3165);
and U4274 (N_4274,N_3160,N_3076);
nor U4275 (N_4275,N_3808,N_3088);
and U4276 (N_4276,N_3579,N_3694);
xor U4277 (N_4277,N_3567,N_3237);
nor U4278 (N_4278,N_3863,N_3250);
or U4279 (N_4279,N_3746,N_3046);
nor U4280 (N_4280,N_3393,N_3325);
and U4281 (N_4281,N_3802,N_3056);
or U4282 (N_4282,N_3347,N_3671);
nor U4283 (N_4283,N_3118,N_3901);
xnor U4284 (N_4284,N_3288,N_3436);
and U4285 (N_4285,N_3896,N_3494);
and U4286 (N_4286,N_3892,N_3667);
or U4287 (N_4287,N_3630,N_3903);
or U4288 (N_4288,N_3732,N_3004);
nor U4289 (N_4289,N_3992,N_3817);
nand U4290 (N_4290,N_3405,N_3517);
and U4291 (N_4291,N_3175,N_3993);
or U4292 (N_4292,N_3136,N_3372);
xor U4293 (N_4293,N_3523,N_3423);
nand U4294 (N_4294,N_3246,N_3765);
nor U4295 (N_4295,N_3256,N_3295);
or U4296 (N_4296,N_3612,N_3300);
or U4297 (N_4297,N_3724,N_3240);
nand U4298 (N_4298,N_3986,N_3028);
nand U4299 (N_4299,N_3735,N_3530);
and U4300 (N_4300,N_3570,N_3197);
nor U4301 (N_4301,N_3110,N_3444);
nand U4302 (N_4302,N_3572,N_3215);
nand U4303 (N_4303,N_3282,N_3585);
or U4304 (N_4304,N_3819,N_3401);
and U4305 (N_4305,N_3080,N_3860);
or U4306 (N_4306,N_3824,N_3315);
xor U4307 (N_4307,N_3284,N_3445);
and U4308 (N_4308,N_3582,N_3864);
xnor U4309 (N_4309,N_3645,N_3171);
or U4310 (N_4310,N_3970,N_3637);
nor U4311 (N_4311,N_3509,N_3311);
nand U4312 (N_4312,N_3141,N_3784);
xnor U4313 (N_4313,N_3828,N_3994);
xnor U4314 (N_4314,N_3879,N_3974);
or U4315 (N_4315,N_3758,N_3382);
nand U4316 (N_4316,N_3490,N_3722);
and U4317 (N_4317,N_3450,N_3367);
xor U4318 (N_4318,N_3087,N_3021);
nand U4319 (N_4319,N_3335,N_3633);
or U4320 (N_4320,N_3761,N_3362);
xor U4321 (N_4321,N_3727,N_3301);
xnor U4322 (N_4322,N_3913,N_3886);
xnor U4323 (N_4323,N_3920,N_3406);
and U4324 (N_4324,N_3790,N_3797);
xor U4325 (N_4325,N_3608,N_3638);
and U4326 (N_4326,N_3559,N_3403);
xnor U4327 (N_4327,N_3067,N_3228);
nor U4328 (N_4328,N_3869,N_3815);
or U4329 (N_4329,N_3692,N_3730);
or U4330 (N_4330,N_3887,N_3827);
and U4331 (N_4331,N_3685,N_3127);
or U4332 (N_4332,N_3924,N_3621);
nor U4333 (N_4333,N_3838,N_3741);
xor U4334 (N_4334,N_3398,N_3043);
and U4335 (N_4335,N_3310,N_3659);
nor U4336 (N_4336,N_3386,N_3700);
and U4337 (N_4337,N_3969,N_3738);
nor U4338 (N_4338,N_3911,N_3365);
xnor U4339 (N_4339,N_3807,N_3275);
or U4340 (N_4340,N_3097,N_3333);
and U4341 (N_4341,N_3470,N_3451);
nand U4342 (N_4342,N_3550,N_3255);
nand U4343 (N_4343,N_3485,N_3234);
and U4344 (N_4344,N_3060,N_3181);
or U4345 (N_4345,N_3983,N_3935);
nand U4346 (N_4346,N_3955,N_3604);
xor U4347 (N_4347,N_3430,N_3279);
or U4348 (N_4348,N_3369,N_3737);
nand U4349 (N_4349,N_3180,N_3984);
or U4350 (N_4350,N_3299,N_3617);
or U4351 (N_4351,N_3126,N_3862);
nor U4352 (N_4352,N_3244,N_3281);
xor U4353 (N_4353,N_3985,N_3927);
or U4354 (N_4354,N_3829,N_3089);
nor U4355 (N_4355,N_3014,N_3705);
nor U4356 (N_4356,N_3041,N_3113);
and U4357 (N_4357,N_3419,N_3654);
or U4358 (N_4358,N_3656,N_3643);
xor U4359 (N_4359,N_3602,N_3407);
or U4360 (N_4360,N_3837,N_3090);
or U4361 (N_4361,N_3032,N_3242);
xor U4362 (N_4362,N_3938,N_3921);
nor U4363 (N_4363,N_3042,N_3019);
nor U4364 (N_4364,N_3107,N_3239);
nand U4365 (N_4365,N_3904,N_3159);
nor U4366 (N_4366,N_3739,N_3040);
or U4367 (N_4367,N_3548,N_3231);
and U4368 (N_4368,N_3134,N_3411);
or U4369 (N_4369,N_3721,N_3878);
and U4370 (N_4370,N_3326,N_3373);
nor U4371 (N_4371,N_3387,N_3998);
nand U4372 (N_4372,N_3681,N_3319);
nand U4373 (N_4373,N_3399,N_3262);
or U4374 (N_4374,N_3842,N_3294);
or U4375 (N_4375,N_3893,N_3498);
xor U4376 (N_4376,N_3193,N_3410);
nor U4377 (N_4377,N_3662,N_3755);
nand U4378 (N_4378,N_3519,N_3476);
and U4379 (N_4379,N_3812,N_3013);
or U4380 (N_4380,N_3711,N_3486);
or U4381 (N_4381,N_3573,N_3614);
and U4382 (N_4382,N_3888,N_3513);
xnor U4383 (N_4383,N_3663,N_3375);
or U4384 (N_4384,N_3640,N_3657);
and U4385 (N_4385,N_3341,N_3277);
or U4386 (N_4386,N_3361,N_3116);
xor U4387 (N_4387,N_3588,N_3873);
or U4388 (N_4388,N_3167,N_3471);
xor U4389 (N_4389,N_3851,N_3022);
and U4390 (N_4390,N_3791,N_3933);
and U4391 (N_4391,N_3413,N_3562);
and U4392 (N_4392,N_3458,N_3589);
nand U4393 (N_4393,N_3781,N_3980);
xnor U4394 (N_4394,N_3767,N_3183);
or U4395 (N_4395,N_3409,N_3825);
nor U4396 (N_4396,N_3546,N_3806);
nand U4397 (N_4397,N_3106,N_3650);
and U4398 (N_4398,N_3428,N_3477);
or U4399 (N_4399,N_3404,N_3757);
and U4400 (N_4400,N_3217,N_3388);
nand U4401 (N_4401,N_3426,N_3634);
or U4402 (N_4402,N_3130,N_3963);
and U4403 (N_4403,N_3818,N_3212);
and U4404 (N_4404,N_3460,N_3396);
nor U4405 (N_4405,N_3769,N_3596);
nor U4406 (N_4406,N_3185,N_3581);
nor U4407 (N_4407,N_3763,N_3811);
or U4408 (N_4408,N_3148,N_3226);
and U4409 (N_4409,N_3620,N_3624);
nor U4410 (N_4410,N_3902,N_3030);
and U4411 (N_4411,N_3743,N_3461);
and U4412 (N_4412,N_3355,N_3641);
xnor U4413 (N_4413,N_3352,N_3547);
nand U4414 (N_4414,N_3704,N_3597);
and U4415 (N_4415,N_3272,N_3906);
or U4416 (N_4416,N_3149,N_3932);
nor U4417 (N_4417,N_3625,N_3198);
xor U4418 (N_4418,N_3764,N_3499);
nor U4419 (N_4419,N_3285,N_3108);
nand U4420 (N_4420,N_3978,N_3975);
and U4421 (N_4421,N_3532,N_3003);
nand U4422 (N_4422,N_3472,N_3096);
xor U4423 (N_4423,N_3948,N_3059);
nor U4424 (N_4424,N_3675,N_3497);
and U4425 (N_4425,N_3100,N_3846);
nand U4426 (N_4426,N_3233,N_3034);
or U4427 (N_4427,N_3564,N_3008);
and U4428 (N_4428,N_3883,N_3176);
xor U4429 (N_4429,N_3563,N_3861);
nor U4430 (N_4430,N_3712,N_3402);
nor U4431 (N_4431,N_3794,N_3990);
nand U4432 (N_4432,N_3219,N_3111);
or U4433 (N_4433,N_3910,N_3363);
nor U4434 (N_4434,N_3642,N_3568);
nand U4435 (N_4435,N_3204,N_3169);
nor U4436 (N_4436,N_3805,N_3527);
xor U4437 (N_4437,N_3351,N_3252);
nor U4438 (N_4438,N_3063,N_3554);
and U4439 (N_4439,N_3002,N_3020);
xnor U4440 (N_4440,N_3344,N_3937);
xnor U4441 (N_4441,N_3698,N_3379);
or U4442 (N_4442,N_3009,N_3408);
and U4443 (N_4443,N_3158,N_3725);
nor U4444 (N_4444,N_3480,N_3745);
xnor U4445 (N_4445,N_3576,N_3987);
and U4446 (N_4446,N_3615,N_3391);
nor U4447 (N_4447,N_3082,N_3314);
xor U4448 (N_4448,N_3504,N_3557);
nor U4449 (N_4449,N_3316,N_3786);
xor U4450 (N_4450,N_3437,N_3928);
xnor U4451 (N_4451,N_3307,N_3412);
xnor U4452 (N_4452,N_3434,N_3977);
nor U4453 (N_4453,N_3782,N_3753);
or U4454 (N_4454,N_3422,N_3447);
xor U4455 (N_4455,N_3505,N_3777);
nor U4456 (N_4456,N_3854,N_3961);
nand U4457 (N_4457,N_3636,N_3894);
and U4458 (N_4458,N_3001,N_3203);
or U4459 (N_4459,N_3865,N_3154);
or U4460 (N_4460,N_3991,N_3427);
or U4461 (N_4461,N_3876,N_3330);
nor U4462 (N_4462,N_3286,N_3025);
or U4463 (N_4463,N_3385,N_3206);
and U4464 (N_4464,N_3680,N_3334);
or U4465 (N_4465,N_3514,N_3338);
xnor U4466 (N_4466,N_3155,N_3655);
nand U4467 (N_4467,N_3780,N_3569);
or U4468 (N_4468,N_3161,N_3037);
nand U4469 (N_4469,N_3031,N_3071);
xnor U4470 (N_4470,N_3075,N_3179);
nor U4471 (N_4471,N_3000,N_3598);
and U4472 (N_4472,N_3354,N_3202);
and U4473 (N_4473,N_3661,N_3696);
nand U4474 (N_4474,N_3858,N_3500);
nor U4475 (N_4475,N_3452,N_3195);
xnor U4476 (N_4476,N_3701,N_3525);
xor U4477 (N_4477,N_3038,N_3015);
nor U4478 (N_4478,N_3462,N_3610);
and U4479 (N_4479,N_3007,N_3062);
xor U4480 (N_4480,N_3956,N_3440);
and U4481 (N_4481,N_3742,N_3380);
nor U4482 (N_4482,N_3194,N_3368);
and U4483 (N_4483,N_3439,N_3109);
or U4484 (N_4484,N_3122,N_3152);
xnor U4485 (N_4485,N_3229,N_3456);
or U4486 (N_4486,N_3397,N_3714);
xnor U4487 (N_4487,N_3174,N_3770);
xnor U4488 (N_4488,N_3200,N_3188);
and U4489 (N_4489,N_3717,N_3142);
or U4490 (N_4490,N_3950,N_3482);
nor U4491 (N_4491,N_3809,N_3178);
nor U4492 (N_4492,N_3072,N_3976);
nor U4493 (N_4493,N_3939,N_3804);
nand U4494 (N_4494,N_3522,N_3626);
nand U4495 (N_4495,N_3356,N_3789);
xor U4496 (N_4496,N_3389,N_3213);
and U4497 (N_4497,N_3102,N_3792);
nor U4498 (N_4498,N_3678,N_3571);
xnor U4499 (N_4499,N_3536,N_3756);
and U4500 (N_4500,N_3826,N_3842);
nor U4501 (N_4501,N_3651,N_3001);
nand U4502 (N_4502,N_3040,N_3573);
or U4503 (N_4503,N_3578,N_3561);
or U4504 (N_4504,N_3812,N_3179);
nor U4505 (N_4505,N_3224,N_3243);
nand U4506 (N_4506,N_3237,N_3276);
or U4507 (N_4507,N_3108,N_3101);
nand U4508 (N_4508,N_3966,N_3816);
xor U4509 (N_4509,N_3754,N_3507);
or U4510 (N_4510,N_3503,N_3797);
or U4511 (N_4511,N_3483,N_3381);
or U4512 (N_4512,N_3901,N_3760);
or U4513 (N_4513,N_3857,N_3080);
xnor U4514 (N_4514,N_3419,N_3327);
and U4515 (N_4515,N_3587,N_3954);
and U4516 (N_4516,N_3522,N_3863);
or U4517 (N_4517,N_3904,N_3636);
xor U4518 (N_4518,N_3800,N_3810);
nor U4519 (N_4519,N_3181,N_3847);
xor U4520 (N_4520,N_3649,N_3889);
and U4521 (N_4521,N_3843,N_3092);
and U4522 (N_4522,N_3519,N_3565);
xnor U4523 (N_4523,N_3013,N_3731);
xor U4524 (N_4524,N_3917,N_3031);
xor U4525 (N_4525,N_3082,N_3001);
xnor U4526 (N_4526,N_3134,N_3645);
or U4527 (N_4527,N_3806,N_3339);
or U4528 (N_4528,N_3535,N_3884);
and U4529 (N_4529,N_3146,N_3224);
nor U4530 (N_4530,N_3789,N_3501);
xnor U4531 (N_4531,N_3098,N_3925);
or U4532 (N_4532,N_3792,N_3279);
nand U4533 (N_4533,N_3129,N_3229);
and U4534 (N_4534,N_3283,N_3298);
nor U4535 (N_4535,N_3917,N_3411);
or U4536 (N_4536,N_3266,N_3319);
and U4537 (N_4537,N_3987,N_3691);
and U4538 (N_4538,N_3213,N_3317);
nor U4539 (N_4539,N_3777,N_3206);
xor U4540 (N_4540,N_3583,N_3383);
and U4541 (N_4541,N_3295,N_3856);
xor U4542 (N_4542,N_3497,N_3600);
xor U4543 (N_4543,N_3834,N_3793);
nand U4544 (N_4544,N_3592,N_3423);
nand U4545 (N_4545,N_3877,N_3287);
nand U4546 (N_4546,N_3400,N_3211);
xnor U4547 (N_4547,N_3026,N_3368);
or U4548 (N_4548,N_3572,N_3040);
xor U4549 (N_4549,N_3634,N_3892);
and U4550 (N_4550,N_3544,N_3229);
xor U4551 (N_4551,N_3533,N_3146);
nor U4552 (N_4552,N_3468,N_3222);
or U4553 (N_4553,N_3786,N_3957);
nor U4554 (N_4554,N_3434,N_3517);
or U4555 (N_4555,N_3144,N_3798);
or U4556 (N_4556,N_3534,N_3161);
and U4557 (N_4557,N_3149,N_3092);
nor U4558 (N_4558,N_3420,N_3786);
or U4559 (N_4559,N_3819,N_3707);
xor U4560 (N_4560,N_3094,N_3902);
and U4561 (N_4561,N_3487,N_3690);
or U4562 (N_4562,N_3599,N_3420);
xor U4563 (N_4563,N_3408,N_3825);
xor U4564 (N_4564,N_3857,N_3968);
nor U4565 (N_4565,N_3063,N_3033);
nor U4566 (N_4566,N_3131,N_3531);
nand U4567 (N_4567,N_3025,N_3398);
nand U4568 (N_4568,N_3413,N_3984);
nor U4569 (N_4569,N_3932,N_3170);
nand U4570 (N_4570,N_3703,N_3551);
and U4571 (N_4571,N_3741,N_3777);
xor U4572 (N_4572,N_3526,N_3846);
and U4573 (N_4573,N_3708,N_3377);
or U4574 (N_4574,N_3984,N_3017);
or U4575 (N_4575,N_3414,N_3987);
or U4576 (N_4576,N_3823,N_3918);
or U4577 (N_4577,N_3155,N_3829);
nor U4578 (N_4578,N_3436,N_3548);
nor U4579 (N_4579,N_3160,N_3220);
and U4580 (N_4580,N_3961,N_3035);
and U4581 (N_4581,N_3886,N_3385);
and U4582 (N_4582,N_3278,N_3810);
nand U4583 (N_4583,N_3494,N_3053);
nand U4584 (N_4584,N_3098,N_3663);
and U4585 (N_4585,N_3789,N_3139);
nand U4586 (N_4586,N_3007,N_3257);
xor U4587 (N_4587,N_3929,N_3586);
xor U4588 (N_4588,N_3983,N_3944);
and U4589 (N_4589,N_3397,N_3810);
or U4590 (N_4590,N_3920,N_3264);
xnor U4591 (N_4591,N_3504,N_3934);
or U4592 (N_4592,N_3426,N_3063);
nor U4593 (N_4593,N_3587,N_3794);
or U4594 (N_4594,N_3414,N_3181);
nand U4595 (N_4595,N_3376,N_3787);
or U4596 (N_4596,N_3925,N_3780);
nor U4597 (N_4597,N_3951,N_3054);
nand U4598 (N_4598,N_3610,N_3807);
or U4599 (N_4599,N_3135,N_3534);
or U4600 (N_4600,N_3090,N_3898);
nor U4601 (N_4601,N_3926,N_3932);
nand U4602 (N_4602,N_3450,N_3785);
nor U4603 (N_4603,N_3414,N_3643);
nand U4604 (N_4604,N_3794,N_3407);
xnor U4605 (N_4605,N_3279,N_3886);
nor U4606 (N_4606,N_3368,N_3631);
nand U4607 (N_4607,N_3100,N_3102);
nand U4608 (N_4608,N_3287,N_3288);
nor U4609 (N_4609,N_3306,N_3168);
and U4610 (N_4610,N_3790,N_3553);
or U4611 (N_4611,N_3406,N_3576);
nand U4612 (N_4612,N_3841,N_3175);
nor U4613 (N_4613,N_3728,N_3612);
or U4614 (N_4614,N_3374,N_3206);
xor U4615 (N_4615,N_3413,N_3502);
xor U4616 (N_4616,N_3019,N_3169);
nand U4617 (N_4617,N_3124,N_3123);
xnor U4618 (N_4618,N_3013,N_3092);
nor U4619 (N_4619,N_3217,N_3531);
and U4620 (N_4620,N_3290,N_3156);
or U4621 (N_4621,N_3086,N_3570);
and U4622 (N_4622,N_3172,N_3263);
xor U4623 (N_4623,N_3897,N_3372);
and U4624 (N_4624,N_3513,N_3250);
or U4625 (N_4625,N_3295,N_3101);
nor U4626 (N_4626,N_3349,N_3018);
or U4627 (N_4627,N_3364,N_3840);
xor U4628 (N_4628,N_3240,N_3543);
and U4629 (N_4629,N_3670,N_3915);
nor U4630 (N_4630,N_3995,N_3426);
nand U4631 (N_4631,N_3266,N_3593);
xnor U4632 (N_4632,N_3726,N_3655);
xor U4633 (N_4633,N_3592,N_3574);
xor U4634 (N_4634,N_3551,N_3268);
nand U4635 (N_4635,N_3156,N_3904);
xnor U4636 (N_4636,N_3061,N_3148);
or U4637 (N_4637,N_3658,N_3898);
nand U4638 (N_4638,N_3886,N_3082);
and U4639 (N_4639,N_3589,N_3117);
nor U4640 (N_4640,N_3432,N_3755);
and U4641 (N_4641,N_3042,N_3470);
or U4642 (N_4642,N_3413,N_3937);
nand U4643 (N_4643,N_3220,N_3623);
nor U4644 (N_4644,N_3098,N_3445);
xor U4645 (N_4645,N_3031,N_3231);
xor U4646 (N_4646,N_3687,N_3828);
and U4647 (N_4647,N_3845,N_3818);
nor U4648 (N_4648,N_3457,N_3298);
and U4649 (N_4649,N_3850,N_3982);
and U4650 (N_4650,N_3759,N_3080);
or U4651 (N_4651,N_3151,N_3796);
nand U4652 (N_4652,N_3385,N_3739);
nand U4653 (N_4653,N_3559,N_3989);
nand U4654 (N_4654,N_3405,N_3095);
nand U4655 (N_4655,N_3427,N_3685);
xnor U4656 (N_4656,N_3965,N_3008);
nand U4657 (N_4657,N_3997,N_3231);
xnor U4658 (N_4658,N_3816,N_3917);
nand U4659 (N_4659,N_3634,N_3850);
nand U4660 (N_4660,N_3657,N_3919);
nand U4661 (N_4661,N_3116,N_3560);
nor U4662 (N_4662,N_3919,N_3958);
nand U4663 (N_4663,N_3057,N_3810);
and U4664 (N_4664,N_3689,N_3741);
nor U4665 (N_4665,N_3109,N_3539);
or U4666 (N_4666,N_3047,N_3558);
nor U4667 (N_4667,N_3523,N_3670);
or U4668 (N_4668,N_3575,N_3249);
and U4669 (N_4669,N_3630,N_3500);
nor U4670 (N_4670,N_3551,N_3849);
nand U4671 (N_4671,N_3260,N_3489);
and U4672 (N_4672,N_3952,N_3317);
or U4673 (N_4673,N_3746,N_3698);
and U4674 (N_4674,N_3638,N_3363);
and U4675 (N_4675,N_3734,N_3362);
xnor U4676 (N_4676,N_3343,N_3556);
xnor U4677 (N_4677,N_3933,N_3328);
nand U4678 (N_4678,N_3065,N_3798);
or U4679 (N_4679,N_3774,N_3624);
nand U4680 (N_4680,N_3835,N_3285);
nor U4681 (N_4681,N_3529,N_3743);
xnor U4682 (N_4682,N_3842,N_3262);
nand U4683 (N_4683,N_3570,N_3758);
and U4684 (N_4684,N_3732,N_3813);
xnor U4685 (N_4685,N_3668,N_3162);
nand U4686 (N_4686,N_3037,N_3086);
nor U4687 (N_4687,N_3654,N_3849);
nor U4688 (N_4688,N_3155,N_3630);
or U4689 (N_4689,N_3221,N_3824);
nor U4690 (N_4690,N_3503,N_3717);
nand U4691 (N_4691,N_3938,N_3584);
nor U4692 (N_4692,N_3246,N_3412);
or U4693 (N_4693,N_3956,N_3599);
and U4694 (N_4694,N_3331,N_3818);
and U4695 (N_4695,N_3076,N_3658);
nor U4696 (N_4696,N_3620,N_3912);
nor U4697 (N_4697,N_3336,N_3095);
nor U4698 (N_4698,N_3306,N_3531);
nand U4699 (N_4699,N_3964,N_3825);
and U4700 (N_4700,N_3141,N_3410);
or U4701 (N_4701,N_3002,N_3876);
nor U4702 (N_4702,N_3289,N_3699);
xnor U4703 (N_4703,N_3537,N_3125);
nor U4704 (N_4704,N_3064,N_3905);
nor U4705 (N_4705,N_3538,N_3397);
or U4706 (N_4706,N_3120,N_3871);
and U4707 (N_4707,N_3706,N_3978);
nand U4708 (N_4708,N_3468,N_3252);
and U4709 (N_4709,N_3554,N_3361);
xnor U4710 (N_4710,N_3061,N_3191);
nand U4711 (N_4711,N_3545,N_3840);
nand U4712 (N_4712,N_3254,N_3543);
nand U4713 (N_4713,N_3997,N_3745);
nor U4714 (N_4714,N_3931,N_3818);
nand U4715 (N_4715,N_3474,N_3636);
nand U4716 (N_4716,N_3623,N_3625);
or U4717 (N_4717,N_3512,N_3579);
or U4718 (N_4718,N_3307,N_3367);
xnor U4719 (N_4719,N_3098,N_3686);
and U4720 (N_4720,N_3114,N_3273);
nand U4721 (N_4721,N_3967,N_3166);
or U4722 (N_4722,N_3507,N_3652);
xnor U4723 (N_4723,N_3181,N_3519);
nor U4724 (N_4724,N_3804,N_3963);
xor U4725 (N_4725,N_3488,N_3210);
or U4726 (N_4726,N_3310,N_3969);
nor U4727 (N_4727,N_3569,N_3873);
xor U4728 (N_4728,N_3926,N_3471);
or U4729 (N_4729,N_3820,N_3016);
and U4730 (N_4730,N_3044,N_3555);
nor U4731 (N_4731,N_3262,N_3635);
nand U4732 (N_4732,N_3718,N_3869);
nand U4733 (N_4733,N_3576,N_3580);
xnor U4734 (N_4734,N_3628,N_3079);
or U4735 (N_4735,N_3429,N_3079);
or U4736 (N_4736,N_3082,N_3587);
and U4737 (N_4737,N_3099,N_3611);
xor U4738 (N_4738,N_3446,N_3848);
nor U4739 (N_4739,N_3714,N_3108);
and U4740 (N_4740,N_3868,N_3092);
nand U4741 (N_4741,N_3297,N_3407);
and U4742 (N_4742,N_3644,N_3396);
nor U4743 (N_4743,N_3487,N_3421);
and U4744 (N_4744,N_3245,N_3973);
and U4745 (N_4745,N_3467,N_3337);
nand U4746 (N_4746,N_3167,N_3781);
or U4747 (N_4747,N_3706,N_3661);
and U4748 (N_4748,N_3923,N_3833);
and U4749 (N_4749,N_3318,N_3857);
nor U4750 (N_4750,N_3426,N_3074);
xnor U4751 (N_4751,N_3690,N_3410);
nor U4752 (N_4752,N_3788,N_3706);
nor U4753 (N_4753,N_3509,N_3196);
or U4754 (N_4754,N_3463,N_3142);
nand U4755 (N_4755,N_3107,N_3961);
or U4756 (N_4756,N_3168,N_3202);
or U4757 (N_4757,N_3461,N_3509);
nand U4758 (N_4758,N_3447,N_3353);
nor U4759 (N_4759,N_3815,N_3843);
nand U4760 (N_4760,N_3649,N_3642);
nor U4761 (N_4761,N_3626,N_3974);
and U4762 (N_4762,N_3683,N_3982);
xor U4763 (N_4763,N_3434,N_3198);
nand U4764 (N_4764,N_3757,N_3562);
xnor U4765 (N_4765,N_3088,N_3426);
or U4766 (N_4766,N_3651,N_3905);
nor U4767 (N_4767,N_3938,N_3465);
nor U4768 (N_4768,N_3717,N_3884);
or U4769 (N_4769,N_3696,N_3002);
nand U4770 (N_4770,N_3540,N_3279);
nor U4771 (N_4771,N_3621,N_3647);
or U4772 (N_4772,N_3934,N_3599);
and U4773 (N_4773,N_3280,N_3833);
xor U4774 (N_4774,N_3123,N_3458);
nand U4775 (N_4775,N_3003,N_3036);
or U4776 (N_4776,N_3767,N_3049);
xnor U4777 (N_4777,N_3715,N_3821);
nor U4778 (N_4778,N_3592,N_3310);
xnor U4779 (N_4779,N_3746,N_3772);
and U4780 (N_4780,N_3878,N_3646);
xnor U4781 (N_4781,N_3295,N_3953);
and U4782 (N_4782,N_3640,N_3330);
and U4783 (N_4783,N_3207,N_3441);
nand U4784 (N_4784,N_3436,N_3157);
nand U4785 (N_4785,N_3033,N_3124);
xor U4786 (N_4786,N_3077,N_3216);
xor U4787 (N_4787,N_3282,N_3846);
or U4788 (N_4788,N_3119,N_3312);
xnor U4789 (N_4789,N_3479,N_3693);
nand U4790 (N_4790,N_3867,N_3998);
nor U4791 (N_4791,N_3540,N_3119);
and U4792 (N_4792,N_3078,N_3612);
or U4793 (N_4793,N_3245,N_3949);
nand U4794 (N_4794,N_3941,N_3606);
and U4795 (N_4795,N_3891,N_3261);
nor U4796 (N_4796,N_3825,N_3056);
nor U4797 (N_4797,N_3980,N_3404);
nand U4798 (N_4798,N_3511,N_3148);
or U4799 (N_4799,N_3388,N_3577);
nor U4800 (N_4800,N_3916,N_3411);
and U4801 (N_4801,N_3655,N_3764);
or U4802 (N_4802,N_3352,N_3541);
and U4803 (N_4803,N_3339,N_3321);
or U4804 (N_4804,N_3249,N_3682);
nand U4805 (N_4805,N_3684,N_3028);
nor U4806 (N_4806,N_3832,N_3412);
and U4807 (N_4807,N_3037,N_3586);
and U4808 (N_4808,N_3769,N_3623);
or U4809 (N_4809,N_3605,N_3553);
nand U4810 (N_4810,N_3072,N_3872);
nor U4811 (N_4811,N_3391,N_3366);
and U4812 (N_4812,N_3855,N_3415);
nor U4813 (N_4813,N_3879,N_3251);
nor U4814 (N_4814,N_3313,N_3675);
xor U4815 (N_4815,N_3075,N_3122);
nor U4816 (N_4816,N_3068,N_3004);
nor U4817 (N_4817,N_3938,N_3708);
xnor U4818 (N_4818,N_3794,N_3709);
and U4819 (N_4819,N_3863,N_3139);
or U4820 (N_4820,N_3741,N_3796);
nor U4821 (N_4821,N_3239,N_3761);
or U4822 (N_4822,N_3610,N_3752);
and U4823 (N_4823,N_3748,N_3775);
nor U4824 (N_4824,N_3397,N_3371);
and U4825 (N_4825,N_3836,N_3791);
or U4826 (N_4826,N_3169,N_3147);
and U4827 (N_4827,N_3776,N_3219);
xor U4828 (N_4828,N_3000,N_3281);
xnor U4829 (N_4829,N_3372,N_3260);
and U4830 (N_4830,N_3408,N_3154);
nand U4831 (N_4831,N_3562,N_3751);
xnor U4832 (N_4832,N_3003,N_3844);
nor U4833 (N_4833,N_3064,N_3760);
nor U4834 (N_4834,N_3303,N_3158);
nand U4835 (N_4835,N_3334,N_3056);
and U4836 (N_4836,N_3071,N_3127);
and U4837 (N_4837,N_3893,N_3532);
or U4838 (N_4838,N_3976,N_3971);
or U4839 (N_4839,N_3678,N_3426);
xor U4840 (N_4840,N_3026,N_3877);
or U4841 (N_4841,N_3330,N_3788);
nor U4842 (N_4842,N_3680,N_3232);
or U4843 (N_4843,N_3048,N_3530);
nand U4844 (N_4844,N_3068,N_3300);
and U4845 (N_4845,N_3768,N_3542);
and U4846 (N_4846,N_3962,N_3055);
or U4847 (N_4847,N_3819,N_3920);
and U4848 (N_4848,N_3899,N_3950);
or U4849 (N_4849,N_3713,N_3015);
nor U4850 (N_4850,N_3196,N_3807);
nand U4851 (N_4851,N_3875,N_3545);
nor U4852 (N_4852,N_3517,N_3745);
xor U4853 (N_4853,N_3441,N_3378);
nor U4854 (N_4854,N_3974,N_3256);
or U4855 (N_4855,N_3115,N_3532);
nand U4856 (N_4856,N_3576,N_3379);
nor U4857 (N_4857,N_3025,N_3534);
xnor U4858 (N_4858,N_3300,N_3767);
or U4859 (N_4859,N_3476,N_3508);
and U4860 (N_4860,N_3389,N_3185);
and U4861 (N_4861,N_3716,N_3266);
xnor U4862 (N_4862,N_3180,N_3174);
or U4863 (N_4863,N_3038,N_3431);
nand U4864 (N_4864,N_3024,N_3319);
and U4865 (N_4865,N_3600,N_3403);
nor U4866 (N_4866,N_3679,N_3845);
and U4867 (N_4867,N_3845,N_3821);
nand U4868 (N_4868,N_3615,N_3837);
nand U4869 (N_4869,N_3501,N_3004);
nand U4870 (N_4870,N_3732,N_3113);
or U4871 (N_4871,N_3374,N_3849);
nand U4872 (N_4872,N_3718,N_3806);
or U4873 (N_4873,N_3534,N_3093);
xor U4874 (N_4874,N_3346,N_3023);
xor U4875 (N_4875,N_3352,N_3687);
xnor U4876 (N_4876,N_3243,N_3323);
and U4877 (N_4877,N_3973,N_3856);
or U4878 (N_4878,N_3790,N_3455);
or U4879 (N_4879,N_3425,N_3643);
or U4880 (N_4880,N_3273,N_3965);
nand U4881 (N_4881,N_3061,N_3883);
xnor U4882 (N_4882,N_3500,N_3022);
or U4883 (N_4883,N_3277,N_3848);
nor U4884 (N_4884,N_3583,N_3974);
xnor U4885 (N_4885,N_3243,N_3903);
nor U4886 (N_4886,N_3964,N_3165);
xnor U4887 (N_4887,N_3771,N_3859);
nand U4888 (N_4888,N_3417,N_3087);
nor U4889 (N_4889,N_3401,N_3706);
and U4890 (N_4890,N_3183,N_3662);
nand U4891 (N_4891,N_3099,N_3642);
xnor U4892 (N_4892,N_3614,N_3966);
nor U4893 (N_4893,N_3356,N_3898);
or U4894 (N_4894,N_3493,N_3983);
or U4895 (N_4895,N_3307,N_3852);
nand U4896 (N_4896,N_3811,N_3800);
or U4897 (N_4897,N_3622,N_3726);
nand U4898 (N_4898,N_3552,N_3498);
xnor U4899 (N_4899,N_3776,N_3971);
nand U4900 (N_4900,N_3777,N_3572);
xnor U4901 (N_4901,N_3268,N_3556);
nor U4902 (N_4902,N_3855,N_3009);
nor U4903 (N_4903,N_3516,N_3375);
xnor U4904 (N_4904,N_3461,N_3702);
or U4905 (N_4905,N_3458,N_3648);
or U4906 (N_4906,N_3029,N_3869);
or U4907 (N_4907,N_3003,N_3576);
or U4908 (N_4908,N_3369,N_3148);
xor U4909 (N_4909,N_3128,N_3983);
or U4910 (N_4910,N_3305,N_3574);
xor U4911 (N_4911,N_3825,N_3368);
or U4912 (N_4912,N_3019,N_3466);
nand U4913 (N_4913,N_3080,N_3828);
xnor U4914 (N_4914,N_3195,N_3123);
xnor U4915 (N_4915,N_3338,N_3718);
xor U4916 (N_4916,N_3734,N_3970);
nor U4917 (N_4917,N_3933,N_3081);
xnor U4918 (N_4918,N_3410,N_3937);
xnor U4919 (N_4919,N_3625,N_3404);
xor U4920 (N_4920,N_3014,N_3152);
xor U4921 (N_4921,N_3809,N_3294);
and U4922 (N_4922,N_3741,N_3103);
nand U4923 (N_4923,N_3778,N_3382);
xnor U4924 (N_4924,N_3092,N_3090);
nand U4925 (N_4925,N_3533,N_3383);
xnor U4926 (N_4926,N_3558,N_3894);
nor U4927 (N_4927,N_3311,N_3914);
or U4928 (N_4928,N_3948,N_3455);
xnor U4929 (N_4929,N_3631,N_3838);
nor U4930 (N_4930,N_3305,N_3429);
and U4931 (N_4931,N_3518,N_3563);
nor U4932 (N_4932,N_3115,N_3746);
and U4933 (N_4933,N_3700,N_3960);
or U4934 (N_4934,N_3149,N_3541);
and U4935 (N_4935,N_3984,N_3566);
nor U4936 (N_4936,N_3876,N_3834);
xor U4937 (N_4937,N_3465,N_3898);
xor U4938 (N_4938,N_3184,N_3642);
xor U4939 (N_4939,N_3957,N_3883);
or U4940 (N_4940,N_3487,N_3234);
xor U4941 (N_4941,N_3965,N_3285);
and U4942 (N_4942,N_3766,N_3559);
xnor U4943 (N_4943,N_3497,N_3933);
xor U4944 (N_4944,N_3003,N_3557);
nor U4945 (N_4945,N_3518,N_3013);
nor U4946 (N_4946,N_3683,N_3781);
or U4947 (N_4947,N_3969,N_3105);
and U4948 (N_4948,N_3628,N_3383);
xnor U4949 (N_4949,N_3272,N_3546);
nor U4950 (N_4950,N_3457,N_3916);
nand U4951 (N_4951,N_3250,N_3965);
xnor U4952 (N_4952,N_3181,N_3259);
and U4953 (N_4953,N_3310,N_3398);
nand U4954 (N_4954,N_3855,N_3124);
or U4955 (N_4955,N_3475,N_3001);
or U4956 (N_4956,N_3202,N_3094);
or U4957 (N_4957,N_3207,N_3909);
nand U4958 (N_4958,N_3427,N_3390);
and U4959 (N_4959,N_3676,N_3113);
nor U4960 (N_4960,N_3976,N_3186);
xnor U4961 (N_4961,N_3566,N_3442);
or U4962 (N_4962,N_3523,N_3204);
xnor U4963 (N_4963,N_3242,N_3165);
xor U4964 (N_4964,N_3448,N_3915);
nand U4965 (N_4965,N_3578,N_3340);
xor U4966 (N_4966,N_3671,N_3819);
nor U4967 (N_4967,N_3573,N_3413);
or U4968 (N_4968,N_3111,N_3894);
nand U4969 (N_4969,N_3314,N_3534);
xor U4970 (N_4970,N_3030,N_3905);
and U4971 (N_4971,N_3855,N_3333);
nand U4972 (N_4972,N_3158,N_3004);
nand U4973 (N_4973,N_3978,N_3795);
nor U4974 (N_4974,N_3319,N_3988);
and U4975 (N_4975,N_3070,N_3481);
xnor U4976 (N_4976,N_3446,N_3198);
and U4977 (N_4977,N_3970,N_3004);
nand U4978 (N_4978,N_3267,N_3819);
or U4979 (N_4979,N_3511,N_3408);
nor U4980 (N_4980,N_3826,N_3312);
or U4981 (N_4981,N_3705,N_3837);
or U4982 (N_4982,N_3087,N_3953);
nor U4983 (N_4983,N_3046,N_3695);
nand U4984 (N_4984,N_3266,N_3555);
nand U4985 (N_4985,N_3917,N_3022);
and U4986 (N_4986,N_3373,N_3409);
nand U4987 (N_4987,N_3564,N_3973);
nor U4988 (N_4988,N_3406,N_3573);
or U4989 (N_4989,N_3524,N_3046);
nor U4990 (N_4990,N_3290,N_3059);
nand U4991 (N_4991,N_3656,N_3210);
nand U4992 (N_4992,N_3149,N_3538);
and U4993 (N_4993,N_3407,N_3070);
nand U4994 (N_4994,N_3281,N_3736);
and U4995 (N_4995,N_3728,N_3497);
and U4996 (N_4996,N_3222,N_3563);
and U4997 (N_4997,N_3029,N_3941);
and U4998 (N_4998,N_3596,N_3036);
nand U4999 (N_4999,N_3564,N_3116);
and U5000 (N_5000,N_4053,N_4161);
and U5001 (N_5001,N_4360,N_4195);
or U5002 (N_5002,N_4820,N_4952);
nor U5003 (N_5003,N_4887,N_4476);
or U5004 (N_5004,N_4328,N_4213);
xnor U5005 (N_5005,N_4078,N_4098);
xnor U5006 (N_5006,N_4569,N_4060);
nor U5007 (N_5007,N_4624,N_4600);
nand U5008 (N_5008,N_4287,N_4025);
nand U5009 (N_5009,N_4933,N_4826);
nand U5010 (N_5010,N_4253,N_4095);
xnor U5011 (N_5011,N_4712,N_4246);
nand U5012 (N_5012,N_4059,N_4064);
xnor U5013 (N_5013,N_4736,N_4668);
xnor U5014 (N_5014,N_4359,N_4400);
and U5015 (N_5015,N_4941,N_4097);
and U5016 (N_5016,N_4200,N_4319);
nor U5017 (N_5017,N_4088,N_4588);
nand U5018 (N_5018,N_4983,N_4613);
or U5019 (N_5019,N_4960,N_4144);
nor U5020 (N_5020,N_4462,N_4849);
and U5021 (N_5021,N_4667,N_4912);
nor U5022 (N_5022,N_4114,N_4922);
or U5023 (N_5023,N_4857,N_4858);
xor U5024 (N_5024,N_4762,N_4115);
or U5025 (N_5025,N_4555,N_4765);
nor U5026 (N_5026,N_4527,N_4640);
nand U5027 (N_5027,N_4474,N_4615);
and U5028 (N_5028,N_4785,N_4589);
and U5029 (N_5029,N_4152,N_4629);
or U5030 (N_5030,N_4422,N_4111);
and U5031 (N_5031,N_4065,N_4222);
or U5032 (N_5032,N_4998,N_4595);
nand U5033 (N_5033,N_4276,N_4548);
nor U5034 (N_5034,N_4930,N_4583);
or U5035 (N_5035,N_4671,N_4086);
and U5036 (N_5036,N_4986,N_4259);
and U5037 (N_5037,N_4051,N_4610);
nor U5038 (N_5038,N_4010,N_4232);
nand U5039 (N_5039,N_4057,N_4190);
xnor U5040 (N_5040,N_4893,N_4333);
and U5041 (N_5041,N_4974,N_4719);
nor U5042 (N_5042,N_4850,N_4755);
nand U5043 (N_5043,N_4054,N_4718);
xnor U5044 (N_5044,N_4967,N_4137);
nand U5045 (N_5045,N_4158,N_4280);
xnor U5046 (N_5046,N_4894,N_4566);
nand U5047 (N_5047,N_4947,N_4266);
nand U5048 (N_5048,N_4368,N_4380);
nand U5049 (N_5049,N_4677,N_4969);
nand U5050 (N_5050,N_4302,N_4109);
nand U5051 (N_5051,N_4616,N_4028);
and U5052 (N_5052,N_4648,N_4292);
xor U5053 (N_5053,N_4423,N_4140);
xor U5054 (N_5054,N_4305,N_4403);
nor U5055 (N_5055,N_4726,N_4408);
or U5056 (N_5056,N_4920,N_4622);
and U5057 (N_5057,N_4199,N_4759);
xor U5058 (N_5058,N_4714,N_4134);
and U5059 (N_5059,N_4007,N_4508);
and U5060 (N_5060,N_4991,N_4009);
xnor U5061 (N_5061,N_4468,N_4020);
nor U5062 (N_5062,N_4171,N_4662);
or U5063 (N_5063,N_4224,N_4187);
or U5064 (N_5064,N_4744,N_4128);
and U5065 (N_5065,N_4029,N_4657);
nor U5066 (N_5066,N_4901,N_4479);
or U5067 (N_5067,N_4427,N_4963);
nand U5068 (N_5068,N_4632,N_4571);
and U5069 (N_5069,N_4814,N_4483);
and U5070 (N_5070,N_4363,N_4107);
nor U5071 (N_5071,N_4908,N_4611);
nor U5072 (N_5072,N_4383,N_4767);
xnor U5073 (N_5073,N_4532,N_4220);
and U5074 (N_5074,N_4557,N_4037);
xor U5075 (N_5075,N_4943,N_4932);
nand U5076 (N_5076,N_4340,N_4031);
nor U5077 (N_5077,N_4273,N_4663);
or U5078 (N_5078,N_4542,N_4768);
or U5079 (N_5079,N_4560,N_4812);
or U5080 (N_5080,N_4766,N_4900);
xnor U5081 (N_5081,N_4938,N_4829);
nor U5082 (N_5082,N_4233,N_4596);
nor U5083 (N_5083,N_4375,N_4939);
xnor U5084 (N_5084,N_4689,N_4397);
or U5085 (N_5085,N_4732,N_4565);
or U5086 (N_5086,N_4157,N_4590);
or U5087 (N_5087,N_4848,N_4544);
nor U5088 (N_5088,N_4729,N_4416);
xor U5089 (N_5089,N_4819,N_4515);
nand U5090 (N_5090,N_4047,N_4455);
xor U5091 (N_5091,N_4045,N_4904);
and U5092 (N_5092,N_4043,N_4439);
nand U5093 (N_5093,N_4870,N_4646);
and U5094 (N_5094,N_4000,N_4637);
nor U5095 (N_5095,N_4921,N_4772);
nor U5096 (N_5096,N_4521,N_4338);
xnor U5097 (N_5097,N_4722,N_4669);
xor U5098 (N_5098,N_4678,N_4541);
xor U5099 (N_5099,N_4295,N_4499);
xor U5100 (N_5100,N_4618,N_4076);
nor U5101 (N_5101,N_4891,N_4433);
nand U5102 (N_5102,N_4883,N_4916);
nand U5103 (N_5103,N_4309,N_4805);
nor U5104 (N_5104,N_4628,N_4742);
and U5105 (N_5105,N_4582,N_4339);
nor U5106 (N_5106,N_4411,N_4019);
nor U5107 (N_5107,N_4815,N_4807);
nand U5108 (N_5108,N_4334,N_4165);
xnor U5109 (N_5109,N_4531,N_4230);
xnor U5110 (N_5110,N_4208,N_4131);
nor U5111 (N_5111,N_4924,N_4886);
and U5112 (N_5112,N_4080,N_4973);
nand U5113 (N_5113,N_4350,N_4730);
xnor U5114 (N_5114,N_4022,N_4124);
and U5115 (N_5115,N_4591,N_4626);
and U5116 (N_5116,N_4656,N_4189);
and U5117 (N_5117,N_4215,N_4331);
or U5118 (N_5118,N_4166,N_4907);
and U5119 (N_5119,N_4971,N_4804);
nand U5120 (N_5120,N_4257,N_4004);
or U5121 (N_5121,N_4504,N_4281);
nand U5122 (N_5122,N_4523,N_4546);
or U5123 (N_5123,N_4556,N_4659);
and U5124 (N_5124,N_4776,N_4415);
or U5125 (N_5125,N_4688,N_4643);
and U5126 (N_5126,N_4428,N_4371);
nand U5127 (N_5127,N_4855,N_4094);
nor U5128 (N_5128,N_4448,N_4852);
xor U5129 (N_5129,N_4181,N_4306);
xnor U5130 (N_5130,N_4308,N_4242);
and U5131 (N_5131,N_4254,N_4420);
xnor U5132 (N_5132,N_4216,N_4132);
nand U5133 (N_5133,N_4062,N_4313);
nand U5134 (N_5134,N_4261,N_4399);
xor U5135 (N_5135,N_4652,N_4609);
xnor U5136 (N_5136,N_4351,N_4482);
xnor U5137 (N_5137,N_4183,N_4279);
or U5138 (N_5138,N_4364,N_4748);
xnor U5139 (N_5139,N_4035,N_4743);
xor U5140 (N_5140,N_4160,N_4454);
or U5141 (N_5141,N_4405,N_4789);
and U5142 (N_5142,N_4436,N_4223);
or U5143 (N_5143,N_4392,N_4984);
nor U5144 (N_5144,N_4205,N_4593);
xor U5145 (N_5145,N_4617,N_4968);
nand U5146 (N_5146,N_4390,N_4553);
nand U5147 (N_5147,N_4987,N_4075);
nor U5148 (N_5148,N_4877,N_4471);
or U5149 (N_5149,N_4844,N_4191);
or U5150 (N_5150,N_4554,N_4749);
xor U5151 (N_5151,N_4018,N_4002);
and U5152 (N_5152,N_4466,N_4185);
or U5153 (N_5153,N_4015,N_4518);
and U5154 (N_5154,N_4248,N_4388);
nand U5155 (N_5155,N_4690,N_4116);
and U5156 (N_5156,N_4834,N_4642);
nand U5157 (N_5157,N_4150,N_4342);
nand U5158 (N_5158,N_4524,N_4354);
or U5159 (N_5159,N_4070,N_4153);
nor U5160 (N_5160,N_4781,N_4926);
or U5161 (N_5161,N_4243,N_4925);
or U5162 (N_5162,N_4460,N_4937);
nand U5163 (N_5163,N_4437,N_4143);
xnor U5164 (N_5164,N_4089,N_4184);
and U5165 (N_5165,N_4746,N_4434);
xnor U5166 (N_5166,N_4449,N_4394);
nor U5167 (N_5167,N_4135,N_4839);
xnor U5168 (N_5168,N_4809,N_4833);
xnor U5169 (N_5169,N_4911,N_4458);
nor U5170 (N_5170,N_4666,N_4965);
nand U5171 (N_5171,N_4535,N_4847);
xnor U5172 (N_5172,N_4110,N_4816);
nand U5173 (N_5173,N_4811,N_4563);
and U5174 (N_5174,N_4516,N_4083);
or U5175 (N_5175,N_4370,N_4251);
nand U5176 (N_5176,N_4180,N_4284);
or U5177 (N_5177,N_4500,N_4239);
nand U5178 (N_5178,N_4039,N_4585);
nor U5179 (N_5179,N_4813,N_4367);
and U5180 (N_5180,N_4151,N_4021);
nor U5181 (N_5181,N_4564,N_4970);
and U5182 (N_5182,N_4827,N_4576);
and U5183 (N_5183,N_4092,N_4934);
nor U5184 (N_5184,N_4465,N_4487);
xnor U5185 (N_5185,N_4793,N_4587);
nor U5186 (N_5186,N_4303,N_4892);
nor U5187 (N_5187,N_4386,N_4707);
nor U5188 (N_5188,N_4317,N_4994);
or U5189 (N_5189,N_4898,N_4341);
xor U5190 (N_5190,N_4361,N_4602);
xor U5191 (N_5191,N_4505,N_4327);
and U5192 (N_5192,N_4055,N_4771);
xor U5193 (N_5193,N_4325,N_4639);
or U5194 (N_5194,N_4956,N_4369);
and U5195 (N_5195,N_4155,N_4824);
or U5196 (N_5196,N_4096,N_4066);
xnor U5197 (N_5197,N_4985,N_4577);
xor U5198 (N_5198,N_4352,N_4867);
or U5199 (N_5199,N_4896,N_4372);
and U5200 (N_5200,N_4362,N_4227);
and U5201 (N_5201,N_4846,N_4903);
and U5202 (N_5202,N_4606,N_4473);
nand U5203 (N_5203,N_4653,N_4514);
or U5204 (N_5204,N_4869,N_4127);
xor U5205 (N_5205,N_4498,N_4272);
nor U5206 (N_5206,N_4450,N_4806);
nor U5207 (N_5207,N_4296,N_4752);
and U5208 (N_5208,N_4958,N_4463);
and U5209 (N_5209,N_4121,N_4580);
xnor U5210 (N_5210,N_4597,N_4562);
xnor U5211 (N_5211,N_4196,N_4620);
xor U5212 (N_5212,N_4413,N_4927);
nand U5213 (N_5213,N_4972,N_4573);
or U5214 (N_5214,N_4796,N_4263);
and U5215 (N_5215,N_4977,N_4679);
or U5216 (N_5216,N_4130,N_4770);
and U5217 (N_5217,N_4429,N_4214);
nor U5218 (N_5218,N_4779,N_4760);
or U5219 (N_5219,N_4989,N_4838);
nor U5220 (N_5220,N_4120,N_4699);
and U5221 (N_5221,N_4245,N_4778);
nor U5222 (N_5222,N_4490,N_4032);
nand U5223 (N_5223,N_4410,N_4701);
xnor U5224 (N_5224,N_4988,N_4536);
and U5225 (N_5225,N_4440,N_4265);
nor U5226 (N_5226,N_4285,N_4438);
nand U5227 (N_5227,N_4865,N_4337);
nor U5228 (N_5228,N_4997,N_4859);
or U5229 (N_5229,N_4962,N_4212);
xnor U5230 (N_5230,N_4262,N_4145);
and U5231 (N_5231,N_4172,N_4170);
and U5232 (N_5232,N_4188,N_4348);
and U5233 (N_5233,N_4426,N_4698);
xnor U5234 (N_5234,N_4651,N_4286);
and U5235 (N_5235,N_4494,N_4638);
and U5236 (N_5236,N_4421,N_4102);
and U5237 (N_5237,N_4836,N_4747);
xor U5238 (N_5238,N_4530,N_4533);
nor U5239 (N_5239,N_4919,N_4966);
or U5240 (N_5240,N_4040,N_4126);
nand U5241 (N_5241,N_4023,N_4326);
or U5242 (N_5242,N_4978,N_4267);
nand U5243 (N_5243,N_4957,N_4299);
nand U5244 (N_5244,N_4792,N_4680);
nor U5245 (N_5245,N_4357,N_4906);
or U5246 (N_5246,N_4154,N_4148);
nor U5247 (N_5247,N_4407,N_4992);
or U5248 (N_5248,N_4840,N_4751);
xor U5249 (N_5249,N_4905,N_4417);
and U5250 (N_5250,N_4802,N_4349);
nor U5251 (N_5251,N_4928,N_4537);
and U5252 (N_5252,N_4168,N_4122);
or U5253 (N_5253,N_4457,N_4027);
or U5254 (N_5254,N_4353,N_4876);
xnor U5255 (N_5255,N_4141,N_4703);
or U5256 (N_5256,N_4676,N_4129);
nor U5257 (N_5257,N_4228,N_4079);
or U5258 (N_5258,N_4123,N_4721);
nand U5259 (N_5259,N_4159,N_4761);
or U5260 (N_5260,N_4377,N_4226);
or U5261 (N_5261,N_4206,N_4513);
and U5262 (N_5262,N_4330,N_4854);
nand U5263 (N_5263,N_4125,N_4347);
xnor U5264 (N_5264,N_4842,N_4142);
nand U5265 (N_5265,N_4830,N_4885);
xor U5266 (N_5266,N_4660,N_4822);
nand U5267 (N_5267,N_4355,N_4061);
nor U5268 (N_5268,N_4136,N_4627);
xor U5269 (N_5269,N_4645,N_4512);
nand U5270 (N_5270,N_4258,N_4982);
nand U5271 (N_5271,N_4268,N_4745);
or U5272 (N_5272,N_4485,N_4431);
xor U5273 (N_5273,N_4547,N_4255);
nand U5274 (N_5274,N_4697,N_4598);
nor U5275 (N_5275,N_4194,N_4649);
and U5276 (N_5276,N_4739,N_4048);
xor U5277 (N_5277,N_4786,N_4841);
or U5278 (N_5278,N_4241,N_4733);
nor U5279 (N_5279,N_4393,N_4345);
nand U5280 (N_5280,N_4817,N_4495);
and U5281 (N_5281,N_4607,N_4346);
or U5282 (N_5282,N_4260,N_4944);
xnor U5283 (N_5283,N_4418,N_4209);
nor U5284 (N_5284,N_4310,N_4800);
and U5285 (N_5285,N_4492,N_4794);
xor U5286 (N_5286,N_4723,N_4949);
or U5287 (N_5287,N_4594,N_4502);
and U5288 (N_5288,N_4837,N_4534);
nand U5289 (N_5289,N_4307,N_4067);
or U5290 (N_5290,N_4993,N_4808);
xor U5291 (N_5291,N_4551,N_4682);
xor U5292 (N_5292,N_4391,N_4387);
nor U5293 (N_5293,N_4396,N_4236);
and U5294 (N_5294,N_4112,N_4481);
xnor U5295 (N_5295,N_4675,N_4783);
nand U5296 (N_5296,N_4373,N_4953);
nor U5297 (N_5297,N_4452,N_4491);
xnor U5298 (N_5298,N_4979,N_4167);
or U5299 (N_5299,N_4318,N_4278);
or U5300 (N_5300,N_4108,N_4731);
nor U5301 (N_5301,N_4681,N_4630);
nor U5302 (N_5302,N_4843,N_4975);
and U5303 (N_5303,N_4091,N_4204);
nand U5304 (N_5304,N_4511,N_4480);
nor U5305 (N_5305,N_4082,N_4173);
and U5306 (N_5306,N_4612,N_4274);
xnor U5307 (N_5307,N_4758,N_4461);
xor U5308 (N_5308,N_4177,N_4851);
nand U5309 (N_5309,N_4954,N_4113);
nor U5310 (N_5310,N_4999,N_4702);
xnor U5311 (N_5311,N_4052,N_4753);
nand U5312 (N_5312,N_4456,N_4250);
nand U5313 (N_5313,N_4614,N_4754);
or U5314 (N_5314,N_4828,N_4382);
or U5315 (N_5315,N_4486,N_4655);
nand U5316 (N_5316,N_4780,N_4832);
and U5317 (N_5317,N_4981,N_4074);
nand U5318 (N_5318,N_4738,N_4378);
nor U5319 (N_5319,N_4049,N_4146);
nand U5320 (N_5320,N_4713,N_4395);
and U5321 (N_5321,N_4401,N_4138);
and U5322 (N_5322,N_4316,N_4791);
nor U5323 (N_5323,N_4878,N_4720);
nor U5324 (N_5324,N_4315,N_4484);
and U5325 (N_5325,N_4210,N_4716);
nor U5326 (N_5326,N_4202,N_4203);
nor U5327 (N_5327,N_4488,N_4875);
and U5328 (N_5328,N_4631,N_4085);
nand U5329 (N_5329,N_4725,N_4178);
or U5330 (N_5330,N_4175,N_4687);
and U5331 (N_5331,N_4030,N_4990);
xnor U5332 (N_5332,N_4522,N_4249);
nor U5333 (N_5333,N_4866,N_4011);
nand U5334 (N_5334,N_4750,N_4298);
nor U5335 (N_5335,N_4231,N_4654);
and U5336 (N_5336,N_4575,N_4519);
xnor U5337 (N_5337,N_4795,N_4414);
or U5338 (N_5338,N_4568,N_4374);
xnor U5339 (N_5339,N_4225,N_4756);
and U5340 (N_5340,N_4003,N_4586);
xnor U5341 (N_5341,N_4578,N_4099);
or U5342 (N_5342,N_4528,N_4529);
nand U5343 (N_5343,N_4710,N_4856);
nor U5344 (N_5344,N_4520,N_4071);
nand U5345 (N_5345,N_4621,N_4543);
or U5346 (N_5346,N_4741,N_4868);
nor U5347 (N_5347,N_4163,N_4803);
nor U5348 (N_5348,N_4674,N_4946);
and U5349 (N_5349,N_4976,N_4186);
and U5350 (N_5350,N_4013,N_4757);
nor U5351 (N_5351,N_4955,N_4940);
or U5352 (N_5352,N_4936,N_4219);
and U5353 (N_5353,N_4951,N_4006);
xor U5354 (N_5354,N_4633,N_4493);
and U5355 (N_5355,N_4635,N_4782);
or U5356 (N_5356,N_4950,N_4100);
and U5357 (N_5357,N_4650,N_4169);
nand U5358 (N_5358,N_4889,N_4608);
and U5359 (N_5359,N_4445,N_4695);
nand U5360 (N_5360,N_4322,N_4881);
nor U5361 (N_5361,N_4412,N_4406);
or U5362 (N_5362,N_4093,N_4017);
nand U5363 (N_5363,N_4320,N_4909);
or U5364 (N_5364,N_4717,N_4244);
and U5365 (N_5365,N_4882,N_4773);
nand U5366 (N_5366,N_4913,N_4435);
nor U5367 (N_5367,N_4379,N_4694);
xnor U5368 (N_5368,N_4636,N_4237);
and U5369 (N_5369,N_4890,N_4294);
and U5370 (N_5370,N_4540,N_4162);
and U5371 (N_5371,N_4715,N_4693);
nand U5372 (N_5372,N_4684,N_4197);
nand U5373 (N_5373,N_4005,N_4871);
xor U5374 (N_5374,N_4873,N_4727);
nor U5375 (N_5375,N_4923,N_4507);
or U5376 (N_5376,N_4475,N_4996);
nand U5377 (N_5377,N_4942,N_4469);
nand U5378 (N_5378,N_4641,N_4321);
nor U5379 (N_5379,N_4365,N_4324);
nor U5380 (N_5380,N_4329,N_4358);
and U5381 (N_5381,N_4910,N_4312);
nor U5382 (N_5382,N_4344,N_4240);
nand U5383 (N_5383,N_4539,N_4432);
nand U5384 (N_5384,N_4935,N_4447);
and U5385 (N_5385,N_4271,N_4304);
xor U5386 (N_5386,N_4073,N_4961);
or U5387 (N_5387,N_4853,N_4902);
or U5388 (N_5388,N_4036,N_4275);
and U5389 (N_5389,N_4728,N_4798);
and U5390 (N_5390,N_4691,N_4104);
nand U5391 (N_5391,N_4147,N_4106);
xnor U5392 (N_5392,N_4179,N_4489);
nor U5393 (N_5393,N_4538,N_4918);
nor U5394 (N_5394,N_4673,N_4558);
or U5395 (N_5395,N_4026,N_4101);
xnor U5396 (N_5396,N_4451,N_4050);
nor U5397 (N_5397,N_4323,N_4777);
nand U5398 (N_5398,N_4300,N_4545);
nand U5399 (N_5399,N_4424,N_4058);
and U5400 (N_5400,N_4235,N_4552);
and U5401 (N_5401,N_4567,N_4477);
and U5402 (N_5402,N_4763,N_4705);
xnor U5403 (N_5403,N_4425,N_4117);
or U5404 (N_5404,N_4277,N_4385);
xor U5405 (N_5405,N_4453,N_4198);
nand U5406 (N_5406,N_4459,N_4139);
and U5407 (N_5407,N_4464,N_4605);
xor U5408 (N_5408,N_4895,N_4164);
xor U5409 (N_5409,N_4603,N_4389);
nor U5410 (N_5410,N_4084,N_4818);
nand U5411 (N_5411,N_4821,N_4526);
nor U5412 (N_5412,N_4874,N_4525);
and U5413 (N_5413,N_4398,N_4343);
xor U5414 (N_5414,N_4282,N_4218);
nand U5415 (N_5415,N_4581,N_4446);
nor U5416 (N_5416,N_4033,N_4234);
xor U5417 (N_5417,N_4297,N_4041);
xor U5418 (N_5418,N_4174,N_4872);
nor U5419 (N_5419,N_4332,N_4899);
nor U5420 (N_5420,N_4863,N_4784);
xor U5421 (N_5421,N_4579,N_4879);
xnor U5422 (N_5422,N_4497,N_4264);
nor U5423 (N_5423,N_4931,N_4366);
and U5424 (N_5424,N_4012,N_4735);
nand U5425 (N_5425,N_4256,N_4193);
nand U5426 (N_5426,N_4501,N_4845);
nor U5427 (N_5427,N_4269,N_4700);
xor U5428 (N_5428,N_4634,N_4708);
xnor U5429 (N_5429,N_4442,N_4862);
or U5430 (N_5430,N_4880,N_4402);
nor U5431 (N_5431,N_4376,N_4584);
nand U5432 (N_5432,N_4570,N_4917);
and U5433 (N_5433,N_4409,N_4959);
xor U5434 (N_5434,N_4192,N_4478);
xnor U5435 (N_5435,N_4574,N_4787);
xnor U5436 (N_5436,N_4443,N_4467);
nand U5437 (N_5437,N_4711,N_4801);
nor U5438 (N_5438,N_4221,N_4156);
nand U5439 (N_5439,N_4270,N_4034);
or U5440 (N_5440,N_4592,N_4509);
nor U5441 (N_5441,N_4044,N_4510);
nand U5442 (N_5442,N_4356,N_4087);
nor U5443 (N_5443,N_4470,N_4119);
and U5444 (N_5444,N_4503,N_4623);
or U5445 (N_5445,N_4314,N_4252);
xnor U5446 (N_5446,N_4238,N_4550);
xor U5447 (N_5447,N_4182,N_4737);
and U5448 (N_5448,N_4038,N_4517);
or U5449 (N_5449,N_4625,N_4797);
and U5450 (N_5450,N_4670,N_4335);
nand U5451 (N_5451,N_4090,N_4915);
xor U5452 (N_5452,N_4661,N_4561);
or U5453 (N_5453,N_4081,N_4685);
and U5454 (N_5454,N_4686,N_4149);
and U5455 (N_5455,N_4217,N_4247);
or U5456 (N_5456,N_4734,N_4790);
nor U5457 (N_5457,N_4229,N_4860);
or U5458 (N_5458,N_4683,N_4823);
xnor U5459 (N_5459,N_4384,N_4001);
xnor U5460 (N_5460,N_4506,N_4572);
nand U5461 (N_5461,N_4288,N_4914);
nor U5462 (N_5462,N_4672,N_4105);
nor U5463 (N_5463,N_4664,N_4619);
xnor U5464 (N_5464,N_4103,N_4709);
or U5465 (N_5465,N_4948,N_4430);
nand U5466 (N_5466,N_4995,N_4980);
or U5467 (N_5467,N_4769,N_4549);
nand U5468 (N_5468,N_4381,N_4788);
xor U5469 (N_5469,N_4444,N_4404);
nand U5470 (N_5470,N_4176,N_4133);
and U5471 (N_5471,N_4211,N_4696);
nor U5472 (N_5472,N_4647,N_4024);
nand U5473 (N_5473,N_4764,N_4291);
and U5474 (N_5474,N_4441,N_4704);
nor U5475 (N_5475,N_4016,N_4601);
and U5476 (N_5476,N_4072,N_4658);
xnor U5477 (N_5477,N_4559,N_4644);
xor U5478 (N_5478,N_4283,N_4825);
nor U5479 (N_5479,N_4289,N_4888);
or U5480 (N_5480,N_4293,N_4884);
nand U5481 (N_5481,N_4063,N_4301);
or U5482 (N_5482,N_4068,N_4897);
or U5483 (N_5483,N_4831,N_4864);
xnor U5484 (N_5484,N_4692,N_4740);
nand U5485 (N_5485,N_4861,N_4835);
nor U5486 (N_5486,N_4604,N_4599);
nor U5487 (N_5487,N_4336,N_4774);
nor U5488 (N_5488,N_4419,N_4496);
nor U5489 (N_5489,N_4945,N_4311);
and U5490 (N_5490,N_4046,N_4201);
nand U5491 (N_5491,N_4042,N_4472);
or U5492 (N_5492,N_4069,N_4929);
nand U5493 (N_5493,N_4706,N_4665);
xor U5494 (N_5494,N_4056,N_4008);
or U5495 (N_5495,N_4810,N_4077);
and U5496 (N_5496,N_4290,N_4118);
xnor U5497 (N_5497,N_4775,N_4207);
and U5498 (N_5498,N_4964,N_4799);
or U5499 (N_5499,N_4724,N_4014);
and U5500 (N_5500,N_4929,N_4059);
nand U5501 (N_5501,N_4441,N_4007);
nand U5502 (N_5502,N_4463,N_4656);
nor U5503 (N_5503,N_4286,N_4683);
and U5504 (N_5504,N_4057,N_4712);
nor U5505 (N_5505,N_4607,N_4862);
nor U5506 (N_5506,N_4084,N_4759);
nor U5507 (N_5507,N_4430,N_4328);
xnor U5508 (N_5508,N_4339,N_4644);
and U5509 (N_5509,N_4915,N_4505);
or U5510 (N_5510,N_4687,N_4022);
nor U5511 (N_5511,N_4653,N_4614);
or U5512 (N_5512,N_4258,N_4009);
or U5513 (N_5513,N_4539,N_4135);
and U5514 (N_5514,N_4839,N_4390);
xor U5515 (N_5515,N_4164,N_4929);
nand U5516 (N_5516,N_4439,N_4856);
or U5517 (N_5517,N_4052,N_4234);
nand U5518 (N_5518,N_4185,N_4293);
and U5519 (N_5519,N_4358,N_4528);
nor U5520 (N_5520,N_4776,N_4178);
or U5521 (N_5521,N_4880,N_4600);
or U5522 (N_5522,N_4285,N_4529);
and U5523 (N_5523,N_4750,N_4430);
xnor U5524 (N_5524,N_4169,N_4007);
and U5525 (N_5525,N_4139,N_4872);
nor U5526 (N_5526,N_4489,N_4275);
nor U5527 (N_5527,N_4496,N_4935);
nor U5528 (N_5528,N_4860,N_4871);
or U5529 (N_5529,N_4040,N_4667);
and U5530 (N_5530,N_4261,N_4618);
nand U5531 (N_5531,N_4380,N_4526);
nand U5532 (N_5532,N_4694,N_4212);
nand U5533 (N_5533,N_4649,N_4599);
nor U5534 (N_5534,N_4783,N_4454);
nor U5535 (N_5535,N_4251,N_4508);
and U5536 (N_5536,N_4546,N_4762);
and U5537 (N_5537,N_4648,N_4837);
xnor U5538 (N_5538,N_4891,N_4880);
nor U5539 (N_5539,N_4805,N_4774);
nand U5540 (N_5540,N_4312,N_4576);
nand U5541 (N_5541,N_4263,N_4041);
nor U5542 (N_5542,N_4647,N_4370);
xnor U5543 (N_5543,N_4195,N_4446);
nor U5544 (N_5544,N_4900,N_4573);
and U5545 (N_5545,N_4050,N_4661);
xor U5546 (N_5546,N_4851,N_4928);
and U5547 (N_5547,N_4703,N_4230);
nand U5548 (N_5548,N_4804,N_4587);
nand U5549 (N_5549,N_4520,N_4739);
and U5550 (N_5550,N_4994,N_4966);
nor U5551 (N_5551,N_4337,N_4869);
nor U5552 (N_5552,N_4997,N_4459);
nand U5553 (N_5553,N_4978,N_4968);
or U5554 (N_5554,N_4611,N_4092);
or U5555 (N_5555,N_4691,N_4755);
nand U5556 (N_5556,N_4702,N_4232);
nand U5557 (N_5557,N_4195,N_4623);
xnor U5558 (N_5558,N_4490,N_4862);
nand U5559 (N_5559,N_4502,N_4742);
nand U5560 (N_5560,N_4413,N_4950);
or U5561 (N_5561,N_4982,N_4788);
or U5562 (N_5562,N_4761,N_4940);
or U5563 (N_5563,N_4587,N_4015);
xnor U5564 (N_5564,N_4085,N_4030);
nor U5565 (N_5565,N_4108,N_4277);
and U5566 (N_5566,N_4187,N_4617);
xnor U5567 (N_5567,N_4479,N_4734);
nor U5568 (N_5568,N_4296,N_4162);
or U5569 (N_5569,N_4493,N_4065);
or U5570 (N_5570,N_4263,N_4607);
or U5571 (N_5571,N_4432,N_4715);
or U5572 (N_5572,N_4981,N_4893);
nor U5573 (N_5573,N_4718,N_4530);
xor U5574 (N_5574,N_4852,N_4753);
and U5575 (N_5575,N_4697,N_4450);
and U5576 (N_5576,N_4180,N_4735);
xnor U5577 (N_5577,N_4889,N_4252);
or U5578 (N_5578,N_4308,N_4930);
nand U5579 (N_5579,N_4845,N_4747);
and U5580 (N_5580,N_4981,N_4678);
nor U5581 (N_5581,N_4267,N_4310);
or U5582 (N_5582,N_4000,N_4656);
nand U5583 (N_5583,N_4446,N_4067);
or U5584 (N_5584,N_4400,N_4621);
xor U5585 (N_5585,N_4533,N_4101);
xnor U5586 (N_5586,N_4448,N_4060);
and U5587 (N_5587,N_4976,N_4121);
and U5588 (N_5588,N_4089,N_4864);
xnor U5589 (N_5589,N_4536,N_4795);
or U5590 (N_5590,N_4437,N_4133);
or U5591 (N_5591,N_4384,N_4281);
xor U5592 (N_5592,N_4527,N_4696);
nand U5593 (N_5593,N_4123,N_4200);
xor U5594 (N_5594,N_4085,N_4088);
nand U5595 (N_5595,N_4965,N_4583);
nand U5596 (N_5596,N_4542,N_4243);
xor U5597 (N_5597,N_4641,N_4919);
nor U5598 (N_5598,N_4587,N_4425);
and U5599 (N_5599,N_4219,N_4365);
xor U5600 (N_5600,N_4721,N_4226);
or U5601 (N_5601,N_4279,N_4455);
nor U5602 (N_5602,N_4408,N_4974);
nor U5603 (N_5603,N_4843,N_4525);
nand U5604 (N_5604,N_4006,N_4484);
nand U5605 (N_5605,N_4710,N_4201);
nand U5606 (N_5606,N_4073,N_4963);
nand U5607 (N_5607,N_4750,N_4420);
or U5608 (N_5608,N_4901,N_4048);
xnor U5609 (N_5609,N_4359,N_4350);
and U5610 (N_5610,N_4761,N_4997);
and U5611 (N_5611,N_4295,N_4251);
or U5612 (N_5612,N_4567,N_4988);
nor U5613 (N_5613,N_4016,N_4946);
or U5614 (N_5614,N_4909,N_4731);
and U5615 (N_5615,N_4657,N_4470);
nor U5616 (N_5616,N_4397,N_4938);
xor U5617 (N_5617,N_4759,N_4836);
xnor U5618 (N_5618,N_4533,N_4649);
nand U5619 (N_5619,N_4550,N_4593);
xnor U5620 (N_5620,N_4474,N_4674);
or U5621 (N_5621,N_4763,N_4964);
or U5622 (N_5622,N_4456,N_4432);
nor U5623 (N_5623,N_4815,N_4450);
xnor U5624 (N_5624,N_4369,N_4651);
nand U5625 (N_5625,N_4873,N_4976);
nor U5626 (N_5626,N_4323,N_4959);
nand U5627 (N_5627,N_4728,N_4434);
nor U5628 (N_5628,N_4740,N_4371);
nand U5629 (N_5629,N_4927,N_4761);
and U5630 (N_5630,N_4166,N_4707);
nand U5631 (N_5631,N_4218,N_4232);
and U5632 (N_5632,N_4775,N_4798);
xnor U5633 (N_5633,N_4154,N_4893);
xor U5634 (N_5634,N_4496,N_4511);
xnor U5635 (N_5635,N_4715,N_4488);
or U5636 (N_5636,N_4854,N_4462);
or U5637 (N_5637,N_4886,N_4342);
or U5638 (N_5638,N_4485,N_4863);
nor U5639 (N_5639,N_4212,N_4140);
nor U5640 (N_5640,N_4591,N_4422);
xnor U5641 (N_5641,N_4766,N_4741);
nand U5642 (N_5642,N_4903,N_4613);
xor U5643 (N_5643,N_4416,N_4098);
and U5644 (N_5644,N_4954,N_4499);
xnor U5645 (N_5645,N_4834,N_4246);
nand U5646 (N_5646,N_4756,N_4541);
and U5647 (N_5647,N_4021,N_4037);
xnor U5648 (N_5648,N_4569,N_4344);
nand U5649 (N_5649,N_4743,N_4327);
or U5650 (N_5650,N_4960,N_4903);
nand U5651 (N_5651,N_4296,N_4224);
xor U5652 (N_5652,N_4122,N_4910);
nor U5653 (N_5653,N_4806,N_4854);
or U5654 (N_5654,N_4376,N_4442);
nor U5655 (N_5655,N_4747,N_4180);
or U5656 (N_5656,N_4984,N_4708);
nor U5657 (N_5657,N_4056,N_4349);
nand U5658 (N_5658,N_4521,N_4628);
nand U5659 (N_5659,N_4133,N_4245);
or U5660 (N_5660,N_4100,N_4720);
nor U5661 (N_5661,N_4568,N_4887);
nor U5662 (N_5662,N_4454,N_4999);
nand U5663 (N_5663,N_4865,N_4135);
and U5664 (N_5664,N_4566,N_4246);
nand U5665 (N_5665,N_4539,N_4661);
nand U5666 (N_5666,N_4809,N_4163);
nor U5667 (N_5667,N_4240,N_4918);
nor U5668 (N_5668,N_4143,N_4110);
xor U5669 (N_5669,N_4666,N_4988);
or U5670 (N_5670,N_4876,N_4162);
nand U5671 (N_5671,N_4728,N_4228);
and U5672 (N_5672,N_4872,N_4305);
xor U5673 (N_5673,N_4385,N_4565);
nor U5674 (N_5674,N_4085,N_4795);
xnor U5675 (N_5675,N_4749,N_4184);
nand U5676 (N_5676,N_4350,N_4324);
nand U5677 (N_5677,N_4734,N_4729);
xor U5678 (N_5678,N_4866,N_4180);
nand U5679 (N_5679,N_4034,N_4683);
and U5680 (N_5680,N_4785,N_4889);
nor U5681 (N_5681,N_4561,N_4728);
xnor U5682 (N_5682,N_4048,N_4451);
xnor U5683 (N_5683,N_4858,N_4608);
nor U5684 (N_5684,N_4483,N_4315);
nor U5685 (N_5685,N_4128,N_4168);
nor U5686 (N_5686,N_4568,N_4336);
nor U5687 (N_5687,N_4297,N_4646);
and U5688 (N_5688,N_4782,N_4435);
nand U5689 (N_5689,N_4889,N_4496);
nand U5690 (N_5690,N_4529,N_4714);
nand U5691 (N_5691,N_4579,N_4635);
nor U5692 (N_5692,N_4527,N_4252);
xor U5693 (N_5693,N_4828,N_4399);
nor U5694 (N_5694,N_4463,N_4247);
nand U5695 (N_5695,N_4059,N_4279);
and U5696 (N_5696,N_4134,N_4921);
nand U5697 (N_5697,N_4763,N_4837);
nand U5698 (N_5698,N_4257,N_4056);
nand U5699 (N_5699,N_4344,N_4053);
or U5700 (N_5700,N_4104,N_4918);
nand U5701 (N_5701,N_4523,N_4568);
nor U5702 (N_5702,N_4269,N_4871);
nor U5703 (N_5703,N_4959,N_4774);
xor U5704 (N_5704,N_4893,N_4801);
xnor U5705 (N_5705,N_4306,N_4355);
and U5706 (N_5706,N_4256,N_4911);
or U5707 (N_5707,N_4267,N_4749);
and U5708 (N_5708,N_4876,N_4688);
nor U5709 (N_5709,N_4609,N_4389);
nor U5710 (N_5710,N_4699,N_4479);
xor U5711 (N_5711,N_4499,N_4855);
or U5712 (N_5712,N_4495,N_4490);
and U5713 (N_5713,N_4941,N_4613);
nor U5714 (N_5714,N_4186,N_4647);
xor U5715 (N_5715,N_4035,N_4151);
nand U5716 (N_5716,N_4759,N_4529);
xnor U5717 (N_5717,N_4593,N_4272);
xor U5718 (N_5718,N_4632,N_4346);
nand U5719 (N_5719,N_4774,N_4360);
nor U5720 (N_5720,N_4639,N_4596);
or U5721 (N_5721,N_4915,N_4527);
and U5722 (N_5722,N_4433,N_4482);
nand U5723 (N_5723,N_4233,N_4474);
nand U5724 (N_5724,N_4332,N_4576);
nor U5725 (N_5725,N_4883,N_4330);
nand U5726 (N_5726,N_4005,N_4865);
nor U5727 (N_5727,N_4250,N_4710);
nor U5728 (N_5728,N_4760,N_4052);
or U5729 (N_5729,N_4523,N_4264);
nand U5730 (N_5730,N_4799,N_4638);
or U5731 (N_5731,N_4817,N_4257);
nor U5732 (N_5732,N_4114,N_4488);
and U5733 (N_5733,N_4349,N_4204);
xnor U5734 (N_5734,N_4519,N_4463);
or U5735 (N_5735,N_4124,N_4743);
or U5736 (N_5736,N_4858,N_4105);
or U5737 (N_5737,N_4131,N_4890);
and U5738 (N_5738,N_4955,N_4989);
xor U5739 (N_5739,N_4541,N_4584);
nand U5740 (N_5740,N_4327,N_4268);
nor U5741 (N_5741,N_4499,N_4986);
nand U5742 (N_5742,N_4511,N_4917);
nand U5743 (N_5743,N_4148,N_4096);
nand U5744 (N_5744,N_4921,N_4545);
nor U5745 (N_5745,N_4196,N_4323);
or U5746 (N_5746,N_4546,N_4832);
xor U5747 (N_5747,N_4352,N_4223);
xor U5748 (N_5748,N_4549,N_4620);
nand U5749 (N_5749,N_4348,N_4039);
nand U5750 (N_5750,N_4129,N_4737);
and U5751 (N_5751,N_4354,N_4412);
and U5752 (N_5752,N_4530,N_4986);
nand U5753 (N_5753,N_4031,N_4014);
and U5754 (N_5754,N_4017,N_4264);
and U5755 (N_5755,N_4281,N_4177);
xnor U5756 (N_5756,N_4889,N_4759);
or U5757 (N_5757,N_4749,N_4425);
nand U5758 (N_5758,N_4377,N_4738);
or U5759 (N_5759,N_4425,N_4030);
xnor U5760 (N_5760,N_4293,N_4279);
nor U5761 (N_5761,N_4898,N_4121);
nand U5762 (N_5762,N_4244,N_4495);
xnor U5763 (N_5763,N_4556,N_4655);
nor U5764 (N_5764,N_4779,N_4464);
xnor U5765 (N_5765,N_4967,N_4015);
and U5766 (N_5766,N_4180,N_4586);
nor U5767 (N_5767,N_4887,N_4837);
nand U5768 (N_5768,N_4957,N_4178);
or U5769 (N_5769,N_4923,N_4375);
nor U5770 (N_5770,N_4128,N_4843);
nand U5771 (N_5771,N_4132,N_4277);
or U5772 (N_5772,N_4832,N_4141);
or U5773 (N_5773,N_4644,N_4539);
and U5774 (N_5774,N_4756,N_4205);
nand U5775 (N_5775,N_4368,N_4561);
nor U5776 (N_5776,N_4356,N_4423);
nand U5777 (N_5777,N_4248,N_4291);
nand U5778 (N_5778,N_4615,N_4833);
nor U5779 (N_5779,N_4293,N_4367);
or U5780 (N_5780,N_4733,N_4991);
xnor U5781 (N_5781,N_4790,N_4997);
xnor U5782 (N_5782,N_4135,N_4301);
xnor U5783 (N_5783,N_4157,N_4221);
xnor U5784 (N_5784,N_4692,N_4002);
nor U5785 (N_5785,N_4963,N_4184);
or U5786 (N_5786,N_4978,N_4346);
nand U5787 (N_5787,N_4921,N_4769);
nor U5788 (N_5788,N_4520,N_4810);
xor U5789 (N_5789,N_4658,N_4753);
xor U5790 (N_5790,N_4330,N_4121);
or U5791 (N_5791,N_4125,N_4737);
and U5792 (N_5792,N_4084,N_4878);
xor U5793 (N_5793,N_4474,N_4943);
or U5794 (N_5794,N_4975,N_4984);
nor U5795 (N_5795,N_4203,N_4007);
xnor U5796 (N_5796,N_4897,N_4905);
or U5797 (N_5797,N_4647,N_4833);
or U5798 (N_5798,N_4059,N_4508);
or U5799 (N_5799,N_4888,N_4910);
xor U5800 (N_5800,N_4411,N_4120);
xor U5801 (N_5801,N_4916,N_4081);
nand U5802 (N_5802,N_4211,N_4997);
nand U5803 (N_5803,N_4445,N_4123);
and U5804 (N_5804,N_4014,N_4601);
and U5805 (N_5805,N_4946,N_4083);
nor U5806 (N_5806,N_4268,N_4145);
xor U5807 (N_5807,N_4349,N_4260);
and U5808 (N_5808,N_4553,N_4055);
xnor U5809 (N_5809,N_4604,N_4788);
xnor U5810 (N_5810,N_4848,N_4659);
nand U5811 (N_5811,N_4184,N_4397);
nor U5812 (N_5812,N_4499,N_4504);
and U5813 (N_5813,N_4226,N_4154);
nor U5814 (N_5814,N_4603,N_4899);
or U5815 (N_5815,N_4134,N_4089);
and U5816 (N_5816,N_4076,N_4347);
or U5817 (N_5817,N_4968,N_4100);
or U5818 (N_5818,N_4971,N_4024);
or U5819 (N_5819,N_4566,N_4538);
xor U5820 (N_5820,N_4051,N_4254);
nor U5821 (N_5821,N_4334,N_4576);
xor U5822 (N_5822,N_4200,N_4950);
and U5823 (N_5823,N_4069,N_4280);
nand U5824 (N_5824,N_4016,N_4712);
or U5825 (N_5825,N_4008,N_4222);
nand U5826 (N_5826,N_4530,N_4024);
xnor U5827 (N_5827,N_4054,N_4339);
xor U5828 (N_5828,N_4929,N_4941);
xnor U5829 (N_5829,N_4052,N_4684);
nand U5830 (N_5830,N_4567,N_4254);
nor U5831 (N_5831,N_4803,N_4644);
xnor U5832 (N_5832,N_4214,N_4739);
xnor U5833 (N_5833,N_4374,N_4556);
nor U5834 (N_5834,N_4698,N_4411);
xor U5835 (N_5835,N_4927,N_4911);
xnor U5836 (N_5836,N_4752,N_4720);
and U5837 (N_5837,N_4417,N_4788);
nor U5838 (N_5838,N_4639,N_4688);
and U5839 (N_5839,N_4956,N_4532);
xnor U5840 (N_5840,N_4778,N_4223);
nor U5841 (N_5841,N_4204,N_4205);
and U5842 (N_5842,N_4112,N_4587);
nor U5843 (N_5843,N_4967,N_4125);
nor U5844 (N_5844,N_4242,N_4236);
xnor U5845 (N_5845,N_4883,N_4812);
xor U5846 (N_5846,N_4784,N_4088);
xnor U5847 (N_5847,N_4850,N_4039);
xnor U5848 (N_5848,N_4500,N_4579);
nor U5849 (N_5849,N_4480,N_4182);
or U5850 (N_5850,N_4170,N_4090);
nand U5851 (N_5851,N_4432,N_4515);
xor U5852 (N_5852,N_4756,N_4610);
nor U5853 (N_5853,N_4304,N_4819);
nand U5854 (N_5854,N_4172,N_4396);
xor U5855 (N_5855,N_4132,N_4279);
xor U5856 (N_5856,N_4533,N_4726);
nor U5857 (N_5857,N_4589,N_4093);
or U5858 (N_5858,N_4241,N_4181);
and U5859 (N_5859,N_4954,N_4912);
or U5860 (N_5860,N_4518,N_4609);
xnor U5861 (N_5861,N_4876,N_4662);
or U5862 (N_5862,N_4301,N_4274);
xor U5863 (N_5863,N_4219,N_4186);
and U5864 (N_5864,N_4966,N_4475);
xor U5865 (N_5865,N_4866,N_4099);
nor U5866 (N_5866,N_4530,N_4913);
nand U5867 (N_5867,N_4004,N_4649);
or U5868 (N_5868,N_4962,N_4870);
or U5869 (N_5869,N_4701,N_4086);
nand U5870 (N_5870,N_4737,N_4238);
nor U5871 (N_5871,N_4126,N_4638);
nand U5872 (N_5872,N_4054,N_4795);
and U5873 (N_5873,N_4192,N_4214);
xor U5874 (N_5874,N_4751,N_4597);
xor U5875 (N_5875,N_4117,N_4630);
nand U5876 (N_5876,N_4287,N_4434);
nand U5877 (N_5877,N_4885,N_4573);
or U5878 (N_5878,N_4173,N_4408);
xor U5879 (N_5879,N_4005,N_4785);
and U5880 (N_5880,N_4761,N_4290);
xnor U5881 (N_5881,N_4104,N_4432);
nand U5882 (N_5882,N_4820,N_4597);
nand U5883 (N_5883,N_4908,N_4065);
nand U5884 (N_5884,N_4573,N_4949);
and U5885 (N_5885,N_4742,N_4884);
xor U5886 (N_5886,N_4608,N_4366);
and U5887 (N_5887,N_4245,N_4970);
nand U5888 (N_5888,N_4355,N_4236);
or U5889 (N_5889,N_4296,N_4181);
nand U5890 (N_5890,N_4602,N_4621);
xnor U5891 (N_5891,N_4929,N_4938);
or U5892 (N_5892,N_4085,N_4620);
nor U5893 (N_5893,N_4486,N_4639);
nor U5894 (N_5894,N_4897,N_4821);
nor U5895 (N_5895,N_4852,N_4029);
nand U5896 (N_5896,N_4582,N_4120);
or U5897 (N_5897,N_4181,N_4119);
nor U5898 (N_5898,N_4303,N_4285);
and U5899 (N_5899,N_4571,N_4417);
or U5900 (N_5900,N_4571,N_4849);
xor U5901 (N_5901,N_4638,N_4869);
nor U5902 (N_5902,N_4257,N_4726);
and U5903 (N_5903,N_4864,N_4443);
or U5904 (N_5904,N_4260,N_4293);
xnor U5905 (N_5905,N_4545,N_4740);
nand U5906 (N_5906,N_4339,N_4637);
or U5907 (N_5907,N_4366,N_4895);
nor U5908 (N_5908,N_4972,N_4242);
or U5909 (N_5909,N_4453,N_4101);
or U5910 (N_5910,N_4613,N_4909);
nand U5911 (N_5911,N_4659,N_4983);
xnor U5912 (N_5912,N_4064,N_4236);
xnor U5913 (N_5913,N_4957,N_4644);
or U5914 (N_5914,N_4792,N_4159);
nand U5915 (N_5915,N_4854,N_4711);
or U5916 (N_5916,N_4875,N_4274);
nand U5917 (N_5917,N_4839,N_4466);
xor U5918 (N_5918,N_4043,N_4158);
nand U5919 (N_5919,N_4555,N_4576);
nor U5920 (N_5920,N_4401,N_4692);
nor U5921 (N_5921,N_4084,N_4710);
nand U5922 (N_5922,N_4311,N_4609);
or U5923 (N_5923,N_4612,N_4870);
or U5924 (N_5924,N_4180,N_4978);
xor U5925 (N_5925,N_4191,N_4651);
nand U5926 (N_5926,N_4419,N_4128);
nor U5927 (N_5927,N_4907,N_4937);
xnor U5928 (N_5928,N_4446,N_4494);
nor U5929 (N_5929,N_4416,N_4498);
and U5930 (N_5930,N_4455,N_4276);
or U5931 (N_5931,N_4482,N_4769);
and U5932 (N_5932,N_4487,N_4964);
nor U5933 (N_5933,N_4412,N_4624);
nor U5934 (N_5934,N_4179,N_4285);
or U5935 (N_5935,N_4901,N_4704);
or U5936 (N_5936,N_4029,N_4034);
or U5937 (N_5937,N_4524,N_4575);
or U5938 (N_5938,N_4000,N_4707);
xor U5939 (N_5939,N_4829,N_4096);
or U5940 (N_5940,N_4765,N_4443);
or U5941 (N_5941,N_4471,N_4422);
or U5942 (N_5942,N_4533,N_4106);
xor U5943 (N_5943,N_4364,N_4495);
and U5944 (N_5944,N_4706,N_4943);
nor U5945 (N_5945,N_4098,N_4113);
xor U5946 (N_5946,N_4151,N_4616);
nor U5947 (N_5947,N_4664,N_4013);
xnor U5948 (N_5948,N_4997,N_4983);
and U5949 (N_5949,N_4089,N_4367);
xor U5950 (N_5950,N_4197,N_4382);
and U5951 (N_5951,N_4796,N_4662);
xnor U5952 (N_5952,N_4988,N_4327);
nand U5953 (N_5953,N_4724,N_4686);
and U5954 (N_5954,N_4297,N_4568);
and U5955 (N_5955,N_4668,N_4393);
nand U5956 (N_5956,N_4588,N_4976);
nand U5957 (N_5957,N_4194,N_4975);
and U5958 (N_5958,N_4596,N_4276);
xor U5959 (N_5959,N_4907,N_4332);
and U5960 (N_5960,N_4751,N_4401);
nand U5961 (N_5961,N_4243,N_4325);
and U5962 (N_5962,N_4979,N_4373);
nand U5963 (N_5963,N_4225,N_4624);
nor U5964 (N_5964,N_4794,N_4175);
or U5965 (N_5965,N_4088,N_4410);
nor U5966 (N_5966,N_4361,N_4409);
nor U5967 (N_5967,N_4080,N_4245);
xnor U5968 (N_5968,N_4140,N_4532);
or U5969 (N_5969,N_4665,N_4173);
or U5970 (N_5970,N_4166,N_4508);
and U5971 (N_5971,N_4122,N_4812);
nand U5972 (N_5972,N_4606,N_4891);
or U5973 (N_5973,N_4878,N_4450);
nand U5974 (N_5974,N_4133,N_4432);
xnor U5975 (N_5975,N_4067,N_4962);
nand U5976 (N_5976,N_4310,N_4660);
or U5977 (N_5977,N_4555,N_4635);
xor U5978 (N_5978,N_4969,N_4288);
xor U5979 (N_5979,N_4269,N_4333);
nor U5980 (N_5980,N_4330,N_4043);
or U5981 (N_5981,N_4118,N_4723);
nand U5982 (N_5982,N_4506,N_4798);
and U5983 (N_5983,N_4817,N_4528);
or U5984 (N_5984,N_4136,N_4787);
or U5985 (N_5985,N_4295,N_4112);
and U5986 (N_5986,N_4141,N_4359);
and U5987 (N_5987,N_4239,N_4356);
and U5988 (N_5988,N_4188,N_4418);
and U5989 (N_5989,N_4875,N_4347);
nand U5990 (N_5990,N_4953,N_4622);
nand U5991 (N_5991,N_4795,N_4746);
or U5992 (N_5992,N_4423,N_4136);
nand U5993 (N_5993,N_4548,N_4872);
and U5994 (N_5994,N_4562,N_4607);
nor U5995 (N_5995,N_4122,N_4372);
nand U5996 (N_5996,N_4879,N_4872);
nand U5997 (N_5997,N_4361,N_4310);
or U5998 (N_5998,N_4896,N_4234);
or U5999 (N_5999,N_4034,N_4003);
and U6000 (N_6000,N_5308,N_5093);
nor U6001 (N_6001,N_5259,N_5020);
or U6002 (N_6002,N_5380,N_5948);
or U6003 (N_6003,N_5954,N_5088);
or U6004 (N_6004,N_5518,N_5435);
nand U6005 (N_6005,N_5075,N_5237);
xnor U6006 (N_6006,N_5058,N_5289);
nand U6007 (N_6007,N_5723,N_5735);
xnor U6008 (N_6008,N_5270,N_5655);
and U6009 (N_6009,N_5038,N_5727);
and U6010 (N_6010,N_5324,N_5149);
xnor U6011 (N_6011,N_5654,N_5448);
or U6012 (N_6012,N_5214,N_5756);
nand U6013 (N_6013,N_5597,N_5783);
nor U6014 (N_6014,N_5244,N_5957);
xor U6015 (N_6015,N_5011,N_5072);
nor U6016 (N_6016,N_5901,N_5496);
nand U6017 (N_6017,N_5123,N_5992);
xor U6018 (N_6018,N_5771,N_5577);
or U6019 (N_6019,N_5708,N_5223);
and U6020 (N_6020,N_5154,N_5995);
nand U6021 (N_6021,N_5725,N_5478);
xor U6022 (N_6022,N_5543,N_5079);
or U6023 (N_6023,N_5297,N_5379);
nor U6024 (N_6024,N_5494,N_5489);
nand U6025 (N_6025,N_5200,N_5357);
and U6026 (N_6026,N_5348,N_5017);
and U6027 (N_6027,N_5918,N_5211);
nor U6028 (N_6028,N_5636,N_5552);
nand U6029 (N_6029,N_5943,N_5016);
or U6030 (N_6030,N_5061,N_5547);
nor U6031 (N_6031,N_5526,N_5871);
or U6032 (N_6032,N_5103,N_5599);
and U6033 (N_6033,N_5483,N_5978);
and U6034 (N_6034,N_5553,N_5907);
xnor U6035 (N_6035,N_5836,N_5902);
nand U6036 (N_6036,N_5680,N_5962);
xnor U6037 (N_6037,N_5492,N_5293);
xor U6038 (N_6038,N_5777,N_5831);
nand U6039 (N_6039,N_5356,N_5290);
nand U6040 (N_6040,N_5117,N_5609);
xnor U6041 (N_6041,N_5516,N_5094);
nor U6042 (N_6042,N_5544,N_5828);
nor U6043 (N_6043,N_5911,N_5732);
xor U6044 (N_6044,N_5841,N_5386);
or U6045 (N_6045,N_5999,N_5459);
nand U6046 (N_6046,N_5268,N_5743);
and U6047 (N_6047,N_5177,N_5082);
xor U6048 (N_6048,N_5051,N_5022);
xor U6049 (N_6049,N_5908,N_5003);
or U6050 (N_6050,N_5903,N_5315);
or U6051 (N_6051,N_5261,N_5277);
nand U6052 (N_6052,N_5984,N_5173);
and U6053 (N_6053,N_5452,N_5833);
and U6054 (N_6054,N_5640,N_5165);
and U6055 (N_6055,N_5081,N_5970);
or U6056 (N_6056,N_5114,N_5747);
and U6057 (N_6057,N_5624,N_5646);
and U6058 (N_6058,N_5586,N_5398);
xor U6059 (N_6059,N_5759,N_5784);
xnor U6060 (N_6060,N_5899,N_5741);
or U6061 (N_6061,N_5717,N_5955);
and U6062 (N_6062,N_5536,N_5920);
nand U6063 (N_6063,N_5569,N_5998);
and U6064 (N_6064,N_5721,N_5730);
or U6065 (N_6065,N_5449,N_5420);
nor U6066 (N_6066,N_5990,N_5115);
and U6067 (N_6067,N_5855,N_5442);
nor U6068 (N_6068,N_5795,N_5642);
and U6069 (N_6069,N_5931,N_5753);
and U6070 (N_6070,N_5385,N_5749);
or U6071 (N_6071,N_5568,N_5222);
and U6072 (N_6072,N_5235,N_5085);
or U6073 (N_6073,N_5711,N_5703);
xor U6074 (N_6074,N_5037,N_5378);
or U6075 (N_6075,N_5965,N_5921);
xor U6076 (N_6076,N_5362,N_5869);
nor U6077 (N_6077,N_5824,N_5738);
nor U6078 (N_6078,N_5505,N_5197);
or U6079 (N_6079,N_5272,N_5258);
or U6080 (N_6080,N_5034,N_5458);
xor U6081 (N_6081,N_5584,N_5558);
and U6082 (N_6082,N_5335,N_5986);
nand U6083 (N_6083,N_5201,N_5195);
nor U6084 (N_6084,N_5819,N_5572);
xnor U6085 (N_6085,N_5212,N_5292);
nor U6086 (N_6086,N_5215,N_5065);
xnor U6087 (N_6087,N_5626,N_5856);
or U6088 (N_6088,N_5439,N_5161);
nor U6089 (N_6089,N_5073,N_5612);
nor U6090 (N_6090,N_5470,N_5371);
xor U6091 (N_6091,N_5410,N_5347);
xnor U6092 (N_6092,N_5790,N_5092);
nor U6093 (N_6093,N_5789,N_5909);
or U6094 (N_6094,N_5438,N_5787);
nand U6095 (N_6095,N_5893,N_5502);
nor U6096 (N_6096,N_5987,N_5567);
and U6097 (N_6097,N_5677,N_5321);
xnor U6098 (N_6098,N_5664,N_5613);
nor U6099 (N_6099,N_5469,N_5676);
xnor U6100 (N_6100,N_5495,N_5110);
or U6101 (N_6101,N_5155,N_5375);
xnor U6102 (N_6102,N_5415,N_5178);
xnor U6103 (N_6103,N_5394,N_5830);
nor U6104 (N_6104,N_5129,N_5762);
and U6105 (N_6105,N_5157,N_5620);
nor U6106 (N_6106,N_5766,N_5808);
nor U6107 (N_6107,N_5576,N_5694);
or U6108 (N_6108,N_5773,N_5108);
or U6109 (N_6109,N_5089,N_5528);
xor U6110 (N_6110,N_5910,N_5596);
nand U6111 (N_6111,N_5797,N_5167);
and U6112 (N_6112,N_5997,N_5994);
or U6113 (N_6113,N_5281,N_5062);
xnor U6114 (N_6114,N_5132,N_5228);
and U6115 (N_6115,N_5772,N_5653);
or U6116 (N_6116,N_5846,N_5419);
and U6117 (N_6117,N_5594,N_5447);
nor U6118 (N_6118,N_5305,N_5796);
nand U6119 (N_6119,N_5809,N_5971);
nand U6120 (N_6120,N_5794,N_5045);
nand U6121 (N_6121,N_5360,N_5206);
nor U6122 (N_6122,N_5414,N_5296);
nor U6123 (N_6123,N_5387,N_5174);
and U6124 (N_6124,N_5951,N_5639);
and U6125 (N_6125,N_5358,N_5896);
nand U6126 (N_6126,N_5456,N_5504);
nand U6127 (N_6127,N_5002,N_5040);
nor U6128 (N_6128,N_5928,N_5905);
nand U6129 (N_6129,N_5813,N_5012);
or U6130 (N_6130,N_5121,N_5059);
nor U6131 (N_6131,N_5637,N_5183);
xor U6132 (N_6132,N_5162,N_5629);
or U6133 (N_6133,N_5670,N_5473);
nor U6134 (N_6134,N_5499,N_5712);
nor U6135 (N_6135,N_5158,N_5980);
or U6136 (N_6136,N_5417,N_5254);
nor U6137 (N_6137,N_5327,N_5926);
or U6138 (N_6138,N_5118,N_5932);
and U6139 (N_6139,N_5207,N_5399);
xor U6140 (N_6140,N_5878,N_5803);
xor U6141 (N_6141,N_5649,N_5275);
or U6142 (N_6142,N_5539,N_5825);
nand U6143 (N_6143,N_5815,N_5311);
or U6144 (N_6144,N_5648,N_5390);
and U6145 (N_6145,N_5798,N_5243);
nand U6146 (N_6146,N_5940,N_5843);
or U6147 (N_6147,N_5616,N_5203);
nand U6148 (N_6148,N_5729,N_5904);
nand U6149 (N_6149,N_5491,N_5559);
nand U6150 (N_6150,N_5239,N_5780);
xor U6151 (N_6151,N_5184,N_5355);
nor U6152 (N_6152,N_5601,N_5872);
nand U6153 (N_6153,N_5310,N_5128);
nand U6154 (N_6154,N_5287,N_5106);
xor U6155 (N_6155,N_5044,N_5460);
nand U6156 (N_6156,N_5508,N_5800);
xnor U6157 (N_6157,N_5169,N_5067);
and U6158 (N_6158,N_5334,N_5615);
nor U6159 (N_6159,N_5715,N_5295);
and U6160 (N_6160,N_5963,N_5163);
nor U6161 (N_6161,N_5823,N_5849);
and U6162 (N_6162,N_5506,N_5028);
xnor U6163 (N_6163,N_5860,N_5430);
and U6164 (N_6164,N_5500,N_5710);
nand U6165 (N_6165,N_5929,N_5959);
nor U6166 (N_6166,N_5561,N_5775);
or U6167 (N_6167,N_5168,N_5472);
and U6168 (N_6168,N_5534,N_5036);
and U6169 (N_6169,N_5481,N_5428);
or U6170 (N_6170,N_5373,N_5190);
or U6171 (N_6171,N_5352,N_5033);
and U6172 (N_6172,N_5070,N_5592);
xor U6173 (N_6173,N_5486,N_5488);
nand U6174 (N_6174,N_5923,N_5706);
nand U6175 (N_6175,N_5066,N_5441);
nor U6176 (N_6176,N_5328,N_5540);
nor U6177 (N_6177,N_5274,N_5213);
nand U6178 (N_6178,N_5917,N_5793);
or U6179 (N_6179,N_5194,N_5216);
nor U6180 (N_6180,N_5988,N_5053);
nand U6181 (N_6181,N_5052,N_5048);
nor U6182 (N_6182,N_5811,N_5925);
xor U6183 (N_6183,N_5827,N_5152);
nor U6184 (N_6184,N_5665,N_5098);
xnor U6185 (N_6185,N_5886,N_5989);
nand U6186 (N_6186,N_5076,N_5018);
or U6187 (N_6187,N_5331,N_5768);
xnor U6188 (N_6188,N_5231,N_5208);
or U6189 (N_6189,N_5429,N_5468);
nor U6190 (N_6190,N_5060,N_5588);
nand U6191 (N_6191,N_5204,N_5443);
xnor U6192 (N_6192,N_5047,N_5069);
xor U6193 (N_6193,N_5234,N_5175);
xnor U6194 (N_6194,N_5884,N_5031);
nand U6195 (N_6195,N_5090,N_5550);
or U6196 (N_6196,N_5143,N_5832);
nor U6197 (N_6197,N_5890,N_5366);
nor U6198 (N_6198,N_5564,N_5638);
xnor U6199 (N_6199,N_5202,N_5377);
nor U6200 (N_6200,N_5936,N_5196);
nand U6201 (N_6201,N_5474,N_5546);
nand U6202 (N_6202,N_5865,N_5912);
and U6203 (N_6203,N_5320,N_5264);
nor U6204 (N_6204,N_5977,N_5961);
xor U6205 (N_6205,N_5151,N_5139);
or U6206 (N_6206,N_5960,N_5107);
or U6207 (N_6207,N_5482,N_5937);
nand U6208 (N_6208,N_5218,N_5187);
nand U6209 (N_6209,N_5758,N_5513);
nand U6210 (N_6210,N_5510,N_5792);
xor U6211 (N_6211,N_5341,N_5454);
nor U6212 (N_6212,N_5266,N_5050);
nand U6213 (N_6213,N_5545,N_5217);
xor U6214 (N_6214,N_5691,N_5906);
xnor U6215 (N_6215,N_5019,N_5185);
or U6216 (N_6216,N_5278,N_5120);
nor U6217 (N_6217,N_5681,N_5240);
and U6218 (N_6218,N_5463,N_5126);
nand U6219 (N_6219,N_5520,N_5384);
and U6220 (N_6220,N_5563,N_5063);
nand U6221 (N_6221,N_5844,N_5104);
and U6222 (N_6222,N_5186,N_5628);
nor U6223 (N_6223,N_5260,N_5299);
nor U6224 (N_6224,N_5336,N_5351);
or U6225 (N_6225,N_5140,N_5845);
nor U6226 (N_6226,N_5249,N_5630);
nand U6227 (N_6227,N_5300,N_5156);
xor U6228 (N_6228,N_5535,N_5317);
xnor U6229 (N_6229,N_5400,N_5560);
xnor U6230 (N_6230,N_5892,N_5924);
xnor U6231 (N_6231,N_5647,N_5096);
nand U6232 (N_6232,N_5226,N_5898);
nand U6233 (N_6233,N_5256,N_5403);
xnor U6234 (N_6234,N_5130,N_5382);
xnor U6235 (N_6235,N_5074,N_5407);
xnor U6236 (N_6236,N_5661,N_5799);
and U6237 (N_6237,N_5250,N_5507);
xnor U6238 (N_6238,N_5742,N_5303);
xnor U6239 (N_6239,N_5698,N_5883);
and U6240 (N_6240,N_5575,N_5457);
nand U6241 (N_6241,N_5580,N_5779);
nor U6242 (N_6242,N_5286,N_5137);
nand U6243 (N_6243,N_5097,N_5982);
or U6244 (N_6244,N_5748,N_5643);
or U6245 (N_6245,N_5557,N_5531);
or U6246 (N_6246,N_5595,N_5659);
and U6247 (N_6247,N_5182,N_5555);
nor U6248 (N_6248,N_5881,N_5556);
nor U6249 (N_6249,N_5273,N_5949);
or U6250 (N_6250,N_5330,N_5985);
or U6251 (N_6251,N_5025,N_5326);
or U6252 (N_6252,N_5125,N_5876);
or U6253 (N_6253,N_5861,N_5238);
or U6254 (N_6254,N_5867,N_5422);
nor U6255 (N_6255,N_5440,N_5975);
nand U6256 (N_6256,N_5105,N_5271);
and U6257 (N_6257,N_5100,N_5688);
xnor U6258 (N_6258,N_5391,N_5645);
nand U6259 (N_6259,N_5078,N_5683);
and U6260 (N_6260,N_5532,N_5523);
xnor U6261 (N_6261,N_5512,N_5029);
xnor U6262 (N_6262,N_5786,N_5820);
nand U6263 (N_6263,N_5685,N_5068);
and U6264 (N_6264,N_5170,N_5605);
or U6265 (N_6265,N_5004,N_5578);
nand U6266 (N_6266,N_5342,N_5702);
nand U6267 (N_6267,N_5119,N_5947);
and U6268 (N_6268,N_5493,N_5774);
nand U6269 (N_6269,N_5421,N_5247);
xnor U6270 (N_6270,N_5604,N_5080);
or U6271 (N_6271,N_5434,N_5229);
nor U6272 (N_6272,N_5625,N_5205);
nand U6273 (N_6273,N_5848,N_5858);
and U6274 (N_6274,N_5144,N_5622);
nor U6275 (N_6275,N_5739,N_5445);
nor U6276 (N_6276,N_5188,N_5381);
or U6277 (N_6277,N_5581,N_5301);
nor U6278 (N_6278,N_5087,N_5109);
and U6279 (N_6279,N_5245,N_5122);
xnor U6280 (N_6280,N_5635,N_5304);
and U6281 (N_6281,N_5209,N_5726);
nor U6282 (N_6282,N_5953,N_5866);
and U6283 (N_6283,N_5674,N_5746);
nand U6284 (N_6284,N_5695,N_5363);
or U6285 (N_6285,N_5714,N_5853);
xor U6286 (N_6286,N_5554,N_5590);
and U6287 (N_6287,N_5537,N_5424);
xnor U6288 (N_6288,N_5367,N_5525);
or U6289 (N_6289,N_5210,N_5340);
nor U6290 (N_6290,N_5383,N_5690);
nand U6291 (N_6291,N_5043,N_5733);
xnor U6292 (N_6292,N_5322,N_5225);
nand U6293 (N_6293,N_5810,N_5147);
and U6294 (N_6294,N_5538,N_5964);
and U6295 (N_6295,N_5574,N_5704);
xor U6296 (N_6296,N_5579,N_5166);
nand U6297 (N_6297,N_5847,N_5198);
or U6298 (N_6298,N_5319,N_5687);
xor U6299 (N_6299,N_5333,N_5376);
and U6300 (N_6300,N_5679,N_5111);
xor U6301 (N_6301,N_5142,N_5306);
xnor U6302 (N_6302,N_5600,N_5889);
nand U6303 (N_6303,N_5973,N_5877);
and U6304 (N_6304,N_5408,N_5541);
or U6305 (N_6305,N_5781,N_5611);
xor U6306 (N_6306,N_5433,N_5956);
and U6307 (N_6307,N_5934,N_5669);
nand U6308 (N_6308,N_5406,N_5263);
nor U6309 (N_6309,N_5055,N_5436);
and U6310 (N_6310,N_5700,N_5979);
or U6311 (N_6311,N_5221,N_5475);
nand U6312 (N_6312,N_5551,N_5148);
and U6313 (N_6313,N_5049,N_5870);
nand U6314 (N_6314,N_5112,N_5631);
xnor U6315 (N_6315,N_5945,N_5701);
or U6316 (N_6316,N_5778,N_5752);
xor U6317 (N_6317,N_5427,N_5927);
or U6318 (N_6318,N_5246,N_5967);
xnor U6319 (N_6319,N_5007,N_5042);
or U6320 (N_6320,N_5302,N_5232);
nor U6321 (N_6321,N_5252,N_5672);
nand U6322 (N_6322,N_5852,N_5193);
or U6323 (N_6323,N_5369,N_5818);
and U6324 (N_6324,N_5822,N_5915);
nand U6325 (N_6325,N_5757,N_5423);
nor U6326 (N_6326,N_5192,N_5750);
xor U6327 (N_6327,N_5533,N_5318);
and U6328 (N_6328,N_5969,N_5325);
xnor U6329 (N_6329,N_5807,N_5431);
and U6330 (N_6330,N_5737,N_5751);
or U6331 (N_6331,N_5868,N_5933);
and U6332 (N_6332,N_5656,N_5220);
nor U6333 (N_6333,N_5313,N_5393);
xnor U6334 (N_6334,N_5498,N_5501);
nor U6335 (N_6335,N_5077,N_5996);
nand U6336 (N_6336,N_5233,N_5451);
nand U6337 (N_6337,N_5138,N_5851);
or U6338 (N_6338,N_5337,N_5895);
nor U6339 (N_6339,N_5692,N_5983);
xnor U6340 (N_6340,N_5740,N_5663);
nand U6341 (N_6341,N_5864,N_5562);
nand U6342 (N_6342,N_5136,N_5859);
or U6343 (N_6343,N_5345,N_5124);
nor U6344 (N_6344,N_5548,N_5972);
nor U6345 (N_6345,N_5484,N_5368);
or U6346 (N_6346,N_5842,N_5039);
xor U6347 (N_6347,N_5279,N_5689);
xor U6348 (N_6348,N_5280,N_5718);
or U6349 (N_6349,N_5135,N_5455);
nor U6350 (N_6350,N_5409,N_5432);
xor U6351 (N_6351,N_5662,N_5976);
xor U6352 (N_6352,N_5660,N_5159);
and U6353 (N_6353,N_5879,N_5658);
xnor U6354 (N_6354,N_5461,N_5573);
xnor U6355 (N_6355,N_5941,N_5641);
nor U6356 (N_6356,N_5064,N_5854);
or U6357 (N_6357,N_5744,N_5071);
nand U6358 (N_6358,N_5897,N_5265);
xor U6359 (N_6359,N_5791,N_5565);
nor U6360 (N_6360,N_5219,N_5008);
nand U6361 (N_6361,N_5444,N_5816);
nand U6362 (N_6362,N_5000,N_5767);
or U6363 (N_6363,N_5010,N_5462);
or U6364 (N_6364,N_5530,N_5521);
xor U6365 (N_6365,N_5465,N_5009);
xor U6366 (N_6366,N_5402,N_5316);
and U6367 (N_6367,N_5527,N_5453);
or U6368 (N_6368,N_5764,N_5919);
or U6369 (N_6369,N_5644,N_5682);
or U6370 (N_6370,N_5479,N_5607);
nand U6371 (N_6371,N_5671,N_5770);
and U6372 (N_6372,N_5916,N_5763);
nand U6373 (N_6373,N_5623,N_5805);
xor U6374 (N_6374,N_5519,N_5046);
xnor U6375 (N_6375,N_5614,N_5814);
and U6376 (N_6376,N_5511,N_5283);
xor U6377 (N_6377,N_5248,N_5591);
or U6378 (N_6378,N_5392,N_5678);
or U6379 (N_6379,N_5801,N_5728);
nand U6380 (N_6380,N_5617,N_5696);
and U6381 (N_6381,N_5372,N_5418);
or U6382 (N_6382,N_5838,N_5875);
or U6383 (N_6383,N_5935,N_5922);
nor U6384 (N_6384,N_5298,N_5282);
and U6385 (N_6385,N_5888,N_5338);
nand U6386 (N_6386,N_5788,N_5515);
xor U6387 (N_6387,N_5891,N_5359);
nand U6388 (N_6388,N_5632,N_5862);
nor U6389 (N_6389,N_5610,N_5745);
and U6390 (N_6390,N_5146,N_5404);
and U6391 (N_6391,N_5131,N_5736);
nor U6392 (N_6392,N_5666,N_5285);
nor U6393 (N_6393,N_5015,N_5765);
nor U6394 (N_6394,N_5307,N_5191);
nand U6395 (N_6395,N_5834,N_5621);
xnor U6396 (N_6396,N_5388,N_5199);
xnor U6397 (N_6397,N_5769,N_5113);
xor U6398 (N_6398,N_5241,N_5724);
or U6399 (N_6399,N_5413,N_5716);
and U6400 (N_6400,N_5652,N_5668);
and U6401 (N_6401,N_5583,N_5412);
nor U6402 (N_6402,N_5312,N_5755);
nor U6403 (N_6403,N_5958,N_5099);
nand U6404 (N_6404,N_5180,N_5024);
and U6405 (N_6405,N_5026,N_5942);
nor U6406 (N_6406,N_5880,N_5056);
or U6407 (N_6407,N_5734,N_5806);
nor U6408 (N_6408,N_5343,N_5731);
and U6409 (N_6409,N_5582,N_5657);
or U6410 (N_6410,N_5837,N_5840);
or U6411 (N_6411,N_5450,N_5416);
and U6412 (N_6412,N_5032,N_5314);
or U6413 (N_6413,N_5405,N_5116);
xor U6414 (N_6414,N_5464,N_5346);
nor U6415 (N_6415,N_5164,N_5587);
nor U6416 (N_6416,N_5160,N_5517);
nand U6417 (N_6417,N_5618,N_5329);
nand U6418 (N_6418,N_5236,N_5914);
nor U6419 (N_6419,N_5471,N_5005);
or U6420 (N_6420,N_5598,N_5633);
nand U6421 (N_6421,N_5882,N_5821);
or U6422 (N_6422,N_5086,N_5585);
xor U6423 (N_6423,N_5467,N_5176);
xor U6424 (N_6424,N_5608,N_5485);
xnor U6425 (N_6425,N_5013,N_5411);
and U6426 (N_6426,N_5675,N_5361);
or U6427 (N_6427,N_5030,N_5476);
xnor U6428 (N_6428,N_5968,N_5401);
or U6429 (N_6429,N_5446,N_5057);
nand U6430 (N_6430,N_5269,N_5145);
and U6431 (N_6431,N_5571,N_5257);
or U6432 (N_6432,N_5593,N_5171);
nor U6433 (N_6433,N_5857,N_5006);
nor U6434 (N_6434,N_5150,N_5522);
nand U6435 (N_6435,N_5466,N_5251);
nand U6436 (N_6436,N_5619,N_5686);
or U6437 (N_6437,N_5389,N_5021);
or U6438 (N_6438,N_5802,N_5242);
nor U6439 (N_6439,N_5885,N_5570);
xor U6440 (N_6440,N_5874,N_5894);
nand U6441 (N_6441,N_5276,N_5761);
or U6442 (N_6442,N_5966,N_5760);
xnor U6443 (N_6443,N_5817,N_5697);
and U6444 (N_6444,N_5364,N_5722);
and U6445 (N_6445,N_5027,N_5395);
xor U6446 (N_6446,N_5323,N_5374);
nand U6447 (N_6447,N_5487,N_5913);
xor U6448 (N_6448,N_5850,N_5284);
nand U6449 (N_6449,N_5804,N_5101);
and U6450 (N_6450,N_5720,N_5035);
nor U6451 (N_6451,N_5253,N_5709);
or U6452 (N_6452,N_5776,N_5344);
nor U6453 (N_6453,N_5602,N_5981);
or U6454 (N_6454,N_5684,N_5397);
and U6455 (N_6455,N_5782,N_5529);
xnor U6456 (N_6456,N_5084,N_5349);
nor U6457 (N_6457,N_5603,N_5255);
xor U6458 (N_6458,N_5227,N_5503);
xor U6459 (N_6459,N_5353,N_5946);
nand U6460 (N_6460,N_5974,N_5288);
nor U6461 (N_6461,N_5091,N_5339);
nor U6462 (N_6462,N_5634,N_5054);
and U6463 (N_6463,N_5524,N_5944);
or U6464 (N_6464,N_5179,N_5887);
or U6465 (N_6465,N_5102,N_5693);
nor U6466 (N_6466,N_5707,N_5354);
or U6467 (N_6467,N_5396,N_5497);
xor U6468 (N_6468,N_5230,N_5673);
nor U6469 (N_6469,N_5950,N_5350);
and U6470 (N_6470,N_5549,N_5812);
or U6471 (N_6471,N_5873,N_5606);
nand U6472 (N_6472,N_5627,N_5023);
or U6473 (N_6473,N_5993,N_5332);
nor U6474 (N_6474,N_5542,N_5713);
or U6475 (N_6475,N_5667,N_5719);
or U6476 (N_6476,N_5224,N_5425);
and U6477 (N_6477,N_5083,N_5189);
or U6478 (N_6478,N_5754,N_5835);
nor U6479 (N_6479,N_5370,N_5426);
nand U6480 (N_6480,N_5365,N_5477);
nand U6481 (N_6481,N_5589,N_5514);
and U6482 (N_6482,N_5127,N_5181);
or U6483 (N_6483,N_5938,N_5826);
nor U6484 (N_6484,N_5863,N_5509);
and U6485 (N_6485,N_5014,N_5651);
xor U6486 (N_6486,N_5309,N_5294);
and U6487 (N_6487,N_5172,N_5291);
nand U6488 (N_6488,N_5095,N_5041);
or U6489 (N_6489,N_5699,N_5650);
nor U6490 (N_6490,N_5134,N_5267);
or U6491 (N_6491,N_5262,N_5566);
nor U6492 (N_6492,N_5939,N_5930);
nand U6493 (N_6493,N_5829,N_5480);
or U6494 (N_6494,N_5437,N_5900);
nor U6495 (N_6495,N_5785,N_5001);
or U6496 (N_6496,N_5952,N_5490);
nor U6497 (N_6497,N_5705,N_5133);
and U6498 (N_6498,N_5153,N_5141);
nor U6499 (N_6499,N_5839,N_5991);
or U6500 (N_6500,N_5175,N_5014);
nor U6501 (N_6501,N_5397,N_5295);
or U6502 (N_6502,N_5282,N_5127);
or U6503 (N_6503,N_5041,N_5974);
or U6504 (N_6504,N_5422,N_5959);
and U6505 (N_6505,N_5458,N_5203);
nand U6506 (N_6506,N_5091,N_5469);
and U6507 (N_6507,N_5952,N_5141);
xor U6508 (N_6508,N_5187,N_5383);
and U6509 (N_6509,N_5642,N_5893);
and U6510 (N_6510,N_5353,N_5294);
nand U6511 (N_6511,N_5294,N_5091);
or U6512 (N_6512,N_5021,N_5837);
nand U6513 (N_6513,N_5396,N_5233);
nand U6514 (N_6514,N_5041,N_5259);
and U6515 (N_6515,N_5195,N_5956);
nand U6516 (N_6516,N_5915,N_5973);
or U6517 (N_6517,N_5461,N_5129);
xnor U6518 (N_6518,N_5320,N_5018);
nand U6519 (N_6519,N_5461,N_5786);
nor U6520 (N_6520,N_5378,N_5577);
nor U6521 (N_6521,N_5011,N_5721);
nand U6522 (N_6522,N_5245,N_5331);
nand U6523 (N_6523,N_5337,N_5601);
nand U6524 (N_6524,N_5714,N_5411);
nand U6525 (N_6525,N_5553,N_5454);
or U6526 (N_6526,N_5133,N_5074);
nand U6527 (N_6527,N_5639,N_5070);
xnor U6528 (N_6528,N_5162,N_5054);
nand U6529 (N_6529,N_5854,N_5536);
xnor U6530 (N_6530,N_5189,N_5625);
nor U6531 (N_6531,N_5891,N_5064);
xnor U6532 (N_6532,N_5894,N_5264);
or U6533 (N_6533,N_5987,N_5436);
or U6534 (N_6534,N_5266,N_5610);
nand U6535 (N_6535,N_5447,N_5914);
nand U6536 (N_6536,N_5329,N_5364);
nor U6537 (N_6537,N_5636,N_5483);
or U6538 (N_6538,N_5301,N_5468);
and U6539 (N_6539,N_5725,N_5265);
nor U6540 (N_6540,N_5855,N_5386);
and U6541 (N_6541,N_5389,N_5557);
xor U6542 (N_6542,N_5255,N_5935);
and U6543 (N_6543,N_5944,N_5812);
and U6544 (N_6544,N_5436,N_5905);
and U6545 (N_6545,N_5649,N_5928);
nor U6546 (N_6546,N_5563,N_5614);
xnor U6547 (N_6547,N_5177,N_5470);
nand U6548 (N_6548,N_5705,N_5497);
or U6549 (N_6549,N_5846,N_5673);
and U6550 (N_6550,N_5100,N_5884);
xnor U6551 (N_6551,N_5762,N_5635);
or U6552 (N_6552,N_5954,N_5172);
nor U6553 (N_6553,N_5486,N_5491);
nand U6554 (N_6554,N_5982,N_5126);
or U6555 (N_6555,N_5177,N_5655);
xor U6556 (N_6556,N_5489,N_5701);
xnor U6557 (N_6557,N_5386,N_5259);
nand U6558 (N_6558,N_5310,N_5598);
nor U6559 (N_6559,N_5405,N_5652);
or U6560 (N_6560,N_5517,N_5487);
or U6561 (N_6561,N_5330,N_5727);
xor U6562 (N_6562,N_5845,N_5604);
or U6563 (N_6563,N_5915,N_5009);
xnor U6564 (N_6564,N_5395,N_5938);
and U6565 (N_6565,N_5489,N_5742);
or U6566 (N_6566,N_5718,N_5258);
nand U6567 (N_6567,N_5420,N_5405);
and U6568 (N_6568,N_5531,N_5662);
nand U6569 (N_6569,N_5739,N_5528);
nand U6570 (N_6570,N_5214,N_5448);
nor U6571 (N_6571,N_5330,N_5506);
nor U6572 (N_6572,N_5124,N_5043);
and U6573 (N_6573,N_5072,N_5260);
nor U6574 (N_6574,N_5876,N_5093);
and U6575 (N_6575,N_5135,N_5750);
and U6576 (N_6576,N_5957,N_5418);
and U6577 (N_6577,N_5799,N_5285);
nor U6578 (N_6578,N_5493,N_5205);
or U6579 (N_6579,N_5779,N_5418);
xnor U6580 (N_6580,N_5482,N_5024);
and U6581 (N_6581,N_5924,N_5649);
nor U6582 (N_6582,N_5713,N_5216);
xnor U6583 (N_6583,N_5598,N_5772);
or U6584 (N_6584,N_5709,N_5956);
and U6585 (N_6585,N_5120,N_5624);
or U6586 (N_6586,N_5773,N_5184);
nor U6587 (N_6587,N_5076,N_5513);
and U6588 (N_6588,N_5782,N_5170);
xnor U6589 (N_6589,N_5733,N_5272);
or U6590 (N_6590,N_5174,N_5266);
nor U6591 (N_6591,N_5879,N_5593);
xnor U6592 (N_6592,N_5407,N_5332);
xnor U6593 (N_6593,N_5930,N_5375);
xor U6594 (N_6594,N_5057,N_5095);
nand U6595 (N_6595,N_5599,N_5959);
and U6596 (N_6596,N_5193,N_5137);
xnor U6597 (N_6597,N_5782,N_5862);
nor U6598 (N_6598,N_5958,N_5357);
or U6599 (N_6599,N_5125,N_5993);
and U6600 (N_6600,N_5663,N_5569);
nand U6601 (N_6601,N_5183,N_5840);
nor U6602 (N_6602,N_5614,N_5968);
xor U6603 (N_6603,N_5311,N_5717);
or U6604 (N_6604,N_5168,N_5756);
xnor U6605 (N_6605,N_5967,N_5656);
nor U6606 (N_6606,N_5177,N_5304);
xnor U6607 (N_6607,N_5536,N_5876);
xor U6608 (N_6608,N_5963,N_5532);
and U6609 (N_6609,N_5364,N_5374);
nand U6610 (N_6610,N_5747,N_5317);
and U6611 (N_6611,N_5732,N_5087);
xor U6612 (N_6612,N_5400,N_5456);
nand U6613 (N_6613,N_5100,N_5908);
nor U6614 (N_6614,N_5885,N_5808);
nor U6615 (N_6615,N_5738,N_5202);
and U6616 (N_6616,N_5107,N_5627);
nand U6617 (N_6617,N_5945,N_5417);
nor U6618 (N_6618,N_5829,N_5335);
nor U6619 (N_6619,N_5775,N_5693);
nor U6620 (N_6620,N_5905,N_5528);
nand U6621 (N_6621,N_5526,N_5321);
or U6622 (N_6622,N_5422,N_5057);
xnor U6623 (N_6623,N_5097,N_5008);
or U6624 (N_6624,N_5425,N_5840);
or U6625 (N_6625,N_5629,N_5715);
or U6626 (N_6626,N_5912,N_5628);
and U6627 (N_6627,N_5119,N_5409);
xor U6628 (N_6628,N_5503,N_5027);
nand U6629 (N_6629,N_5652,N_5965);
and U6630 (N_6630,N_5867,N_5459);
and U6631 (N_6631,N_5064,N_5118);
xnor U6632 (N_6632,N_5359,N_5134);
nor U6633 (N_6633,N_5606,N_5727);
xor U6634 (N_6634,N_5436,N_5616);
or U6635 (N_6635,N_5056,N_5594);
nor U6636 (N_6636,N_5488,N_5379);
or U6637 (N_6637,N_5942,N_5568);
or U6638 (N_6638,N_5747,N_5807);
and U6639 (N_6639,N_5203,N_5188);
nand U6640 (N_6640,N_5926,N_5796);
and U6641 (N_6641,N_5705,N_5896);
nor U6642 (N_6642,N_5876,N_5802);
nand U6643 (N_6643,N_5950,N_5515);
or U6644 (N_6644,N_5604,N_5492);
and U6645 (N_6645,N_5511,N_5901);
or U6646 (N_6646,N_5590,N_5598);
nand U6647 (N_6647,N_5484,N_5958);
nand U6648 (N_6648,N_5669,N_5460);
nor U6649 (N_6649,N_5742,N_5928);
xnor U6650 (N_6650,N_5277,N_5589);
nand U6651 (N_6651,N_5837,N_5397);
or U6652 (N_6652,N_5298,N_5986);
nand U6653 (N_6653,N_5686,N_5178);
xor U6654 (N_6654,N_5106,N_5225);
nand U6655 (N_6655,N_5707,N_5990);
nor U6656 (N_6656,N_5693,N_5002);
or U6657 (N_6657,N_5290,N_5740);
or U6658 (N_6658,N_5830,N_5149);
nand U6659 (N_6659,N_5963,N_5833);
or U6660 (N_6660,N_5929,N_5224);
and U6661 (N_6661,N_5352,N_5497);
or U6662 (N_6662,N_5802,N_5020);
and U6663 (N_6663,N_5101,N_5636);
xnor U6664 (N_6664,N_5708,N_5270);
nor U6665 (N_6665,N_5634,N_5840);
nand U6666 (N_6666,N_5316,N_5719);
nor U6667 (N_6667,N_5923,N_5573);
nand U6668 (N_6668,N_5658,N_5625);
xnor U6669 (N_6669,N_5786,N_5243);
nand U6670 (N_6670,N_5146,N_5190);
nand U6671 (N_6671,N_5352,N_5094);
and U6672 (N_6672,N_5882,N_5303);
xnor U6673 (N_6673,N_5397,N_5775);
and U6674 (N_6674,N_5343,N_5216);
nand U6675 (N_6675,N_5976,N_5460);
and U6676 (N_6676,N_5183,N_5835);
xnor U6677 (N_6677,N_5779,N_5083);
nor U6678 (N_6678,N_5795,N_5242);
nand U6679 (N_6679,N_5900,N_5537);
and U6680 (N_6680,N_5384,N_5924);
nor U6681 (N_6681,N_5555,N_5655);
nor U6682 (N_6682,N_5284,N_5799);
nor U6683 (N_6683,N_5768,N_5710);
nand U6684 (N_6684,N_5739,N_5362);
or U6685 (N_6685,N_5146,N_5552);
xnor U6686 (N_6686,N_5666,N_5427);
or U6687 (N_6687,N_5822,N_5441);
nor U6688 (N_6688,N_5579,N_5094);
or U6689 (N_6689,N_5187,N_5304);
nor U6690 (N_6690,N_5696,N_5829);
nor U6691 (N_6691,N_5293,N_5295);
xnor U6692 (N_6692,N_5122,N_5036);
nor U6693 (N_6693,N_5206,N_5795);
xnor U6694 (N_6694,N_5063,N_5920);
xnor U6695 (N_6695,N_5243,N_5909);
nand U6696 (N_6696,N_5974,N_5218);
xor U6697 (N_6697,N_5309,N_5270);
nand U6698 (N_6698,N_5976,N_5979);
or U6699 (N_6699,N_5707,N_5893);
or U6700 (N_6700,N_5176,N_5792);
nand U6701 (N_6701,N_5200,N_5474);
nand U6702 (N_6702,N_5617,N_5304);
nand U6703 (N_6703,N_5588,N_5679);
and U6704 (N_6704,N_5746,N_5673);
or U6705 (N_6705,N_5422,N_5564);
or U6706 (N_6706,N_5652,N_5859);
or U6707 (N_6707,N_5856,N_5051);
nand U6708 (N_6708,N_5596,N_5784);
or U6709 (N_6709,N_5454,N_5456);
nor U6710 (N_6710,N_5619,N_5413);
or U6711 (N_6711,N_5372,N_5927);
nand U6712 (N_6712,N_5468,N_5088);
or U6713 (N_6713,N_5958,N_5310);
and U6714 (N_6714,N_5646,N_5230);
and U6715 (N_6715,N_5512,N_5556);
or U6716 (N_6716,N_5668,N_5392);
and U6717 (N_6717,N_5095,N_5725);
or U6718 (N_6718,N_5610,N_5660);
and U6719 (N_6719,N_5739,N_5843);
or U6720 (N_6720,N_5431,N_5117);
xnor U6721 (N_6721,N_5135,N_5390);
nor U6722 (N_6722,N_5921,N_5228);
xnor U6723 (N_6723,N_5497,N_5032);
nor U6724 (N_6724,N_5254,N_5889);
xor U6725 (N_6725,N_5616,N_5700);
nor U6726 (N_6726,N_5759,N_5412);
xnor U6727 (N_6727,N_5728,N_5341);
nand U6728 (N_6728,N_5403,N_5977);
or U6729 (N_6729,N_5833,N_5742);
and U6730 (N_6730,N_5814,N_5451);
or U6731 (N_6731,N_5505,N_5103);
or U6732 (N_6732,N_5937,N_5763);
nor U6733 (N_6733,N_5939,N_5026);
and U6734 (N_6734,N_5535,N_5635);
nor U6735 (N_6735,N_5803,N_5714);
nand U6736 (N_6736,N_5177,N_5130);
xor U6737 (N_6737,N_5963,N_5490);
and U6738 (N_6738,N_5913,N_5404);
xnor U6739 (N_6739,N_5562,N_5497);
xor U6740 (N_6740,N_5202,N_5204);
xnor U6741 (N_6741,N_5899,N_5481);
or U6742 (N_6742,N_5424,N_5514);
nor U6743 (N_6743,N_5222,N_5486);
nor U6744 (N_6744,N_5672,N_5479);
or U6745 (N_6745,N_5407,N_5996);
or U6746 (N_6746,N_5333,N_5353);
xor U6747 (N_6747,N_5190,N_5045);
or U6748 (N_6748,N_5469,N_5462);
xor U6749 (N_6749,N_5735,N_5733);
and U6750 (N_6750,N_5904,N_5666);
or U6751 (N_6751,N_5539,N_5099);
or U6752 (N_6752,N_5899,N_5111);
and U6753 (N_6753,N_5783,N_5664);
xnor U6754 (N_6754,N_5133,N_5109);
nand U6755 (N_6755,N_5210,N_5902);
nand U6756 (N_6756,N_5600,N_5819);
or U6757 (N_6757,N_5427,N_5875);
nor U6758 (N_6758,N_5466,N_5960);
and U6759 (N_6759,N_5568,N_5369);
and U6760 (N_6760,N_5474,N_5138);
nand U6761 (N_6761,N_5290,N_5089);
nor U6762 (N_6762,N_5605,N_5319);
or U6763 (N_6763,N_5155,N_5295);
and U6764 (N_6764,N_5520,N_5181);
xor U6765 (N_6765,N_5143,N_5934);
and U6766 (N_6766,N_5169,N_5383);
or U6767 (N_6767,N_5551,N_5336);
nor U6768 (N_6768,N_5379,N_5247);
xor U6769 (N_6769,N_5279,N_5551);
nor U6770 (N_6770,N_5445,N_5515);
or U6771 (N_6771,N_5418,N_5226);
nand U6772 (N_6772,N_5206,N_5422);
or U6773 (N_6773,N_5699,N_5074);
or U6774 (N_6774,N_5038,N_5718);
nor U6775 (N_6775,N_5849,N_5800);
nor U6776 (N_6776,N_5566,N_5307);
xor U6777 (N_6777,N_5776,N_5897);
or U6778 (N_6778,N_5144,N_5766);
xor U6779 (N_6779,N_5652,N_5665);
xor U6780 (N_6780,N_5752,N_5511);
or U6781 (N_6781,N_5161,N_5431);
or U6782 (N_6782,N_5572,N_5705);
and U6783 (N_6783,N_5520,N_5215);
or U6784 (N_6784,N_5138,N_5542);
and U6785 (N_6785,N_5236,N_5604);
xnor U6786 (N_6786,N_5700,N_5439);
xor U6787 (N_6787,N_5094,N_5419);
xor U6788 (N_6788,N_5411,N_5761);
and U6789 (N_6789,N_5910,N_5866);
and U6790 (N_6790,N_5540,N_5806);
nor U6791 (N_6791,N_5397,N_5559);
nor U6792 (N_6792,N_5500,N_5292);
xor U6793 (N_6793,N_5166,N_5918);
nand U6794 (N_6794,N_5842,N_5172);
and U6795 (N_6795,N_5767,N_5550);
nor U6796 (N_6796,N_5660,N_5622);
nand U6797 (N_6797,N_5287,N_5505);
xor U6798 (N_6798,N_5202,N_5742);
nand U6799 (N_6799,N_5672,N_5188);
and U6800 (N_6800,N_5854,N_5899);
xnor U6801 (N_6801,N_5767,N_5133);
or U6802 (N_6802,N_5657,N_5121);
and U6803 (N_6803,N_5809,N_5171);
and U6804 (N_6804,N_5617,N_5261);
or U6805 (N_6805,N_5447,N_5731);
nor U6806 (N_6806,N_5233,N_5379);
nand U6807 (N_6807,N_5801,N_5459);
and U6808 (N_6808,N_5852,N_5772);
or U6809 (N_6809,N_5295,N_5139);
nand U6810 (N_6810,N_5252,N_5422);
and U6811 (N_6811,N_5699,N_5492);
and U6812 (N_6812,N_5300,N_5702);
nand U6813 (N_6813,N_5475,N_5292);
or U6814 (N_6814,N_5865,N_5827);
nor U6815 (N_6815,N_5807,N_5982);
nand U6816 (N_6816,N_5968,N_5974);
xor U6817 (N_6817,N_5789,N_5357);
nor U6818 (N_6818,N_5117,N_5514);
and U6819 (N_6819,N_5633,N_5484);
nor U6820 (N_6820,N_5848,N_5859);
or U6821 (N_6821,N_5529,N_5641);
and U6822 (N_6822,N_5566,N_5484);
and U6823 (N_6823,N_5643,N_5825);
or U6824 (N_6824,N_5918,N_5097);
or U6825 (N_6825,N_5677,N_5191);
and U6826 (N_6826,N_5803,N_5089);
nand U6827 (N_6827,N_5192,N_5782);
and U6828 (N_6828,N_5006,N_5288);
nand U6829 (N_6829,N_5570,N_5355);
nor U6830 (N_6830,N_5586,N_5317);
nor U6831 (N_6831,N_5175,N_5869);
nor U6832 (N_6832,N_5615,N_5610);
nor U6833 (N_6833,N_5778,N_5657);
or U6834 (N_6834,N_5728,N_5639);
nor U6835 (N_6835,N_5018,N_5922);
nand U6836 (N_6836,N_5839,N_5369);
nor U6837 (N_6837,N_5218,N_5964);
and U6838 (N_6838,N_5991,N_5249);
and U6839 (N_6839,N_5581,N_5568);
nand U6840 (N_6840,N_5988,N_5537);
or U6841 (N_6841,N_5889,N_5833);
and U6842 (N_6842,N_5725,N_5411);
nor U6843 (N_6843,N_5962,N_5748);
and U6844 (N_6844,N_5033,N_5032);
nor U6845 (N_6845,N_5916,N_5679);
nor U6846 (N_6846,N_5188,N_5408);
and U6847 (N_6847,N_5461,N_5594);
or U6848 (N_6848,N_5213,N_5758);
nand U6849 (N_6849,N_5703,N_5851);
nor U6850 (N_6850,N_5731,N_5120);
nand U6851 (N_6851,N_5148,N_5922);
nand U6852 (N_6852,N_5483,N_5386);
xnor U6853 (N_6853,N_5825,N_5126);
nor U6854 (N_6854,N_5880,N_5317);
or U6855 (N_6855,N_5877,N_5631);
and U6856 (N_6856,N_5560,N_5557);
xnor U6857 (N_6857,N_5887,N_5894);
xor U6858 (N_6858,N_5816,N_5899);
nor U6859 (N_6859,N_5717,N_5118);
and U6860 (N_6860,N_5252,N_5215);
nor U6861 (N_6861,N_5977,N_5484);
xnor U6862 (N_6862,N_5743,N_5206);
or U6863 (N_6863,N_5447,N_5202);
or U6864 (N_6864,N_5324,N_5031);
and U6865 (N_6865,N_5073,N_5901);
or U6866 (N_6866,N_5059,N_5498);
nand U6867 (N_6867,N_5115,N_5800);
nor U6868 (N_6868,N_5273,N_5696);
and U6869 (N_6869,N_5025,N_5037);
xor U6870 (N_6870,N_5279,N_5957);
nor U6871 (N_6871,N_5906,N_5916);
or U6872 (N_6872,N_5492,N_5952);
nor U6873 (N_6873,N_5284,N_5697);
and U6874 (N_6874,N_5946,N_5974);
or U6875 (N_6875,N_5696,N_5687);
xor U6876 (N_6876,N_5580,N_5170);
or U6877 (N_6877,N_5003,N_5837);
nor U6878 (N_6878,N_5388,N_5093);
xor U6879 (N_6879,N_5945,N_5796);
or U6880 (N_6880,N_5790,N_5245);
and U6881 (N_6881,N_5863,N_5508);
nor U6882 (N_6882,N_5980,N_5254);
nor U6883 (N_6883,N_5204,N_5759);
or U6884 (N_6884,N_5951,N_5873);
xnor U6885 (N_6885,N_5416,N_5530);
xnor U6886 (N_6886,N_5547,N_5960);
nand U6887 (N_6887,N_5525,N_5053);
xnor U6888 (N_6888,N_5388,N_5914);
and U6889 (N_6889,N_5618,N_5731);
nor U6890 (N_6890,N_5896,N_5153);
nor U6891 (N_6891,N_5754,N_5626);
and U6892 (N_6892,N_5057,N_5718);
nand U6893 (N_6893,N_5798,N_5737);
and U6894 (N_6894,N_5356,N_5478);
nor U6895 (N_6895,N_5399,N_5779);
nand U6896 (N_6896,N_5950,N_5078);
nand U6897 (N_6897,N_5584,N_5978);
nor U6898 (N_6898,N_5730,N_5927);
nand U6899 (N_6899,N_5416,N_5524);
and U6900 (N_6900,N_5870,N_5515);
or U6901 (N_6901,N_5454,N_5576);
or U6902 (N_6902,N_5820,N_5806);
nand U6903 (N_6903,N_5574,N_5815);
or U6904 (N_6904,N_5495,N_5974);
and U6905 (N_6905,N_5748,N_5844);
nand U6906 (N_6906,N_5793,N_5970);
nor U6907 (N_6907,N_5698,N_5213);
nor U6908 (N_6908,N_5972,N_5514);
xnor U6909 (N_6909,N_5786,N_5207);
or U6910 (N_6910,N_5585,N_5562);
or U6911 (N_6911,N_5127,N_5791);
or U6912 (N_6912,N_5796,N_5588);
nor U6913 (N_6913,N_5441,N_5707);
and U6914 (N_6914,N_5134,N_5450);
nor U6915 (N_6915,N_5439,N_5359);
or U6916 (N_6916,N_5369,N_5622);
or U6917 (N_6917,N_5085,N_5838);
or U6918 (N_6918,N_5748,N_5269);
or U6919 (N_6919,N_5464,N_5455);
nand U6920 (N_6920,N_5928,N_5975);
nor U6921 (N_6921,N_5594,N_5662);
and U6922 (N_6922,N_5561,N_5362);
or U6923 (N_6923,N_5134,N_5696);
or U6924 (N_6924,N_5034,N_5473);
nand U6925 (N_6925,N_5977,N_5701);
nor U6926 (N_6926,N_5956,N_5575);
and U6927 (N_6927,N_5802,N_5640);
or U6928 (N_6928,N_5015,N_5214);
nand U6929 (N_6929,N_5161,N_5988);
and U6930 (N_6930,N_5804,N_5828);
xnor U6931 (N_6931,N_5148,N_5565);
and U6932 (N_6932,N_5885,N_5838);
xnor U6933 (N_6933,N_5934,N_5635);
or U6934 (N_6934,N_5103,N_5288);
or U6935 (N_6935,N_5385,N_5149);
xnor U6936 (N_6936,N_5612,N_5134);
and U6937 (N_6937,N_5269,N_5410);
nor U6938 (N_6938,N_5342,N_5775);
or U6939 (N_6939,N_5282,N_5573);
xor U6940 (N_6940,N_5549,N_5613);
nor U6941 (N_6941,N_5016,N_5351);
nor U6942 (N_6942,N_5454,N_5106);
xnor U6943 (N_6943,N_5063,N_5917);
nand U6944 (N_6944,N_5210,N_5367);
nand U6945 (N_6945,N_5645,N_5800);
nor U6946 (N_6946,N_5244,N_5229);
nand U6947 (N_6947,N_5877,N_5299);
and U6948 (N_6948,N_5049,N_5805);
nor U6949 (N_6949,N_5937,N_5524);
nand U6950 (N_6950,N_5739,N_5232);
xor U6951 (N_6951,N_5659,N_5262);
or U6952 (N_6952,N_5806,N_5158);
nand U6953 (N_6953,N_5196,N_5216);
and U6954 (N_6954,N_5077,N_5568);
xnor U6955 (N_6955,N_5941,N_5404);
xnor U6956 (N_6956,N_5532,N_5172);
and U6957 (N_6957,N_5874,N_5609);
nor U6958 (N_6958,N_5583,N_5742);
xnor U6959 (N_6959,N_5786,N_5298);
nor U6960 (N_6960,N_5288,N_5852);
nand U6961 (N_6961,N_5100,N_5811);
and U6962 (N_6962,N_5421,N_5179);
nand U6963 (N_6963,N_5377,N_5549);
xnor U6964 (N_6964,N_5746,N_5378);
and U6965 (N_6965,N_5212,N_5540);
or U6966 (N_6966,N_5539,N_5939);
nand U6967 (N_6967,N_5741,N_5272);
or U6968 (N_6968,N_5139,N_5718);
xnor U6969 (N_6969,N_5548,N_5815);
nand U6970 (N_6970,N_5498,N_5486);
or U6971 (N_6971,N_5139,N_5076);
nor U6972 (N_6972,N_5329,N_5971);
nor U6973 (N_6973,N_5033,N_5471);
nor U6974 (N_6974,N_5213,N_5260);
xor U6975 (N_6975,N_5780,N_5216);
nor U6976 (N_6976,N_5986,N_5647);
xor U6977 (N_6977,N_5656,N_5579);
nor U6978 (N_6978,N_5755,N_5471);
xnor U6979 (N_6979,N_5943,N_5050);
nor U6980 (N_6980,N_5940,N_5599);
and U6981 (N_6981,N_5251,N_5328);
nand U6982 (N_6982,N_5742,N_5562);
nand U6983 (N_6983,N_5084,N_5103);
or U6984 (N_6984,N_5121,N_5252);
or U6985 (N_6985,N_5525,N_5501);
or U6986 (N_6986,N_5985,N_5296);
xor U6987 (N_6987,N_5046,N_5949);
or U6988 (N_6988,N_5180,N_5727);
xor U6989 (N_6989,N_5800,N_5586);
xnor U6990 (N_6990,N_5020,N_5284);
nor U6991 (N_6991,N_5386,N_5459);
xnor U6992 (N_6992,N_5856,N_5741);
or U6993 (N_6993,N_5798,N_5120);
nor U6994 (N_6994,N_5650,N_5884);
and U6995 (N_6995,N_5208,N_5270);
nor U6996 (N_6996,N_5762,N_5207);
and U6997 (N_6997,N_5748,N_5394);
nor U6998 (N_6998,N_5361,N_5759);
or U6999 (N_6999,N_5838,N_5080);
xnor U7000 (N_7000,N_6149,N_6144);
and U7001 (N_7001,N_6557,N_6194);
nand U7002 (N_7002,N_6212,N_6406);
xor U7003 (N_7003,N_6056,N_6115);
nor U7004 (N_7004,N_6847,N_6333);
xnor U7005 (N_7005,N_6186,N_6733);
nand U7006 (N_7006,N_6527,N_6600);
nor U7007 (N_7007,N_6199,N_6261);
and U7008 (N_7008,N_6266,N_6647);
nor U7009 (N_7009,N_6592,N_6454);
nor U7010 (N_7010,N_6417,N_6483);
and U7011 (N_7011,N_6955,N_6951);
xor U7012 (N_7012,N_6973,N_6168);
or U7013 (N_7013,N_6792,N_6879);
nor U7014 (N_7014,N_6257,N_6931);
xor U7015 (N_7015,N_6443,N_6609);
xnor U7016 (N_7016,N_6669,N_6095);
or U7017 (N_7017,N_6552,N_6368);
nand U7018 (N_7018,N_6660,N_6240);
nand U7019 (N_7019,N_6601,N_6227);
and U7020 (N_7020,N_6356,N_6793);
or U7021 (N_7021,N_6743,N_6263);
or U7022 (N_7022,N_6907,N_6626);
or U7023 (N_7023,N_6890,N_6964);
nor U7024 (N_7024,N_6332,N_6902);
nor U7025 (N_7025,N_6587,N_6362);
nand U7026 (N_7026,N_6710,N_6039);
and U7027 (N_7027,N_6739,N_6585);
and U7028 (N_7028,N_6838,N_6146);
and U7029 (N_7029,N_6046,N_6352);
nor U7030 (N_7030,N_6289,N_6512);
and U7031 (N_7031,N_6595,N_6041);
and U7032 (N_7032,N_6258,N_6155);
nand U7033 (N_7033,N_6496,N_6657);
or U7034 (N_7034,N_6022,N_6843);
nand U7035 (N_7035,N_6249,N_6223);
nand U7036 (N_7036,N_6325,N_6250);
nor U7037 (N_7037,N_6556,N_6510);
and U7038 (N_7038,N_6016,N_6132);
nor U7039 (N_7039,N_6324,N_6775);
or U7040 (N_7040,N_6081,N_6184);
xnor U7041 (N_7041,N_6282,N_6499);
xnor U7042 (N_7042,N_6900,N_6012);
or U7043 (N_7043,N_6028,N_6208);
xor U7044 (N_7044,N_6667,N_6230);
or U7045 (N_7045,N_6845,N_6596);
nor U7046 (N_7046,N_6681,N_6017);
nor U7047 (N_7047,N_6069,N_6063);
nor U7048 (N_7048,N_6606,N_6237);
nor U7049 (N_7049,N_6941,N_6372);
nor U7050 (N_7050,N_6757,N_6914);
nand U7051 (N_7051,N_6815,N_6287);
nor U7052 (N_7052,N_6448,N_6942);
xnor U7053 (N_7053,N_6807,N_6059);
nand U7054 (N_7054,N_6755,N_6937);
or U7055 (N_7055,N_6108,N_6383);
xnor U7056 (N_7056,N_6818,N_6415);
nand U7057 (N_7057,N_6154,N_6272);
nand U7058 (N_7058,N_6997,N_6286);
xor U7059 (N_7059,N_6814,N_6192);
nand U7060 (N_7060,N_6005,N_6961);
nand U7061 (N_7061,N_6304,N_6607);
nand U7062 (N_7062,N_6539,N_6173);
xor U7063 (N_7063,N_6099,N_6713);
or U7064 (N_7064,N_6288,N_6989);
and U7065 (N_7065,N_6088,N_6629);
or U7066 (N_7066,N_6447,N_6414);
xor U7067 (N_7067,N_6096,N_6954);
or U7068 (N_7068,N_6746,N_6070);
nand U7069 (N_7069,N_6598,N_6238);
or U7070 (N_7070,N_6917,N_6980);
nor U7071 (N_7071,N_6072,N_6891);
or U7072 (N_7072,N_6759,N_6178);
or U7073 (N_7073,N_6611,N_6283);
and U7074 (N_7074,N_6767,N_6800);
nand U7075 (N_7075,N_6180,N_6541);
or U7076 (N_7076,N_6200,N_6861);
and U7077 (N_7077,N_6153,N_6094);
nand U7078 (N_7078,N_6066,N_6213);
nor U7079 (N_7079,N_6472,N_6720);
xnor U7080 (N_7080,N_6080,N_6579);
nor U7081 (N_7081,N_6299,N_6399);
nand U7082 (N_7082,N_6277,N_6489);
nor U7083 (N_7083,N_6544,N_6328);
and U7084 (N_7084,N_6365,N_6018);
and U7085 (N_7085,N_6816,N_6124);
xor U7086 (N_7086,N_6032,N_6130);
xnor U7087 (N_7087,N_6337,N_6811);
or U7088 (N_7088,N_6623,N_6741);
nand U7089 (N_7089,N_6307,N_6226);
or U7090 (N_7090,N_6174,N_6978);
and U7091 (N_7091,N_6666,N_6225);
xnor U7092 (N_7092,N_6523,N_6463);
xnor U7093 (N_7093,N_6247,N_6382);
xor U7094 (N_7094,N_6116,N_6806);
nor U7095 (N_7095,N_6262,N_6561);
or U7096 (N_7096,N_6458,N_6380);
xnor U7097 (N_7097,N_6576,N_6311);
or U7098 (N_7098,N_6122,N_6885);
xnor U7099 (N_7099,N_6172,N_6461);
nand U7100 (N_7100,N_6419,N_6948);
nand U7101 (N_7101,N_6634,N_6752);
or U7102 (N_7102,N_6594,N_6664);
or U7103 (N_7103,N_6179,N_6668);
or U7104 (N_7104,N_6404,N_6197);
or U7105 (N_7105,N_6407,N_6428);
nand U7106 (N_7106,N_6737,N_6047);
xor U7107 (N_7107,N_6930,N_6217);
and U7108 (N_7108,N_6500,N_6825);
or U7109 (N_7109,N_6260,N_6363);
xor U7110 (N_7110,N_6170,N_6791);
nand U7111 (N_7111,N_6052,N_6724);
xnor U7112 (N_7112,N_6011,N_6873);
nand U7113 (N_7113,N_6703,N_6345);
or U7114 (N_7114,N_6850,N_6492);
xor U7115 (N_7115,N_6974,N_6706);
nand U7116 (N_7116,N_6450,N_6677);
or U7117 (N_7117,N_6353,N_6797);
xnor U7118 (N_7118,N_6156,N_6473);
nor U7119 (N_7119,N_6318,N_6529);
nand U7120 (N_7120,N_6698,N_6371);
and U7121 (N_7121,N_6034,N_6769);
or U7122 (N_7122,N_6319,N_6103);
nand U7123 (N_7123,N_6358,N_6469);
and U7124 (N_7124,N_6214,N_6620);
nor U7125 (N_7125,N_6812,N_6418);
nor U7126 (N_7126,N_6008,N_6118);
and U7127 (N_7127,N_6366,N_6152);
or U7128 (N_7128,N_6785,N_6763);
or U7129 (N_7129,N_6140,N_6905);
nand U7130 (N_7130,N_6295,N_6922);
and U7131 (N_7131,N_6548,N_6782);
and U7132 (N_7132,N_6568,N_6903);
nor U7133 (N_7133,N_6136,N_6462);
nand U7134 (N_7134,N_6264,N_6756);
xor U7135 (N_7135,N_6738,N_6646);
or U7136 (N_7136,N_6564,N_6187);
nand U7137 (N_7137,N_6679,N_6639);
nand U7138 (N_7138,N_6497,N_6910);
nor U7139 (N_7139,N_6452,N_6312);
nand U7140 (N_7140,N_6166,N_6532);
xnor U7141 (N_7141,N_6700,N_6425);
nand U7142 (N_7142,N_6235,N_6615);
or U7143 (N_7143,N_6965,N_6940);
nor U7144 (N_7144,N_6894,N_6293);
nand U7145 (N_7145,N_6520,N_6621);
nor U7146 (N_7146,N_6384,N_6993);
nor U7147 (N_7147,N_6430,N_6608);
or U7148 (N_7148,N_6723,N_6549);
xor U7149 (N_7149,N_6685,N_6374);
or U7150 (N_7150,N_6364,N_6882);
and U7151 (N_7151,N_6019,N_6939);
and U7152 (N_7152,N_6431,N_6836);
and U7153 (N_7153,N_6360,N_6962);
nand U7154 (N_7154,N_6165,N_6866);
and U7155 (N_7155,N_6765,N_6521);
nor U7156 (N_7156,N_6886,N_6751);
xor U7157 (N_7157,N_6986,N_6129);
nand U7158 (N_7158,N_6928,N_6898);
nand U7159 (N_7159,N_6842,N_6758);
nor U7160 (N_7160,N_6109,N_6901);
and U7161 (N_7161,N_6602,N_6423);
nor U7162 (N_7162,N_6061,N_6160);
nand U7163 (N_7163,N_6342,N_6958);
and U7164 (N_7164,N_6291,N_6856);
or U7165 (N_7165,N_6844,N_6762);
nand U7166 (N_7166,N_6622,N_6542);
nand U7167 (N_7167,N_6717,N_6983);
nand U7168 (N_7168,N_6446,N_6031);
nor U7169 (N_7169,N_6869,N_6317);
and U7170 (N_7170,N_6068,N_6540);
nand U7171 (N_7171,N_6676,N_6693);
and U7172 (N_7172,N_6935,N_6871);
nand U7173 (N_7173,N_6092,N_6486);
nand U7174 (N_7174,N_6967,N_6895);
nand U7175 (N_7175,N_6916,N_6003);
or U7176 (N_7176,N_6281,N_6709);
nor U7177 (N_7177,N_6728,N_6078);
xor U7178 (N_7178,N_6329,N_6605);
nor U7179 (N_7179,N_6987,N_6426);
or U7180 (N_7180,N_6137,N_6773);
and U7181 (N_7181,N_6141,N_6531);
xnor U7182 (N_7182,N_6488,N_6390);
or U7183 (N_7183,N_6270,N_6347);
nand U7184 (N_7184,N_6829,N_6221);
or U7185 (N_7185,N_6672,N_6401);
xor U7186 (N_7186,N_6701,N_6887);
and U7187 (N_7187,N_6188,N_6934);
nor U7188 (N_7188,N_6010,N_6563);
xor U7189 (N_7189,N_6004,N_6956);
or U7190 (N_7190,N_6259,N_6025);
nand U7191 (N_7191,N_6851,N_6645);
nand U7192 (N_7192,N_6480,N_6210);
nand U7193 (N_7193,N_6267,N_6754);
nand U7194 (N_7194,N_6794,N_6968);
nor U7195 (N_7195,N_6175,N_6550);
nand U7196 (N_7196,N_6193,N_6766);
and U7197 (N_7197,N_6176,N_6897);
xnor U7198 (N_7198,N_6920,N_6904);
nand U7199 (N_7199,N_6359,N_6429);
nand U7200 (N_7200,N_6157,N_6921);
or U7201 (N_7201,N_6860,N_6490);
or U7202 (N_7202,N_6553,N_6727);
or U7203 (N_7203,N_6239,N_6831);
xor U7204 (N_7204,N_6373,N_6933);
or U7205 (N_7205,N_6035,N_6632);
and U7206 (N_7206,N_6091,N_6945);
xnor U7207 (N_7207,N_6841,N_6551);
nor U7208 (N_7208,N_6637,N_6938);
or U7209 (N_7209,N_6231,N_6734);
and U7210 (N_7210,N_6460,N_6798);
nand U7211 (N_7211,N_6705,N_6134);
nor U7212 (N_7212,N_6453,N_6673);
or U7213 (N_7213,N_6086,N_6519);
xnor U7214 (N_7214,N_6659,N_6749);
nor U7215 (N_7215,N_6114,N_6718);
or U7216 (N_7216,N_6327,N_6315);
nand U7217 (N_7217,N_6219,N_6688);
or U7218 (N_7218,N_6670,N_6991);
nand U7219 (N_7219,N_6889,N_6641);
nor U7220 (N_7220,N_6278,N_6138);
xor U7221 (N_7221,N_6880,N_6222);
xnor U7222 (N_7222,N_6369,N_6305);
nand U7223 (N_7223,N_6308,N_6100);
nand U7224 (N_7224,N_6397,N_6216);
and U7225 (N_7225,N_6105,N_6925);
and U7226 (N_7226,N_6236,N_6878);
xor U7227 (N_7227,N_6378,N_6135);
xor U7228 (N_7228,N_6950,N_6121);
or U7229 (N_7229,N_6946,N_6344);
or U7230 (N_7230,N_6823,N_6899);
or U7231 (N_7231,N_6159,N_6248);
nand U7232 (N_7232,N_6392,N_6120);
xor U7233 (N_7233,N_6171,N_6779);
nand U7234 (N_7234,N_6582,N_6470);
nand U7235 (N_7235,N_6143,N_6674);
and U7236 (N_7236,N_6631,N_6457);
or U7237 (N_7237,N_6442,N_6830);
xnor U7238 (N_7238,N_6725,N_6977);
xnor U7239 (N_7239,N_6719,N_6142);
or U7240 (N_7240,N_6926,N_6953);
nor U7241 (N_7241,N_6348,N_6630);
or U7242 (N_7242,N_6777,N_6648);
or U7243 (N_7243,N_6218,N_6000);
nor U7244 (N_7244,N_6837,N_6433);
xor U7245 (N_7245,N_6876,N_6888);
or U7246 (N_7246,N_6826,N_6655);
or U7247 (N_7247,N_6689,N_6432);
xor U7248 (N_7248,N_6870,N_6255);
nand U7249 (N_7249,N_6854,N_6535);
nand U7250 (N_7250,N_6616,N_6273);
nor U7251 (N_7251,N_6245,N_6824);
nor U7252 (N_7252,N_6808,N_6229);
nor U7253 (N_7253,N_6776,N_6436);
xnor U7254 (N_7254,N_6501,N_6191);
nor U7255 (N_7255,N_6906,N_6821);
and U7256 (N_7256,N_6996,N_6456);
nand U7257 (N_7257,N_6139,N_6195);
and U7258 (N_7258,N_6618,N_6874);
xor U7259 (N_7259,N_6150,N_6745);
nor U7260 (N_7260,N_6909,N_6786);
nor U7261 (N_7261,N_6297,N_6377);
xor U7262 (N_7262,N_6482,N_6799);
xor U7263 (N_7263,N_6735,N_6361);
nand U7264 (N_7264,N_6686,N_6809);
xor U7265 (N_7265,N_6466,N_6098);
xor U7266 (N_7266,N_6403,N_6044);
xor U7267 (N_7267,N_6336,N_6636);
and U7268 (N_7268,N_6196,N_6864);
xor U7269 (N_7269,N_6451,N_6590);
nand U7270 (N_7270,N_6638,N_6203);
xnor U7271 (N_7271,N_6960,N_6051);
xnor U7272 (N_7272,N_6065,N_6424);
and U7273 (N_7273,N_6538,N_6554);
and U7274 (N_7274,N_6164,N_6511);
or U7275 (N_7275,N_6543,N_6546);
or U7276 (N_7276,N_6127,N_6694);
nor U7277 (N_7277,N_6682,N_6613);
nor U7278 (N_7278,N_6834,N_6084);
and U7279 (N_7279,N_6349,N_6148);
xnor U7280 (N_7280,N_6370,N_6729);
or U7281 (N_7281,N_6002,N_6848);
xor U7282 (N_7282,N_6079,N_6445);
nor U7283 (N_7283,N_6449,N_6015);
and U7284 (N_7284,N_6586,N_6479);
and U7285 (N_7285,N_6665,N_6274);
and U7286 (N_7286,N_6768,N_6995);
or U7287 (N_7287,N_6627,N_6678);
xnor U7288 (N_7288,N_6998,N_6692);
nand U7289 (N_7289,N_6650,N_6514);
or U7290 (N_7290,N_6947,N_6232);
xor U7291 (N_7291,N_6201,N_6220);
and U7292 (N_7292,N_6093,N_6721);
nand U7293 (N_7293,N_6772,N_6865);
or U7294 (N_7294,N_6427,N_6589);
or U7295 (N_7295,N_6253,N_6963);
and U7296 (N_7296,N_6764,N_6014);
nor U7297 (N_7297,N_6969,N_6316);
xnor U7298 (N_7298,N_6562,N_6813);
nor U7299 (N_7299,N_6509,N_6064);
nand U7300 (N_7300,N_6254,N_6420);
nor U7301 (N_7301,N_6009,N_6675);
and U7302 (N_7302,N_6057,N_6984);
nor U7303 (N_7303,N_6832,N_6400);
xor U7304 (N_7304,N_6732,N_6872);
and U7305 (N_7305,N_6023,N_6007);
xnor U7306 (N_7306,N_6224,N_6972);
nand U7307 (N_7307,N_6029,N_6441);
or U7308 (N_7308,N_6133,N_6073);
or U7309 (N_7309,N_6715,N_6204);
nand U7310 (N_7310,N_6413,N_6128);
and U7311 (N_7311,N_6558,N_6858);
and U7312 (N_7312,N_6584,N_6952);
or U7313 (N_7313,N_6102,N_6614);
nand U7314 (N_7314,N_6908,N_6284);
and U7315 (N_7315,N_6687,N_6591);
nor U7316 (N_7316,N_6911,N_6280);
and U7317 (N_7317,N_6388,N_6367);
nand U7318 (N_7318,N_6524,N_6714);
nand U7319 (N_7319,N_6747,N_6487);
xnor U7320 (N_7320,N_6742,N_6045);
xor U7321 (N_7321,N_6256,N_6990);
nor U7322 (N_7322,N_6503,N_6038);
xnor U7323 (N_7323,N_6409,N_6985);
xnor U7324 (N_7324,N_6533,N_6516);
nor U7325 (N_7325,N_6913,N_6748);
or U7326 (N_7326,N_6040,N_6313);
nand U7327 (N_7327,N_6508,N_6321);
and U7328 (N_7328,N_6435,N_6619);
nor U7329 (N_7329,N_6411,N_6583);
xor U7330 (N_7330,N_6444,N_6357);
nor U7331 (N_7331,N_6774,N_6919);
nand U7332 (N_7332,N_6241,N_6033);
xnor U7333 (N_7333,N_6296,N_6859);
xnor U7334 (N_7334,N_6465,N_6566);
xor U7335 (N_7335,N_6567,N_6625);
xnor U7336 (N_7336,N_6690,N_6402);
nor U7337 (N_7337,N_6581,N_6269);
and U7338 (N_7338,N_6234,N_6205);
nand U7339 (N_7339,N_6736,N_6744);
nor U7340 (N_7340,N_6599,N_6405);
xnor U7341 (N_7341,N_6923,N_6320);
nand U7342 (N_7342,N_6537,N_6107);
nand U7343 (N_7343,N_6617,N_6300);
nand U7344 (N_7344,N_6464,N_6635);
nor U7345 (N_7345,N_6053,N_6309);
nor U7346 (N_7346,N_6013,N_6338);
and U7347 (N_7347,N_6074,N_6001);
or U7348 (N_7348,N_6699,N_6498);
or U7349 (N_7349,N_6857,N_6588);
nand U7350 (N_7350,N_6408,N_6351);
and U7351 (N_7351,N_6438,N_6265);
xnor U7352 (N_7352,N_6478,N_6206);
nand U7353 (N_7353,N_6055,N_6957);
and U7354 (N_7354,N_6396,N_6242);
nand U7355 (N_7355,N_6545,N_6927);
or U7356 (N_7356,N_6375,N_6485);
nand U7357 (N_7357,N_6787,N_6030);
or U7358 (N_7358,N_6228,N_6580);
nor U7359 (N_7359,N_6912,N_6043);
nor U7360 (N_7360,N_6680,N_6802);
or U7361 (N_7361,N_6702,N_6350);
nor U7362 (N_7362,N_6663,N_6471);
xor U7363 (N_7363,N_6387,N_6119);
xor U7364 (N_7364,N_6711,N_6391);
nor U7365 (N_7365,N_6112,N_6167);
nor U7366 (N_7366,N_6083,N_6513);
nor U7367 (N_7367,N_6726,N_6573);
and U7368 (N_7368,N_6493,N_6612);
xor U7369 (N_7369,N_6355,N_6569);
nand U7370 (N_7370,N_6817,N_6306);
and U7371 (N_7371,N_6393,N_6707);
or U7372 (N_7372,N_6394,N_6656);
xnor U7373 (N_7373,N_6944,N_6555);
xor U7374 (N_7374,N_6788,N_6572);
and U7375 (N_7375,N_6323,N_6243);
xor U7376 (N_7376,N_6185,N_6181);
nand U7377 (N_7377,N_6839,N_6559);
xnor U7378 (N_7378,N_6949,N_6202);
or U7379 (N_7379,N_6932,N_6302);
xor U7380 (N_7380,N_6671,N_6077);
nor U7381 (N_7381,N_6994,N_6976);
xnor U7382 (N_7382,N_6021,N_6893);
nand U7383 (N_7383,N_6593,N_6868);
and U7384 (N_7384,N_6104,N_6416);
nand U7385 (N_7385,N_6803,N_6849);
nand U7386 (N_7386,N_6691,N_6145);
nor U7387 (N_7387,N_6036,N_6294);
nor U7388 (N_7388,N_6644,N_6658);
xor U7389 (N_7389,N_6026,N_6640);
and U7390 (N_7390,N_6090,N_6918);
nor U7391 (N_7391,N_6504,N_6507);
or U7392 (N_7392,N_6314,N_6796);
xor U7393 (N_7393,N_6125,N_6481);
nor U7394 (N_7394,N_6840,N_6207);
and U7395 (N_7395,N_6131,N_6805);
or U7396 (N_7396,N_6440,N_6177);
xor U7397 (N_7397,N_6684,N_6783);
xor U7398 (N_7398,N_6704,N_6183);
nand U7399 (N_7399,N_6604,N_6476);
nand U7400 (N_7400,N_6525,N_6975);
nor U7401 (N_7401,N_6505,N_6082);
and U7402 (N_7402,N_6731,N_6067);
or U7403 (N_7403,N_6292,N_6271);
or U7404 (N_7404,N_6395,N_6827);
xnor U7405 (N_7405,N_6780,N_6042);
xor U7406 (N_7406,N_6058,N_6389);
nor U7407 (N_7407,N_6712,N_6169);
and U7408 (N_7408,N_6049,N_6771);
nand U7409 (N_7409,N_6422,N_6722);
nand U7410 (N_7410,N_6828,N_6804);
or U7411 (N_7411,N_6892,N_6867);
xnor U7412 (N_7412,N_6233,N_6182);
nor U7413 (N_7413,N_6575,N_6740);
nand U7414 (N_7414,N_6346,N_6881);
or U7415 (N_7415,N_6101,N_6877);
nor U7416 (N_7416,N_6494,N_6477);
or U7417 (N_7417,N_6896,N_6298);
nand U7418 (N_7418,N_6190,N_6822);
nor U7419 (N_7419,N_6381,N_6060);
or U7420 (N_7420,N_6603,N_6385);
nand U7421 (N_7421,N_6853,N_6578);
or U7422 (N_7422,N_6695,N_6833);
and U7423 (N_7423,N_6502,N_6966);
nor U7424 (N_7424,N_6111,N_6971);
and U7425 (N_7425,N_6117,N_6534);
and U7426 (N_7426,N_6379,N_6113);
xnor U7427 (N_7427,N_6484,N_6303);
nand U7428 (N_7428,N_6276,N_6943);
and U7429 (N_7429,N_6339,N_6158);
nand U7430 (N_7430,N_6642,N_6760);
nand U7431 (N_7431,N_6696,N_6784);
xor U7432 (N_7432,N_6341,N_6439);
nand U7433 (N_7433,N_6565,N_6126);
nor U7434 (N_7434,N_6970,N_6123);
xor U7435 (N_7435,N_6790,N_6301);
or U7436 (N_7436,N_6097,N_6819);
nor U7437 (N_7437,N_6560,N_6628);
nor U7438 (N_7438,N_6246,N_6795);
nor U7439 (N_7439,N_6597,N_6801);
xor U7440 (N_7440,N_6506,N_6653);
xnor U7441 (N_7441,N_6434,N_6037);
nor U7442 (N_7442,N_6661,N_6981);
or U7443 (N_7443,N_6863,N_6855);
xnor U7444 (N_7444,N_6526,N_6062);
nor U7445 (N_7445,N_6340,N_6761);
and U7446 (N_7446,N_6884,N_6770);
nand U7447 (N_7447,N_6020,N_6110);
and U7448 (N_7448,N_6810,N_6334);
xnor U7449 (N_7449,N_6050,N_6085);
xor U7450 (N_7450,N_6468,N_6982);
xor U7451 (N_7451,N_6354,N_6883);
or U7452 (N_7452,N_6054,N_6147);
or U7453 (N_7453,N_6310,N_6515);
and U7454 (N_7454,N_6209,N_6571);
and U7455 (N_7455,N_6753,N_6275);
xnor U7456 (N_7456,N_6643,N_6024);
and U7457 (N_7457,N_6279,N_6536);
or U7458 (N_7458,N_6215,N_6376);
nand U7459 (N_7459,N_6189,N_6087);
nor U7460 (N_7460,N_6862,N_6386);
and U7461 (N_7461,N_6654,N_6789);
xnor U7462 (N_7462,N_6517,N_6089);
or U7463 (N_7463,N_6852,N_6161);
nand U7464 (N_7464,N_6716,N_6198);
nand U7465 (N_7465,N_6915,N_6652);
or U7466 (N_7466,N_6491,N_6467);
nand U7467 (N_7467,N_6518,N_6076);
nor U7468 (N_7468,N_6421,N_6330);
and U7469 (N_7469,N_6335,N_6662);
nand U7470 (N_7470,N_6781,N_6528);
xnor U7471 (N_7471,N_6251,N_6027);
and U7472 (N_7472,N_6326,N_6495);
xnor U7473 (N_7473,N_6979,N_6268);
nand U7474 (N_7474,N_6846,N_6162);
nor U7475 (N_7475,N_6455,N_6071);
xnor U7476 (N_7476,N_6530,N_6331);
and U7477 (N_7477,N_6048,N_6708);
xnor U7478 (N_7478,N_6547,N_6290);
nand U7479 (N_7479,N_6522,N_6610);
nor U7480 (N_7480,N_6475,N_6936);
and U7481 (N_7481,N_6343,N_6285);
and U7482 (N_7482,N_6577,N_6999);
xnor U7483 (N_7483,N_6992,N_6633);
and U7484 (N_7484,N_6211,N_6835);
xnor U7485 (N_7485,N_6252,N_6624);
nor U7486 (N_7486,N_6006,N_6778);
xnor U7487 (N_7487,N_6683,N_6244);
and U7488 (N_7488,N_6163,N_6437);
xor U7489 (N_7489,N_6474,N_6075);
and U7490 (N_7490,N_6649,N_6651);
nor U7491 (N_7491,N_6875,N_6929);
or U7492 (N_7492,N_6574,N_6322);
nand U7493 (N_7493,N_6750,N_6924);
and U7494 (N_7494,N_6697,N_6988);
and U7495 (N_7495,N_6106,N_6459);
xnor U7496 (N_7496,N_6398,N_6570);
xnor U7497 (N_7497,N_6410,N_6412);
or U7498 (N_7498,N_6959,N_6730);
and U7499 (N_7499,N_6151,N_6820);
nor U7500 (N_7500,N_6511,N_6583);
xnor U7501 (N_7501,N_6729,N_6408);
xor U7502 (N_7502,N_6987,N_6435);
nand U7503 (N_7503,N_6895,N_6073);
nor U7504 (N_7504,N_6186,N_6330);
xor U7505 (N_7505,N_6628,N_6936);
nor U7506 (N_7506,N_6346,N_6409);
nand U7507 (N_7507,N_6129,N_6223);
and U7508 (N_7508,N_6964,N_6421);
nor U7509 (N_7509,N_6119,N_6939);
and U7510 (N_7510,N_6185,N_6303);
or U7511 (N_7511,N_6417,N_6980);
nor U7512 (N_7512,N_6884,N_6225);
and U7513 (N_7513,N_6869,N_6176);
xnor U7514 (N_7514,N_6294,N_6989);
nand U7515 (N_7515,N_6998,N_6686);
xnor U7516 (N_7516,N_6111,N_6048);
nor U7517 (N_7517,N_6730,N_6114);
or U7518 (N_7518,N_6109,N_6545);
nor U7519 (N_7519,N_6315,N_6572);
nor U7520 (N_7520,N_6649,N_6789);
xor U7521 (N_7521,N_6496,N_6484);
nand U7522 (N_7522,N_6897,N_6483);
xnor U7523 (N_7523,N_6351,N_6477);
nand U7524 (N_7524,N_6736,N_6334);
xor U7525 (N_7525,N_6635,N_6059);
nor U7526 (N_7526,N_6756,N_6375);
nand U7527 (N_7527,N_6439,N_6108);
and U7528 (N_7528,N_6907,N_6276);
xor U7529 (N_7529,N_6791,N_6905);
xnor U7530 (N_7530,N_6767,N_6826);
and U7531 (N_7531,N_6453,N_6601);
or U7532 (N_7532,N_6890,N_6154);
nand U7533 (N_7533,N_6384,N_6415);
nor U7534 (N_7534,N_6902,N_6403);
nand U7535 (N_7535,N_6639,N_6383);
or U7536 (N_7536,N_6542,N_6737);
nor U7537 (N_7537,N_6539,N_6047);
and U7538 (N_7538,N_6726,N_6038);
and U7539 (N_7539,N_6188,N_6092);
nand U7540 (N_7540,N_6525,N_6000);
and U7541 (N_7541,N_6090,N_6863);
nor U7542 (N_7542,N_6406,N_6126);
nor U7543 (N_7543,N_6563,N_6760);
nand U7544 (N_7544,N_6930,N_6778);
and U7545 (N_7545,N_6978,N_6215);
and U7546 (N_7546,N_6497,N_6682);
and U7547 (N_7547,N_6947,N_6630);
or U7548 (N_7548,N_6921,N_6199);
and U7549 (N_7549,N_6460,N_6090);
or U7550 (N_7550,N_6293,N_6371);
or U7551 (N_7551,N_6838,N_6083);
nand U7552 (N_7552,N_6910,N_6745);
nand U7553 (N_7553,N_6104,N_6434);
nor U7554 (N_7554,N_6117,N_6834);
and U7555 (N_7555,N_6293,N_6601);
nor U7556 (N_7556,N_6563,N_6944);
and U7557 (N_7557,N_6402,N_6146);
and U7558 (N_7558,N_6177,N_6663);
nand U7559 (N_7559,N_6899,N_6665);
and U7560 (N_7560,N_6926,N_6947);
xor U7561 (N_7561,N_6645,N_6623);
and U7562 (N_7562,N_6043,N_6127);
nand U7563 (N_7563,N_6676,N_6845);
or U7564 (N_7564,N_6854,N_6529);
nand U7565 (N_7565,N_6914,N_6084);
and U7566 (N_7566,N_6728,N_6917);
nand U7567 (N_7567,N_6253,N_6225);
nand U7568 (N_7568,N_6710,N_6498);
nand U7569 (N_7569,N_6926,N_6184);
or U7570 (N_7570,N_6007,N_6613);
nand U7571 (N_7571,N_6367,N_6844);
xor U7572 (N_7572,N_6123,N_6401);
xor U7573 (N_7573,N_6161,N_6234);
nor U7574 (N_7574,N_6767,N_6711);
and U7575 (N_7575,N_6538,N_6853);
xnor U7576 (N_7576,N_6815,N_6879);
or U7577 (N_7577,N_6991,N_6315);
or U7578 (N_7578,N_6683,N_6772);
nand U7579 (N_7579,N_6273,N_6407);
and U7580 (N_7580,N_6311,N_6689);
nor U7581 (N_7581,N_6785,N_6313);
xnor U7582 (N_7582,N_6400,N_6687);
nand U7583 (N_7583,N_6251,N_6423);
or U7584 (N_7584,N_6627,N_6800);
xor U7585 (N_7585,N_6969,N_6700);
xnor U7586 (N_7586,N_6567,N_6237);
xor U7587 (N_7587,N_6162,N_6275);
nand U7588 (N_7588,N_6391,N_6076);
and U7589 (N_7589,N_6902,N_6301);
xor U7590 (N_7590,N_6248,N_6477);
or U7591 (N_7591,N_6718,N_6217);
nand U7592 (N_7592,N_6512,N_6610);
xor U7593 (N_7593,N_6518,N_6550);
or U7594 (N_7594,N_6432,N_6235);
nor U7595 (N_7595,N_6299,N_6539);
or U7596 (N_7596,N_6223,N_6036);
xor U7597 (N_7597,N_6391,N_6031);
nor U7598 (N_7598,N_6130,N_6241);
nand U7599 (N_7599,N_6694,N_6376);
and U7600 (N_7600,N_6173,N_6039);
nor U7601 (N_7601,N_6200,N_6529);
and U7602 (N_7602,N_6660,N_6221);
nor U7603 (N_7603,N_6753,N_6028);
xor U7604 (N_7604,N_6892,N_6291);
or U7605 (N_7605,N_6724,N_6570);
nand U7606 (N_7606,N_6318,N_6725);
nand U7607 (N_7607,N_6411,N_6190);
or U7608 (N_7608,N_6287,N_6325);
and U7609 (N_7609,N_6221,N_6644);
or U7610 (N_7610,N_6698,N_6312);
xnor U7611 (N_7611,N_6038,N_6081);
nand U7612 (N_7612,N_6281,N_6835);
nor U7613 (N_7613,N_6026,N_6477);
or U7614 (N_7614,N_6655,N_6903);
nor U7615 (N_7615,N_6985,N_6427);
xor U7616 (N_7616,N_6984,N_6250);
nor U7617 (N_7617,N_6163,N_6594);
nor U7618 (N_7618,N_6111,N_6333);
nand U7619 (N_7619,N_6160,N_6449);
nand U7620 (N_7620,N_6182,N_6550);
or U7621 (N_7621,N_6033,N_6489);
xor U7622 (N_7622,N_6385,N_6625);
nor U7623 (N_7623,N_6907,N_6791);
nor U7624 (N_7624,N_6295,N_6062);
and U7625 (N_7625,N_6252,N_6470);
xor U7626 (N_7626,N_6024,N_6595);
or U7627 (N_7627,N_6382,N_6296);
xnor U7628 (N_7628,N_6942,N_6630);
nor U7629 (N_7629,N_6265,N_6677);
nand U7630 (N_7630,N_6114,N_6268);
or U7631 (N_7631,N_6358,N_6459);
nand U7632 (N_7632,N_6720,N_6320);
or U7633 (N_7633,N_6721,N_6798);
xnor U7634 (N_7634,N_6684,N_6359);
and U7635 (N_7635,N_6740,N_6783);
nor U7636 (N_7636,N_6867,N_6757);
or U7637 (N_7637,N_6976,N_6638);
nand U7638 (N_7638,N_6941,N_6507);
and U7639 (N_7639,N_6205,N_6438);
nand U7640 (N_7640,N_6419,N_6416);
or U7641 (N_7641,N_6986,N_6441);
nor U7642 (N_7642,N_6946,N_6250);
nand U7643 (N_7643,N_6258,N_6396);
and U7644 (N_7644,N_6315,N_6095);
xor U7645 (N_7645,N_6905,N_6892);
nor U7646 (N_7646,N_6034,N_6257);
and U7647 (N_7647,N_6578,N_6678);
and U7648 (N_7648,N_6030,N_6836);
nand U7649 (N_7649,N_6048,N_6644);
xor U7650 (N_7650,N_6495,N_6411);
or U7651 (N_7651,N_6335,N_6844);
nand U7652 (N_7652,N_6252,N_6370);
nand U7653 (N_7653,N_6803,N_6523);
xor U7654 (N_7654,N_6941,N_6555);
xnor U7655 (N_7655,N_6793,N_6338);
nand U7656 (N_7656,N_6203,N_6944);
xor U7657 (N_7657,N_6046,N_6684);
or U7658 (N_7658,N_6906,N_6914);
nor U7659 (N_7659,N_6629,N_6215);
nand U7660 (N_7660,N_6870,N_6029);
and U7661 (N_7661,N_6163,N_6217);
xnor U7662 (N_7662,N_6135,N_6241);
or U7663 (N_7663,N_6820,N_6477);
xor U7664 (N_7664,N_6527,N_6523);
nor U7665 (N_7665,N_6721,N_6176);
nand U7666 (N_7666,N_6042,N_6851);
nand U7667 (N_7667,N_6441,N_6791);
xor U7668 (N_7668,N_6889,N_6946);
xnor U7669 (N_7669,N_6442,N_6014);
or U7670 (N_7670,N_6031,N_6621);
nor U7671 (N_7671,N_6347,N_6912);
nor U7672 (N_7672,N_6217,N_6354);
xnor U7673 (N_7673,N_6707,N_6921);
and U7674 (N_7674,N_6460,N_6547);
and U7675 (N_7675,N_6166,N_6110);
and U7676 (N_7676,N_6473,N_6030);
and U7677 (N_7677,N_6748,N_6508);
nand U7678 (N_7678,N_6182,N_6986);
and U7679 (N_7679,N_6965,N_6605);
nor U7680 (N_7680,N_6121,N_6231);
xor U7681 (N_7681,N_6537,N_6989);
xnor U7682 (N_7682,N_6363,N_6319);
xnor U7683 (N_7683,N_6025,N_6000);
nor U7684 (N_7684,N_6799,N_6711);
nand U7685 (N_7685,N_6578,N_6259);
nand U7686 (N_7686,N_6756,N_6964);
or U7687 (N_7687,N_6284,N_6415);
or U7688 (N_7688,N_6394,N_6293);
or U7689 (N_7689,N_6222,N_6835);
xor U7690 (N_7690,N_6818,N_6541);
or U7691 (N_7691,N_6859,N_6981);
nand U7692 (N_7692,N_6063,N_6216);
xnor U7693 (N_7693,N_6806,N_6873);
nand U7694 (N_7694,N_6071,N_6643);
or U7695 (N_7695,N_6857,N_6238);
or U7696 (N_7696,N_6175,N_6842);
or U7697 (N_7697,N_6394,N_6758);
or U7698 (N_7698,N_6369,N_6752);
or U7699 (N_7699,N_6478,N_6951);
nand U7700 (N_7700,N_6660,N_6214);
and U7701 (N_7701,N_6751,N_6986);
or U7702 (N_7702,N_6376,N_6236);
nor U7703 (N_7703,N_6769,N_6125);
nand U7704 (N_7704,N_6972,N_6403);
nand U7705 (N_7705,N_6221,N_6456);
and U7706 (N_7706,N_6378,N_6346);
or U7707 (N_7707,N_6144,N_6898);
nor U7708 (N_7708,N_6319,N_6918);
xnor U7709 (N_7709,N_6871,N_6491);
xnor U7710 (N_7710,N_6966,N_6421);
nor U7711 (N_7711,N_6256,N_6423);
or U7712 (N_7712,N_6748,N_6504);
or U7713 (N_7713,N_6855,N_6429);
or U7714 (N_7714,N_6796,N_6086);
nor U7715 (N_7715,N_6495,N_6809);
or U7716 (N_7716,N_6601,N_6215);
nor U7717 (N_7717,N_6626,N_6563);
nor U7718 (N_7718,N_6332,N_6257);
xnor U7719 (N_7719,N_6896,N_6319);
and U7720 (N_7720,N_6309,N_6373);
xnor U7721 (N_7721,N_6908,N_6048);
or U7722 (N_7722,N_6222,N_6619);
nand U7723 (N_7723,N_6683,N_6913);
nand U7724 (N_7724,N_6504,N_6294);
or U7725 (N_7725,N_6489,N_6421);
xnor U7726 (N_7726,N_6411,N_6231);
or U7727 (N_7727,N_6883,N_6413);
xnor U7728 (N_7728,N_6742,N_6675);
nor U7729 (N_7729,N_6023,N_6870);
and U7730 (N_7730,N_6181,N_6770);
or U7731 (N_7731,N_6004,N_6743);
and U7732 (N_7732,N_6877,N_6001);
and U7733 (N_7733,N_6586,N_6232);
or U7734 (N_7734,N_6280,N_6579);
xnor U7735 (N_7735,N_6987,N_6747);
xor U7736 (N_7736,N_6779,N_6558);
xor U7737 (N_7737,N_6217,N_6682);
and U7738 (N_7738,N_6365,N_6686);
or U7739 (N_7739,N_6240,N_6350);
xor U7740 (N_7740,N_6709,N_6008);
nand U7741 (N_7741,N_6308,N_6517);
nand U7742 (N_7742,N_6651,N_6858);
nor U7743 (N_7743,N_6951,N_6015);
and U7744 (N_7744,N_6893,N_6168);
nand U7745 (N_7745,N_6665,N_6825);
nand U7746 (N_7746,N_6366,N_6589);
and U7747 (N_7747,N_6414,N_6551);
xor U7748 (N_7748,N_6399,N_6800);
nand U7749 (N_7749,N_6359,N_6167);
and U7750 (N_7750,N_6856,N_6433);
or U7751 (N_7751,N_6619,N_6710);
nor U7752 (N_7752,N_6088,N_6996);
or U7753 (N_7753,N_6870,N_6474);
nand U7754 (N_7754,N_6201,N_6788);
nand U7755 (N_7755,N_6175,N_6973);
xor U7756 (N_7756,N_6796,N_6672);
nand U7757 (N_7757,N_6055,N_6395);
and U7758 (N_7758,N_6990,N_6598);
xnor U7759 (N_7759,N_6937,N_6281);
and U7760 (N_7760,N_6147,N_6415);
nor U7761 (N_7761,N_6240,N_6806);
xor U7762 (N_7762,N_6622,N_6363);
xnor U7763 (N_7763,N_6176,N_6682);
xor U7764 (N_7764,N_6091,N_6432);
nand U7765 (N_7765,N_6024,N_6149);
and U7766 (N_7766,N_6552,N_6267);
or U7767 (N_7767,N_6997,N_6904);
and U7768 (N_7768,N_6664,N_6890);
nor U7769 (N_7769,N_6747,N_6447);
and U7770 (N_7770,N_6633,N_6107);
or U7771 (N_7771,N_6393,N_6058);
or U7772 (N_7772,N_6579,N_6414);
nor U7773 (N_7773,N_6287,N_6986);
and U7774 (N_7774,N_6206,N_6647);
and U7775 (N_7775,N_6425,N_6214);
nor U7776 (N_7776,N_6581,N_6535);
or U7777 (N_7777,N_6843,N_6143);
xnor U7778 (N_7778,N_6926,N_6283);
or U7779 (N_7779,N_6860,N_6157);
and U7780 (N_7780,N_6875,N_6591);
nor U7781 (N_7781,N_6662,N_6466);
nor U7782 (N_7782,N_6006,N_6679);
xnor U7783 (N_7783,N_6256,N_6126);
nor U7784 (N_7784,N_6856,N_6143);
or U7785 (N_7785,N_6961,N_6608);
or U7786 (N_7786,N_6796,N_6782);
or U7787 (N_7787,N_6944,N_6878);
nand U7788 (N_7788,N_6990,N_6314);
nor U7789 (N_7789,N_6111,N_6565);
and U7790 (N_7790,N_6264,N_6714);
and U7791 (N_7791,N_6079,N_6777);
or U7792 (N_7792,N_6636,N_6908);
nor U7793 (N_7793,N_6347,N_6501);
nor U7794 (N_7794,N_6465,N_6417);
nor U7795 (N_7795,N_6406,N_6409);
nor U7796 (N_7796,N_6570,N_6403);
xor U7797 (N_7797,N_6780,N_6984);
and U7798 (N_7798,N_6209,N_6915);
xnor U7799 (N_7799,N_6286,N_6683);
xnor U7800 (N_7800,N_6075,N_6040);
and U7801 (N_7801,N_6107,N_6892);
or U7802 (N_7802,N_6955,N_6136);
nand U7803 (N_7803,N_6167,N_6222);
xnor U7804 (N_7804,N_6125,N_6087);
nand U7805 (N_7805,N_6258,N_6280);
xnor U7806 (N_7806,N_6270,N_6062);
nor U7807 (N_7807,N_6068,N_6326);
and U7808 (N_7808,N_6304,N_6273);
xnor U7809 (N_7809,N_6895,N_6074);
and U7810 (N_7810,N_6977,N_6733);
nor U7811 (N_7811,N_6925,N_6657);
xnor U7812 (N_7812,N_6749,N_6716);
or U7813 (N_7813,N_6104,N_6469);
or U7814 (N_7814,N_6935,N_6587);
or U7815 (N_7815,N_6574,N_6616);
or U7816 (N_7816,N_6343,N_6618);
nor U7817 (N_7817,N_6833,N_6181);
nor U7818 (N_7818,N_6771,N_6087);
or U7819 (N_7819,N_6329,N_6874);
and U7820 (N_7820,N_6471,N_6837);
or U7821 (N_7821,N_6214,N_6645);
xnor U7822 (N_7822,N_6023,N_6744);
nand U7823 (N_7823,N_6091,N_6816);
xor U7824 (N_7824,N_6152,N_6492);
and U7825 (N_7825,N_6583,N_6090);
or U7826 (N_7826,N_6451,N_6736);
nor U7827 (N_7827,N_6380,N_6063);
or U7828 (N_7828,N_6123,N_6074);
and U7829 (N_7829,N_6670,N_6296);
nor U7830 (N_7830,N_6507,N_6359);
or U7831 (N_7831,N_6554,N_6685);
or U7832 (N_7832,N_6486,N_6277);
xor U7833 (N_7833,N_6416,N_6480);
and U7834 (N_7834,N_6066,N_6856);
or U7835 (N_7835,N_6516,N_6671);
or U7836 (N_7836,N_6651,N_6491);
nand U7837 (N_7837,N_6132,N_6071);
and U7838 (N_7838,N_6457,N_6404);
and U7839 (N_7839,N_6899,N_6245);
nor U7840 (N_7840,N_6218,N_6261);
or U7841 (N_7841,N_6539,N_6940);
nand U7842 (N_7842,N_6184,N_6118);
nor U7843 (N_7843,N_6118,N_6510);
nand U7844 (N_7844,N_6889,N_6880);
or U7845 (N_7845,N_6432,N_6220);
xnor U7846 (N_7846,N_6504,N_6991);
nand U7847 (N_7847,N_6793,N_6795);
xor U7848 (N_7848,N_6716,N_6162);
or U7849 (N_7849,N_6021,N_6579);
xor U7850 (N_7850,N_6116,N_6510);
or U7851 (N_7851,N_6598,N_6745);
xor U7852 (N_7852,N_6933,N_6543);
nand U7853 (N_7853,N_6201,N_6078);
nor U7854 (N_7854,N_6595,N_6317);
or U7855 (N_7855,N_6529,N_6883);
xnor U7856 (N_7856,N_6420,N_6186);
nor U7857 (N_7857,N_6316,N_6448);
nor U7858 (N_7858,N_6591,N_6444);
nand U7859 (N_7859,N_6886,N_6265);
nand U7860 (N_7860,N_6155,N_6918);
and U7861 (N_7861,N_6615,N_6937);
or U7862 (N_7862,N_6876,N_6363);
nor U7863 (N_7863,N_6441,N_6267);
nand U7864 (N_7864,N_6020,N_6508);
or U7865 (N_7865,N_6072,N_6450);
xnor U7866 (N_7866,N_6363,N_6617);
or U7867 (N_7867,N_6930,N_6515);
nor U7868 (N_7868,N_6909,N_6649);
nor U7869 (N_7869,N_6035,N_6514);
nand U7870 (N_7870,N_6623,N_6212);
xnor U7871 (N_7871,N_6124,N_6965);
xor U7872 (N_7872,N_6636,N_6460);
or U7873 (N_7873,N_6003,N_6376);
and U7874 (N_7874,N_6384,N_6506);
and U7875 (N_7875,N_6586,N_6735);
nor U7876 (N_7876,N_6742,N_6895);
and U7877 (N_7877,N_6072,N_6464);
xnor U7878 (N_7878,N_6278,N_6543);
nor U7879 (N_7879,N_6706,N_6043);
xor U7880 (N_7880,N_6946,N_6864);
and U7881 (N_7881,N_6356,N_6054);
xor U7882 (N_7882,N_6587,N_6533);
nor U7883 (N_7883,N_6913,N_6036);
nand U7884 (N_7884,N_6145,N_6994);
nand U7885 (N_7885,N_6561,N_6139);
and U7886 (N_7886,N_6218,N_6589);
nand U7887 (N_7887,N_6717,N_6913);
xor U7888 (N_7888,N_6494,N_6070);
xnor U7889 (N_7889,N_6015,N_6155);
nand U7890 (N_7890,N_6573,N_6337);
and U7891 (N_7891,N_6433,N_6763);
and U7892 (N_7892,N_6489,N_6276);
nand U7893 (N_7893,N_6282,N_6528);
xor U7894 (N_7894,N_6060,N_6338);
and U7895 (N_7895,N_6340,N_6656);
or U7896 (N_7896,N_6709,N_6303);
nand U7897 (N_7897,N_6672,N_6352);
and U7898 (N_7898,N_6670,N_6333);
nor U7899 (N_7899,N_6841,N_6082);
nand U7900 (N_7900,N_6576,N_6378);
xor U7901 (N_7901,N_6689,N_6981);
nand U7902 (N_7902,N_6256,N_6018);
nor U7903 (N_7903,N_6359,N_6697);
xor U7904 (N_7904,N_6777,N_6019);
xnor U7905 (N_7905,N_6376,N_6290);
nand U7906 (N_7906,N_6276,N_6283);
and U7907 (N_7907,N_6730,N_6197);
xor U7908 (N_7908,N_6855,N_6222);
nor U7909 (N_7909,N_6979,N_6252);
xor U7910 (N_7910,N_6036,N_6917);
or U7911 (N_7911,N_6642,N_6078);
nor U7912 (N_7912,N_6458,N_6203);
nor U7913 (N_7913,N_6632,N_6627);
and U7914 (N_7914,N_6981,N_6109);
or U7915 (N_7915,N_6912,N_6116);
xnor U7916 (N_7916,N_6607,N_6552);
xor U7917 (N_7917,N_6756,N_6502);
or U7918 (N_7918,N_6854,N_6760);
nand U7919 (N_7919,N_6080,N_6011);
or U7920 (N_7920,N_6886,N_6049);
and U7921 (N_7921,N_6906,N_6518);
nand U7922 (N_7922,N_6462,N_6614);
nand U7923 (N_7923,N_6650,N_6658);
xor U7924 (N_7924,N_6253,N_6571);
nor U7925 (N_7925,N_6212,N_6772);
xor U7926 (N_7926,N_6614,N_6303);
xor U7927 (N_7927,N_6599,N_6301);
and U7928 (N_7928,N_6543,N_6071);
and U7929 (N_7929,N_6794,N_6100);
nor U7930 (N_7930,N_6833,N_6636);
xnor U7931 (N_7931,N_6503,N_6419);
or U7932 (N_7932,N_6469,N_6625);
xor U7933 (N_7933,N_6315,N_6376);
and U7934 (N_7934,N_6899,N_6714);
xor U7935 (N_7935,N_6150,N_6834);
or U7936 (N_7936,N_6170,N_6704);
nand U7937 (N_7937,N_6158,N_6423);
nand U7938 (N_7938,N_6017,N_6831);
xnor U7939 (N_7939,N_6980,N_6481);
nor U7940 (N_7940,N_6370,N_6345);
nand U7941 (N_7941,N_6032,N_6199);
nand U7942 (N_7942,N_6002,N_6746);
or U7943 (N_7943,N_6875,N_6711);
or U7944 (N_7944,N_6512,N_6242);
nor U7945 (N_7945,N_6327,N_6979);
xnor U7946 (N_7946,N_6453,N_6475);
nor U7947 (N_7947,N_6312,N_6678);
and U7948 (N_7948,N_6993,N_6050);
xnor U7949 (N_7949,N_6703,N_6539);
nand U7950 (N_7950,N_6215,N_6367);
xnor U7951 (N_7951,N_6944,N_6760);
nand U7952 (N_7952,N_6172,N_6020);
and U7953 (N_7953,N_6670,N_6257);
xor U7954 (N_7954,N_6090,N_6298);
or U7955 (N_7955,N_6383,N_6840);
or U7956 (N_7956,N_6641,N_6326);
xnor U7957 (N_7957,N_6864,N_6087);
and U7958 (N_7958,N_6190,N_6933);
xnor U7959 (N_7959,N_6327,N_6167);
nand U7960 (N_7960,N_6105,N_6126);
or U7961 (N_7961,N_6280,N_6110);
or U7962 (N_7962,N_6119,N_6609);
nor U7963 (N_7963,N_6634,N_6050);
nand U7964 (N_7964,N_6112,N_6645);
and U7965 (N_7965,N_6080,N_6196);
nand U7966 (N_7966,N_6021,N_6367);
xor U7967 (N_7967,N_6782,N_6297);
nor U7968 (N_7968,N_6574,N_6409);
nor U7969 (N_7969,N_6100,N_6451);
nand U7970 (N_7970,N_6726,N_6836);
nand U7971 (N_7971,N_6125,N_6696);
xnor U7972 (N_7972,N_6796,N_6542);
and U7973 (N_7973,N_6904,N_6533);
nand U7974 (N_7974,N_6508,N_6833);
or U7975 (N_7975,N_6196,N_6052);
nor U7976 (N_7976,N_6270,N_6186);
nand U7977 (N_7977,N_6025,N_6525);
nand U7978 (N_7978,N_6134,N_6366);
and U7979 (N_7979,N_6707,N_6415);
or U7980 (N_7980,N_6628,N_6997);
nand U7981 (N_7981,N_6125,N_6455);
nor U7982 (N_7982,N_6192,N_6139);
nor U7983 (N_7983,N_6560,N_6475);
xor U7984 (N_7984,N_6224,N_6995);
nor U7985 (N_7985,N_6855,N_6728);
and U7986 (N_7986,N_6703,N_6582);
and U7987 (N_7987,N_6397,N_6176);
nor U7988 (N_7988,N_6786,N_6571);
and U7989 (N_7989,N_6654,N_6924);
xor U7990 (N_7990,N_6145,N_6151);
or U7991 (N_7991,N_6397,N_6016);
and U7992 (N_7992,N_6946,N_6688);
xor U7993 (N_7993,N_6090,N_6485);
xor U7994 (N_7994,N_6936,N_6696);
or U7995 (N_7995,N_6993,N_6302);
and U7996 (N_7996,N_6100,N_6311);
nor U7997 (N_7997,N_6666,N_6369);
nor U7998 (N_7998,N_6312,N_6816);
nor U7999 (N_7999,N_6281,N_6997);
xnor U8000 (N_8000,N_7009,N_7965);
and U8001 (N_8001,N_7938,N_7243);
or U8002 (N_8002,N_7337,N_7699);
nor U8003 (N_8003,N_7176,N_7486);
xnor U8004 (N_8004,N_7940,N_7906);
xnor U8005 (N_8005,N_7682,N_7917);
and U8006 (N_8006,N_7663,N_7128);
nand U8007 (N_8007,N_7905,N_7999);
and U8008 (N_8008,N_7186,N_7133);
xnor U8009 (N_8009,N_7469,N_7509);
nor U8010 (N_8010,N_7560,N_7242);
nor U8011 (N_8011,N_7972,N_7416);
xor U8012 (N_8012,N_7209,N_7245);
nand U8013 (N_8013,N_7419,N_7830);
nor U8014 (N_8014,N_7949,N_7646);
xnor U8015 (N_8015,N_7867,N_7052);
or U8016 (N_8016,N_7527,N_7078);
or U8017 (N_8017,N_7692,N_7013);
xnor U8018 (N_8018,N_7430,N_7409);
xor U8019 (N_8019,N_7195,N_7281);
nor U8020 (N_8020,N_7293,N_7642);
nor U8021 (N_8021,N_7810,N_7444);
or U8022 (N_8022,N_7320,N_7029);
xnor U8023 (N_8023,N_7945,N_7261);
nor U8024 (N_8024,N_7708,N_7177);
and U8025 (N_8025,N_7066,N_7207);
xnor U8026 (N_8026,N_7196,N_7655);
nor U8027 (N_8027,N_7923,N_7382);
nand U8028 (N_8028,N_7262,N_7422);
and U8029 (N_8029,N_7350,N_7057);
and U8030 (N_8030,N_7908,N_7211);
and U8031 (N_8031,N_7820,N_7408);
or U8032 (N_8032,N_7405,N_7815);
nor U8033 (N_8033,N_7055,N_7662);
or U8034 (N_8034,N_7926,N_7226);
and U8035 (N_8035,N_7421,N_7754);
nor U8036 (N_8036,N_7983,N_7311);
nor U8037 (N_8037,N_7377,N_7324);
and U8038 (N_8038,N_7470,N_7204);
or U8039 (N_8039,N_7121,N_7755);
nor U8040 (N_8040,N_7499,N_7330);
and U8041 (N_8041,N_7929,N_7158);
or U8042 (N_8042,N_7963,N_7156);
and U8043 (N_8043,N_7877,N_7436);
xor U8044 (N_8044,N_7956,N_7290);
nand U8045 (N_8045,N_7059,N_7417);
nor U8046 (N_8046,N_7076,N_7615);
or U8047 (N_8047,N_7811,N_7855);
and U8048 (N_8048,N_7305,N_7455);
nand U8049 (N_8049,N_7414,N_7643);
xnor U8050 (N_8050,N_7959,N_7909);
xor U8051 (N_8051,N_7145,N_7309);
xor U8052 (N_8052,N_7619,N_7691);
nor U8053 (N_8053,N_7545,N_7611);
or U8054 (N_8054,N_7171,N_7928);
nor U8055 (N_8055,N_7550,N_7962);
or U8056 (N_8056,N_7501,N_7990);
and U8057 (N_8057,N_7448,N_7939);
nor U8058 (N_8058,N_7315,N_7716);
and U8059 (N_8059,N_7944,N_7771);
and U8060 (N_8060,N_7367,N_7572);
or U8061 (N_8061,N_7236,N_7331);
or U8062 (N_8062,N_7368,N_7825);
nand U8063 (N_8063,N_7342,N_7732);
and U8064 (N_8064,N_7707,N_7061);
or U8065 (N_8065,N_7056,N_7102);
and U8066 (N_8066,N_7362,N_7542);
xnor U8067 (N_8067,N_7523,N_7679);
or U8068 (N_8068,N_7048,N_7996);
or U8069 (N_8069,N_7286,N_7757);
xnor U8070 (N_8070,N_7849,N_7902);
nor U8071 (N_8071,N_7396,N_7374);
nand U8072 (N_8072,N_7510,N_7473);
or U8073 (N_8073,N_7298,N_7080);
or U8074 (N_8074,N_7168,N_7987);
nor U8075 (N_8075,N_7897,N_7182);
or U8076 (N_8076,N_7622,N_7117);
and U8077 (N_8077,N_7528,N_7150);
or U8078 (N_8078,N_7251,N_7552);
nand U8079 (N_8079,N_7788,N_7887);
nand U8080 (N_8080,N_7934,N_7793);
and U8081 (N_8081,N_7652,N_7975);
or U8082 (N_8082,N_7860,N_7265);
or U8083 (N_8083,N_7138,N_7508);
and U8084 (N_8084,N_7296,N_7600);
or U8085 (N_8085,N_7210,N_7667);
nand U8086 (N_8086,N_7152,N_7673);
or U8087 (N_8087,N_7427,N_7933);
or U8088 (N_8088,N_7014,N_7759);
and U8089 (N_8089,N_7961,N_7481);
nand U8090 (N_8090,N_7323,N_7719);
or U8091 (N_8091,N_7852,N_7203);
nor U8092 (N_8092,N_7651,N_7641);
nor U8093 (N_8093,N_7912,N_7060);
and U8094 (N_8094,N_7636,N_7760);
nor U8095 (N_8095,N_7037,N_7482);
and U8096 (N_8096,N_7118,N_7162);
and U8097 (N_8097,N_7503,N_7273);
and U8098 (N_8098,N_7089,N_7927);
or U8099 (N_8099,N_7697,N_7573);
or U8100 (N_8100,N_7595,N_7774);
nor U8101 (N_8101,N_7984,N_7023);
nand U8102 (N_8102,N_7005,N_7558);
and U8103 (N_8103,N_7058,N_7395);
nand U8104 (N_8104,N_7034,N_7618);
or U8105 (N_8105,N_7986,N_7846);
nor U8106 (N_8106,N_7890,N_7025);
and U8107 (N_8107,N_7252,N_7365);
nand U8108 (N_8108,N_7488,N_7456);
and U8109 (N_8109,N_7935,N_7590);
nand U8110 (N_8110,N_7791,N_7910);
nor U8111 (N_8111,N_7522,N_7921);
or U8112 (N_8112,N_7106,N_7109);
xnor U8113 (N_8113,N_7340,N_7457);
or U8114 (N_8114,N_7865,N_7792);
xnor U8115 (N_8115,N_7997,N_7690);
or U8116 (N_8116,N_7178,N_7828);
nand U8117 (N_8117,N_7267,N_7954);
nand U8118 (N_8118,N_7586,N_7404);
nor U8119 (N_8119,N_7659,N_7274);
or U8120 (N_8120,N_7842,N_7863);
nand U8121 (N_8121,N_7534,N_7838);
nor U8122 (N_8122,N_7982,N_7310);
xnor U8123 (N_8123,N_7447,N_7010);
nor U8124 (N_8124,N_7445,N_7706);
nand U8125 (N_8125,N_7442,N_7571);
xor U8126 (N_8126,N_7094,N_7597);
and U8127 (N_8127,N_7313,N_7151);
or U8128 (N_8128,N_7717,N_7072);
nor U8129 (N_8129,N_7533,N_7745);
nand U8130 (N_8130,N_7208,N_7360);
nand U8131 (N_8131,N_7466,N_7785);
nor U8132 (N_8132,N_7988,N_7345);
xor U8133 (N_8133,N_7153,N_7547);
xor U8134 (N_8134,N_7389,N_7705);
or U8135 (N_8135,N_7570,N_7750);
nor U8136 (N_8136,N_7016,N_7770);
and U8137 (N_8137,N_7981,N_7976);
and U8138 (N_8138,N_7191,N_7036);
nor U8139 (N_8139,N_7798,N_7143);
nand U8140 (N_8140,N_7175,N_7278);
and U8141 (N_8141,N_7915,N_7853);
xnor U8142 (N_8142,N_7703,N_7285);
nand U8143 (N_8143,N_7260,N_7380);
nor U8144 (N_8144,N_7901,N_7064);
nor U8145 (N_8145,N_7288,N_7583);
or U8146 (N_8146,N_7730,N_7603);
or U8147 (N_8147,N_7955,N_7598);
nor U8148 (N_8148,N_7322,N_7539);
xor U8149 (N_8149,N_7739,N_7189);
and U8150 (N_8150,N_7063,N_7644);
nand U8151 (N_8151,N_7392,N_7731);
or U8152 (N_8152,N_7647,N_7297);
nand U8153 (N_8153,N_7379,N_7454);
and U8154 (N_8154,N_7049,N_7140);
and U8155 (N_8155,N_7301,N_7067);
and U8156 (N_8156,N_7683,N_7230);
nand U8157 (N_8157,N_7007,N_7361);
and U8158 (N_8158,N_7631,N_7300);
nand U8159 (N_8159,N_7904,N_7526);
or U8160 (N_8160,N_7681,N_7213);
nor U8161 (N_8161,N_7784,N_7824);
or U8162 (N_8162,N_7781,N_7462);
or U8163 (N_8163,N_7876,N_7335);
nor U8164 (N_8164,N_7639,N_7507);
xnor U8165 (N_8165,N_7174,N_7864);
and U8166 (N_8166,N_7347,N_7835);
nor U8167 (N_8167,N_7868,N_7500);
and U8168 (N_8168,N_7778,N_7530);
xor U8169 (N_8169,N_7812,N_7188);
xor U8170 (N_8170,N_7856,N_7587);
xnor U8171 (N_8171,N_7660,N_7329);
or U8172 (N_8172,N_7187,N_7390);
nand U8173 (N_8173,N_7479,N_7450);
or U8174 (N_8174,N_7726,N_7870);
nor U8175 (N_8175,N_7688,N_7371);
xor U8176 (N_8176,N_7967,N_7718);
or U8177 (N_8177,N_7748,N_7913);
nor U8178 (N_8178,N_7201,N_7391);
or U8179 (N_8179,N_7253,N_7773);
nor U8180 (N_8180,N_7093,N_7991);
or U8181 (N_8181,N_7665,N_7775);
or U8182 (N_8182,N_7139,N_7666);
or U8183 (N_8183,N_7544,N_7831);
nand U8184 (N_8184,N_7410,N_7294);
and U8185 (N_8185,N_7752,N_7766);
nor U8186 (N_8186,N_7426,N_7376);
and U8187 (N_8187,N_7515,N_7104);
nand U8188 (N_8188,N_7763,N_7875);
or U8189 (N_8189,N_7432,N_7556);
or U8190 (N_8190,N_7847,N_7483);
xnor U8191 (N_8191,N_7234,N_7433);
and U8192 (N_8192,N_7053,N_7979);
nor U8193 (N_8193,N_7817,N_7964);
or U8194 (N_8194,N_7202,N_7924);
nand U8195 (N_8195,N_7489,N_7497);
xnor U8196 (N_8196,N_7585,N_7649);
or U8197 (N_8197,N_7369,N_7768);
xnor U8198 (N_8198,N_7993,N_7415);
and U8199 (N_8199,N_7710,N_7640);
xnor U8200 (N_8200,N_7460,N_7446);
or U8201 (N_8201,N_7173,N_7412);
xor U8202 (N_8202,N_7024,N_7711);
xnor U8203 (N_8203,N_7263,N_7630);
nor U8204 (N_8204,N_7065,N_7635);
nand U8205 (N_8205,N_7363,N_7217);
and U8206 (N_8206,N_7492,N_7687);
or U8207 (N_8207,N_7018,N_7169);
nand U8208 (N_8208,N_7357,N_7882);
nor U8209 (N_8209,N_7941,N_7095);
nor U8210 (N_8210,N_7004,N_7519);
and U8211 (N_8211,N_7762,N_7308);
nor U8212 (N_8212,N_7678,N_7664);
nor U8213 (N_8213,N_7127,N_7696);
nand U8214 (N_8214,N_7712,N_7073);
xor U8215 (N_8215,N_7850,N_7468);
and U8216 (N_8216,N_7077,N_7126);
and U8217 (N_8217,N_7969,N_7931);
or U8218 (N_8218,N_7998,N_7657);
or U8219 (N_8219,N_7675,N_7465);
or U8220 (N_8220,N_7453,N_7616);
and U8221 (N_8221,N_7799,N_7062);
nand U8222 (N_8222,N_7898,N_7353);
nor U8223 (N_8223,N_7818,N_7802);
and U8224 (N_8224,N_7193,N_7992);
or U8225 (N_8225,N_7304,N_7540);
or U8226 (N_8226,N_7861,N_7306);
nand U8227 (N_8227,N_7449,N_7038);
nand U8228 (N_8228,N_7943,N_7275);
xnor U8229 (N_8229,N_7319,N_7536);
or U8230 (N_8230,N_7741,N_7676);
or U8231 (N_8231,N_7756,N_7366);
or U8232 (N_8232,N_7030,N_7554);
and U8233 (N_8233,N_7411,N_7922);
or U8234 (N_8234,N_7235,N_7378);
and U8235 (N_8235,N_7223,N_7241);
or U8236 (N_8236,N_7420,N_7521);
nor U8237 (N_8237,N_7645,N_7028);
nor U8238 (N_8238,N_7255,N_7008);
or U8239 (N_8239,N_7561,N_7478);
or U8240 (N_8240,N_7787,N_7406);
xnor U8241 (N_8241,N_7511,N_7129);
nand U8242 (N_8242,N_7776,N_7686);
or U8243 (N_8243,N_7567,N_7936);
or U8244 (N_8244,N_7364,N_7295);
and U8245 (N_8245,N_7238,N_7985);
xor U8246 (N_8246,N_7822,N_7441);
nor U8247 (N_8247,N_7167,N_7989);
nor U8248 (N_8248,N_7225,N_7740);
or U8249 (N_8249,N_7035,N_7485);
and U8250 (N_8250,N_7249,N_7866);
or U8251 (N_8251,N_7183,N_7702);
or U8252 (N_8252,N_7518,N_7612);
and U8253 (N_8253,N_7862,N_7170);
and U8254 (N_8254,N_7351,N_7907);
nand U8255 (N_8255,N_7885,N_7809);
xnor U8256 (N_8256,N_7020,N_7881);
or U8257 (N_8257,N_7769,N_7327);
and U8258 (N_8258,N_7565,N_7385);
or U8259 (N_8259,N_7834,N_7423);
or U8260 (N_8260,N_7474,N_7086);
and U8261 (N_8261,N_7532,N_7596);
xnor U8262 (N_8262,N_7487,N_7475);
nor U8263 (N_8263,N_7840,N_7484);
nand U8264 (N_8264,N_7107,N_7247);
xnor U8265 (N_8265,N_7617,N_7805);
nor U8266 (N_8266,N_7312,N_7685);
or U8267 (N_8267,N_7514,N_7950);
nor U8268 (N_8268,N_7591,N_7480);
xnor U8269 (N_8269,N_7701,N_7393);
xor U8270 (N_8270,N_7054,N_7689);
xor U8271 (N_8271,N_7092,N_7650);
nand U8272 (N_8272,N_7179,N_7033);
nor U8273 (N_8273,N_7733,N_7859);
nor U8274 (N_8274,N_7000,N_7797);
xnor U8275 (N_8275,N_7398,N_7535);
nand U8276 (N_8276,N_7264,N_7738);
or U8277 (N_8277,N_7088,N_7477);
nand U8278 (N_8278,N_7737,N_7800);
nor U8279 (N_8279,N_7397,N_7704);
nand U8280 (N_8280,N_7872,N_7370);
and U8281 (N_8281,N_7506,N_7541);
nand U8282 (N_8282,N_7592,N_7011);
xor U8283 (N_8283,N_7914,N_7628);
xnor U8284 (N_8284,N_7043,N_7873);
or U8285 (N_8285,N_7761,N_7584);
nand U8286 (N_8286,N_7458,N_7464);
or U8287 (N_8287,N_7021,N_7579);
nor U8288 (N_8288,N_7075,N_7874);
and U8289 (N_8289,N_7266,N_7589);
nand U8290 (N_8290,N_7157,N_7123);
xor U8291 (N_8291,N_7283,N_7082);
or U8292 (N_8292,N_7957,N_7538);
xnor U8293 (N_8293,N_7715,N_7125);
nor U8294 (N_8294,N_7400,N_7698);
and U8295 (N_8295,N_7978,N_7149);
xor U8296 (N_8296,N_7858,N_7229);
and U8297 (N_8297,N_7299,N_7851);
nor U8298 (N_8298,N_7105,N_7947);
and U8299 (N_8299,N_7120,N_7879);
nor U8300 (N_8300,N_7142,N_7884);
nand U8301 (N_8301,N_7747,N_7974);
nor U8302 (N_8302,N_7973,N_7594);
and U8303 (N_8303,N_7661,N_7680);
xor U8304 (N_8304,N_7517,N_7493);
nor U8305 (N_8305,N_7399,N_7823);
nand U8306 (N_8306,N_7440,N_7601);
xnor U8307 (N_8307,N_7557,N_7581);
and U8308 (N_8308,N_7767,N_7531);
xnor U8309 (N_8309,N_7165,N_7069);
nor U8310 (N_8310,N_7184,N_7279);
xor U8311 (N_8311,N_7130,N_7746);
nand U8312 (N_8312,N_7548,N_7796);
and U8313 (N_8313,N_7880,N_7816);
nand U8314 (N_8314,N_7231,N_7958);
or U8315 (N_8315,N_7632,N_7513);
and U8316 (N_8316,N_7192,N_7359);
nand U8317 (N_8317,N_7046,N_7111);
or U8318 (N_8318,N_7735,N_7491);
or U8319 (N_8319,N_7566,N_7224);
nor U8320 (N_8320,N_7610,N_7228);
xnor U8321 (N_8321,N_7837,N_7103);
nor U8322 (N_8322,N_7751,N_7257);
and U8323 (N_8323,N_7633,N_7159);
nor U8324 (N_8324,N_7424,N_7833);
nor U8325 (N_8325,N_7505,N_7790);
nand U8326 (N_8326,N_7725,N_7002);
or U8327 (N_8327,N_7205,N_7578);
or U8328 (N_8328,N_7083,N_7339);
nand U8329 (N_8329,N_7219,N_7119);
or U8330 (N_8330,N_7071,N_7100);
or U8331 (N_8331,N_7074,N_7047);
nor U8332 (N_8332,N_7878,N_7749);
and U8333 (N_8333,N_7693,N_7670);
xnor U8334 (N_8334,N_7272,N_7222);
nand U8335 (N_8335,N_7250,N_7714);
xnor U8336 (N_8336,N_7172,N_7218);
nand U8337 (N_8337,N_7634,N_7808);
and U8338 (N_8338,N_7434,N_7899);
nand U8339 (N_8339,N_7626,N_7081);
nor U8340 (N_8340,N_7141,N_7180);
and U8341 (N_8341,N_7942,N_7888);
nand U8342 (N_8342,N_7124,N_7525);
nand U8343 (N_8343,N_7467,N_7032);
and U8344 (N_8344,N_7580,N_7318);
and U8345 (N_8345,N_7268,N_7431);
xnor U8346 (N_8346,N_7215,N_7709);
nor U8347 (N_8347,N_7144,N_7895);
nand U8348 (N_8348,N_7779,N_7326);
nor U8349 (N_8349,N_7786,N_7780);
or U8350 (N_8350,N_7871,N_7804);
nor U8351 (N_8351,N_7349,N_7848);
and U8352 (N_8352,N_7017,N_7328);
nand U8353 (N_8353,N_7953,N_7101);
nor U8354 (N_8354,N_7256,N_7896);
nand U8355 (N_8355,N_7232,N_7614);
and U8356 (N_8356,N_7317,N_7108);
nand U8357 (N_8357,N_7543,N_7199);
nand U8358 (N_8358,N_7443,N_7045);
nand U8359 (N_8359,N_7325,N_7971);
or U8360 (N_8360,N_7827,N_7653);
and U8361 (N_8361,N_7951,N_7096);
xor U8362 (N_8362,N_7970,N_7553);
nand U8363 (N_8363,N_7677,N_7729);
or U8364 (N_8364,N_7734,N_7147);
or U8365 (N_8365,N_7051,N_7112);
nor U8366 (N_8366,N_7244,N_7044);
xor U8367 (N_8367,N_7821,N_7181);
nor U8368 (N_8368,N_7302,N_7602);
and U8369 (N_8369,N_7995,N_7384);
and U8370 (N_8370,N_7930,N_7980);
nand U8371 (N_8371,N_7041,N_7402);
xnor U8372 (N_8372,N_7606,N_7190);
nor U8373 (N_8373,N_7425,N_7916);
nand U8374 (N_8374,N_7569,N_7358);
nand U8375 (N_8375,N_7629,N_7352);
and U8376 (N_8376,N_7814,N_7968);
or U8377 (N_8377,N_7599,N_7918);
xnor U8378 (N_8378,N_7605,N_7844);
nand U8379 (N_8379,N_7476,N_7588);
nor U8380 (N_8380,N_7607,N_7490);
nor U8381 (N_8381,N_7461,N_7197);
xor U8382 (N_8382,N_7394,N_7338);
nand U8383 (N_8383,N_7559,N_7254);
and U8384 (N_8384,N_7806,N_7206);
xor U8385 (N_8385,N_7136,N_7994);
nor U8386 (N_8386,N_7627,N_7568);
nor U8387 (N_8387,N_7372,N_7504);
xnor U8388 (N_8388,N_7085,N_7332);
xnor U8389 (N_8389,N_7403,N_7723);
or U8390 (N_8390,N_7562,N_7713);
xor U8391 (N_8391,N_7303,N_7282);
nand U8392 (N_8392,N_7892,N_7068);
nand U8393 (N_8393,N_7154,N_7829);
or U8394 (N_8394,N_7114,N_7087);
and U8395 (N_8395,N_7341,N_7439);
or U8396 (N_8396,N_7551,N_7819);
and U8397 (N_8397,N_7292,N_7131);
or U8398 (N_8398,N_7012,N_7134);
nor U8399 (N_8399,N_7654,N_7658);
xnor U8400 (N_8400,N_7672,N_7276);
and U8401 (N_8401,N_7155,N_7623);
xnor U8402 (N_8402,N_7216,N_7593);
xor U8403 (N_8403,N_7070,N_7050);
and U8404 (N_8404,N_7137,N_7459);
and U8405 (N_8405,N_7280,N_7516);
or U8406 (N_8406,N_7031,N_7502);
nand U8407 (N_8407,N_7843,N_7920);
and U8408 (N_8408,N_7212,N_7269);
xnor U8409 (N_8409,N_7783,N_7237);
xnor U8410 (N_8410,N_7006,N_7496);
xnor U8411 (N_8411,N_7015,N_7116);
nand U8412 (N_8412,N_7163,N_7079);
nand U8413 (N_8413,N_7132,N_7724);
nand U8414 (N_8414,N_7161,N_7753);
nor U8415 (N_8415,N_7684,N_7722);
xnor U8416 (N_8416,N_7233,N_7373);
or U8417 (N_8417,N_7289,N_7529);
xor U8418 (N_8418,N_7695,N_7546);
nor U8419 (N_8419,N_7084,N_7344);
xnor U8420 (N_8420,N_7777,N_7428);
nor U8421 (N_8421,N_7334,N_7039);
and U8422 (N_8422,N_7259,N_7900);
and U8423 (N_8423,N_7883,N_7577);
or U8424 (N_8424,N_7287,N_7932);
and U8425 (N_8425,N_7637,N_7135);
nand U8426 (N_8426,N_7463,N_7429);
and U8427 (N_8427,N_7911,N_7512);
or U8428 (N_8428,N_7937,N_7795);
and U8429 (N_8429,N_7625,N_7383);
and U8430 (N_8430,N_7764,N_7122);
xnor U8431 (N_8431,N_7407,N_7782);
and U8432 (N_8432,N_7495,N_7221);
nand U8433 (N_8433,N_7624,N_7564);
nand U8434 (N_8434,N_7946,N_7903);
or U8435 (N_8435,N_7758,N_7674);
xor U8436 (N_8436,N_7613,N_7343);
nand U8437 (N_8437,N_7333,N_7027);
or U8438 (N_8438,N_7381,N_7194);
and U8439 (N_8439,N_7401,N_7807);
or U8440 (N_8440,N_7549,N_7246);
nor U8441 (N_8441,N_7894,N_7555);
and U8442 (N_8442,N_7869,N_7270);
nor U8443 (N_8443,N_7721,N_7314);
nand U8444 (N_8444,N_7115,N_7277);
xnor U8445 (N_8445,N_7386,N_7889);
or U8446 (N_8446,N_7387,N_7891);
or U8447 (N_8447,N_7841,N_7919);
nand U8448 (N_8448,N_7160,N_7977);
and U8449 (N_8449,N_7091,N_7966);
nor U8450 (N_8450,N_7742,N_7451);
nor U8451 (N_8451,N_7582,N_7952);
nor U8452 (N_8452,N_7604,N_7826);
nand U8453 (N_8453,N_7097,N_7524);
xnor U8454 (N_8454,N_7845,N_7099);
xor U8455 (N_8455,N_7348,N_7418);
nand U8456 (N_8456,N_7854,N_7437);
or U8457 (N_8457,N_7727,N_7472);
and U8458 (N_8458,N_7227,N_7671);
xor U8459 (N_8459,N_7435,N_7960);
nand U8460 (N_8460,N_7146,N_7042);
xnor U8461 (N_8461,N_7575,N_7258);
and U8462 (N_8462,N_7239,N_7886);
or U8463 (N_8463,N_7813,N_7438);
or U8464 (N_8464,N_7164,N_7090);
nand U8465 (N_8465,N_7728,N_7836);
nor U8466 (N_8466,N_7498,N_7656);
nand U8467 (N_8467,N_7608,N_7291);
nor U8468 (N_8468,N_7765,N_7248);
xor U8469 (N_8469,N_7744,N_7789);
and U8470 (N_8470,N_7925,N_7893);
xnor U8471 (N_8471,N_7648,N_7857);
xnor U8472 (N_8472,N_7803,N_7271);
and U8473 (N_8473,N_7001,N_7148);
or U8474 (N_8474,N_7355,N_7284);
and U8475 (N_8475,N_7743,N_7948);
xor U8476 (N_8476,N_7113,N_7537);
nand U8477 (N_8477,N_7801,N_7356);
xnor U8478 (N_8478,N_7574,N_7471);
nand U8479 (N_8479,N_7022,N_7668);
nand U8480 (N_8480,N_7772,N_7576);
xnor U8481 (N_8481,N_7316,N_7669);
or U8482 (N_8482,N_7620,N_7026);
xor U8483 (N_8483,N_7413,N_7839);
xnor U8484 (N_8484,N_7694,N_7321);
xor U8485 (N_8485,N_7040,N_7494);
nor U8486 (N_8486,N_7336,N_7638);
nand U8487 (N_8487,N_7720,N_7563);
nand U8488 (N_8488,N_7736,N_7240);
nand U8489 (N_8489,N_7307,N_7346);
nand U8490 (N_8490,N_7214,N_7609);
xor U8491 (N_8491,N_7520,N_7452);
or U8492 (N_8492,N_7166,N_7700);
or U8493 (N_8493,N_7098,N_7354);
xnor U8494 (N_8494,N_7200,N_7832);
and U8495 (N_8495,N_7794,N_7185);
xor U8496 (N_8496,N_7375,N_7198);
xnor U8497 (N_8497,N_7220,N_7388);
and U8498 (N_8498,N_7110,N_7019);
or U8499 (N_8499,N_7621,N_7003);
nor U8500 (N_8500,N_7324,N_7675);
nor U8501 (N_8501,N_7604,N_7895);
or U8502 (N_8502,N_7786,N_7316);
nand U8503 (N_8503,N_7947,N_7835);
xor U8504 (N_8504,N_7181,N_7325);
or U8505 (N_8505,N_7068,N_7972);
xnor U8506 (N_8506,N_7909,N_7762);
nand U8507 (N_8507,N_7099,N_7306);
nand U8508 (N_8508,N_7466,N_7328);
nor U8509 (N_8509,N_7106,N_7332);
nand U8510 (N_8510,N_7469,N_7263);
nor U8511 (N_8511,N_7039,N_7233);
xnor U8512 (N_8512,N_7199,N_7738);
or U8513 (N_8513,N_7888,N_7487);
and U8514 (N_8514,N_7917,N_7510);
xor U8515 (N_8515,N_7679,N_7394);
or U8516 (N_8516,N_7283,N_7746);
nor U8517 (N_8517,N_7284,N_7015);
nand U8518 (N_8518,N_7008,N_7214);
xor U8519 (N_8519,N_7647,N_7861);
and U8520 (N_8520,N_7179,N_7877);
xor U8521 (N_8521,N_7911,N_7689);
nand U8522 (N_8522,N_7824,N_7120);
and U8523 (N_8523,N_7684,N_7927);
xor U8524 (N_8524,N_7997,N_7026);
nand U8525 (N_8525,N_7354,N_7207);
or U8526 (N_8526,N_7922,N_7107);
or U8527 (N_8527,N_7289,N_7716);
and U8528 (N_8528,N_7158,N_7822);
and U8529 (N_8529,N_7343,N_7410);
xnor U8530 (N_8530,N_7806,N_7198);
and U8531 (N_8531,N_7643,N_7647);
xor U8532 (N_8532,N_7377,N_7834);
nand U8533 (N_8533,N_7662,N_7065);
and U8534 (N_8534,N_7129,N_7958);
or U8535 (N_8535,N_7866,N_7626);
xor U8536 (N_8536,N_7569,N_7728);
nand U8537 (N_8537,N_7817,N_7314);
or U8538 (N_8538,N_7681,N_7562);
nor U8539 (N_8539,N_7328,N_7731);
and U8540 (N_8540,N_7865,N_7852);
and U8541 (N_8541,N_7756,N_7993);
nand U8542 (N_8542,N_7842,N_7422);
and U8543 (N_8543,N_7814,N_7732);
xnor U8544 (N_8544,N_7053,N_7145);
or U8545 (N_8545,N_7031,N_7347);
and U8546 (N_8546,N_7223,N_7777);
nor U8547 (N_8547,N_7609,N_7662);
and U8548 (N_8548,N_7378,N_7029);
nand U8549 (N_8549,N_7669,N_7131);
or U8550 (N_8550,N_7477,N_7882);
nor U8551 (N_8551,N_7541,N_7467);
nand U8552 (N_8552,N_7285,N_7692);
or U8553 (N_8553,N_7078,N_7860);
nor U8554 (N_8554,N_7482,N_7089);
nor U8555 (N_8555,N_7638,N_7853);
xor U8556 (N_8556,N_7389,N_7900);
or U8557 (N_8557,N_7127,N_7012);
nand U8558 (N_8558,N_7924,N_7276);
and U8559 (N_8559,N_7421,N_7117);
xor U8560 (N_8560,N_7781,N_7842);
or U8561 (N_8561,N_7335,N_7056);
nor U8562 (N_8562,N_7894,N_7095);
or U8563 (N_8563,N_7837,N_7460);
nand U8564 (N_8564,N_7871,N_7560);
and U8565 (N_8565,N_7968,N_7245);
nor U8566 (N_8566,N_7934,N_7575);
or U8567 (N_8567,N_7441,N_7823);
and U8568 (N_8568,N_7686,N_7660);
and U8569 (N_8569,N_7850,N_7858);
nand U8570 (N_8570,N_7910,N_7464);
xnor U8571 (N_8571,N_7788,N_7729);
and U8572 (N_8572,N_7822,N_7193);
or U8573 (N_8573,N_7079,N_7273);
and U8574 (N_8574,N_7813,N_7790);
and U8575 (N_8575,N_7612,N_7893);
nor U8576 (N_8576,N_7362,N_7883);
or U8577 (N_8577,N_7572,N_7341);
or U8578 (N_8578,N_7024,N_7193);
nor U8579 (N_8579,N_7912,N_7525);
and U8580 (N_8580,N_7979,N_7837);
and U8581 (N_8581,N_7951,N_7380);
xnor U8582 (N_8582,N_7378,N_7645);
and U8583 (N_8583,N_7413,N_7094);
or U8584 (N_8584,N_7792,N_7545);
and U8585 (N_8585,N_7975,N_7369);
nor U8586 (N_8586,N_7173,N_7569);
nand U8587 (N_8587,N_7604,N_7187);
or U8588 (N_8588,N_7309,N_7683);
nand U8589 (N_8589,N_7985,N_7648);
nor U8590 (N_8590,N_7580,N_7751);
nand U8591 (N_8591,N_7726,N_7995);
nand U8592 (N_8592,N_7412,N_7940);
nand U8593 (N_8593,N_7239,N_7094);
or U8594 (N_8594,N_7723,N_7414);
and U8595 (N_8595,N_7169,N_7220);
nor U8596 (N_8596,N_7160,N_7828);
xor U8597 (N_8597,N_7570,N_7262);
xor U8598 (N_8598,N_7649,N_7807);
nor U8599 (N_8599,N_7772,N_7476);
nor U8600 (N_8600,N_7844,N_7575);
or U8601 (N_8601,N_7395,N_7319);
nand U8602 (N_8602,N_7215,N_7401);
xor U8603 (N_8603,N_7449,N_7649);
xnor U8604 (N_8604,N_7729,N_7122);
xor U8605 (N_8605,N_7756,N_7435);
nor U8606 (N_8606,N_7045,N_7236);
or U8607 (N_8607,N_7814,N_7007);
nand U8608 (N_8608,N_7799,N_7285);
nor U8609 (N_8609,N_7760,N_7711);
or U8610 (N_8610,N_7446,N_7156);
xor U8611 (N_8611,N_7501,N_7282);
or U8612 (N_8612,N_7575,N_7336);
nor U8613 (N_8613,N_7933,N_7613);
and U8614 (N_8614,N_7030,N_7357);
nand U8615 (N_8615,N_7308,N_7572);
xnor U8616 (N_8616,N_7394,N_7508);
or U8617 (N_8617,N_7135,N_7396);
or U8618 (N_8618,N_7893,N_7577);
xnor U8619 (N_8619,N_7933,N_7686);
nand U8620 (N_8620,N_7590,N_7752);
nand U8621 (N_8621,N_7768,N_7585);
nand U8622 (N_8622,N_7595,N_7605);
xnor U8623 (N_8623,N_7946,N_7675);
or U8624 (N_8624,N_7653,N_7032);
nor U8625 (N_8625,N_7520,N_7980);
nand U8626 (N_8626,N_7086,N_7738);
nand U8627 (N_8627,N_7659,N_7347);
nand U8628 (N_8628,N_7106,N_7053);
nor U8629 (N_8629,N_7184,N_7948);
nor U8630 (N_8630,N_7679,N_7629);
nand U8631 (N_8631,N_7098,N_7647);
and U8632 (N_8632,N_7512,N_7923);
nand U8633 (N_8633,N_7739,N_7115);
xnor U8634 (N_8634,N_7856,N_7946);
or U8635 (N_8635,N_7331,N_7636);
xor U8636 (N_8636,N_7876,N_7509);
or U8637 (N_8637,N_7337,N_7477);
nand U8638 (N_8638,N_7779,N_7191);
or U8639 (N_8639,N_7185,N_7832);
or U8640 (N_8640,N_7481,N_7134);
and U8641 (N_8641,N_7888,N_7822);
nand U8642 (N_8642,N_7972,N_7899);
nand U8643 (N_8643,N_7035,N_7537);
nor U8644 (N_8644,N_7829,N_7254);
and U8645 (N_8645,N_7144,N_7456);
xnor U8646 (N_8646,N_7013,N_7271);
or U8647 (N_8647,N_7532,N_7080);
or U8648 (N_8648,N_7134,N_7240);
and U8649 (N_8649,N_7447,N_7345);
nand U8650 (N_8650,N_7889,N_7366);
nand U8651 (N_8651,N_7628,N_7018);
or U8652 (N_8652,N_7376,N_7674);
nand U8653 (N_8653,N_7912,N_7232);
xnor U8654 (N_8654,N_7600,N_7286);
nor U8655 (N_8655,N_7026,N_7758);
nor U8656 (N_8656,N_7000,N_7172);
and U8657 (N_8657,N_7422,N_7047);
nand U8658 (N_8658,N_7005,N_7542);
nor U8659 (N_8659,N_7733,N_7427);
or U8660 (N_8660,N_7304,N_7379);
nor U8661 (N_8661,N_7871,N_7169);
or U8662 (N_8662,N_7806,N_7480);
nor U8663 (N_8663,N_7846,N_7668);
xor U8664 (N_8664,N_7877,N_7769);
xor U8665 (N_8665,N_7084,N_7717);
and U8666 (N_8666,N_7669,N_7970);
xor U8667 (N_8667,N_7222,N_7397);
or U8668 (N_8668,N_7769,N_7044);
nand U8669 (N_8669,N_7157,N_7932);
xnor U8670 (N_8670,N_7012,N_7904);
or U8671 (N_8671,N_7719,N_7593);
nor U8672 (N_8672,N_7639,N_7905);
nor U8673 (N_8673,N_7798,N_7492);
xor U8674 (N_8674,N_7650,N_7865);
or U8675 (N_8675,N_7561,N_7120);
and U8676 (N_8676,N_7398,N_7712);
or U8677 (N_8677,N_7449,N_7022);
nor U8678 (N_8678,N_7141,N_7233);
xnor U8679 (N_8679,N_7344,N_7978);
nand U8680 (N_8680,N_7936,N_7989);
nand U8681 (N_8681,N_7973,N_7060);
and U8682 (N_8682,N_7489,N_7158);
or U8683 (N_8683,N_7162,N_7734);
and U8684 (N_8684,N_7616,N_7406);
xor U8685 (N_8685,N_7465,N_7516);
nand U8686 (N_8686,N_7379,N_7596);
nor U8687 (N_8687,N_7472,N_7276);
xnor U8688 (N_8688,N_7705,N_7162);
nand U8689 (N_8689,N_7403,N_7495);
nand U8690 (N_8690,N_7099,N_7768);
xor U8691 (N_8691,N_7972,N_7329);
or U8692 (N_8692,N_7102,N_7931);
or U8693 (N_8693,N_7032,N_7914);
nand U8694 (N_8694,N_7758,N_7110);
or U8695 (N_8695,N_7704,N_7482);
xor U8696 (N_8696,N_7698,N_7442);
or U8697 (N_8697,N_7927,N_7411);
and U8698 (N_8698,N_7442,N_7137);
nand U8699 (N_8699,N_7917,N_7597);
nor U8700 (N_8700,N_7240,N_7687);
or U8701 (N_8701,N_7215,N_7907);
nor U8702 (N_8702,N_7478,N_7172);
nor U8703 (N_8703,N_7775,N_7322);
or U8704 (N_8704,N_7343,N_7543);
nor U8705 (N_8705,N_7798,N_7195);
nor U8706 (N_8706,N_7588,N_7133);
nor U8707 (N_8707,N_7507,N_7442);
nand U8708 (N_8708,N_7591,N_7642);
nand U8709 (N_8709,N_7052,N_7992);
and U8710 (N_8710,N_7108,N_7225);
xor U8711 (N_8711,N_7712,N_7151);
nand U8712 (N_8712,N_7663,N_7136);
xnor U8713 (N_8713,N_7275,N_7380);
xnor U8714 (N_8714,N_7642,N_7806);
nor U8715 (N_8715,N_7093,N_7795);
and U8716 (N_8716,N_7173,N_7822);
and U8717 (N_8717,N_7171,N_7785);
nor U8718 (N_8718,N_7087,N_7918);
nand U8719 (N_8719,N_7245,N_7692);
xnor U8720 (N_8720,N_7018,N_7017);
xnor U8721 (N_8721,N_7999,N_7500);
or U8722 (N_8722,N_7461,N_7699);
nand U8723 (N_8723,N_7161,N_7520);
xor U8724 (N_8724,N_7916,N_7066);
nand U8725 (N_8725,N_7430,N_7994);
or U8726 (N_8726,N_7693,N_7032);
nand U8727 (N_8727,N_7991,N_7128);
and U8728 (N_8728,N_7398,N_7413);
or U8729 (N_8729,N_7411,N_7118);
and U8730 (N_8730,N_7374,N_7678);
xnor U8731 (N_8731,N_7641,N_7083);
nand U8732 (N_8732,N_7515,N_7125);
xor U8733 (N_8733,N_7554,N_7607);
nor U8734 (N_8734,N_7697,N_7241);
nor U8735 (N_8735,N_7158,N_7008);
nand U8736 (N_8736,N_7907,N_7470);
and U8737 (N_8737,N_7281,N_7342);
or U8738 (N_8738,N_7580,N_7232);
xor U8739 (N_8739,N_7602,N_7656);
nor U8740 (N_8740,N_7096,N_7619);
xnor U8741 (N_8741,N_7001,N_7280);
nor U8742 (N_8742,N_7020,N_7402);
and U8743 (N_8743,N_7524,N_7794);
or U8744 (N_8744,N_7448,N_7349);
and U8745 (N_8745,N_7543,N_7592);
nor U8746 (N_8746,N_7522,N_7912);
nor U8747 (N_8747,N_7693,N_7236);
nor U8748 (N_8748,N_7588,N_7810);
nor U8749 (N_8749,N_7528,N_7027);
and U8750 (N_8750,N_7411,N_7944);
nand U8751 (N_8751,N_7377,N_7511);
or U8752 (N_8752,N_7775,N_7115);
and U8753 (N_8753,N_7781,N_7798);
nand U8754 (N_8754,N_7117,N_7579);
and U8755 (N_8755,N_7897,N_7825);
xor U8756 (N_8756,N_7038,N_7048);
nor U8757 (N_8757,N_7478,N_7601);
nand U8758 (N_8758,N_7386,N_7185);
nand U8759 (N_8759,N_7869,N_7073);
nand U8760 (N_8760,N_7374,N_7265);
or U8761 (N_8761,N_7278,N_7543);
nor U8762 (N_8762,N_7211,N_7217);
and U8763 (N_8763,N_7043,N_7182);
or U8764 (N_8764,N_7995,N_7674);
and U8765 (N_8765,N_7978,N_7317);
nor U8766 (N_8766,N_7525,N_7425);
xor U8767 (N_8767,N_7251,N_7260);
or U8768 (N_8768,N_7784,N_7174);
xor U8769 (N_8769,N_7271,N_7509);
and U8770 (N_8770,N_7357,N_7609);
or U8771 (N_8771,N_7648,N_7144);
and U8772 (N_8772,N_7352,N_7961);
xor U8773 (N_8773,N_7713,N_7131);
xor U8774 (N_8774,N_7283,N_7940);
xor U8775 (N_8775,N_7498,N_7355);
nand U8776 (N_8776,N_7844,N_7400);
and U8777 (N_8777,N_7157,N_7206);
xnor U8778 (N_8778,N_7833,N_7384);
nand U8779 (N_8779,N_7947,N_7577);
xor U8780 (N_8780,N_7617,N_7634);
nor U8781 (N_8781,N_7958,N_7694);
or U8782 (N_8782,N_7605,N_7066);
nand U8783 (N_8783,N_7531,N_7476);
and U8784 (N_8784,N_7632,N_7293);
xor U8785 (N_8785,N_7382,N_7927);
and U8786 (N_8786,N_7743,N_7373);
or U8787 (N_8787,N_7830,N_7676);
xor U8788 (N_8788,N_7679,N_7853);
xor U8789 (N_8789,N_7699,N_7122);
nor U8790 (N_8790,N_7813,N_7223);
nor U8791 (N_8791,N_7794,N_7040);
xnor U8792 (N_8792,N_7710,N_7942);
and U8793 (N_8793,N_7792,N_7616);
or U8794 (N_8794,N_7307,N_7984);
xnor U8795 (N_8795,N_7279,N_7149);
and U8796 (N_8796,N_7945,N_7055);
xnor U8797 (N_8797,N_7607,N_7227);
nand U8798 (N_8798,N_7151,N_7908);
or U8799 (N_8799,N_7579,N_7760);
nor U8800 (N_8800,N_7417,N_7290);
nand U8801 (N_8801,N_7805,N_7283);
xnor U8802 (N_8802,N_7219,N_7069);
xnor U8803 (N_8803,N_7847,N_7947);
or U8804 (N_8804,N_7694,N_7446);
and U8805 (N_8805,N_7571,N_7753);
nand U8806 (N_8806,N_7856,N_7006);
nor U8807 (N_8807,N_7685,N_7678);
nor U8808 (N_8808,N_7635,N_7459);
nand U8809 (N_8809,N_7120,N_7817);
or U8810 (N_8810,N_7566,N_7348);
nor U8811 (N_8811,N_7444,N_7070);
or U8812 (N_8812,N_7661,N_7084);
nor U8813 (N_8813,N_7866,N_7463);
and U8814 (N_8814,N_7797,N_7746);
xnor U8815 (N_8815,N_7498,N_7178);
nor U8816 (N_8816,N_7253,N_7673);
xor U8817 (N_8817,N_7918,N_7876);
nand U8818 (N_8818,N_7312,N_7645);
nand U8819 (N_8819,N_7312,N_7188);
and U8820 (N_8820,N_7594,N_7280);
and U8821 (N_8821,N_7634,N_7739);
nand U8822 (N_8822,N_7455,N_7194);
xnor U8823 (N_8823,N_7595,N_7929);
and U8824 (N_8824,N_7524,N_7051);
nor U8825 (N_8825,N_7820,N_7762);
nor U8826 (N_8826,N_7342,N_7363);
nor U8827 (N_8827,N_7183,N_7967);
xnor U8828 (N_8828,N_7777,N_7484);
xnor U8829 (N_8829,N_7200,N_7045);
and U8830 (N_8830,N_7329,N_7135);
nor U8831 (N_8831,N_7482,N_7259);
nand U8832 (N_8832,N_7382,N_7911);
xor U8833 (N_8833,N_7739,N_7057);
xor U8834 (N_8834,N_7467,N_7330);
and U8835 (N_8835,N_7683,N_7706);
xnor U8836 (N_8836,N_7834,N_7910);
nand U8837 (N_8837,N_7648,N_7193);
nand U8838 (N_8838,N_7369,N_7499);
xnor U8839 (N_8839,N_7322,N_7856);
and U8840 (N_8840,N_7808,N_7424);
or U8841 (N_8841,N_7374,N_7531);
nor U8842 (N_8842,N_7091,N_7863);
or U8843 (N_8843,N_7616,N_7903);
nand U8844 (N_8844,N_7218,N_7022);
nand U8845 (N_8845,N_7719,N_7499);
and U8846 (N_8846,N_7071,N_7155);
nand U8847 (N_8847,N_7652,N_7207);
xor U8848 (N_8848,N_7476,N_7925);
xor U8849 (N_8849,N_7638,N_7412);
and U8850 (N_8850,N_7800,N_7872);
nand U8851 (N_8851,N_7467,N_7121);
nand U8852 (N_8852,N_7106,N_7692);
nand U8853 (N_8853,N_7103,N_7132);
xnor U8854 (N_8854,N_7044,N_7619);
nor U8855 (N_8855,N_7353,N_7129);
or U8856 (N_8856,N_7684,N_7815);
nor U8857 (N_8857,N_7200,N_7584);
nand U8858 (N_8858,N_7698,N_7460);
nand U8859 (N_8859,N_7199,N_7937);
nor U8860 (N_8860,N_7607,N_7089);
nand U8861 (N_8861,N_7004,N_7671);
and U8862 (N_8862,N_7412,N_7040);
and U8863 (N_8863,N_7347,N_7195);
or U8864 (N_8864,N_7020,N_7144);
nand U8865 (N_8865,N_7048,N_7152);
and U8866 (N_8866,N_7780,N_7064);
or U8867 (N_8867,N_7072,N_7427);
or U8868 (N_8868,N_7355,N_7132);
xor U8869 (N_8869,N_7240,N_7236);
nor U8870 (N_8870,N_7210,N_7825);
or U8871 (N_8871,N_7304,N_7841);
xnor U8872 (N_8872,N_7869,N_7016);
or U8873 (N_8873,N_7011,N_7601);
nor U8874 (N_8874,N_7050,N_7232);
and U8875 (N_8875,N_7938,N_7094);
and U8876 (N_8876,N_7588,N_7270);
nor U8877 (N_8877,N_7925,N_7402);
nor U8878 (N_8878,N_7663,N_7183);
and U8879 (N_8879,N_7696,N_7983);
nand U8880 (N_8880,N_7160,N_7838);
or U8881 (N_8881,N_7694,N_7549);
nand U8882 (N_8882,N_7624,N_7687);
nor U8883 (N_8883,N_7414,N_7135);
or U8884 (N_8884,N_7265,N_7595);
or U8885 (N_8885,N_7232,N_7161);
xnor U8886 (N_8886,N_7857,N_7441);
and U8887 (N_8887,N_7256,N_7119);
nand U8888 (N_8888,N_7495,N_7900);
nand U8889 (N_8889,N_7839,N_7932);
and U8890 (N_8890,N_7922,N_7277);
xor U8891 (N_8891,N_7314,N_7419);
xor U8892 (N_8892,N_7024,N_7137);
xnor U8893 (N_8893,N_7040,N_7366);
nand U8894 (N_8894,N_7706,N_7009);
nand U8895 (N_8895,N_7135,N_7702);
nand U8896 (N_8896,N_7967,N_7519);
xnor U8897 (N_8897,N_7102,N_7704);
nor U8898 (N_8898,N_7869,N_7681);
or U8899 (N_8899,N_7346,N_7018);
and U8900 (N_8900,N_7529,N_7501);
xor U8901 (N_8901,N_7988,N_7275);
nand U8902 (N_8902,N_7359,N_7792);
and U8903 (N_8903,N_7523,N_7816);
xnor U8904 (N_8904,N_7685,N_7776);
or U8905 (N_8905,N_7034,N_7401);
and U8906 (N_8906,N_7136,N_7631);
or U8907 (N_8907,N_7795,N_7702);
nand U8908 (N_8908,N_7876,N_7077);
xnor U8909 (N_8909,N_7192,N_7591);
xor U8910 (N_8910,N_7422,N_7949);
xor U8911 (N_8911,N_7203,N_7643);
or U8912 (N_8912,N_7161,N_7300);
and U8913 (N_8913,N_7846,N_7467);
xnor U8914 (N_8914,N_7533,N_7592);
and U8915 (N_8915,N_7456,N_7885);
or U8916 (N_8916,N_7383,N_7421);
and U8917 (N_8917,N_7134,N_7513);
or U8918 (N_8918,N_7280,N_7660);
nand U8919 (N_8919,N_7233,N_7558);
or U8920 (N_8920,N_7827,N_7073);
nor U8921 (N_8921,N_7964,N_7456);
or U8922 (N_8922,N_7995,N_7681);
nor U8923 (N_8923,N_7722,N_7967);
nor U8924 (N_8924,N_7527,N_7887);
xnor U8925 (N_8925,N_7665,N_7228);
xor U8926 (N_8926,N_7673,N_7607);
or U8927 (N_8927,N_7822,N_7687);
and U8928 (N_8928,N_7803,N_7855);
and U8929 (N_8929,N_7026,N_7372);
or U8930 (N_8930,N_7882,N_7563);
nor U8931 (N_8931,N_7402,N_7779);
and U8932 (N_8932,N_7475,N_7413);
or U8933 (N_8933,N_7286,N_7638);
nor U8934 (N_8934,N_7690,N_7861);
or U8935 (N_8935,N_7200,N_7634);
xnor U8936 (N_8936,N_7060,N_7273);
nor U8937 (N_8937,N_7523,N_7527);
or U8938 (N_8938,N_7650,N_7106);
xnor U8939 (N_8939,N_7534,N_7903);
nor U8940 (N_8940,N_7021,N_7826);
nand U8941 (N_8941,N_7846,N_7725);
or U8942 (N_8942,N_7775,N_7009);
xor U8943 (N_8943,N_7689,N_7078);
nor U8944 (N_8944,N_7647,N_7543);
nand U8945 (N_8945,N_7946,N_7692);
and U8946 (N_8946,N_7817,N_7636);
xnor U8947 (N_8947,N_7047,N_7318);
nand U8948 (N_8948,N_7165,N_7679);
or U8949 (N_8949,N_7424,N_7327);
and U8950 (N_8950,N_7663,N_7716);
or U8951 (N_8951,N_7130,N_7316);
nand U8952 (N_8952,N_7546,N_7415);
or U8953 (N_8953,N_7896,N_7103);
nor U8954 (N_8954,N_7801,N_7312);
nand U8955 (N_8955,N_7609,N_7263);
nand U8956 (N_8956,N_7320,N_7892);
or U8957 (N_8957,N_7007,N_7456);
nor U8958 (N_8958,N_7413,N_7661);
or U8959 (N_8959,N_7359,N_7422);
nand U8960 (N_8960,N_7743,N_7035);
or U8961 (N_8961,N_7551,N_7680);
nor U8962 (N_8962,N_7672,N_7909);
nor U8963 (N_8963,N_7894,N_7917);
nand U8964 (N_8964,N_7041,N_7662);
xnor U8965 (N_8965,N_7459,N_7458);
and U8966 (N_8966,N_7318,N_7107);
and U8967 (N_8967,N_7646,N_7365);
xnor U8968 (N_8968,N_7710,N_7086);
and U8969 (N_8969,N_7634,N_7232);
nand U8970 (N_8970,N_7405,N_7063);
and U8971 (N_8971,N_7343,N_7985);
and U8972 (N_8972,N_7045,N_7736);
and U8973 (N_8973,N_7752,N_7928);
nand U8974 (N_8974,N_7859,N_7792);
xor U8975 (N_8975,N_7972,N_7950);
and U8976 (N_8976,N_7226,N_7866);
or U8977 (N_8977,N_7136,N_7968);
and U8978 (N_8978,N_7487,N_7884);
or U8979 (N_8979,N_7958,N_7833);
xnor U8980 (N_8980,N_7783,N_7188);
nand U8981 (N_8981,N_7741,N_7720);
nor U8982 (N_8982,N_7816,N_7459);
or U8983 (N_8983,N_7309,N_7164);
xor U8984 (N_8984,N_7767,N_7206);
xnor U8985 (N_8985,N_7372,N_7421);
and U8986 (N_8986,N_7485,N_7048);
and U8987 (N_8987,N_7473,N_7453);
or U8988 (N_8988,N_7963,N_7985);
and U8989 (N_8989,N_7118,N_7695);
xor U8990 (N_8990,N_7731,N_7636);
and U8991 (N_8991,N_7438,N_7811);
nand U8992 (N_8992,N_7026,N_7580);
nor U8993 (N_8993,N_7982,N_7357);
and U8994 (N_8994,N_7348,N_7559);
or U8995 (N_8995,N_7071,N_7705);
or U8996 (N_8996,N_7984,N_7434);
xnor U8997 (N_8997,N_7972,N_7586);
nand U8998 (N_8998,N_7197,N_7703);
nor U8999 (N_8999,N_7615,N_7249);
or U9000 (N_9000,N_8400,N_8313);
nand U9001 (N_9001,N_8492,N_8139);
nor U9002 (N_9002,N_8303,N_8582);
nand U9003 (N_9003,N_8832,N_8002);
nor U9004 (N_9004,N_8914,N_8606);
and U9005 (N_9005,N_8770,N_8245);
or U9006 (N_9006,N_8676,N_8273);
nand U9007 (N_9007,N_8939,N_8306);
and U9008 (N_9008,N_8763,N_8120);
nand U9009 (N_9009,N_8357,N_8250);
xor U9010 (N_9010,N_8370,N_8550);
nand U9011 (N_9011,N_8869,N_8500);
nand U9012 (N_9012,N_8508,N_8957);
and U9013 (N_9013,N_8873,N_8092);
or U9014 (N_9014,N_8008,N_8575);
nand U9015 (N_9015,N_8523,N_8865);
and U9016 (N_9016,N_8056,N_8312);
or U9017 (N_9017,N_8542,N_8617);
and U9018 (N_9018,N_8178,N_8891);
nor U9019 (N_9019,N_8862,N_8408);
xor U9020 (N_9020,N_8997,N_8307);
and U9021 (N_9021,N_8905,N_8212);
nand U9022 (N_9022,N_8427,N_8177);
and U9023 (N_9023,N_8986,N_8554);
and U9024 (N_9024,N_8601,N_8126);
nor U9025 (N_9025,N_8634,N_8830);
or U9026 (N_9026,N_8387,N_8852);
xor U9027 (N_9027,N_8300,N_8052);
or U9028 (N_9028,N_8181,N_8931);
xor U9029 (N_9029,N_8261,N_8741);
nor U9030 (N_9030,N_8722,N_8467);
or U9031 (N_9031,N_8879,N_8156);
nand U9032 (N_9032,N_8125,N_8607);
and U9033 (N_9033,N_8291,N_8924);
xnor U9034 (N_9034,N_8683,N_8235);
and U9035 (N_9035,N_8505,N_8328);
nand U9036 (N_9036,N_8710,N_8790);
or U9037 (N_9037,N_8585,N_8149);
and U9038 (N_9038,N_8082,N_8968);
nor U9039 (N_9039,N_8541,N_8014);
nor U9040 (N_9040,N_8440,N_8006);
nor U9041 (N_9041,N_8119,N_8202);
and U9042 (N_9042,N_8208,N_8735);
and U9043 (N_9043,N_8123,N_8641);
nand U9044 (N_9044,N_8987,N_8749);
xnor U9045 (N_9045,N_8824,N_8209);
or U9046 (N_9046,N_8128,N_8108);
nand U9047 (N_9047,N_8112,N_8622);
or U9048 (N_9048,N_8376,N_8583);
and U9049 (N_9049,N_8875,N_8952);
or U9050 (N_9050,N_8906,N_8455);
xnor U9051 (N_9051,N_8154,N_8662);
nor U9052 (N_9052,N_8984,N_8979);
xor U9053 (N_9053,N_8761,N_8613);
nor U9054 (N_9054,N_8480,N_8724);
and U9055 (N_9055,N_8829,N_8766);
xnor U9056 (N_9056,N_8336,N_8342);
or U9057 (N_9057,N_8439,N_8731);
xor U9058 (N_9058,N_8949,N_8309);
and U9059 (N_9059,N_8220,N_8354);
nand U9060 (N_9060,N_8743,N_8451);
xnor U9061 (N_9061,N_8897,N_8791);
nor U9062 (N_9062,N_8061,N_8848);
xor U9063 (N_9063,N_8825,N_8765);
nand U9064 (N_9064,N_8925,N_8597);
nand U9065 (N_9065,N_8394,N_8780);
nor U9066 (N_9066,N_8927,N_8104);
nor U9067 (N_9067,N_8758,N_8134);
xnor U9068 (N_9068,N_8611,N_8109);
or U9069 (N_9069,N_8165,N_8549);
xor U9070 (N_9070,N_8027,N_8893);
xnor U9071 (N_9071,N_8544,N_8750);
xor U9072 (N_9072,N_8584,N_8371);
nand U9073 (N_9073,N_8563,N_8373);
or U9074 (N_9074,N_8753,N_8302);
xor U9075 (N_9075,N_8163,N_8754);
xor U9076 (N_9076,N_8147,N_8262);
xor U9077 (N_9077,N_8459,N_8518);
xnor U9078 (N_9078,N_8351,N_8067);
nor U9079 (N_9079,N_8643,N_8828);
nand U9080 (N_9080,N_8434,N_8093);
xor U9081 (N_9081,N_8624,N_8991);
nor U9082 (N_9082,N_8231,N_8880);
xnor U9083 (N_9083,N_8454,N_8921);
or U9084 (N_9084,N_8343,N_8918);
or U9085 (N_9085,N_8833,N_8422);
xnor U9086 (N_9086,N_8205,N_8332);
xor U9087 (N_9087,N_8680,N_8962);
xnor U9088 (N_9088,N_8771,N_8048);
and U9089 (N_9089,N_8269,N_8071);
nor U9090 (N_9090,N_8477,N_8647);
xor U9091 (N_9091,N_8864,N_8041);
and U9092 (N_9092,N_8928,N_8456);
or U9093 (N_9093,N_8000,N_8407);
or U9094 (N_9094,N_8548,N_8026);
or U9095 (N_9095,N_8981,N_8274);
xnor U9096 (N_9096,N_8238,N_8369);
or U9097 (N_9097,N_8276,N_8497);
nand U9098 (N_9098,N_8160,N_8232);
or U9099 (N_9099,N_8169,N_8805);
nor U9100 (N_9100,N_8755,N_8446);
or U9101 (N_9101,N_8364,N_8210);
xor U9102 (N_9102,N_8519,N_8756);
xor U9103 (N_9103,N_8520,N_8999);
and U9104 (N_9104,N_8267,N_8331);
nor U9105 (N_9105,N_8396,N_8815);
or U9106 (N_9106,N_8510,N_8916);
xor U9107 (N_9107,N_8857,N_8063);
xnor U9108 (N_9108,N_8608,N_8097);
xor U9109 (N_9109,N_8428,N_8083);
or U9110 (N_9110,N_8535,N_8907);
or U9111 (N_9111,N_8615,N_8671);
and U9112 (N_9112,N_8747,N_8404);
or U9113 (N_9113,N_8337,N_8389);
xnor U9114 (N_9114,N_8666,N_8385);
nand U9115 (N_9115,N_8806,N_8064);
xor U9116 (N_9116,N_8195,N_8431);
or U9117 (N_9117,N_8507,N_8118);
nand U9118 (N_9118,N_8689,N_8562);
and U9119 (N_9119,N_8863,N_8383);
nor U9120 (N_9120,N_8487,N_8340);
and U9121 (N_9121,N_8397,N_8580);
and U9122 (N_9122,N_8240,N_8764);
or U9123 (N_9123,N_8482,N_8329);
nand U9124 (N_9124,N_8684,N_8499);
or U9125 (N_9125,N_8708,N_8560);
xnor U9126 (N_9126,N_8531,N_8860);
or U9127 (N_9127,N_8416,N_8271);
and U9128 (N_9128,N_8589,N_8457);
or U9129 (N_9129,N_8961,N_8474);
and U9130 (N_9130,N_8567,N_8425);
nor U9131 (N_9131,N_8078,N_8890);
nor U9132 (N_9132,N_8511,N_8781);
xor U9133 (N_9133,N_8522,N_8760);
and U9134 (N_9134,N_8292,N_8596);
or U9135 (N_9135,N_8729,N_8651);
and U9136 (N_9136,N_8900,N_8066);
xor U9137 (N_9137,N_8105,N_8200);
nand U9138 (N_9138,N_8198,N_8776);
or U9139 (N_9139,N_8138,N_8317);
xor U9140 (N_9140,N_8035,N_8909);
or U9141 (N_9141,N_8490,N_8223);
and U9142 (N_9142,N_8024,N_8812);
nor U9143 (N_9143,N_8219,N_8712);
xnor U9144 (N_9144,N_8171,N_8222);
xor U9145 (N_9145,N_8659,N_8571);
nor U9146 (N_9146,N_8588,N_8516);
xnor U9147 (N_9147,N_8967,N_8032);
nor U9148 (N_9148,N_8076,N_8950);
xor U9149 (N_9149,N_8088,N_8665);
or U9150 (N_9150,N_8941,N_8784);
nor U9151 (N_9151,N_8029,N_8166);
and U9152 (N_9152,N_8556,N_8405);
nor U9153 (N_9153,N_8850,N_8144);
nand U9154 (N_9154,N_8287,N_8242);
xnor U9155 (N_9155,N_8578,N_8688);
xnor U9156 (N_9156,N_8971,N_8954);
nand U9157 (N_9157,N_8384,N_8996);
xor U9158 (N_9158,N_8311,N_8473);
nor U9159 (N_9159,N_8546,N_8218);
xnor U9160 (N_9160,N_8183,N_8895);
and U9161 (N_9161,N_8642,N_8573);
or U9162 (N_9162,N_8837,N_8819);
or U9163 (N_9163,N_8524,N_8868);
or U9164 (N_9164,N_8877,N_8377);
nor U9165 (N_9165,N_8707,N_8650);
nor U9166 (N_9166,N_8072,N_8491);
nand U9167 (N_9167,N_8243,N_8226);
and U9168 (N_9168,N_8060,N_8586);
nand U9169 (N_9169,N_8424,N_8324);
and U9170 (N_9170,N_8789,N_8813);
xor U9171 (N_9171,N_8362,N_8823);
nor U9172 (N_9172,N_8995,N_8039);
xnor U9173 (N_9173,N_8721,N_8009);
or U9174 (N_9174,N_8752,N_8983);
xor U9175 (N_9175,N_8536,N_8807);
and U9176 (N_9176,N_8687,N_8577);
or U9177 (N_9177,N_8881,N_8594);
nand U9178 (N_9178,N_8975,N_8561);
xnor U9179 (N_9179,N_8746,N_8839);
xnor U9180 (N_9180,N_8472,N_8265);
nor U9181 (N_9181,N_8512,N_8327);
xnor U9182 (N_9182,N_8803,N_8059);
nor U9183 (N_9183,N_8551,N_8559);
nor U9184 (N_9184,N_8378,N_8736);
nor U9185 (N_9185,N_8135,N_8055);
or U9186 (N_9186,N_8566,N_8898);
or U9187 (N_9187,N_8834,N_8237);
nor U9188 (N_9188,N_8442,N_8678);
or U9189 (N_9189,N_8911,N_8751);
xnor U9190 (N_9190,N_8934,N_8161);
nand U9191 (N_9191,N_8528,N_8192);
nand U9192 (N_9192,N_8587,N_8783);
xnor U9193 (N_9193,N_8019,N_8867);
nor U9194 (N_9194,N_8447,N_8841);
xor U9195 (N_9195,N_8234,N_8915);
or U9196 (N_9196,N_8185,N_8375);
and U9197 (N_9197,N_8363,N_8347);
nand U9198 (N_9198,N_8951,N_8669);
or U9199 (N_9199,N_8919,N_8395);
or U9200 (N_9200,N_8025,N_8013);
nand U9201 (N_9201,N_8290,N_8252);
nand U9202 (N_9202,N_8663,N_8976);
nand U9203 (N_9203,N_8233,N_8581);
and U9204 (N_9204,N_8127,N_8018);
or U9205 (N_9205,N_8334,N_8186);
nor U9206 (N_9206,N_8525,N_8441);
or U9207 (N_9207,N_8858,N_8640);
nand U9208 (N_9208,N_8162,N_8316);
xor U9209 (N_9209,N_8657,N_8846);
or U9210 (N_9210,N_8885,N_8638);
xor U9211 (N_9211,N_8325,N_8326);
nand U9212 (N_9212,N_8412,N_8576);
nand U9213 (N_9213,N_8011,N_8155);
nor U9214 (N_9214,N_8856,N_8374);
or U9215 (N_9215,N_8103,N_8948);
nand U9216 (N_9216,N_8674,N_8552);
or U9217 (N_9217,N_8050,N_8004);
nand U9218 (N_9218,N_8164,N_8279);
nor U9219 (N_9219,N_8229,N_8475);
and U9220 (N_9220,N_8143,N_8462);
nand U9221 (N_9221,N_8849,N_8379);
or U9222 (N_9222,N_8053,N_8122);
xnor U9223 (N_9223,N_8703,N_8744);
and U9224 (N_9224,N_8196,N_8521);
or U9225 (N_9225,N_8221,N_8028);
xor U9226 (N_9226,N_8793,N_8621);
or U9227 (N_9227,N_8132,N_8699);
and U9228 (N_9228,N_8217,N_8727);
or U9229 (N_9229,N_8759,N_8140);
or U9230 (N_9230,N_8653,N_8636);
or U9231 (N_9231,N_8224,N_8782);
xor U9232 (N_9232,N_8565,N_8946);
and U9233 (N_9233,N_8007,N_8538);
or U9234 (N_9234,N_8692,N_8453);
nor U9235 (N_9235,N_8655,N_8664);
nor U9236 (N_9236,N_8157,N_8835);
and U9237 (N_9237,N_8871,N_8940);
nor U9238 (N_9238,N_8215,N_8206);
xnor U9239 (N_9239,N_8798,N_8152);
xor U9240 (N_9240,N_8859,N_8845);
xor U9241 (N_9241,N_8023,N_8042);
nand U9242 (N_9242,N_8517,N_8094);
and U9243 (N_9243,N_8945,N_8310);
and U9244 (N_9244,N_8504,N_8757);
xnor U9245 (N_9245,N_8172,N_8988);
nor U9246 (N_9246,N_8449,N_8872);
nor U9247 (N_9247,N_8286,N_8180);
and U9248 (N_9248,N_8073,N_8547);
nor U9249 (N_9249,N_8677,N_8115);
and U9250 (N_9250,N_8506,N_8133);
or U9251 (N_9251,N_8333,N_8670);
nand U9252 (N_9252,N_8579,N_8726);
and U9253 (N_9253,N_8058,N_8775);
nand U9254 (N_9254,N_8352,N_8284);
xor U9255 (N_9255,N_8820,N_8483);
or U9256 (N_9256,N_8515,N_8705);
xor U9257 (N_9257,N_8977,N_8479);
nand U9258 (N_9258,N_8772,N_8811);
nor U9259 (N_9259,N_8124,N_8495);
nor U9260 (N_9260,N_8718,N_8188);
nor U9261 (N_9261,N_8501,N_8494);
nor U9262 (N_9262,N_8896,N_8894);
and U9263 (N_9263,N_8920,N_8629);
nand U9264 (N_9264,N_8016,N_8433);
and U9265 (N_9265,N_8673,N_8840);
and U9266 (N_9266,N_8341,N_8623);
or U9267 (N_9267,N_8958,N_8346);
nor U9268 (N_9268,N_8353,N_8870);
or U9269 (N_9269,N_8484,N_8251);
or U9270 (N_9270,N_8658,N_8168);
nor U9271 (N_9271,N_8116,N_8367);
or U9272 (N_9272,N_8074,N_8003);
nand U9273 (N_9273,N_8301,N_8197);
nand U9274 (N_9274,N_8532,N_8972);
nand U9275 (N_9275,N_8295,N_8216);
or U9276 (N_9276,N_8953,N_8420);
nor U9277 (N_9277,N_8630,N_8738);
nand U9278 (N_9278,N_8190,N_8944);
nor U9279 (N_9279,N_8498,N_8452);
and U9280 (N_9280,N_8675,N_8627);
or U9281 (N_9281,N_8034,N_8762);
nor U9282 (N_9282,N_8569,N_8963);
or U9283 (N_9283,N_8769,N_8600);
nand U9284 (N_9284,N_8804,N_8349);
or U9285 (N_9285,N_8737,N_8633);
nand U9286 (N_9286,N_8418,N_8465);
xor U9287 (N_9287,N_8365,N_8788);
nand U9288 (N_9288,N_8866,N_8359);
and U9289 (N_9289,N_8099,N_8381);
and U9290 (N_9290,N_8553,N_8145);
and U9291 (N_9291,N_8701,N_8244);
and U9292 (N_9292,N_8184,N_8010);
and U9293 (N_9293,N_8372,N_8130);
and U9294 (N_9294,N_8393,N_8632);
or U9295 (N_9295,N_8667,N_8767);
xor U9296 (N_9296,N_8414,N_8929);
xnor U9297 (N_9297,N_8430,N_8654);
or U9298 (N_9298,N_8450,N_8368);
nor U9299 (N_9299,N_8922,N_8888);
xnor U9300 (N_9300,N_8037,N_8020);
nand U9301 (N_9301,N_8982,N_8847);
xor U9302 (N_9302,N_8777,N_8142);
or U9303 (N_9303,N_8779,N_8942);
or U9304 (N_9304,N_8739,N_8411);
and U9305 (N_9305,N_8278,N_8696);
xnor U9306 (N_9306,N_8502,N_8421);
or U9307 (N_9307,N_8213,N_8610);
and U9308 (N_9308,N_8795,N_8296);
nand U9309 (N_9309,N_8543,N_8970);
and U9310 (N_9310,N_8493,N_8545);
nand U9311 (N_9311,N_8682,N_8913);
and U9312 (N_9312,N_8173,N_8398);
and U9313 (N_9313,N_8827,N_8285);
nor U9314 (N_9314,N_8275,N_8360);
nor U9315 (N_9315,N_8253,N_8711);
nor U9316 (N_9316,N_8980,N_8903);
nand U9317 (N_9317,N_8399,N_8668);
xnor U9318 (N_9318,N_8255,N_8964);
and U9319 (N_9319,N_8260,N_8614);
xor U9320 (N_9320,N_8153,N_8137);
nor U9321 (N_9321,N_8992,N_8356);
xor U9322 (N_9322,N_8170,N_8201);
nand U9323 (N_9323,N_8794,N_8555);
nor U9324 (N_9324,N_8257,N_8426);
or U9325 (N_9325,N_8854,N_8644);
nand U9326 (N_9326,N_8338,N_8047);
and U9327 (N_9327,N_8258,N_8478);
or U9328 (N_9328,N_8470,N_8489);
nor U9329 (N_9329,N_8413,N_8810);
or U9330 (N_9330,N_8592,N_8635);
and U9331 (N_9331,N_8836,N_8994);
nor U9332 (N_9332,N_8616,N_8646);
and U9333 (N_9333,N_8734,N_8593);
nor U9334 (N_9334,N_8778,N_8626);
xor U9335 (N_9335,N_8792,N_8339);
nand U9336 (N_9336,N_8148,N_8415);
xor U9337 (N_9337,N_8693,N_8021);
nand U9338 (N_9338,N_8661,N_8001);
xor U9339 (N_9339,N_8203,N_8247);
nor U9340 (N_9340,N_8969,N_8717);
or U9341 (N_9341,N_8748,N_8388);
or U9342 (N_9342,N_8038,N_8409);
nor U9343 (N_9343,N_8445,N_8604);
and U9344 (N_9344,N_8323,N_8706);
nand U9345 (N_9345,N_8620,N_8809);
and U9346 (N_9346,N_8851,N_8159);
nor U9347 (N_9347,N_8080,N_8281);
xor U9348 (N_9348,N_8466,N_8179);
nor U9349 (N_9349,N_8876,N_8904);
and U9350 (N_9350,N_8838,N_8787);
nor U9351 (N_9351,N_8193,N_8732);
nand U9352 (N_9352,N_8797,N_8831);
xnor U9353 (N_9353,N_8702,N_8086);
and U9354 (N_9354,N_8084,N_8685);
nor U9355 (N_9355,N_8488,N_8297);
nand U9356 (N_9356,N_8917,N_8033);
nor U9357 (N_9357,N_8017,N_8628);
nand U9358 (N_9358,N_8637,N_8051);
nand U9359 (N_9359,N_8526,N_8656);
and U9360 (N_9360,N_8207,N_8402);
nor U9361 (N_9361,N_8228,N_8887);
or U9362 (N_9362,N_8625,N_8649);
xor U9363 (N_9363,N_8391,N_8978);
xnor U9364 (N_9364,N_8974,N_8537);
or U9365 (N_9365,N_8102,N_8861);
nor U9366 (N_9366,N_8277,N_8246);
nand U9367 (N_9367,N_8098,N_8719);
nand U9368 (N_9368,N_8936,N_8476);
or U9369 (N_9369,N_8111,N_8716);
and U9370 (N_9370,N_8176,N_8619);
nand U9371 (N_9371,N_8167,N_8539);
or U9372 (N_9372,N_8121,N_8085);
xnor U9373 (N_9373,N_8015,N_8249);
nand U9374 (N_9374,N_8272,N_8800);
xor U9375 (N_9375,N_8631,N_8355);
and U9376 (N_9376,N_8335,N_8882);
nor U9377 (N_9377,N_8382,N_8818);
or U9378 (N_9378,N_8283,N_8417);
nand U9379 (N_9379,N_8527,N_8802);
and U9380 (N_9380,N_8117,N_8639);
xor U9381 (N_9381,N_8513,N_8932);
nand U9382 (N_9382,N_8087,N_8101);
xor U9383 (N_9383,N_8568,N_8723);
or U9384 (N_9384,N_8289,N_8348);
xnor U9385 (N_9385,N_8270,N_8304);
nand U9386 (N_9386,N_8540,N_8293);
and U9387 (N_9387,N_8204,N_8403);
and U9388 (N_9388,N_8330,N_8923);
xor U9389 (N_9389,N_8728,N_8530);
or U9390 (N_9390,N_8443,N_8129);
nor U9391 (N_9391,N_8182,N_8715);
nand U9392 (N_9392,N_8406,N_8239);
xnor U9393 (N_9393,N_8429,N_8486);
nor U9394 (N_9394,N_8886,N_8030);
or U9395 (N_9395,N_8503,N_8005);
or U9396 (N_9396,N_8318,N_8256);
or U9397 (N_9397,N_8366,N_8801);
and U9398 (N_9398,N_8874,N_8912);
or U9399 (N_9399,N_8043,N_8298);
and U9400 (N_9400,N_8187,N_8826);
nand U9401 (N_9401,N_8602,N_8199);
xnor U9402 (N_9402,N_8816,N_8690);
or U9403 (N_9403,N_8054,N_8100);
nand U9404 (N_9404,N_8211,N_8843);
or U9405 (N_9405,N_8151,N_8965);
or U9406 (N_9406,N_8514,N_8943);
or U9407 (N_9407,N_8471,N_8444);
and U9408 (N_9408,N_8305,N_8745);
nand U9409 (N_9409,N_8468,N_8822);
xnor U9410 (N_9410,N_8853,N_8704);
xnor U9411 (N_9411,N_8652,N_8266);
xor U9412 (N_9412,N_8344,N_8090);
xor U9413 (N_9413,N_8679,N_8095);
nand U9414 (N_9414,N_8225,N_8648);
or U9415 (N_9415,N_8268,N_8740);
nand U9416 (N_9416,N_8817,N_8079);
nand U9417 (N_9417,N_8742,N_8463);
xnor U9418 (N_9418,N_8350,N_8591);
and U9419 (N_9419,N_8786,N_8844);
xnor U9420 (N_9420,N_8469,N_8892);
nand U9421 (N_9421,N_8150,N_8436);
nand U9422 (N_9422,N_8227,N_8131);
nand U9423 (N_9423,N_8214,N_8609);
nand U9424 (N_9424,N_8574,N_8572);
or U9425 (N_9425,N_8570,N_8533);
nor U9426 (N_9426,N_8174,N_8908);
nor U9427 (N_9427,N_8959,N_8796);
and U9428 (N_9428,N_8605,N_8036);
and U9429 (N_9429,N_8282,N_8768);
nor U9430 (N_9430,N_8423,N_8448);
nor U9431 (N_9431,N_8299,N_8938);
or U9432 (N_9432,N_8821,N_8158);
xor U9433 (N_9433,N_8599,N_8899);
nor U9434 (N_9434,N_8814,N_8590);
and U9435 (N_9435,N_8081,N_8065);
xnor U9436 (N_9436,N_8259,N_8438);
xor U9437 (N_9437,N_8189,N_8280);
and U9438 (N_9438,N_8902,N_8419);
xor U9439 (N_9439,N_8889,N_8785);
nor U9440 (N_9440,N_8068,N_8194);
or U9441 (N_9441,N_8392,N_8774);
xnor U9442 (N_9442,N_8697,N_8534);
or U9443 (N_9443,N_8595,N_8107);
nand U9444 (N_9444,N_8713,N_8933);
xnor U9445 (N_9445,N_8990,N_8681);
or U9446 (N_9446,N_8618,N_8236);
or U9447 (N_9447,N_8686,N_8709);
nor U9448 (N_9448,N_8031,N_8612);
and U9449 (N_9449,N_8985,N_8096);
or U9450 (N_9450,N_8485,N_8319);
nor U9451 (N_9451,N_8089,N_8937);
nand U9452 (N_9452,N_8077,N_8294);
nor U9453 (N_9453,N_8380,N_8698);
and U9454 (N_9454,N_8714,N_8930);
nand U9455 (N_9455,N_8146,N_8110);
xnor U9456 (N_9456,N_8557,N_8645);
or U9457 (N_9457,N_8496,N_8926);
nand U9458 (N_9458,N_8935,N_8091);
or U9459 (N_9459,N_8910,N_8730);
xnor U9460 (N_9460,N_8321,N_8012);
nand U9461 (N_9461,N_8460,N_8390);
nor U9462 (N_9462,N_8106,N_8799);
nand U9463 (N_9463,N_8075,N_8461);
xor U9464 (N_9464,N_8070,N_8046);
nand U9465 (N_9465,N_8998,N_8045);
nand U9466 (N_9466,N_8264,N_8481);
nand U9467 (N_9467,N_8288,N_8114);
xnor U9468 (N_9468,N_8720,N_8700);
nor U9469 (N_9469,N_8966,N_8386);
xnor U9470 (N_9470,N_8509,N_8773);
xor U9471 (N_9471,N_8598,N_8437);
xor U9472 (N_9472,N_8956,N_8993);
xor U9473 (N_9473,N_8241,N_8694);
or U9474 (N_9474,N_8401,N_8883);
and U9475 (N_9475,N_8733,N_8136);
and U9476 (N_9476,N_8884,N_8960);
nand U9477 (N_9477,N_8315,N_8842);
nand U9478 (N_9478,N_8230,N_8432);
nor U9479 (N_9479,N_8248,N_8308);
nand U9480 (N_9480,N_8057,N_8022);
or U9481 (N_9481,N_8695,N_8435);
xnor U9482 (N_9482,N_8049,N_8878);
or U9483 (N_9483,N_8113,N_8458);
nor U9484 (N_9484,N_8410,N_8345);
nor U9485 (N_9485,N_8322,N_8808);
and U9486 (N_9486,N_8358,N_8263);
nor U9487 (N_9487,N_8660,N_8691);
and U9488 (N_9488,N_8672,N_8044);
and U9489 (N_9489,N_8040,N_8901);
and U9490 (N_9490,N_8725,N_8069);
nand U9491 (N_9491,N_8464,N_8564);
nor U9492 (N_9492,N_8529,N_8254);
xnor U9493 (N_9493,N_8141,N_8361);
nor U9494 (N_9494,N_8989,N_8973);
nor U9495 (N_9495,N_8955,N_8855);
or U9496 (N_9496,N_8191,N_8558);
xnor U9497 (N_9497,N_8320,N_8062);
or U9498 (N_9498,N_8603,N_8314);
nor U9499 (N_9499,N_8175,N_8947);
xnor U9500 (N_9500,N_8696,N_8829);
or U9501 (N_9501,N_8575,N_8149);
nor U9502 (N_9502,N_8843,N_8066);
or U9503 (N_9503,N_8483,N_8534);
nor U9504 (N_9504,N_8077,N_8413);
nand U9505 (N_9505,N_8469,N_8465);
nand U9506 (N_9506,N_8036,N_8177);
xor U9507 (N_9507,N_8345,N_8139);
or U9508 (N_9508,N_8500,N_8153);
nor U9509 (N_9509,N_8790,N_8124);
xnor U9510 (N_9510,N_8292,N_8029);
or U9511 (N_9511,N_8815,N_8814);
xnor U9512 (N_9512,N_8110,N_8494);
nand U9513 (N_9513,N_8227,N_8163);
and U9514 (N_9514,N_8153,N_8508);
nand U9515 (N_9515,N_8750,N_8453);
xnor U9516 (N_9516,N_8099,N_8326);
and U9517 (N_9517,N_8030,N_8455);
or U9518 (N_9518,N_8330,N_8005);
nor U9519 (N_9519,N_8131,N_8569);
and U9520 (N_9520,N_8650,N_8854);
and U9521 (N_9521,N_8136,N_8155);
xor U9522 (N_9522,N_8497,N_8935);
nor U9523 (N_9523,N_8927,N_8644);
or U9524 (N_9524,N_8872,N_8041);
or U9525 (N_9525,N_8567,N_8342);
nor U9526 (N_9526,N_8907,N_8204);
nand U9527 (N_9527,N_8812,N_8785);
nor U9528 (N_9528,N_8317,N_8661);
or U9529 (N_9529,N_8408,N_8685);
and U9530 (N_9530,N_8108,N_8364);
nand U9531 (N_9531,N_8276,N_8978);
nor U9532 (N_9532,N_8846,N_8664);
xnor U9533 (N_9533,N_8474,N_8929);
nand U9534 (N_9534,N_8484,N_8687);
xor U9535 (N_9535,N_8962,N_8434);
and U9536 (N_9536,N_8769,N_8489);
nor U9537 (N_9537,N_8225,N_8498);
and U9538 (N_9538,N_8934,N_8812);
nand U9539 (N_9539,N_8722,N_8438);
or U9540 (N_9540,N_8443,N_8426);
and U9541 (N_9541,N_8457,N_8507);
and U9542 (N_9542,N_8978,N_8890);
nor U9543 (N_9543,N_8462,N_8027);
nor U9544 (N_9544,N_8234,N_8549);
nand U9545 (N_9545,N_8666,N_8155);
or U9546 (N_9546,N_8265,N_8140);
xor U9547 (N_9547,N_8438,N_8138);
or U9548 (N_9548,N_8134,N_8257);
or U9549 (N_9549,N_8400,N_8974);
and U9550 (N_9550,N_8310,N_8603);
xor U9551 (N_9551,N_8048,N_8994);
and U9552 (N_9552,N_8029,N_8538);
nand U9553 (N_9553,N_8204,N_8289);
and U9554 (N_9554,N_8165,N_8147);
and U9555 (N_9555,N_8847,N_8578);
nand U9556 (N_9556,N_8169,N_8234);
xnor U9557 (N_9557,N_8699,N_8258);
xnor U9558 (N_9558,N_8686,N_8881);
nand U9559 (N_9559,N_8393,N_8061);
and U9560 (N_9560,N_8211,N_8894);
nand U9561 (N_9561,N_8986,N_8630);
nand U9562 (N_9562,N_8283,N_8710);
xor U9563 (N_9563,N_8626,N_8507);
xnor U9564 (N_9564,N_8309,N_8545);
or U9565 (N_9565,N_8438,N_8593);
nor U9566 (N_9566,N_8934,N_8540);
nand U9567 (N_9567,N_8917,N_8020);
nor U9568 (N_9568,N_8356,N_8587);
xnor U9569 (N_9569,N_8897,N_8102);
and U9570 (N_9570,N_8718,N_8340);
xnor U9571 (N_9571,N_8540,N_8495);
and U9572 (N_9572,N_8201,N_8248);
or U9573 (N_9573,N_8420,N_8333);
or U9574 (N_9574,N_8010,N_8282);
xor U9575 (N_9575,N_8205,N_8040);
and U9576 (N_9576,N_8259,N_8450);
and U9577 (N_9577,N_8878,N_8036);
and U9578 (N_9578,N_8342,N_8053);
and U9579 (N_9579,N_8304,N_8195);
nand U9580 (N_9580,N_8045,N_8424);
and U9581 (N_9581,N_8831,N_8212);
or U9582 (N_9582,N_8137,N_8465);
or U9583 (N_9583,N_8779,N_8376);
nand U9584 (N_9584,N_8444,N_8334);
nand U9585 (N_9585,N_8153,N_8453);
nand U9586 (N_9586,N_8123,N_8353);
and U9587 (N_9587,N_8803,N_8981);
xor U9588 (N_9588,N_8966,N_8107);
xor U9589 (N_9589,N_8250,N_8732);
xnor U9590 (N_9590,N_8898,N_8236);
nand U9591 (N_9591,N_8769,N_8599);
nand U9592 (N_9592,N_8325,N_8717);
nor U9593 (N_9593,N_8560,N_8321);
xor U9594 (N_9594,N_8853,N_8857);
nor U9595 (N_9595,N_8083,N_8487);
xnor U9596 (N_9596,N_8359,N_8514);
or U9597 (N_9597,N_8349,N_8956);
nand U9598 (N_9598,N_8326,N_8727);
or U9599 (N_9599,N_8709,N_8129);
or U9600 (N_9600,N_8314,N_8225);
xor U9601 (N_9601,N_8353,N_8035);
nand U9602 (N_9602,N_8736,N_8021);
nor U9603 (N_9603,N_8951,N_8384);
and U9604 (N_9604,N_8228,N_8215);
xor U9605 (N_9605,N_8272,N_8410);
and U9606 (N_9606,N_8375,N_8208);
and U9607 (N_9607,N_8441,N_8811);
nand U9608 (N_9608,N_8884,N_8540);
nand U9609 (N_9609,N_8080,N_8715);
xor U9610 (N_9610,N_8389,N_8510);
and U9611 (N_9611,N_8646,N_8042);
or U9612 (N_9612,N_8432,N_8736);
xnor U9613 (N_9613,N_8895,N_8187);
or U9614 (N_9614,N_8662,N_8733);
nor U9615 (N_9615,N_8168,N_8928);
nand U9616 (N_9616,N_8257,N_8006);
xor U9617 (N_9617,N_8109,N_8307);
or U9618 (N_9618,N_8462,N_8689);
or U9619 (N_9619,N_8516,N_8035);
and U9620 (N_9620,N_8503,N_8312);
nand U9621 (N_9621,N_8297,N_8683);
or U9622 (N_9622,N_8174,N_8659);
and U9623 (N_9623,N_8835,N_8105);
and U9624 (N_9624,N_8438,N_8271);
nand U9625 (N_9625,N_8349,N_8316);
nor U9626 (N_9626,N_8848,N_8779);
nor U9627 (N_9627,N_8304,N_8409);
nand U9628 (N_9628,N_8284,N_8451);
xor U9629 (N_9629,N_8659,N_8937);
nor U9630 (N_9630,N_8991,N_8813);
and U9631 (N_9631,N_8108,N_8969);
nand U9632 (N_9632,N_8313,N_8736);
and U9633 (N_9633,N_8057,N_8804);
nand U9634 (N_9634,N_8398,N_8245);
nand U9635 (N_9635,N_8971,N_8509);
nand U9636 (N_9636,N_8109,N_8857);
or U9637 (N_9637,N_8542,N_8160);
and U9638 (N_9638,N_8520,N_8815);
or U9639 (N_9639,N_8813,N_8008);
nor U9640 (N_9640,N_8236,N_8006);
and U9641 (N_9641,N_8189,N_8224);
or U9642 (N_9642,N_8789,N_8403);
nand U9643 (N_9643,N_8532,N_8217);
nand U9644 (N_9644,N_8299,N_8453);
nand U9645 (N_9645,N_8293,N_8904);
and U9646 (N_9646,N_8233,N_8277);
or U9647 (N_9647,N_8642,N_8033);
nor U9648 (N_9648,N_8949,N_8414);
xor U9649 (N_9649,N_8521,N_8708);
or U9650 (N_9650,N_8394,N_8165);
xor U9651 (N_9651,N_8941,N_8819);
nand U9652 (N_9652,N_8856,N_8687);
xor U9653 (N_9653,N_8836,N_8946);
and U9654 (N_9654,N_8641,N_8873);
xor U9655 (N_9655,N_8747,N_8355);
or U9656 (N_9656,N_8601,N_8054);
xnor U9657 (N_9657,N_8047,N_8749);
nand U9658 (N_9658,N_8153,N_8039);
xor U9659 (N_9659,N_8579,N_8341);
nor U9660 (N_9660,N_8721,N_8099);
or U9661 (N_9661,N_8021,N_8484);
xor U9662 (N_9662,N_8795,N_8624);
or U9663 (N_9663,N_8872,N_8578);
nor U9664 (N_9664,N_8142,N_8072);
and U9665 (N_9665,N_8107,N_8136);
xor U9666 (N_9666,N_8929,N_8125);
xnor U9667 (N_9667,N_8776,N_8770);
nor U9668 (N_9668,N_8414,N_8702);
nor U9669 (N_9669,N_8387,N_8206);
nor U9670 (N_9670,N_8172,N_8466);
nor U9671 (N_9671,N_8935,N_8516);
xor U9672 (N_9672,N_8519,N_8642);
nor U9673 (N_9673,N_8847,N_8957);
nor U9674 (N_9674,N_8848,N_8071);
or U9675 (N_9675,N_8906,N_8066);
nand U9676 (N_9676,N_8949,N_8079);
xnor U9677 (N_9677,N_8878,N_8752);
nor U9678 (N_9678,N_8128,N_8136);
nand U9679 (N_9679,N_8476,N_8719);
nor U9680 (N_9680,N_8174,N_8088);
or U9681 (N_9681,N_8077,N_8881);
nand U9682 (N_9682,N_8705,N_8683);
or U9683 (N_9683,N_8281,N_8738);
nand U9684 (N_9684,N_8799,N_8154);
nor U9685 (N_9685,N_8171,N_8481);
and U9686 (N_9686,N_8796,N_8690);
and U9687 (N_9687,N_8246,N_8932);
nor U9688 (N_9688,N_8272,N_8436);
nand U9689 (N_9689,N_8584,N_8365);
and U9690 (N_9690,N_8182,N_8839);
nor U9691 (N_9691,N_8466,N_8424);
nor U9692 (N_9692,N_8735,N_8610);
and U9693 (N_9693,N_8604,N_8018);
and U9694 (N_9694,N_8602,N_8702);
and U9695 (N_9695,N_8537,N_8774);
or U9696 (N_9696,N_8687,N_8069);
nor U9697 (N_9697,N_8022,N_8206);
and U9698 (N_9698,N_8061,N_8831);
xor U9699 (N_9699,N_8617,N_8562);
xnor U9700 (N_9700,N_8303,N_8475);
nand U9701 (N_9701,N_8040,N_8483);
nor U9702 (N_9702,N_8695,N_8905);
nand U9703 (N_9703,N_8104,N_8946);
nand U9704 (N_9704,N_8268,N_8704);
and U9705 (N_9705,N_8990,N_8747);
nand U9706 (N_9706,N_8461,N_8521);
nor U9707 (N_9707,N_8964,N_8326);
xor U9708 (N_9708,N_8750,N_8631);
nor U9709 (N_9709,N_8229,N_8908);
nand U9710 (N_9710,N_8068,N_8358);
nor U9711 (N_9711,N_8544,N_8799);
nand U9712 (N_9712,N_8721,N_8340);
nor U9713 (N_9713,N_8376,N_8056);
or U9714 (N_9714,N_8547,N_8136);
xnor U9715 (N_9715,N_8769,N_8869);
or U9716 (N_9716,N_8045,N_8642);
xnor U9717 (N_9717,N_8136,N_8477);
xor U9718 (N_9718,N_8364,N_8427);
and U9719 (N_9719,N_8861,N_8910);
nand U9720 (N_9720,N_8029,N_8076);
and U9721 (N_9721,N_8161,N_8378);
and U9722 (N_9722,N_8641,N_8689);
and U9723 (N_9723,N_8576,N_8958);
and U9724 (N_9724,N_8046,N_8676);
or U9725 (N_9725,N_8616,N_8936);
nor U9726 (N_9726,N_8088,N_8845);
or U9727 (N_9727,N_8433,N_8085);
and U9728 (N_9728,N_8254,N_8439);
xor U9729 (N_9729,N_8598,N_8753);
xnor U9730 (N_9730,N_8325,N_8907);
and U9731 (N_9731,N_8765,N_8545);
or U9732 (N_9732,N_8464,N_8050);
or U9733 (N_9733,N_8680,N_8541);
and U9734 (N_9734,N_8852,N_8571);
and U9735 (N_9735,N_8067,N_8885);
nand U9736 (N_9736,N_8181,N_8095);
nor U9737 (N_9737,N_8265,N_8771);
nor U9738 (N_9738,N_8144,N_8143);
xnor U9739 (N_9739,N_8700,N_8264);
nor U9740 (N_9740,N_8537,N_8352);
xor U9741 (N_9741,N_8693,N_8216);
and U9742 (N_9742,N_8794,N_8360);
nor U9743 (N_9743,N_8061,N_8577);
nor U9744 (N_9744,N_8824,N_8969);
nor U9745 (N_9745,N_8882,N_8326);
xnor U9746 (N_9746,N_8322,N_8150);
and U9747 (N_9747,N_8291,N_8690);
and U9748 (N_9748,N_8673,N_8252);
nand U9749 (N_9749,N_8833,N_8249);
nor U9750 (N_9750,N_8374,N_8177);
xnor U9751 (N_9751,N_8176,N_8517);
and U9752 (N_9752,N_8613,N_8975);
and U9753 (N_9753,N_8718,N_8383);
nand U9754 (N_9754,N_8190,N_8392);
and U9755 (N_9755,N_8382,N_8286);
nand U9756 (N_9756,N_8577,N_8542);
nand U9757 (N_9757,N_8997,N_8761);
or U9758 (N_9758,N_8891,N_8938);
nor U9759 (N_9759,N_8295,N_8669);
xor U9760 (N_9760,N_8136,N_8479);
xnor U9761 (N_9761,N_8834,N_8282);
or U9762 (N_9762,N_8598,N_8296);
or U9763 (N_9763,N_8452,N_8776);
or U9764 (N_9764,N_8166,N_8634);
xor U9765 (N_9765,N_8782,N_8312);
or U9766 (N_9766,N_8018,N_8983);
and U9767 (N_9767,N_8529,N_8988);
and U9768 (N_9768,N_8574,N_8079);
or U9769 (N_9769,N_8224,N_8519);
or U9770 (N_9770,N_8856,N_8861);
nor U9771 (N_9771,N_8516,N_8539);
xor U9772 (N_9772,N_8549,N_8426);
nor U9773 (N_9773,N_8987,N_8567);
and U9774 (N_9774,N_8539,N_8775);
xor U9775 (N_9775,N_8243,N_8541);
xnor U9776 (N_9776,N_8287,N_8837);
or U9777 (N_9777,N_8900,N_8112);
or U9778 (N_9778,N_8635,N_8505);
or U9779 (N_9779,N_8296,N_8592);
nor U9780 (N_9780,N_8366,N_8979);
xnor U9781 (N_9781,N_8016,N_8349);
xnor U9782 (N_9782,N_8637,N_8072);
nand U9783 (N_9783,N_8420,N_8573);
and U9784 (N_9784,N_8347,N_8822);
xor U9785 (N_9785,N_8265,N_8751);
or U9786 (N_9786,N_8067,N_8032);
or U9787 (N_9787,N_8213,N_8446);
nand U9788 (N_9788,N_8184,N_8812);
nor U9789 (N_9789,N_8444,N_8886);
and U9790 (N_9790,N_8286,N_8141);
xnor U9791 (N_9791,N_8981,N_8805);
xor U9792 (N_9792,N_8237,N_8530);
or U9793 (N_9793,N_8496,N_8048);
and U9794 (N_9794,N_8727,N_8565);
xnor U9795 (N_9795,N_8212,N_8976);
nor U9796 (N_9796,N_8067,N_8385);
and U9797 (N_9797,N_8287,N_8244);
nand U9798 (N_9798,N_8070,N_8321);
nor U9799 (N_9799,N_8381,N_8822);
and U9800 (N_9800,N_8858,N_8545);
or U9801 (N_9801,N_8770,N_8743);
or U9802 (N_9802,N_8194,N_8337);
or U9803 (N_9803,N_8167,N_8199);
and U9804 (N_9804,N_8167,N_8776);
xnor U9805 (N_9805,N_8675,N_8638);
or U9806 (N_9806,N_8719,N_8739);
nor U9807 (N_9807,N_8520,N_8056);
xnor U9808 (N_9808,N_8496,N_8190);
nand U9809 (N_9809,N_8134,N_8645);
and U9810 (N_9810,N_8990,N_8722);
xor U9811 (N_9811,N_8147,N_8806);
nand U9812 (N_9812,N_8060,N_8158);
or U9813 (N_9813,N_8659,N_8991);
nor U9814 (N_9814,N_8845,N_8370);
or U9815 (N_9815,N_8536,N_8651);
nand U9816 (N_9816,N_8384,N_8340);
or U9817 (N_9817,N_8858,N_8091);
or U9818 (N_9818,N_8359,N_8288);
nand U9819 (N_9819,N_8230,N_8812);
or U9820 (N_9820,N_8972,N_8808);
nor U9821 (N_9821,N_8640,N_8666);
and U9822 (N_9822,N_8806,N_8107);
or U9823 (N_9823,N_8915,N_8012);
nor U9824 (N_9824,N_8527,N_8836);
or U9825 (N_9825,N_8633,N_8383);
xnor U9826 (N_9826,N_8907,N_8580);
nand U9827 (N_9827,N_8495,N_8483);
nor U9828 (N_9828,N_8855,N_8727);
nor U9829 (N_9829,N_8593,N_8640);
xnor U9830 (N_9830,N_8298,N_8979);
xnor U9831 (N_9831,N_8792,N_8411);
or U9832 (N_9832,N_8739,N_8294);
and U9833 (N_9833,N_8411,N_8989);
and U9834 (N_9834,N_8488,N_8864);
nor U9835 (N_9835,N_8119,N_8198);
and U9836 (N_9836,N_8666,N_8607);
nand U9837 (N_9837,N_8837,N_8757);
nand U9838 (N_9838,N_8406,N_8534);
xor U9839 (N_9839,N_8600,N_8704);
xor U9840 (N_9840,N_8537,N_8431);
nand U9841 (N_9841,N_8620,N_8478);
nor U9842 (N_9842,N_8698,N_8981);
or U9843 (N_9843,N_8417,N_8913);
xnor U9844 (N_9844,N_8243,N_8169);
or U9845 (N_9845,N_8403,N_8961);
xnor U9846 (N_9846,N_8009,N_8922);
or U9847 (N_9847,N_8558,N_8805);
xor U9848 (N_9848,N_8418,N_8537);
or U9849 (N_9849,N_8882,N_8464);
xnor U9850 (N_9850,N_8614,N_8211);
and U9851 (N_9851,N_8759,N_8295);
and U9852 (N_9852,N_8406,N_8383);
nand U9853 (N_9853,N_8407,N_8425);
or U9854 (N_9854,N_8783,N_8021);
xnor U9855 (N_9855,N_8203,N_8822);
and U9856 (N_9856,N_8892,N_8900);
nand U9857 (N_9857,N_8292,N_8003);
xor U9858 (N_9858,N_8151,N_8587);
or U9859 (N_9859,N_8624,N_8043);
and U9860 (N_9860,N_8445,N_8974);
nand U9861 (N_9861,N_8846,N_8453);
nand U9862 (N_9862,N_8169,N_8472);
xor U9863 (N_9863,N_8244,N_8766);
xor U9864 (N_9864,N_8052,N_8768);
or U9865 (N_9865,N_8193,N_8114);
and U9866 (N_9866,N_8445,N_8592);
nor U9867 (N_9867,N_8381,N_8228);
or U9868 (N_9868,N_8354,N_8147);
nor U9869 (N_9869,N_8349,N_8025);
or U9870 (N_9870,N_8031,N_8609);
or U9871 (N_9871,N_8883,N_8350);
and U9872 (N_9872,N_8685,N_8670);
and U9873 (N_9873,N_8810,N_8452);
xnor U9874 (N_9874,N_8557,N_8868);
nor U9875 (N_9875,N_8149,N_8209);
xor U9876 (N_9876,N_8499,N_8660);
or U9877 (N_9877,N_8784,N_8915);
nor U9878 (N_9878,N_8075,N_8762);
nand U9879 (N_9879,N_8219,N_8646);
and U9880 (N_9880,N_8036,N_8438);
nand U9881 (N_9881,N_8567,N_8228);
xnor U9882 (N_9882,N_8445,N_8494);
nand U9883 (N_9883,N_8194,N_8662);
nand U9884 (N_9884,N_8210,N_8930);
and U9885 (N_9885,N_8737,N_8538);
xor U9886 (N_9886,N_8182,N_8211);
nand U9887 (N_9887,N_8412,N_8229);
nor U9888 (N_9888,N_8792,N_8342);
or U9889 (N_9889,N_8763,N_8779);
or U9890 (N_9890,N_8543,N_8545);
and U9891 (N_9891,N_8422,N_8029);
and U9892 (N_9892,N_8742,N_8110);
nor U9893 (N_9893,N_8335,N_8003);
nor U9894 (N_9894,N_8079,N_8905);
or U9895 (N_9895,N_8688,N_8528);
or U9896 (N_9896,N_8929,N_8869);
and U9897 (N_9897,N_8487,N_8846);
xnor U9898 (N_9898,N_8489,N_8571);
xor U9899 (N_9899,N_8022,N_8335);
and U9900 (N_9900,N_8716,N_8785);
xor U9901 (N_9901,N_8662,N_8602);
and U9902 (N_9902,N_8600,N_8094);
and U9903 (N_9903,N_8337,N_8229);
nand U9904 (N_9904,N_8227,N_8921);
xor U9905 (N_9905,N_8285,N_8554);
nor U9906 (N_9906,N_8290,N_8652);
nand U9907 (N_9907,N_8170,N_8552);
or U9908 (N_9908,N_8680,N_8626);
or U9909 (N_9909,N_8926,N_8201);
and U9910 (N_9910,N_8524,N_8434);
nand U9911 (N_9911,N_8401,N_8515);
nand U9912 (N_9912,N_8771,N_8671);
and U9913 (N_9913,N_8451,N_8486);
nor U9914 (N_9914,N_8724,N_8192);
nor U9915 (N_9915,N_8514,N_8109);
nand U9916 (N_9916,N_8367,N_8877);
and U9917 (N_9917,N_8087,N_8631);
or U9918 (N_9918,N_8757,N_8323);
nor U9919 (N_9919,N_8923,N_8602);
nand U9920 (N_9920,N_8095,N_8741);
nor U9921 (N_9921,N_8646,N_8834);
nor U9922 (N_9922,N_8601,N_8304);
nand U9923 (N_9923,N_8562,N_8491);
and U9924 (N_9924,N_8429,N_8791);
nor U9925 (N_9925,N_8510,N_8518);
or U9926 (N_9926,N_8209,N_8295);
nand U9927 (N_9927,N_8650,N_8831);
nor U9928 (N_9928,N_8481,N_8501);
and U9929 (N_9929,N_8188,N_8712);
xor U9930 (N_9930,N_8825,N_8185);
or U9931 (N_9931,N_8864,N_8037);
xor U9932 (N_9932,N_8442,N_8783);
nand U9933 (N_9933,N_8383,N_8628);
xor U9934 (N_9934,N_8225,N_8487);
and U9935 (N_9935,N_8343,N_8199);
and U9936 (N_9936,N_8657,N_8658);
or U9937 (N_9937,N_8599,N_8507);
nor U9938 (N_9938,N_8380,N_8290);
xor U9939 (N_9939,N_8522,N_8143);
nor U9940 (N_9940,N_8512,N_8172);
or U9941 (N_9941,N_8193,N_8267);
or U9942 (N_9942,N_8580,N_8276);
and U9943 (N_9943,N_8233,N_8528);
and U9944 (N_9944,N_8478,N_8906);
nor U9945 (N_9945,N_8771,N_8701);
nor U9946 (N_9946,N_8556,N_8926);
or U9947 (N_9947,N_8571,N_8213);
nand U9948 (N_9948,N_8023,N_8549);
nor U9949 (N_9949,N_8073,N_8628);
nor U9950 (N_9950,N_8802,N_8654);
and U9951 (N_9951,N_8920,N_8698);
nand U9952 (N_9952,N_8248,N_8262);
xnor U9953 (N_9953,N_8088,N_8495);
or U9954 (N_9954,N_8540,N_8131);
and U9955 (N_9955,N_8006,N_8203);
nand U9956 (N_9956,N_8554,N_8333);
nor U9957 (N_9957,N_8278,N_8406);
or U9958 (N_9958,N_8204,N_8860);
nor U9959 (N_9959,N_8755,N_8161);
xor U9960 (N_9960,N_8753,N_8952);
nor U9961 (N_9961,N_8879,N_8318);
and U9962 (N_9962,N_8243,N_8266);
or U9963 (N_9963,N_8879,N_8343);
xor U9964 (N_9964,N_8040,N_8268);
xnor U9965 (N_9965,N_8678,N_8166);
xnor U9966 (N_9966,N_8731,N_8766);
xnor U9967 (N_9967,N_8240,N_8664);
nor U9968 (N_9968,N_8568,N_8753);
nor U9969 (N_9969,N_8951,N_8998);
xnor U9970 (N_9970,N_8256,N_8721);
and U9971 (N_9971,N_8650,N_8729);
and U9972 (N_9972,N_8589,N_8289);
nand U9973 (N_9973,N_8178,N_8430);
or U9974 (N_9974,N_8361,N_8032);
or U9975 (N_9975,N_8882,N_8306);
and U9976 (N_9976,N_8358,N_8212);
xor U9977 (N_9977,N_8395,N_8427);
or U9978 (N_9978,N_8420,N_8356);
or U9979 (N_9979,N_8060,N_8054);
xnor U9980 (N_9980,N_8377,N_8127);
xnor U9981 (N_9981,N_8858,N_8265);
and U9982 (N_9982,N_8806,N_8075);
nor U9983 (N_9983,N_8165,N_8732);
nor U9984 (N_9984,N_8470,N_8822);
and U9985 (N_9985,N_8833,N_8811);
or U9986 (N_9986,N_8629,N_8344);
nand U9987 (N_9987,N_8305,N_8526);
nand U9988 (N_9988,N_8011,N_8878);
or U9989 (N_9989,N_8969,N_8348);
xor U9990 (N_9990,N_8800,N_8702);
nor U9991 (N_9991,N_8483,N_8113);
nor U9992 (N_9992,N_8572,N_8467);
xor U9993 (N_9993,N_8246,N_8875);
or U9994 (N_9994,N_8266,N_8992);
nor U9995 (N_9995,N_8551,N_8799);
nand U9996 (N_9996,N_8405,N_8718);
or U9997 (N_9997,N_8685,N_8837);
and U9998 (N_9998,N_8887,N_8459);
xnor U9999 (N_9999,N_8249,N_8076);
and U10000 (N_10000,N_9918,N_9012);
nand U10001 (N_10001,N_9287,N_9372);
nand U10002 (N_10002,N_9333,N_9415);
or U10003 (N_10003,N_9029,N_9110);
and U10004 (N_10004,N_9246,N_9574);
or U10005 (N_10005,N_9152,N_9185);
or U10006 (N_10006,N_9221,N_9472);
nand U10007 (N_10007,N_9857,N_9627);
and U10008 (N_10008,N_9102,N_9626);
and U10009 (N_10009,N_9463,N_9760);
xnor U10010 (N_10010,N_9800,N_9780);
xor U10011 (N_10011,N_9389,N_9986);
xor U10012 (N_10012,N_9452,N_9514);
xnor U10013 (N_10013,N_9314,N_9925);
xor U10014 (N_10014,N_9190,N_9488);
xnor U10015 (N_10015,N_9787,N_9891);
and U10016 (N_10016,N_9070,N_9873);
and U10017 (N_10017,N_9090,N_9080);
nor U10018 (N_10018,N_9635,N_9535);
nor U10019 (N_10019,N_9837,N_9318);
or U10020 (N_10020,N_9100,N_9946);
or U10021 (N_10021,N_9822,N_9607);
and U10022 (N_10022,N_9099,N_9790);
nand U10023 (N_10023,N_9832,N_9570);
xor U10024 (N_10024,N_9376,N_9276);
xor U10025 (N_10025,N_9758,N_9244);
or U10026 (N_10026,N_9293,N_9004);
xnor U10027 (N_10027,N_9138,N_9763);
nand U10028 (N_10028,N_9727,N_9936);
xnor U10029 (N_10029,N_9159,N_9157);
nand U10030 (N_10030,N_9002,N_9878);
nor U10031 (N_10031,N_9056,N_9967);
nor U10032 (N_10032,N_9529,N_9236);
nand U10033 (N_10033,N_9059,N_9641);
or U10034 (N_10034,N_9091,N_9541);
or U10035 (N_10035,N_9632,N_9782);
and U10036 (N_10036,N_9567,N_9937);
xor U10037 (N_10037,N_9438,N_9904);
nor U10038 (N_10038,N_9669,N_9829);
and U10039 (N_10039,N_9137,N_9629);
and U10040 (N_10040,N_9752,N_9382);
xnor U10041 (N_10041,N_9944,N_9818);
or U10042 (N_10042,N_9815,N_9942);
or U10043 (N_10043,N_9660,N_9571);
and U10044 (N_10044,N_9951,N_9261);
and U10045 (N_10045,N_9850,N_9473);
or U10046 (N_10046,N_9860,N_9493);
and U10047 (N_10047,N_9969,N_9442);
nand U10048 (N_10048,N_9528,N_9028);
nand U10049 (N_10049,N_9653,N_9055);
nand U10050 (N_10050,N_9612,N_9062);
and U10051 (N_10051,N_9783,N_9882);
and U10052 (N_10052,N_9801,N_9714);
or U10053 (N_10053,N_9726,N_9699);
and U10054 (N_10054,N_9677,N_9756);
or U10055 (N_10055,N_9953,N_9998);
xnor U10056 (N_10056,N_9344,N_9411);
nor U10057 (N_10057,N_9409,N_9482);
xnor U10058 (N_10058,N_9458,N_9484);
nor U10059 (N_10059,N_9156,N_9527);
nor U10060 (N_10060,N_9712,N_9875);
nand U10061 (N_10061,N_9720,N_9419);
xor U10062 (N_10062,N_9604,N_9810);
and U10063 (N_10063,N_9087,N_9025);
nor U10064 (N_10064,N_9692,N_9863);
or U10065 (N_10065,N_9310,N_9922);
nand U10066 (N_10066,N_9346,N_9499);
and U10067 (N_10067,N_9022,N_9196);
nand U10068 (N_10068,N_9864,N_9417);
nand U10069 (N_10069,N_9716,N_9877);
nand U10070 (N_10070,N_9271,N_9189);
and U10071 (N_10071,N_9869,N_9279);
xor U10072 (N_10072,N_9448,N_9521);
nor U10073 (N_10073,N_9885,N_9048);
nand U10074 (N_10074,N_9114,N_9562);
nand U10075 (N_10075,N_9708,N_9956);
nand U10076 (N_10076,N_9399,N_9961);
or U10077 (N_10077,N_9556,N_9664);
xor U10078 (N_10078,N_9609,N_9950);
nor U10079 (N_10079,N_9693,N_9021);
and U10080 (N_10080,N_9470,N_9757);
nor U10081 (N_10081,N_9454,N_9578);
or U10082 (N_10082,N_9487,N_9146);
or U10083 (N_10083,N_9921,N_9777);
xnor U10084 (N_10084,N_9565,N_9175);
xor U10085 (N_10085,N_9642,N_9453);
xnor U10086 (N_10086,N_9665,N_9394);
xor U10087 (N_10087,N_9687,N_9744);
and U10088 (N_10088,N_9148,N_9806);
and U10089 (N_10089,N_9977,N_9823);
nor U10090 (N_10090,N_9990,N_9019);
xnor U10091 (N_10091,N_9902,N_9077);
nor U10092 (N_10092,N_9064,N_9218);
nor U10093 (N_10093,N_9151,N_9180);
nand U10094 (N_10094,N_9930,N_9229);
xnor U10095 (N_10095,N_9351,N_9281);
nand U10096 (N_10096,N_9395,N_9037);
xor U10097 (N_10097,N_9948,N_9150);
and U10098 (N_10098,N_9549,N_9427);
nand U10099 (N_10099,N_9054,N_9282);
or U10100 (N_10100,N_9928,N_9174);
and U10101 (N_10101,N_9347,N_9187);
nor U10102 (N_10102,N_9000,N_9781);
or U10103 (N_10103,N_9809,N_9836);
xnor U10104 (N_10104,N_9721,N_9071);
and U10105 (N_10105,N_9994,N_9509);
nand U10106 (N_10106,N_9081,N_9234);
xor U10107 (N_10107,N_9126,N_9910);
nor U10108 (N_10108,N_9589,N_9413);
or U10109 (N_10109,N_9980,N_9602);
and U10110 (N_10110,N_9648,N_9290);
or U10111 (N_10111,N_9769,N_9416);
or U10112 (N_10112,N_9742,N_9033);
xor U10113 (N_10113,N_9212,N_9981);
nor U10114 (N_10114,N_9608,N_9125);
and U10115 (N_10115,N_9865,N_9779);
nor U10116 (N_10116,N_9663,N_9030);
nor U10117 (N_10117,N_9817,N_9265);
nand U10118 (N_10118,N_9480,N_9251);
nor U10119 (N_10119,N_9294,N_9119);
and U10120 (N_10120,N_9704,N_9886);
nor U10121 (N_10121,N_9661,N_9729);
and U10122 (N_10122,N_9407,N_9354);
nor U10123 (N_10123,N_9222,N_9406);
xnor U10124 (N_10124,N_9034,N_9084);
nand U10125 (N_10125,N_9547,N_9459);
or U10126 (N_10126,N_9598,N_9935);
nand U10127 (N_10127,N_9031,N_9974);
nand U10128 (N_10128,N_9469,N_9610);
or U10129 (N_10129,N_9239,N_9437);
and U10130 (N_10130,N_9106,N_9444);
and U10131 (N_10131,N_9775,N_9724);
nand U10132 (N_10132,N_9447,N_9205);
and U10133 (N_10133,N_9941,N_9590);
xnor U10134 (N_10134,N_9804,N_9041);
nor U10135 (N_10135,N_9555,N_9262);
and U10136 (N_10136,N_9923,N_9300);
xor U10137 (N_10137,N_9580,N_9995);
xnor U10138 (N_10138,N_9361,N_9621);
xor U10139 (N_10139,N_9552,N_9073);
nand U10140 (N_10140,N_9101,N_9924);
nand U10141 (N_10141,N_9206,N_9349);
nand U10142 (N_10142,N_9434,N_9465);
or U10143 (N_10143,N_9975,N_9063);
or U10144 (N_10144,N_9622,N_9979);
nor U10145 (N_10145,N_9519,N_9847);
xnor U10146 (N_10146,N_9518,N_9467);
nor U10147 (N_10147,N_9583,N_9136);
and U10148 (N_10148,N_9008,N_9027);
and U10149 (N_10149,N_9320,N_9841);
nand U10150 (N_10150,N_9410,N_9855);
nor U10151 (N_10151,N_9121,N_9304);
xnor U10152 (N_10152,N_9182,N_9732);
nand U10153 (N_10153,N_9184,N_9620);
or U10154 (N_10154,N_9939,N_9365);
nor U10155 (N_10155,N_9132,N_9384);
or U10156 (N_10156,N_9984,N_9581);
xor U10157 (N_10157,N_9036,N_9165);
nor U10158 (N_10158,N_9844,N_9539);
or U10159 (N_10159,N_9173,N_9796);
or U10160 (N_10160,N_9501,N_9371);
and U10161 (N_10161,N_9713,N_9826);
xnor U10162 (N_10162,N_9795,N_9163);
nor U10163 (N_10163,N_9507,N_9671);
xnor U10164 (N_10164,N_9883,N_9614);
and U10165 (N_10165,N_9049,N_9741);
xor U10166 (N_10166,N_9778,N_9353);
and U10167 (N_10167,N_9658,N_9587);
and U10168 (N_10168,N_9147,N_9605);
nand U10169 (N_10169,N_9814,N_9845);
nand U10170 (N_10170,N_9531,N_9217);
or U10171 (N_10171,N_9412,N_9495);
xnor U10172 (N_10172,N_9647,N_9340);
xnor U10173 (N_10173,N_9312,N_9242);
xor U10174 (N_10174,N_9171,N_9633);
and U10175 (N_10175,N_9973,N_9588);
nand U10176 (N_10176,N_9464,N_9505);
xor U10177 (N_10177,N_9490,N_9966);
or U10178 (N_10178,N_9914,N_9997);
or U10179 (N_10179,N_9247,N_9140);
nor U10180 (N_10180,N_9375,N_9848);
nor U10181 (N_10181,N_9897,N_9696);
xor U10182 (N_10182,N_9425,N_9792);
nor U10183 (N_10183,N_9717,N_9420);
or U10184 (N_10184,N_9178,N_9856);
xor U10185 (N_10185,N_9748,N_9751);
nor U10186 (N_10186,N_9770,N_9485);
or U10187 (N_10187,N_9153,N_9166);
nand U10188 (N_10188,N_9116,N_9443);
xor U10189 (N_10189,N_9985,N_9083);
xnor U10190 (N_10190,N_9168,N_9306);
xor U10191 (N_10191,N_9141,N_9249);
or U10192 (N_10192,N_9144,N_9093);
nand U10193 (N_10193,N_9003,N_9903);
xor U10194 (N_10194,N_9253,N_9707);
or U10195 (N_10195,N_9295,N_9009);
nand U10196 (N_10196,N_9380,N_9972);
nor U10197 (N_10197,N_9989,N_9695);
xor U10198 (N_10198,N_9646,N_9435);
nor U10199 (N_10199,N_9825,N_9548);
and U10200 (N_10200,N_9970,N_9731);
nor U10201 (N_10201,N_9534,N_9978);
and U10202 (N_10202,N_9390,N_9103);
or U10203 (N_10203,N_9201,N_9193);
or U10204 (N_10204,N_9569,N_9332);
nor U10205 (N_10205,N_9208,N_9250);
or U10206 (N_10206,N_9761,N_9651);
nor U10207 (N_10207,N_9593,N_9636);
nor U10208 (N_10208,N_9486,N_9920);
xor U10209 (N_10209,N_9776,N_9355);
xnor U10210 (N_10210,N_9913,N_9667);
nand U10211 (N_10211,N_9849,N_9710);
nand U10212 (N_10212,N_9931,N_9285);
or U10213 (N_10213,N_9266,N_9591);
nand U10214 (N_10214,N_9572,N_9112);
or U10215 (N_10215,N_9400,N_9728);
nand U10216 (N_10216,N_9013,N_9337);
and U10217 (N_10217,N_9449,N_9224);
nor U10218 (N_10218,N_9808,N_9793);
nor U10219 (N_10219,N_9619,N_9703);
or U10220 (N_10220,N_9367,N_9403);
nand U10221 (N_10221,N_9592,N_9305);
xor U10222 (N_10222,N_9672,N_9738);
and U10223 (N_10223,N_9900,N_9476);
nand U10224 (N_10224,N_9500,N_9945);
and U10225 (N_10225,N_9074,N_9283);
and U10226 (N_10226,N_9026,N_9299);
nand U10227 (N_10227,N_9754,N_9128);
or U10228 (N_10228,N_9839,N_9957);
and U10229 (N_10229,N_9329,N_9197);
nand U10230 (N_10230,N_9391,N_9876);
nor U10231 (N_10231,N_9450,N_9040);
or U10232 (N_10232,N_9740,N_9940);
nor U10233 (N_10233,N_9585,N_9524);
and U10234 (N_10234,N_9225,N_9615);
or U10235 (N_10235,N_9649,N_9919);
and U10236 (N_10236,N_9254,N_9601);
or U10237 (N_10237,N_9336,N_9124);
xor U10238 (N_10238,N_9094,N_9043);
and U10239 (N_10239,N_9192,N_9260);
nor U10240 (N_10240,N_9131,N_9772);
nor U10241 (N_10241,N_9474,N_9297);
nor U10242 (N_10242,N_9164,N_9824);
nor U10243 (N_10243,N_9701,N_9630);
nor U10244 (N_10244,N_9813,N_9705);
xnor U10245 (N_10245,N_9183,N_9652);
or U10246 (N_10246,N_9958,N_9516);
or U10247 (N_10247,N_9542,N_9342);
nand U10248 (N_10248,N_9933,N_9475);
nand U10249 (N_10249,N_9846,N_9335);
or U10250 (N_10250,N_9943,N_9659);
nor U10251 (N_10251,N_9538,N_9827);
nor U10252 (N_10252,N_9111,N_9017);
and U10253 (N_10253,N_9235,N_9785);
and U10254 (N_10254,N_9440,N_9368);
and U10255 (N_10255,N_9001,N_9983);
nor U10256 (N_10256,N_9893,N_9700);
nand U10257 (N_10257,N_9082,N_9268);
nand U10258 (N_10258,N_9053,N_9142);
nand U10259 (N_10259,N_9263,N_9668);
nand U10260 (N_10260,N_9523,N_9264);
nor U10261 (N_10261,N_9227,N_9816);
and U10262 (N_10262,N_9926,N_9993);
and U10263 (N_10263,N_9095,N_9862);
or U10264 (N_10264,N_9035,N_9868);
nor U10265 (N_10265,N_9730,N_9645);
nor U10266 (N_10266,N_9820,N_9145);
xnor U10267 (N_10267,N_9952,N_9456);
xnor U10268 (N_10268,N_9654,N_9759);
xnor U10269 (N_10269,N_9960,N_9853);
and U10270 (N_10270,N_9962,N_9965);
xor U10271 (N_10271,N_9613,N_9309);
or U10272 (N_10272,N_9558,N_9564);
or U10273 (N_10273,N_9898,N_9167);
nand U10274 (N_10274,N_9155,N_9096);
and U10275 (N_10275,N_9331,N_9108);
and U10276 (N_10276,N_9388,N_9418);
and U10277 (N_10277,N_9471,N_9553);
xor U10278 (N_10278,N_9277,N_9430);
and U10279 (N_10279,N_9198,N_9135);
nand U10280 (N_10280,N_9679,N_9330);
xor U10281 (N_10281,N_9088,N_9828);
and U10282 (N_10282,N_9422,N_9402);
xor U10283 (N_10283,N_9369,N_9323);
nor U10284 (N_10284,N_9489,N_9214);
xnor U10285 (N_10285,N_9195,N_9510);
nor U10286 (N_10286,N_9755,N_9326);
xor U10287 (N_10287,N_9508,N_9999);
nand U10288 (N_10288,N_9308,N_9097);
or U10289 (N_10289,N_9870,N_9018);
and U10290 (N_10290,N_9216,N_9842);
and U10291 (N_10291,N_9982,N_9520);
or U10292 (N_10292,N_9007,N_9327);
nand U10293 (N_10293,N_9536,N_9895);
nand U10294 (N_10294,N_9280,N_9143);
nand U10295 (N_10295,N_9582,N_9303);
nand U10296 (N_10296,N_9888,N_9934);
and U10297 (N_10297,N_9020,N_9511);
xor U10298 (N_10298,N_9803,N_9006);
xnor U10299 (N_10299,N_9530,N_9494);
and U10300 (N_10300,N_9032,N_9603);
xor U10301 (N_10301,N_9697,N_9955);
xnor U10302 (N_10302,N_9874,N_9324);
xnor U10303 (N_10303,N_9328,N_9052);
and U10304 (N_10304,N_9455,N_9258);
xor U10305 (N_10305,N_9680,N_9243);
nand U10306 (N_10306,N_9867,N_9194);
or U10307 (N_10307,N_9750,N_9496);
or U10308 (N_10308,N_9676,N_9799);
nor U10309 (N_10309,N_9595,N_9624);
nand U10310 (N_10310,N_9691,N_9871);
and U10311 (N_10311,N_9515,N_9718);
xor U10312 (N_10312,N_9573,N_9107);
nor U10313 (N_10313,N_9011,N_9267);
and U10314 (N_10314,N_9259,N_9805);
nand U10315 (N_10315,N_9773,N_9360);
xnor U10316 (N_10316,N_9971,N_9492);
nand U10317 (N_10317,N_9915,N_9325);
nor U10318 (N_10318,N_9579,N_9057);
nor U10319 (N_10319,N_9838,N_9466);
or U10320 (N_10320,N_9764,N_9311);
or U10321 (N_10321,N_9563,N_9843);
and U10322 (N_10322,N_9789,N_9479);
nor U10323 (N_10323,N_9015,N_9852);
and U10324 (N_10324,N_9540,N_9460);
and U10325 (N_10325,N_9678,N_9872);
nor U10326 (N_10326,N_9719,N_9533);
nand U10327 (N_10327,N_9784,N_9996);
xnor U10328 (N_10328,N_9042,N_9105);
or U10329 (N_10329,N_9386,N_9181);
or U10330 (N_10330,N_9457,N_9139);
or U10331 (N_10331,N_9272,N_9566);
xnor U10332 (N_10332,N_9341,N_9207);
nor U10333 (N_10333,N_9628,N_9359);
nand U10334 (N_10334,N_9546,N_9373);
nand U10335 (N_10335,N_9606,N_9477);
xor U10336 (N_10336,N_9357,N_9045);
and U10337 (N_10337,N_9289,N_9513);
nor U10338 (N_10338,N_9115,N_9010);
and U10339 (N_10339,N_9640,N_9237);
or U10340 (N_10340,N_9016,N_9988);
xnor U10341 (N_10341,N_9334,N_9774);
or U10342 (N_10342,N_9879,N_9256);
and U10343 (N_10343,N_9113,N_9638);
and U10344 (N_10344,N_9274,N_9684);
or U10345 (N_10345,N_9835,N_9446);
or U10346 (N_10346,N_9269,N_9768);
nand U10347 (N_10347,N_9130,N_9067);
nand U10348 (N_10348,N_9186,N_9230);
nor U10349 (N_10349,N_9445,N_9798);
xor U10350 (N_10350,N_9424,N_9050);
nor U10351 (N_10351,N_9639,N_9321);
and U10352 (N_10352,N_9611,N_9656);
nor U10353 (N_10353,N_9436,N_9286);
nand U10354 (N_10354,N_9199,N_9840);
nor U10355 (N_10355,N_9431,N_9377);
or U10356 (N_10356,N_9912,N_9092);
and U10357 (N_10357,N_9120,N_9315);
and U10358 (N_10358,N_9385,N_9599);
and U10359 (N_10359,N_9356,N_9414);
nor U10360 (N_10360,N_9075,N_9428);
xnor U10361 (N_10361,N_9383,N_9735);
nor U10362 (N_10362,N_9949,N_9149);
and U10363 (N_10363,N_9273,N_9169);
nor U10364 (N_10364,N_9709,N_9623);
xnor U10365 (N_10365,N_9597,N_9502);
xnor U10366 (N_10366,N_9288,N_9685);
or U10367 (N_10367,N_9014,N_9532);
or U10368 (N_10368,N_9118,N_9370);
and U10369 (N_10369,N_9404,N_9561);
xor U10370 (N_10370,N_9233,N_9392);
nand U10371 (N_10371,N_9226,N_9743);
nor U10372 (N_10372,N_9172,N_9644);
or U10373 (N_10373,N_9702,N_9338);
and U10374 (N_10374,N_9917,N_9954);
nand U10375 (N_10375,N_9426,N_9858);
or U10376 (N_10376,N_9047,N_9405);
nor U10377 (N_10377,N_9987,N_9123);
nand U10378 (N_10378,N_9176,N_9767);
or U10379 (N_10379,N_9023,N_9317);
xnor U10380 (N_10380,N_9248,N_9398);
and U10381 (N_10381,N_9762,N_9739);
and U10382 (N_10382,N_9560,N_9889);
and U10383 (N_10383,N_9617,N_9526);
nand U10384 (N_10384,N_9177,N_9594);
nand U10385 (N_10385,N_9512,N_9733);
and U10386 (N_10386,N_9322,N_9284);
or U10387 (N_10387,N_9498,N_9162);
and U10388 (N_10388,N_9905,N_9378);
xnor U10389 (N_10389,N_9046,N_9098);
nand U10390 (N_10390,N_9964,N_9210);
or U10391 (N_10391,N_9899,N_9786);
or U10392 (N_10392,N_9880,N_9491);
or U10393 (N_10393,N_9497,N_9746);
nor U10394 (N_10394,N_9584,N_9127);
or U10395 (N_10395,N_9302,N_9929);
xnor U10396 (N_10396,N_9833,N_9711);
nor U10397 (N_10397,N_9352,N_9545);
and U10398 (N_10398,N_9749,N_9722);
nor U10399 (N_10399,N_9723,N_9129);
nand U10400 (N_10400,N_9675,N_9932);
xnor U10401 (N_10401,N_9160,N_9892);
or U10402 (N_10402,N_9851,N_9379);
nand U10403 (N_10403,N_9634,N_9896);
xor U10404 (N_10404,N_9947,N_9557);
or U10405 (N_10405,N_9408,N_9252);
or U10406 (N_10406,N_9223,N_9963);
nor U10407 (N_10407,N_9747,N_9866);
or U10408 (N_10408,N_9161,N_9421);
nand U10409 (N_10409,N_9643,N_9791);
nand U10410 (N_10410,N_9807,N_9830);
nor U10411 (N_10411,N_9278,N_9232);
xor U10412 (N_10412,N_9066,N_9483);
nor U10413 (N_10413,N_9525,N_9686);
nor U10414 (N_10414,N_9812,N_9433);
xnor U10415 (N_10415,N_9058,N_9203);
nor U10416 (N_10416,N_9076,N_9451);
nor U10417 (N_10417,N_9343,N_9069);
nor U10418 (N_10418,N_9117,N_9211);
and U10419 (N_10419,N_9976,N_9209);
nor U10420 (N_10420,N_9204,N_9202);
or U10421 (N_10421,N_9038,N_9245);
or U10422 (N_10422,N_9596,N_9618);
or U10423 (N_10423,N_9397,N_9559);
nor U10424 (N_10424,N_9462,N_9364);
or U10425 (N_10425,N_9655,N_9366);
nor U10426 (N_10426,N_9698,N_9358);
nand U10427 (N_10427,N_9670,N_9690);
or U10428 (N_10428,N_9362,N_9432);
nand U10429 (N_10429,N_9959,N_9068);
xnor U10430 (N_10430,N_9220,N_9215);
nor U10431 (N_10431,N_9291,N_9307);
xor U10432 (N_10432,N_9797,N_9550);
nor U10433 (N_10433,N_9298,N_9908);
nor U10434 (N_10434,N_9241,N_9736);
nand U10435 (N_10435,N_9683,N_9766);
xor U10436 (N_10436,N_9788,N_9881);
xnor U10437 (N_10437,N_9737,N_9831);
and U10438 (N_10438,N_9517,N_9554);
nor U10439 (N_10439,N_9387,N_9715);
or U10440 (N_10440,N_9854,N_9078);
nand U10441 (N_10441,N_9577,N_9901);
and U10442 (N_10442,N_9154,N_9350);
or U10443 (N_10443,N_9348,N_9079);
xnor U10444 (N_10444,N_9191,N_9706);
nor U10445 (N_10445,N_9794,N_9104);
nand U10446 (N_10446,N_9522,N_9228);
and U10447 (N_10447,N_9631,N_9133);
xor U10448 (N_10448,N_9504,N_9503);
xor U10449 (N_10449,N_9170,N_9393);
nand U10450 (N_10450,N_9657,N_9396);
nor U10451 (N_10451,N_9231,N_9666);
or U10452 (N_10452,N_9765,N_9821);
nand U10453 (N_10453,N_9551,N_9345);
xnor U10454 (N_10454,N_9429,N_9319);
xnor U10455 (N_10455,N_9616,N_9834);
xnor U10456 (N_10456,N_9381,N_9158);
xnor U10457 (N_10457,N_9909,N_9745);
nand U10458 (N_10458,N_9861,N_9461);
xnor U10459 (N_10459,N_9694,N_9005);
xnor U10460 (N_10460,N_9725,N_9927);
or U10461 (N_10461,N_9802,N_9109);
or U10462 (N_10462,N_9044,N_9255);
nor U10463 (N_10463,N_9401,N_9339);
nand U10464 (N_10464,N_9219,N_9674);
or U10465 (N_10465,N_9884,N_9024);
nand U10466 (N_10466,N_9916,N_9363);
nor U10467 (N_10467,N_9296,N_9441);
nand U10468 (N_10468,N_9637,N_9200);
nor U10469 (N_10469,N_9859,N_9600);
xor U10470 (N_10470,N_9894,N_9673);
xor U10471 (N_10471,N_9072,N_9689);
and U10472 (N_10472,N_9907,N_9576);
or U10473 (N_10473,N_9061,N_9060);
nor U10474 (N_10474,N_9544,N_9238);
nor U10475 (N_10475,N_9575,N_9478);
or U10476 (N_10476,N_9275,N_9586);
and U10477 (N_10477,N_9906,N_9681);
xnor U10478 (N_10478,N_9134,N_9650);
or U10479 (N_10479,N_9890,N_9301);
or U10480 (N_10480,N_9662,N_9811);
and U10481 (N_10481,N_9682,N_9179);
or U10482 (N_10482,N_9753,N_9292);
and U10483 (N_10483,N_9992,N_9240);
or U10484 (N_10484,N_9543,N_9688);
and U10485 (N_10485,N_9051,N_9313);
nand U10486 (N_10486,N_9213,N_9734);
xnor U10487 (N_10487,N_9089,N_9911);
or U10488 (N_10488,N_9188,N_9506);
nor U10489 (N_10489,N_9039,N_9085);
xnor U10490 (N_10490,N_9991,N_9938);
nor U10491 (N_10491,N_9374,N_9423);
nor U10492 (N_10492,N_9625,N_9968);
or U10493 (N_10493,N_9887,N_9468);
or U10494 (N_10494,N_9568,N_9257);
and U10495 (N_10495,N_9771,N_9270);
nor U10496 (N_10496,N_9065,N_9537);
nor U10497 (N_10497,N_9316,N_9819);
nor U10498 (N_10498,N_9122,N_9481);
nand U10499 (N_10499,N_9439,N_9086);
nand U10500 (N_10500,N_9715,N_9591);
or U10501 (N_10501,N_9736,N_9452);
nor U10502 (N_10502,N_9320,N_9361);
and U10503 (N_10503,N_9873,N_9289);
or U10504 (N_10504,N_9344,N_9386);
nor U10505 (N_10505,N_9199,N_9188);
and U10506 (N_10506,N_9315,N_9933);
nor U10507 (N_10507,N_9367,N_9122);
xnor U10508 (N_10508,N_9502,N_9254);
and U10509 (N_10509,N_9749,N_9361);
and U10510 (N_10510,N_9276,N_9741);
or U10511 (N_10511,N_9901,N_9799);
nor U10512 (N_10512,N_9489,N_9671);
and U10513 (N_10513,N_9332,N_9942);
and U10514 (N_10514,N_9177,N_9807);
and U10515 (N_10515,N_9117,N_9194);
nand U10516 (N_10516,N_9998,N_9714);
nand U10517 (N_10517,N_9222,N_9397);
nand U10518 (N_10518,N_9446,N_9863);
nor U10519 (N_10519,N_9181,N_9275);
nand U10520 (N_10520,N_9268,N_9753);
and U10521 (N_10521,N_9706,N_9001);
nand U10522 (N_10522,N_9452,N_9116);
xnor U10523 (N_10523,N_9807,N_9220);
nor U10524 (N_10524,N_9087,N_9692);
or U10525 (N_10525,N_9962,N_9339);
nor U10526 (N_10526,N_9832,N_9684);
and U10527 (N_10527,N_9212,N_9728);
or U10528 (N_10528,N_9663,N_9335);
nor U10529 (N_10529,N_9740,N_9422);
xor U10530 (N_10530,N_9492,N_9735);
nor U10531 (N_10531,N_9991,N_9752);
nand U10532 (N_10532,N_9832,N_9628);
or U10533 (N_10533,N_9852,N_9148);
nor U10534 (N_10534,N_9595,N_9011);
nand U10535 (N_10535,N_9031,N_9028);
nand U10536 (N_10536,N_9673,N_9796);
nor U10537 (N_10537,N_9103,N_9870);
xor U10538 (N_10538,N_9236,N_9314);
nand U10539 (N_10539,N_9025,N_9760);
xnor U10540 (N_10540,N_9767,N_9485);
and U10541 (N_10541,N_9945,N_9609);
and U10542 (N_10542,N_9111,N_9471);
xor U10543 (N_10543,N_9896,N_9727);
and U10544 (N_10544,N_9404,N_9958);
nand U10545 (N_10545,N_9259,N_9563);
nor U10546 (N_10546,N_9120,N_9132);
xor U10547 (N_10547,N_9071,N_9133);
nand U10548 (N_10548,N_9832,N_9836);
nand U10549 (N_10549,N_9636,N_9311);
nor U10550 (N_10550,N_9318,N_9964);
nor U10551 (N_10551,N_9988,N_9082);
and U10552 (N_10552,N_9153,N_9242);
or U10553 (N_10553,N_9178,N_9525);
nand U10554 (N_10554,N_9586,N_9844);
nand U10555 (N_10555,N_9272,N_9109);
nor U10556 (N_10556,N_9369,N_9482);
xnor U10557 (N_10557,N_9935,N_9134);
nor U10558 (N_10558,N_9694,N_9733);
or U10559 (N_10559,N_9509,N_9905);
xnor U10560 (N_10560,N_9247,N_9098);
or U10561 (N_10561,N_9295,N_9429);
or U10562 (N_10562,N_9436,N_9780);
and U10563 (N_10563,N_9105,N_9395);
nor U10564 (N_10564,N_9573,N_9344);
nand U10565 (N_10565,N_9371,N_9235);
nor U10566 (N_10566,N_9026,N_9758);
or U10567 (N_10567,N_9123,N_9594);
and U10568 (N_10568,N_9342,N_9169);
and U10569 (N_10569,N_9541,N_9608);
or U10570 (N_10570,N_9332,N_9730);
nand U10571 (N_10571,N_9817,N_9289);
nor U10572 (N_10572,N_9507,N_9340);
nor U10573 (N_10573,N_9549,N_9841);
nor U10574 (N_10574,N_9180,N_9855);
xnor U10575 (N_10575,N_9678,N_9895);
nor U10576 (N_10576,N_9326,N_9559);
xnor U10577 (N_10577,N_9947,N_9414);
xor U10578 (N_10578,N_9042,N_9632);
or U10579 (N_10579,N_9264,N_9881);
and U10580 (N_10580,N_9991,N_9370);
nor U10581 (N_10581,N_9949,N_9202);
nor U10582 (N_10582,N_9235,N_9746);
nor U10583 (N_10583,N_9605,N_9097);
nor U10584 (N_10584,N_9032,N_9012);
nand U10585 (N_10585,N_9416,N_9145);
xor U10586 (N_10586,N_9307,N_9145);
nor U10587 (N_10587,N_9119,N_9193);
nand U10588 (N_10588,N_9980,N_9213);
and U10589 (N_10589,N_9895,N_9403);
xnor U10590 (N_10590,N_9136,N_9240);
and U10591 (N_10591,N_9905,N_9422);
xor U10592 (N_10592,N_9647,N_9184);
nor U10593 (N_10593,N_9744,N_9510);
nand U10594 (N_10594,N_9505,N_9307);
nor U10595 (N_10595,N_9398,N_9350);
xnor U10596 (N_10596,N_9914,N_9200);
xor U10597 (N_10597,N_9079,N_9724);
nand U10598 (N_10598,N_9887,N_9546);
and U10599 (N_10599,N_9202,N_9258);
xor U10600 (N_10600,N_9569,N_9924);
and U10601 (N_10601,N_9974,N_9819);
nor U10602 (N_10602,N_9276,N_9817);
xnor U10603 (N_10603,N_9370,N_9096);
nand U10604 (N_10604,N_9519,N_9238);
nand U10605 (N_10605,N_9026,N_9837);
or U10606 (N_10606,N_9069,N_9475);
or U10607 (N_10607,N_9732,N_9649);
and U10608 (N_10608,N_9952,N_9906);
nand U10609 (N_10609,N_9893,N_9940);
or U10610 (N_10610,N_9247,N_9751);
nor U10611 (N_10611,N_9894,N_9476);
nor U10612 (N_10612,N_9104,N_9159);
or U10613 (N_10613,N_9593,N_9322);
nand U10614 (N_10614,N_9812,N_9757);
xnor U10615 (N_10615,N_9286,N_9895);
and U10616 (N_10616,N_9101,N_9864);
or U10617 (N_10617,N_9338,N_9561);
nand U10618 (N_10618,N_9709,N_9376);
or U10619 (N_10619,N_9319,N_9548);
nand U10620 (N_10620,N_9849,N_9679);
or U10621 (N_10621,N_9540,N_9929);
nand U10622 (N_10622,N_9128,N_9657);
nand U10623 (N_10623,N_9320,N_9918);
nand U10624 (N_10624,N_9460,N_9263);
nand U10625 (N_10625,N_9927,N_9643);
xnor U10626 (N_10626,N_9621,N_9892);
xor U10627 (N_10627,N_9959,N_9957);
xnor U10628 (N_10628,N_9455,N_9636);
and U10629 (N_10629,N_9547,N_9125);
and U10630 (N_10630,N_9340,N_9911);
nand U10631 (N_10631,N_9414,N_9326);
nand U10632 (N_10632,N_9676,N_9430);
nand U10633 (N_10633,N_9514,N_9232);
and U10634 (N_10634,N_9182,N_9769);
nor U10635 (N_10635,N_9778,N_9766);
nor U10636 (N_10636,N_9549,N_9468);
nor U10637 (N_10637,N_9881,N_9774);
xnor U10638 (N_10638,N_9059,N_9067);
xnor U10639 (N_10639,N_9390,N_9379);
nand U10640 (N_10640,N_9727,N_9072);
xor U10641 (N_10641,N_9503,N_9669);
nor U10642 (N_10642,N_9067,N_9742);
nand U10643 (N_10643,N_9663,N_9651);
or U10644 (N_10644,N_9159,N_9846);
nor U10645 (N_10645,N_9813,N_9533);
nand U10646 (N_10646,N_9146,N_9478);
and U10647 (N_10647,N_9074,N_9610);
nand U10648 (N_10648,N_9658,N_9076);
and U10649 (N_10649,N_9979,N_9989);
and U10650 (N_10650,N_9153,N_9351);
nand U10651 (N_10651,N_9611,N_9644);
nor U10652 (N_10652,N_9882,N_9115);
or U10653 (N_10653,N_9564,N_9808);
nor U10654 (N_10654,N_9481,N_9739);
nand U10655 (N_10655,N_9644,N_9683);
nand U10656 (N_10656,N_9661,N_9995);
nand U10657 (N_10657,N_9603,N_9189);
and U10658 (N_10658,N_9686,N_9058);
and U10659 (N_10659,N_9268,N_9712);
or U10660 (N_10660,N_9773,N_9532);
or U10661 (N_10661,N_9359,N_9052);
and U10662 (N_10662,N_9768,N_9548);
nor U10663 (N_10663,N_9950,N_9981);
and U10664 (N_10664,N_9127,N_9291);
xnor U10665 (N_10665,N_9781,N_9595);
and U10666 (N_10666,N_9916,N_9753);
or U10667 (N_10667,N_9482,N_9257);
nor U10668 (N_10668,N_9998,N_9834);
and U10669 (N_10669,N_9437,N_9662);
nand U10670 (N_10670,N_9715,N_9140);
nand U10671 (N_10671,N_9190,N_9820);
or U10672 (N_10672,N_9247,N_9422);
or U10673 (N_10673,N_9480,N_9262);
or U10674 (N_10674,N_9473,N_9689);
nand U10675 (N_10675,N_9330,N_9860);
xor U10676 (N_10676,N_9064,N_9184);
nand U10677 (N_10677,N_9153,N_9275);
or U10678 (N_10678,N_9224,N_9809);
nor U10679 (N_10679,N_9886,N_9797);
and U10680 (N_10680,N_9221,N_9835);
or U10681 (N_10681,N_9628,N_9960);
or U10682 (N_10682,N_9559,N_9525);
xnor U10683 (N_10683,N_9510,N_9039);
and U10684 (N_10684,N_9253,N_9079);
or U10685 (N_10685,N_9590,N_9118);
or U10686 (N_10686,N_9251,N_9421);
nand U10687 (N_10687,N_9571,N_9739);
and U10688 (N_10688,N_9696,N_9145);
and U10689 (N_10689,N_9825,N_9044);
nand U10690 (N_10690,N_9152,N_9829);
or U10691 (N_10691,N_9789,N_9821);
nor U10692 (N_10692,N_9916,N_9991);
and U10693 (N_10693,N_9665,N_9379);
and U10694 (N_10694,N_9166,N_9488);
nor U10695 (N_10695,N_9185,N_9933);
nor U10696 (N_10696,N_9343,N_9799);
and U10697 (N_10697,N_9804,N_9291);
nor U10698 (N_10698,N_9980,N_9753);
or U10699 (N_10699,N_9978,N_9975);
xnor U10700 (N_10700,N_9121,N_9053);
and U10701 (N_10701,N_9897,N_9369);
and U10702 (N_10702,N_9674,N_9569);
xor U10703 (N_10703,N_9494,N_9597);
nor U10704 (N_10704,N_9581,N_9979);
or U10705 (N_10705,N_9898,N_9668);
nor U10706 (N_10706,N_9083,N_9635);
nor U10707 (N_10707,N_9427,N_9173);
or U10708 (N_10708,N_9265,N_9453);
or U10709 (N_10709,N_9476,N_9668);
nor U10710 (N_10710,N_9760,N_9858);
xnor U10711 (N_10711,N_9129,N_9442);
and U10712 (N_10712,N_9474,N_9227);
and U10713 (N_10713,N_9766,N_9135);
and U10714 (N_10714,N_9155,N_9433);
nand U10715 (N_10715,N_9201,N_9994);
and U10716 (N_10716,N_9118,N_9834);
and U10717 (N_10717,N_9730,N_9506);
xor U10718 (N_10718,N_9662,N_9312);
and U10719 (N_10719,N_9174,N_9830);
and U10720 (N_10720,N_9951,N_9131);
nand U10721 (N_10721,N_9645,N_9021);
nor U10722 (N_10722,N_9012,N_9159);
nor U10723 (N_10723,N_9187,N_9001);
nand U10724 (N_10724,N_9459,N_9226);
or U10725 (N_10725,N_9110,N_9748);
nand U10726 (N_10726,N_9778,N_9943);
xor U10727 (N_10727,N_9845,N_9397);
nor U10728 (N_10728,N_9174,N_9531);
or U10729 (N_10729,N_9777,N_9463);
nor U10730 (N_10730,N_9090,N_9193);
nor U10731 (N_10731,N_9401,N_9379);
or U10732 (N_10732,N_9425,N_9467);
and U10733 (N_10733,N_9542,N_9245);
nand U10734 (N_10734,N_9850,N_9353);
and U10735 (N_10735,N_9999,N_9930);
nor U10736 (N_10736,N_9137,N_9951);
nor U10737 (N_10737,N_9964,N_9469);
nor U10738 (N_10738,N_9867,N_9503);
nand U10739 (N_10739,N_9435,N_9377);
nor U10740 (N_10740,N_9362,N_9475);
or U10741 (N_10741,N_9155,N_9700);
xnor U10742 (N_10742,N_9904,N_9571);
and U10743 (N_10743,N_9429,N_9767);
and U10744 (N_10744,N_9654,N_9777);
xnor U10745 (N_10745,N_9133,N_9823);
nand U10746 (N_10746,N_9553,N_9232);
nor U10747 (N_10747,N_9604,N_9748);
nor U10748 (N_10748,N_9323,N_9931);
nand U10749 (N_10749,N_9974,N_9567);
xor U10750 (N_10750,N_9422,N_9643);
xnor U10751 (N_10751,N_9817,N_9446);
xor U10752 (N_10752,N_9950,N_9852);
nand U10753 (N_10753,N_9265,N_9201);
nor U10754 (N_10754,N_9083,N_9155);
nor U10755 (N_10755,N_9280,N_9124);
xor U10756 (N_10756,N_9528,N_9770);
xnor U10757 (N_10757,N_9397,N_9624);
nor U10758 (N_10758,N_9569,N_9603);
nand U10759 (N_10759,N_9828,N_9599);
xnor U10760 (N_10760,N_9604,N_9149);
nor U10761 (N_10761,N_9204,N_9224);
and U10762 (N_10762,N_9771,N_9943);
xnor U10763 (N_10763,N_9425,N_9056);
xor U10764 (N_10764,N_9132,N_9842);
nand U10765 (N_10765,N_9398,N_9925);
xnor U10766 (N_10766,N_9782,N_9163);
nor U10767 (N_10767,N_9726,N_9700);
xnor U10768 (N_10768,N_9668,N_9436);
or U10769 (N_10769,N_9350,N_9152);
and U10770 (N_10770,N_9677,N_9726);
nor U10771 (N_10771,N_9129,N_9703);
xnor U10772 (N_10772,N_9566,N_9867);
xnor U10773 (N_10773,N_9962,N_9017);
and U10774 (N_10774,N_9257,N_9977);
and U10775 (N_10775,N_9589,N_9208);
nand U10776 (N_10776,N_9421,N_9794);
and U10777 (N_10777,N_9670,N_9803);
nand U10778 (N_10778,N_9023,N_9385);
or U10779 (N_10779,N_9653,N_9910);
nand U10780 (N_10780,N_9578,N_9518);
or U10781 (N_10781,N_9923,N_9727);
or U10782 (N_10782,N_9002,N_9908);
xnor U10783 (N_10783,N_9116,N_9985);
xnor U10784 (N_10784,N_9097,N_9307);
nand U10785 (N_10785,N_9077,N_9414);
nand U10786 (N_10786,N_9940,N_9706);
or U10787 (N_10787,N_9532,N_9316);
or U10788 (N_10788,N_9336,N_9140);
nand U10789 (N_10789,N_9347,N_9881);
or U10790 (N_10790,N_9551,N_9377);
nand U10791 (N_10791,N_9187,N_9503);
or U10792 (N_10792,N_9902,N_9258);
nor U10793 (N_10793,N_9481,N_9366);
nand U10794 (N_10794,N_9874,N_9047);
nor U10795 (N_10795,N_9079,N_9847);
nand U10796 (N_10796,N_9114,N_9954);
nor U10797 (N_10797,N_9950,N_9681);
xnor U10798 (N_10798,N_9170,N_9502);
nor U10799 (N_10799,N_9005,N_9212);
xnor U10800 (N_10800,N_9635,N_9170);
xnor U10801 (N_10801,N_9230,N_9407);
nor U10802 (N_10802,N_9007,N_9916);
nand U10803 (N_10803,N_9174,N_9610);
nor U10804 (N_10804,N_9601,N_9080);
nand U10805 (N_10805,N_9989,N_9211);
xnor U10806 (N_10806,N_9207,N_9050);
nor U10807 (N_10807,N_9475,N_9229);
xnor U10808 (N_10808,N_9077,N_9574);
nor U10809 (N_10809,N_9051,N_9977);
nand U10810 (N_10810,N_9293,N_9168);
and U10811 (N_10811,N_9160,N_9316);
nor U10812 (N_10812,N_9774,N_9191);
nand U10813 (N_10813,N_9376,N_9726);
xor U10814 (N_10814,N_9075,N_9395);
and U10815 (N_10815,N_9312,N_9299);
nor U10816 (N_10816,N_9109,N_9490);
xor U10817 (N_10817,N_9651,N_9174);
xnor U10818 (N_10818,N_9981,N_9149);
nor U10819 (N_10819,N_9749,N_9740);
nand U10820 (N_10820,N_9108,N_9477);
xnor U10821 (N_10821,N_9949,N_9229);
or U10822 (N_10822,N_9732,N_9613);
xnor U10823 (N_10823,N_9256,N_9247);
xor U10824 (N_10824,N_9368,N_9920);
or U10825 (N_10825,N_9834,N_9748);
nand U10826 (N_10826,N_9430,N_9871);
nand U10827 (N_10827,N_9117,N_9060);
xor U10828 (N_10828,N_9973,N_9923);
nand U10829 (N_10829,N_9538,N_9599);
xnor U10830 (N_10830,N_9440,N_9238);
nor U10831 (N_10831,N_9165,N_9283);
nand U10832 (N_10832,N_9013,N_9474);
xnor U10833 (N_10833,N_9464,N_9402);
and U10834 (N_10834,N_9879,N_9358);
and U10835 (N_10835,N_9050,N_9101);
or U10836 (N_10836,N_9740,N_9451);
or U10837 (N_10837,N_9722,N_9170);
or U10838 (N_10838,N_9265,N_9830);
or U10839 (N_10839,N_9289,N_9029);
and U10840 (N_10840,N_9794,N_9704);
xnor U10841 (N_10841,N_9443,N_9091);
xor U10842 (N_10842,N_9851,N_9291);
or U10843 (N_10843,N_9442,N_9025);
xor U10844 (N_10844,N_9783,N_9761);
or U10845 (N_10845,N_9255,N_9121);
nor U10846 (N_10846,N_9072,N_9071);
or U10847 (N_10847,N_9378,N_9601);
or U10848 (N_10848,N_9297,N_9949);
or U10849 (N_10849,N_9800,N_9804);
nand U10850 (N_10850,N_9366,N_9457);
xor U10851 (N_10851,N_9937,N_9805);
or U10852 (N_10852,N_9608,N_9815);
and U10853 (N_10853,N_9776,N_9434);
and U10854 (N_10854,N_9213,N_9271);
nand U10855 (N_10855,N_9613,N_9920);
or U10856 (N_10856,N_9523,N_9260);
or U10857 (N_10857,N_9591,N_9262);
xor U10858 (N_10858,N_9573,N_9153);
nand U10859 (N_10859,N_9228,N_9452);
and U10860 (N_10860,N_9138,N_9292);
nor U10861 (N_10861,N_9213,N_9909);
nand U10862 (N_10862,N_9261,N_9524);
xnor U10863 (N_10863,N_9549,N_9402);
nand U10864 (N_10864,N_9784,N_9360);
xnor U10865 (N_10865,N_9631,N_9141);
nand U10866 (N_10866,N_9877,N_9239);
and U10867 (N_10867,N_9380,N_9644);
xor U10868 (N_10868,N_9886,N_9779);
nand U10869 (N_10869,N_9022,N_9543);
nand U10870 (N_10870,N_9273,N_9384);
nand U10871 (N_10871,N_9545,N_9437);
nand U10872 (N_10872,N_9244,N_9765);
or U10873 (N_10873,N_9693,N_9524);
nor U10874 (N_10874,N_9413,N_9244);
and U10875 (N_10875,N_9292,N_9116);
nor U10876 (N_10876,N_9093,N_9830);
xor U10877 (N_10877,N_9069,N_9245);
nor U10878 (N_10878,N_9985,N_9450);
nor U10879 (N_10879,N_9005,N_9999);
and U10880 (N_10880,N_9891,N_9935);
and U10881 (N_10881,N_9177,N_9140);
and U10882 (N_10882,N_9169,N_9732);
nand U10883 (N_10883,N_9851,N_9832);
nor U10884 (N_10884,N_9863,N_9155);
nor U10885 (N_10885,N_9471,N_9297);
and U10886 (N_10886,N_9088,N_9183);
or U10887 (N_10887,N_9630,N_9572);
xor U10888 (N_10888,N_9590,N_9233);
nand U10889 (N_10889,N_9398,N_9954);
or U10890 (N_10890,N_9257,N_9843);
nand U10891 (N_10891,N_9338,N_9649);
or U10892 (N_10892,N_9797,N_9026);
or U10893 (N_10893,N_9708,N_9478);
xnor U10894 (N_10894,N_9423,N_9411);
or U10895 (N_10895,N_9551,N_9727);
and U10896 (N_10896,N_9369,N_9314);
or U10897 (N_10897,N_9340,N_9152);
xnor U10898 (N_10898,N_9782,N_9697);
nand U10899 (N_10899,N_9101,N_9905);
xnor U10900 (N_10900,N_9885,N_9720);
xor U10901 (N_10901,N_9537,N_9117);
nor U10902 (N_10902,N_9038,N_9446);
xnor U10903 (N_10903,N_9080,N_9767);
xnor U10904 (N_10904,N_9324,N_9291);
nor U10905 (N_10905,N_9081,N_9396);
xor U10906 (N_10906,N_9993,N_9830);
xnor U10907 (N_10907,N_9267,N_9547);
and U10908 (N_10908,N_9957,N_9736);
nand U10909 (N_10909,N_9315,N_9775);
and U10910 (N_10910,N_9200,N_9688);
nor U10911 (N_10911,N_9995,N_9407);
or U10912 (N_10912,N_9432,N_9577);
nand U10913 (N_10913,N_9338,N_9113);
and U10914 (N_10914,N_9805,N_9736);
or U10915 (N_10915,N_9686,N_9913);
nand U10916 (N_10916,N_9408,N_9966);
or U10917 (N_10917,N_9911,N_9589);
nor U10918 (N_10918,N_9277,N_9623);
and U10919 (N_10919,N_9275,N_9478);
nand U10920 (N_10920,N_9776,N_9318);
nand U10921 (N_10921,N_9900,N_9025);
nand U10922 (N_10922,N_9102,N_9314);
and U10923 (N_10923,N_9371,N_9938);
and U10924 (N_10924,N_9764,N_9941);
and U10925 (N_10925,N_9365,N_9404);
nand U10926 (N_10926,N_9854,N_9884);
or U10927 (N_10927,N_9735,N_9942);
xnor U10928 (N_10928,N_9497,N_9028);
nor U10929 (N_10929,N_9778,N_9831);
nand U10930 (N_10930,N_9840,N_9672);
nand U10931 (N_10931,N_9336,N_9353);
and U10932 (N_10932,N_9190,N_9297);
nor U10933 (N_10933,N_9814,N_9964);
and U10934 (N_10934,N_9574,N_9646);
xnor U10935 (N_10935,N_9999,N_9461);
xnor U10936 (N_10936,N_9525,N_9779);
nor U10937 (N_10937,N_9643,N_9027);
xor U10938 (N_10938,N_9251,N_9511);
and U10939 (N_10939,N_9251,N_9452);
xnor U10940 (N_10940,N_9336,N_9900);
nor U10941 (N_10941,N_9681,N_9123);
or U10942 (N_10942,N_9111,N_9030);
xnor U10943 (N_10943,N_9323,N_9849);
nand U10944 (N_10944,N_9990,N_9185);
nand U10945 (N_10945,N_9930,N_9518);
xor U10946 (N_10946,N_9019,N_9239);
xnor U10947 (N_10947,N_9209,N_9711);
nand U10948 (N_10948,N_9276,N_9597);
and U10949 (N_10949,N_9670,N_9779);
nor U10950 (N_10950,N_9762,N_9168);
nor U10951 (N_10951,N_9932,N_9166);
or U10952 (N_10952,N_9816,N_9400);
and U10953 (N_10953,N_9240,N_9819);
or U10954 (N_10954,N_9578,N_9824);
nand U10955 (N_10955,N_9582,N_9091);
or U10956 (N_10956,N_9016,N_9408);
and U10957 (N_10957,N_9805,N_9664);
and U10958 (N_10958,N_9147,N_9615);
or U10959 (N_10959,N_9147,N_9636);
nand U10960 (N_10960,N_9511,N_9010);
xnor U10961 (N_10961,N_9540,N_9720);
and U10962 (N_10962,N_9919,N_9279);
or U10963 (N_10963,N_9709,N_9484);
nand U10964 (N_10964,N_9136,N_9758);
nand U10965 (N_10965,N_9504,N_9362);
nand U10966 (N_10966,N_9228,N_9955);
and U10967 (N_10967,N_9865,N_9366);
and U10968 (N_10968,N_9193,N_9837);
nand U10969 (N_10969,N_9199,N_9029);
or U10970 (N_10970,N_9250,N_9636);
nand U10971 (N_10971,N_9979,N_9544);
xor U10972 (N_10972,N_9612,N_9817);
nor U10973 (N_10973,N_9850,N_9231);
xnor U10974 (N_10974,N_9206,N_9176);
nand U10975 (N_10975,N_9342,N_9806);
or U10976 (N_10976,N_9004,N_9660);
nand U10977 (N_10977,N_9392,N_9521);
and U10978 (N_10978,N_9348,N_9155);
and U10979 (N_10979,N_9343,N_9847);
xnor U10980 (N_10980,N_9316,N_9931);
xnor U10981 (N_10981,N_9467,N_9595);
or U10982 (N_10982,N_9740,N_9604);
xor U10983 (N_10983,N_9805,N_9935);
xnor U10984 (N_10984,N_9472,N_9178);
or U10985 (N_10985,N_9589,N_9112);
xnor U10986 (N_10986,N_9818,N_9494);
xnor U10987 (N_10987,N_9959,N_9492);
and U10988 (N_10988,N_9075,N_9308);
nand U10989 (N_10989,N_9218,N_9326);
and U10990 (N_10990,N_9016,N_9721);
xor U10991 (N_10991,N_9238,N_9138);
or U10992 (N_10992,N_9351,N_9752);
or U10993 (N_10993,N_9342,N_9242);
nor U10994 (N_10994,N_9347,N_9208);
nand U10995 (N_10995,N_9603,N_9878);
xor U10996 (N_10996,N_9927,N_9887);
xnor U10997 (N_10997,N_9114,N_9228);
and U10998 (N_10998,N_9581,N_9584);
or U10999 (N_10999,N_9588,N_9077);
nor U11000 (N_11000,N_10565,N_10526);
or U11001 (N_11001,N_10627,N_10569);
xor U11002 (N_11002,N_10897,N_10820);
and U11003 (N_11003,N_10032,N_10338);
nand U11004 (N_11004,N_10872,N_10893);
and U11005 (N_11005,N_10774,N_10036);
xor U11006 (N_11006,N_10207,N_10388);
xnor U11007 (N_11007,N_10042,N_10723);
xnor U11008 (N_11008,N_10462,N_10489);
nor U11009 (N_11009,N_10266,N_10403);
nor U11010 (N_11010,N_10096,N_10621);
nand U11011 (N_11011,N_10105,N_10140);
nor U11012 (N_11012,N_10732,N_10878);
and U11013 (N_11013,N_10252,N_10260);
xor U11014 (N_11014,N_10862,N_10559);
xor U11015 (N_11015,N_10743,N_10496);
xor U11016 (N_11016,N_10104,N_10329);
xor U11017 (N_11017,N_10461,N_10320);
xor U11018 (N_11018,N_10106,N_10278);
nand U11019 (N_11019,N_10458,N_10024);
nand U11020 (N_11020,N_10999,N_10448);
nor U11021 (N_11021,N_10112,N_10285);
xnor U11022 (N_11022,N_10875,N_10865);
xor U11023 (N_11023,N_10275,N_10750);
xor U11024 (N_11024,N_10794,N_10988);
xor U11025 (N_11025,N_10372,N_10057);
nor U11026 (N_11026,N_10141,N_10836);
xor U11027 (N_11027,N_10188,N_10917);
nand U11028 (N_11028,N_10799,N_10321);
nand U11029 (N_11029,N_10305,N_10715);
or U11030 (N_11030,N_10068,N_10775);
nor U11031 (N_11031,N_10089,N_10813);
or U11032 (N_11032,N_10877,N_10229);
or U11033 (N_11033,N_10473,N_10707);
and U11034 (N_11034,N_10409,N_10322);
xnor U11035 (N_11035,N_10861,N_10198);
nor U11036 (N_11036,N_10664,N_10438);
or U11037 (N_11037,N_10401,N_10589);
nor U11038 (N_11038,N_10560,N_10746);
nand U11039 (N_11039,N_10588,N_10922);
or U11040 (N_11040,N_10823,N_10349);
and U11041 (N_11041,N_10725,N_10827);
xnor U11042 (N_11042,N_10779,N_10186);
and U11043 (N_11043,N_10471,N_10040);
nor U11044 (N_11044,N_10015,N_10716);
nor U11045 (N_11045,N_10478,N_10705);
nor U11046 (N_11046,N_10889,N_10689);
nor U11047 (N_11047,N_10181,N_10807);
or U11048 (N_11048,N_10619,N_10272);
nor U11049 (N_11049,N_10607,N_10671);
nor U11050 (N_11050,N_10702,N_10019);
nor U11051 (N_11051,N_10695,N_10751);
and U11052 (N_11052,N_10833,N_10916);
or U11053 (N_11053,N_10262,N_10302);
and U11054 (N_11054,N_10975,N_10578);
and U11055 (N_11055,N_10124,N_10282);
and U11056 (N_11056,N_10234,N_10626);
xor U11057 (N_11057,N_10356,N_10642);
or U11058 (N_11058,N_10789,N_10660);
nor U11059 (N_11059,N_10797,N_10668);
and U11060 (N_11060,N_10811,N_10687);
xnor U11061 (N_11061,N_10265,N_10097);
and U11062 (N_11062,N_10523,N_10939);
or U11063 (N_11063,N_10063,N_10784);
nand U11064 (N_11064,N_10834,N_10162);
nor U11065 (N_11065,N_10021,N_10263);
and U11066 (N_11066,N_10452,N_10955);
and U11067 (N_11067,N_10535,N_10371);
or U11068 (N_11068,N_10390,N_10859);
nor U11069 (N_11069,N_10787,N_10035);
nand U11070 (N_11070,N_10635,N_10481);
and U11071 (N_11071,N_10107,N_10798);
or U11072 (N_11072,N_10623,N_10638);
xnor U11073 (N_11073,N_10992,N_10968);
xor U11074 (N_11074,N_10056,N_10803);
nor U11075 (N_11075,N_10038,N_10914);
nor U11076 (N_11076,N_10700,N_10777);
nand U11077 (N_11077,N_10080,N_10355);
nor U11078 (N_11078,N_10210,N_10016);
xnor U11079 (N_11079,N_10520,N_10501);
nor U11080 (N_11080,N_10656,N_10271);
nor U11081 (N_11081,N_10896,N_10366);
or U11082 (N_11082,N_10413,N_10628);
and U11083 (N_11083,N_10394,N_10079);
and U11084 (N_11084,N_10555,N_10849);
nor U11085 (N_11085,N_10690,N_10201);
or U11086 (N_11086,N_10399,N_10256);
xnor U11087 (N_11087,N_10821,N_10518);
or U11088 (N_11088,N_10957,N_10945);
nand U11089 (N_11089,N_10749,N_10719);
nand U11090 (N_11090,N_10143,N_10611);
or U11091 (N_11091,N_10848,N_10146);
xor U11092 (N_11092,N_10236,N_10476);
nor U11093 (N_11093,N_10130,N_10450);
nor U11094 (N_11094,N_10013,N_10663);
and U11095 (N_11095,N_10582,N_10241);
nor U11096 (N_11096,N_10192,N_10088);
nor U11097 (N_11097,N_10453,N_10340);
or U11098 (N_11098,N_10730,N_10070);
or U11099 (N_11099,N_10752,N_10328);
xnor U11100 (N_11100,N_10362,N_10822);
nor U11101 (N_11101,N_10185,N_10944);
xnor U11102 (N_11102,N_10318,N_10864);
nand U11103 (N_11103,N_10091,N_10919);
nand U11104 (N_11104,N_10081,N_10658);
nand U11105 (N_11105,N_10326,N_10030);
and U11106 (N_11106,N_10243,N_10629);
xor U11107 (N_11107,N_10488,N_10325);
nor U11108 (N_11108,N_10899,N_10397);
xor U11109 (N_11109,N_10921,N_10269);
nor U11110 (N_11110,N_10984,N_10457);
nor U11111 (N_11111,N_10041,N_10906);
or U11112 (N_11112,N_10762,N_10844);
xnor U11113 (N_11113,N_10773,N_10590);
nor U11114 (N_11114,N_10824,N_10545);
xnor U11115 (N_11115,N_10926,N_10101);
or U11116 (N_11116,N_10404,N_10684);
nor U11117 (N_11117,N_10856,N_10986);
nor U11118 (N_11118,N_10484,N_10115);
or U11119 (N_11119,N_10317,N_10486);
nand U11120 (N_11120,N_10503,N_10539);
xor U11121 (N_11121,N_10910,N_10995);
nand U11122 (N_11122,N_10697,N_10247);
nor U11123 (N_11123,N_10092,N_10159);
and U11124 (N_11124,N_10354,N_10729);
xnor U11125 (N_11125,N_10434,N_10993);
xnor U11126 (N_11126,N_10128,N_10625);
or U11127 (N_11127,N_10522,N_10954);
nand U11128 (N_11128,N_10853,N_10116);
or U11129 (N_11129,N_10157,N_10277);
nand U11130 (N_11130,N_10538,N_10492);
nor U11131 (N_11131,N_10962,N_10598);
nor U11132 (N_11132,N_10246,N_10907);
or U11133 (N_11133,N_10432,N_10838);
and U11134 (N_11134,N_10802,N_10614);
xnor U11135 (N_11135,N_10742,N_10396);
nand U11136 (N_11136,N_10854,N_10111);
or U11137 (N_11137,N_10810,N_10994);
and U11138 (N_11138,N_10965,N_10395);
xnor U11139 (N_11139,N_10055,N_10973);
nand U11140 (N_11140,N_10612,N_10977);
xnor U11141 (N_11141,N_10459,N_10710);
or U11142 (N_11142,N_10309,N_10220);
xor U11143 (N_11143,N_10067,N_10677);
or U11144 (N_11144,N_10873,N_10901);
or U11145 (N_11145,N_10972,N_10706);
or U11146 (N_11146,N_10536,N_10693);
xnor U11147 (N_11147,N_10123,N_10604);
nor U11148 (N_11148,N_10547,N_10912);
and U11149 (N_11149,N_10874,N_10190);
nor U11150 (N_11150,N_10920,N_10238);
nand U11151 (N_11151,N_10126,N_10332);
or U11152 (N_11152,N_10913,N_10661);
or U11153 (N_11153,N_10348,N_10044);
and U11154 (N_11154,N_10734,N_10259);
nand U11155 (N_11155,N_10662,N_10624);
nand U11156 (N_11156,N_10370,N_10205);
nor U11157 (N_11157,N_10782,N_10433);
and U11158 (N_11158,N_10681,N_10483);
or U11159 (N_11159,N_10368,N_10437);
and U11160 (N_11160,N_10781,N_10943);
nand U11161 (N_11161,N_10064,N_10659);
and U11162 (N_11162,N_10998,N_10026);
xor U11163 (N_11163,N_10699,N_10713);
nor U11164 (N_11164,N_10618,N_10825);
xnor U11165 (N_11165,N_10981,N_10655);
nor U11166 (N_11166,N_10391,N_10209);
nor U11167 (N_11167,N_10225,N_10020);
nand U11168 (N_11168,N_10704,N_10631);
nand U11169 (N_11169,N_10414,N_10745);
or U11170 (N_11170,N_10172,N_10846);
nand U11171 (N_11171,N_10712,N_10449);
and U11172 (N_11172,N_10600,N_10435);
nor U11173 (N_11173,N_10540,N_10963);
xor U11174 (N_11174,N_10860,N_10170);
nand U11175 (N_11175,N_10867,N_10307);
nand U11176 (N_11176,N_10632,N_10224);
nand U11177 (N_11177,N_10076,N_10250);
nor U11178 (N_11178,N_10273,N_10525);
or U11179 (N_11179,N_10180,N_10398);
nor U11180 (N_11180,N_10940,N_10194);
nand U11181 (N_11181,N_10378,N_10286);
xnor U11182 (N_11182,N_10242,N_10310);
and U11183 (N_11183,N_10747,N_10937);
or U11184 (N_11184,N_10454,N_10208);
nand U11185 (N_11185,N_10330,N_10189);
and U11186 (N_11186,N_10650,N_10230);
nand U11187 (N_11187,N_10543,N_10423);
and U11188 (N_11188,N_10424,N_10583);
or U11189 (N_11189,N_10025,N_10384);
or U11190 (N_11190,N_10237,N_10908);
nor U11191 (N_11191,N_10460,N_10319);
nor U11192 (N_11192,N_10466,N_10649);
or U11193 (N_11193,N_10129,N_10426);
or U11194 (N_11194,N_10616,N_10755);
and U11195 (N_11195,N_10200,N_10610);
and U11196 (N_11196,N_10174,N_10144);
nor U11197 (N_11197,N_10411,N_10770);
and U11198 (N_11198,N_10563,N_10283);
nand U11199 (N_11199,N_10793,N_10887);
and U11200 (N_11200,N_10548,N_10744);
and U11201 (N_11201,N_10685,N_10508);
nor U11202 (N_11202,N_10280,N_10045);
xor U11203 (N_11203,N_10139,N_10670);
and U11204 (N_11204,N_10367,N_10580);
xnor U11205 (N_11205,N_10087,N_10287);
xor U11206 (N_11206,N_10477,N_10211);
nor U11207 (N_11207,N_10575,N_10176);
and U11208 (N_11208,N_10410,N_10674);
nand U11209 (N_11209,N_10613,N_10534);
nand U11210 (N_11210,N_10930,N_10979);
xor U11211 (N_11211,N_10043,N_10617);
and U11212 (N_11212,N_10009,N_10869);
xor U11213 (N_11213,N_10152,N_10791);
and U11214 (N_11214,N_10982,N_10008);
xor U11215 (N_11215,N_10915,N_10427);
and U11216 (N_11216,N_10728,N_10584);
and U11217 (N_11217,N_10643,N_10002);
nand U11218 (N_11218,N_10905,N_10669);
nand U11219 (N_11219,N_10383,N_10808);
nand U11220 (N_11220,N_10108,N_10469);
xnor U11221 (N_11221,N_10007,N_10961);
or U11222 (N_11222,N_10254,N_10133);
nand U11223 (N_11223,N_10487,N_10335);
nor U11224 (N_11224,N_10720,N_10717);
or U11225 (N_11225,N_10066,N_10216);
xnor U11226 (N_11226,N_10421,N_10997);
nand U11227 (N_11227,N_10974,N_10953);
nand U11228 (N_11228,N_10154,N_10933);
or U11229 (N_11229,N_10620,N_10533);
nand U11230 (N_11230,N_10761,N_10160);
and U11231 (N_11231,N_10499,N_10516);
nand U11232 (N_11232,N_10805,N_10837);
or U11233 (N_11233,N_10806,N_10722);
nor U11234 (N_11234,N_10608,N_10183);
nand U11235 (N_11235,N_10351,N_10258);
or U11236 (N_11236,N_10463,N_10357);
nand U11237 (N_11237,N_10316,N_10479);
nor U11238 (N_11238,N_10592,N_10771);
nor U11239 (N_11239,N_10857,N_10757);
nand U11240 (N_11240,N_10490,N_10000);
and U11241 (N_11241,N_10001,N_10731);
and U11242 (N_11242,N_10850,N_10726);
nand U11243 (N_11243,N_10698,N_10402);
or U11244 (N_11244,N_10835,N_10885);
nor U11245 (N_11245,N_10102,N_10602);
or U11246 (N_11246,N_10554,N_10507);
or U11247 (N_11247,N_10970,N_10918);
xor U11248 (N_11248,N_10891,N_10958);
nor U11249 (N_11249,N_10082,N_10339);
nand U11250 (N_11250,N_10514,N_10541);
nor U11251 (N_11251,N_10267,N_10692);
nand U11252 (N_11252,N_10222,N_10050);
xnor U11253 (N_11253,N_10217,N_10502);
and U11254 (N_11254,N_10888,N_10117);
and U11255 (N_11255,N_10171,N_10585);
xor U11256 (N_11256,N_10778,N_10428);
or U11257 (N_11257,N_10515,N_10125);
or U11258 (N_11258,N_10168,N_10196);
nor U11259 (N_11259,N_10892,N_10003);
nor U11260 (N_11260,N_10828,N_10084);
and U11261 (N_11261,N_10809,N_10830);
nor U11262 (N_11262,N_10240,N_10047);
or U11263 (N_11263,N_10493,N_10881);
nor U11264 (N_11264,N_10826,N_10517);
xnor U11265 (N_11265,N_10058,N_10149);
and U11266 (N_11266,N_10817,N_10178);
nand U11267 (N_11267,N_10415,N_10333);
or U11268 (N_11268,N_10739,N_10193);
nand U11269 (N_11269,N_10218,N_10166);
or U11270 (N_11270,N_10736,N_10377);
nand U11271 (N_11271,N_10298,N_10566);
or U11272 (N_11272,N_10132,N_10297);
xnor U11273 (N_11273,N_10071,N_10253);
nand U11274 (N_11274,N_10936,N_10852);
xnor U11275 (N_11275,N_10676,N_10911);
nand U11276 (N_11276,N_10155,N_10296);
nand U11277 (N_11277,N_10870,N_10637);
xor U11278 (N_11278,N_10161,N_10407);
and U11279 (N_11279,N_10416,N_10299);
or U11280 (N_11280,N_10754,N_10195);
nor U11281 (N_11281,N_10197,N_10879);
nor U11282 (N_11282,N_10644,N_10480);
or U11283 (N_11283,N_10199,N_10346);
or U11284 (N_11284,N_10667,N_10855);
and U11285 (N_11285,N_10264,N_10495);
or U11286 (N_11286,N_10562,N_10763);
nand U11287 (N_11287,N_10672,N_10831);
xnor U11288 (N_11288,N_10500,N_10701);
xor U11289 (N_11289,N_10135,N_10345);
and U11290 (N_11290,N_10599,N_10094);
and U11291 (N_11291,N_10039,N_10145);
or U11292 (N_11292,N_10959,N_10430);
or U11293 (N_11293,N_10683,N_10680);
and U11294 (N_11294,N_10796,N_10311);
and U11295 (N_11295,N_10284,N_10233);
or U11296 (N_11296,N_10924,N_10923);
and U11297 (N_11297,N_10549,N_10591);
nor U11298 (N_11298,N_10895,N_10093);
and U11299 (N_11299,N_10336,N_10389);
and U11300 (N_11300,N_10948,N_10052);
nand U11301 (N_11301,N_10202,N_10767);
nor U11302 (N_11302,N_10086,N_10095);
xnor U11303 (N_11303,N_10313,N_10561);
nor U11304 (N_11304,N_10675,N_10227);
or U11305 (N_11305,N_10439,N_10967);
or U11306 (N_11306,N_10090,N_10709);
nor U11307 (N_11307,N_10651,N_10653);
xor U11308 (N_11308,N_10441,N_10509);
xnor U11309 (N_11309,N_10950,N_10866);
or U11310 (N_11310,N_10898,N_10327);
nand U11311 (N_11311,N_10350,N_10567);
xnor U11312 (N_11312,N_10110,N_10274);
or U11313 (N_11313,N_10361,N_10691);
or U11314 (N_11314,N_10184,N_10839);
or U11315 (N_11315,N_10903,N_10576);
xor U11316 (N_11316,N_10446,N_10978);
and U11317 (N_11317,N_10293,N_10932);
xor U11318 (N_11318,N_10475,N_10942);
or U11319 (N_11319,N_10051,N_10902);
or U11320 (N_11320,N_10647,N_10759);
xor U11321 (N_11321,N_10011,N_10657);
or U11322 (N_11322,N_10785,N_10738);
nor U11323 (N_11323,N_10577,N_10360);
nand U11324 (N_11324,N_10344,N_10894);
nor U11325 (N_11325,N_10890,N_10615);
nand U11326 (N_11326,N_10422,N_10380);
and U11327 (N_11327,N_10927,N_10630);
nor U11328 (N_11328,N_10639,N_10581);
xnor U11329 (N_11329,N_10871,N_10136);
or U11330 (N_11330,N_10214,N_10158);
xnor U11331 (N_11331,N_10290,N_10255);
nor U11332 (N_11332,N_10060,N_10506);
and U11333 (N_11333,N_10418,N_10028);
and U11334 (N_11334,N_10818,N_10303);
nand U11335 (N_11335,N_10363,N_10570);
or U11336 (N_11336,N_10840,N_10727);
or U11337 (N_11337,N_10098,N_10289);
nand U11338 (N_11338,N_10443,N_10491);
nor U11339 (N_11339,N_10552,N_10551);
xnor U11340 (N_11340,N_10379,N_10884);
or U11341 (N_11341,N_10279,N_10510);
and U11342 (N_11342,N_10369,N_10938);
or U11343 (N_11343,N_10696,N_10100);
nor U11344 (N_11344,N_10029,N_10597);
xor U11345 (N_11345,N_10470,N_10990);
and U11346 (N_11346,N_10324,N_10851);
nor U11347 (N_11347,N_10364,N_10783);
nor U11348 (N_11348,N_10027,N_10231);
or U11349 (N_11349,N_10334,N_10504);
nand U11350 (N_11350,N_10249,N_10177);
nand U11351 (N_11351,N_10315,N_10595);
and U11352 (N_11352,N_10956,N_10530);
nand U11353 (N_11353,N_10381,N_10665);
or U11354 (N_11354,N_10935,N_10594);
and U11355 (N_11355,N_10472,N_10724);
nor U11356 (N_11356,N_10109,N_10646);
and U11357 (N_11357,N_10167,N_10138);
nand U11358 (N_11358,N_10593,N_10281);
nor U11359 (N_11359,N_10308,N_10529);
and U11360 (N_11360,N_10634,N_10292);
nand U11361 (N_11361,N_10679,N_10103);
and U11362 (N_11362,N_10099,N_10455);
or U11363 (N_11363,N_10987,N_10012);
xnor U11364 (N_11364,N_10251,N_10572);
or U11365 (N_11365,N_10023,N_10314);
nor U11366 (N_11366,N_10711,N_10641);
nor U11367 (N_11367,N_10776,N_10587);
and U11368 (N_11368,N_10966,N_10694);
xnor U11369 (N_11369,N_10412,N_10931);
xnor U11370 (N_11370,N_10758,N_10083);
or U11371 (N_11371,N_10886,N_10341);
and U11372 (N_11372,N_10393,N_10445);
nor U11373 (N_11373,N_10405,N_10521);
nand U11374 (N_11374,N_10772,N_10312);
nand U11375 (N_11375,N_10257,N_10417);
nor U11376 (N_11376,N_10121,N_10880);
nor U11377 (N_11377,N_10976,N_10682);
or U11378 (N_11378,N_10358,N_10842);
nor U11379 (N_11379,N_10429,N_10800);
xor U11380 (N_11380,N_10553,N_10733);
and U11381 (N_11381,N_10568,N_10373);
xnor U11382 (N_11382,N_10816,N_10941);
xor U11383 (N_11383,N_10465,N_10175);
or U11384 (N_11384,N_10832,N_10034);
xor U11385 (N_11385,N_10980,N_10498);
nand U11386 (N_11386,N_10431,N_10519);
and U11387 (N_11387,N_10863,N_10347);
nor U11388 (N_11388,N_10239,N_10142);
xnor U11389 (N_11389,N_10323,N_10542);
or U11390 (N_11390,N_10219,N_10010);
nor U11391 (N_11391,N_10163,N_10137);
or U11392 (N_11392,N_10512,N_10118);
nor U11393 (N_11393,N_10564,N_10686);
nor U11394 (N_11394,N_10065,N_10127);
and U11395 (N_11395,N_10300,N_10947);
nor U11396 (N_11396,N_10636,N_10069);
xnor U11397 (N_11397,N_10983,N_10147);
nor U11398 (N_11398,N_10114,N_10928);
and U11399 (N_11399,N_10819,N_10374);
and U11400 (N_11400,N_10688,N_10814);
xnor U11401 (N_11401,N_10946,N_10037);
nand U11402 (N_11402,N_10425,N_10708);
or U11403 (N_11403,N_10215,N_10558);
and U11404 (N_11404,N_10485,N_10294);
xnor U11405 (N_11405,N_10033,N_10841);
and U11406 (N_11406,N_10061,N_10603);
nor U11407 (N_11407,N_10022,N_10703);
nand U11408 (N_11408,N_10546,N_10245);
or U11409 (N_11409,N_10187,N_10005);
and U11410 (N_11410,N_10969,N_10444);
nand U11411 (N_11411,N_10596,N_10666);
nor U11412 (N_11412,N_10801,N_10400);
nand U11413 (N_11413,N_10606,N_10574);
or U11414 (N_11414,N_10756,N_10964);
and U11415 (N_11415,N_10971,N_10847);
and U11416 (N_11416,N_10531,N_10795);
and U11417 (N_11417,N_10059,N_10829);
nor U11418 (N_11418,N_10248,N_10226);
nand U11419 (N_11419,N_10482,N_10556);
nor U11420 (N_11420,N_10544,N_10904);
xnor U11421 (N_11421,N_10735,N_10223);
xor U11422 (N_11422,N_10232,N_10165);
xnor U11423 (N_11423,N_10153,N_10376);
or U11424 (N_11424,N_10342,N_10392);
and U11425 (N_11425,N_10601,N_10929);
nand U11426 (N_11426,N_10815,N_10764);
nor U11427 (N_11427,N_10419,N_10276);
nand U11428 (N_11428,N_10053,N_10718);
nor U11429 (N_11429,N_10843,N_10845);
nand U11430 (N_11430,N_10301,N_10622);
nor U11431 (N_11431,N_10440,N_10812);
nand U11432 (N_11432,N_10451,N_10075);
nor U11433 (N_11433,N_10288,N_10952);
or U11434 (N_11434,N_10550,N_10766);
xor U11435 (N_11435,N_10261,N_10270);
or U11436 (N_11436,N_10046,N_10513);
or U11437 (N_11437,N_10385,N_10447);
and U11438 (N_11438,N_10528,N_10985);
nand U11439 (N_11439,N_10408,N_10648);
nor U11440 (N_11440,N_10120,N_10150);
and U11441 (N_11441,N_10573,N_10951);
or U11442 (N_11442,N_10131,N_10382);
or U11443 (N_11443,N_10031,N_10304);
xnor U11444 (N_11444,N_10740,N_10306);
or U11445 (N_11445,N_10173,N_10268);
nand U11446 (N_11446,N_10678,N_10586);
and U11447 (N_11447,N_10714,N_10900);
nand U11448 (N_11448,N_10456,N_10353);
nor U11449 (N_11449,N_10122,N_10868);
or U11450 (N_11450,N_10352,N_10203);
nor U11451 (N_11451,N_10925,N_10991);
nand U11452 (N_11452,N_10934,N_10221);
nor U11453 (N_11453,N_10737,N_10077);
or U11454 (N_11454,N_10537,N_10073);
xor U11455 (N_11455,N_10996,N_10468);
or U11456 (N_11456,N_10511,N_10640);
or U11457 (N_11457,N_10467,N_10387);
or U11458 (N_11458,N_10228,N_10464);
nand U11459 (N_11459,N_10645,N_10164);
xor U11460 (N_11460,N_10788,N_10018);
or U11461 (N_11461,N_10406,N_10062);
and U11462 (N_11462,N_10386,N_10579);
xnor U11463 (N_11463,N_10004,N_10295);
nor U11464 (N_11464,N_10442,N_10119);
xor U11465 (N_11465,N_10769,N_10191);
nor U11466 (N_11466,N_10760,N_10182);
and U11467 (N_11467,N_10571,N_10786);
xor U11468 (N_11468,N_10949,N_10049);
xor U11469 (N_11469,N_10085,N_10721);
nand U11470 (N_11470,N_10213,N_10858);
and U11471 (N_11471,N_10343,N_10780);
or U11472 (N_11472,N_10212,N_10017);
nor U11473 (N_11473,N_10748,N_10605);
or U11474 (N_11474,N_10876,N_10804);
and U11475 (N_11475,N_10006,N_10497);
or U11476 (N_11476,N_10048,N_10291);
and U11477 (N_11477,N_10375,N_10960);
nor U11478 (N_11478,N_10078,N_10673);
nor U11479 (N_11479,N_10532,N_10156);
nand U11480 (N_11480,N_10113,N_10882);
nand U11481 (N_11481,N_10633,N_10989);
and U11482 (N_11482,N_10790,N_10337);
and U11483 (N_11483,N_10179,N_10883);
xor U11484 (N_11484,N_10652,N_10204);
or U11485 (N_11485,N_10148,N_10365);
nor U11486 (N_11486,N_10169,N_10206);
xnor U11487 (N_11487,N_10792,N_10768);
nor U11488 (N_11488,N_10753,N_10054);
nor U11489 (N_11489,N_10151,N_10765);
or U11490 (N_11490,N_10244,N_10527);
and U11491 (N_11491,N_10557,N_10074);
nand U11492 (N_11492,N_10072,N_10505);
nand U11493 (N_11493,N_10420,N_10359);
and U11494 (N_11494,N_10014,N_10654);
and U11495 (N_11495,N_10474,N_10494);
xor U11496 (N_11496,N_10331,N_10909);
or U11497 (N_11497,N_10524,N_10741);
xor U11498 (N_11498,N_10609,N_10134);
or U11499 (N_11499,N_10235,N_10436);
nand U11500 (N_11500,N_10092,N_10973);
nand U11501 (N_11501,N_10546,N_10769);
xnor U11502 (N_11502,N_10928,N_10397);
nor U11503 (N_11503,N_10817,N_10233);
and U11504 (N_11504,N_10498,N_10792);
nor U11505 (N_11505,N_10700,N_10758);
and U11506 (N_11506,N_10735,N_10229);
and U11507 (N_11507,N_10595,N_10090);
and U11508 (N_11508,N_10099,N_10412);
or U11509 (N_11509,N_10037,N_10249);
nor U11510 (N_11510,N_10926,N_10777);
nand U11511 (N_11511,N_10769,N_10754);
nand U11512 (N_11512,N_10009,N_10787);
xor U11513 (N_11513,N_10439,N_10685);
or U11514 (N_11514,N_10005,N_10599);
and U11515 (N_11515,N_10189,N_10651);
xnor U11516 (N_11516,N_10954,N_10923);
and U11517 (N_11517,N_10201,N_10406);
xor U11518 (N_11518,N_10554,N_10637);
and U11519 (N_11519,N_10588,N_10199);
or U11520 (N_11520,N_10804,N_10847);
and U11521 (N_11521,N_10892,N_10384);
nand U11522 (N_11522,N_10340,N_10680);
nand U11523 (N_11523,N_10980,N_10110);
or U11524 (N_11524,N_10377,N_10435);
nor U11525 (N_11525,N_10470,N_10638);
or U11526 (N_11526,N_10187,N_10354);
xnor U11527 (N_11527,N_10430,N_10541);
nor U11528 (N_11528,N_10632,N_10496);
and U11529 (N_11529,N_10502,N_10591);
nor U11530 (N_11530,N_10972,N_10795);
nand U11531 (N_11531,N_10206,N_10476);
or U11532 (N_11532,N_10248,N_10704);
or U11533 (N_11533,N_10995,N_10665);
xor U11534 (N_11534,N_10837,N_10146);
xor U11535 (N_11535,N_10276,N_10689);
nand U11536 (N_11536,N_10443,N_10196);
or U11537 (N_11537,N_10092,N_10183);
and U11538 (N_11538,N_10101,N_10275);
nor U11539 (N_11539,N_10780,N_10254);
and U11540 (N_11540,N_10129,N_10582);
nor U11541 (N_11541,N_10780,N_10441);
and U11542 (N_11542,N_10136,N_10383);
xor U11543 (N_11543,N_10121,N_10595);
nor U11544 (N_11544,N_10101,N_10244);
and U11545 (N_11545,N_10557,N_10129);
and U11546 (N_11546,N_10625,N_10528);
nand U11547 (N_11547,N_10473,N_10179);
nand U11548 (N_11548,N_10659,N_10214);
and U11549 (N_11549,N_10939,N_10863);
nand U11550 (N_11550,N_10523,N_10241);
nor U11551 (N_11551,N_10049,N_10522);
xor U11552 (N_11552,N_10861,N_10027);
and U11553 (N_11553,N_10114,N_10984);
xnor U11554 (N_11554,N_10930,N_10942);
xnor U11555 (N_11555,N_10777,N_10981);
or U11556 (N_11556,N_10003,N_10896);
nor U11557 (N_11557,N_10411,N_10142);
and U11558 (N_11558,N_10282,N_10079);
nand U11559 (N_11559,N_10891,N_10080);
or U11560 (N_11560,N_10448,N_10872);
xor U11561 (N_11561,N_10373,N_10554);
xor U11562 (N_11562,N_10405,N_10602);
and U11563 (N_11563,N_10663,N_10614);
or U11564 (N_11564,N_10475,N_10996);
xor U11565 (N_11565,N_10730,N_10827);
xnor U11566 (N_11566,N_10359,N_10865);
or U11567 (N_11567,N_10794,N_10774);
xor U11568 (N_11568,N_10565,N_10738);
and U11569 (N_11569,N_10232,N_10512);
xor U11570 (N_11570,N_10623,N_10223);
and U11571 (N_11571,N_10820,N_10866);
nor U11572 (N_11572,N_10015,N_10181);
nor U11573 (N_11573,N_10066,N_10137);
and U11574 (N_11574,N_10981,N_10710);
xnor U11575 (N_11575,N_10602,N_10814);
and U11576 (N_11576,N_10968,N_10951);
nand U11577 (N_11577,N_10659,N_10570);
nor U11578 (N_11578,N_10971,N_10445);
nor U11579 (N_11579,N_10852,N_10401);
or U11580 (N_11580,N_10020,N_10995);
and U11581 (N_11581,N_10381,N_10220);
nor U11582 (N_11582,N_10395,N_10206);
or U11583 (N_11583,N_10484,N_10827);
and U11584 (N_11584,N_10015,N_10037);
xnor U11585 (N_11585,N_10268,N_10562);
and U11586 (N_11586,N_10666,N_10152);
or U11587 (N_11587,N_10578,N_10080);
nor U11588 (N_11588,N_10007,N_10166);
and U11589 (N_11589,N_10366,N_10494);
and U11590 (N_11590,N_10254,N_10320);
nor U11591 (N_11591,N_10838,N_10968);
nor U11592 (N_11592,N_10831,N_10095);
xnor U11593 (N_11593,N_10438,N_10166);
and U11594 (N_11594,N_10806,N_10326);
and U11595 (N_11595,N_10252,N_10230);
nor U11596 (N_11596,N_10712,N_10620);
or U11597 (N_11597,N_10550,N_10194);
or U11598 (N_11598,N_10060,N_10129);
xnor U11599 (N_11599,N_10064,N_10030);
nand U11600 (N_11600,N_10830,N_10802);
nor U11601 (N_11601,N_10768,N_10685);
xor U11602 (N_11602,N_10141,N_10708);
and U11603 (N_11603,N_10644,N_10157);
xnor U11604 (N_11604,N_10761,N_10746);
xor U11605 (N_11605,N_10376,N_10089);
nand U11606 (N_11606,N_10564,N_10814);
nand U11607 (N_11607,N_10566,N_10485);
xor U11608 (N_11608,N_10698,N_10984);
xnor U11609 (N_11609,N_10608,N_10207);
and U11610 (N_11610,N_10490,N_10854);
nor U11611 (N_11611,N_10258,N_10921);
nand U11612 (N_11612,N_10119,N_10703);
nand U11613 (N_11613,N_10174,N_10853);
nor U11614 (N_11614,N_10683,N_10315);
xnor U11615 (N_11615,N_10747,N_10745);
xnor U11616 (N_11616,N_10835,N_10785);
xnor U11617 (N_11617,N_10616,N_10585);
xnor U11618 (N_11618,N_10785,N_10479);
xnor U11619 (N_11619,N_10579,N_10133);
nand U11620 (N_11620,N_10559,N_10755);
nand U11621 (N_11621,N_10301,N_10499);
nand U11622 (N_11622,N_10701,N_10142);
or U11623 (N_11623,N_10173,N_10634);
nor U11624 (N_11624,N_10222,N_10472);
and U11625 (N_11625,N_10774,N_10795);
xnor U11626 (N_11626,N_10403,N_10312);
nand U11627 (N_11627,N_10729,N_10511);
and U11628 (N_11628,N_10460,N_10409);
or U11629 (N_11629,N_10372,N_10489);
nor U11630 (N_11630,N_10654,N_10821);
xnor U11631 (N_11631,N_10852,N_10515);
nand U11632 (N_11632,N_10340,N_10947);
xnor U11633 (N_11633,N_10706,N_10328);
nor U11634 (N_11634,N_10615,N_10196);
or U11635 (N_11635,N_10786,N_10735);
xor U11636 (N_11636,N_10308,N_10757);
xnor U11637 (N_11637,N_10559,N_10162);
nor U11638 (N_11638,N_10514,N_10232);
or U11639 (N_11639,N_10270,N_10373);
and U11640 (N_11640,N_10668,N_10429);
xor U11641 (N_11641,N_10906,N_10152);
or U11642 (N_11642,N_10036,N_10705);
xnor U11643 (N_11643,N_10762,N_10485);
and U11644 (N_11644,N_10090,N_10914);
xor U11645 (N_11645,N_10167,N_10627);
nor U11646 (N_11646,N_10720,N_10446);
and U11647 (N_11647,N_10211,N_10676);
xnor U11648 (N_11648,N_10206,N_10543);
nand U11649 (N_11649,N_10461,N_10410);
and U11650 (N_11650,N_10314,N_10455);
nor U11651 (N_11651,N_10956,N_10637);
and U11652 (N_11652,N_10381,N_10732);
xnor U11653 (N_11653,N_10747,N_10465);
nand U11654 (N_11654,N_10208,N_10301);
and U11655 (N_11655,N_10385,N_10128);
nand U11656 (N_11656,N_10504,N_10984);
nand U11657 (N_11657,N_10896,N_10525);
nor U11658 (N_11658,N_10795,N_10763);
and U11659 (N_11659,N_10061,N_10030);
or U11660 (N_11660,N_10023,N_10390);
or U11661 (N_11661,N_10017,N_10513);
and U11662 (N_11662,N_10238,N_10688);
and U11663 (N_11663,N_10641,N_10991);
and U11664 (N_11664,N_10981,N_10407);
or U11665 (N_11665,N_10042,N_10399);
nand U11666 (N_11666,N_10472,N_10304);
and U11667 (N_11667,N_10320,N_10323);
nor U11668 (N_11668,N_10502,N_10704);
and U11669 (N_11669,N_10301,N_10325);
nand U11670 (N_11670,N_10374,N_10762);
and U11671 (N_11671,N_10048,N_10830);
nor U11672 (N_11672,N_10071,N_10320);
nor U11673 (N_11673,N_10537,N_10072);
nor U11674 (N_11674,N_10699,N_10880);
and U11675 (N_11675,N_10910,N_10833);
xnor U11676 (N_11676,N_10788,N_10320);
and U11677 (N_11677,N_10711,N_10922);
or U11678 (N_11678,N_10213,N_10149);
xnor U11679 (N_11679,N_10875,N_10957);
and U11680 (N_11680,N_10604,N_10536);
or U11681 (N_11681,N_10446,N_10279);
xor U11682 (N_11682,N_10115,N_10045);
xor U11683 (N_11683,N_10483,N_10437);
or U11684 (N_11684,N_10407,N_10314);
nor U11685 (N_11685,N_10601,N_10041);
nand U11686 (N_11686,N_10452,N_10016);
nor U11687 (N_11687,N_10116,N_10158);
nand U11688 (N_11688,N_10698,N_10863);
xnor U11689 (N_11689,N_10455,N_10022);
and U11690 (N_11690,N_10563,N_10191);
and U11691 (N_11691,N_10313,N_10655);
xnor U11692 (N_11692,N_10029,N_10333);
and U11693 (N_11693,N_10143,N_10327);
or U11694 (N_11694,N_10658,N_10195);
or U11695 (N_11695,N_10977,N_10314);
and U11696 (N_11696,N_10521,N_10056);
xnor U11697 (N_11697,N_10726,N_10403);
and U11698 (N_11698,N_10848,N_10928);
nand U11699 (N_11699,N_10959,N_10561);
nor U11700 (N_11700,N_10146,N_10326);
xnor U11701 (N_11701,N_10114,N_10383);
xnor U11702 (N_11702,N_10416,N_10091);
xnor U11703 (N_11703,N_10681,N_10697);
and U11704 (N_11704,N_10367,N_10690);
nor U11705 (N_11705,N_10433,N_10199);
nor U11706 (N_11706,N_10285,N_10315);
and U11707 (N_11707,N_10405,N_10304);
and U11708 (N_11708,N_10349,N_10580);
nand U11709 (N_11709,N_10812,N_10543);
or U11710 (N_11710,N_10644,N_10230);
or U11711 (N_11711,N_10629,N_10166);
nor U11712 (N_11712,N_10507,N_10439);
nand U11713 (N_11713,N_10200,N_10591);
nand U11714 (N_11714,N_10217,N_10163);
and U11715 (N_11715,N_10196,N_10864);
or U11716 (N_11716,N_10192,N_10771);
nor U11717 (N_11717,N_10747,N_10176);
and U11718 (N_11718,N_10770,N_10497);
nand U11719 (N_11719,N_10814,N_10302);
or U11720 (N_11720,N_10632,N_10378);
xnor U11721 (N_11721,N_10696,N_10361);
nand U11722 (N_11722,N_10538,N_10993);
nand U11723 (N_11723,N_10102,N_10317);
nand U11724 (N_11724,N_10358,N_10438);
or U11725 (N_11725,N_10231,N_10576);
xor U11726 (N_11726,N_10469,N_10104);
nor U11727 (N_11727,N_10603,N_10545);
and U11728 (N_11728,N_10990,N_10271);
nand U11729 (N_11729,N_10766,N_10159);
or U11730 (N_11730,N_10697,N_10051);
xor U11731 (N_11731,N_10304,N_10906);
xor U11732 (N_11732,N_10597,N_10799);
xnor U11733 (N_11733,N_10978,N_10036);
and U11734 (N_11734,N_10681,N_10657);
xor U11735 (N_11735,N_10821,N_10989);
nand U11736 (N_11736,N_10347,N_10500);
or U11737 (N_11737,N_10299,N_10241);
and U11738 (N_11738,N_10961,N_10086);
nor U11739 (N_11739,N_10405,N_10616);
nor U11740 (N_11740,N_10637,N_10893);
nand U11741 (N_11741,N_10055,N_10214);
and U11742 (N_11742,N_10210,N_10966);
nor U11743 (N_11743,N_10149,N_10124);
nor U11744 (N_11744,N_10818,N_10429);
xor U11745 (N_11745,N_10758,N_10869);
and U11746 (N_11746,N_10020,N_10545);
and U11747 (N_11747,N_10267,N_10491);
or U11748 (N_11748,N_10537,N_10237);
nor U11749 (N_11749,N_10699,N_10689);
nand U11750 (N_11750,N_10364,N_10431);
or U11751 (N_11751,N_10405,N_10436);
nor U11752 (N_11752,N_10502,N_10995);
nor U11753 (N_11753,N_10042,N_10305);
xor U11754 (N_11754,N_10082,N_10085);
xnor U11755 (N_11755,N_10325,N_10065);
or U11756 (N_11756,N_10375,N_10142);
nor U11757 (N_11757,N_10383,N_10347);
and U11758 (N_11758,N_10057,N_10592);
xor U11759 (N_11759,N_10644,N_10571);
nor U11760 (N_11760,N_10493,N_10955);
or U11761 (N_11761,N_10898,N_10661);
xor U11762 (N_11762,N_10327,N_10330);
nand U11763 (N_11763,N_10759,N_10643);
nand U11764 (N_11764,N_10954,N_10991);
nor U11765 (N_11765,N_10096,N_10254);
or U11766 (N_11766,N_10129,N_10451);
nand U11767 (N_11767,N_10264,N_10560);
nor U11768 (N_11768,N_10566,N_10986);
nor U11769 (N_11769,N_10292,N_10811);
nand U11770 (N_11770,N_10950,N_10446);
nand U11771 (N_11771,N_10347,N_10322);
nor U11772 (N_11772,N_10671,N_10391);
and U11773 (N_11773,N_10757,N_10558);
nor U11774 (N_11774,N_10537,N_10382);
nand U11775 (N_11775,N_10188,N_10781);
nor U11776 (N_11776,N_10765,N_10600);
nor U11777 (N_11777,N_10492,N_10074);
and U11778 (N_11778,N_10337,N_10238);
or U11779 (N_11779,N_10053,N_10188);
nand U11780 (N_11780,N_10514,N_10210);
or U11781 (N_11781,N_10413,N_10509);
nand U11782 (N_11782,N_10360,N_10700);
xor U11783 (N_11783,N_10139,N_10880);
and U11784 (N_11784,N_10208,N_10750);
or U11785 (N_11785,N_10811,N_10920);
nor U11786 (N_11786,N_10317,N_10320);
xor U11787 (N_11787,N_10527,N_10826);
and U11788 (N_11788,N_10921,N_10711);
nor U11789 (N_11789,N_10514,N_10215);
and U11790 (N_11790,N_10847,N_10919);
or U11791 (N_11791,N_10902,N_10146);
and U11792 (N_11792,N_10534,N_10635);
nand U11793 (N_11793,N_10649,N_10562);
nand U11794 (N_11794,N_10333,N_10091);
xnor U11795 (N_11795,N_10442,N_10957);
nand U11796 (N_11796,N_10886,N_10480);
or U11797 (N_11797,N_10944,N_10947);
or U11798 (N_11798,N_10902,N_10791);
and U11799 (N_11799,N_10383,N_10147);
nor U11800 (N_11800,N_10824,N_10479);
and U11801 (N_11801,N_10574,N_10732);
nand U11802 (N_11802,N_10474,N_10287);
nor U11803 (N_11803,N_10686,N_10535);
nand U11804 (N_11804,N_10889,N_10935);
or U11805 (N_11805,N_10394,N_10176);
nor U11806 (N_11806,N_10074,N_10623);
nand U11807 (N_11807,N_10395,N_10476);
nand U11808 (N_11808,N_10590,N_10424);
or U11809 (N_11809,N_10119,N_10488);
xnor U11810 (N_11810,N_10035,N_10678);
nand U11811 (N_11811,N_10639,N_10274);
and U11812 (N_11812,N_10794,N_10840);
or U11813 (N_11813,N_10455,N_10698);
xnor U11814 (N_11814,N_10019,N_10120);
nand U11815 (N_11815,N_10767,N_10259);
nor U11816 (N_11816,N_10647,N_10163);
xnor U11817 (N_11817,N_10256,N_10066);
and U11818 (N_11818,N_10284,N_10314);
or U11819 (N_11819,N_10030,N_10855);
nor U11820 (N_11820,N_10841,N_10849);
xor U11821 (N_11821,N_10393,N_10645);
or U11822 (N_11822,N_10842,N_10258);
nand U11823 (N_11823,N_10944,N_10746);
xnor U11824 (N_11824,N_10456,N_10227);
nand U11825 (N_11825,N_10711,N_10864);
nand U11826 (N_11826,N_10990,N_10596);
nand U11827 (N_11827,N_10257,N_10218);
nand U11828 (N_11828,N_10858,N_10689);
and U11829 (N_11829,N_10496,N_10926);
or U11830 (N_11830,N_10472,N_10691);
nor U11831 (N_11831,N_10209,N_10110);
xor U11832 (N_11832,N_10766,N_10475);
or U11833 (N_11833,N_10271,N_10095);
nand U11834 (N_11834,N_10599,N_10146);
xnor U11835 (N_11835,N_10017,N_10068);
nor U11836 (N_11836,N_10709,N_10987);
nor U11837 (N_11837,N_10877,N_10670);
xnor U11838 (N_11838,N_10857,N_10780);
and U11839 (N_11839,N_10199,N_10539);
and U11840 (N_11840,N_10952,N_10649);
xnor U11841 (N_11841,N_10665,N_10230);
xnor U11842 (N_11842,N_10065,N_10424);
xnor U11843 (N_11843,N_10977,N_10981);
xnor U11844 (N_11844,N_10564,N_10746);
nor U11845 (N_11845,N_10228,N_10788);
or U11846 (N_11846,N_10961,N_10879);
nand U11847 (N_11847,N_10811,N_10824);
or U11848 (N_11848,N_10387,N_10413);
and U11849 (N_11849,N_10449,N_10719);
or U11850 (N_11850,N_10625,N_10383);
nand U11851 (N_11851,N_10020,N_10213);
nor U11852 (N_11852,N_10895,N_10577);
xnor U11853 (N_11853,N_10201,N_10206);
nand U11854 (N_11854,N_10467,N_10276);
and U11855 (N_11855,N_10095,N_10565);
nand U11856 (N_11856,N_10579,N_10892);
nand U11857 (N_11857,N_10353,N_10211);
nor U11858 (N_11858,N_10991,N_10057);
or U11859 (N_11859,N_10539,N_10202);
nand U11860 (N_11860,N_10018,N_10482);
nor U11861 (N_11861,N_10865,N_10302);
xor U11862 (N_11862,N_10016,N_10040);
nor U11863 (N_11863,N_10027,N_10582);
xnor U11864 (N_11864,N_10365,N_10941);
nor U11865 (N_11865,N_10585,N_10539);
or U11866 (N_11866,N_10355,N_10282);
nor U11867 (N_11867,N_10977,N_10439);
and U11868 (N_11868,N_10783,N_10918);
xnor U11869 (N_11869,N_10857,N_10309);
nand U11870 (N_11870,N_10366,N_10760);
and U11871 (N_11871,N_10189,N_10993);
xnor U11872 (N_11872,N_10377,N_10437);
nor U11873 (N_11873,N_10600,N_10927);
nand U11874 (N_11874,N_10941,N_10240);
or U11875 (N_11875,N_10850,N_10718);
xnor U11876 (N_11876,N_10401,N_10975);
nor U11877 (N_11877,N_10499,N_10156);
nor U11878 (N_11878,N_10999,N_10796);
nor U11879 (N_11879,N_10839,N_10175);
and U11880 (N_11880,N_10201,N_10420);
xor U11881 (N_11881,N_10514,N_10135);
xor U11882 (N_11882,N_10915,N_10108);
and U11883 (N_11883,N_10716,N_10752);
or U11884 (N_11884,N_10789,N_10688);
and U11885 (N_11885,N_10781,N_10273);
nor U11886 (N_11886,N_10941,N_10805);
nor U11887 (N_11887,N_10013,N_10290);
and U11888 (N_11888,N_10265,N_10826);
nand U11889 (N_11889,N_10912,N_10899);
or U11890 (N_11890,N_10203,N_10897);
xnor U11891 (N_11891,N_10531,N_10551);
nand U11892 (N_11892,N_10466,N_10079);
nor U11893 (N_11893,N_10806,N_10592);
nand U11894 (N_11894,N_10093,N_10056);
xor U11895 (N_11895,N_10129,N_10323);
and U11896 (N_11896,N_10903,N_10744);
nand U11897 (N_11897,N_10546,N_10617);
or U11898 (N_11898,N_10808,N_10877);
nor U11899 (N_11899,N_10689,N_10164);
nor U11900 (N_11900,N_10935,N_10179);
xor U11901 (N_11901,N_10324,N_10368);
nand U11902 (N_11902,N_10063,N_10352);
nand U11903 (N_11903,N_10045,N_10735);
nand U11904 (N_11904,N_10721,N_10575);
and U11905 (N_11905,N_10323,N_10994);
and U11906 (N_11906,N_10476,N_10138);
or U11907 (N_11907,N_10939,N_10528);
nor U11908 (N_11908,N_10123,N_10945);
xnor U11909 (N_11909,N_10078,N_10798);
xnor U11910 (N_11910,N_10138,N_10871);
nand U11911 (N_11911,N_10095,N_10376);
or U11912 (N_11912,N_10731,N_10662);
nor U11913 (N_11913,N_10664,N_10935);
or U11914 (N_11914,N_10545,N_10731);
nor U11915 (N_11915,N_10241,N_10360);
nor U11916 (N_11916,N_10179,N_10856);
or U11917 (N_11917,N_10863,N_10365);
nand U11918 (N_11918,N_10142,N_10978);
and U11919 (N_11919,N_10944,N_10213);
and U11920 (N_11920,N_10407,N_10872);
nand U11921 (N_11921,N_10247,N_10565);
and U11922 (N_11922,N_10541,N_10993);
and U11923 (N_11923,N_10275,N_10747);
or U11924 (N_11924,N_10506,N_10018);
xnor U11925 (N_11925,N_10784,N_10164);
xor U11926 (N_11926,N_10250,N_10118);
and U11927 (N_11927,N_10783,N_10508);
xnor U11928 (N_11928,N_10318,N_10231);
and U11929 (N_11929,N_10502,N_10864);
or U11930 (N_11930,N_10744,N_10367);
or U11931 (N_11931,N_10992,N_10212);
and U11932 (N_11932,N_10725,N_10797);
and U11933 (N_11933,N_10822,N_10876);
or U11934 (N_11934,N_10837,N_10067);
nand U11935 (N_11935,N_10158,N_10776);
or U11936 (N_11936,N_10586,N_10417);
and U11937 (N_11937,N_10123,N_10428);
xnor U11938 (N_11938,N_10921,N_10601);
nand U11939 (N_11939,N_10160,N_10747);
nand U11940 (N_11940,N_10729,N_10587);
nand U11941 (N_11941,N_10909,N_10114);
or U11942 (N_11942,N_10858,N_10940);
or U11943 (N_11943,N_10912,N_10237);
nor U11944 (N_11944,N_10020,N_10788);
nor U11945 (N_11945,N_10928,N_10410);
nor U11946 (N_11946,N_10052,N_10193);
nand U11947 (N_11947,N_10399,N_10336);
nor U11948 (N_11948,N_10585,N_10694);
xnor U11949 (N_11949,N_10930,N_10149);
and U11950 (N_11950,N_10652,N_10194);
nor U11951 (N_11951,N_10442,N_10432);
nand U11952 (N_11952,N_10781,N_10695);
nor U11953 (N_11953,N_10600,N_10170);
or U11954 (N_11954,N_10134,N_10212);
and U11955 (N_11955,N_10696,N_10375);
or U11956 (N_11956,N_10060,N_10451);
nand U11957 (N_11957,N_10984,N_10465);
nor U11958 (N_11958,N_10799,N_10040);
xnor U11959 (N_11959,N_10004,N_10679);
nor U11960 (N_11960,N_10723,N_10919);
and U11961 (N_11961,N_10050,N_10080);
or U11962 (N_11962,N_10318,N_10363);
nand U11963 (N_11963,N_10474,N_10996);
nor U11964 (N_11964,N_10899,N_10647);
and U11965 (N_11965,N_10190,N_10494);
xnor U11966 (N_11966,N_10614,N_10914);
nor U11967 (N_11967,N_10948,N_10707);
nand U11968 (N_11968,N_10861,N_10974);
and U11969 (N_11969,N_10509,N_10490);
nand U11970 (N_11970,N_10728,N_10218);
and U11971 (N_11971,N_10616,N_10118);
nand U11972 (N_11972,N_10687,N_10252);
xor U11973 (N_11973,N_10592,N_10944);
or U11974 (N_11974,N_10589,N_10931);
xnor U11975 (N_11975,N_10745,N_10035);
nand U11976 (N_11976,N_10374,N_10133);
xor U11977 (N_11977,N_10976,N_10704);
nand U11978 (N_11978,N_10095,N_10349);
nand U11979 (N_11979,N_10356,N_10545);
nor U11980 (N_11980,N_10528,N_10189);
or U11981 (N_11981,N_10844,N_10117);
and U11982 (N_11982,N_10669,N_10382);
xnor U11983 (N_11983,N_10964,N_10186);
or U11984 (N_11984,N_10533,N_10840);
and U11985 (N_11985,N_10406,N_10485);
xor U11986 (N_11986,N_10786,N_10280);
nor U11987 (N_11987,N_10337,N_10283);
and U11988 (N_11988,N_10382,N_10356);
nor U11989 (N_11989,N_10085,N_10535);
xor U11990 (N_11990,N_10151,N_10576);
nor U11991 (N_11991,N_10420,N_10146);
xnor U11992 (N_11992,N_10067,N_10254);
nor U11993 (N_11993,N_10144,N_10233);
nor U11994 (N_11994,N_10521,N_10499);
xnor U11995 (N_11995,N_10368,N_10768);
and U11996 (N_11996,N_10354,N_10649);
nor U11997 (N_11997,N_10342,N_10333);
and U11998 (N_11998,N_10045,N_10713);
and U11999 (N_11999,N_10501,N_10852);
nand U12000 (N_12000,N_11970,N_11533);
nor U12001 (N_12001,N_11485,N_11556);
nor U12002 (N_12002,N_11255,N_11842);
or U12003 (N_12003,N_11264,N_11840);
xnor U12004 (N_12004,N_11861,N_11890);
nor U12005 (N_12005,N_11241,N_11321);
nor U12006 (N_12006,N_11636,N_11425);
and U12007 (N_12007,N_11333,N_11590);
or U12008 (N_12008,N_11178,N_11462);
and U12009 (N_12009,N_11597,N_11516);
and U12010 (N_12010,N_11390,N_11375);
nand U12011 (N_12011,N_11608,N_11641);
and U12012 (N_12012,N_11669,N_11719);
nand U12013 (N_12013,N_11739,N_11176);
or U12014 (N_12014,N_11549,N_11077);
nand U12015 (N_12015,N_11596,N_11272);
xor U12016 (N_12016,N_11878,N_11023);
or U12017 (N_12017,N_11835,N_11013);
or U12018 (N_12018,N_11459,N_11155);
xnor U12019 (N_12019,N_11100,N_11429);
nand U12020 (N_12020,N_11771,N_11406);
nor U12021 (N_12021,N_11723,N_11611);
or U12022 (N_12022,N_11296,N_11256);
or U12023 (N_12023,N_11607,N_11610);
nor U12024 (N_12024,N_11804,N_11671);
nor U12025 (N_12025,N_11331,N_11754);
or U12026 (N_12026,N_11644,N_11779);
nor U12027 (N_12027,N_11547,N_11986);
and U12028 (N_12028,N_11961,N_11686);
nor U12029 (N_12029,N_11589,N_11504);
xnor U12030 (N_12030,N_11713,N_11833);
nor U12031 (N_12031,N_11123,N_11904);
nor U12032 (N_12032,N_11034,N_11867);
and U12033 (N_12033,N_11768,N_11481);
or U12034 (N_12034,N_11870,N_11548);
nor U12035 (N_12035,N_11653,N_11679);
nand U12036 (N_12036,N_11287,N_11758);
nand U12037 (N_12037,N_11344,N_11220);
or U12038 (N_12038,N_11352,N_11917);
nor U12039 (N_12039,N_11216,N_11612);
nor U12040 (N_12040,N_11638,N_11434);
xor U12041 (N_12041,N_11475,N_11985);
nor U12042 (N_12042,N_11422,N_11588);
nor U12043 (N_12043,N_11524,N_11347);
xor U12044 (N_12044,N_11138,N_11189);
nand U12045 (N_12045,N_11722,N_11351);
and U12046 (N_12046,N_11319,N_11677);
nand U12047 (N_12047,N_11634,N_11091);
or U12048 (N_12048,N_11799,N_11205);
xor U12049 (N_12049,N_11260,N_11693);
or U12050 (N_12050,N_11909,N_11057);
nand U12051 (N_12051,N_11831,N_11322);
nand U12052 (N_12052,N_11295,N_11177);
nor U12053 (N_12053,N_11194,N_11349);
nor U12054 (N_12054,N_11281,N_11223);
or U12055 (N_12055,N_11912,N_11106);
nor U12056 (N_12056,N_11685,N_11619);
nor U12057 (N_12057,N_11578,N_11594);
nand U12058 (N_12058,N_11926,N_11795);
or U12059 (N_12059,N_11030,N_11164);
and U12060 (N_12060,N_11550,N_11838);
and U12061 (N_12061,N_11440,N_11311);
xnor U12062 (N_12062,N_11740,N_11149);
xor U12063 (N_12063,N_11665,N_11412);
nand U12064 (N_12064,N_11134,N_11334);
nand U12065 (N_12065,N_11435,N_11101);
and U12066 (N_12066,N_11121,N_11217);
or U12067 (N_12067,N_11797,N_11328);
and U12068 (N_12068,N_11206,N_11666);
nor U12069 (N_12069,N_11947,N_11345);
or U12070 (N_12070,N_11169,N_11744);
nand U12071 (N_12071,N_11512,N_11212);
or U12072 (N_12072,N_11284,N_11600);
nor U12073 (N_12073,N_11315,N_11496);
nand U12074 (N_12074,N_11561,N_11704);
and U12075 (N_12075,N_11125,N_11983);
nor U12076 (N_12076,N_11268,N_11239);
xor U12077 (N_12077,N_11989,N_11336);
nand U12078 (N_12078,N_11866,N_11881);
and U12079 (N_12079,N_11160,N_11076);
and U12080 (N_12080,N_11577,N_11625);
xor U12081 (N_12081,N_11183,N_11477);
and U12082 (N_12082,N_11772,N_11718);
and U12083 (N_12083,N_11522,N_11729);
and U12084 (N_12084,N_11844,N_11828);
or U12085 (N_12085,N_11752,N_11492);
and U12086 (N_12086,N_11252,N_11409);
and U12087 (N_12087,N_11497,N_11676);
nor U12088 (N_12088,N_11499,N_11179);
and U12089 (N_12089,N_11014,N_11171);
or U12090 (N_12090,N_11895,N_11364);
nand U12091 (N_12091,N_11692,N_11456);
nor U12092 (N_12092,N_11040,N_11506);
or U12093 (N_12093,N_11716,N_11660);
xnor U12094 (N_12094,N_11300,N_11438);
or U12095 (N_12095,N_11308,N_11172);
or U12096 (N_12096,N_11789,N_11130);
nand U12097 (N_12097,N_11952,N_11615);
and U12098 (N_12098,N_11996,N_11568);
or U12099 (N_12099,N_11663,N_11508);
xnor U12100 (N_12100,N_11051,N_11025);
nor U12101 (N_12101,N_11544,N_11717);
nand U12102 (N_12102,N_11529,N_11817);
and U12103 (N_12103,N_11307,N_11855);
nor U12104 (N_12104,N_11363,N_11543);
or U12105 (N_12105,N_11756,N_11994);
and U12106 (N_12106,N_11736,N_11628);
xnor U12107 (N_12107,N_11055,N_11312);
nor U12108 (N_12108,N_11401,N_11063);
or U12109 (N_12109,N_11118,N_11960);
xnor U12110 (N_12110,N_11237,N_11498);
xnor U12111 (N_12111,N_11436,N_11503);
and U12112 (N_12112,N_11525,N_11876);
and U12113 (N_12113,N_11320,N_11127);
and U12114 (N_12114,N_11251,N_11187);
xor U12115 (N_12115,N_11366,N_11270);
or U12116 (N_12116,N_11073,N_11111);
or U12117 (N_12117,N_11203,N_11813);
and U12118 (N_12118,N_11210,N_11579);
or U12119 (N_12119,N_11786,N_11208);
nor U12120 (N_12120,N_11727,N_11493);
or U12121 (N_12121,N_11099,N_11166);
or U12122 (N_12122,N_11301,N_11119);
nand U12123 (N_12123,N_11884,N_11468);
and U12124 (N_12124,N_11648,N_11185);
xnor U12125 (N_12125,N_11621,N_11816);
xor U12126 (N_12126,N_11937,N_11690);
nor U12127 (N_12127,N_11879,N_11293);
xnor U12128 (N_12128,N_11053,N_11068);
or U12129 (N_12129,N_11150,N_11583);
nor U12130 (N_12130,N_11658,N_11822);
nor U12131 (N_12131,N_11473,N_11773);
nand U12132 (N_12132,N_11661,N_11152);
xor U12133 (N_12133,N_11464,N_11193);
or U12134 (N_12134,N_11195,N_11829);
and U12135 (N_12135,N_11248,N_11888);
nand U12136 (N_12136,N_11931,N_11291);
nand U12137 (N_12137,N_11065,N_11467);
nand U12138 (N_12138,N_11234,N_11274);
or U12139 (N_12139,N_11219,N_11017);
xor U12140 (N_12140,N_11389,N_11749);
nand U12141 (N_12141,N_11624,N_11142);
or U12142 (N_12142,N_11998,N_11601);
nor U12143 (N_12143,N_11755,N_11081);
nand U12144 (N_12144,N_11592,N_11342);
nor U12145 (N_12145,N_11942,N_11980);
or U12146 (N_12146,N_11928,N_11972);
or U12147 (N_12147,N_11458,N_11002);
nand U12148 (N_12148,N_11957,N_11886);
nor U12149 (N_12149,N_11113,N_11827);
nand U12150 (N_12150,N_11896,N_11188);
nor U12151 (N_12151,N_11585,N_11026);
xor U12152 (N_12152,N_11446,N_11262);
nand U12153 (N_12153,N_11447,N_11486);
and U12154 (N_12154,N_11104,N_11376);
nor U12155 (N_12155,N_11997,N_11096);
and U12156 (N_12156,N_11557,N_11297);
nor U12157 (N_12157,N_11213,N_11442);
nor U12158 (N_12158,N_11482,N_11891);
nand U12159 (N_12159,N_11403,N_11286);
nand U12160 (N_12160,N_11863,N_11837);
nand U12161 (N_12161,N_11108,N_11606);
or U12162 (N_12162,N_11011,N_11684);
nand U12163 (N_12163,N_11805,N_11654);
or U12164 (N_12164,N_11292,N_11480);
and U12165 (N_12165,N_11581,N_11043);
and U12166 (N_12166,N_11027,N_11536);
and U12167 (N_12167,N_11747,N_11484);
or U12168 (N_12168,N_11427,N_11028);
xnor U12169 (N_12169,N_11703,N_11354);
or U12170 (N_12170,N_11472,N_11453);
xnor U12171 (N_12171,N_11925,N_11775);
nand U12172 (N_12172,N_11316,N_11818);
and U12173 (N_12173,N_11132,N_11538);
nor U12174 (N_12174,N_11507,N_11770);
or U12175 (N_12175,N_11198,N_11211);
nand U12176 (N_12176,N_11318,N_11602);
xor U12177 (N_12177,N_11964,N_11117);
or U12178 (N_12178,N_11563,N_11276);
xnor U12179 (N_12179,N_11680,N_11725);
nand U12180 (N_12180,N_11258,N_11359);
xnor U12181 (N_12181,N_11204,N_11079);
nand U12182 (N_12182,N_11593,N_11921);
xor U12183 (N_12183,N_11324,N_11042);
nand U12184 (N_12184,N_11552,N_11672);
xnor U12185 (N_12185,N_11901,N_11558);
nor U12186 (N_12186,N_11800,N_11097);
or U12187 (N_12187,N_11167,N_11109);
nand U12188 (N_12188,N_11854,N_11760);
xor U12189 (N_12189,N_11992,N_11706);
xnor U12190 (N_12190,N_11977,N_11987);
nor U12191 (N_12191,N_11033,N_11869);
and U12192 (N_12192,N_11708,N_11646);
nand U12193 (N_12193,N_11174,N_11820);
xnor U12194 (N_12194,N_11218,N_11378);
nor U12195 (N_12195,N_11728,N_11629);
xnor U12196 (N_12196,N_11790,N_11133);
xnor U12197 (N_12197,N_11059,N_11801);
xor U12198 (N_12198,N_11072,N_11807);
or U12199 (N_12199,N_11955,N_11124);
and U12200 (N_12200,N_11720,N_11207);
and U12201 (N_12201,N_11882,N_11959);
or U12202 (N_12202,N_11225,N_11061);
nand U12203 (N_12203,N_11031,N_11979);
or U12204 (N_12204,N_11787,N_11044);
nor U12205 (N_12205,N_11340,N_11916);
and U12206 (N_12206,N_11085,N_11929);
nor U12207 (N_12207,N_11698,N_11022);
xnor U12208 (N_12208,N_11735,N_11452);
nand U12209 (N_12209,N_11365,N_11696);
and U12210 (N_12210,N_11656,N_11982);
or U12211 (N_12211,N_11060,N_11834);
xor U12212 (N_12212,N_11510,N_11443);
xor U12213 (N_12213,N_11938,N_11299);
nand U12214 (N_12214,N_11711,N_11399);
and U12215 (N_12215,N_11785,N_11338);
nand U12216 (N_12216,N_11353,N_11930);
nand U12217 (N_12217,N_11794,N_11415);
or U12218 (N_12218,N_11701,N_11488);
nor U12219 (N_12219,N_11247,N_11675);
xnor U12220 (N_12220,N_11466,N_11039);
nand U12221 (N_12221,N_11843,N_11531);
xnor U12222 (N_12222,N_11457,N_11521);
nor U12223 (N_12223,N_11657,N_11010);
or U12224 (N_12224,N_11250,N_11131);
xnor U12225 (N_12225,N_11962,N_11483);
nand U12226 (N_12226,N_11846,N_11971);
nor U12227 (N_12227,N_11240,N_11872);
or U12228 (N_12228,N_11215,N_11433);
nor U12229 (N_12229,N_11598,N_11518);
or U12230 (N_12230,N_11086,N_11991);
and U12231 (N_12231,N_11190,N_11731);
nand U12232 (N_12232,N_11377,N_11271);
nor U12233 (N_12233,N_11224,N_11070);
nand U12234 (N_12234,N_11859,N_11393);
or U12235 (N_12235,N_11753,N_11877);
xnor U12236 (N_12236,N_11571,N_11249);
nor U12237 (N_12237,N_11988,N_11927);
and U12238 (N_12238,N_11082,N_11186);
nor U12239 (N_12239,N_11047,N_11586);
or U12240 (N_12240,N_11120,N_11562);
xor U12241 (N_12241,N_11226,N_11003);
and U12242 (N_12242,N_11535,N_11802);
xor U12243 (N_12243,N_11726,N_11936);
xor U12244 (N_12244,N_11759,N_11280);
nor U12245 (N_12245,N_11058,N_11180);
or U12246 (N_12246,N_11900,N_11932);
and U12247 (N_12247,N_11724,N_11441);
nor U12248 (N_12248,N_11181,N_11575);
and U12249 (N_12249,N_11490,N_11954);
or U12250 (N_12250,N_11647,N_11574);
and U12251 (N_12251,N_11655,N_11437);
and U12252 (N_12252,N_11761,N_11098);
nand U12253 (N_12253,N_11545,N_11275);
and U12254 (N_12254,N_11361,N_11856);
nand U12255 (N_12255,N_11981,N_11871);
nor U12256 (N_12256,N_11192,N_11815);
nand U12257 (N_12257,N_11537,N_11089);
and U12258 (N_12258,N_11469,N_11559);
or U12259 (N_12259,N_11920,N_11470);
nand U12260 (N_12260,N_11824,N_11384);
xor U12261 (N_12261,N_11501,N_11388);
and U12262 (N_12262,N_11071,N_11000);
and U12263 (N_12263,N_11107,N_11635);
or U12264 (N_12264,N_11963,N_11967);
and U12265 (N_12265,N_11673,N_11652);
nor U12266 (N_12266,N_11509,N_11862);
nand U12267 (N_12267,N_11054,N_11392);
nand U12268 (N_12268,N_11062,N_11742);
nor U12269 (N_12269,N_11569,N_11128);
or U12270 (N_12270,N_11709,N_11745);
nor U12271 (N_12271,N_11200,N_11806);
nand U12272 (N_12272,N_11683,N_11451);
xnor U12273 (N_12273,N_11651,N_11605);
nand U12274 (N_12274,N_11329,N_11623);
and U12275 (N_12275,N_11848,N_11001);
or U12276 (N_12276,N_11715,N_11781);
nor U12277 (N_12277,N_11630,N_11631);
nand U12278 (N_12278,N_11956,N_11554);
nor U12279 (N_12279,N_11514,N_11139);
and U12280 (N_12280,N_11609,N_11461);
xnor U12281 (N_12281,N_11893,N_11784);
xnor U12282 (N_12282,N_11305,N_11924);
and U12283 (N_12283,N_11943,N_11694);
nand U12284 (N_12284,N_11935,N_11236);
or U12285 (N_12285,N_11933,N_11905);
nor U12286 (N_12286,N_11515,N_11094);
xor U12287 (N_12287,N_11404,N_11821);
xor U12288 (N_12288,N_11774,N_11337);
and U12289 (N_12289,N_11748,N_11019);
or U12290 (N_12290,N_11009,N_11021);
or U12291 (N_12291,N_11148,N_11112);
and U12292 (N_12292,N_11809,N_11595);
or U12293 (N_12293,N_11135,N_11478);
and U12294 (N_12294,N_11587,N_11910);
nor U12295 (N_12295,N_11162,N_11463);
or U12296 (N_12296,N_11783,N_11491);
nor U12297 (N_12297,N_11542,N_11147);
or U12298 (N_12298,N_11012,N_11432);
and U12299 (N_12299,N_11914,N_11369);
nor U12300 (N_12300,N_11494,N_11778);
or U12301 (N_12301,N_11941,N_11650);
xnor U12302 (N_12302,N_11093,N_11165);
nand U12303 (N_12303,N_11883,N_11505);
and U12304 (N_12304,N_11567,N_11479);
xnor U12305 (N_12305,N_11279,N_11145);
and U12306 (N_12306,N_11540,N_11911);
xnor U12307 (N_12307,N_11243,N_11046);
or U12308 (N_12308,N_11413,N_11898);
nor U12309 (N_12309,N_11004,N_11944);
nand U12310 (N_12310,N_11035,N_11371);
or U12311 (N_12311,N_11143,N_11343);
xnor U12312 (N_12312,N_11974,N_11632);
nand U12313 (N_12313,N_11394,N_11776);
xnor U12314 (N_12314,N_11417,N_11370);
nand U12315 (N_12315,N_11868,N_11122);
and U12316 (N_12316,N_11024,N_11897);
nor U12317 (N_12317,N_11730,N_11126);
or U12318 (N_12318,N_11572,N_11330);
xor U12319 (N_12319,N_11140,N_11990);
or U12320 (N_12320,N_11945,N_11313);
xnor U12321 (N_12321,N_11519,N_11083);
and U12322 (N_12322,N_11793,N_11923);
nand U12323 (N_12323,N_11700,N_11721);
and U12324 (N_12324,N_11699,N_11277);
xor U12325 (N_12325,N_11476,N_11254);
or U12326 (N_12326,N_11845,N_11282);
or U12327 (N_12327,N_11428,N_11555);
and U12328 (N_12328,N_11408,N_11880);
nand U12329 (N_12329,N_11642,N_11407);
nor U12330 (N_12330,N_11908,N_11431);
xor U12331 (N_12331,N_11667,N_11156);
nand U12332 (N_12332,N_11095,N_11391);
and U12333 (N_12333,N_11853,N_11018);
or U12334 (N_12334,N_11858,N_11674);
nand U12335 (N_12335,N_11530,N_11064);
and U12336 (N_12336,N_11873,N_11450);
nand U12337 (N_12337,N_11424,N_11633);
or U12338 (N_12338,N_11751,N_11439);
nand U12339 (N_12339,N_11278,N_11887);
nand U12340 (N_12340,N_11373,N_11227);
or U12341 (N_12341,N_11015,N_11687);
nand U12342 (N_12342,N_11528,N_11103);
and U12343 (N_12343,N_11154,N_11310);
nor U12344 (N_12344,N_11714,N_11067);
nor U12345 (N_12345,N_11416,N_11546);
or U12346 (N_12346,N_11420,N_11688);
nor U12347 (N_12347,N_11743,N_11454);
xor U12348 (N_12348,N_11993,N_11426);
nor U12349 (N_12349,N_11852,N_11105);
xor U12350 (N_12350,N_11288,N_11201);
or U12351 (N_12351,N_11539,N_11746);
nor U12352 (N_12352,N_11196,N_11520);
xor U12353 (N_12353,N_11839,N_11153);
xnor U12354 (N_12354,N_11966,N_11697);
or U12355 (N_12355,N_11640,N_11173);
or U12356 (N_12356,N_11814,N_11832);
or U12357 (N_12357,N_11137,N_11048);
xnor U12358 (N_12358,N_11526,N_11757);
nor U12359 (N_12359,N_11209,N_11616);
or U12360 (N_12360,N_11163,N_11517);
nand U12361 (N_12361,N_11007,N_11362);
and U12362 (N_12362,N_11235,N_11622);
nor U12363 (N_12363,N_11037,N_11907);
xor U12364 (N_12364,N_11626,N_11769);
xnor U12365 (N_12365,N_11591,N_11681);
xnor U12366 (N_12366,N_11005,N_11245);
nor U12367 (N_12367,N_11965,N_11639);
xor U12368 (N_12368,N_11702,N_11599);
or U12369 (N_12369,N_11474,N_11242);
or U12370 (N_12370,N_11874,N_11302);
or U12371 (N_12371,N_11500,N_11144);
and U12372 (N_12372,N_11682,N_11885);
xnor U12373 (N_12373,N_11341,N_11306);
or U12374 (N_12374,N_11662,N_11823);
nor U12375 (N_12375,N_11032,N_11949);
nand U12376 (N_12376,N_11903,N_11129);
nand U12377 (N_12377,N_11875,N_11465);
nor U12378 (N_12378,N_11762,N_11382);
nand U12379 (N_12379,N_11819,N_11946);
nand U12380 (N_12380,N_11267,N_11767);
xnor U12381 (N_12381,N_11304,N_11527);
nand U12382 (N_12382,N_11290,N_11159);
nor U12383 (N_12383,N_11049,N_11455);
nor U12384 (N_12384,N_11976,N_11738);
and U12385 (N_12385,N_11798,N_11263);
nand U12386 (N_12386,N_11741,N_11826);
nand U12387 (N_12387,N_11939,N_11289);
xnor U12388 (N_12388,N_11020,N_11202);
xnor U12389 (N_12389,N_11421,N_11614);
nor U12390 (N_12390,N_11968,N_11008);
nor U12391 (N_12391,N_11116,N_11448);
nand U12392 (N_12392,N_11618,N_11511);
nand U12393 (N_12393,N_11471,N_11765);
and U12394 (N_12394,N_11849,N_11184);
xnor U12395 (N_12395,N_11732,N_11582);
or U12396 (N_12396,N_11847,N_11913);
nor U12397 (N_12397,N_11782,N_11906);
nor U12398 (N_12398,N_11788,N_11750);
and U12399 (N_12399,N_11995,N_11273);
nand U12400 (N_12400,N_11360,N_11984);
nand U12401 (N_12401,N_11553,N_11229);
or U12402 (N_12402,N_11405,N_11707);
and U12403 (N_12403,N_11257,N_11523);
nand U12404 (N_12404,N_11006,N_11951);
and U12405 (N_12405,N_11764,N_11418);
and U12406 (N_12406,N_11102,N_11411);
and U12407 (N_12407,N_11052,N_11825);
and U12408 (N_12408,N_11573,N_11266);
or U12409 (N_12409,N_11170,N_11830);
nor U12410 (N_12410,N_11811,N_11691);
xor U12411 (N_12411,N_11565,N_11075);
nand U12412 (N_12412,N_11269,N_11386);
or U12413 (N_12413,N_11689,N_11380);
nand U12414 (N_12414,N_11069,N_11078);
and U12415 (N_12415,N_11766,N_11038);
xnor U12416 (N_12416,N_11230,N_11576);
nand U12417 (N_12417,N_11357,N_11780);
and U12418 (N_12418,N_11645,N_11368);
and U12419 (N_12419,N_11265,N_11036);
or U12420 (N_12420,N_11950,N_11110);
nand U12421 (N_12421,N_11402,N_11090);
or U12422 (N_12422,N_11733,N_11080);
nand U12423 (N_12423,N_11566,N_11796);
and U12424 (N_12424,N_11383,N_11151);
xnor U12425 (N_12425,N_11953,N_11710);
or U12426 (N_12426,N_11041,N_11604);
nand U12427 (N_12427,N_11356,N_11191);
and U12428 (N_12428,N_11303,N_11620);
or U12429 (N_12429,N_11367,N_11643);
nand U12430 (N_12430,N_11763,N_11808);
or U12431 (N_12431,N_11670,N_11734);
and U12432 (N_12432,N_11973,N_11836);
and U12433 (N_12433,N_11294,N_11915);
xor U12434 (N_12434,N_11326,N_11850);
xor U12435 (N_12435,N_11232,N_11355);
or U12436 (N_12436,N_11387,N_11812);
nand U12437 (N_12437,N_11864,N_11902);
nor U12438 (N_12438,N_11146,N_11199);
or U12439 (N_12439,N_11115,N_11580);
nand U12440 (N_12440,N_11397,N_11214);
nand U12441 (N_12441,N_11114,N_11841);
xor U12442 (N_12442,N_11627,N_11016);
nand U12443 (N_12443,N_11705,N_11975);
nand U12444 (N_12444,N_11637,N_11560);
nor U12445 (N_12445,N_11158,N_11233);
or U12446 (N_12446,N_11074,N_11737);
nand U12447 (N_12447,N_11851,N_11430);
nand U12448 (N_12448,N_11541,N_11374);
nand U12449 (N_12449,N_11379,N_11892);
or U12450 (N_12450,N_11045,N_11958);
xnor U12451 (N_12451,N_11396,N_11253);
nand U12452 (N_12452,N_11285,N_11414);
and U12453 (N_12453,N_11502,N_11584);
nand U12454 (N_12454,N_11445,N_11029);
nand U12455 (N_12455,N_11810,N_11860);
xor U12456 (N_12456,N_11978,N_11712);
and U12457 (N_12457,N_11066,N_11603);
nand U12458 (N_12458,N_11792,N_11317);
xnor U12459 (N_12459,N_11400,N_11613);
xor U12460 (N_12460,N_11259,N_11157);
or U12461 (N_12461,N_11570,N_11261);
nor U12462 (N_12462,N_11350,N_11934);
nand U12463 (N_12463,N_11136,N_11088);
and U12464 (N_12464,N_11668,N_11327);
xor U12465 (N_12465,N_11050,N_11948);
nand U12466 (N_12466,N_11339,N_11298);
xnor U12467 (N_12467,N_11649,N_11084);
or U12468 (N_12468,N_11513,N_11564);
xor U12469 (N_12469,N_11495,N_11919);
nor U12470 (N_12470,N_11395,N_11161);
and U12471 (N_12471,N_11175,N_11419);
xnor U12472 (N_12472,N_11894,N_11940);
nand U12473 (N_12473,N_11332,N_11489);
and U12474 (N_12474,N_11664,N_11056);
nor U12475 (N_12475,N_11534,N_11325);
nor U12476 (N_12476,N_11410,N_11969);
and U12477 (N_12477,N_11791,N_11182);
nor U12478 (N_12478,N_11551,N_11449);
xnor U12479 (N_12479,N_11857,N_11348);
nor U12480 (N_12480,N_11889,N_11777);
nand U12481 (N_12481,N_11358,N_11246);
nand U12482 (N_12482,N_11398,N_11228);
and U12483 (N_12483,N_11346,N_11087);
xor U12484 (N_12484,N_11423,N_11238);
nor U12485 (N_12485,N_11381,N_11918);
nand U12486 (N_12486,N_11283,N_11922);
nand U12487 (N_12487,N_11231,N_11309);
nand U12488 (N_12488,N_11617,N_11659);
nor U12489 (N_12489,N_11487,N_11372);
or U12490 (N_12490,N_11244,N_11865);
or U12491 (N_12491,N_11221,N_11695);
and U12492 (N_12492,N_11168,N_11323);
xor U12493 (N_12493,N_11899,N_11678);
and U12494 (N_12494,N_11222,N_11803);
nand U12495 (N_12495,N_11197,N_11460);
nand U12496 (N_12496,N_11385,N_11314);
and U12497 (N_12497,N_11444,N_11092);
xor U12498 (N_12498,N_11335,N_11141);
nand U12499 (N_12499,N_11999,N_11532);
xnor U12500 (N_12500,N_11356,N_11371);
nor U12501 (N_12501,N_11002,N_11584);
xnor U12502 (N_12502,N_11716,N_11439);
and U12503 (N_12503,N_11307,N_11025);
or U12504 (N_12504,N_11100,N_11673);
nand U12505 (N_12505,N_11927,N_11150);
xnor U12506 (N_12506,N_11632,N_11840);
xnor U12507 (N_12507,N_11418,N_11718);
nand U12508 (N_12508,N_11152,N_11465);
nand U12509 (N_12509,N_11862,N_11944);
xnor U12510 (N_12510,N_11091,N_11895);
nand U12511 (N_12511,N_11880,N_11667);
nand U12512 (N_12512,N_11369,N_11131);
xnor U12513 (N_12513,N_11058,N_11017);
nor U12514 (N_12514,N_11705,N_11417);
xnor U12515 (N_12515,N_11146,N_11945);
and U12516 (N_12516,N_11020,N_11302);
nand U12517 (N_12517,N_11508,N_11630);
xor U12518 (N_12518,N_11780,N_11086);
and U12519 (N_12519,N_11979,N_11680);
or U12520 (N_12520,N_11175,N_11028);
xor U12521 (N_12521,N_11499,N_11044);
or U12522 (N_12522,N_11046,N_11584);
nand U12523 (N_12523,N_11531,N_11713);
nand U12524 (N_12524,N_11764,N_11154);
nand U12525 (N_12525,N_11279,N_11913);
or U12526 (N_12526,N_11012,N_11078);
nor U12527 (N_12527,N_11135,N_11466);
nor U12528 (N_12528,N_11395,N_11524);
and U12529 (N_12529,N_11020,N_11050);
nand U12530 (N_12530,N_11586,N_11085);
and U12531 (N_12531,N_11485,N_11887);
and U12532 (N_12532,N_11230,N_11441);
or U12533 (N_12533,N_11124,N_11462);
and U12534 (N_12534,N_11045,N_11215);
or U12535 (N_12535,N_11028,N_11412);
and U12536 (N_12536,N_11645,N_11432);
and U12537 (N_12537,N_11560,N_11814);
nand U12538 (N_12538,N_11182,N_11121);
or U12539 (N_12539,N_11800,N_11108);
nor U12540 (N_12540,N_11638,N_11142);
nor U12541 (N_12541,N_11463,N_11968);
nand U12542 (N_12542,N_11969,N_11752);
nand U12543 (N_12543,N_11373,N_11854);
and U12544 (N_12544,N_11888,N_11157);
xnor U12545 (N_12545,N_11450,N_11565);
or U12546 (N_12546,N_11272,N_11420);
xor U12547 (N_12547,N_11968,N_11098);
and U12548 (N_12548,N_11888,N_11005);
and U12549 (N_12549,N_11118,N_11861);
and U12550 (N_12550,N_11750,N_11254);
and U12551 (N_12551,N_11760,N_11809);
and U12552 (N_12552,N_11227,N_11277);
and U12553 (N_12553,N_11458,N_11282);
nand U12554 (N_12554,N_11673,N_11775);
and U12555 (N_12555,N_11280,N_11365);
nand U12556 (N_12556,N_11786,N_11133);
nor U12557 (N_12557,N_11850,N_11958);
xor U12558 (N_12558,N_11190,N_11786);
or U12559 (N_12559,N_11046,N_11746);
nor U12560 (N_12560,N_11573,N_11206);
nor U12561 (N_12561,N_11591,N_11528);
nor U12562 (N_12562,N_11007,N_11662);
xnor U12563 (N_12563,N_11864,N_11559);
nor U12564 (N_12564,N_11202,N_11171);
xor U12565 (N_12565,N_11633,N_11396);
and U12566 (N_12566,N_11994,N_11641);
or U12567 (N_12567,N_11697,N_11239);
nand U12568 (N_12568,N_11428,N_11436);
nor U12569 (N_12569,N_11663,N_11024);
and U12570 (N_12570,N_11693,N_11227);
or U12571 (N_12571,N_11353,N_11732);
nor U12572 (N_12572,N_11365,N_11418);
nor U12573 (N_12573,N_11776,N_11161);
and U12574 (N_12574,N_11072,N_11116);
xnor U12575 (N_12575,N_11314,N_11479);
nand U12576 (N_12576,N_11294,N_11843);
or U12577 (N_12577,N_11937,N_11535);
xor U12578 (N_12578,N_11210,N_11792);
nor U12579 (N_12579,N_11406,N_11994);
nor U12580 (N_12580,N_11972,N_11396);
xnor U12581 (N_12581,N_11257,N_11186);
or U12582 (N_12582,N_11045,N_11201);
xor U12583 (N_12583,N_11337,N_11910);
xor U12584 (N_12584,N_11535,N_11234);
nand U12585 (N_12585,N_11722,N_11256);
or U12586 (N_12586,N_11855,N_11550);
nand U12587 (N_12587,N_11664,N_11860);
nor U12588 (N_12588,N_11550,N_11108);
xor U12589 (N_12589,N_11674,N_11604);
and U12590 (N_12590,N_11218,N_11978);
xnor U12591 (N_12591,N_11948,N_11929);
and U12592 (N_12592,N_11586,N_11204);
xnor U12593 (N_12593,N_11264,N_11905);
xor U12594 (N_12594,N_11184,N_11042);
and U12595 (N_12595,N_11430,N_11762);
xor U12596 (N_12596,N_11898,N_11877);
xor U12597 (N_12597,N_11337,N_11176);
xor U12598 (N_12598,N_11056,N_11793);
or U12599 (N_12599,N_11855,N_11889);
or U12600 (N_12600,N_11077,N_11999);
nor U12601 (N_12601,N_11701,N_11639);
and U12602 (N_12602,N_11423,N_11606);
xnor U12603 (N_12603,N_11614,N_11623);
or U12604 (N_12604,N_11249,N_11803);
or U12605 (N_12605,N_11546,N_11150);
and U12606 (N_12606,N_11833,N_11093);
or U12607 (N_12607,N_11040,N_11333);
nor U12608 (N_12608,N_11936,N_11850);
nor U12609 (N_12609,N_11501,N_11902);
and U12610 (N_12610,N_11630,N_11400);
and U12611 (N_12611,N_11441,N_11081);
nor U12612 (N_12612,N_11311,N_11222);
nand U12613 (N_12613,N_11961,N_11081);
xor U12614 (N_12614,N_11481,N_11082);
nand U12615 (N_12615,N_11420,N_11704);
nor U12616 (N_12616,N_11253,N_11354);
nor U12617 (N_12617,N_11243,N_11789);
xnor U12618 (N_12618,N_11556,N_11913);
nor U12619 (N_12619,N_11900,N_11407);
nand U12620 (N_12620,N_11638,N_11125);
nand U12621 (N_12621,N_11692,N_11484);
xnor U12622 (N_12622,N_11712,N_11154);
nand U12623 (N_12623,N_11786,N_11776);
and U12624 (N_12624,N_11982,N_11019);
xor U12625 (N_12625,N_11975,N_11790);
or U12626 (N_12626,N_11725,N_11545);
nand U12627 (N_12627,N_11448,N_11089);
xnor U12628 (N_12628,N_11719,N_11000);
xnor U12629 (N_12629,N_11998,N_11944);
nand U12630 (N_12630,N_11898,N_11436);
xnor U12631 (N_12631,N_11828,N_11398);
or U12632 (N_12632,N_11787,N_11382);
and U12633 (N_12633,N_11715,N_11608);
or U12634 (N_12634,N_11549,N_11308);
or U12635 (N_12635,N_11856,N_11921);
nand U12636 (N_12636,N_11382,N_11465);
or U12637 (N_12637,N_11821,N_11630);
xnor U12638 (N_12638,N_11612,N_11953);
xnor U12639 (N_12639,N_11089,N_11011);
nor U12640 (N_12640,N_11559,N_11113);
nor U12641 (N_12641,N_11118,N_11457);
nor U12642 (N_12642,N_11846,N_11083);
or U12643 (N_12643,N_11450,N_11629);
nand U12644 (N_12644,N_11085,N_11579);
or U12645 (N_12645,N_11430,N_11188);
xnor U12646 (N_12646,N_11030,N_11341);
and U12647 (N_12647,N_11527,N_11861);
xnor U12648 (N_12648,N_11791,N_11613);
or U12649 (N_12649,N_11843,N_11670);
or U12650 (N_12650,N_11928,N_11777);
xnor U12651 (N_12651,N_11386,N_11080);
or U12652 (N_12652,N_11001,N_11463);
or U12653 (N_12653,N_11930,N_11064);
nand U12654 (N_12654,N_11255,N_11797);
xnor U12655 (N_12655,N_11482,N_11495);
nand U12656 (N_12656,N_11305,N_11390);
and U12657 (N_12657,N_11927,N_11604);
and U12658 (N_12658,N_11342,N_11078);
nor U12659 (N_12659,N_11373,N_11151);
nand U12660 (N_12660,N_11166,N_11141);
nand U12661 (N_12661,N_11570,N_11360);
or U12662 (N_12662,N_11573,N_11402);
nor U12663 (N_12663,N_11467,N_11296);
nand U12664 (N_12664,N_11912,N_11245);
or U12665 (N_12665,N_11205,N_11865);
and U12666 (N_12666,N_11372,N_11763);
and U12667 (N_12667,N_11101,N_11154);
xor U12668 (N_12668,N_11498,N_11649);
nand U12669 (N_12669,N_11590,N_11081);
nor U12670 (N_12670,N_11571,N_11306);
xnor U12671 (N_12671,N_11689,N_11166);
nand U12672 (N_12672,N_11334,N_11229);
or U12673 (N_12673,N_11357,N_11756);
and U12674 (N_12674,N_11787,N_11764);
and U12675 (N_12675,N_11644,N_11783);
nand U12676 (N_12676,N_11722,N_11123);
nor U12677 (N_12677,N_11220,N_11478);
and U12678 (N_12678,N_11881,N_11878);
xnor U12679 (N_12679,N_11064,N_11082);
xor U12680 (N_12680,N_11526,N_11225);
nor U12681 (N_12681,N_11924,N_11772);
and U12682 (N_12682,N_11541,N_11466);
xor U12683 (N_12683,N_11905,N_11731);
nor U12684 (N_12684,N_11881,N_11613);
nand U12685 (N_12685,N_11062,N_11705);
or U12686 (N_12686,N_11302,N_11089);
nand U12687 (N_12687,N_11744,N_11610);
nor U12688 (N_12688,N_11273,N_11326);
or U12689 (N_12689,N_11234,N_11177);
or U12690 (N_12690,N_11437,N_11859);
xnor U12691 (N_12691,N_11523,N_11600);
nand U12692 (N_12692,N_11395,N_11054);
or U12693 (N_12693,N_11626,N_11583);
xor U12694 (N_12694,N_11215,N_11670);
or U12695 (N_12695,N_11756,N_11637);
nand U12696 (N_12696,N_11214,N_11915);
nand U12697 (N_12697,N_11870,N_11451);
nor U12698 (N_12698,N_11675,N_11955);
or U12699 (N_12699,N_11546,N_11689);
and U12700 (N_12700,N_11229,N_11805);
and U12701 (N_12701,N_11243,N_11417);
and U12702 (N_12702,N_11774,N_11204);
nor U12703 (N_12703,N_11980,N_11589);
nor U12704 (N_12704,N_11951,N_11257);
and U12705 (N_12705,N_11479,N_11311);
nor U12706 (N_12706,N_11377,N_11765);
and U12707 (N_12707,N_11941,N_11785);
xor U12708 (N_12708,N_11860,N_11419);
or U12709 (N_12709,N_11545,N_11637);
nand U12710 (N_12710,N_11149,N_11817);
or U12711 (N_12711,N_11830,N_11690);
or U12712 (N_12712,N_11503,N_11210);
nand U12713 (N_12713,N_11385,N_11996);
xnor U12714 (N_12714,N_11655,N_11439);
and U12715 (N_12715,N_11536,N_11231);
nor U12716 (N_12716,N_11113,N_11567);
nor U12717 (N_12717,N_11425,N_11818);
nor U12718 (N_12718,N_11323,N_11607);
and U12719 (N_12719,N_11023,N_11802);
xor U12720 (N_12720,N_11268,N_11920);
nand U12721 (N_12721,N_11154,N_11427);
and U12722 (N_12722,N_11025,N_11283);
nand U12723 (N_12723,N_11565,N_11097);
and U12724 (N_12724,N_11366,N_11884);
nor U12725 (N_12725,N_11460,N_11643);
xor U12726 (N_12726,N_11925,N_11912);
nand U12727 (N_12727,N_11562,N_11225);
xor U12728 (N_12728,N_11925,N_11333);
nand U12729 (N_12729,N_11072,N_11675);
nor U12730 (N_12730,N_11750,N_11798);
and U12731 (N_12731,N_11222,N_11539);
nand U12732 (N_12732,N_11087,N_11269);
nor U12733 (N_12733,N_11869,N_11857);
and U12734 (N_12734,N_11996,N_11115);
xnor U12735 (N_12735,N_11966,N_11629);
nand U12736 (N_12736,N_11223,N_11412);
nor U12737 (N_12737,N_11043,N_11009);
and U12738 (N_12738,N_11068,N_11633);
or U12739 (N_12739,N_11693,N_11453);
xor U12740 (N_12740,N_11047,N_11088);
or U12741 (N_12741,N_11835,N_11310);
nand U12742 (N_12742,N_11348,N_11951);
nand U12743 (N_12743,N_11851,N_11265);
nor U12744 (N_12744,N_11813,N_11929);
xnor U12745 (N_12745,N_11823,N_11252);
and U12746 (N_12746,N_11232,N_11241);
or U12747 (N_12747,N_11223,N_11947);
and U12748 (N_12748,N_11627,N_11341);
nor U12749 (N_12749,N_11289,N_11082);
xnor U12750 (N_12750,N_11064,N_11381);
nor U12751 (N_12751,N_11982,N_11380);
nor U12752 (N_12752,N_11474,N_11772);
or U12753 (N_12753,N_11075,N_11643);
or U12754 (N_12754,N_11850,N_11915);
xor U12755 (N_12755,N_11073,N_11402);
nor U12756 (N_12756,N_11595,N_11138);
and U12757 (N_12757,N_11471,N_11382);
and U12758 (N_12758,N_11001,N_11227);
nand U12759 (N_12759,N_11838,N_11813);
and U12760 (N_12760,N_11685,N_11571);
or U12761 (N_12761,N_11563,N_11843);
xnor U12762 (N_12762,N_11291,N_11438);
or U12763 (N_12763,N_11787,N_11214);
nor U12764 (N_12764,N_11487,N_11660);
nand U12765 (N_12765,N_11251,N_11171);
and U12766 (N_12766,N_11169,N_11547);
nand U12767 (N_12767,N_11753,N_11090);
nand U12768 (N_12768,N_11580,N_11513);
xnor U12769 (N_12769,N_11098,N_11442);
and U12770 (N_12770,N_11393,N_11005);
xnor U12771 (N_12771,N_11811,N_11699);
xnor U12772 (N_12772,N_11157,N_11204);
nor U12773 (N_12773,N_11626,N_11174);
xnor U12774 (N_12774,N_11796,N_11670);
or U12775 (N_12775,N_11489,N_11393);
or U12776 (N_12776,N_11524,N_11580);
nor U12777 (N_12777,N_11540,N_11429);
nor U12778 (N_12778,N_11288,N_11000);
and U12779 (N_12779,N_11214,N_11626);
xor U12780 (N_12780,N_11767,N_11046);
and U12781 (N_12781,N_11884,N_11515);
or U12782 (N_12782,N_11733,N_11087);
nor U12783 (N_12783,N_11746,N_11025);
nand U12784 (N_12784,N_11271,N_11768);
nand U12785 (N_12785,N_11286,N_11399);
nor U12786 (N_12786,N_11086,N_11881);
nand U12787 (N_12787,N_11242,N_11942);
and U12788 (N_12788,N_11456,N_11219);
and U12789 (N_12789,N_11144,N_11157);
xnor U12790 (N_12790,N_11896,N_11588);
xor U12791 (N_12791,N_11185,N_11264);
and U12792 (N_12792,N_11231,N_11374);
nand U12793 (N_12793,N_11586,N_11858);
nor U12794 (N_12794,N_11531,N_11314);
or U12795 (N_12795,N_11620,N_11059);
nand U12796 (N_12796,N_11843,N_11562);
and U12797 (N_12797,N_11556,N_11637);
and U12798 (N_12798,N_11554,N_11363);
nor U12799 (N_12799,N_11170,N_11934);
nand U12800 (N_12800,N_11028,N_11306);
nand U12801 (N_12801,N_11927,N_11993);
and U12802 (N_12802,N_11374,N_11446);
or U12803 (N_12803,N_11252,N_11360);
nand U12804 (N_12804,N_11573,N_11423);
nand U12805 (N_12805,N_11317,N_11575);
and U12806 (N_12806,N_11918,N_11086);
and U12807 (N_12807,N_11778,N_11457);
nand U12808 (N_12808,N_11581,N_11546);
nor U12809 (N_12809,N_11673,N_11007);
nand U12810 (N_12810,N_11761,N_11366);
and U12811 (N_12811,N_11957,N_11511);
or U12812 (N_12812,N_11642,N_11088);
and U12813 (N_12813,N_11581,N_11215);
nand U12814 (N_12814,N_11747,N_11375);
nand U12815 (N_12815,N_11562,N_11769);
nand U12816 (N_12816,N_11783,N_11888);
nor U12817 (N_12817,N_11924,N_11749);
xor U12818 (N_12818,N_11229,N_11416);
nand U12819 (N_12819,N_11268,N_11498);
and U12820 (N_12820,N_11779,N_11299);
and U12821 (N_12821,N_11791,N_11913);
nand U12822 (N_12822,N_11381,N_11395);
xnor U12823 (N_12823,N_11340,N_11333);
nand U12824 (N_12824,N_11203,N_11508);
or U12825 (N_12825,N_11507,N_11300);
nand U12826 (N_12826,N_11277,N_11263);
nand U12827 (N_12827,N_11443,N_11840);
nor U12828 (N_12828,N_11193,N_11343);
nand U12829 (N_12829,N_11265,N_11460);
nor U12830 (N_12830,N_11201,N_11709);
nor U12831 (N_12831,N_11550,N_11469);
or U12832 (N_12832,N_11064,N_11592);
nand U12833 (N_12833,N_11393,N_11743);
or U12834 (N_12834,N_11140,N_11114);
nand U12835 (N_12835,N_11374,N_11654);
xnor U12836 (N_12836,N_11634,N_11276);
nand U12837 (N_12837,N_11950,N_11797);
nor U12838 (N_12838,N_11123,N_11862);
or U12839 (N_12839,N_11931,N_11313);
nor U12840 (N_12840,N_11165,N_11836);
xnor U12841 (N_12841,N_11564,N_11658);
and U12842 (N_12842,N_11873,N_11188);
nand U12843 (N_12843,N_11037,N_11328);
and U12844 (N_12844,N_11815,N_11717);
xnor U12845 (N_12845,N_11079,N_11242);
nor U12846 (N_12846,N_11475,N_11698);
nor U12847 (N_12847,N_11971,N_11625);
and U12848 (N_12848,N_11448,N_11368);
or U12849 (N_12849,N_11764,N_11464);
xnor U12850 (N_12850,N_11267,N_11394);
or U12851 (N_12851,N_11004,N_11221);
xor U12852 (N_12852,N_11297,N_11057);
or U12853 (N_12853,N_11012,N_11647);
nor U12854 (N_12854,N_11427,N_11467);
and U12855 (N_12855,N_11502,N_11097);
or U12856 (N_12856,N_11786,N_11473);
xor U12857 (N_12857,N_11033,N_11905);
xor U12858 (N_12858,N_11787,N_11042);
nor U12859 (N_12859,N_11625,N_11153);
and U12860 (N_12860,N_11612,N_11013);
or U12861 (N_12861,N_11405,N_11377);
nand U12862 (N_12862,N_11894,N_11929);
nor U12863 (N_12863,N_11320,N_11865);
or U12864 (N_12864,N_11691,N_11315);
or U12865 (N_12865,N_11337,N_11161);
and U12866 (N_12866,N_11574,N_11360);
xnor U12867 (N_12867,N_11574,N_11706);
nor U12868 (N_12868,N_11513,N_11164);
and U12869 (N_12869,N_11613,N_11957);
or U12870 (N_12870,N_11897,N_11400);
or U12871 (N_12871,N_11112,N_11626);
nand U12872 (N_12872,N_11978,N_11727);
nand U12873 (N_12873,N_11941,N_11841);
xnor U12874 (N_12874,N_11770,N_11098);
nor U12875 (N_12875,N_11342,N_11588);
or U12876 (N_12876,N_11493,N_11709);
nor U12877 (N_12877,N_11349,N_11253);
xor U12878 (N_12878,N_11760,N_11524);
nor U12879 (N_12879,N_11618,N_11448);
and U12880 (N_12880,N_11304,N_11941);
and U12881 (N_12881,N_11134,N_11779);
or U12882 (N_12882,N_11690,N_11152);
nand U12883 (N_12883,N_11025,N_11319);
xor U12884 (N_12884,N_11229,N_11663);
and U12885 (N_12885,N_11553,N_11773);
nand U12886 (N_12886,N_11561,N_11286);
xor U12887 (N_12887,N_11772,N_11014);
and U12888 (N_12888,N_11430,N_11138);
xnor U12889 (N_12889,N_11519,N_11469);
nor U12890 (N_12890,N_11411,N_11948);
nor U12891 (N_12891,N_11448,N_11561);
nand U12892 (N_12892,N_11765,N_11175);
nor U12893 (N_12893,N_11193,N_11421);
and U12894 (N_12894,N_11580,N_11648);
xor U12895 (N_12895,N_11144,N_11748);
xnor U12896 (N_12896,N_11276,N_11612);
nor U12897 (N_12897,N_11361,N_11380);
xor U12898 (N_12898,N_11835,N_11389);
xnor U12899 (N_12899,N_11184,N_11511);
nor U12900 (N_12900,N_11833,N_11164);
nand U12901 (N_12901,N_11931,N_11417);
and U12902 (N_12902,N_11486,N_11922);
nor U12903 (N_12903,N_11939,N_11169);
or U12904 (N_12904,N_11343,N_11294);
xor U12905 (N_12905,N_11310,N_11296);
nand U12906 (N_12906,N_11539,N_11188);
xor U12907 (N_12907,N_11166,N_11342);
and U12908 (N_12908,N_11476,N_11349);
nand U12909 (N_12909,N_11867,N_11182);
or U12910 (N_12910,N_11688,N_11100);
and U12911 (N_12911,N_11331,N_11209);
nand U12912 (N_12912,N_11982,N_11637);
and U12913 (N_12913,N_11653,N_11386);
nor U12914 (N_12914,N_11210,N_11605);
and U12915 (N_12915,N_11848,N_11076);
xnor U12916 (N_12916,N_11988,N_11050);
nand U12917 (N_12917,N_11023,N_11183);
or U12918 (N_12918,N_11916,N_11194);
xor U12919 (N_12919,N_11935,N_11800);
nand U12920 (N_12920,N_11612,N_11625);
nor U12921 (N_12921,N_11917,N_11643);
nand U12922 (N_12922,N_11029,N_11816);
nor U12923 (N_12923,N_11105,N_11288);
nor U12924 (N_12924,N_11537,N_11535);
and U12925 (N_12925,N_11398,N_11406);
nor U12926 (N_12926,N_11841,N_11704);
or U12927 (N_12927,N_11489,N_11144);
or U12928 (N_12928,N_11560,N_11818);
and U12929 (N_12929,N_11017,N_11740);
nor U12930 (N_12930,N_11388,N_11424);
xnor U12931 (N_12931,N_11096,N_11251);
and U12932 (N_12932,N_11372,N_11851);
nor U12933 (N_12933,N_11120,N_11520);
or U12934 (N_12934,N_11281,N_11581);
nand U12935 (N_12935,N_11017,N_11682);
xnor U12936 (N_12936,N_11697,N_11371);
xor U12937 (N_12937,N_11412,N_11187);
nand U12938 (N_12938,N_11756,N_11918);
nand U12939 (N_12939,N_11727,N_11234);
xor U12940 (N_12940,N_11532,N_11371);
and U12941 (N_12941,N_11610,N_11350);
xnor U12942 (N_12942,N_11185,N_11459);
and U12943 (N_12943,N_11054,N_11899);
nor U12944 (N_12944,N_11253,N_11639);
xor U12945 (N_12945,N_11210,N_11275);
nor U12946 (N_12946,N_11231,N_11753);
nor U12947 (N_12947,N_11051,N_11472);
nand U12948 (N_12948,N_11457,N_11891);
xor U12949 (N_12949,N_11121,N_11583);
nand U12950 (N_12950,N_11561,N_11184);
and U12951 (N_12951,N_11033,N_11000);
or U12952 (N_12952,N_11843,N_11707);
or U12953 (N_12953,N_11931,N_11594);
or U12954 (N_12954,N_11756,N_11220);
and U12955 (N_12955,N_11245,N_11327);
nor U12956 (N_12956,N_11980,N_11160);
and U12957 (N_12957,N_11165,N_11473);
nand U12958 (N_12958,N_11336,N_11210);
nor U12959 (N_12959,N_11654,N_11799);
and U12960 (N_12960,N_11225,N_11788);
or U12961 (N_12961,N_11792,N_11776);
and U12962 (N_12962,N_11642,N_11895);
and U12963 (N_12963,N_11017,N_11300);
or U12964 (N_12964,N_11584,N_11566);
nor U12965 (N_12965,N_11326,N_11885);
nor U12966 (N_12966,N_11627,N_11489);
or U12967 (N_12967,N_11035,N_11405);
nor U12968 (N_12968,N_11099,N_11867);
and U12969 (N_12969,N_11718,N_11719);
nor U12970 (N_12970,N_11055,N_11321);
nand U12971 (N_12971,N_11527,N_11054);
and U12972 (N_12972,N_11213,N_11973);
nand U12973 (N_12973,N_11570,N_11028);
or U12974 (N_12974,N_11651,N_11193);
nor U12975 (N_12975,N_11880,N_11612);
or U12976 (N_12976,N_11478,N_11223);
and U12977 (N_12977,N_11936,N_11828);
or U12978 (N_12978,N_11562,N_11857);
or U12979 (N_12979,N_11893,N_11989);
or U12980 (N_12980,N_11842,N_11667);
xor U12981 (N_12981,N_11105,N_11535);
nand U12982 (N_12982,N_11666,N_11611);
nor U12983 (N_12983,N_11575,N_11247);
nand U12984 (N_12984,N_11245,N_11059);
xor U12985 (N_12985,N_11453,N_11636);
nor U12986 (N_12986,N_11597,N_11767);
nor U12987 (N_12987,N_11723,N_11873);
or U12988 (N_12988,N_11599,N_11925);
and U12989 (N_12989,N_11623,N_11913);
nand U12990 (N_12990,N_11284,N_11724);
nor U12991 (N_12991,N_11750,N_11793);
nor U12992 (N_12992,N_11798,N_11276);
or U12993 (N_12993,N_11731,N_11760);
and U12994 (N_12994,N_11029,N_11763);
or U12995 (N_12995,N_11549,N_11841);
nand U12996 (N_12996,N_11093,N_11579);
and U12997 (N_12997,N_11400,N_11670);
nand U12998 (N_12998,N_11230,N_11795);
and U12999 (N_12999,N_11280,N_11117);
and U13000 (N_13000,N_12979,N_12941);
nand U13001 (N_13001,N_12609,N_12408);
and U13002 (N_13002,N_12395,N_12095);
xor U13003 (N_13003,N_12694,N_12615);
or U13004 (N_13004,N_12624,N_12810);
xnor U13005 (N_13005,N_12799,N_12210);
and U13006 (N_13006,N_12018,N_12113);
and U13007 (N_13007,N_12480,N_12500);
nor U13008 (N_13008,N_12312,N_12604);
nand U13009 (N_13009,N_12372,N_12432);
or U13010 (N_13010,N_12848,N_12525);
xnor U13011 (N_13011,N_12171,N_12011);
xor U13012 (N_13012,N_12722,N_12928);
or U13013 (N_13013,N_12476,N_12428);
xor U13014 (N_13014,N_12429,N_12735);
and U13015 (N_13015,N_12055,N_12237);
and U13016 (N_13016,N_12073,N_12310);
nand U13017 (N_13017,N_12339,N_12990);
and U13018 (N_13018,N_12384,N_12587);
and U13019 (N_13019,N_12635,N_12797);
nand U13020 (N_13020,N_12398,N_12571);
nand U13021 (N_13021,N_12366,N_12352);
or U13022 (N_13022,N_12707,N_12324);
or U13023 (N_13023,N_12281,N_12047);
nand U13024 (N_13024,N_12924,N_12071);
xnor U13025 (N_13025,N_12056,N_12637);
nand U13026 (N_13026,N_12871,N_12331);
nor U13027 (N_13027,N_12667,N_12961);
and U13028 (N_13028,N_12917,N_12894);
and U13029 (N_13029,N_12440,N_12484);
and U13030 (N_13030,N_12962,N_12856);
or U13031 (N_13031,N_12613,N_12463);
or U13032 (N_13032,N_12666,N_12948);
nand U13033 (N_13033,N_12037,N_12016);
xnor U13034 (N_13034,N_12329,N_12744);
xor U13035 (N_13035,N_12473,N_12247);
nand U13036 (N_13036,N_12345,N_12414);
and U13037 (N_13037,N_12616,N_12994);
nor U13038 (N_13038,N_12387,N_12751);
and U13039 (N_13039,N_12173,N_12892);
and U13040 (N_13040,N_12779,N_12364);
xnor U13041 (N_13041,N_12176,N_12721);
nand U13042 (N_13042,N_12365,N_12021);
and U13043 (N_13043,N_12253,N_12864);
xnor U13044 (N_13044,N_12711,N_12900);
or U13045 (N_13045,N_12193,N_12317);
xor U13046 (N_13046,N_12868,N_12040);
or U13047 (N_13047,N_12293,N_12791);
nor U13048 (N_13048,N_12377,N_12517);
xnor U13049 (N_13049,N_12893,N_12318);
or U13050 (N_13050,N_12456,N_12148);
or U13051 (N_13051,N_12001,N_12241);
or U13052 (N_13052,N_12921,N_12708);
nand U13053 (N_13053,N_12438,N_12570);
and U13054 (N_13054,N_12728,N_12454);
nand U13055 (N_13055,N_12922,N_12147);
or U13056 (N_13056,N_12959,N_12514);
xor U13057 (N_13057,N_12131,N_12788);
and U13058 (N_13058,N_12025,N_12431);
and U13059 (N_13059,N_12772,N_12907);
nand U13060 (N_13060,N_12986,N_12160);
and U13061 (N_13061,N_12705,N_12211);
xor U13062 (N_13062,N_12134,N_12421);
xnor U13063 (N_13063,N_12305,N_12044);
xor U13064 (N_13064,N_12939,N_12695);
or U13065 (N_13065,N_12209,N_12789);
or U13066 (N_13066,N_12337,N_12261);
nor U13067 (N_13067,N_12409,N_12181);
and U13068 (N_13068,N_12611,N_12837);
or U13069 (N_13069,N_12862,N_12307);
or U13070 (N_13070,N_12822,N_12684);
nor U13071 (N_13071,N_12970,N_12085);
nor U13072 (N_13072,N_12869,N_12692);
nand U13073 (N_13073,N_12703,N_12243);
nand U13074 (N_13074,N_12698,N_12851);
or U13075 (N_13075,N_12487,N_12841);
and U13076 (N_13076,N_12760,N_12642);
nand U13077 (N_13077,N_12075,N_12726);
nand U13078 (N_13078,N_12010,N_12522);
xnor U13079 (N_13079,N_12644,N_12424);
xnor U13080 (N_13080,N_12200,N_12993);
and U13081 (N_13081,N_12397,N_12375);
xnor U13082 (N_13082,N_12966,N_12688);
nand U13083 (N_13083,N_12027,N_12087);
xor U13084 (N_13084,N_12320,N_12518);
and U13085 (N_13085,N_12739,N_12566);
and U13086 (N_13086,N_12043,N_12254);
nor U13087 (N_13087,N_12787,N_12098);
or U13088 (N_13088,N_12081,N_12283);
or U13089 (N_13089,N_12065,N_12296);
nor U13090 (N_13090,N_12887,N_12236);
xnor U13091 (N_13091,N_12673,N_12733);
nand U13092 (N_13092,N_12466,N_12139);
nor U13093 (N_13093,N_12468,N_12945);
or U13094 (N_13094,N_12763,N_12671);
nor U13095 (N_13095,N_12836,N_12441);
xnor U13096 (N_13096,N_12141,N_12094);
xnor U13097 (N_13097,N_12538,N_12641);
and U13098 (N_13098,N_12839,N_12942);
or U13099 (N_13099,N_12104,N_12342);
nand U13100 (N_13100,N_12818,N_12082);
nor U13101 (N_13101,N_12042,N_12031);
and U13102 (N_13102,N_12294,N_12453);
nor U13103 (N_13103,N_12062,N_12649);
nand U13104 (N_13104,N_12861,N_12008);
and U13105 (N_13105,N_12954,N_12239);
and U13106 (N_13106,N_12656,N_12479);
and U13107 (N_13107,N_12413,N_12101);
or U13108 (N_13108,N_12060,N_12731);
xor U13109 (N_13109,N_12632,N_12497);
nor U13110 (N_13110,N_12164,N_12678);
and U13111 (N_13111,N_12547,N_12277);
or U13112 (N_13112,N_12334,N_12447);
and U13113 (N_13113,N_12314,N_12817);
xnor U13114 (N_13114,N_12880,N_12890);
nor U13115 (N_13115,N_12508,N_12588);
and U13116 (N_13116,N_12813,N_12423);
nor U13117 (N_13117,N_12149,N_12410);
nor U13118 (N_13118,N_12156,N_12406);
or U13119 (N_13119,N_12560,N_12316);
xor U13120 (N_13120,N_12114,N_12255);
nor U13121 (N_13121,N_12765,N_12713);
nor U13122 (N_13122,N_12309,N_12912);
nor U13123 (N_13123,N_12589,N_12984);
nor U13124 (N_13124,N_12079,N_12761);
and U13125 (N_13125,N_12555,N_12106);
nand U13126 (N_13126,N_12554,N_12226);
nor U13127 (N_13127,N_12842,N_12449);
nand U13128 (N_13128,N_12205,N_12600);
nor U13129 (N_13129,N_12038,N_12299);
or U13130 (N_13130,N_12544,N_12991);
and U13131 (N_13131,N_12415,N_12778);
nor U13132 (N_13132,N_12605,N_12121);
nand U13133 (N_13133,N_12552,N_12284);
nor U13134 (N_13134,N_12373,N_12458);
xor U13135 (N_13135,N_12483,N_12883);
nor U13136 (N_13136,N_12157,N_12475);
nand U13137 (N_13137,N_12831,N_12670);
xor U13138 (N_13138,N_12578,N_12385);
nand U13139 (N_13139,N_12242,N_12512);
nor U13140 (N_13140,N_12800,N_12825);
or U13141 (N_13141,N_12950,N_12911);
xor U13142 (N_13142,N_12072,N_12807);
and U13143 (N_13143,N_12776,N_12145);
or U13144 (N_13144,N_12658,N_12865);
nor U13145 (N_13145,N_12461,N_12919);
and U13146 (N_13146,N_12889,N_12235);
or U13147 (N_13147,N_12981,N_12505);
nand U13148 (N_13148,N_12834,N_12103);
and U13149 (N_13149,N_12492,N_12433);
or U13150 (N_13150,N_12380,N_12257);
nand U13151 (N_13151,N_12361,N_12151);
nand U13152 (N_13152,N_12940,N_12606);
and U13153 (N_13153,N_12457,N_12786);
or U13154 (N_13154,N_12402,N_12964);
or U13155 (N_13155,N_12266,N_12186);
and U13156 (N_13156,N_12576,N_12974);
nand U13157 (N_13157,N_12099,N_12541);
or U13158 (N_13158,N_12353,N_12022);
and U13159 (N_13159,N_12654,N_12163);
nor U13160 (N_13160,N_12832,N_12549);
xnor U13161 (N_13161,N_12798,N_12218);
nor U13162 (N_13162,N_12740,N_12960);
or U13163 (N_13163,N_12059,N_12464);
xnor U13164 (N_13164,N_12017,N_12596);
or U13165 (N_13165,N_12973,N_12404);
nor U13166 (N_13166,N_12371,N_12773);
and U13167 (N_13167,N_12762,N_12363);
nand U13168 (N_13168,N_12450,N_12640);
and U13169 (N_13169,N_12203,N_12199);
and U13170 (N_13170,N_12680,N_12197);
xnor U13171 (N_13171,N_12348,N_12448);
nand U13172 (N_13172,N_12853,N_12282);
or U13173 (N_13173,N_12125,N_12625);
nor U13174 (N_13174,N_12982,N_12399);
nor U13175 (N_13175,N_12225,N_12191);
nand U13176 (N_13176,N_12224,N_12873);
or U13177 (N_13177,N_12565,N_12679);
or U13178 (N_13178,N_12699,N_12881);
nor U13179 (N_13179,N_12485,N_12168);
nor U13180 (N_13180,N_12933,N_12947);
and U13181 (N_13181,N_12574,N_12367);
nand U13182 (N_13182,N_12368,N_12080);
nand U13183 (N_13183,N_12411,N_12621);
nand U13184 (N_13184,N_12929,N_12128);
nand U13185 (N_13185,N_12231,N_12478);
or U13186 (N_13186,N_12488,N_12581);
xor U13187 (N_13187,N_12845,N_12407);
nor U13188 (N_13188,N_12298,N_12550);
nand U13189 (N_13189,N_12091,N_12774);
xnor U13190 (N_13190,N_12290,N_12758);
and U13191 (N_13191,N_12591,N_12516);
nor U13192 (N_13192,N_12327,N_12129);
nor U13193 (N_13193,N_12801,N_12906);
or U13194 (N_13194,N_12166,N_12957);
and U13195 (N_13195,N_12819,N_12246);
or U13196 (N_13196,N_12196,N_12418);
nor U13197 (N_13197,N_12304,N_12455);
or U13198 (N_13198,N_12972,N_12738);
nand U13199 (N_13199,N_12852,N_12035);
nor U13200 (N_13200,N_12556,N_12741);
nor U13201 (N_13201,N_12401,N_12378);
and U13202 (N_13202,N_12002,N_12201);
or U13203 (N_13203,N_12746,N_12700);
xor U13204 (N_13204,N_12150,N_12288);
nor U13205 (N_13205,N_12169,N_12771);
nand U13206 (N_13206,N_12102,N_12618);
and U13207 (N_13207,N_12383,N_12357);
or U13208 (N_13208,N_12221,N_12612);
xnor U13209 (N_13209,N_12360,N_12041);
xnor U13210 (N_13210,N_12736,N_12144);
or U13211 (N_13211,N_12351,N_12162);
nor U13212 (N_13212,N_12195,N_12474);
xor U13213 (N_13213,N_12730,N_12926);
and U13214 (N_13214,N_12527,N_12105);
xor U13215 (N_13215,N_12058,N_12523);
nand U13216 (N_13216,N_12562,N_12628);
nor U13217 (N_13217,N_12061,N_12084);
or U13218 (N_13218,N_12215,N_12267);
and U13219 (N_13219,N_12491,N_12559);
or U13220 (N_13220,N_12392,N_12070);
and U13221 (N_13221,N_12586,N_12054);
nor U13222 (N_13222,N_12835,N_12108);
nor U13223 (N_13223,N_12036,N_12498);
xor U13224 (N_13224,N_12117,N_12083);
or U13225 (N_13225,N_12668,N_12119);
nand U13226 (N_13226,N_12875,N_12952);
nor U13227 (N_13227,N_12369,N_12706);
xnor U13228 (N_13228,N_12968,N_12391);
nand U13229 (N_13229,N_12719,N_12386);
nand U13230 (N_13230,N_12750,N_12734);
xor U13231 (N_13231,N_12451,N_12965);
nor U13232 (N_13232,N_12285,N_12066);
and U13233 (N_13233,N_12426,N_12340);
or U13234 (N_13234,N_12422,N_12886);
xor U13235 (N_13235,N_12443,N_12459);
nor U13236 (N_13236,N_12536,N_12526);
nand U13237 (N_13237,N_12127,N_12009);
xor U13238 (N_13238,N_12471,N_12617);
or U13239 (N_13239,N_12557,N_12821);
nor U13240 (N_13240,N_12638,N_12100);
nand U13241 (N_13241,N_12724,N_12495);
and U13242 (N_13242,N_12400,N_12003);
xor U13243 (N_13243,N_12276,N_12252);
nand U13244 (N_13244,N_12382,N_12077);
or U13245 (N_13245,N_12158,N_12244);
nor U13246 (N_13246,N_12292,N_12093);
xnor U13247 (N_13247,N_12826,N_12086);
and U13248 (N_13248,N_12496,N_12208);
and U13249 (N_13249,N_12785,N_12165);
nor U13250 (N_13250,N_12696,N_12969);
nand U13251 (N_13251,N_12756,N_12109);
xor U13252 (N_13252,N_12238,N_12659);
xnor U13253 (N_13253,N_12946,N_12812);
nand U13254 (N_13254,N_12133,N_12472);
xor U13255 (N_13255,N_12573,N_12506);
nand U13256 (N_13256,N_12828,N_12511);
and U13257 (N_13257,N_12301,N_12716);
and U13258 (N_13258,N_12805,N_12202);
xnor U13259 (N_13259,N_12824,N_12806);
or U13260 (N_13260,N_12569,N_12877);
xnor U13261 (N_13261,N_12983,N_12938);
and U13262 (N_13262,N_12174,N_12546);
nand U13263 (N_13263,N_12216,N_12178);
and U13264 (N_13264,N_12913,N_12350);
nor U13265 (N_13265,N_12590,N_12850);
and U13266 (N_13266,N_12660,N_12614);
nand U13267 (N_13267,N_12888,N_12452);
or U13268 (N_13268,N_12985,N_12325);
or U13269 (N_13269,N_12521,N_12995);
xnor U13270 (N_13270,N_12602,N_12814);
nor U13271 (N_13271,N_12295,N_12980);
nor U13272 (N_13272,N_12030,N_12359);
or U13273 (N_13273,N_12619,N_12006);
xor U13274 (N_13274,N_12757,N_12580);
xor U13275 (N_13275,N_12494,N_12122);
or U13276 (N_13276,N_12855,N_12405);
nor U13277 (N_13277,N_12015,N_12185);
nand U13278 (N_13278,N_12172,N_12394);
nor U13279 (N_13279,N_12245,N_12034);
xor U13280 (N_13280,N_12647,N_12194);
xnor U13281 (N_13281,N_12096,N_12112);
nand U13282 (N_13282,N_12650,N_12182);
xnor U13283 (N_13283,N_12575,N_12437);
xnor U13284 (N_13284,N_12228,N_12553);
nand U13285 (N_13285,N_12572,N_12847);
nand U13286 (N_13286,N_12795,N_12998);
and U13287 (N_13287,N_12748,N_12233);
nand U13288 (N_13288,N_12681,N_12430);
xnor U13289 (N_13289,N_12265,N_12090);
nand U13290 (N_13290,N_12901,N_12727);
or U13291 (N_13291,N_12783,N_12362);
nor U13292 (N_13292,N_12997,N_12420);
nor U13293 (N_13293,N_12446,N_12223);
nand U13294 (N_13294,N_12709,N_12212);
nand U13295 (N_13295,N_12005,N_12833);
xor U13296 (N_13296,N_12214,N_12291);
nor U13297 (N_13297,N_12780,N_12050);
or U13298 (N_13298,N_12271,N_12766);
nor U13299 (N_13299,N_12802,N_12608);
xor U13300 (N_13300,N_12934,N_12840);
and U13301 (N_13301,N_12250,N_12794);
nand U13302 (N_13302,N_12460,N_12045);
xnor U13303 (N_13303,N_12545,N_12595);
and U13304 (N_13304,N_12768,N_12672);
nand U13305 (N_13305,N_12273,N_12412);
and U13306 (N_13306,N_12583,N_12425);
and U13307 (N_13307,N_12051,N_12558);
or U13308 (N_13308,N_12923,N_12515);
nand U13309 (N_13309,N_12676,N_12823);
nand U13310 (N_13310,N_12607,N_12280);
or U13311 (N_13311,N_12623,N_12319);
nor U13312 (N_13312,N_12770,N_12490);
xor U13313 (N_13313,N_12229,N_12704);
nand U13314 (N_13314,N_12445,N_12076);
xnor U13315 (N_13315,N_12723,N_12020);
or U13316 (N_13316,N_12662,N_12519);
xor U13317 (N_13317,N_12916,N_12978);
nor U13318 (N_13318,N_12355,N_12220);
and U13319 (N_13319,N_12146,N_12338);
nand U13320 (N_13320,N_12563,N_12321);
and U13321 (N_13321,N_12349,N_12665);
nor U13322 (N_13322,N_12192,N_12326);
xnor U13323 (N_13323,N_12315,N_12669);
xnor U13324 (N_13324,N_12715,N_12636);
and U13325 (N_13325,N_12657,N_12531);
nand U13326 (N_13326,N_12393,N_12743);
xnor U13327 (N_13327,N_12198,N_12300);
xor U13328 (N_13328,N_12249,N_12720);
nor U13329 (N_13329,N_12564,N_12026);
nand U13330 (N_13330,N_12567,N_12753);
and U13331 (N_13331,N_12701,N_12918);
and U13332 (N_13332,N_12520,N_12535);
nor U13333 (N_13333,N_12092,N_12956);
and U13334 (N_13334,N_12126,N_12804);
nand U13335 (N_13335,N_12328,N_12863);
nor U13336 (N_13336,N_12811,N_12534);
or U13337 (N_13337,N_12661,N_12330);
and U13338 (N_13338,N_12937,N_12436);
or U13339 (N_13339,N_12504,N_12486);
or U13340 (N_13340,N_12416,N_12908);
nand U13341 (N_13341,N_12876,N_12502);
nand U13342 (N_13342,N_12975,N_12376);
and U13343 (N_13343,N_12270,N_12333);
xor U13344 (N_13344,N_12130,N_12381);
nor U13345 (N_13345,N_12354,N_12389);
or U13346 (N_13346,N_12467,N_12815);
nand U13347 (N_13347,N_12944,N_12039);
xnor U13348 (N_13348,N_12529,N_12159);
nand U13349 (N_13349,N_12603,N_12167);
and U13350 (N_13350,N_12138,N_12878);
nand U13351 (N_13351,N_12909,N_12259);
nand U13352 (N_13352,N_12227,N_12336);
and U13353 (N_13353,N_12882,N_12434);
or U13354 (N_13354,N_12925,N_12577);
nor U13355 (N_13355,N_12183,N_12594);
or U13356 (N_13356,N_12513,N_12207);
nor U13357 (N_13357,N_12442,N_12630);
xnor U13358 (N_13358,N_12601,N_12999);
xnor U13359 (N_13359,N_12470,N_12691);
nand U13360 (N_13360,N_12803,N_12417);
xor U13361 (N_13361,N_12593,N_12097);
xnor U13362 (N_13362,N_12530,N_12914);
nand U13363 (N_13363,N_12439,N_12289);
nor U13364 (N_13364,N_12052,N_12714);
and U13365 (N_13365,N_12809,N_12078);
nor U13366 (N_13366,N_12633,N_12874);
xor U13367 (N_13367,N_12343,N_12967);
nand U13368 (N_13368,N_12932,N_12648);
xor U13369 (N_13369,N_12626,N_12915);
and U13370 (N_13370,N_12256,N_12689);
xnor U13371 (N_13371,N_12248,N_12346);
and U13372 (N_13372,N_12507,N_12493);
nor U13373 (N_13373,N_12275,N_12322);
and U13374 (N_13374,N_12793,N_12528);
xnor U13375 (N_13375,N_12896,N_12177);
nand U13376 (N_13376,N_12987,N_12323);
nand U13377 (N_13377,N_12663,N_12068);
or U13378 (N_13378,N_12949,N_12028);
nand U13379 (N_13379,N_12717,N_12769);
nand U13380 (N_13380,N_12548,N_12465);
and U13381 (N_13381,N_12118,N_12755);
xor U13382 (N_13382,N_12189,N_12023);
nand U13383 (N_13383,N_12920,N_12585);
nor U13384 (N_13384,N_12781,N_12561);
nand U13385 (N_13385,N_12069,N_12057);
or U13386 (N_13386,N_12955,N_12370);
or U13387 (N_13387,N_12885,N_12143);
nand U13388 (N_13388,N_12686,N_12115);
or U13389 (N_13389,N_12796,N_12462);
xor U13390 (N_13390,N_12963,N_12792);
nand U13391 (N_13391,N_12857,N_12046);
and U13392 (N_13392,N_12014,N_12971);
or U13393 (N_13393,N_12808,N_12844);
xor U13394 (N_13394,N_12142,N_12132);
xor U13395 (N_13395,N_12992,N_12693);
nand U13396 (N_13396,N_12219,N_12931);
xor U13397 (N_13397,N_12286,N_12866);
xnor U13398 (N_13398,N_12652,N_12107);
and U13399 (N_13399,N_12674,N_12390);
nor U13400 (N_13400,N_12419,N_12899);
or U13401 (N_13401,N_12599,N_12444);
nor U13402 (N_13402,N_12867,N_12745);
xnor U13403 (N_13403,N_12677,N_12532);
or U13404 (N_13404,N_12136,N_12024);
and U13405 (N_13405,N_12388,N_12204);
nor U13406 (N_13406,N_12631,N_12435);
nor U13407 (N_13407,N_12622,N_12344);
nand U13408 (N_13408,N_12120,N_12905);
and U13409 (N_13409,N_12777,N_12958);
xnor U13410 (N_13410,N_12664,N_12634);
nand U13411 (N_13411,N_12152,N_12332);
and U13412 (N_13412,N_12568,N_12188);
or U13413 (N_13413,N_12651,N_12579);
nand U13414 (N_13414,N_12379,N_12891);
or U13415 (N_13415,N_12499,N_12903);
nor U13416 (N_13416,N_12213,N_12175);
and U13417 (N_13417,N_12927,N_12935);
nor U13418 (N_13418,N_12048,N_12222);
or U13419 (N_13419,N_12161,N_12627);
and U13420 (N_13420,N_12049,N_12187);
and U13421 (N_13421,N_12272,N_12645);
and U13422 (N_13422,N_12584,N_12258);
nor U13423 (N_13423,N_12358,N_12764);
nand U13424 (N_13424,N_12019,N_12610);
and U13425 (N_13425,N_12629,N_12240);
nor U13426 (N_13426,N_12729,N_12895);
and U13427 (N_13427,N_12543,N_12598);
or U13428 (N_13428,N_12217,N_12064);
nor U13429 (N_13429,N_12951,N_12790);
xnor U13430 (N_13430,N_12302,N_12074);
xnor U13431 (N_13431,N_12509,N_12004);
xnor U13432 (N_13432,N_12816,N_12718);
or U13433 (N_13433,N_12737,N_12341);
xnor U13434 (N_13434,N_12190,N_12697);
xnor U13435 (N_13435,N_12110,N_12013);
and U13436 (N_13436,N_12303,N_12347);
and U13437 (N_13437,N_12170,N_12481);
nand U13438 (N_13438,N_12859,N_12725);
nor U13439 (N_13439,N_12264,N_12989);
nor U13440 (N_13440,N_12124,N_12858);
or U13441 (N_13441,N_12592,N_12653);
nor U13442 (N_13442,N_12269,N_12469);
xnor U13443 (N_13443,N_12687,N_12838);
or U13444 (N_13444,N_12830,N_12732);
nand U13445 (N_13445,N_12311,N_12710);
nor U13446 (N_13446,N_12137,N_12278);
and U13447 (N_13447,N_12033,N_12232);
and U13448 (N_13448,N_12053,N_12335);
nor U13449 (N_13449,N_12533,N_12872);
xnor U13450 (N_13450,N_12029,N_12287);
and U13451 (N_13451,N_12184,N_12306);
or U13452 (N_13452,N_12690,N_12775);
or U13453 (N_13453,N_12374,N_12988);
and U13454 (N_13454,N_12260,N_12489);
nand U13455 (N_13455,N_12943,N_12234);
and U13456 (N_13456,N_12759,N_12089);
or U13457 (N_13457,N_12827,N_12682);
xnor U13458 (N_13458,N_12297,N_12620);
nand U13459 (N_13459,N_12206,N_12860);
or U13460 (N_13460,N_12884,N_12313);
nand U13461 (N_13461,N_12012,N_12754);
or U13462 (N_13462,N_12356,N_12902);
xnor U13463 (N_13463,N_12251,N_12179);
nand U13464 (N_13464,N_12477,N_12849);
and U13465 (N_13465,N_12140,N_12482);
nand U13466 (N_13466,N_12646,N_12843);
and U13467 (N_13467,N_12675,N_12930);
or U13468 (N_13468,N_12782,N_12274);
nand U13469 (N_13469,N_12180,N_12829);
and U13470 (N_13470,N_12032,N_12904);
nor U13471 (N_13471,N_12007,N_12154);
or U13472 (N_13472,N_12854,N_12897);
or U13473 (N_13473,N_12702,N_12501);
and U13474 (N_13474,N_12597,N_12155);
or U13475 (N_13475,N_12898,N_12116);
or U13476 (N_13476,N_12153,N_12712);
xnor U13477 (N_13477,N_12643,N_12000);
or U13478 (N_13478,N_12540,N_12551);
nor U13479 (N_13479,N_12111,N_12742);
xor U13480 (N_13480,N_12262,N_12976);
and U13481 (N_13481,N_12953,N_12279);
or U13482 (N_13482,N_12977,N_12539);
nand U13483 (N_13483,N_12996,N_12683);
xor U13484 (N_13484,N_12542,N_12767);
nor U13485 (N_13485,N_12685,N_12910);
xor U13486 (N_13486,N_12308,N_12582);
or U13487 (N_13487,N_12403,N_12268);
xor U13488 (N_13488,N_12537,N_12503);
nand U13489 (N_13489,N_12524,N_12784);
xor U13490 (N_13490,N_12135,N_12936);
nand U13491 (N_13491,N_12263,N_12870);
or U13492 (N_13492,N_12820,N_12752);
xor U13493 (N_13493,N_12123,N_12088);
nand U13494 (N_13494,N_12063,N_12396);
nand U13495 (N_13495,N_12879,N_12747);
xor U13496 (N_13496,N_12510,N_12427);
nor U13497 (N_13497,N_12749,N_12230);
nand U13498 (N_13498,N_12067,N_12639);
nand U13499 (N_13499,N_12846,N_12655);
nand U13500 (N_13500,N_12468,N_12993);
nor U13501 (N_13501,N_12792,N_12820);
or U13502 (N_13502,N_12950,N_12290);
nand U13503 (N_13503,N_12797,N_12398);
or U13504 (N_13504,N_12624,N_12502);
nor U13505 (N_13505,N_12094,N_12144);
or U13506 (N_13506,N_12507,N_12038);
or U13507 (N_13507,N_12967,N_12114);
and U13508 (N_13508,N_12684,N_12927);
or U13509 (N_13509,N_12878,N_12697);
xnor U13510 (N_13510,N_12631,N_12580);
nor U13511 (N_13511,N_12648,N_12530);
nand U13512 (N_13512,N_12381,N_12315);
or U13513 (N_13513,N_12907,N_12222);
nor U13514 (N_13514,N_12785,N_12422);
or U13515 (N_13515,N_12586,N_12611);
or U13516 (N_13516,N_12279,N_12917);
nand U13517 (N_13517,N_12566,N_12034);
nor U13518 (N_13518,N_12302,N_12511);
nand U13519 (N_13519,N_12630,N_12020);
nand U13520 (N_13520,N_12317,N_12236);
nand U13521 (N_13521,N_12975,N_12685);
nand U13522 (N_13522,N_12024,N_12160);
nor U13523 (N_13523,N_12569,N_12614);
nand U13524 (N_13524,N_12460,N_12933);
nor U13525 (N_13525,N_12423,N_12113);
nand U13526 (N_13526,N_12640,N_12695);
nand U13527 (N_13527,N_12708,N_12256);
xor U13528 (N_13528,N_12363,N_12944);
or U13529 (N_13529,N_12720,N_12479);
nand U13530 (N_13530,N_12070,N_12416);
nor U13531 (N_13531,N_12564,N_12224);
and U13532 (N_13532,N_12498,N_12888);
nand U13533 (N_13533,N_12742,N_12454);
xor U13534 (N_13534,N_12502,N_12332);
or U13535 (N_13535,N_12471,N_12322);
nor U13536 (N_13536,N_12341,N_12927);
nand U13537 (N_13537,N_12768,N_12397);
and U13538 (N_13538,N_12529,N_12850);
nand U13539 (N_13539,N_12781,N_12240);
nand U13540 (N_13540,N_12363,N_12572);
and U13541 (N_13541,N_12872,N_12081);
nor U13542 (N_13542,N_12287,N_12447);
nand U13543 (N_13543,N_12274,N_12386);
nand U13544 (N_13544,N_12823,N_12680);
and U13545 (N_13545,N_12845,N_12606);
or U13546 (N_13546,N_12046,N_12136);
nor U13547 (N_13547,N_12882,N_12498);
xor U13548 (N_13548,N_12241,N_12028);
nand U13549 (N_13549,N_12448,N_12428);
nor U13550 (N_13550,N_12866,N_12073);
nor U13551 (N_13551,N_12599,N_12224);
and U13552 (N_13552,N_12679,N_12308);
and U13553 (N_13553,N_12553,N_12663);
nor U13554 (N_13554,N_12835,N_12116);
nor U13555 (N_13555,N_12000,N_12456);
nor U13556 (N_13556,N_12959,N_12738);
or U13557 (N_13557,N_12250,N_12579);
or U13558 (N_13558,N_12583,N_12132);
or U13559 (N_13559,N_12718,N_12358);
nor U13560 (N_13560,N_12404,N_12912);
or U13561 (N_13561,N_12617,N_12318);
xor U13562 (N_13562,N_12477,N_12060);
and U13563 (N_13563,N_12257,N_12222);
or U13564 (N_13564,N_12921,N_12640);
nor U13565 (N_13565,N_12861,N_12013);
and U13566 (N_13566,N_12595,N_12908);
nand U13567 (N_13567,N_12326,N_12963);
nor U13568 (N_13568,N_12502,N_12203);
nor U13569 (N_13569,N_12936,N_12416);
or U13570 (N_13570,N_12021,N_12715);
xor U13571 (N_13571,N_12498,N_12375);
xnor U13572 (N_13572,N_12757,N_12840);
or U13573 (N_13573,N_12977,N_12728);
and U13574 (N_13574,N_12278,N_12094);
and U13575 (N_13575,N_12829,N_12167);
xnor U13576 (N_13576,N_12670,N_12402);
or U13577 (N_13577,N_12410,N_12671);
or U13578 (N_13578,N_12586,N_12827);
or U13579 (N_13579,N_12166,N_12296);
nor U13580 (N_13580,N_12327,N_12187);
nand U13581 (N_13581,N_12370,N_12703);
or U13582 (N_13582,N_12115,N_12809);
nand U13583 (N_13583,N_12210,N_12861);
nand U13584 (N_13584,N_12870,N_12055);
nand U13585 (N_13585,N_12362,N_12489);
or U13586 (N_13586,N_12474,N_12727);
xor U13587 (N_13587,N_12507,N_12101);
nor U13588 (N_13588,N_12075,N_12823);
nor U13589 (N_13589,N_12309,N_12837);
and U13590 (N_13590,N_12945,N_12026);
xor U13591 (N_13591,N_12717,N_12601);
xnor U13592 (N_13592,N_12468,N_12991);
or U13593 (N_13593,N_12187,N_12650);
xnor U13594 (N_13594,N_12863,N_12884);
nand U13595 (N_13595,N_12913,N_12844);
and U13596 (N_13596,N_12158,N_12421);
xnor U13597 (N_13597,N_12426,N_12225);
xnor U13598 (N_13598,N_12527,N_12409);
and U13599 (N_13599,N_12248,N_12595);
xnor U13600 (N_13600,N_12472,N_12018);
nand U13601 (N_13601,N_12019,N_12604);
and U13602 (N_13602,N_12899,N_12019);
nand U13603 (N_13603,N_12144,N_12253);
nand U13604 (N_13604,N_12443,N_12946);
or U13605 (N_13605,N_12940,N_12740);
nor U13606 (N_13606,N_12899,N_12190);
and U13607 (N_13607,N_12996,N_12037);
or U13608 (N_13608,N_12751,N_12307);
or U13609 (N_13609,N_12064,N_12463);
xnor U13610 (N_13610,N_12545,N_12280);
xnor U13611 (N_13611,N_12171,N_12987);
xnor U13612 (N_13612,N_12338,N_12130);
nor U13613 (N_13613,N_12133,N_12688);
or U13614 (N_13614,N_12247,N_12442);
or U13615 (N_13615,N_12152,N_12319);
or U13616 (N_13616,N_12889,N_12121);
or U13617 (N_13617,N_12194,N_12237);
nor U13618 (N_13618,N_12616,N_12333);
nor U13619 (N_13619,N_12017,N_12634);
nor U13620 (N_13620,N_12215,N_12075);
xor U13621 (N_13621,N_12338,N_12623);
or U13622 (N_13622,N_12311,N_12483);
or U13623 (N_13623,N_12887,N_12029);
or U13624 (N_13624,N_12521,N_12945);
nand U13625 (N_13625,N_12379,N_12717);
and U13626 (N_13626,N_12363,N_12859);
nor U13627 (N_13627,N_12819,N_12161);
nor U13628 (N_13628,N_12118,N_12767);
and U13629 (N_13629,N_12506,N_12023);
nor U13630 (N_13630,N_12311,N_12692);
nor U13631 (N_13631,N_12924,N_12905);
xor U13632 (N_13632,N_12489,N_12428);
and U13633 (N_13633,N_12107,N_12619);
or U13634 (N_13634,N_12247,N_12831);
or U13635 (N_13635,N_12206,N_12232);
or U13636 (N_13636,N_12157,N_12632);
or U13637 (N_13637,N_12157,N_12198);
nand U13638 (N_13638,N_12123,N_12511);
nor U13639 (N_13639,N_12693,N_12321);
nand U13640 (N_13640,N_12453,N_12474);
nand U13641 (N_13641,N_12252,N_12163);
nand U13642 (N_13642,N_12575,N_12703);
nand U13643 (N_13643,N_12814,N_12857);
and U13644 (N_13644,N_12517,N_12305);
and U13645 (N_13645,N_12145,N_12972);
or U13646 (N_13646,N_12430,N_12057);
nand U13647 (N_13647,N_12631,N_12852);
xor U13648 (N_13648,N_12684,N_12952);
nor U13649 (N_13649,N_12718,N_12540);
and U13650 (N_13650,N_12630,N_12160);
nand U13651 (N_13651,N_12913,N_12150);
xor U13652 (N_13652,N_12974,N_12593);
and U13653 (N_13653,N_12116,N_12013);
nand U13654 (N_13654,N_12142,N_12636);
nor U13655 (N_13655,N_12527,N_12666);
nand U13656 (N_13656,N_12915,N_12610);
or U13657 (N_13657,N_12116,N_12378);
nor U13658 (N_13658,N_12214,N_12731);
and U13659 (N_13659,N_12121,N_12372);
xnor U13660 (N_13660,N_12978,N_12577);
xnor U13661 (N_13661,N_12251,N_12809);
nor U13662 (N_13662,N_12898,N_12514);
nor U13663 (N_13663,N_12795,N_12782);
nand U13664 (N_13664,N_12101,N_12698);
nor U13665 (N_13665,N_12551,N_12479);
xnor U13666 (N_13666,N_12244,N_12035);
and U13667 (N_13667,N_12158,N_12203);
nand U13668 (N_13668,N_12496,N_12262);
or U13669 (N_13669,N_12297,N_12974);
and U13670 (N_13670,N_12351,N_12589);
nand U13671 (N_13671,N_12324,N_12131);
and U13672 (N_13672,N_12613,N_12164);
xor U13673 (N_13673,N_12438,N_12988);
xor U13674 (N_13674,N_12832,N_12778);
nand U13675 (N_13675,N_12266,N_12411);
xor U13676 (N_13676,N_12488,N_12478);
or U13677 (N_13677,N_12323,N_12656);
xor U13678 (N_13678,N_12522,N_12239);
nand U13679 (N_13679,N_12476,N_12013);
nor U13680 (N_13680,N_12832,N_12080);
or U13681 (N_13681,N_12025,N_12570);
and U13682 (N_13682,N_12388,N_12487);
xnor U13683 (N_13683,N_12348,N_12672);
or U13684 (N_13684,N_12762,N_12385);
or U13685 (N_13685,N_12934,N_12414);
and U13686 (N_13686,N_12453,N_12402);
xor U13687 (N_13687,N_12529,N_12717);
nor U13688 (N_13688,N_12356,N_12305);
or U13689 (N_13689,N_12654,N_12768);
and U13690 (N_13690,N_12123,N_12522);
nor U13691 (N_13691,N_12722,N_12315);
xor U13692 (N_13692,N_12290,N_12573);
or U13693 (N_13693,N_12378,N_12125);
and U13694 (N_13694,N_12181,N_12567);
nor U13695 (N_13695,N_12644,N_12734);
nor U13696 (N_13696,N_12751,N_12573);
and U13697 (N_13697,N_12428,N_12243);
nand U13698 (N_13698,N_12645,N_12807);
and U13699 (N_13699,N_12823,N_12635);
nand U13700 (N_13700,N_12694,N_12137);
and U13701 (N_13701,N_12791,N_12112);
xnor U13702 (N_13702,N_12574,N_12344);
xnor U13703 (N_13703,N_12095,N_12264);
xor U13704 (N_13704,N_12445,N_12228);
or U13705 (N_13705,N_12892,N_12470);
or U13706 (N_13706,N_12392,N_12554);
or U13707 (N_13707,N_12295,N_12159);
and U13708 (N_13708,N_12349,N_12653);
and U13709 (N_13709,N_12842,N_12991);
and U13710 (N_13710,N_12122,N_12866);
nor U13711 (N_13711,N_12073,N_12559);
or U13712 (N_13712,N_12798,N_12168);
and U13713 (N_13713,N_12655,N_12352);
or U13714 (N_13714,N_12875,N_12633);
or U13715 (N_13715,N_12677,N_12754);
nand U13716 (N_13716,N_12238,N_12827);
and U13717 (N_13717,N_12820,N_12882);
xor U13718 (N_13718,N_12198,N_12033);
and U13719 (N_13719,N_12530,N_12617);
nor U13720 (N_13720,N_12907,N_12602);
xor U13721 (N_13721,N_12725,N_12107);
nand U13722 (N_13722,N_12320,N_12535);
and U13723 (N_13723,N_12902,N_12672);
nor U13724 (N_13724,N_12708,N_12000);
and U13725 (N_13725,N_12397,N_12977);
xor U13726 (N_13726,N_12223,N_12751);
and U13727 (N_13727,N_12488,N_12607);
nand U13728 (N_13728,N_12435,N_12024);
and U13729 (N_13729,N_12199,N_12174);
nand U13730 (N_13730,N_12932,N_12960);
nor U13731 (N_13731,N_12010,N_12652);
nor U13732 (N_13732,N_12593,N_12034);
or U13733 (N_13733,N_12810,N_12844);
nor U13734 (N_13734,N_12230,N_12406);
xnor U13735 (N_13735,N_12000,N_12488);
nand U13736 (N_13736,N_12529,N_12820);
and U13737 (N_13737,N_12949,N_12737);
and U13738 (N_13738,N_12573,N_12249);
xnor U13739 (N_13739,N_12513,N_12327);
nor U13740 (N_13740,N_12783,N_12285);
nand U13741 (N_13741,N_12140,N_12057);
nor U13742 (N_13742,N_12405,N_12224);
nor U13743 (N_13743,N_12941,N_12211);
or U13744 (N_13744,N_12380,N_12265);
nand U13745 (N_13745,N_12407,N_12435);
xor U13746 (N_13746,N_12632,N_12502);
xnor U13747 (N_13747,N_12322,N_12034);
nand U13748 (N_13748,N_12270,N_12184);
nand U13749 (N_13749,N_12396,N_12982);
xor U13750 (N_13750,N_12451,N_12050);
or U13751 (N_13751,N_12883,N_12647);
or U13752 (N_13752,N_12141,N_12001);
nor U13753 (N_13753,N_12777,N_12406);
or U13754 (N_13754,N_12983,N_12548);
nand U13755 (N_13755,N_12638,N_12546);
xor U13756 (N_13756,N_12256,N_12451);
and U13757 (N_13757,N_12148,N_12863);
nand U13758 (N_13758,N_12811,N_12315);
xnor U13759 (N_13759,N_12766,N_12952);
xor U13760 (N_13760,N_12406,N_12101);
xnor U13761 (N_13761,N_12960,N_12312);
nor U13762 (N_13762,N_12146,N_12164);
and U13763 (N_13763,N_12135,N_12341);
and U13764 (N_13764,N_12192,N_12461);
nand U13765 (N_13765,N_12744,N_12591);
and U13766 (N_13766,N_12457,N_12790);
nand U13767 (N_13767,N_12483,N_12167);
or U13768 (N_13768,N_12888,N_12634);
and U13769 (N_13769,N_12064,N_12900);
and U13770 (N_13770,N_12578,N_12278);
or U13771 (N_13771,N_12959,N_12078);
xnor U13772 (N_13772,N_12267,N_12523);
or U13773 (N_13773,N_12413,N_12816);
nand U13774 (N_13774,N_12800,N_12136);
nand U13775 (N_13775,N_12150,N_12600);
nand U13776 (N_13776,N_12550,N_12183);
xor U13777 (N_13777,N_12677,N_12709);
and U13778 (N_13778,N_12819,N_12077);
nand U13779 (N_13779,N_12146,N_12762);
xor U13780 (N_13780,N_12888,N_12097);
nor U13781 (N_13781,N_12169,N_12399);
nor U13782 (N_13782,N_12149,N_12842);
xor U13783 (N_13783,N_12591,N_12460);
and U13784 (N_13784,N_12407,N_12888);
or U13785 (N_13785,N_12418,N_12025);
nor U13786 (N_13786,N_12297,N_12619);
or U13787 (N_13787,N_12803,N_12621);
nand U13788 (N_13788,N_12406,N_12838);
nor U13789 (N_13789,N_12687,N_12337);
and U13790 (N_13790,N_12847,N_12223);
nand U13791 (N_13791,N_12408,N_12847);
or U13792 (N_13792,N_12470,N_12309);
xnor U13793 (N_13793,N_12876,N_12713);
nand U13794 (N_13794,N_12461,N_12454);
and U13795 (N_13795,N_12243,N_12065);
and U13796 (N_13796,N_12861,N_12345);
nor U13797 (N_13797,N_12711,N_12998);
xor U13798 (N_13798,N_12076,N_12682);
or U13799 (N_13799,N_12801,N_12876);
xor U13800 (N_13800,N_12096,N_12363);
nand U13801 (N_13801,N_12567,N_12778);
and U13802 (N_13802,N_12915,N_12977);
xor U13803 (N_13803,N_12741,N_12998);
and U13804 (N_13804,N_12568,N_12111);
or U13805 (N_13805,N_12250,N_12649);
nor U13806 (N_13806,N_12651,N_12737);
nor U13807 (N_13807,N_12694,N_12777);
or U13808 (N_13808,N_12109,N_12616);
nand U13809 (N_13809,N_12147,N_12269);
or U13810 (N_13810,N_12139,N_12591);
or U13811 (N_13811,N_12841,N_12496);
or U13812 (N_13812,N_12305,N_12395);
or U13813 (N_13813,N_12033,N_12956);
xor U13814 (N_13814,N_12203,N_12648);
or U13815 (N_13815,N_12613,N_12939);
and U13816 (N_13816,N_12738,N_12609);
or U13817 (N_13817,N_12952,N_12176);
or U13818 (N_13818,N_12662,N_12131);
xor U13819 (N_13819,N_12384,N_12536);
nand U13820 (N_13820,N_12292,N_12203);
and U13821 (N_13821,N_12486,N_12580);
xor U13822 (N_13822,N_12619,N_12709);
nor U13823 (N_13823,N_12109,N_12358);
nand U13824 (N_13824,N_12782,N_12847);
or U13825 (N_13825,N_12135,N_12460);
nor U13826 (N_13826,N_12736,N_12897);
xnor U13827 (N_13827,N_12289,N_12495);
nor U13828 (N_13828,N_12570,N_12381);
and U13829 (N_13829,N_12952,N_12296);
or U13830 (N_13830,N_12039,N_12336);
or U13831 (N_13831,N_12912,N_12268);
or U13832 (N_13832,N_12256,N_12427);
and U13833 (N_13833,N_12598,N_12365);
nor U13834 (N_13834,N_12875,N_12210);
nand U13835 (N_13835,N_12002,N_12919);
nor U13836 (N_13836,N_12767,N_12450);
and U13837 (N_13837,N_12602,N_12246);
xor U13838 (N_13838,N_12789,N_12679);
nor U13839 (N_13839,N_12041,N_12336);
nand U13840 (N_13840,N_12465,N_12070);
nand U13841 (N_13841,N_12309,N_12370);
or U13842 (N_13842,N_12385,N_12422);
nand U13843 (N_13843,N_12373,N_12718);
xnor U13844 (N_13844,N_12841,N_12060);
and U13845 (N_13845,N_12535,N_12991);
nand U13846 (N_13846,N_12478,N_12595);
or U13847 (N_13847,N_12066,N_12475);
nand U13848 (N_13848,N_12842,N_12024);
nand U13849 (N_13849,N_12047,N_12343);
or U13850 (N_13850,N_12090,N_12299);
nand U13851 (N_13851,N_12965,N_12627);
xor U13852 (N_13852,N_12138,N_12773);
and U13853 (N_13853,N_12548,N_12367);
or U13854 (N_13854,N_12763,N_12192);
nand U13855 (N_13855,N_12621,N_12687);
xor U13856 (N_13856,N_12623,N_12351);
nand U13857 (N_13857,N_12619,N_12325);
nor U13858 (N_13858,N_12236,N_12951);
and U13859 (N_13859,N_12298,N_12024);
nor U13860 (N_13860,N_12738,N_12473);
nand U13861 (N_13861,N_12710,N_12515);
nor U13862 (N_13862,N_12791,N_12582);
nand U13863 (N_13863,N_12407,N_12421);
xor U13864 (N_13864,N_12185,N_12077);
nor U13865 (N_13865,N_12134,N_12565);
xnor U13866 (N_13866,N_12180,N_12434);
or U13867 (N_13867,N_12502,N_12906);
nand U13868 (N_13868,N_12285,N_12697);
or U13869 (N_13869,N_12942,N_12861);
nor U13870 (N_13870,N_12252,N_12208);
nor U13871 (N_13871,N_12833,N_12254);
and U13872 (N_13872,N_12116,N_12971);
nand U13873 (N_13873,N_12876,N_12989);
xnor U13874 (N_13874,N_12766,N_12901);
nor U13875 (N_13875,N_12085,N_12994);
nand U13876 (N_13876,N_12826,N_12788);
or U13877 (N_13877,N_12556,N_12175);
and U13878 (N_13878,N_12681,N_12910);
nor U13879 (N_13879,N_12134,N_12208);
nor U13880 (N_13880,N_12732,N_12357);
nor U13881 (N_13881,N_12670,N_12150);
and U13882 (N_13882,N_12563,N_12492);
nor U13883 (N_13883,N_12069,N_12678);
and U13884 (N_13884,N_12297,N_12970);
or U13885 (N_13885,N_12988,N_12803);
xnor U13886 (N_13886,N_12192,N_12702);
nand U13887 (N_13887,N_12053,N_12566);
xnor U13888 (N_13888,N_12986,N_12961);
and U13889 (N_13889,N_12718,N_12444);
nor U13890 (N_13890,N_12776,N_12224);
and U13891 (N_13891,N_12770,N_12802);
and U13892 (N_13892,N_12231,N_12816);
xor U13893 (N_13893,N_12382,N_12747);
or U13894 (N_13894,N_12980,N_12076);
xnor U13895 (N_13895,N_12469,N_12231);
nor U13896 (N_13896,N_12640,N_12618);
xor U13897 (N_13897,N_12415,N_12201);
and U13898 (N_13898,N_12329,N_12923);
and U13899 (N_13899,N_12485,N_12982);
nand U13900 (N_13900,N_12170,N_12552);
and U13901 (N_13901,N_12141,N_12089);
and U13902 (N_13902,N_12222,N_12389);
xor U13903 (N_13903,N_12468,N_12629);
nor U13904 (N_13904,N_12383,N_12706);
and U13905 (N_13905,N_12657,N_12847);
and U13906 (N_13906,N_12727,N_12460);
or U13907 (N_13907,N_12804,N_12648);
or U13908 (N_13908,N_12645,N_12131);
and U13909 (N_13909,N_12282,N_12521);
nand U13910 (N_13910,N_12123,N_12862);
xnor U13911 (N_13911,N_12415,N_12747);
nand U13912 (N_13912,N_12163,N_12801);
xor U13913 (N_13913,N_12872,N_12499);
xnor U13914 (N_13914,N_12734,N_12555);
or U13915 (N_13915,N_12070,N_12632);
nand U13916 (N_13916,N_12005,N_12414);
and U13917 (N_13917,N_12065,N_12910);
nor U13918 (N_13918,N_12993,N_12339);
xor U13919 (N_13919,N_12602,N_12804);
nor U13920 (N_13920,N_12779,N_12170);
nor U13921 (N_13921,N_12711,N_12704);
nor U13922 (N_13922,N_12586,N_12334);
and U13923 (N_13923,N_12903,N_12478);
nor U13924 (N_13924,N_12950,N_12851);
or U13925 (N_13925,N_12262,N_12223);
nand U13926 (N_13926,N_12918,N_12433);
xor U13927 (N_13927,N_12723,N_12773);
xor U13928 (N_13928,N_12448,N_12456);
nor U13929 (N_13929,N_12131,N_12937);
xor U13930 (N_13930,N_12199,N_12212);
and U13931 (N_13931,N_12085,N_12484);
nor U13932 (N_13932,N_12954,N_12905);
and U13933 (N_13933,N_12955,N_12602);
or U13934 (N_13934,N_12456,N_12227);
nand U13935 (N_13935,N_12922,N_12950);
or U13936 (N_13936,N_12985,N_12048);
or U13937 (N_13937,N_12831,N_12302);
nor U13938 (N_13938,N_12058,N_12156);
nand U13939 (N_13939,N_12815,N_12791);
and U13940 (N_13940,N_12983,N_12145);
nor U13941 (N_13941,N_12559,N_12428);
nand U13942 (N_13942,N_12834,N_12066);
nand U13943 (N_13943,N_12602,N_12344);
nor U13944 (N_13944,N_12462,N_12106);
nand U13945 (N_13945,N_12059,N_12935);
xor U13946 (N_13946,N_12769,N_12737);
nor U13947 (N_13947,N_12338,N_12937);
nand U13948 (N_13948,N_12766,N_12919);
or U13949 (N_13949,N_12417,N_12635);
xor U13950 (N_13950,N_12314,N_12342);
or U13951 (N_13951,N_12270,N_12906);
and U13952 (N_13952,N_12477,N_12304);
nor U13953 (N_13953,N_12235,N_12329);
or U13954 (N_13954,N_12771,N_12129);
nor U13955 (N_13955,N_12566,N_12353);
or U13956 (N_13956,N_12862,N_12806);
nor U13957 (N_13957,N_12865,N_12272);
xor U13958 (N_13958,N_12714,N_12209);
and U13959 (N_13959,N_12048,N_12247);
xor U13960 (N_13960,N_12098,N_12783);
nand U13961 (N_13961,N_12974,N_12975);
and U13962 (N_13962,N_12712,N_12035);
nor U13963 (N_13963,N_12525,N_12703);
and U13964 (N_13964,N_12175,N_12025);
xor U13965 (N_13965,N_12227,N_12846);
xor U13966 (N_13966,N_12180,N_12610);
xor U13967 (N_13967,N_12716,N_12934);
xnor U13968 (N_13968,N_12840,N_12043);
nor U13969 (N_13969,N_12511,N_12035);
and U13970 (N_13970,N_12468,N_12294);
xnor U13971 (N_13971,N_12721,N_12175);
and U13972 (N_13972,N_12830,N_12282);
nand U13973 (N_13973,N_12859,N_12391);
nand U13974 (N_13974,N_12018,N_12079);
or U13975 (N_13975,N_12336,N_12865);
nand U13976 (N_13976,N_12771,N_12130);
xnor U13977 (N_13977,N_12579,N_12655);
and U13978 (N_13978,N_12171,N_12911);
or U13979 (N_13979,N_12991,N_12812);
and U13980 (N_13980,N_12979,N_12115);
nor U13981 (N_13981,N_12898,N_12656);
nor U13982 (N_13982,N_12201,N_12363);
xor U13983 (N_13983,N_12177,N_12851);
nor U13984 (N_13984,N_12429,N_12970);
nor U13985 (N_13985,N_12851,N_12689);
xnor U13986 (N_13986,N_12895,N_12941);
xnor U13987 (N_13987,N_12537,N_12553);
nor U13988 (N_13988,N_12696,N_12192);
and U13989 (N_13989,N_12185,N_12415);
nor U13990 (N_13990,N_12958,N_12856);
xnor U13991 (N_13991,N_12388,N_12634);
nand U13992 (N_13992,N_12610,N_12886);
nand U13993 (N_13993,N_12342,N_12398);
or U13994 (N_13994,N_12433,N_12507);
or U13995 (N_13995,N_12178,N_12729);
nor U13996 (N_13996,N_12483,N_12135);
nor U13997 (N_13997,N_12527,N_12732);
xnor U13998 (N_13998,N_12341,N_12273);
and U13999 (N_13999,N_12718,N_12311);
xnor U14000 (N_14000,N_13060,N_13304);
or U14001 (N_14001,N_13821,N_13401);
nand U14002 (N_14002,N_13800,N_13273);
and U14003 (N_14003,N_13012,N_13965);
xnor U14004 (N_14004,N_13994,N_13698);
nand U14005 (N_14005,N_13468,N_13536);
or U14006 (N_14006,N_13601,N_13000);
nor U14007 (N_14007,N_13515,N_13549);
nand U14008 (N_14008,N_13688,N_13371);
nor U14009 (N_14009,N_13096,N_13015);
nand U14010 (N_14010,N_13827,N_13560);
and U14011 (N_14011,N_13807,N_13646);
and U14012 (N_14012,N_13850,N_13322);
xor U14013 (N_14013,N_13610,N_13219);
or U14014 (N_14014,N_13491,N_13106);
nor U14015 (N_14015,N_13317,N_13641);
xor U14016 (N_14016,N_13482,N_13848);
or U14017 (N_14017,N_13225,N_13064);
xnor U14018 (N_14018,N_13768,N_13962);
or U14019 (N_14019,N_13525,N_13657);
nand U14020 (N_14020,N_13707,N_13624);
nor U14021 (N_14021,N_13861,N_13543);
and U14022 (N_14022,N_13414,N_13142);
nor U14023 (N_14023,N_13160,N_13739);
nand U14024 (N_14024,N_13383,N_13891);
nand U14025 (N_14025,N_13443,N_13576);
xnor U14026 (N_14026,N_13280,N_13464);
nand U14027 (N_14027,N_13944,N_13666);
xnor U14028 (N_14028,N_13897,N_13833);
or U14029 (N_14029,N_13025,N_13094);
nand U14030 (N_14030,N_13871,N_13867);
nand U14031 (N_14031,N_13539,N_13481);
nor U14032 (N_14032,N_13282,N_13089);
nor U14033 (N_14033,N_13928,N_13356);
or U14034 (N_14034,N_13756,N_13039);
or U14035 (N_14035,N_13426,N_13895);
nor U14036 (N_14036,N_13979,N_13830);
xnor U14037 (N_14037,N_13817,N_13763);
or U14038 (N_14038,N_13520,N_13375);
or U14039 (N_14039,N_13990,N_13785);
nor U14040 (N_14040,N_13099,N_13198);
nand U14041 (N_14041,N_13090,N_13981);
and U14042 (N_14042,N_13831,N_13595);
or U14043 (N_14043,N_13622,N_13287);
nor U14044 (N_14044,N_13795,N_13163);
and U14045 (N_14045,N_13521,N_13858);
xnor U14046 (N_14046,N_13700,N_13947);
nor U14047 (N_14047,N_13672,N_13948);
nand U14048 (N_14048,N_13853,N_13669);
nand U14049 (N_14049,N_13145,N_13769);
or U14050 (N_14050,N_13903,N_13792);
and U14051 (N_14051,N_13321,N_13194);
nor U14052 (N_14052,N_13983,N_13725);
or U14053 (N_14053,N_13599,N_13136);
nand U14054 (N_14054,N_13139,N_13936);
xor U14055 (N_14055,N_13483,N_13606);
nand U14056 (N_14056,N_13146,N_13774);
nor U14057 (N_14057,N_13271,N_13393);
nand U14058 (N_14058,N_13233,N_13899);
nor U14059 (N_14059,N_13221,N_13002);
xor U14060 (N_14060,N_13682,N_13333);
and U14061 (N_14061,N_13737,N_13016);
nor U14062 (N_14062,N_13202,N_13806);
or U14063 (N_14063,N_13373,N_13938);
nand U14064 (N_14064,N_13721,N_13924);
and U14065 (N_14065,N_13722,N_13809);
xor U14066 (N_14066,N_13068,N_13926);
xnor U14067 (N_14067,N_13603,N_13093);
or U14068 (N_14068,N_13746,N_13476);
or U14069 (N_14069,N_13592,N_13578);
nand U14070 (N_14070,N_13971,N_13961);
or U14071 (N_14071,N_13442,N_13751);
xnor U14072 (N_14072,N_13253,N_13241);
nor U14073 (N_14073,N_13034,N_13446);
nor U14074 (N_14074,N_13913,N_13767);
xnor U14075 (N_14075,N_13571,N_13638);
and U14076 (N_14076,N_13863,N_13656);
xnor U14077 (N_14077,N_13609,N_13151);
or U14078 (N_14078,N_13019,N_13797);
and U14079 (N_14079,N_13449,N_13305);
nand U14080 (N_14080,N_13963,N_13229);
and U14081 (N_14081,N_13480,N_13881);
and U14082 (N_14082,N_13055,N_13101);
nand U14083 (N_14083,N_13862,N_13598);
xor U14084 (N_14084,N_13250,N_13900);
nand U14085 (N_14085,N_13613,N_13181);
or U14086 (N_14086,N_13020,N_13479);
xnor U14087 (N_14087,N_13615,N_13484);
xor U14088 (N_14088,N_13757,N_13411);
nor U14089 (N_14089,N_13402,N_13995);
or U14090 (N_14090,N_13395,N_13906);
or U14091 (N_14091,N_13380,N_13868);
or U14092 (N_14092,N_13196,N_13980);
or U14093 (N_14093,N_13689,N_13943);
xor U14094 (N_14094,N_13041,N_13759);
and U14095 (N_14095,N_13619,N_13355);
or U14096 (N_14096,N_13193,N_13950);
and U14097 (N_14097,N_13789,N_13206);
xor U14098 (N_14098,N_13550,N_13318);
nor U14099 (N_14099,N_13132,N_13937);
nand U14100 (N_14100,N_13120,N_13665);
and U14101 (N_14101,N_13554,N_13008);
xnor U14102 (N_14102,N_13410,N_13274);
nand U14103 (N_14103,N_13220,N_13859);
or U14104 (N_14104,N_13372,N_13922);
xnor U14105 (N_14105,N_13191,N_13330);
or U14106 (N_14106,N_13964,N_13458);
nand U14107 (N_14107,N_13643,N_13088);
or U14108 (N_14108,N_13137,N_13880);
nand U14109 (N_14109,N_13738,N_13557);
and U14110 (N_14110,N_13057,N_13566);
xor U14111 (N_14111,N_13231,N_13061);
and U14112 (N_14112,N_13620,N_13664);
nand U14113 (N_14113,N_13329,N_13532);
nand U14114 (N_14114,N_13832,N_13600);
xnor U14115 (N_14115,N_13676,N_13349);
nor U14116 (N_14116,N_13546,N_13882);
or U14117 (N_14117,N_13284,N_13517);
or U14118 (N_14118,N_13626,N_13267);
nand U14119 (N_14119,N_13234,N_13720);
nor U14120 (N_14120,N_13201,N_13487);
xor U14121 (N_14121,N_13714,N_13819);
nor U14122 (N_14122,N_13248,N_13133);
and U14123 (N_14123,N_13946,N_13416);
xnor U14124 (N_14124,N_13929,N_13421);
and U14125 (N_14125,N_13548,N_13045);
xnor U14126 (N_14126,N_13417,N_13149);
nand U14127 (N_14127,N_13004,N_13156);
and U14128 (N_14128,N_13205,N_13199);
xnor U14129 (N_14129,N_13846,N_13864);
xnor U14130 (N_14130,N_13105,N_13810);
and U14131 (N_14131,N_13408,N_13392);
or U14132 (N_14132,N_13433,N_13171);
xor U14133 (N_14133,N_13912,N_13298);
and U14134 (N_14134,N_13777,N_13823);
or U14135 (N_14135,N_13790,N_13628);
xor U14136 (N_14136,N_13908,N_13813);
nor U14137 (N_14137,N_13308,N_13625);
nand U14138 (N_14138,N_13915,N_13854);
or U14139 (N_14139,N_13942,N_13818);
and U14140 (N_14140,N_13904,N_13118);
nor U14141 (N_14141,N_13424,N_13510);
nor U14142 (N_14142,N_13453,N_13377);
and U14143 (N_14143,N_13545,N_13765);
nand U14144 (N_14144,N_13358,N_13736);
nand U14145 (N_14145,N_13278,N_13100);
nand U14146 (N_14146,N_13635,N_13455);
and U14147 (N_14147,N_13050,N_13989);
nor U14148 (N_14148,N_13843,N_13754);
xnor U14149 (N_14149,N_13387,N_13583);
or U14150 (N_14150,N_13627,N_13243);
or U14151 (N_14151,N_13940,N_13300);
xnor U14152 (N_14152,N_13386,N_13214);
or U14153 (N_14153,N_13988,N_13872);
nand U14154 (N_14154,N_13239,N_13796);
nand U14155 (N_14155,N_13621,N_13452);
and U14156 (N_14156,N_13888,N_13388);
and U14157 (N_14157,N_13342,N_13072);
xor U14158 (N_14158,N_13430,N_13461);
and U14159 (N_14159,N_13423,N_13771);
nand U14160 (N_14160,N_13530,N_13135);
nor U14161 (N_14161,N_13091,N_13702);
or U14162 (N_14162,N_13037,N_13876);
or U14163 (N_14163,N_13889,N_13690);
nor U14164 (N_14164,N_13001,N_13884);
and U14165 (N_14165,N_13917,N_13164);
or U14166 (N_14166,N_13652,N_13561);
and U14167 (N_14167,N_13175,N_13814);
nand U14168 (N_14168,N_13230,N_13920);
nand U14169 (N_14169,N_13745,N_13028);
and U14170 (N_14170,N_13316,N_13828);
or U14171 (N_14171,N_13901,N_13459);
xnor U14172 (N_14172,N_13495,N_13324);
and U14173 (N_14173,N_13092,N_13653);
xnor U14174 (N_14174,N_13281,N_13679);
nand U14175 (N_14175,N_13974,N_13212);
nand U14176 (N_14176,N_13109,N_13159);
or U14177 (N_14177,N_13085,N_13634);
nand U14178 (N_14178,N_13123,N_13747);
and U14179 (N_14179,N_13066,N_13183);
nor U14180 (N_14180,N_13266,N_13617);
xnor U14181 (N_14181,N_13803,N_13017);
nor U14182 (N_14182,N_13121,N_13772);
nor U14183 (N_14183,N_13674,N_13647);
nand U14184 (N_14184,N_13079,N_13049);
or U14185 (N_14185,N_13435,N_13251);
xor U14186 (N_14186,N_13396,N_13701);
and U14187 (N_14187,N_13413,N_13187);
nor U14188 (N_14188,N_13293,N_13749);
nand U14189 (N_14189,N_13892,N_13642);
nor U14190 (N_14190,N_13629,N_13334);
xnor U14191 (N_14191,N_13492,N_13357);
or U14192 (N_14192,N_13633,N_13503);
nand U14193 (N_14193,N_13122,N_13933);
nand U14194 (N_14194,N_13462,N_13254);
or U14195 (N_14195,N_13894,N_13589);
nor U14196 (N_14196,N_13390,N_13501);
nor U14197 (N_14197,N_13706,N_13352);
xor U14198 (N_14198,N_13836,N_13051);
xor U14199 (N_14199,N_13125,N_13129);
and U14200 (N_14200,N_13968,N_13496);
or U14201 (N_14201,N_13153,N_13343);
and U14202 (N_14202,N_13215,N_13256);
nor U14203 (N_14203,N_13572,N_13580);
or U14204 (N_14204,N_13662,N_13987);
and U14205 (N_14205,N_13555,N_13842);
xor U14206 (N_14206,N_13941,N_13328);
nor U14207 (N_14207,N_13724,N_13457);
or U14208 (N_14208,N_13026,N_13385);
nand U14209 (N_14209,N_13607,N_13655);
xor U14210 (N_14210,N_13742,N_13338);
xor U14211 (N_14211,N_13602,N_13046);
nand U14212 (N_14212,N_13207,N_13346);
or U14213 (N_14213,N_13006,N_13313);
nand U14214 (N_14214,N_13162,N_13909);
nor U14215 (N_14215,N_13493,N_13568);
or U14216 (N_14216,N_13374,N_13053);
nor U14217 (N_14217,N_13570,N_13781);
and U14218 (N_14218,N_13031,N_13540);
and U14219 (N_14219,N_13878,N_13378);
or U14220 (N_14220,N_13058,N_13528);
or U14221 (N_14221,N_13584,N_13516);
nor U14222 (N_14222,N_13069,N_13154);
nand U14223 (N_14223,N_13114,N_13671);
nand U14224 (N_14224,N_13029,N_13363);
xor U14225 (N_14225,N_13873,N_13640);
nand U14226 (N_14226,N_13816,N_13575);
xor U14227 (N_14227,N_13509,N_13117);
nor U14228 (N_14228,N_13704,N_13518);
and U14229 (N_14229,N_13381,N_13222);
and U14230 (N_14230,N_13052,N_13727);
nor U14231 (N_14231,N_13477,N_13535);
nor U14232 (N_14232,N_13784,N_13422);
and U14233 (N_14233,N_13911,N_13348);
nor U14234 (N_14234,N_13223,N_13030);
or U14235 (N_14235,N_13276,N_13242);
or U14236 (N_14236,N_13717,N_13102);
nand U14237 (N_14237,N_13286,N_13003);
xor U14238 (N_14238,N_13531,N_13261);
and U14239 (N_14239,N_13519,N_13726);
xnor U14240 (N_14240,N_13775,N_13463);
nor U14241 (N_14241,N_13840,N_13984);
xnor U14242 (N_14242,N_13710,N_13070);
nor U14243 (N_14243,N_13131,N_13172);
nand U14244 (N_14244,N_13551,N_13793);
nor U14245 (N_14245,N_13692,N_13195);
nand U14246 (N_14246,N_13081,N_13986);
and U14247 (N_14247,N_13112,N_13699);
nor U14248 (N_14248,N_13982,N_13326);
xnor U14249 (N_14249,N_13779,N_13719);
nor U14250 (N_14250,N_13451,N_13712);
nand U14251 (N_14251,N_13812,N_13890);
nor U14252 (N_14252,N_13534,N_13958);
nand U14253 (N_14253,N_13921,N_13910);
and U14254 (N_14254,N_13246,N_13038);
xnor U14255 (N_14255,N_13320,N_13311);
xor U14256 (N_14256,N_13444,N_13157);
nand U14257 (N_14257,N_13847,N_13425);
or U14258 (N_14258,N_13384,N_13552);
xnor U14259 (N_14259,N_13167,N_13902);
or U14260 (N_14260,N_13932,N_13734);
or U14261 (N_14261,N_13299,N_13347);
or U14262 (N_14262,N_13776,N_13558);
xor U14263 (N_14263,N_13359,N_13748);
or U14264 (N_14264,N_13758,N_13778);
or U14265 (N_14265,N_13178,N_13339);
nor U14266 (N_14266,N_13954,N_13588);
nor U14267 (N_14267,N_13143,N_13465);
nand U14268 (N_14268,N_13428,N_13898);
nand U14269 (N_14269,N_13696,N_13024);
or U14270 (N_14270,N_13460,N_13930);
nor U14271 (N_14271,N_13504,N_13325);
and U14272 (N_14272,N_13907,N_13649);
xnor U14273 (N_14273,N_13885,N_13366);
xnor U14274 (N_14274,N_13547,N_13705);
and U14275 (N_14275,N_13997,N_13791);
or U14276 (N_14276,N_13750,N_13826);
and U14277 (N_14277,N_13508,N_13639);
xor U14278 (N_14278,N_13860,N_13432);
xor U14279 (N_14279,N_13730,N_13753);
nand U14280 (N_14280,N_13977,N_13469);
and U14281 (N_14281,N_13119,N_13200);
and U14282 (N_14282,N_13297,N_13337);
nor U14283 (N_14283,N_13269,N_13773);
and U14284 (N_14284,N_13086,N_13935);
and U14285 (N_14285,N_13309,N_13703);
or U14286 (N_14286,N_13232,N_13967);
xor U14287 (N_14287,N_13567,N_13927);
nand U14288 (N_14288,N_13562,N_13650);
xnor U14289 (N_14289,N_13755,N_13808);
nor U14290 (N_14290,N_13174,N_13033);
xnor U14291 (N_14291,N_13541,N_13802);
nor U14292 (N_14292,N_13953,N_13553);
and U14293 (N_14293,N_13027,N_13708);
or U14294 (N_14294,N_13593,N_13184);
xnor U14295 (N_14295,N_13694,N_13996);
xnor U14296 (N_14296,N_13668,N_13340);
and U14297 (N_14297,N_13467,N_13078);
xnor U14298 (N_14298,N_13506,N_13611);
and U14299 (N_14299,N_13262,N_13345);
and U14300 (N_14300,N_13713,N_13152);
or U14301 (N_14301,N_13365,N_13849);
xor U14302 (N_14302,N_13970,N_13569);
xor U14303 (N_14303,N_13059,N_13957);
and U14304 (N_14304,N_13955,N_13485);
and U14305 (N_14305,N_13018,N_13332);
nor U14306 (N_14306,N_13658,N_13914);
nand U14307 (N_14307,N_13080,N_13168);
xnor U14308 (N_14308,N_13400,N_13344);
or U14309 (N_14309,N_13670,N_13204);
or U14310 (N_14310,N_13361,N_13255);
or U14311 (N_14311,N_13277,N_13265);
nand U14312 (N_14312,N_13237,N_13073);
xnor U14313 (N_14313,N_13475,N_13845);
xnor U14314 (N_14314,N_13470,N_13923);
or U14315 (N_14315,N_13307,N_13667);
or U14316 (N_14316,N_13005,N_13040);
and U14317 (N_14317,N_13165,N_13407);
xnor U14318 (N_14318,N_13866,N_13839);
nand U14319 (N_14319,N_13811,N_13978);
nor U14320 (N_14320,N_13084,N_13675);
nor U14321 (N_14321,N_13939,N_13258);
xnor U14322 (N_14322,N_13870,N_13240);
nand U14323 (N_14323,N_13527,N_13244);
or U14324 (N_14324,N_13054,N_13208);
or U14325 (N_14325,N_13141,N_13973);
xor U14326 (N_14326,N_13382,N_13419);
and U14327 (N_14327,N_13283,N_13036);
nand U14328 (N_14328,N_13169,N_13764);
xor U14329 (N_14329,N_13681,N_13762);
nor U14330 (N_14330,N_13687,N_13404);
and U14331 (N_14331,N_13415,N_13011);
or U14332 (N_14332,N_13636,N_13966);
nand U14333 (N_14333,N_13732,N_13350);
xor U14334 (N_14334,N_13203,N_13454);
and U14335 (N_14335,N_13403,N_13450);
nor U14336 (N_14336,N_13429,N_13960);
or U14337 (N_14337,N_13216,N_13035);
or U14338 (N_14338,N_13585,N_13770);
xor U14339 (N_14339,N_13486,N_13440);
nand U14340 (N_14340,N_13209,N_13412);
and U14341 (N_14341,N_13507,N_13992);
or U14342 (N_14342,N_13150,N_13197);
nand U14343 (N_14343,N_13279,N_13362);
nand U14344 (N_14344,N_13677,N_13581);
nand U14345 (N_14345,N_13786,N_13113);
nand U14346 (N_14346,N_13218,N_13760);
and U14347 (N_14347,N_13788,N_13798);
xor U14348 (N_14348,N_13228,N_13761);
and U14349 (N_14349,N_13685,N_13499);
xor U14350 (N_14350,N_13632,N_13155);
xnor U14351 (N_14351,N_13680,N_13182);
nand U14352 (N_14352,N_13673,N_13063);
or U14353 (N_14353,N_13857,N_13161);
nor U14354 (N_14354,N_13740,N_13289);
xor U14355 (N_14355,N_13379,N_13735);
nor U14356 (N_14356,N_13787,N_13360);
nand U14357 (N_14357,N_13931,N_13693);
and U14358 (N_14358,N_13743,N_13124);
nand U14359 (N_14359,N_13918,N_13247);
nor U14360 (N_14360,N_13993,N_13841);
and U14361 (N_14361,N_13353,N_13292);
and U14362 (N_14362,N_13494,N_13166);
nor U14363 (N_14363,N_13523,N_13952);
nor U14364 (N_14364,N_13303,N_13447);
nand U14365 (N_14365,N_13341,N_13533);
or U14366 (N_14366,N_13822,N_13728);
xnor U14367 (N_14367,N_13076,N_13879);
xor U14368 (N_14368,N_13376,N_13563);
nand U14369 (N_14369,N_13513,N_13331);
and U14370 (N_14370,N_13586,N_13062);
nor U14371 (N_14371,N_13180,N_13043);
or U14372 (N_14372,N_13327,N_13731);
nand U14373 (N_14373,N_13874,N_13177);
nand U14374 (N_14374,N_13473,N_13236);
nor U14375 (N_14375,N_13288,N_13013);
or U14376 (N_14376,N_13559,N_13097);
nor U14377 (N_14377,N_13217,N_13522);
and U14378 (N_14378,N_13210,N_13556);
xnor U14379 (N_14379,N_13565,N_13009);
and U14380 (N_14380,N_13835,N_13956);
and U14381 (N_14381,N_13173,N_13301);
xor U14382 (N_14382,N_13082,N_13022);
and U14383 (N_14383,N_13014,N_13856);
xor U14384 (N_14384,N_13213,N_13498);
or U14385 (N_14385,N_13976,N_13893);
nand U14386 (N_14386,N_13110,N_13711);
and U14387 (N_14387,N_13295,N_13659);
nor U14388 (N_14388,N_13290,N_13252);
nor U14389 (N_14389,N_13466,N_13564);
nand U14390 (N_14390,N_13263,N_13896);
xor U14391 (N_14391,N_13147,N_13648);
xor U14392 (N_14392,N_13766,N_13654);
nand U14393 (N_14393,N_13975,N_13799);
nand U14394 (N_14394,N_13067,N_13075);
or U14395 (N_14395,N_13582,N_13820);
nand U14396 (N_14396,N_13406,N_13077);
nand U14397 (N_14397,N_13718,N_13354);
and U14398 (N_14398,N_13612,N_13695);
and U14399 (N_14399,N_13249,N_13644);
or U14400 (N_14400,N_13972,N_13691);
nand U14401 (N_14401,N_13837,N_13684);
nand U14402 (N_14402,N_13804,N_13497);
nand U14403 (N_14403,N_13637,N_13844);
and U14404 (N_14404,N_13431,N_13397);
xor U14405 (N_14405,N_13351,N_13886);
or U14406 (N_14406,N_13951,N_13056);
nor U14407 (N_14407,N_13597,N_13127);
and U14408 (N_14408,N_13716,N_13170);
nand U14409 (N_14409,N_13438,N_13529);
xnor U14410 (N_14410,N_13663,N_13919);
nand U14411 (N_14411,N_13176,N_13590);
and U14412 (N_14412,N_13591,N_13875);
nand U14413 (N_14413,N_13645,N_13264);
or U14414 (N_14414,N_13126,N_13370);
or U14415 (N_14415,N_13189,N_13852);
xnor U14416 (N_14416,N_13245,N_13065);
xor U14417 (N_14417,N_13969,N_13226);
nand U14418 (N_14418,N_13441,N_13103);
and U14419 (N_14419,N_13437,N_13587);
xor U14420 (N_14420,N_13855,N_13573);
and U14421 (N_14421,N_13021,N_13192);
nand U14422 (N_14422,N_13144,N_13047);
nand U14423 (N_14423,N_13185,N_13294);
or U14424 (N_14424,N_13405,N_13825);
nand U14425 (N_14425,N_13211,N_13445);
xor U14426 (N_14426,N_13782,N_13115);
and U14427 (N_14427,N_13511,N_13291);
xor U14428 (N_14428,N_13998,N_13098);
nand U14429 (N_14429,N_13780,N_13389);
or U14430 (N_14430,N_13474,N_13335);
nor U14431 (N_14431,N_13594,N_13869);
xor U14432 (N_14432,N_13733,N_13661);
nand U14433 (N_14433,N_13238,N_13614);
or U14434 (N_14434,N_13272,N_13715);
nor U14435 (N_14435,N_13887,N_13824);
nand U14436 (N_14436,N_13368,N_13838);
or U14437 (N_14437,N_13505,N_13427);
xnor U14438 (N_14438,N_13138,N_13783);
xnor U14439 (N_14439,N_13436,N_13865);
xor U14440 (N_14440,N_13829,N_13999);
and U14441 (N_14441,N_13116,N_13959);
nor U14442 (N_14442,N_13032,N_13805);
nand U14443 (N_14443,N_13631,N_13489);
and U14444 (N_14444,N_13851,N_13111);
nor U14445 (N_14445,N_13514,N_13394);
xnor U14446 (N_14446,N_13044,N_13439);
nor U14447 (N_14447,N_13456,N_13224);
and U14448 (N_14448,N_13490,N_13314);
or U14449 (N_14449,N_13618,N_13623);
xnor U14450 (N_14450,N_13678,N_13577);
nor U14451 (N_14451,N_13630,N_13128);
and U14452 (N_14452,N_13542,N_13296);
nor U14453 (N_14453,N_13660,N_13500);
nand U14454 (N_14454,N_13186,N_13148);
nor U14455 (N_14455,N_13190,N_13179);
nand U14456 (N_14456,N_13409,N_13596);
or U14457 (N_14457,N_13310,N_13537);
and U14458 (N_14458,N_13448,N_13488);
nor U14459 (N_14459,N_13158,N_13275);
and U14460 (N_14460,N_13399,N_13605);
nand U14461 (N_14461,N_13526,N_13877);
nor U14462 (N_14462,N_13709,N_13729);
or U14463 (N_14463,N_13834,N_13512);
nor U14464 (N_14464,N_13883,N_13323);
or U14465 (N_14465,N_13270,N_13074);
and U14466 (N_14466,N_13418,N_13235);
xor U14467 (N_14467,N_13188,N_13905);
nand U14468 (N_14468,N_13815,N_13130);
and U14469 (N_14469,N_13398,N_13471);
nand U14470 (N_14470,N_13794,N_13651);
nand U14471 (N_14471,N_13697,N_13524);
or U14472 (N_14472,N_13259,N_13312);
nor U14473 (N_14473,N_13007,N_13140);
or U14474 (N_14474,N_13744,N_13134);
nand U14475 (N_14475,N_13087,N_13574);
or U14476 (N_14476,N_13095,N_13604);
and U14477 (N_14477,N_13934,N_13420);
and U14478 (N_14478,N_13319,N_13391);
nand U14479 (N_14479,N_13925,N_13071);
nand U14480 (N_14480,N_13048,N_13579);
or U14481 (N_14481,N_13108,N_13916);
xnor U14482 (N_14482,N_13945,N_13741);
and U14483 (N_14483,N_13991,N_13538);
nor U14484 (N_14484,N_13502,N_13260);
and U14485 (N_14485,N_13801,N_13752);
or U14486 (N_14486,N_13949,N_13306);
nor U14487 (N_14487,N_13302,N_13478);
nor U14488 (N_14488,N_13616,N_13683);
or U14489 (N_14489,N_13083,N_13723);
nor U14490 (N_14490,N_13268,N_13104);
xor U14491 (N_14491,N_13364,N_13227);
and U14492 (N_14492,N_13023,N_13608);
nor U14493 (N_14493,N_13315,N_13686);
and U14494 (N_14494,N_13010,N_13042);
or U14495 (N_14495,N_13367,N_13544);
xnor U14496 (N_14496,N_13257,N_13472);
nand U14497 (N_14497,N_13285,N_13434);
nor U14498 (N_14498,N_13336,N_13369);
nor U14499 (N_14499,N_13985,N_13107);
nand U14500 (N_14500,N_13080,N_13473);
xor U14501 (N_14501,N_13139,N_13339);
xnor U14502 (N_14502,N_13050,N_13247);
xor U14503 (N_14503,N_13185,N_13135);
xnor U14504 (N_14504,N_13871,N_13866);
nor U14505 (N_14505,N_13336,N_13182);
nand U14506 (N_14506,N_13583,N_13761);
nand U14507 (N_14507,N_13712,N_13074);
nor U14508 (N_14508,N_13089,N_13655);
and U14509 (N_14509,N_13201,N_13296);
nand U14510 (N_14510,N_13803,N_13117);
nor U14511 (N_14511,N_13842,N_13582);
or U14512 (N_14512,N_13681,N_13160);
nor U14513 (N_14513,N_13938,N_13249);
or U14514 (N_14514,N_13725,N_13415);
and U14515 (N_14515,N_13753,N_13762);
or U14516 (N_14516,N_13394,N_13706);
nor U14517 (N_14517,N_13625,N_13046);
and U14518 (N_14518,N_13244,N_13606);
or U14519 (N_14519,N_13698,N_13493);
nand U14520 (N_14520,N_13468,N_13621);
xor U14521 (N_14521,N_13832,N_13304);
and U14522 (N_14522,N_13055,N_13941);
xnor U14523 (N_14523,N_13820,N_13991);
nand U14524 (N_14524,N_13510,N_13291);
and U14525 (N_14525,N_13052,N_13811);
xnor U14526 (N_14526,N_13724,N_13527);
and U14527 (N_14527,N_13849,N_13200);
or U14528 (N_14528,N_13292,N_13674);
xnor U14529 (N_14529,N_13261,N_13119);
nor U14530 (N_14530,N_13188,N_13630);
or U14531 (N_14531,N_13067,N_13129);
and U14532 (N_14532,N_13443,N_13434);
nor U14533 (N_14533,N_13022,N_13519);
nand U14534 (N_14534,N_13800,N_13289);
and U14535 (N_14535,N_13738,N_13623);
or U14536 (N_14536,N_13679,N_13006);
nand U14537 (N_14537,N_13531,N_13864);
xnor U14538 (N_14538,N_13936,N_13941);
or U14539 (N_14539,N_13268,N_13208);
xor U14540 (N_14540,N_13856,N_13976);
and U14541 (N_14541,N_13248,N_13851);
xor U14542 (N_14542,N_13760,N_13559);
and U14543 (N_14543,N_13578,N_13576);
nand U14544 (N_14544,N_13072,N_13805);
and U14545 (N_14545,N_13010,N_13095);
and U14546 (N_14546,N_13489,N_13685);
or U14547 (N_14547,N_13367,N_13725);
nand U14548 (N_14548,N_13157,N_13828);
nand U14549 (N_14549,N_13838,N_13151);
nor U14550 (N_14550,N_13387,N_13090);
nor U14551 (N_14551,N_13659,N_13052);
and U14552 (N_14552,N_13595,N_13647);
nand U14553 (N_14553,N_13885,N_13549);
nand U14554 (N_14554,N_13061,N_13271);
and U14555 (N_14555,N_13511,N_13998);
and U14556 (N_14556,N_13425,N_13492);
and U14557 (N_14557,N_13560,N_13639);
or U14558 (N_14558,N_13507,N_13610);
or U14559 (N_14559,N_13185,N_13577);
xnor U14560 (N_14560,N_13842,N_13471);
and U14561 (N_14561,N_13377,N_13489);
or U14562 (N_14562,N_13699,N_13618);
nor U14563 (N_14563,N_13133,N_13323);
or U14564 (N_14564,N_13966,N_13640);
nor U14565 (N_14565,N_13518,N_13989);
or U14566 (N_14566,N_13268,N_13138);
and U14567 (N_14567,N_13343,N_13665);
or U14568 (N_14568,N_13874,N_13239);
or U14569 (N_14569,N_13222,N_13646);
and U14570 (N_14570,N_13053,N_13991);
and U14571 (N_14571,N_13058,N_13998);
or U14572 (N_14572,N_13065,N_13448);
or U14573 (N_14573,N_13884,N_13268);
and U14574 (N_14574,N_13990,N_13079);
or U14575 (N_14575,N_13653,N_13277);
xor U14576 (N_14576,N_13617,N_13878);
xnor U14577 (N_14577,N_13080,N_13086);
nor U14578 (N_14578,N_13368,N_13966);
nand U14579 (N_14579,N_13216,N_13544);
and U14580 (N_14580,N_13537,N_13165);
or U14581 (N_14581,N_13922,N_13755);
nor U14582 (N_14582,N_13069,N_13376);
nor U14583 (N_14583,N_13754,N_13095);
nor U14584 (N_14584,N_13399,N_13470);
xor U14585 (N_14585,N_13236,N_13556);
xnor U14586 (N_14586,N_13460,N_13986);
nor U14587 (N_14587,N_13269,N_13016);
nor U14588 (N_14588,N_13496,N_13044);
nor U14589 (N_14589,N_13996,N_13726);
or U14590 (N_14590,N_13657,N_13741);
and U14591 (N_14591,N_13258,N_13225);
xnor U14592 (N_14592,N_13250,N_13724);
and U14593 (N_14593,N_13067,N_13108);
or U14594 (N_14594,N_13739,N_13223);
nand U14595 (N_14595,N_13483,N_13238);
xor U14596 (N_14596,N_13576,N_13313);
and U14597 (N_14597,N_13504,N_13256);
or U14598 (N_14598,N_13547,N_13320);
xor U14599 (N_14599,N_13075,N_13589);
or U14600 (N_14600,N_13557,N_13058);
xnor U14601 (N_14601,N_13337,N_13265);
or U14602 (N_14602,N_13181,N_13002);
or U14603 (N_14603,N_13648,N_13796);
nand U14604 (N_14604,N_13177,N_13977);
and U14605 (N_14605,N_13723,N_13010);
xnor U14606 (N_14606,N_13746,N_13106);
xor U14607 (N_14607,N_13730,N_13838);
xnor U14608 (N_14608,N_13467,N_13200);
and U14609 (N_14609,N_13591,N_13408);
nand U14610 (N_14610,N_13159,N_13821);
or U14611 (N_14611,N_13962,N_13670);
xor U14612 (N_14612,N_13867,N_13845);
nand U14613 (N_14613,N_13416,N_13900);
xnor U14614 (N_14614,N_13829,N_13329);
nor U14615 (N_14615,N_13820,N_13254);
nand U14616 (N_14616,N_13285,N_13546);
or U14617 (N_14617,N_13768,N_13054);
and U14618 (N_14618,N_13862,N_13461);
nor U14619 (N_14619,N_13475,N_13836);
nand U14620 (N_14620,N_13178,N_13215);
nor U14621 (N_14621,N_13429,N_13813);
xnor U14622 (N_14622,N_13286,N_13305);
xnor U14623 (N_14623,N_13876,N_13073);
nor U14624 (N_14624,N_13575,N_13866);
nor U14625 (N_14625,N_13649,N_13485);
and U14626 (N_14626,N_13150,N_13554);
or U14627 (N_14627,N_13084,N_13876);
nor U14628 (N_14628,N_13433,N_13190);
nand U14629 (N_14629,N_13193,N_13738);
and U14630 (N_14630,N_13343,N_13841);
and U14631 (N_14631,N_13873,N_13385);
xor U14632 (N_14632,N_13963,N_13701);
and U14633 (N_14633,N_13425,N_13950);
or U14634 (N_14634,N_13308,N_13585);
or U14635 (N_14635,N_13584,N_13874);
xnor U14636 (N_14636,N_13458,N_13220);
xor U14637 (N_14637,N_13570,N_13759);
nor U14638 (N_14638,N_13389,N_13206);
nand U14639 (N_14639,N_13631,N_13667);
xnor U14640 (N_14640,N_13576,N_13745);
nand U14641 (N_14641,N_13207,N_13710);
xnor U14642 (N_14642,N_13500,N_13598);
xor U14643 (N_14643,N_13798,N_13406);
xor U14644 (N_14644,N_13516,N_13166);
xor U14645 (N_14645,N_13568,N_13311);
and U14646 (N_14646,N_13212,N_13033);
nor U14647 (N_14647,N_13563,N_13718);
and U14648 (N_14648,N_13331,N_13134);
or U14649 (N_14649,N_13911,N_13602);
and U14650 (N_14650,N_13639,N_13482);
and U14651 (N_14651,N_13545,N_13835);
and U14652 (N_14652,N_13357,N_13404);
nand U14653 (N_14653,N_13667,N_13755);
and U14654 (N_14654,N_13640,N_13283);
nor U14655 (N_14655,N_13872,N_13579);
nand U14656 (N_14656,N_13163,N_13591);
xnor U14657 (N_14657,N_13428,N_13718);
nand U14658 (N_14658,N_13847,N_13569);
nor U14659 (N_14659,N_13421,N_13079);
or U14660 (N_14660,N_13336,N_13370);
and U14661 (N_14661,N_13628,N_13935);
nor U14662 (N_14662,N_13931,N_13395);
xor U14663 (N_14663,N_13408,N_13571);
and U14664 (N_14664,N_13264,N_13060);
xor U14665 (N_14665,N_13913,N_13617);
xnor U14666 (N_14666,N_13733,N_13444);
xnor U14667 (N_14667,N_13141,N_13440);
or U14668 (N_14668,N_13069,N_13441);
xnor U14669 (N_14669,N_13582,N_13733);
and U14670 (N_14670,N_13891,N_13157);
xnor U14671 (N_14671,N_13142,N_13736);
xnor U14672 (N_14672,N_13711,N_13405);
xnor U14673 (N_14673,N_13383,N_13845);
xor U14674 (N_14674,N_13591,N_13318);
xor U14675 (N_14675,N_13678,N_13384);
nor U14676 (N_14676,N_13601,N_13504);
nand U14677 (N_14677,N_13456,N_13193);
nor U14678 (N_14678,N_13281,N_13805);
and U14679 (N_14679,N_13294,N_13547);
and U14680 (N_14680,N_13897,N_13708);
or U14681 (N_14681,N_13834,N_13862);
and U14682 (N_14682,N_13073,N_13740);
and U14683 (N_14683,N_13409,N_13818);
nor U14684 (N_14684,N_13954,N_13672);
nor U14685 (N_14685,N_13865,N_13716);
or U14686 (N_14686,N_13026,N_13619);
and U14687 (N_14687,N_13833,N_13494);
or U14688 (N_14688,N_13994,N_13015);
xor U14689 (N_14689,N_13538,N_13701);
nor U14690 (N_14690,N_13431,N_13160);
xnor U14691 (N_14691,N_13257,N_13059);
or U14692 (N_14692,N_13159,N_13275);
xor U14693 (N_14693,N_13560,N_13052);
and U14694 (N_14694,N_13017,N_13204);
nor U14695 (N_14695,N_13195,N_13411);
nand U14696 (N_14696,N_13685,N_13020);
or U14697 (N_14697,N_13516,N_13134);
nand U14698 (N_14698,N_13393,N_13923);
nand U14699 (N_14699,N_13244,N_13229);
nand U14700 (N_14700,N_13954,N_13756);
xnor U14701 (N_14701,N_13110,N_13813);
and U14702 (N_14702,N_13933,N_13348);
nand U14703 (N_14703,N_13057,N_13042);
or U14704 (N_14704,N_13634,N_13979);
or U14705 (N_14705,N_13880,N_13976);
nand U14706 (N_14706,N_13728,N_13758);
nand U14707 (N_14707,N_13564,N_13768);
nand U14708 (N_14708,N_13504,N_13432);
and U14709 (N_14709,N_13106,N_13363);
and U14710 (N_14710,N_13830,N_13235);
xor U14711 (N_14711,N_13613,N_13316);
or U14712 (N_14712,N_13767,N_13351);
nand U14713 (N_14713,N_13005,N_13782);
nand U14714 (N_14714,N_13458,N_13658);
nand U14715 (N_14715,N_13351,N_13891);
nand U14716 (N_14716,N_13154,N_13941);
nand U14717 (N_14717,N_13607,N_13322);
xnor U14718 (N_14718,N_13208,N_13927);
nand U14719 (N_14719,N_13628,N_13728);
and U14720 (N_14720,N_13937,N_13987);
nor U14721 (N_14721,N_13218,N_13841);
or U14722 (N_14722,N_13590,N_13132);
and U14723 (N_14723,N_13079,N_13278);
or U14724 (N_14724,N_13992,N_13862);
or U14725 (N_14725,N_13011,N_13236);
nor U14726 (N_14726,N_13309,N_13976);
nand U14727 (N_14727,N_13480,N_13114);
xor U14728 (N_14728,N_13083,N_13655);
nand U14729 (N_14729,N_13566,N_13097);
xor U14730 (N_14730,N_13950,N_13829);
xor U14731 (N_14731,N_13065,N_13284);
and U14732 (N_14732,N_13381,N_13944);
nor U14733 (N_14733,N_13968,N_13010);
xnor U14734 (N_14734,N_13310,N_13783);
and U14735 (N_14735,N_13729,N_13800);
nor U14736 (N_14736,N_13879,N_13543);
or U14737 (N_14737,N_13446,N_13207);
nand U14738 (N_14738,N_13530,N_13086);
or U14739 (N_14739,N_13096,N_13759);
xnor U14740 (N_14740,N_13791,N_13470);
nor U14741 (N_14741,N_13264,N_13820);
and U14742 (N_14742,N_13008,N_13856);
nor U14743 (N_14743,N_13077,N_13893);
nor U14744 (N_14744,N_13811,N_13918);
nor U14745 (N_14745,N_13326,N_13985);
or U14746 (N_14746,N_13197,N_13381);
nor U14747 (N_14747,N_13126,N_13907);
nand U14748 (N_14748,N_13531,N_13745);
nand U14749 (N_14749,N_13286,N_13440);
and U14750 (N_14750,N_13009,N_13610);
or U14751 (N_14751,N_13315,N_13041);
xnor U14752 (N_14752,N_13608,N_13692);
or U14753 (N_14753,N_13141,N_13362);
or U14754 (N_14754,N_13810,N_13272);
nand U14755 (N_14755,N_13532,N_13572);
or U14756 (N_14756,N_13280,N_13483);
or U14757 (N_14757,N_13137,N_13013);
or U14758 (N_14758,N_13696,N_13510);
xor U14759 (N_14759,N_13275,N_13584);
and U14760 (N_14760,N_13319,N_13284);
nand U14761 (N_14761,N_13415,N_13625);
nand U14762 (N_14762,N_13193,N_13060);
nand U14763 (N_14763,N_13134,N_13532);
nor U14764 (N_14764,N_13269,N_13120);
nand U14765 (N_14765,N_13972,N_13989);
or U14766 (N_14766,N_13524,N_13049);
xnor U14767 (N_14767,N_13986,N_13670);
or U14768 (N_14768,N_13420,N_13143);
or U14769 (N_14769,N_13738,N_13426);
nor U14770 (N_14770,N_13591,N_13778);
xnor U14771 (N_14771,N_13409,N_13369);
nand U14772 (N_14772,N_13025,N_13682);
nor U14773 (N_14773,N_13144,N_13089);
and U14774 (N_14774,N_13182,N_13913);
xor U14775 (N_14775,N_13476,N_13779);
nor U14776 (N_14776,N_13697,N_13194);
nor U14777 (N_14777,N_13026,N_13267);
or U14778 (N_14778,N_13345,N_13327);
and U14779 (N_14779,N_13996,N_13216);
or U14780 (N_14780,N_13676,N_13991);
xnor U14781 (N_14781,N_13927,N_13291);
and U14782 (N_14782,N_13900,N_13537);
nor U14783 (N_14783,N_13504,N_13684);
and U14784 (N_14784,N_13770,N_13506);
and U14785 (N_14785,N_13990,N_13480);
nand U14786 (N_14786,N_13301,N_13792);
or U14787 (N_14787,N_13973,N_13171);
nor U14788 (N_14788,N_13131,N_13041);
nand U14789 (N_14789,N_13372,N_13727);
and U14790 (N_14790,N_13160,N_13706);
or U14791 (N_14791,N_13029,N_13938);
xor U14792 (N_14792,N_13059,N_13562);
or U14793 (N_14793,N_13739,N_13347);
and U14794 (N_14794,N_13734,N_13545);
nand U14795 (N_14795,N_13988,N_13171);
xnor U14796 (N_14796,N_13437,N_13364);
nor U14797 (N_14797,N_13952,N_13368);
xnor U14798 (N_14798,N_13918,N_13308);
or U14799 (N_14799,N_13988,N_13948);
xor U14800 (N_14800,N_13714,N_13525);
or U14801 (N_14801,N_13406,N_13272);
nor U14802 (N_14802,N_13886,N_13827);
or U14803 (N_14803,N_13770,N_13168);
xnor U14804 (N_14804,N_13675,N_13132);
and U14805 (N_14805,N_13236,N_13667);
nand U14806 (N_14806,N_13007,N_13660);
and U14807 (N_14807,N_13644,N_13990);
nand U14808 (N_14808,N_13960,N_13657);
and U14809 (N_14809,N_13953,N_13980);
and U14810 (N_14810,N_13954,N_13924);
and U14811 (N_14811,N_13874,N_13534);
xnor U14812 (N_14812,N_13945,N_13622);
nand U14813 (N_14813,N_13612,N_13168);
xor U14814 (N_14814,N_13961,N_13303);
xnor U14815 (N_14815,N_13304,N_13991);
xor U14816 (N_14816,N_13811,N_13981);
or U14817 (N_14817,N_13263,N_13774);
nand U14818 (N_14818,N_13045,N_13518);
or U14819 (N_14819,N_13936,N_13010);
xnor U14820 (N_14820,N_13543,N_13589);
nor U14821 (N_14821,N_13035,N_13129);
nand U14822 (N_14822,N_13436,N_13777);
xnor U14823 (N_14823,N_13493,N_13101);
or U14824 (N_14824,N_13467,N_13155);
nor U14825 (N_14825,N_13484,N_13460);
nor U14826 (N_14826,N_13256,N_13127);
xnor U14827 (N_14827,N_13969,N_13840);
xor U14828 (N_14828,N_13402,N_13291);
nand U14829 (N_14829,N_13222,N_13835);
or U14830 (N_14830,N_13739,N_13323);
nand U14831 (N_14831,N_13384,N_13233);
or U14832 (N_14832,N_13957,N_13866);
nand U14833 (N_14833,N_13208,N_13454);
nand U14834 (N_14834,N_13691,N_13646);
or U14835 (N_14835,N_13462,N_13313);
and U14836 (N_14836,N_13957,N_13994);
xor U14837 (N_14837,N_13463,N_13224);
nand U14838 (N_14838,N_13385,N_13042);
or U14839 (N_14839,N_13218,N_13401);
and U14840 (N_14840,N_13744,N_13789);
nand U14841 (N_14841,N_13790,N_13127);
nor U14842 (N_14842,N_13690,N_13246);
nor U14843 (N_14843,N_13645,N_13361);
or U14844 (N_14844,N_13124,N_13333);
or U14845 (N_14845,N_13318,N_13969);
and U14846 (N_14846,N_13845,N_13985);
nand U14847 (N_14847,N_13880,N_13889);
xor U14848 (N_14848,N_13638,N_13463);
nand U14849 (N_14849,N_13962,N_13764);
nor U14850 (N_14850,N_13604,N_13470);
or U14851 (N_14851,N_13815,N_13254);
and U14852 (N_14852,N_13782,N_13728);
xnor U14853 (N_14853,N_13826,N_13947);
nor U14854 (N_14854,N_13107,N_13070);
nor U14855 (N_14855,N_13725,N_13914);
and U14856 (N_14856,N_13818,N_13811);
xor U14857 (N_14857,N_13966,N_13419);
or U14858 (N_14858,N_13066,N_13247);
nor U14859 (N_14859,N_13340,N_13586);
or U14860 (N_14860,N_13880,N_13661);
nand U14861 (N_14861,N_13448,N_13359);
nand U14862 (N_14862,N_13233,N_13923);
xor U14863 (N_14863,N_13466,N_13806);
or U14864 (N_14864,N_13997,N_13506);
nand U14865 (N_14865,N_13905,N_13006);
or U14866 (N_14866,N_13028,N_13033);
or U14867 (N_14867,N_13888,N_13314);
or U14868 (N_14868,N_13944,N_13997);
and U14869 (N_14869,N_13833,N_13879);
and U14870 (N_14870,N_13923,N_13680);
or U14871 (N_14871,N_13668,N_13128);
and U14872 (N_14872,N_13031,N_13661);
or U14873 (N_14873,N_13418,N_13477);
xnor U14874 (N_14874,N_13387,N_13173);
nor U14875 (N_14875,N_13976,N_13094);
nand U14876 (N_14876,N_13305,N_13412);
nor U14877 (N_14877,N_13187,N_13415);
or U14878 (N_14878,N_13525,N_13967);
nand U14879 (N_14879,N_13435,N_13146);
nor U14880 (N_14880,N_13062,N_13464);
nand U14881 (N_14881,N_13804,N_13634);
nor U14882 (N_14882,N_13816,N_13046);
or U14883 (N_14883,N_13929,N_13930);
nor U14884 (N_14884,N_13566,N_13534);
or U14885 (N_14885,N_13234,N_13118);
or U14886 (N_14886,N_13196,N_13354);
nor U14887 (N_14887,N_13755,N_13078);
and U14888 (N_14888,N_13050,N_13080);
or U14889 (N_14889,N_13282,N_13594);
nor U14890 (N_14890,N_13248,N_13893);
xnor U14891 (N_14891,N_13667,N_13278);
nor U14892 (N_14892,N_13858,N_13900);
nand U14893 (N_14893,N_13366,N_13104);
nand U14894 (N_14894,N_13397,N_13748);
and U14895 (N_14895,N_13217,N_13094);
xnor U14896 (N_14896,N_13435,N_13377);
or U14897 (N_14897,N_13547,N_13485);
nor U14898 (N_14898,N_13821,N_13257);
nand U14899 (N_14899,N_13097,N_13791);
xor U14900 (N_14900,N_13616,N_13442);
and U14901 (N_14901,N_13152,N_13734);
and U14902 (N_14902,N_13276,N_13667);
or U14903 (N_14903,N_13629,N_13840);
nand U14904 (N_14904,N_13946,N_13165);
nor U14905 (N_14905,N_13864,N_13004);
nor U14906 (N_14906,N_13691,N_13039);
and U14907 (N_14907,N_13958,N_13297);
or U14908 (N_14908,N_13167,N_13203);
nor U14909 (N_14909,N_13368,N_13168);
nand U14910 (N_14910,N_13624,N_13291);
nand U14911 (N_14911,N_13091,N_13245);
nand U14912 (N_14912,N_13617,N_13221);
nor U14913 (N_14913,N_13281,N_13212);
or U14914 (N_14914,N_13440,N_13716);
and U14915 (N_14915,N_13873,N_13132);
or U14916 (N_14916,N_13850,N_13650);
nand U14917 (N_14917,N_13252,N_13043);
or U14918 (N_14918,N_13121,N_13299);
nor U14919 (N_14919,N_13762,N_13619);
or U14920 (N_14920,N_13472,N_13102);
and U14921 (N_14921,N_13687,N_13482);
nor U14922 (N_14922,N_13445,N_13292);
or U14923 (N_14923,N_13877,N_13197);
or U14924 (N_14924,N_13300,N_13732);
or U14925 (N_14925,N_13199,N_13686);
and U14926 (N_14926,N_13849,N_13155);
xnor U14927 (N_14927,N_13784,N_13080);
or U14928 (N_14928,N_13522,N_13092);
nor U14929 (N_14929,N_13424,N_13656);
nor U14930 (N_14930,N_13080,N_13150);
nor U14931 (N_14931,N_13885,N_13986);
nor U14932 (N_14932,N_13507,N_13138);
nor U14933 (N_14933,N_13265,N_13842);
nor U14934 (N_14934,N_13474,N_13664);
or U14935 (N_14935,N_13480,N_13165);
and U14936 (N_14936,N_13159,N_13403);
or U14937 (N_14937,N_13323,N_13782);
xor U14938 (N_14938,N_13766,N_13418);
xnor U14939 (N_14939,N_13693,N_13584);
nand U14940 (N_14940,N_13987,N_13836);
nor U14941 (N_14941,N_13443,N_13648);
or U14942 (N_14942,N_13185,N_13121);
nor U14943 (N_14943,N_13090,N_13841);
nand U14944 (N_14944,N_13393,N_13103);
nor U14945 (N_14945,N_13157,N_13390);
xor U14946 (N_14946,N_13412,N_13077);
nand U14947 (N_14947,N_13883,N_13822);
xnor U14948 (N_14948,N_13615,N_13849);
xnor U14949 (N_14949,N_13422,N_13622);
nand U14950 (N_14950,N_13423,N_13550);
xor U14951 (N_14951,N_13326,N_13612);
nand U14952 (N_14952,N_13281,N_13879);
and U14953 (N_14953,N_13997,N_13087);
and U14954 (N_14954,N_13467,N_13893);
and U14955 (N_14955,N_13973,N_13373);
nand U14956 (N_14956,N_13903,N_13221);
or U14957 (N_14957,N_13695,N_13430);
and U14958 (N_14958,N_13561,N_13957);
and U14959 (N_14959,N_13738,N_13968);
or U14960 (N_14960,N_13526,N_13486);
or U14961 (N_14961,N_13216,N_13167);
nor U14962 (N_14962,N_13493,N_13130);
xnor U14963 (N_14963,N_13220,N_13710);
or U14964 (N_14964,N_13875,N_13640);
nor U14965 (N_14965,N_13595,N_13401);
xor U14966 (N_14966,N_13537,N_13440);
nand U14967 (N_14967,N_13989,N_13497);
and U14968 (N_14968,N_13085,N_13274);
nor U14969 (N_14969,N_13089,N_13367);
nor U14970 (N_14970,N_13044,N_13258);
xor U14971 (N_14971,N_13693,N_13018);
nor U14972 (N_14972,N_13788,N_13447);
nand U14973 (N_14973,N_13909,N_13629);
nor U14974 (N_14974,N_13663,N_13736);
and U14975 (N_14975,N_13419,N_13486);
or U14976 (N_14976,N_13050,N_13032);
nor U14977 (N_14977,N_13913,N_13519);
or U14978 (N_14978,N_13658,N_13908);
or U14979 (N_14979,N_13251,N_13012);
and U14980 (N_14980,N_13552,N_13918);
nand U14981 (N_14981,N_13210,N_13126);
nor U14982 (N_14982,N_13328,N_13352);
and U14983 (N_14983,N_13602,N_13651);
or U14984 (N_14984,N_13714,N_13909);
and U14985 (N_14985,N_13967,N_13485);
nor U14986 (N_14986,N_13989,N_13889);
nor U14987 (N_14987,N_13196,N_13181);
and U14988 (N_14988,N_13873,N_13522);
and U14989 (N_14989,N_13555,N_13766);
nand U14990 (N_14990,N_13026,N_13877);
and U14991 (N_14991,N_13450,N_13291);
nor U14992 (N_14992,N_13379,N_13404);
xnor U14993 (N_14993,N_13361,N_13586);
xor U14994 (N_14994,N_13297,N_13125);
and U14995 (N_14995,N_13645,N_13693);
nor U14996 (N_14996,N_13085,N_13557);
and U14997 (N_14997,N_13337,N_13531);
nand U14998 (N_14998,N_13661,N_13970);
nor U14999 (N_14999,N_13632,N_13073);
and UO_0 (O_0,N_14880,N_14986);
and UO_1 (O_1,N_14599,N_14580);
nand UO_2 (O_2,N_14346,N_14250);
nor UO_3 (O_3,N_14710,N_14550);
or UO_4 (O_4,N_14517,N_14872);
and UO_5 (O_5,N_14001,N_14598);
xnor UO_6 (O_6,N_14273,N_14771);
and UO_7 (O_7,N_14094,N_14847);
or UO_8 (O_8,N_14744,N_14991);
xnor UO_9 (O_9,N_14063,N_14307);
and UO_10 (O_10,N_14352,N_14623);
nand UO_11 (O_11,N_14581,N_14306);
and UO_12 (O_12,N_14539,N_14182);
nand UO_13 (O_13,N_14037,N_14265);
nor UO_14 (O_14,N_14054,N_14261);
and UO_15 (O_15,N_14049,N_14120);
and UO_16 (O_16,N_14918,N_14336);
nor UO_17 (O_17,N_14369,N_14842);
or UO_18 (O_18,N_14435,N_14124);
xnor UO_19 (O_19,N_14401,N_14103);
and UO_20 (O_20,N_14209,N_14800);
nor UO_21 (O_21,N_14072,N_14434);
or UO_22 (O_22,N_14846,N_14108);
or UO_23 (O_23,N_14077,N_14560);
nand UO_24 (O_24,N_14805,N_14395);
nor UO_25 (O_25,N_14875,N_14714);
nand UO_26 (O_26,N_14231,N_14594);
nand UO_27 (O_27,N_14674,N_14389);
or UO_28 (O_28,N_14836,N_14948);
nor UO_29 (O_29,N_14184,N_14276);
and UO_30 (O_30,N_14571,N_14690);
nand UO_31 (O_31,N_14553,N_14582);
and UO_32 (O_32,N_14586,N_14126);
and UO_33 (O_33,N_14178,N_14425);
xor UO_34 (O_34,N_14959,N_14385);
or UO_35 (O_35,N_14937,N_14823);
and UO_36 (O_36,N_14953,N_14627);
and UO_37 (O_37,N_14381,N_14048);
nand UO_38 (O_38,N_14059,N_14679);
nor UO_39 (O_39,N_14529,N_14382);
xnor UO_40 (O_40,N_14631,N_14863);
and UO_41 (O_41,N_14018,N_14859);
nor UO_42 (O_42,N_14113,N_14405);
and UO_43 (O_43,N_14324,N_14669);
xor UO_44 (O_44,N_14721,N_14688);
nand UO_45 (O_45,N_14521,N_14082);
nand UO_46 (O_46,N_14839,N_14665);
nor UO_47 (O_47,N_14730,N_14228);
nand UO_48 (O_48,N_14096,N_14264);
or UO_49 (O_49,N_14145,N_14380);
or UO_50 (O_50,N_14466,N_14256);
nand UO_51 (O_51,N_14752,N_14632);
nand UO_52 (O_52,N_14568,N_14468);
nor UO_53 (O_53,N_14944,N_14375);
and UO_54 (O_54,N_14841,N_14007);
and UO_55 (O_55,N_14716,N_14756);
nand UO_56 (O_56,N_14292,N_14268);
nand UO_57 (O_57,N_14128,N_14153);
nand UO_58 (O_58,N_14759,N_14971);
or UO_59 (O_59,N_14777,N_14659);
or UO_60 (O_60,N_14740,N_14766);
nor UO_61 (O_61,N_14414,N_14350);
xnor UO_62 (O_62,N_14440,N_14574);
and UO_63 (O_63,N_14793,N_14232);
nor UO_64 (O_64,N_14281,N_14975);
and UO_65 (O_65,N_14023,N_14940);
xor UO_66 (O_66,N_14086,N_14214);
and UO_67 (O_67,N_14230,N_14984);
nand UO_68 (O_68,N_14957,N_14898);
xnor UO_69 (O_69,N_14300,N_14343);
nand UO_70 (O_70,N_14171,N_14733);
xnor UO_71 (O_71,N_14935,N_14905);
or UO_72 (O_72,N_14446,N_14104);
xor UO_73 (O_73,N_14879,N_14775);
xnor UO_74 (O_74,N_14022,N_14211);
or UO_75 (O_75,N_14004,N_14029);
xor UO_76 (O_76,N_14645,N_14252);
xnor UO_77 (O_77,N_14515,N_14225);
nand UO_78 (O_78,N_14174,N_14287);
nand UO_79 (O_79,N_14198,N_14633);
and UO_80 (O_80,N_14279,N_14199);
xor UO_81 (O_81,N_14203,N_14833);
nor UO_82 (O_82,N_14497,N_14009);
nor UO_83 (O_83,N_14376,N_14500);
nand UO_84 (O_84,N_14662,N_14927);
xor UO_85 (O_85,N_14192,N_14412);
and UO_86 (O_86,N_14938,N_14768);
and UO_87 (O_87,N_14933,N_14297);
xor UO_88 (O_88,N_14920,N_14835);
nand UO_89 (O_89,N_14896,N_14894);
or UO_90 (O_90,N_14578,N_14363);
or UO_91 (O_91,N_14993,N_14782);
or UO_92 (O_92,N_14069,N_14963);
or UO_93 (O_93,N_14206,N_14843);
xor UO_94 (O_94,N_14367,N_14547);
xor UO_95 (O_95,N_14507,N_14526);
xnor UO_96 (O_96,N_14246,N_14949);
nand UO_97 (O_97,N_14538,N_14611);
xor UO_98 (O_98,N_14067,N_14461);
or UO_99 (O_99,N_14567,N_14426);
or UO_100 (O_100,N_14678,N_14871);
nor UO_101 (O_101,N_14387,N_14562);
and UO_102 (O_102,N_14637,N_14436);
or UO_103 (O_103,N_14906,N_14008);
nor UO_104 (O_104,N_14055,N_14015);
or UO_105 (O_105,N_14374,N_14394);
xor UO_106 (O_106,N_14196,N_14162);
and UO_107 (O_107,N_14208,N_14438);
nor UO_108 (O_108,N_14520,N_14703);
or UO_109 (O_109,N_14789,N_14473);
nand UO_110 (O_110,N_14760,N_14460);
nor UO_111 (O_111,N_14071,N_14911);
nor UO_112 (O_112,N_14179,N_14087);
xnor UO_113 (O_113,N_14298,N_14427);
xor UO_114 (O_114,N_14423,N_14654);
nor UO_115 (O_115,N_14869,N_14980);
and UO_116 (O_116,N_14143,N_14221);
nand UO_117 (O_117,N_14195,N_14590);
nor UO_118 (O_118,N_14589,N_14084);
xor UO_119 (O_119,N_14144,N_14779);
and UO_120 (O_120,N_14966,N_14372);
and UO_121 (O_121,N_14432,N_14377);
or UO_122 (O_122,N_14255,N_14135);
xnor UO_123 (O_123,N_14670,N_14328);
xor UO_124 (O_124,N_14105,N_14242);
nor UO_125 (O_125,N_14803,N_14116);
nand UO_126 (O_126,N_14934,N_14844);
nand UO_127 (O_127,N_14236,N_14728);
and UO_128 (O_128,N_14142,N_14459);
and UO_129 (O_129,N_14647,N_14849);
and UO_130 (O_130,N_14990,N_14577);
nand UO_131 (O_131,N_14337,N_14333);
nand UO_132 (O_132,N_14122,N_14806);
nor UO_133 (O_133,N_14615,N_14817);
nor UO_134 (O_134,N_14596,N_14604);
xnor UO_135 (O_135,N_14277,N_14617);
xor UO_136 (O_136,N_14006,N_14982);
nand UO_137 (O_137,N_14204,N_14402);
xor UO_138 (O_138,N_14441,N_14165);
xnor UO_139 (O_139,N_14667,N_14437);
and UO_140 (O_140,N_14262,N_14451);
nor UO_141 (O_141,N_14537,N_14076);
nand UO_142 (O_142,N_14244,N_14684);
xor UO_143 (O_143,N_14757,N_14219);
xnor UO_144 (O_144,N_14233,N_14770);
or UO_145 (O_145,N_14731,N_14341);
and UO_146 (O_146,N_14386,N_14447);
nand UO_147 (O_147,N_14482,N_14326);
nand UO_148 (O_148,N_14146,N_14876);
nand UO_149 (O_149,N_14293,N_14910);
nor UO_150 (O_150,N_14652,N_14780);
nand UO_151 (O_151,N_14677,N_14035);
xnor UO_152 (O_152,N_14640,N_14099);
or UO_153 (O_153,N_14065,N_14098);
or UO_154 (O_154,N_14764,N_14347);
or UO_155 (O_155,N_14315,N_14699);
and UO_156 (O_156,N_14820,N_14490);
nand UO_157 (O_157,N_14344,N_14290);
nor UO_158 (O_158,N_14420,N_14453);
nand UO_159 (O_159,N_14579,N_14433);
nor UO_160 (O_160,N_14117,N_14224);
nand UO_161 (O_161,N_14784,N_14965);
nand UO_162 (O_162,N_14607,N_14561);
and UO_163 (O_163,N_14318,N_14712);
or UO_164 (O_164,N_14646,N_14988);
and UO_165 (O_165,N_14163,N_14137);
nor UO_166 (O_166,N_14053,N_14724);
xnor UO_167 (O_167,N_14945,N_14083);
or UO_168 (O_168,N_14774,N_14593);
or UO_169 (O_169,N_14533,N_14392);
nor UO_170 (O_170,N_14691,N_14235);
and UO_171 (O_171,N_14469,N_14316);
nand UO_172 (O_172,N_14545,N_14751);
nor UO_173 (O_173,N_14860,N_14489);
nor UO_174 (O_174,N_14664,N_14483);
nor UO_175 (O_175,N_14810,N_14907);
xnor UO_176 (O_176,N_14528,N_14886);
nor UO_177 (O_177,N_14892,N_14061);
xnor UO_178 (O_178,N_14422,N_14157);
and UO_179 (O_179,N_14696,N_14111);
nand UO_180 (O_180,N_14330,N_14606);
or UO_181 (O_181,N_14391,N_14003);
nand UO_182 (O_182,N_14253,N_14932);
and UO_183 (O_183,N_14384,N_14033);
or UO_184 (O_184,N_14812,N_14851);
nand UO_185 (O_185,N_14698,N_14176);
and UO_186 (O_186,N_14566,N_14090);
or UO_187 (O_187,N_14958,N_14028);
and UO_188 (O_188,N_14913,N_14946);
nand UO_189 (O_189,N_14686,N_14431);
or UO_190 (O_190,N_14824,N_14240);
or UO_191 (O_191,N_14057,N_14388);
xor UO_192 (O_192,N_14612,N_14857);
or UO_193 (O_193,N_14947,N_14799);
nor UO_194 (O_194,N_14185,N_14419);
nor UO_195 (O_195,N_14666,N_14216);
xor UO_196 (O_196,N_14925,N_14929);
or UO_197 (O_197,N_14583,N_14263);
xor UO_198 (O_198,N_14622,N_14322);
or UO_199 (O_199,N_14160,N_14471);
nor UO_200 (O_200,N_14997,N_14866);
and UO_201 (O_201,N_14406,N_14331);
nand UO_202 (O_202,N_14075,N_14480);
and UO_203 (O_203,N_14428,N_14762);
or UO_204 (O_204,N_14269,N_14854);
nand UO_205 (O_205,N_14074,N_14417);
xor UO_206 (O_206,N_14811,N_14280);
and UO_207 (O_207,N_14070,N_14656);
nand UO_208 (O_208,N_14804,N_14704);
nand UO_209 (O_209,N_14746,N_14822);
nor UO_210 (O_210,N_14251,N_14202);
nor UO_211 (O_211,N_14785,N_14641);
or UO_212 (O_212,N_14418,N_14150);
nor UO_213 (O_213,N_14271,N_14890);
nor UO_214 (O_214,N_14683,N_14969);
xnor UO_215 (O_215,N_14772,N_14828);
and UO_216 (O_216,N_14675,N_14254);
or UO_217 (O_217,N_14295,N_14080);
nor UO_218 (O_218,N_14685,N_14865);
nor UO_219 (O_219,N_14791,N_14005);
or UO_220 (O_220,N_14398,N_14636);
xnor UO_221 (O_221,N_14034,N_14819);
nand UO_222 (O_222,N_14158,N_14056);
or UO_223 (O_223,N_14575,N_14858);
nand UO_224 (O_224,N_14564,N_14701);
and UO_225 (O_225,N_14540,N_14976);
xor UO_226 (O_226,N_14207,N_14016);
xnor UO_227 (O_227,N_14989,N_14706);
xnor UO_228 (O_228,N_14353,N_14831);
nand UO_229 (O_229,N_14868,N_14899);
or UO_230 (O_230,N_14542,N_14802);
nand UO_231 (O_231,N_14546,N_14960);
nand UO_232 (O_232,N_14319,N_14123);
and UO_233 (O_233,N_14465,N_14335);
nand UO_234 (O_234,N_14501,N_14525);
xnor UO_235 (O_235,N_14442,N_14152);
nor UO_236 (O_236,N_14234,N_14634);
or UO_237 (O_237,N_14897,N_14610);
nand UO_238 (O_238,N_14715,N_14272);
nand UO_239 (O_239,N_14608,N_14628);
nand UO_240 (O_240,N_14729,N_14175);
nand UO_241 (O_241,N_14410,N_14977);
or UO_242 (O_242,N_14345,N_14320);
nand UO_243 (O_243,N_14411,N_14464);
and UO_244 (O_244,N_14115,N_14400);
nor UO_245 (O_245,N_14516,N_14304);
nand UO_246 (O_246,N_14642,N_14814);
xnor UO_247 (O_247,N_14895,N_14916);
nor UO_248 (O_248,N_14635,N_14643);
and UO_249 (O_249,N_14481,N_14616);
and UO_250 (O_250,N_14149,N_14747);
nor UO_251 (O_251,N_14031,N_14855);
nand UO_252 (O_252,N_14021,N_14166);
nor UO_253 (O_253,N_14275,N_14217);
nor UO_254 (O_254,N_14870,N_14605);
nor UO_255 (O_255,N_14191,N_14995);
xnor UO_256 (O_256,N_14761,N_14474);
nor UO_257 (O_257,N_14334,N_14439);
nor UO_258 (O_258,N_14514,N_14790);
nor UO_259 (O_259,N_14917,N_14559);
nor UO_260 (O_260,N_14783,N_14286);
nand UO_261 (O_261,N_14639,N_14010);
and UO_262 (O_262,N_14181,N_14188);
xnor UO_263 (O_263,N_14915,N_14161);
nand UO_264 (O_264,N_14725,N_14301);
nand UO_265 (O_265,N_14024,N_14587);
nand UO_266 (O_266,N_14908,N_14223);
nor UO_267 (O_267,N_14558,N_14393);
and UO_268 (O_268,N_14726,N_14338);
nor UO_269 (O_269,N_14722,N_14758);
or UO_270 (O_270,N_14765,N_14073);
and UO_271 (O_271,N_14818,N_14970);
nor UO_272 (O_272,N_14450,N_14794);
nor UO_273 (O_273,N_14707,N_14180);
nor UO_274 (O_274,N_14600,N_14778);
nand UO_275 (O_275,N_14928,N_14060);
or UO_276 (O_276,N_14270,N_14133);
or UO_277 (O_277,N_14522,N_14498);
or UO_278 (O_278,N_14151,N_14883);
xnor UO_279 (O_279,N_14630,N_14457);
nand UO_280 (O_280,N_14541,N_14661);
nor UO_281 (O_281,N_14443,N_14914);
and UO_282 (O_282,N_14364,N_14992);
or UO_283 (O_283,N_14329,N_14827);
xor UO_284 (O_284,N_14213,N_14186);
and UO_285 (O_285,N_14987,N_14257);
and UO_286 (O_286,N_14680,N_14332);
nand UO_287 (O_287,N_14172,N_14570);
and UO_288 (O_288,N_14107,N_14421);
nor UO_289 (O_289,N_14226,N_14554);
nor UO_290 (O_290,N_14648,N_14366);
or UO_291 (O_291,N_14125,N_14106);
nor UO_292 (O_292,N_14815,N_14941);
and UO_293 (O_293,N_14807,N_14968);
and UO_294 (O_294,N_14495,N_14900);
and UO_295 (O_295,N_14026,N_14050);
and UO_296 (O_296,N_14245,N_14565);
or UO_297 (O_297,N_14695,N_14351);
xor UO_298 (O_298,N_14808,N_14536);
nor UO_299 (O_299,N_14237,N_14737);
and UO_300 (O_300,N_14921,N_14739);
or UO_301 (O_301,N_14139,N_14205);
or UO_302 (O_302,N_14700,N_14754);
xnor UO_303 (O_303,N_14379,N_14499);
and UO_304 (O_304,N_14961,N_14413);
nand UO_305 (O_305,N_14569,N_14864);
nor UO_306 (O_306,N_14720,N_14342);
nand UO_307 (O_307,N_14058,N_14092);
nor UO_308 (O_308,N_14472,N_14742);
nand UO_309 (O_309,N_14355,N_14170);
and UO_310 (O_310,N_14629,N_14852);
nor UO_311 (O_311,N_14625,N_14042);
and UO_312 (O_312,N_14002,N_14874);
and UO_313 (O_313,N_14132,N_14278);
nand UO_314 (O_314,N_14266,N_14429);
or UO_315 (O_315,N_14983,N_14882);
nor UO_316 (O_316,N_14902,N_14138);
nor UO_317 (O_317,N_14357,N_14796);
xor UO_318 (O_318,N_14148,N_14430);
xor UO_319 (O_319,N_14717,N_14781);
xor UO_320 (O_320,N_14047,N_14951);
xor UO_321 (O_321,N_14672,N_14508);
or UO_322 (O_322,N_14488,N_14510);
nand UO_323 (O_323,N_14378,N_14749);
or UO_324 (O_324,N_14557,N_14349);
nor UO_325 (O_325,N_14544,N_14030);
nor UO_326 (O_326,N_14014,N_14981);
xnor UO_327 (O_327,N_14502,N_14734);
nand UO_328 (O_328,N_14763,N_14840);
nor UO_329 (O_329,N_14738,N_14626);
or UO_330 (O_330,N_14190,N_14644);
nand UO_331 (O_331,N_14127,N_14039);
and UO_332 (O_332,N_14311,N_14591);
xnor UO_333 (O_333,N_14036,N_14848);
and UO_334 (O_334,N_14543,N_14573);
xnor UO_335 (O_335,N_14651,N_14032);
nand UO_336 (O_336,N_14693,N_14267);
xor UO_337 (O_337,N_14620,N_14052);
xnor UO_338 (O_338,N_14584,N_14173);
nand UO_339 (O_339,N_14702,N_14942);
or UO_340 (O_340,N_14985,N_14100);
nand UO_341 (O_341,N_14850,N_14909);
and UO_342 (O_342,N_14873,N_14129);
and UO_343 (O_343,N_14455,N_14201);
nor UO_344 (O_344,N_14358,N_14931);
and UO_345 (O_345,N_14926,N_14404);
xnor UO_346 (O_346,N_14187,N_14091);
or UO_347 (O_347,N_14614,N_14486);
or UO_348 (O_348,N_14974,N_14215);
nand UO_349 (O_349,N_14792,N_14093);
and UO_350 (O_350,N_14200,N_14505);
or UO_351 (O_351,N_14339,N_14888);
xnor UO_352 (O_352,N_14813,N_14889);
or UO_353 (O_353,N_14618,N_14861);
nand UO_354 (O_354,N_14708,N_14830);
and UO_355 (O_355,N_14081,N_14736);
xor UO_356 (O_356,N_14735,N_14797);
xor UO_357 (O_357,N_14408,N_14924);
or UO_358 (O_358,N_14994,N_14518);
nor UO_359 (O_359,N_14283,N_14321);
and UO_360 (O_360,N_14177,N_14409);
or UO_361 (O_361,N_14110,N_14424);
nor UO_362 (O_362,N_14383,N_14602);
nor UO_363 (O_363,N_14572,N_14979);
nand UO_364 (O_364,N_14011,N_14798);
nor UO_365 (O_365,N_14496,N_14939);
xor UO_366 (O_366,N_14595,N_14197);
and UO_367 (O_367,N_14284,N_14078);
xnor UO_368 (O_368,N_14189,N_14524);
xnor UO_369 (O_369,N_14294,N_14041);
nand UO_370 (O_370,N_14923,N_14671);
and UO_371 (O_371,N_14303,N_14534);
xnor UO_372 (O_372,N_14755,N_14212);
nand UO_373 (O_373,N_14592,N_14013);
xnor UO_374 (O_374,N_14470,N_14445);
xor UO_375 (O_375,N_14973,N_14478);
and UO_376 (O_376,N_14660,N_14891);
xor UO_377 (O_377,N_14689,N_14773);
xor UO_378 (O_378,N_14227,N_14493);
or UO_379 (O_379,N_14837,N_14463);
or UO_380 (O_380,N_14930,N_14282);
or UO_381 (O_381,N_14743,N_14856);
nor UO_382 (O_382,N_14658,N_14360);
nand UO_383 (O_383,N_14448,N_14556);
or UO_384 (O_384,N_14832,N_14609);
or UO_385 (O_385,N_14887,N_14912);
or UO_386 (O_386,N_14694,N_14296);
or UO_387 (O_387,N_14962,N_14130);
nor UO_388 (O_388,N_14362,N_14741);
and UO_389 (O_389,N_14878,N_14085);
and UO_390 (O_390,N_14164,N_14373);
and UO_391 (O_391,N_14248,N_14504);
or UO_392 (O_392,N_14727,N_14485);
or UO_393 (O_393,N_14588,N_14668);
nand UO_394 (O_394,N_14239,N_14051);
nor UO_395 (O_395,N_14118,N_14709);
nand UO_396 (O_396,N_14399,N_14456);
and UO_397 (O_397,N_14901,N_14649);
or UO_398 (O_398,N_14681,N_14167);
nor UO_399 (O_399,N_14323,N_14291);
nand UO_400 (O_400,N_14222,N_14241);
and UO_401 (O_401,N_14952,N_14954);
xor UO_402 (O_402,N_14210,N_14314);
nand UO_403 (O_403,N_14354,N_14390);
xnor UO_404 (O_404,N_14062,N_14655);
xnor UO_405 (O_405,N_14816,N_14452);
or UO_406 (O_406,N_14603,N_14168);
nand UO_407 (O_407,N_14147,N_14317);
nand UO_408 (O_408,N_14312,N_14370);
nand UO_409 (O_409,N_14829,N_14692);
xnor UO_410 (O_410,N_14826,N_14585);
and UO_411 (O_411,N_14068,N_14308);
or UO_412 (O_412,N_14795,N_14853);
and UO_413 (O_413,N_14119,N_14444);
or UO_414 (O_414,N_14102,N_14079);
nand UO_415 (O_415,N_14801,N_14356);
nor UO_416 (O_416,N_14964,N_14719);
nand UO_417 (O_417,N_14000,N_14884);
nand UO_418 (O_418,N_14484,N_14825);
nor UO_419 (O_419,N_14121,N_14285);
nand UO_420 (O_420,N_14624,N_14903);
or UO_421 (O_421,N_14838,N_14972);
nor UO_422 (O_422,N_14359,N_14936);
nor UO_423 (O_423,N_14274,N_14155);
nand UO_424 (O_424,N_14243,N_14046);
xor UO_425 (O_425,N_14998,N_14893);
nand UO_426 (O_426,N_14040,N_14955);
nand UO_427 (O_427,N_14415,N_14732);
nor UO_428 (O_428,N_14950,N_14467);
or UO_429 (O_429,N_14017,N_14136);
and UO_430 (O_430,N_14109,N_14809);
xor UO_431 (O_431,N_14477,N_14956);
nor UO_432 (O_432,N_14967,N_14821);
xnor UO_433 (O_433,N_14697,N_14305);
or UO_434 (O_434,N_14260,N_14512);
and UO_435 (O_435,N_14613,N_14513);
nor UO_436 (O_436,N_14247,N_14881);
nand UO_437 (O_437,N_14340,N_14114);
nand UO_438 (O_438,N_14531,N_14183);
nand UO_439 (O_439,N_14996,N_14141);
nor UO_440 (O_440,N_14025,N_14563);
and UO_441 (O_441,N_14238,N_14361);
and UO_442 (O_442,N_14218,N_14193);
nor UO_443 (O_443,N_14299,N_14548);
nor UO_444 (O_444,N_14788,N_14601);
nand UO_445 (O_445,N_14302,N_14723);
or UO_446 (O_446,N_14687,N_14407);
and UO_447 (O_447,N_14978,N_14638);
nor UO_448 (O_448,N_14095,N_14919);
or UO_449 (O_449,N_14549,N_14479);
or UO_450 (O_450,N_14552,N_14156);
and UO_451 (O_451,N_14750,N_14476);
xnor UO_452 (O_452,N_14506,N_14503);
xnor UO_453 (O_453,N_14309,N_14519);
nand UO_454 (O_454,N_14509,N_14348);
and UO_455 (O_455,N_14530,N_14834);
or UO_456 (O_456,N_14043,N_14713);
xnor UO_457 (O_457,N_14140,N_14194);
xor UO_458 (O_458,N_14229,N_14097);
nor UO_459 (O_459,N_14475,N_14576);
nand UO_460 (O_460,N_14676,N_14066);
nor UO_461 (O_461,N_14020,N_14535);
and UO_462 (O_462,N_14527,N_14064);
nand UO_463 (O_463,N_14159,N_14748);
xor UO_464 (O_464,N_14845,N_14597);
or UO_465 (O_465,N_14259,N_14711);
nor UO_466 (O_466,N_14089,N_14885);
and UO_467 (O_467,N_14027,N_14396);
nor UO_468 (O_468,N_14289,N_14767);
nor UO_469 (O_469,N_14371,N_14487);
or UO_470 (O_470,N_14249,N_14718);
nor UO_471 (O_471,N_14787,N_14999);
and UO_472 (O_472,N_14555,N_14458);
and UO_473 (O_473,N_14657,N_14650);
and UO_474 (O_474,N_14653,N_14220);
or UO_475 (O_475,N_14112,N_14325);
or UO_476 (O_476,N_14045,N_14169);
or UO_477 (O_477,N_14368,N_14491);
nor UO_478 (O_478,N_14904,N_14532);
nand UO_479 (O_479,N_14454,N_14673);
nand UO_480 (O_480,N_14313,N_14551);
and UO_481 (O_481,N_14745,N_14753);
or UO_482 (O_482,N_14416,N_14877);
nand UO_483 (O_483,N_14943,N_14019);
xor UO_484 (O_484,N_14038,N_14088);
and UO_485 (O_485,N_14867,N_14663);
or UO_486 (O_486,N_14494,N_14492);
nor UO_487 (O_487,N_14154,N_14511);
nor UO_488 (O_488,N_14621,N_14134);
nand UO_489 (O_489,N_14523,N_14365);
nand UO_490 (O_490,N_14682,N_14619);
nor UO_491 (O_491,N_14705,N_14786);
nor UO_492 (O_492,N_14462,N_14397);
or UO_493 (O_493,N_14012,N_14769);
xor UO_494 (O_494,N_14862,N_14131);
nor UO_495 (O_495,N_14776,N_14922);
or UO_496 (O_496,N_14403,N_14044);
nor UO_497 (O_497,N_14101,N_14449);
or UO_498 (O_498,N_14327,N_14258);
xor UO_499 (O_499,N_14288,N_14310);
nor UO_500 (O_500,N_14123,N_14041);
or UO_501 (O_501,N_14387,N_14858);
xor UO_502 (O_502,N_14665,N_14459);
nand UO_503 (O_503,N_14413,N_14503);
nor UO_504 (O_504,N_14505,N_14892);
nand UO_505 (O_505,N_14631,N_14993);
nor UO_506 (O_506,N_14863,N_14509);
or UO_507 (O_507,N_14829,N_14146);
and UO_508 (O_508,N_14429,N_14146);
or UO_509 (O_509,N_14725,N_14768);
nand UO_510 (O_510,N_14197,N_14625);
nor UO_511 (O_511,N_14416,N_14125);
nor UO_512 (O_512,N_14457,N_14113);
xor UO_513 (O_513,N_14482,N_14719);
nor UO_514 (O_514,N_14876,N_14833);
and UO_515 (O_515,N_14481,N_14382);
and UO_516 (O_516,N_14516,N_14026);
nor UO_517 (O_517,N_14948,N_14833);
xnor UO_518 (O_518,N_14495,N_14241);
xor UO_519 (O_519,N_14355,N_14357);
xor UO_520 (O_520,N_14189,N_14856);
nor UO_521 (O_521,N_14262,N_14719);
xnor UO_522 (O_522,N_14052,N_14827);
nand UO_523 (O_523,N_14528,N_14223);
nand UO_524 (O_524,N_14596,N_14372);
nand UO_525 (O_525,N_14513,N_14786);
nor UO_526 (O_526,N_14491,N_14094);
and UO_527 (O_527,N_14801,N_14496);
or UO_528 (O_528,N_14487,N_14621);
or UO_529 (O_529,N_14558,N_14482);
nor UO_530 (O_530,N_14088,N_14684);
or UO_531 (O_531,N_14781,N_14544);
or UO_532 (O_532,N_14680,N_14296);
xor UO_533 (O_533,N_14357,N_14294);
nand UO_534 (O_534,N_14142,N_14212);
and UO_535 (O_535,N_14614,N_14385);
nor UO_536 (O_536,N_14362,N_14606);
nand UO_537 (O_537,N_14273,N_14617);
nor UO_538 (O_538,N_14794,N_14392);
nand UO_539 (O_539,N_14919,N_14391);
xor UO_540 (O_540,N_14562,N_14782);
and UO_541 (O_541,N_14097,N_14324);
nand UO_542 (O_542,N_14204,N_14500);
and UO_543 (O_543,N_14615,N_14386);
nor UO_544 (O_544,N_14440,N_14587);
or UO_545 (O_545,N_14959,N_14199);
and UO_546 (O_546,N_14498,N_14152);
or UO_547 (O_547,N_14930,N_14529);
nor UO_548 (O_548,N_14265,N_14495);
xor UO_549 (O_549,N_14764,N_14369);
nand UO_550 (O_550,N_14399,N_14222);
nor UO_551 (O_551,N_14589,N_14774);
xnor UO_552 (O_552,N_14229,N_14429);
or UO_553 (O_553,N_14587,N_14398);
nor UO_554 (O_554,N_14273,N_14282);
or UO_555 (O_555,N_14243,N_14327);
and UO_556 (O_556,N_14292,N_14848);
nor UO_557 (O_557,N_14734,N_14499);
or UO_558 (O_558,N_14906,N_14104);
or UO_559 (O_559,N_14868,N_14509);
nand UO_560 (O_560,N_14209,N_14232);
nor UO_561 (O_561,N_14167,N_14906);
xnor UO_562 (O_562,N_14469,N_14738);
and UO_563 (O_563,N_14756,N_14733);
or UO_564 (O_564,N_14204,N_14358);
xnor UO_565 (O_565,N_14616,N_14499);
nor UO_566 (O_566,N_14688,N_14286);
xnor UO_567 (O_567,N_14947,N_14761);
xor UO_568 (O_568,N_14040,N_14847);
or UO_569 (O_569,N_14886,N_14242);
or UO_570 (O_570,N_14283,N_14349);
or UO_571 (O_571,N_14922,N_14862);
or UO_572 (O_572,N_14385,N_14503);
nand UO_573 (O_573,N_14567,N_14142);
xor UO_574 (O_574,N_14406,N_14449);
or UO_575 (O_575,N_14592,N_14668);
or UO_576 (O_576,N_14712,N_14718);
xor UO_577 (O_577,N_14046,N_14726);
nor UO_578 (O_578,N_14965,N_14365);
and UO_579 (O_579,N_14364,N_14145);
and UO_580 (O_580,N_14121,N_14275);
xor UO_581 (O_581,N_14137,N_14495);
nor UO_582 (O_582,N_14867,N_14456);
nand UO_583 (O_583,N_14319,N_14370);
or UO_584 (O_584,N_14598,N_14290);
nand UO_585 (O_585,N_14769,N_14255);
nand UO_586 (O_586,N_14043,N_14894);
nor UO_587 (O_587,N_14691,N_14834);
and UO_588 (O_588,N_14286,N_14795);
or UO_589 (O_589,N_14625,N_14118);
and UO_590 (O_590,N_14638,N_14121);
and UO_591 (O_591,N_14593,N_14993);
nand UO_592 (O_592,N_14900,N_14496);
and UO_593 (O_593,N_14625,N_14423);
nor UO_594 (O_594,N_14749,N_14472);
and UO_595 (O_595,N_14990,N_14510);
nand UO_596 (O_596,N_14852,N_14443);
xnor UO_597 (O_597,N_14570,N_14395);
nand UO_598 (O_598,N_14806,N_14039);
nand UO_599 (O_599,N_14952,N_14349);
and UO_600 (O_600,N_14835,N_14741);
or UO_601 (O_601,N_14434,N_14388);
nor UO_602 (O_602,N_14269,N_14242);
and UO_603 (O_603,N_14990,N_14908);
nor UO_604 (O_604,N_14737,N_14949);
or UO_605 (O_605,N_14994,N_14783);
or UO_606 (O_606,N_14111,N_14646);
nand UO_607 (O_607,N_14077,N_14054);
or UO_608 (O_608,N_14685,N_14673);
xor UO_609 (O_609,N_14839,N_14802);
and UO_610 (O_610,N_14048,N_14519);
and UO_611 (O_611,N_14542,N_14598);
nand UO_612 (O_612,N_14943,N_14594);
and UO_613 (O_613,N_14218,N_14591);
xnor UO_614 (O_614,N_14659,N_14566);
or UO_615 (O_615,N_14579,N_14068);
nor UO_616 (O_616,N_14739,N_14139);
or UO_617 (O_617,N_14615,N_14787);
xor UO_618 (O_618,N_14856,N_14530);
or UO_619 (O_619,N_14514,N_14644);
or UO_620 (O_620,N_14048,N_14429);
and UO_621 (O_621,N_14847,N_14450);
and UO_622 (O_622,N_14762,N_14366);
and UO_623 (O_623,N_14898,N_14689);
and UO_624 (O_624,N_14792,N_14707);
and UO_625 (O_625,N_14113,N_14091);
nand UO_626 (O_626,N_14015,N_14776);
xor UO_627 (O_627,N_14561,N_14117);
or UO_628 (O_628,N_14752,N_14189);
nor UO_629 (O_629,N_14564,N_14143);
nand UO_630 (O_630,N_14279,N_14106);
nor UO_631 (O_631,N_14761,N_14677);
xor UO_632 (O_632,N_14317,N_14518);
nand UO_633 (O_633,N_14821,N_14007);
or UO_634 (O_634,N_14174,N_14179);
or UO_635 (O_635,N_14393,N_14402);
nand UO_636 (O_636,N_14186,N_14079);
or UO_637 (O_637,N_14147,N_14441);
and UO_638 (O_638,N_14346,N_14924);
and UO_639 (O_639,N_14480,N_14931);
xor UO_640 (O_640,N_14244,N_14855);
nand UO_641 (O_641,N_14779,N_14594);
or UO_642 (O_642,N_14244,N_14374);
nor UO_643 (O_643,N_14397,N_14440);
and UO_644 (O_644,N_14710,N_14396);
or UO_645 (O_645,N_14964,N_14328);
nand UO_646 (O_646,N_14027,N_14182);
nor UO_647 (O_647,N_14275,N_14192);
and UO_648 (O_648,N_14383,N_14512);
nor UO_649 (O_649,N_14314,N_14707);
and UO_650 (O_650,N_14658,N_14182);
nand UO_651 (O_651,N_14576,N_14109);
nor UO_652 (O_652,N_14482,N_14674);
or UO_653 (O_653,N_14129,N_14237);
nor UO_654 (O_654,N_14936,N_14947);
nand UO_655 (O_655,N_14775,N_14436);
or UO_656 (O_656,N_14187,N_14524);
and UO_657 (O_657,N_14976,N_14185);
nand UO_658 (O_658,N_14749,N_14408);
nor UO_659 (O_659,N_14859,N_14281);
or UO_660 (O_660,N_14890,N_14620);
or UO_661 (O_661,N_14040,N_14894);
nand UO_662 (O_662,N_14438,N_14248);
nand UO_663 (O_663,N_14886,N_14125);
xnor UO_664 (O_664,N_14753,N_14979);
xor UO_665 (O_665,N_14403,N_14496);
and UO_666 (O_666,N_14011,N_14157);
xor UO_667 (O_667,N_14706,N_14086);
and UO_668 (O_668,N_14244,N_14108);
and UO_669 (O_669,N_14625,N_14387);
nor UO_670 (O_670,N_14107,N_14378);
and UO_671 (O_671,N_14141,N_14445);
nor UO_672 (O_672,N_14088,N_14968);
nand UO_673 (O_673,N_14295,N_14889);
nand UO_674 (O_674,N_14349,N_14599);
nor UO_675 (O_675,N_14267,N_14405);
and UO_676 (O_676,N_14859,N_14166);
xnor UO_677 (O_677,N_14765,N_14570);
and UO_678 (O_678,N_14008,N_14996);
or UO_679 (O_679,N_14556,N_14196);
and UO_680 (O_680,N_14628,N_14143);
nor UO_681 (O_681,N_14796,N_14784);
xor UO_682 (O_682,N_14148,N_14450);
nand UO_683 (O_683,N_14111,N_14324);
and UO_684 (O_684,N_14575,N_14200);
xor UO_685 (O_685,N_14339,N_14848);
nor UO_686 (O_686,N_14330,N_14627);
or UO_687 (O_687,N_14453,N_14334);
nor UO_688 (O_688,N_14951,N_14337);
or UO_689 (O_689,N_14571,N_14416);
and UO_690 (O_690,N_14064,N_14058);
and UO_691 (O_691,N_14296,N_14831);
nand UO_692 (O_692,N_14488,N_14104);
xnor UO_693 (O_693,N_14002,N_14118);
xor UO_694 (O_694,N_14222,N_14901);
and UO_695 (O_695,N_14481,N_14097);
and UO_696 (O_696,N_14771,N_14191);
and UO_697 (O_697,N_14698,N_14903);
and UO_698 (O_698,N_14017,N_14815);
and UO_699 (O_699,N_14785,N_14505);
nand UO_700 (O_700,N_14811,N_14829);
xnor UO_701 (O_701,N_14219,N_14856);
nand UO_702 (O_702,N_14301,N_14848);
or UO_703 (O_703,N_14557,N_14587);
and UO_704 (O_704,N_14567,N_14494);
or UO_705 (O_705,N_14213,N_14124);
nand UO_706 (O_706,N_14233,N_14789);
nor UO_707 (O_707,N_14225,N_14426);
nor UO_708 (O_708,N_14679,N_14701);
or UO_709 (O_709,N_14994,N_14174);
and UO_710 (O_710,N_14847,N_14741);
xor UO_711 (O_711,N_14449,N_14024);
or UO_712 (O_712,N_14869,N_14160);
xor UO_713 (O_713,N_14627,N_14811);
and UO_714 (O_714,N_14465,N_14861);
nand UO_715 (O_715,N_14544,N_14344);
nor UO_716 (O_716,N_14526,N_14261);
xor UO_717 (O_717,N_14893,N_14102);
nand UO_718 (O_718,N_14901,N_14473);
nor UO_719 (O_719,N_14439,N_14115);
xor UO_720 (O_720,N_14080,N_14704);
nand UO_721 (O_721,N_14247,N_14440);
nand UO_722 (O_722,N_14149,N_14506);
or UO_723 (O_723,N_14296,N_14144);
and UO_724 (O_724,N_14313,N_14260);
nand UO_725 (O_725,N_14456,N_14190);
xnor UO_726 (O_726,N_14804,N_14244);
and UO_727 (O_727,N_14669,N_14304);
nand UO_728 (O_728,N_14806,N_14652);
nand UO_729 (O_729,N_14900,N_14699);
xnor UO_730 (O_730,N_14868,N_14494);
nor UO_731 (O_731,N_14670,N_14485);
nand UO_732 (O_732,N_14467,N_14414);
and UO_733 (O_733,N_14825,N_14539);
or UO_734 (O_734,N_14533,N_14718);
xnor UO_735 (O_735,N_14651,N_14216);
and UO_736 (O_736,N_14031,N_14489);
or UO_737 (O_737,N_14033,N_14460);
nor UO_738 (O_738,N_14832,N_14439);
or UO_739 (O_739,N_14441,N_14507);
xor UO_740 (O_740,N_14709,N_14901);
nor UO_741 (O_741,N_14823,N_14743);
or UO_742 (O_742,N_14611,N_14466);
nor UO_743 (O_743,N_14843,N_14848);
and UO_744 (O_744,N_14866,N_14780);
xnor UO_745 (O_745,N_14668,N_14896);
xor UO_746 (O_746,N_14134,N_14865);
nor UO_747 (O_747,N_14737,N_14064);
nor UO_748 (O_748,N_14956,N_14643);
xor UO_749 (O_749,N_14811,N_14375);
nor UO_750 (O_750,N_14216,N_14877);
or UO_751 (O_751,N_14909,N_14726);
nor UO_752 (O_752,N_14295,N_14110);
nor UO_753 (O_753,N_14001,N_14183);
nand UO_754 (O_754,N_14650,N_14851);
and UO_755 (O_755,N_14681,N_14518);
xnor UO_756 (O_756,N_14434,N_14618);
and UO_757 (O_757,N_14587,N_14508);
nor UO_758 (O_758,N_14831,N_14721);
or UO_759 (O_759,N_14840,N_14743);
and UO_760 (O_760,N_14758,N_14275);
nand UO_761 (O_761,N_14634,N_14651);
or UO_762 (O_762,N_14186,N_14744);
nor UO_763 (O_763,N_14320,N_14774);
or UO_764 (O_764,N_14929,N_14135);
xnor UO_765 (O_765,N_14718,N_14911);
or UO_766 (O_766,N_14212,N_14583);
or UO_767 (O_767,N_14447,N_14367);
xor UO_768 (O_768,N_14182,N_14960);
xor UO_769 (O_769,N_14341,N_14516);
and UO_770 (O_770,N_14801,N_14900);
and UO_771 (O_771,N_14883,N_14837);
and UO_772 (O_772,N_14956,N_14831);
nand UO_773 (O_773,N_14205,N_14504);
or UO_774 (O_774,N_14826,N_14070);
or UO_775 (O_775,N_14619,N_14522);
and UO_776 (O_776,N_14219,N_14974);
and UO_777 (O_777,N_14980,N_14100);
nor UO_778 (O_778,N_14411,N_14489);
and UO_779 (O_779,N_14087,N_14705);
or UO_780 (O_780,N_14831,N_14119);
nand UO_781 (O_781,N_14482,N_14990);
xnor UO_782 (O_782,N_14019,N_14770);
or UO_783 (O_783,N_14510,N_14178);
nor UO_784 (O_784,N_14691,N_14360);
or UO_785 (O_785,N_14794,N_14692);
xor UO_786 (O_786,N_14630,N_14142);
nand UO_787 (O_787,N_14743,N_14634);
and UO_788 (O_788,N_14251,N_14785);
nand UO_789 (O_789,N_14000,N_14439);
nand UO_790 (O_790,N_14313,N_14991);
or UO_791 (O_791,N_14102,N_14542);
xor UO_792 (O_792,N_14463,N_14623);
nand UO_793 (O_793,N_14525,N_14999);
xor UO_794 (O_794,N_14088,N_14473);
xor UO_795 (O_795,N_14820,N_14435);
nor UO_796 (O_796,N_14789,N_14783);
xor UO_797 (O_797,N_14015,N_14207);
and UO_798 (O_798,N_14180,N_14717);
or UO_799 (O_799,N_14851,N_14335);
and UO_800 (O_800,N_14564,N_14444);
nand UO_801 (O_801,N_14604,N_14630);
xor UO_802 (O_802,N_14381,N_14782);
or UO_803 (O_803,N_14865,N_14618);
nand UO_804 (O_804,N_14270,N_14748);
and UO_805 (O_805,N_14589,N_14795);
or UO_806 (O_806,N_14729,N_14104);
nor UO_807 (O_807,N_14854,N_14793);
xor UO_808 (O_808,N_14014,N_14630);
xor UO_809 (O_809,N_14323,N_14792);
nand UO_810 (O_810,N_14965,N_14964);
nand UO_811 (O_811,N_14969,N_14263);
xnor UO_812 (O_812,N_14828,N_14260);
or UO_813 (O_813,N_14327,N_14201);
xor UO_814 (O_814,N_14192,N_14768);
nor UO_815 (O_815,N_14189,N_14630);
and UO_816 (O_816,N_14006,N_14952);
and UO_817 (O_817,N_14488,N_14871);
xor UO_818 (O_818,N_14263,N_14170);
and UO_819 (O_819,N_14217,N_14746);
xor UO_820 (O_820,N_14881,N_14400);
xor UO_821 (O_821,N_14028,N_14124);
xnor UO_822 (O_822,N_14652,N_14986);
nand UO_823 (O_823,N_14450,N_14912);
nor UO_824 (O_824,N_14027,N_14732);
xor UO_825 (O_825,N_14256,N_14608);
nor UO_826 (O_826,N_14744,N_14842);
nand UO_827 (O_827,N_14453,N_14739);
xor UO_828 (O_828,N_14803,N_14635);
xnor UO_829 (O_829,N_14535,N_14956);
xor UO_830 (O_830,N_14347,N_14211);
xor UO_831 (O_831,N_14908,N_14896);
or UO_832 (O_832,N_14408,N_14065);
nand UO_833 (O_833,N_14982,N_14677);
nor UO_834 (O_834,N_14374,N_14005);
and UO_835 (O_835,N_14203,N_14305);
nand UO_836 (O_836,N_14691,N_14130);
or UO_837 (O_837,N_14323,N_14096);
nor UO_838 (O_838,N_14760,N_14621);
and UO_839 (O_839,N_14984,N_14736);
xnor UO_840 (O_840,N_14961,N_14688);
nand UO_841 (O_841,N_14621,N_14888);
or UO_842 (O_842,N_14030,N_14875);
nor UO_843 (O_843,N_14770,N_14350);
nor UO_844 (O_844,N_14245,N_14980);
nand UO_845 (O_845,N_14388,N_14730);
nor UO_846 (O_846,N_14164,N_14206);
xor UO_847 (O_847,N_14192,N_14290);
nor UO_848 (O_848,N_14376,N_14227);
nor UO_849 (O_849,N_14736,N_14640);
or UO_850 (O_850,N_14808,N_14581);
or UO_851 (O_851,N_14649,N_14605);
nor UO_852 (O_852,N_14534,N_14158);
nand UO_853 (O_853,N_14374,N_14727);
nand UO_854 (O_854,N_14420,N_14805);
xnor UO_855 (O_855,N_14304,N_14488);
and UO_856 (O_856,N_14667,N_14492);
nor UO_857 (O_857,N_14629,N_14802);
and UO_858 (O_858,N_14203,N_14434);
nor UO_859 (O_859,N_14504,N_14105);
and UO_860 (O_860,N_14504,N_14119);
or UO_861 (O_861,N_14836,N_14110);
or UO_862 (O_862,N_14310,N_14512);
or UO_863 (O_863,N_14894,N_14041);
xor UO_864 (O_864,N_14945,N_14066);
or UO_865 (O_865,N_14015,N_14222);
or UO_866 (O_866,N_14271,N_14687);
and UO_867 (O_867,N_14482,N_14522);
and UO_868 (O_868,N_14744,N_14080);
or UO_869 (O_869,N_14335,N_14010);
or UO_870 (O_870,N_14041,N_14762);
nand UO_871 (O_871,N_14541,N_14935);
nand UO_872 (O_872,N_14193,N_14342);
nor UO_873 (O_873,N_14019,N_14580);
nor UO_874 (O_874,N_14689,N_14374);
nor UO_875 (O_875,N_14315,N_14221);
xor UO_876 (O_876,N_14382,N_14734);
and UO_877 (O_877,N_14267,N_14962);
and UO_878 (O_878,N_14688,N_14288);
nor UO_879 (O_879,N_14247,N_14319);
nor UO_880 (O_880,N_14709,N_14085);
nand UO_881 (O_881,N_14240,N_14091);
nand UO_882 (O_882,N_14746,N_14814);
nand UO_883 (O_883,N_14611,N_14200);
nand UO_884 (O_884,N_14144,N_14994);
nand UO_885 (O_885,N_14471,N_14679);
nand UO_886 (O_886,N_14618,N_14483);
xor UO_887 (O_887,N_14326,N_14345);
and UO_888 (O_888,N_14426,N_14540);
nand UO_889 (O_889,N_14178,N_14229);
nand UO_890 (O_890,N_14025,N_14949);
nor UO_891 (O_891,N_14564,N_14706);
xnor UO_892 (O_892,N_14219,N_14353);
or UO_893 (O_893,N_14283,N_14570);
xnor UO_894 (O_894,N_14313,N_14907);
nor UO_895 (O_895,N_14677,N_14048);
xor UO_896 (O_896,N_14500,N_14073);
nor UO_897 (O_897,N_14925,N_14357);
xnor UO_898 (O_898,N_14051,N_14237);
nand UO_899 (O_899,N_14713,N_14333);
xnor UO_900 (O_900,N_14917,N_14732);
nand UO_901 (O_901,N_14216,N_14168);
nor UO_902 (O_902,N_14330,N_14112);
xor UO_903 (O_903,N_14934,N_14105);
xnor UO_904 (O_904,N_14056,N_14968);
nor UO_905 (O_905,N_14235,N_14837);
or UO_906 (O_906,N_14242,N_14312);
nand UO_907 (O_907,N_14739,N_14876);
or UO_908 (O_908,N_14734,N_14946);
nor UO_909 (O_909,N_14194,N_14221);
and UO_910 (O_910,N_14512,N_14117);
or UO_911 (O_911,N_14187,N_14148);
or UO_912 (O_912,N_14237,N_14325);
or UO_913 (O_913,N_14950,N_14778);
or UO_914 (O_914,N_14146,N_14505);
xnor UO_915 (O_915,N_14493,N_14854);
and UO_916 (O_916,N_14698,N_14929);
and UO_917 (O_917,N_14417,N_14920);
nor UO_918 (O_918,N_14887,N_14846);
nand UO_919 (O_919,N_14685,N_14011);
and UO_920 (O_920,N_14649,N_14066);
xor UO_921 (O_921,N_14475,N_14372);
nor UO_922 (O_922,N_14777,N_14700);
and UO_923 (O_923,N_14704,N_14637);
nand UO_924 (O_924,N_14152,N_14344);
nor UO_925 (O_925,N_14288,N_14637);
xnor UO_926 (O_926,N_14997,N_14680);
or UO_927 (O_927,N_14304,N_14210);
and UO_928 (O_928,N_14525,N_14207);
xnor UO_929 (O_929,N_14624,N_14288);
and UO_930 (O_930,N_14728,N_14362);
and UO_931 (O_931,N_14017,N_14857);
nor UO_932 (O_932,N_14783,N_14705);
xnor UO_933 (O_933,N_14563,N_14318);
and UO_934 (O_934,N_14124,N_14544);
or UO_935 (O_935,N_14807,N_14021);
or UO_936 (O_936,N_14958,N_14781);
nor UO_937 (O_937,N_14506,N_14421);
nor UO_938 (O_938,N_14957,N_14004);
nor UO_939 (O_939,N_14459,N_14427);
nor UO_940 (O_940,N_14976,N_14814);
nand UO_941 (O_941,N_14235,N_14463);
xnor UO_942 (O_942,N_14333,N_14320);
and UO_943 (O_943,N_14034,N_14793);
or UO_944 (O_944,N_14145,N_14691);
and UO_945 (O_945,N_14166,N_14989);
xor UO_946 (O_946,N_14514,N_14433);
xor UO_947 (O_947,N_14223,N_14982);
nand UO_948 (O_948,N_14782,N_14333);
or UO_949 (O_949,N_14964,N_14060);
or UO_950 (O_950,N_14660,N_14307);
and UO_951 (O_951,N_14983,N_14830);
and UO_952 (O_952,N_14845,N_14919);
or UO_953 (O_953,N_14618,N_14262);
xnor UO_954 (O_954,N_14265,N_14304);
xor UO_955 (O_955,N_14080,N_14479);
or UO_956 (O_956,N_14300,N_14737);
xnor UO_957 (O_957,N_14994,N_14549);
and UO_958 (O_958,N_14660,N_14838);
xnor UO_959 (O_959,N_14282,N_14559);
nand UO_960 (O_960,N_14898,N_14040);
xor UO_961 (O_961,N_14870,N_14433);
and UO_962 (O_962,N_14644,N_14958);
xor UO_963 (O_963,N_14586,N_14655);
nor UO_964 (O_964,N_14540,N_14353);
or UO_965 (O_965,N_14746,N_14197);
nand UO_966 (O_966,N_14137,N_14741);
and UO_967 (O_967,N_14378,N_14083);
nor UO_968 (O_968,N_14259,N_14900);
xor UO_969 (O_969,N_14378,N_14218);
nor UO_970 (O_970,N_14474,N_14274);
or UO_971 (O_971,N_14717,N_14049);
nor UO_972 (O_972,N_14491,N_14294);
and UO_973 (O_973,N_14640,N_14437);
nor UO_974 (O_974,N_14719,N_14847);
and UO_975 (O_975,N_14496,N_14290);
or UO_976 (O_976,N_14882,N_14588);
or UO_977 (O_977,N_14037,N_14184);
nor UO_978 (O_978,N_14425,N_14748);
or UO_979 (O_979,N_14337,N_14990);
nand UO_980 (O_980,N_14576,N_14738);
nand UO_981 (O_981,N_14892,N_14458);
nor UO_982 (O_982,N_14874,N_14109);
nand UO_983 (O_983,N_14846,N_14651);
nor UO_984 (O_984,N_14751,N_14244);
nand UO_985 (O_985,N_14583,N_14177);
or UO_986 (O_986,N_14787,N_14472);
xor UO_987 (O_987,N_14089,N_14641);
xor UO_988 (O_988,N_14073,N_14587);
nand UO_989 (O_989,N_14344,N_14924);
nand UO_990 (O_990,N_14045,N_14352);
and UO_991 (O_991,N_14340,N_14344);
or UO_992 (O_992,N_14400,N_14549);
xor UO_993 (O_993,N_14281,N_14101);
nor UO_994 (O_994,N_14140,N_14314);
xnor UO_995 (O_995,N_14311,N_14945);
or UO_996 (O_996,N_14027,N_14595);
xor UO_997 (O_997,N_14704,N_14352);
nor UO_998 (O_998,N_14572,N_14276);
or UO_999 (O_999,N_14978,N_14285);
nor UO_1000 (O_1000,N_14710,N_14408);
and UO_1001 (O_1001,N_14610,N_14052);
nand UO_1002 (O_1002,N_14122,N_14706);
nor UO_1003 (O_1003,N_14378,N_14356);
or UO_1004 (O_1004,N_14876,N_14440);
and UO_1005 (O_1005,N_14397,N_14583);
and UO_1006 (O_1006,N_14634,N_14707);
or UO_1007 (O_1007,N_14907,N_14325);
nand UO_1008 (O_1008,N_14012,N_14752);
xor UO_1009 (O_1009,N_14317,N_14535);
nor UO_1010 (O_1010,N_14588,N_14727);
xnor UO_1011 (O_1011,N_14377,N_14162);
and UO_1012 (O_1012,N_14113,N_14284);
or UO_1013 (O_1013,N_14299,N_14217);
nor UO_1014 (O_1014,N_14028,N_14312);
or UO_1015 (O_1015,N_14389,N_14427);
nand UO_1016 (O_1016,N_14594,N_14955);
nand UO_1017 (O_1017,N_14649,N_14520);
nand UO_1018 (O_1018,N_14837,N_14590);
or UO_1019 (O_1019,N_14598,N_14637);
and UO_1020 (O_1020,N_14003,N_14295);
or UO_1021 (O_1021,N_14551,N_14397);
or UO_1022 (O_1022,N_14949,N_14453);
and UO_1023 (O_1023,N_14458,N_14103);
xnor UO_1024 (O_1024,N_14216,N_14823);
and UO_1025 (O_1025,N_14964,N_14821);
nor UO_1026 (O_1026,N_14979,N_14606);
xnor UO_1027 (O_1027,N_14807,N_14210);
nand UO_1028 (O_1028,N_14323,N_14581);
or UO_1029 (O_1029,N_14257,N_14255);
or UO_1030 (O_1030,N_14443,N_14469);
or UO_1031 (O_1031,N_14129,N_14756);
xor UO_1032 (O_1032,N_14007,N_14345);
nand UO_1033 (O_1033,N_14745,N_14989);
nor UO_1034 (O_1034,N_14958,N_14304);
and UO_1035 (O_1035,N_14143,N_14684);
nor UO_1036 (O_1036,N_14313,N_14143);
or UO_1037 (O_1037,N_14541,N_14815);
or UO_1038 (O_1038,N_14720,N_14377);
and UO_1039 (O_1039,N_14299,N_14958);
nor UO_1040 (O_1040,N_14887,N_14521);
or UO_1041 (O_1041,N_14164,N_14934);
and UO_1042 (O_1042,N_14736,N_14202);
nand UO_1043 (O_1043,N_14549,N_14398);
nor UO_1044 (O_1044,N_14511,N_14077);
and UO_1045 (O_1045,N_14645,N_14363);
and UO_1046 (O_1046,N_14266,N_14640);
nand UO_1047 (O_1047,N_14322,N_14004);
and UO_1048 (O_1048,N_14999,N_14478);
nor UO_1049 (O_1049,N_14614,N_14867);
and UO_1050 (O_1050,N_14621,N_14908);
xor UO_1051 (O_1051,N_14763,N_14145);
and UO_1052 (O_1052,N_14132,N_14291);
nand UO_1053 (O_1053,N_14149,N_14378);
xor UO_1054 (O_1054,N_14636,N_14521);
nor UO_1055 (O_1055,N_14498,N_14863);
and UO_1056 (O_1056,N_14831,N_14135);
and UO_1057 (O_1057,N_14507,N_14879);
or UO_1058 (O_1058,N_14170,N_14554);
or UO_1059 (O_1059,N_14046,N_14097);
xnor UO_1060 (O_1060,N_14254,N_14345);
xor UO_1061 (O_1061,N_14628,N_14464);
or UO_1062 (O_1062,N_14213,N_14362);
and UO_1063 (O_1063,N_14874,N_14679);
xor UO_1064 (O_1064,N_14168,N_14129);
and UO_1065 (O_1065,N_14534,N_14069);
and UO_1066 (O_1066,N_14534,N_14599);
nand UO_1067 (O_1067,N_14784,N_14413);
and UO_1068 (O_1068,N_14386,N_14369);
nand UO_1069 (O_1069,N_14709,N_14390);
xor UO_1070 (O_1070,N_14723,N_14577);
nor UO_1071 (O_1071,N_14299,N_14816);
or UO_1072 (O_1072,N_14241,N_14414);
nor UO_1073 (O_1073,N_14687,N_14857);
nand UO_1074 (O_1074,N_14265,N_14668);
nor UO_1075 (O_1075,N_14524,N_14872);
nand UO_1076 (O_1076,N_14232,N_14143);
nor UO_1077 (O_1077,N_14484,N_14551);
xnor UO_1078 (O_1078,N_14895,N_14718);
or UO_1079 (O_1079,N_14085,N_14584);
and UO_1080 (O_1080,N_14030,N_14821);
nor UO_1081 (O_1081,N_14518,N_14433);
nor UO_1082 (O_1082,N_14221,N_14258);
or UO_1083 (O_1083,N_14822,N_14380);
nand UO_1084 (O_1084,N_14871,N_14671);
or UO_1085 (O_1085,N_14488,N_14340);
nor UO_1086 (O_1086,N_14391,N_14809);
nand UO_1087 (O_1087,N_14974,N_14541);
nor UO_1088 (O_1088,N_14583,N_14308);
xor UO_1089 (O_1089,N_14277,N_14371);
and UO_1090 (O_1090,N_14726,N_14105);
or UO_1091 (O_1091,N_14549,N_14385);
nand UO_1092 (O_1092,N_14110,N_14815);
nand UO_1093 (O_1093,N_14428,N_14756);
xnor UO_1094 (O_1094,N_14013,N_14579);
xnor UO_1095 (O_1095,N_14497,N_14956);
xnor UO_1096 (O_1096,N_14579,N_14649);
xor UO_1097 (O_1097,N_14166,N_14073);
and UO_1098 (O_1098,N_14105,N_14830);
and UO_1099 (O_1099,N_14222,N_14790);
nand UO_1100 (O_1100,N_14319,N_14435);
and UO_1101 (O_1101,N_14080,N_14656);
or UO_1102 (O_1102,N_14103,N_14770);
and UO_1103 (O_1103,N_14600,N_14693);
xnor UO_1104 (O_1104,N_14336,N_14202);
and UO_1105 (O_1105,N_14449,N_14064);
or UO_1106 (O_1106,N_14214,N_14817);
nor UO_1107 (O_1107,N_14257,N_14332);
nor UO_1108 (O_1108,N_14830,N_14167);
or UO_1109 (O_1109,N_14038,N_14059);
nand UO_1110 (O_1110,N_14573,N_14964);
or UO_1111 (O_1111,N_14295,N_14018);
and UO_1112 (O_1112,N_14441,N_14572);
and UO_1113 (O_1113,N_14650,N_14762);
and UO_1114 (O_1114,N_14438,N_14793);
xnor UO_1115 (O_1115,N_14112,N_14130);
nor UO_1116 (O_1116,N_14349,N_14332);
nand UO_1117 (O_1117,N_14042,N_14680);
or UO_1118 (O_1118,N_14224,N_14609);
xor UO_1119 (O_1119,N_14096,N_14024);
and UO_1120 (O_1120,N_14950,N_14769);
or UO_1121 (O_1121,N_14465,N_14451);
nor UO_1122 (O_1122,N_14910,N_14642);
xor UO_1123 (O_1123,N_14494,N_14819);
nand UO_1124 (O_1124,N_14578,N_14160);
and UO_1125 (O_1125,N_14175,N_14264);
xor UO_1126 (O_1126,N_14579,N_14698);
and UO_1127 (O_1127,N_14669,N_14602);
nand UO_1128 (O_1128,N_14911,N_14189);
nand UO_1129 (O_1129,N_14742,N_14223);
nor UO_1130 (O_1130,N_14942,N_14212);
nor UO_1131 (O_1131,N_14601,N_14056);
xnor UO_1132 (O_1132,N_14628,N_14408);
and UO_1133 (O_1133,N_14377,N_14929);
xor UO_1134 (O_1134,N_14398,N_14196);
nor UO_1135 (O_1135,N_14983,N_14871);
nand UO_1136 (O_1136,N_14974,N_14228);
nand UO_1137 (O_1137,N_14169,N_14363);
nor UO_1138 (O_1138,N_14347,N_14744);
nand UO_1139 (O_1139,N_14557,N_14746);
nor UO_1140 (O_1140,N_14187,N_14756);
nand UO_1141 (O_1141,N_14876,N_14180);
xor UO_1142 (O_1142,N_14191,N_14273);
nor UO_1143 (O_1143,N_14460,N_14839);
nand UO_1144 (O_1144,N_14810,N_14224);
or UO_1145 (O_1145,N_14506,N_14796);
nand UO_1146 (O_1146,N_14794,N_14889);
and UO_1147 (O_1147,N_14623,N_14053);
nand UO_1148 (O_1148,N_14360,N_14475);
xnor UO_1149 (O_1149,N_14042,N_14066);
nor UO_1150 (O_1150,N_14250,N_14594);
nand UO_1151 (O_1151,N_14483,N_14440);
and UO_1152 (O_1152,N_14474,N_14858);
xnor UO_1153 (O_1153,N_14796,N_14876);
or UO_1154 (O_1154,N_14958,N_14999);
xnor UO_1155 (O_1155,N_14826,N_14301);
xnor UO_1156 (O_1156,N_14412,N_14967);
and UO_1157 (O_1157,N_14711,N_14095);
or UO_1158 (O_1158,N_14133,N_14775);
nor UO_1159 (O_1159,N_14637,N_14393);
or UO_1160 (O_1160,N_14829,N_14563);
nor UO_1161 (O_1161,N_14228,N_14637);
or UO_1162 (O_1162,N_14641,N_14234);
nor UO_1163 (O_1163,N_14271,N_14123);
nand UO_1164 (O_1164,N_14438,N_14416);
nor UO_1165 (O_1165,N_14434,N_14379);
nor UO_1166 (O_1166,N_14048,N_14695);
nand UO_1167 (O_1167,N_14256,N_14423);
nor UO_1168 (O_1168,N_14005,N_14328);
nor UO_1169 (O_1169,N_14321,N_14822);
or UO_1170 (O_1170,N_14027,N_14152);
and UO_1171 (O_1171,N_14609,N_14827);
and UO_1172 (O_1172,N_14559,N_14900);
and UO_1173 (O_1173,N_14348,N_14555);
and UO_1174 (O_1174,N_14464,N_14389);
or UO_1175 (O_1175,N_14561,N_14210);
xnor UO_1176 (O_1176,N_14284,N_14291);
or UO_1177 (O_1177,N_14452,N_14720);
or UO_1178 (O_1178,N_14142,N_14278);
and UO_1179 (O_1179,N_14654,N_14414);
xnor UO_1180 (O_1180,N_14829,N_14690);
nor UO_1181 (O_1181,N_14932,N_14428);
and UO_1182 (O_1182,N_14770,N_14766);
xnor UO_1183 (O_1183,N_14057,N_14868);
nor UO_1184 (O_1184,N_14208,N_14408);
and UO_1185 (O_1185,N_14625,N_14400);
and UO_1186 (O_1186,N_14973,N_14750);
and UO_1187 (O_1187,N_14370,N_14795);
and UO_1188 (O_1188,N_14516,N_14514);
or UO_1189 (O_1189,N_14206,N_14909);
nor UO_1190 (O_1190,N_14992,N_14593);
nor UO_1191 (O_1191,N_14911,N_14008);
and UO_1192 (O_1192,N_14316,N_14208);
nor UO_1193 (O_1193,N_14050,N_14152);
and UO_1194 (O_1194,N_14511,N_14286);
xnor UO_1195 (O_1195,N_14322,N_14493);
xnor UO_1196 (O_1196,N_14361,N_14015);
xnor UO_1197 (O_1197,N_14718,N_14232);
or UO_1198 (O_1198,N_14334,N_14048);
or UO_1199 (O_1199,N_14308,N_14941);
or UO_1200 (O_1200,N_14081,N_14612);
nor UO_1201 (O_1201,N_14160,N_14470);
xnor UO_1202 (O_1202,N_14114,N_14423);
and UO_1203 (O_1203,N_14006,N_14323);
nor UO_1204 (O_1204,N_14384,N_14962);
xnor UO_1205 (O_1205,N_14032,N_14277);
or UO_1206 (O_1206,N_14485,N_14651);
nand UO_1207 (O_1207,N_14286,N_14040);
nand UO_1208 (O_1208,N_14359,N_14990);
and UO_1209 (O_1209,N_14181,N_14178);
xnor UO_1210 (O_1210,N_14411,N_14982);
xor UO_1211 (O_1211,N_14433,N_14745);
nand UO_1212 (O_1212,N_14600,N_14924);
and UO_1213 (O_1213,N_14391,N_14338);
nor UO_1214 (O_1214,N_14488,N_14960);
and UO_1215 (O_1215,N_14600,N_14105);
and UO_1216 (O_1216,N_14332,N_14939);
xor UO_1217 (O_1217,N_14406,N_14893);
nand UO_1218 (O_1218,N_14099,N_14460);
xor UO_1219 (O_1219,N_14981,N_14986);
xor UO_1220 (O_1220,N_14377,N_14992);
nor UO_1221 (O_1221,N_14010,N_14728);
nand UO_1222 (O_1222,N_14143,N_14216);
nand UO_1223 (O_1223,N_14202,N_14691);
xnor UO_1224 (O_1224,N_14421,N_14405);
or UO_1225 (O_1225,N_14657,N_14510);
or UO_1226 (O_1226,N_14085,N_14451);
nand UO_1227 (O_1227,N_14536,N_14542);
nor UO_1228 (O_1228,N_14133,N_14139);
and UO_1229 (O_1229,N_14733,N_14603);
and UO_1230 (O_1230,N_14423,N_14566);
xor UO_1231 (O_1231,N_14724,N_14780);
xor UO_1232 (O_1232,N_14532,N_14906);
and UO_1233 (O_1233,N_14411,N_14053);
xnor UO_1234 (O_1234,N_14882,N_14001);
xnor UO_1235 (O_1235,N_14699,N_14138);
nand UO_1236 (O_1236,N_14718,N_14271);
and UO_1237 (O_1237,N_14793,N_14257);
xor UO_1238 (O_1238,N_14887,N_14996);
and UO_1239 (O_1239,N_14997,N_14090);
or UO_1240 (O_1240,N_14893,N_14738);
nand UO_1241 (O_1241,N_14848,N_14220);
and UO_1242 (O_1242,N_14418,N_14728);
xor UO_1243 (O_1243,N_14241,N_14832);
nand UO_1244 (O_1244,N_14782,N_14970);
and UO_1245 (O_1245,N_14261,N_14157);
or UO_1246 (O_1246,N_14250,N_14138);
and UO_1247 (O_1247,N_14835,N_14645);
or UO_1248 (O_1248,N_14041,N_14372);
nor UO_1249 (O_1249,N_14567,N_14173);
and UO_1250 (O_1250,N_14702,N_14286);
and UO_1251 (O_1251,N_14209,N_14339);
nor UO_1252 (O_1252,N_14290,N_14892);
nor UO_1253 (O_1253,N_14538,N_14294);
or UO_1254 (O_1254,N_14992,N_14473);
xor UO_1255 (O_1255,N_14164,N_14299);
and UO_1256 (O_1256,N_14843,N_14935);
nand UO_1257 (O_1257,N_14098,N_14132);
and UO_1258 (O_1258,N_14174,N_14938);
and UO_1259 (O_1259,N_14521,N_14245);
nand UO_1260 (O_1260,N_14071,N_14456);
and UO_1261 (O_1261,N_14143,N_14854);
nor UO_1262 (O_1262,N_14930,N_14101);
xnor UO_1263 (O_1263,N_14349,N_14342);
nor UO_1264 (O_1264,N_14048,N_14417);
nand UO_1265 (O_1265,N_14712,N_14966);
xor UO_1266 (O_1266,N_14066,N_14339);
nand UO_1267 (O_1267,N_14091,N_14987);
nand UO_1268 (O_1268,N_14822,N_14423);
nor UO_1269 (O_1269,N_14952,N_14728);
nor UO_1270 (O_1270,N_14062,N_14502);
and UO_1271 (O_1271,N_14861,N_14796);
nor UO_1272 (O_1272,N_14030,N_14466);
nor UO_1273 (O_1273,N_14830,N_14979);
and UO_1274 (O_1274,N_14508,N_14107);
nor UO_1275 (O_1275,N_14809,N_14236);
xor UO_1276 (O_1276,N_14464,N_14674);
nand UO_1277 (O_1277,N_14747,N_14860);
xor UO_1278 (O_1278,N_14173,N_14880);
nand UO_1279 (O_1279,N_14954,N_14059);
and UO_1280 (O_1280,N_14328,N_14492);
nand UO_1281 (O_1281,N_14994,N_14700);
or UO_1282 (O_1282,N_14854,N_14747);
and UO_1283 (O_1283,N_14908,N_14985);
or UO_1284 (O_1284,N_14301,N_14345);
or UO_1285 (O_1285,N_14131,N_14331);
nand UO_1286 (O_1286,N_14896,N_14263);
nand UO_1287 (O_1287,N_14641,N_14141);
or UO_1288 (O_1288,N_14061,N_14672);
nor UO_1289 (O_1289,N_14478,N_14266);
nand UO_1290 (O_1290,N_14341,N_14966);
xor UO_1291 (O_1291,N_14628,N_14553);
and UO_1292 (O_1292,N_14629,N_14332);
nor UO_1293 (O_1293,N_14503,N_14066);
nand UO_1294 (O_1294,N_14547,N_14056);
or UO_1295 (O_1295,N_14192,N_14234);
or UO_1296 (O_1296,N_14438,N_14320);
nor UO_1297 (O_1297,N_14732,N_14358);
nand UO_1298 (O_1298,N_14308,N_14073);
or UO_1299 (O_1299,N_14492,N_14389);
or UO_1300 (O_1300,N_14006,N_14381);
xor UO_1301 (O_1301,N_14489,N_14693);
and UO_1302 (O_1302,N_14231,N_14754);
or UO_1303 (O_1303,N_14281,N_14074);
or UO_1304 (O_1304,N_14913,N_14519);
nor UO_1305 (O_1305,N_14988,N_14800);
and UO_1306 (O_1306,N_14389,N_14157);
or UO_1307 (O_1307,N_14851,N_14686);
and UO_1308 (O_1308,N_14640,N_14381);
xor UO_1309 (O_1309,N_14962,N_14233);
nand UO_1310 (O_1310,N_14595,N_14599);
xor UO_1311 (O_1311,N_14188,N_14326);
and UO_1312 (O_1312,N_14889,N_14717);
nor UO_1313 (O_1313,N_14996,N_14466);
nor UO_1314 (O_1314,N_14058,N_14460);
and UO_1315 (O_1315,N_14460,N_14558);
and UO_1316 (O_1316,N_14008,N_14307);
or UO_1317 (O_1317,N_14305,N_14592);
nand UO_1318 (O_1318,N_14794,N_14026);
nor UO_1319 (O_1319,N_14992,N_14858);
or UO_1320 (O_1320,N_14243,N_14115);
nand UO_1321 (O_1321,N_14197,N_14519);
and UO_1322 (O_1322,N_14304,N_14694);
nand UO_1323 (O_1323,N_14822,N_14968);
and UO_1324 (O_1324,N_14827,N_14535);
or UO_1325 (O_1325,N_14840,N_14128);
xor UO_1326 (O_1326,N_14313,N_14416);
nor UO_1327 (O_1327,N_14208,N_14913);
nand UO_1328 (O_1328,N_14013,N_14569);
xor UO_1329 (O_1329,N_14120,N_14964);
xnor UO_1330 (O_1330,N_14159,N_14657);
and UO_1331 (O_1331,N_14269,N_14947);
xor UO_1332 (O_1332,N_14125,N_14279);
nand UO_1333 (O_1333,N_14638,N_14324);
or UO_1334 (O_1334,N_14959,N_14939);
xor UO_1335 (O_1335,N_14009,N_14811);
xor UO_1336 (O_1336,N_14968,N_14906);
nor UO_1337 (O_1337,N_14444,N_14936);
xnor UO_1338 (O_1338,N_14049,N_14469);
nor UO_1339 (O_1339,N_14550,N_14488);
and UO_1340 (O_1340,N_14951,N_14815);
nor UO_1341 (O_1341,N_14487,N_14261);
and UO_1342 (O_1342,N_14003,N_14070);
and UO_1343 (O_1343,N_14585,N_14577);
xnor UO_1344 (O_1344,N_14965,N_14455);
or UO_1345 (O_1345,N_14448,N_14683);
and UO_1346 (O_1346,N_14578,N_14445);
xor UO_1347 (O_1347,N_14608,N_14953);
and UO_1348 (O_1348,N_14357,N_14971);
nor UO_1349 (O_1349,N_14974,N_14399);
or UO_1350 (O_1350,N_14822,N_14887);
and UO_1351 (O_1351,N_14465,N_14757);
xor UO_1352 (O_1352,N_14546,N_14728);
xor UO_1353 (O_1353,N_14125,N_14051);
nand UO_1354 (O_1354,N_14237,N_14254);
nand UO_1355 (O_1355,N_14989,N_14089);
nor UO_1356 (O_1356,N_14251,N_14683);
nor UO_1357 (O_1357,N_14184,N_14296);
and UO_1358 (O_1358,N_14708,N_14140);
and UO_1359 (O_1359,N_14906,N_14931);
xor UO_1360 (O_1360,N_14095,N_14472);
nand UO_1361 (O_1361,N_14158,N_14085);
nor UO_1362 (O_1362,N_14076,N_14678);
xor UO_1363 (O_1363,N_14360,N_14540);
nor UO_1364 (O_1364,N_14605,N_14733);
xor UO_1365 (O_1365,N_14250,N_14074);
and UO_1366 (O_1366,N_14072,N_14524);
or UO_1367 (O_1367,N_14727,N_14924);
nand UO_1368 (O_1368,N_14752,N_14336);
nand UO_1369 (O_1369,N_14202,N_14753);
nand UO_1370 (O_1370,N_14779,N_14954);
xor UO_1371 (O_1371,N_14994,N_14367);
xnor UO_1372 (O_1372,N_14240,N_14414);
nand UO_1373 (O_1373,N_14536,N_14273);
and UO_1374 (O_1374,N_14668,N_14395);
and UO_1375 (O_1375,N_14798,N_14134);
nor UO_1376 (O_1376,N_14308,N_14558);
and UO_1377 (O_1377,N_14449,N_14405);
and UO_1378 (O_1378,N_14792,N_14891);
and UO_1379 (O_1379,N_14591,N_14160);
nor UO_1380 (O_1380,N_14678,N_14964);
nor UO_1381 (O_1381,N_14336,N_14682);
nor UO_1382 (O_1382,N_14230,N_14081);
and UO_1383 (O_1383,N_14046,N_14942);
xor UO_1384 (O_1384,N_14375,N_14535);
nor UO_1385 (O_1385,N_14929,N_14883);
or UO_1386 (O_1386,N_14314,N_14332);
nor UO_1387 (O_1387,N_14613,N_14935);
xnor UO_1388 (O_1388,N_14163,N_14336);
or UO_1389 (O_1389,N_14101,N_14557);
and UO_1390 (O_1390,N_14084,N_14919);
xor UO_1391 (O_1391,N_14064,N_14919);
nand UO_1392 (O_1392,N_14775,N_14912);
and UO_1393 (O_1393,N_14703,N_14844);
xor UO_1394 (O_1394,N_14192,N_14787);
nor UO_1395 (O_1395,N_14944,N_14161);
or UO_1396 (O_1396,N_14298,N_14041);
or UO_1397 (O_1397,N_14916,N_14643);
or UO_1398 (O_1398,N_14416,N_14189);
xor UO_1399 (O_1399,N_14481,N_14774);
xor UO_1400 (O_1400,N_14065,N_14364);
nand UO_1401 (O_1401,N_14729,N_14760);
nor UO_1402 (O_1402,N_14227,N_14706);
nand UO_1403 (O_1403,N_14094,N_14026);
nand UO_1404 (O_1404,N_14299,N_14292);
xor UO_1405 (O_1405,N_14087,N_14972);
nand UO_1406 (O_1406,N_14408,N_14060);
and UO_1407 (O_1407,N_14445,N_14814);
xor UO_1408 (O_1408,N_14787,N_14102);
nand UO_1409 (O_1409,N_14990,N_14095);
nand UO_1410 (O_1410,N_14139,N_14159);
xor UO_1411 (O_1411,N_14272,N_14480);
or UO_1412 (O_1412,N_14693,N_14136);
xnor UO_1413 (O_1413,N_14757,N_14779);
xor UO_1414 (O_1414,N_14346,N_14531);
nor UO_1415 (O_1415,N_14916,N_14953);
xor UO_1416 (O_1416,N_14057,N_14456);
nor UO_1417 (O_1417,N_14503,N_14254);
or UO_1418 (O_1418,N_14711,N_14281);
nor UO_1419 (O_1419,N_14467,N_14583);
xor UO_1420 (O_1420,N_14339,N_14963);
nor UO_1421 (O_1421,N_14981,N_14036);
nor UO_1422 (O_1422,N_14344,N_14381);
xor UO_1423 (O_1423,N_14155,N_14291);
nor UO_1424 (O_1424,N_14778,N_14218);
or UO_1425 (O_1425,N_14960,N_14640);
and UO_1426 (O_1426,N_14258,N_14424);
xor UO_1427 (O_1427,N_14417,N_14352);
nor UO_1428 (O_1428,N_14491,N_14384);
nand UO_1429 (O_1429,N_14978,N_14507);
nor UO_1430 (O_1430,N_14468,N_14383);
and UO_1431 (O_1431,N_14586,N_14100);
nor UO_1432 (O_1432,N_14291,N_14268);
xnor UO_1433 (O_1433,N_14790,N_14380);
and UO_1434 (O_1434,N_14883,N_14947);
xor UO_1435 (O_1435,N_14329,N_14037);
and UO_1436 (O_1436,N_14251,N_14323);
or UO_1437 (O_1437,N_14386,N_14327);
xnor UO_1438 (O_1438,N_14303,N_14890);
nor UO_1439 (O_1439,N_14215,N_14135);
nand UO_1440 (O_1440,N_14325,N_14624);
nor UO_1441 (O_1441,N_14487,N_14907);
xor UO_1442 (O_1442,N_14895,N_14965);
or UO_1443 (O_1443,N_14406,N_14498);
xnor UO_1444 (O_1444,N_14618,N_14677);
nor UO_1445 (O_1445,N_14903,N_14030);
xnor UO_1446 (O_1446,N_14892,N_14835);
or UO_1447 (O_1447,N_14017,N_14754);
and UO_1448 (O_1448,N_14173,N_14396);
and UO_1449 (O_1449,N_14030,N_14225);
nand UO_1450 (O_1450,N_14299,N_14684);
nand UO_1451 (O_1451,N_14829,N_14791);
nor UO_1452 (O_1452,N_14366,N_14890);
nand UO_1453 (O_1453,N_14102,N_14782);
nor UO_1454 (O_1454,N_14241,N_14326);
and UO_1455 (O_1455,N_14217,N_14351);
nor UO_1456 (O_1456,N_14188,N_14828);
or UO_1457 (O_1457,N_14078,N_14396);
or UO_1458 (O_1458,N_14245,N_14485);
xor UO_1459 (O_1459,N_14426,N_14631);
and UO_1460 (O_1460,N_14683,N_14640);
xnor UO_1461 (O_1461,N_14334,N_14164);
xnor UO_1462 (O_1462,N_14911,N_14457);
nor UO_1463 (O_1463,N_14851,N_14361);
nor UO_1464 (O_1464,N_14079,N_14918);
and UO_1465 (O_1465,N_14993,N_14372);
and UO_1466 (O_1466,N_14825,N_14758);
or UO_1467 (O_1467,N_14865,N_14294);
nand UO_1468 (O_1468,N_14470,N_14490);
nor UO_1469 (O_1469,N_14811,N_14977);
nor UO_1470 (O_1470,N_14438,N_14710);
nand UO_1471 (O_1471,N_14054,N_14940);
xor UO_1472 (O_1472,N_14762,N_14818);
nand UO_1473 (O_1473,N_14044,N_14147);
xnor UO_1474 (O_1474,N_14355,N_14043);
nand UO_1475 (O_1475,N_14019,N_14476);
and UO_1476 (O_1476,N_14605,N_14604);
xor UO_1477 (O_1477,N_14327,N_14979);
and UO_1478 (O_1478,N_14612,N_14644);
nor UO_1479 (O_1479,N_14752,N_14936);
xnor UO_1480 (O_1480,N_14951,N_14609);
nor UO_1481 (O_1481,N_14321,N_14605);
and UO_1482 (O_1482,N_14002,N_14368);
nor UO_1483 (O_1483,N_14908,N_14456);
nor UO_1484 (O_1484,N_14873,N_14335);
or UO_1485 (O_1485,N_14092,N_14982);
or UO_1486 (O_1486,N_14486,N_14126);
and UO_1487 (O_1487,N_14814,N_14152);
nand UO_1488 (O_1488,N_14596,N_14784);
xor UO_1489 (O_1489,N_14725,N_14429);
nand UO_1490 (O_1490,N_14700,N_14744);
nor UO_1491 (O_1491,N_14729,N_14108);
nand UO_1492 (O_1492,N_14274,N_14232);
nor UO_1493 (O_1493,N_14151,N_14400);
or UO_1494 (O_1494,N_14882,N_14121);
xor UO_1495 (O_1495,N_14152,N_14670);
xor UO_1496 (O_1496,N_14027,N_14157);
xnor UO_1497 (O_1497,N_14673,N_14963);
nand UO_1498 (O_1498,N_14512,N_14143);
or UO_1499 (O_1499,N_14850,N_14995);
or UO_1500 (O_1500,N_14972,N_14598);
and UO_1501 (O_1501,N_14923,N_14313);
or UO_1502 (O_1502,N_14592,N_14498);
xnor UO_1503 (O_1503,N_14171,N_14649);
xor UO_1504 (O_1504,N_14506,N_14121);
nor UO_1505 (O_1505,N_14987,N_14635);
or UO_1506 (O_1506,N_14503,N_14302);
or UO_1507 (O_1507,N_14511,N_14425);
and UO_1508 (O_1508,N_14480,N_14860);
nor UO_1509 (O_1509,N_14197,N_14107);
and UO_1510 (O_1510,N_14906,N_14215);
nor UO_1511 (O_1511,N_14858,N_14590);
nor UO_1512 (O_1512,N_14156,N_14492);
nand UO_1513 (O_1513,N_14475,N_14788);
or UO_1514 (O_1514,N_14293,N_14704);
and UO_1515 (O_1515,N_14142,N_14110);
and UO_1516 (O_1516,N_14499,N_14991);
nor UO_1517 (O_1517,N_14444,N_14387);
nand UO_1518 (O_1518,N_14962,N_14073);
nor UO_1519 (O_1519,N_14227,N_14087);
and UO_1520 (O_1520,N_14472,N_14242);
nor UO_1521 (O_1521,N_14555,N_14601);
nand UO_1522 (O_1522,N_14312,N_14603);
and UO_1523 (O_1523,N_14980,N_14712);
nor UO_1524 (O_1524,N_14070,N_14153);
or UO_1525 (O_1525,N_14975,N_14840);
and UO_1526 (O_1526,N_14393,N_14073);
and UO_1527 (O_1527,N_14948,N_14708);
nor UO_1528 (O_1528,N_14837,N_14011);
xor UO_1529 (O_1529,N_14039,N_14210);
nor UO_1530 (O_1530,N_14632,N_14942);
nand UO_1531 (O_1531,N_14078,N_14834);
or UO_1532 (O_1532,N_14177,N_14960);
xnor UO_1533 (O_1533,N_14540,N_14014);
nor UO_1534 (O_1534,N_14340,N_14992);
or UO_1535 (O_1535,N_14942,N_14171);
xnor UO_1536 (O_1536,N_14337,N_14215);
and UO_1537 (O_1537,N_14267,N_14216);
or UO_1538 (O_1538,N_14134,N_14643);
nor UO_1539 (O_1539,N_14436,N_14055);
nand UO_1540 (O_1540,N_14825,N_14397);
or UO_1541 (O_1541,N_14569,N_14559);
nand UO_1542 (O_1542,N_14266,N_14618);
and UO_1543 (O_1543,N_14691,N_14421);
xor UO_1544 (O_1544,N_14653,N_14492);
and UO_1545 (O_1545,N_14881,N_14139);
xnor UO_1546 (O_1546,N_14246,N_14420);
or UO_1547 (O_1547,N_14152,N_14133);
nor UO_1548 (O_1548,N_14290,N_14649);
xnor UO_1549 (O_1549,N_14079,N_14133);
nor UO_1550 (O_1550,N_14348,N_14802);
or UO_1551 (O_1551,N_14425,N_14606);
or UO_1552 (O_1552,N_14597,N_14319);
nor UO_1553 (O_1553,N_14920,N_14958);
nand UO_1554 (O_1554,N_14496,N_14072);
nor UO_1555 (O_1555,N_14581,N_14687);
or UO_1556 (O_1556,N_14945,N_14948);
xor UO_1557 (O_1557,N_14808,N_14179);
nand UO_1558 (O_1558,N_14526,N_14604);
and UO_1559 (O_1559,N_14120,N_14643);
and UO_1560 (O_1560,N_14068,N_14267);
or UO_1561 (O_1561,N_14092,N_14572);
and UO_1562 (O_1562,N_14931,N_14134);
and UO_1563 (O_1563,N_14762,N_14078);
nand UO_1564 (O_1564,N_14185,N_14892);
xor UO_1565 (O_1565,N_14753,N_14320);
nor UO_1566 (O_1566,N_14683,N_14727);
nor UO_1567 (O_1567,N_14534,N_14673);
xnor UO_1568 (O_1568,N_14881,N_14758);
or UO_1569 (O_1569,N_14322,N_14609);
and UO_1570 (O_1570,N_14928,N_14672);
nand UO_1571 (O_1571,N_14849,N_14132);
and UO_1572 (O_1572,N_14368,N_14855);
or UO_1573 (O_1573,N_14965,N_14328);
or UO_1574 (O_1574,N_14829,N_14105);
nand UO_1575 (O_1575,N_14397,N_14952);
or UO_1576 (O_1576,N_14050,N_14631);
nor UO_1577 (O_1577,N_14468,N_14078);
and UO_1578 (O_1578,N_14894,N_14280);
nand UO_1579 (O_1579,N_14656,N_14858);
xor UO_1580 (O_1580,N_14874,N_14093);
nor UO_1581 (O_1581,N_14475,N_14736);
nor UO_1582 (O_1582,N_14609,N_14163);
nand UO_1583 (O_1583,N_14438,N_14711);
or UO_1584 (O_1584,N_14941,N_14028);
xnor UO_1585 (O_1585,N_14116,N_14972);
xnor UO_1586 (O_1586,N_14272,N_14401);
xor UO_1587 (O_1587,N_14749,N_14757);
nand UO_1588 (O_1588,N_14286,N_14273);
nand UO_1589 (O_1589,N_14335,N_14528);
nand UO_1590 (O_1590,N_14803,N_14275);
and UO_1591 (O_1591,N_14329,N_14370);
or UO_1592 (O_1592,N_14879,N_14345);
nor UO_1593 (O_1593,N_14323,N_14670);
xnor UO_1594 (O_1594,N_14451,N_14137);
or UO_1595 (O_1595,N_14419,N_14232);
and UO_1596 (O_1596,N_14698,N_14791);
xnor UO_1597 (O_1597,N_14324,N_14622);
xnor UO_1598 (O_1598,N_14077,N_14064);
or UO_1599 (O_1599,N_14821,N_14421);
nor UO_1600 (O_1600,N_14916,N_14417);
and UO_1601 (O_1601,N_14941,N_14736);
or UO_1602 (O_1602,N_14537,N_14269);
or UO_1603 (O_1603,N_14777,N_14350);
xor UO_1604 (O_1604,N_14578,N_14447);
xor UO_1605 (O_1605,N_14224,N_14291);
xnor UO_1606 (O_1606,N_14635,N_14530);
xnor UO_1607 (O_1607,N_14435,N_14588);
nand UO_1608 (O_1608,N_14594,N_14537);
or UO_1609 (O_1609,N_14996,N_14014);
xnor UO_1610 (O_1610,N_14939,N_14189);
or UO_1611 (O_1611,N_14809,N_14430);
nor UO_1612 (O_1612,N_14780,N_14584);
xor UO_1613 (O_1613,N_14850,N_14696);
or UO_1614 (O_1614,N_14077,N_14663);
nor UO_1615 (O_1615,N_14861,N_14315);
nand UO_1616 (O_1616,N_14008,N_14012);
and UO_1617 (O_1617,N_14986,N_14318);
xnor UO_1618 (O_1618,N_14286,N_14800);
and UO_1619 (O_1619,N_14155,N_14310);
or UO_1620 (O_1620,N_14051,N_14835);
nand UO_1621 (O_1621,N_14371,N_14160);
nor UO_1622 (O_1622,N_14166,N_14996);
xor UO_1623 (O_1623,N_14806,N_14965);
xnor UO_1624 (O_1624,N_14207,N_14928);
or UO_1625 (O_1625,N_14062,N_14094);
nand UO_1626 (O_1626,N_14703,N_14103);
nor UO_1627 (O_1627,N_14544,N_14932);
nor UO_1628 (O_1628,N_14218,N_14498);
nand UO_1629 (O_1629,N_14758,N_14419);
and UO_1630 (O_1630,N_14338,N_14967);
xor UO_1631 (O_1631,N_14917,N_14821);
or UO_1632 (O_1632,N_14010,N_14321);
or UO_1633 (O_1633,N_14836,N_14205);
nor UO_1634 (O_1634,N_14636,N_14125);
nor UO_1635 (O_1635,N_14374,N_14699);
nand UO_1636 (O_1636,N_14217,N_14809);
nor UO_1637 (O_1637,N_14138,N_14832);
and UO_1638 (O_1638,N_14962,N_14612);
and UO_1639 (O_1639,N_14887,N_14641);
nor UO_1640 (O_1640,N_14839,N_14155);
nand UO_1641 (O_1641,N_14376,N_14534);
nand UO_1642 (O_1642,N_14930,N_14826);
nand UO_1643 (O_1643,N_14345,N_14442);
xnor UO_1644 (O_1644,N_14219,N_14584);
nand UO_1645 (O_1645,N_14620,N_14494);
nand UO_1646 (O_1646,N_14749,N_14695);
or UO_1647 (O_1647,N_14526,N_14052);
nand UO_1648 (O_1648,N_14840,N_14045);
nand UO_1649 (O_1649,N_14745,N_14476);
and UO_1650 (O_1650,N_14371,N_14492);
or UO_1651 (O_1651,N_14368,N_14075);
nor UO_1652 (O_1652,N_14551,N_14780);
nor UO_1653 (O_1653,N_14153,N_14557);
and UO_1654 (O_1654,N_14144,N_14132);
nand UO_1655 (O_1655,N_14551,N_14261);
and UO_1656 (O_1656,N_14476,N_14899);
and UO_1657 (O_1657,N_14489,N_14137);
nand UO_1658 (O_1658,N_14436,N_14565);
or UO_1659 (O_1659,N_14307,N_14618);
and UO_1660 (O_1660,N_14347,N_14726);
or UO_1661 (O_1661,N_14038,N_14775);
xor UO_1662 (O_1662,N_14752,N_14571);
nor UO_1663 (O_1663,N_14478,N_14702);
or UO_1664 (O_1664,N_14070,N_14759);
xor UO_1665 (O_1665,N_14426,N_14028);
nor UO_1666 (O_1666,N_14834,N_14399);
and UO_1667 (O_1667,N_14567,N_14431);
or UO_1668 (O_1668,N_14781,N_14428);
xnor UO_1669 (O_1669,N_14974,N_14408);
xnor UO_1670 (O_1670,N_14616,N_14009);
or UO_1671 (O_1671,N_14033,N_14235);
and UO_1672 (O_1672,N_14191,N_14523);
or UO_1673 (O_1673,N_14419,N_14913);
or UO_1674 (O_1674,N_14314,N_14166);
xnor UO_1675 (O_1675,N_14593,N_14199);
xnor UO_1676 (O_1676,N_14409,N_14978);
nand UO_1677 (O_1677,N_14032,N_14033);
nor UO_1678 (O_1678,N_14144,N_14440);
nor UO_1679 (O_1679,N_14146,N_14148);
xnor UO_1680 (O_1680,N_14026,N_14240);
and UO_1681 (O_1681,N_14691,N_14046);
nor UO_1682 (O_1682,N_14991,N_14583);
and UO_1683 (O_1683,N_14899,N_14489);
nor UO_1684 (O_1684,N_14695,N_14890);
or UO_1685 (O_1685,N_14794,N_14988);
nand UO_1686 (O_1686,N_14219,N_14836);
and UO_1687 (O_1687,N_14776,N_14041);
or UO_1688 (O_1688,N_14717,N_14513);
and UO_1689 (O_1689,N_14102,N_14964);
nor UO_1690 (O_1690,N_14136,N_14382);
xor UO_1691 (O_1691,N_14409,N_14551);
nor UO_1692 (O_1692,N_14850,N_14793);
or UO_1693 (O_1693,N_14381,N_14143);
xor UO_1694 (O_1694,N_14229,N_14237);
nor UO_1695 (O_1695,N_14488,N_14354);
nor UO_1696 (O_1696,N_14515,N_14625);
and UO_1697 (O_1697,N_14303,N_14175);
xnor UO_1698 (O_1698,N_14045,N_14457);
nand UO_1699 (O_1699,N_14718,N_14426);
and UO_1700 (O_1700,N_14345,N_14583);
nand UO_1701 (O_1701,N_14124,N_14378);
or UO_1702 (O_1702,N_14124,N_14298);
nor UO_1703 (O_1703,N_14498,N_14221);
and UO_1704 (O_1704,N_14926,N_14035);
nand UO_1705 (O_1705,N_14018,N_14207);
nor UO_1706 (O_1706,N_14942,N_14646);
xor UO_1707 (O_1707,N_14467,N_14755);
nor UO_1708 (O_1708,N_14363,N_14778);
nand UO_1709 (O_1709,N_14075,N_14301);
nor UO_1710 (O_1710,N_14052,N_14705);
nand UO_1711 (O_1711,N_14337,N_14564);
nand UO_1712 (O_1712,N_14462,N_14368);
xor UO_1713 (O_1713,N_14013,N_14831);
xnor UO_1714 (O_1714,N_14566,N_14581);
xor UO_1715 (O_1715,N_14437,N_14315);
xnor UO_1716 (O_1716,N_14847,N_14732);
or UO_1717 (O_1717,N_14150,N_14646);
or UO_1718 (O_1718,N_14603,N_14342);
nand UO_1719 (O_1719,N_14071,N_14762);
and UO_1720 (O_1720,N_14997,N_14905);
nor UO_1721 (O_1721,N_14195,N_14213);
or UO_1722 (O_1722,N_14155,N_14640);
nand UO_1723 (O_1723,N_14891,N_14822);
xor UO_1724 (O_1724,N_14699,N_14251);
or UO_1725 (O_1725,N_14949,N_14757);
nand UO_1726 (O_1726,N_14813,N_14380);
xor UO_1727 (O_1727,N_14840,N_14777);
nand UO_1728 (O_1728,N_14097,N_14204);
nor UO_1729 (O_1729,N_14836,N_14788);
xnor UO_1730 (O_1730,N_14458,N_14475);
nor UO_1731 (O_1731,N_14552,N_14275);
xnor UO_1732 (O_1732,N_14259,N_14816);
xnor UO_1733 (O_1733,N_14722,N_14096);
xnor UO_1734 (O_1734,N_14101,N_14626);
and UO_1735 (O_1735,N_14366,N_14969);
or UO_1736 (O_1736,N_14586,N_14112);
or UO_1737 (O_1737,N_14446,N_14712);
xor UO_1738 (O_1738,N_14260,N_14927);
nor UO_1739 (O_1739,N_14674,N_14426);
and UO_1740 (O_1740,N_14800,N_14772);
nor UO_1741 (O_1741,N_14862,N_14690);
nand UO_1742 (O_1742,N_14547,N_14285);
and UO_1743 (O_1743,N_14891,N_14178);
or UO_1744 (O_1744,N_14032,N_14527);
and UO_1745 (O_1745,N_14890,N_14898);
and UO_1746 (O_1746,N_14516,N_14186);
and UO_1747 (O_1747,N_14091,N_14301);
and UO_1748 (O_1748,N_14769,N_14017);
and UO_1749 (O_1749,N_14375,N_14583);
nor UO_1750 (O_1750,N_14895,N_14494);
nand UO_1751 (O_1751,N_14400,N_14978);
or UO_1752 (O_1752,N_14026,N_14910);
nor UO_1753 (O_1753,N_14512,N_14685);
and UO_1754 (O_1754,N_14352,N_14123);
xnor UO_1755 (O_1755,N_14784,N_14932);
xor UO_1756 (O_1756,N_14512,N_14887);
or UO_1757 (O_1757,N_14461,N_14227);
nand UO_1758 (O_1758,N_14132,N_14211);
xor UO_1759 (O_1759,N_14010,N_14607);
and UO_1760 (O_1760,N_14671,N_14329);
xor UO_1761 (O_1761,N_14824,N_14702);
and UO_1762 (O_1762,N_14035,N_14006);
and UO_1763 (O_1763,N_14395,N_14195);
nand UO_1764 (O_1764,N_14109,N_14135);
and UO_1765 (O_1765,N_14150,N_14091);
or UO_1766 (O_1766,N_14509,N_14188);
xnor UO_1767 (O_1767,N_14593,N_14060);
nor UO_1768 (O_1768,N_14087,N_14205);
xor UO_1769 (O_1769,N_14139,N_14097);
nor UO_1770 (O_1770,N_14372,N_14685);
nor UO_1771 (O_1771,N_14171,N_14092);
nor UO_1772 (O_1772,N_14886,N_14638);
and UO_1773 (O_1773,N_14793,N_14973);
nand UO_1774 (O_1774,N_14576,N_14901);
xnor UO_1775 (O_1775,N_14900,N_14598);
or UO_1776 (O_1776,N_14007,N_14542);
nand UO_1777 (O_1777,N_14363,N_14977);
or UO_1778 (O_1778,N_14706,N_14132);
nor UO_1779 (O_1779,N_14961,N_14544);
xor UO_1780 (O_1780,N_14032,N_14035);
and UO_1781 (O_1781,N_14856,N_14429);
or UO_1782 (O_1782,N_14539,N_14100);
nand UO_1783 (O_1783,N_14075,N_14181);
nand UO_1784 (O_1784,N_14283,N_14628);
or UO_1785 (O_1785,N_14076,N_14072);
xnor UO_1786 (O_1786,N_14449,N_14443);
nand UO_1787 (O_1787,N_14743,N_14956);
nand UO_1788 (O_1788,N_14686,N_14626);
xor UO_1789 (O_1789,N_14068,N_14895);
xnor UO_1790 (O_1790,N_14716,N_14876);
xnor UO_1791 (O_1791,N_14855,N_14077);
xnor UO_1792 (O_1792,N_14207,N_14952);
and UO_1793 (O_1793,N_14945,N_14009);
nor UO_1794 (O_1794,N_14947,N_14877);
nand UO_1795 (O_1795,N_14490,N_14613);
nor UO_1796 (O_1796,N_14199,N_14221);
or UO_1797 (O_1797,N_14654,N_14570);
nand UO_1798 (O_1798,N_14994,N_14749);
nor UO_1799 (O_1799,N_14813,N_14074);
xor UO_1800 (O_1800,N_14535,N_14729);
nor UO_1801 (O_1801,N_14208,N_14814);
nand UO_1802 (O_1802,N_14099,N_14291);
xor UO_1803 (O_1803,N_14418,N_14586);
or UO_1804 (O_1804,N_14862,N_14139);
or UO_1805 (O_1805,N_14060,N_14000);
nand UO_1806 (O_1806,N_14142,N_14324);
xnor UO_1807 (O_1807,N_14433,N_14826);
and UO_1808 (O_1808,N_14464,N_14996);
nand UO_1809 (O_1809,N_14847,N_14134);
nor UO_1810 (O_1810,N_14165,N_14660);
or UO_1811 (O_1811,N_14990,N_14404);
nor UO_1812 (O_1812,N_14582,N_14996);
nand UO_1813 (O_1813,N_14665,N_14526);
nand UO_1814 (O_1814,N_14637,N_14595);
nand UO_1815 (O_1815,N_14159,N_14221);
and UO_1816 (O_1816,N_14752,N_14436);
nor UO_1817 (O_1817,N_14070,N_14012);
or UO_1818 (O_1818,N_14593,N_14394);
xor UO_1819 (O_1819,N_14441,N_14307);
and UO_1820 (O_1820,N_14562,N_14187);
nand UO_1821 (O_1821,N_14215,N_14034);
nor UO_1822 (O_1822,N_14651,N_14187);
nand UO_1823 (O_1823,N_14612,N_14155);
xor UO_1824 (O_1824,N_14280,N_14403);
xor UO_1825 (O_1825,N_14410,N_14843);
or UO_1826 (O_1826,N_14333,N_14140);
and UO_1827 (O_1827,N_14634,N_14433);
or UO_1828 (O_1828,N_14407,N_14098);
or UO_1829 (O_1829,N_14081,N_14663);
xor UO_1830 (O_1830,N_14922,N_14220);
or UO_1831 (O_1831,N_14251,N_14794);
xnor UO_1832 (O_1832,N_14049,N_14192);
nor UO_1833 (O_1833,N_14705,N_14170);
nor UO_1834 (O_1834,N_14320,N_14970);
or UO_1835 (O_1835,N_14218,N_14129);
or UO_1836 (O_1836,N_14599,N_14909);
or UO_1837 (O_1837,N_14367,N_14114);
xor UO_1838 (O_1838,N_14032,N_14977);
nand UO_1839 (O_1839,N_14499,N_14159);
nand UO_1840 (O_1840,N_14912,N_14386);
and UO_1841 (O_1841,N_14457,N_14080);
and UO_1842 (O_1842,N_14574,N_14961);
xnor UO_1843 (O_1843,N_14802,N_14350);
nor UO_1844 (O_1844,N_14369,N_14800);
xor UO_1845 (O_1845,N_14063,N_14793);
and UO_1846 (O_1846,N_14415,N_14124);
and UO_1847 (O_1847,N_14175,N_14714);
or UO_1848 (O_1848,N_14740,N_14125);
or UO_1849 (O_1849,N_14583,N_14709);
nand UO_1850 (O_1850,N_14078,N_14618);
and UO_1851 (O_1851,N_14485,N_14833);
or UO_1852 (O_1852,N_14357,N_14679);
nor UO_1853 (O_1853,N_14034,N_14979);
xnor UO_1854 (O_1854,N_14758,N_14644);
and UO_1855 (O_1855,N_14254,N_14640);
or UO_1856 (O_1856,N_14137,N_14128);
xor UO_1857 (O_1857,N_14442,N_14955);
nor UO_1858 (O_1858,N_14956,N_14079);
or UO_1859 (O_1859,N_14916,N_14702);
xor UO_1860 (O_1860,N_14086,N_14511);
or UO_1861 (O_1861,N_14694,N_14815);
or UO_1862 (O_1862,N_14631,N_14037);
nand UO_1863 (O_1863,N_14980,N_14294);
or UO_1864 (O_1864,N_14512,N_14903);
and UO_1865 (O_1865,N_14198,N_14261);
nor UO_1866 (O_1866,N_14125,N_14334);
and UO_1867 (O_1867,N_14800,N_14426);
or UO_1868 (O_1868,N_14572,N_14337);
xnor UO_1869 (O_1869,N_14802,N_14713);
and UO_1870 (O_1870,N_14839,N_14154);
nand UO_1871 (O_1871,N_14773,N_14038);
or UO_1872 (O_1872,N_14506,N_14742);
nor UO_1873 (O_1873,N_14943,N_14850);
nand UO_1874 (O_1874,N_14948,N_14967);
nand UO_1875 (O_1875,N_14902,N_14807);
or UO_1876 (O_1876,N_14464,N_14998);
nor UO_1877 (O_1877,N_14750,N_14166);
nand UO_1878 (O_1878,N_14899,N_14130);
nor UO_1879 (O_1879,N_14717,N_14242);
xnor UO_1880 (O_1880,N_14648,N_14818);
xnor UO_1881 (O_1881,N_14200,N_14014);
or UO_1882 (O_1882,N_14047,N_14167);
and UO_1883 (O_1883,N_14107,N_14637);
nand UO_1884 (O_1884,N_14626,N_14271);
nor UO_1885 (O_1885,N_14685,N_14364);
and UO_1886 (O_1886,N_14749,N_14696);
nor UO_1887 (O_1887,N_14377,N_14446);
or UO_1888 (O_1888,N_14409,N_14599);
nor UO_1889 (O_1889,N_14243,N_14874);
or UO_1890 (O_1890,N_14317,N_14058);
nand UO_1891 (O_1891,N_14969,N_14102);
nor UO_1892 (O_1892,N_14785,N_14218);
xor UO_1893 (O_1893,N_14241,N_14559);
xor UO_1894 (O_1894,N_14502,N_14184);
nand UO_1895 (O_1895,N_14624,N_14599);
nand UO_1896 (O_1896,N_14071,N_14125);
xnor UO_1897 (O_1897,N_14886,N_14019);
xor UO_1898 (O_1898,N_14002,N_14824);
or UO_1899 (O_1899,N_14010,N_14238);
or UO_1900 (O_1900,N_14859,N_14265);
nand UO_1901 (O_1901,N_14945,N_14697);
or UO_1902 (O_1902,N_14528,N_14465);
and UO_1903 (O_1903,N_14377,N_14487);
nand UO_1904 (O_1904,N_14361,N_14035);
nand UO_1905 (O_1905,N_14973,N_14016);
and UO_1906 (O_1906,N_14768,N_14999);
nor UO_1907 (O_1907,N_14196,N_14958);
nor UO_1908 (O_1908,N_14576,N_14309);
xor UO_1909 (O_1909,N_14684,N_14292);
xor UO_1910 (O_1910,N_14399,N_14487);
and UO_1911 (O_1911,N_14208,N_14891);
and UO_1912 (O_1912,N_14090,N_14376);
or UO_1913 (O_1913,N_14787,N_14258);
xor UO_1914 (O_1914,N_14144,N_14745);
and UO_1915 (O_1915,N_14826,N_14703);
nand UO_1916 (O_1916,N_14176,N_14098);
and UO_1917 (O_1917,N_14729,N_14709);
xnor UO_1918 (O_1918,N_14967,N_14869);
nand UO_1919 (O_1919,N_14151,N_14335);
and UO_1920 (O_1920,N_14432,N_14724);
xor UO_1921 (O_1921,N_14081,N_14366);
nor UO_1922 (O_1922,N_14285,N_14899);
or UO_1923 (O_1923,N_14386,N_14320);
xnor UO_1924 (O_1924,N_14408,N_14277);
or UO_1925 (O_1925,N_14792,N_14773);
and UO_1926 (O_1926,N_14324,N_14004);
xnor UO_1927 (O_1927,N_14157,N_14976);
and UO_1928 (O_1928,N_14138,N_14865);
or UO_1929 (O_1929,N_14729,N_14792);
and UO_1930 (O_1930,N_14047,N_14971);
nor UO_1931 (O_1931,N_14742,N_14561);
and UO_1932 (O_1932,N_14481,N_14813);
nand UO_1933 (O_1933,N_14644,N_14530);
nor UO_1934 (O_1934,N_14200,N_14641);
or UO_1935 (O_1935,N_14584,N_14113);
nor UO_1936 (O_1936,N_14204,N_14805);
xor UO_1937 (O_1937,N_14696,N_14657);
or UO_1938 (O_1938,N_14078,N_14928);
nor UO_1939 (O_1939,N_14746,N_14624);
nor UO_1940 (O_1940,N_14677,N_14188);
xor UO_1941 (O_1941,N_14006,N_14281);
xnor UO_1942 (O_1942,N_14553,N_14277);
nand UO_1943 (O_1943,N_14160,N_14904);
xor UO_1944 (O_1944,N_14312,N_14036);
nor UO_1945 (O_1945,N_14922,N_14875);
xor UO_1946 (O_1946,N_14596,N_14095);
and UO_1947 (O_1947,N_14480,N_14508);
nor UO_1948 (O_1948,N_14280,N_14080);
or UO_1949 (O_1949,N_14603,N_14590);
or UO_1950 (O_1950,N_14813,N_14226);
nand UO_1951 (O_1951,N_14759,N_14017);
xor UO_1952 (O_1952,N_14710,N_14114);
nand UO_1953 (O_1953,N_14847,N_14004);
xnor UO_1954 (O_1954,N_14055,N_14469);
or UO_1955 (O_1955,N_14253,N_14480);
xnor UO_1956 (O_1956,N_14026,N_14067);
nand UO_1957 (O_1957,N_14032,N_14056);
and UO_1958 (O_1958,N_14927,N_14250);
and UO_1959 (O_1959,N_14058,N_14248);
or UO_1960 (O_1960,N_14779,N_14085);
and UO_1961 (O_1961,N_14509,N_14309);
nor UO_1962 (O_1962,N_14947,N_14853);
or UO_1963 (O_1963,N_14342,N_14674);
xnor UO_1964 (O_1964,N_14149,N_14422);
or UO_1965 (O_1965,N_14624,N_14581);
nand UO_1966 (O_1966,N_14820,N_14131);
and UO_1967 (O_1967,N_14641,N_14518);
nand UO_1968 (O_1968,N_14679,N_14076);
nor UO_1969 (O_1969,N_14610,N_14839);
and UO_1970 (O_1970,N_14335,N_14860);
and UO_1971 (O_1971,N_14905,N_14948);
or UO_1972 (O_1972,N_14817,N_14189);
xor UO_1973 (O_1973,N_14260,N_14432);
or UO_1974 (O_1974,N_14398,N_14000);
nor UO_1975 (O_1975,N_14170,N_14735);
xnor UO_1976 (O_1976,N_14634,N_14151);
nor UO_1977 (O_1977,N_14483,N_14802);
xor UO_1978 (O_1978,N_14517,N_14885);
and UO_1979 (O_1979,N_14413,N_14996);
nor UO_1980 (O_1980,N_14665,N_14842);
nand UO_1981 (O_1981,N_14597,N_14556);
or UO_1982 (O_1982,N_14387,N_14653);
nor UO_1983 (O_1983,N_14247,N_14706);
xnor UO_1984 (O_1984,N_14902,N_14488);
and UO_1985 (O_1985,N_14446,N_14470);
xnor UO_1986 (O_1986,N_14183,N_14328);
nor UO_1987 (O_1987,N_14529,N_14293);
or UO_1988 (O_1988,N_14524,N_14119);
nor UO_1989 (O_1989,N_14437,N_14515);
or UO_1990 (O_1990,N_14737,N_14158);
or UO_1991 (O_1991,N_14426,N_14664);
or UO_1992 (O_1992,N_14882,N_14250);
and UO_1993 (O_1993,N_14205,N_14359);
and UO_1994 (O_1994,N_14674,N_14619);
xor UO_1995 (O_1995,N_14068,N_14169);
nor UO_1996 (O_1996,N_14653,N_14794);
and UO_1997 (O_1997,N_14610,N_14901);
xor UO_1998 (O_1998,N_14076,N_14683);
and UO_1999 (O_1999,N_14134,N_14925);
endmodule