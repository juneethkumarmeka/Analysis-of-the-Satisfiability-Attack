module basic_3000_30000_3500_25_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
or U0 (N_0,In_1709,In_1327);
or U1 (N_1,In_7,In_1005);
and U2 (N_2,In_1115,In_491);
or U3 (N_3,In_2870,In_2309);
or U4 (N_4,In_668,In_1239);
and U5 (N_5,In_459,In_1888);
nor U6 (N_6,In_2996,In_1795);
nand U7 (N_7,In_17,In_13);
xor U8 (N_8,In_889,In_1277);
nor U9 (N_9,In_2618,In_1601);
nand U10 (N_10,In_560,In_1539);
or U11 (N_11,In_1272,In_617);
nor U12 (N_12,In_2845,In_2234);
nand U13 (N_13,In_218,In_2276);
nor U14 (N_14,In_481,In_832);
and U15 (N_15,In_1081,In_1054);
xnor U16 (N_16,In_1126,In_2160);
or U17 (N_17,In_672,In_530);
nand U18 (N_18,In_615,In_2075);
nor U19 (N_19,In_1218,In_1171);
xor U20 (N_20,In_574,In_125);
nor U21 (N_21,In_2069,In_2176);
and U22 (N_22,In_1523,In_2694);
nand U23 (N_23,In_1134,In_670);
nand U24 (N_24,In_2366,In_2982);
and U25 (N_25,In_1179,In_1652);
xnor U26 (N_26,In_1075,In_2699);
and U27 (N_27,In_545,In_1465);
xor U28 (N_28,In_980,In_2021);
and U29 (N_29,In_2960,In_1479);
nor U30 (N_30,In_700,In_2641);
nor U31 (N_31,In_922,In_2848);
nor U32 (N_32,In_2859,In_139);
xor U33 (N_33,In_183,In_867);
xnor U34 (N_34,In_859,In_2225);
or U35 (N_35,In_181,In_2296);
nor U36 (N_36,In_418,In_641);
nand U37 (N_37,In_2854,In_2298);
and U38 (N_38,In_2061,In_592);
xnor U39 (N_39,In_1396,In_2408);
or U40 (N_40,In_1278,In_2831);
and U41 (N_41,In_2074,In_2951);
xnor U42 (N_42,In_518,In_444);
and U43 (N_43,In_1297,In_2394);
or U44 (N_44,In_565,In_351);
and U45 (N_45,In_167,In_1873);
nand U46 (N_46,In_886,In_2849);
nand U47 (N_47,In_2168,In_122);
xnor U48 (N_48,In_1003,In_224);
nand U49 (N_49,In_2106,In_1170);
and U50 (N_50,In_1123,In_1289);
xnor U51 (N_51,In_677,In_509);
or U52 (N_52,In_1843,In_1219);
or U53 (N_53,In_2514,In_2112);
nand U54 (N_54,In_2751,In_2059);
and U55 (N_55,In_2524,In_1590);
or U56 (N_56,In_1902,In_1783);
nor U57 (N_57,In_169,In_2601);
or U58 (N_58,In_2447,In_2381);
nand U59 (N_59,In_2661,In_1673);
nand U60 (N_60,In_1603,In_2724);
nand U61 (N_61,In_141,In_1009);
or U62 (N_62,In_875,In_2292);
and U63 (N_63,In_2119,In_1764);
xnor U64 (N_64,In_1934,In_350);
and U65 (N_65,In_730,In_771);
and U66 (N_66,In_2474,In_1419);
nor U67 (N_67,In_1400,In_420);
nor U68 (N_68,In_26,In_748);
and U69 (N_69,In_2738,In_525);
or U70 (N_70,In_877,In_1882);
xnor U71 (N_71,In_1004,In_2765);
or U72 (N_72,In_2277,In_1261);
xnor U73 (N_73,In_2389,In_373);
nor U74 (N_74,In_1267,In_2302);
and U75 (N_75,In_10,In_2020);
and U76 (N_76,In_2100,In_1940);
and U77 (N_77,In_992,In_900);
or U78 (N_78,In_2934,In_2558);
or U79 (N_79,In_655,In_888);
nor U80 (N_80,In_1658,In_1397);
and U81 (N_81,In_1343,In_2241);
xor U82 (N_82,In_2818,In_2926);
nand U83 (N_83,In_1990,In_2211);
nor U84 (N_84,In_1165,In_1384);
or U85 (N_85,In_2792,In_945);
nor U86 (N_86,In_379,In_1513);
nand U87 (N_87,In_2365,In_2864);
nor U88 (N_88,In_507,In_1367);
nand U89 (N_89,In_2534,In_1286);
nand U90 (N_90,In_336,In_2055);
nand U91 (N_91,In_22,In_1895);
or U92 (N_92,In_910,In_1284);
or U93 (N_93,In_1688,In_324);
xor U94 (N_94,In_2651,In_1942);
nand U95 (N_95,In_586,In_61);
nand U96 (N_96,In_281,In_562);
xor U97 (N_97,In_824,In_268);
or U98 (N_98,In_1647,In_413);
nand U99 (N_99,In_1989,In_305);
nand U100 (N_100,In_1352,In_495);
nor U101 (N_101,In_1439,In_2611);
nor U102 (N_102,In_917,In_571);
nand U103 (N_103,In_2930,In_1847);
and U104 (N_104,In_970,In_1329);
nor U105 (N_105,In_2146,In_2598);
xnor U106 (N_106,In_2710,In_1450);
xnor U107 (N_107,In_2489,In_1562);
xnor U108 (N_108,In_1996,In_1095);
or U109 (N_109,In_2925,In_1429);
nor U110 (N_110,In_1721,In_1020);
and U111 (N_111,In_759,In_2583);
nor U112 (N_112,In_925,In_2325);
or U113 (N_113,In_1182,In_2513);
and U114 (N_114,In_2678,In_1470);
nand U115 (N_115,In_1392,In_1924);
nor U116 (N_116,In_1726,In_1798);
xnor U117 (N_117,In_133,In_1089);
nor U118 (N_118,In_1808,In_1270);
xor U119 (N_119,In_544,In_2551);
nor U120 (N_120,In_1860,In_1373);
xor U121 (N_121,In_1130,In_2564);
and U122 (N_122,In_1162,In_750);
xor U123 (N_123,In_2667,In_2689);
xor U124 (N_124,In_703,In_319);
nor U125 (N_125,In_1637,In_393);
or U126 (N_126,In_650,In_1509);
nand U127 (N_127,In_2014,In_2334);
or U128 (N_128,In_2909,In_942);
nor U129 (N_129,In_1443,In_1623);
nand U130 (N_130,In_1019,In_410);
nand U131 (N_131,In_1803,In_1281);
xor U132 (N_132,In_816,In_470);
or U133 (N_133,In_2432,In_2987);
nand U134 (N_134,In_483,In_2581);
nand U135 (N_135,In_430,In_463);
nand U136 (N_136,In_2090,In_1168);
nor U137 (N_137,In_1410,In_101);
nand U138 (N_138,In_2714,In_2361);
nand U139 (N_139,In_2668,In_2826);
xnor U140 (N_140,In_12,In_2774);
and U141 (N_141,In_1264,In_755);
nand U142 (N_142,In_1920,In_2753);
or U143 (N_143,In_515,In_520);
nor U144 (N_144,In_2655,In_2913);
or U145 (N_145,In_2041,In_782);
and U146 (N_146,In_1935,In_2985);
and U147 (N_147,In_2877,In_1156);
nand U148 (N_148,In_1083,In_2585);
nand U149 (N_149,In_1648,In_2786);
xnor U150 (N_150,In_608,In_954);
nor U151 (N_151,In_2917,In_1665);
nand U152 (N_152,In_2093,In_2261);
nand U153 (N_153,In_1306,In_2284);
xnor U154 (N_154,In_557,In_2507);
or U155 (N_155,In_2700,In_1525);
xnor U156 (N_156,In_1823,In_1300);
nand U157 (N_157,In_1697,In_317);
nand U158 (N_158,In_1377,In_477);
or U159 (N_159,In_708,In_1448);
nand U160 (N_160,In_1187,In_433);
xnor U161 (N_161,In_732,In_2869);
xnor U162 (N_162,In_1919,In_778);
or U163 (N_163,In_1326,In_861);
nor U164 (N_164,In_1030,In_665);
and U165 (N_165,In_1451,In_1246);
nand U166 (N_166,In_1540,In_1322);
nor U167 (N_167,In_62,In_2498);
nand U168 (N_168,In_689,In_95);
and U169 (N_169,In_2442,In_2073);
nor U170 (N_170,In_2331,In_1793);
nor U171 (N_171,In_2265,In_607);
and U172 (N_172,In_1129,In_381);
and U173 (N_173,In_362,In_331);
or U174 (N_174,In_2042,In_1640);
xnor U175 (N_175,In_937,In_1946);
xor U176 (N_176,In_831,In_588);
and U177 (N_177,In_146,In_2793);
and U178 (N_178,In_2556,In_763);
and U179 (N_179,In_80,In_2769);
xor U180 (N_180,In_2030,In_1039);
nand U181 (N_181,In_2755,In_929);
nand U182 (N_182,In_2883,In_2255);
nand U183 (N_183,In_1131,In_2048);
nor U184 (N_184,In_1700,In_2892);
or U185 (N_185,In_1045,In_223);
xnor U186 (N_186,In_2968,In_996);
and U187 (N_187,In_1679,In_920);
xor U188 (N_188,In_2579,In_1690);
nand U189 (N_189,In_2227,In_845);
or U190 (N_190,In_448,In_924);
nand U191 (N_191,In_1008,In_153);
and U192 (N_192,In_2981,In_551);
xor U193 (N_193,In_86,In_364);
and U194 (N_194,In_2811,In_713);
nor U195 (N_195,In_871,In_485);
nand U196 (N_196,In_2533,In_1041);
or U197 (N_197,In_1070,In_1909);
nor U198 (N_198,In_1887,In_2025);
xnor U199 (N_199,In_2313,In_538);
or U200 (N_200,In_1176,In_180);
or U201 (N_201,In_243,In_63);
nor U202 (N_202,In_188,In_1702);
nor U203 (N_203,In_603,In_734);
nor U204 (N_204,In_1633,In_220);
or U205 (N_205,In_1038,In_2123);
nand U206 (N_206,In_72,In_1107);
xnor U207 (N_207,In_1093,In_583);
xor U208 (N_208,In_107,In_165);
and U209 (N_209,In_812,In_2310);
or U210 (N_210,In_1105,In_2129);
and U211 (N_211,In_1643,In_2382);
and U212 (N_212,In_2664,In_1617);
xnor U213 (N_213,In_24,In_2721);
nor U214 (N_214,In_2120,In_284);
xor U215 (N_215,In_2695,In_2910);
xnor U216 (N_216,In_452,In_1893);
nand U217 (N_217,In_1196,In_118);
nand U218 (N_218,In_1422,In_1122);
nor U219 (N_219,In_1576,In_994);
or U220 (N_220,In_291,In_2995);
or U221 (N_221,In_2326,In_406);
xnor U222 (N_222,In_1172,In_2360);
or U223 (N_223,In_593,In_175);
nand U224 (N_224,In_2941,In_457);
or U225 (N_225,In_805,In_997);
nand U226 (N_226,In_1490,In_2253);
and U227 (N_227,In_2530,In_814);
nor U228 (N_228,In_2687,In_2392);
and U229 (N_229,In_981,In_2399);
and U230 (N_230,In_2777,In_415);
nor U231 (N_231,In_2354,In_1758);
and U232 (N_232,In_2003,In_2882);
xnor U233 (N_233,In_844,In_642);
xnor U234 (N_234,In_1481,In_1120);
nor U235 (N_235,In_640,In_1427);
or U236 (N_236,In_550,In_913);
and U237 (N_237,In_1420,In_1453);
nand U238 (N_238,In_1280,In_2992);
xor U239 (N_239,In_1828,In_2923);
and U240 (N_240,In_1982,In_1575);
and U241 (N_241,In_2608,In_2084);
or U242 (N_242,In_1854,In_850);
or U243 (N_243,In_348,In_2580);
nor U244 (N_244,In_943,In_1254);
nor U245 (N_245,In_332,In_1613);
or U246 (N_246,In_436,In_1356);
and U247 (N_247,In_2081,In_1699);
and U248 (N_248,In_2764,In_2565);
and U249 (N_249,In_1664,In_772);
and U250 (N_250,In_659,In_589);
xnor U251 (N_251,In_2949,In_32);
nor U252 (N_252,In_721,In_1628);
or U253 (N_253,In_2018,In_1189);
and U254 (N_254,In_1458,In_811);
or U255 (N_255,In_2957,In_630);
or U256 (N_256,In_1884,In_2138);
nor U257 (N_257,In_962,In_1110);
xnor U258 (N_258,In_2140,In_335);
or U259 (N_259,In_2975,In_1135);
or U260 (N_260,In_1723,In_2602);
nor U261 (N_261,In_2756,In_1118);
or U262 (N_262,In_2890,In_2544);
xnor U263 (N_263,In_1761,In_1524);
xor U264 (N_264,In_380,In_2575);
or U265 (N_265,In_693,In_254);
xor U266 (N_266,In_446,In_1475);
or U267 (N_267,In_353,In_534);
nor U268 (N_268,In_2871,In_1896);
and U269 (N_269,In_1065,In_2133);
xnor U270 (N_270,In_978,In_2973);
nand U271 (N_271,In_387,In_756);
and U272 (N_272,In_241,In_621);
nand U273 (N_273,In_1032,In_843);
nor U274 (N_274,In_2062,In_1139);
nand U275 (N_275,In_308,In_1202);
nand U276 (N_276,In_1132,In_2395);
nor U277 (N_277,In_2156,In_1975);
nand U278 (N_278,In_880,In_1413);
or U279 (N_279,In_128,In_2902);
xor U280 (N_280,In_320,In_1023);
nand U281 (N_281,In_625,In_316);
or U282 (N_282,In_2099,In_293);
xnor U283 (N_283,In_602,In_1432);
nor U284 (N_284,In_938,In_2494);
nor U285 (N_285,In_271,In_2587);
xor U286 (N_286,In_178,In_1245);
nand U287 (N_287,In_2315,In_493);
and U288 (N_288,In_1668,In_1155);
nor U289 (N_289,In_1710,In_70);
nand U290 (N_290,In_2485,In_25);
nand U291 (N_291,In_304,In_1500);
nor U292 (N_292,In_769,In_2780);
and U293 (N_293,In_1784,In_1476);
xor U294 (N_294,In_1712,In_1813);
nor U295 (N_295,In_1376,In_573);
xor U296 (N_296,In_842,In_653);
xnor U297 (N_297,In_907,In_522);
and U298 (N_298,In_1301,In_1050);
nand U299 (N_299,In_1347,In_2116);
nor U300 (N_300,In_2184,In_940);
nor U301 (N_301,In_2137,In_1133);
nand U302 (N_302,In_2343,In_911);
or U303 (N_303,In_1591,In_2752);
or U304 (N_304,In_91,In_1938);
or U305 (N_305,In_2153,In_2952);
or U306 (N_306,In_174,In_927);
xor U307 (N_307,In_2159,In_2506);
or U308 (N_308,In_626,In_89);
or U309 (N_309,In_1404,In_1738);
nor U310 (N_310,In_1206,In_777);
nand U311 (N_311,In_510,In_1011);
and U312 (N_312,In_2490,In_2068);
xnor U313 (N_313,In_142,In_1497);
or U314 (N_314,In_930,In_338);
and U315 (N_315,In_1145,In_2427);
and U316 (N_316,In_2672,In_2098);
xor U317 (N_317,In_2496,In_2851);
and U318 (N_318,In_853,In_2188);
or U319 (N_319,In_1158,In_1111);
and U320 (N_320,In_2911,In_2164);
or U321 (N_321,In_2145,In_1867);
and U322 (N_322,In_2701,In_2535);
xor U323 (N_323,In_599,In_1826);
or U324 (N_324,In_2875,In_2237);
and U325 (N_325,In_1234,In_1889);
or U326 (N_326,In_801,In_2036);
nand U327 (N_327,In_2666,In_115);
nor U328 (N_328,In_377,In_1407);
nor U329 (N_329,In_1203,In_1739);
xnor U330 (N_330,In_1510,In_2559);
nand U331 (N_331,In_2333,In_1611);
nand U332 (N_332,In_365,In_1563);
or U333 (N_333,In_2725,In_256);
and U334 (N_334,In_94,In_1102);
xor U335 (N_335,In_1961,In_2676);
nor U336 (N_336,In_2621,In_1237);
nand U337 (N_337,In_982,In_2595);
and U338 (N_338,In_1211,In_2903);
nand U339 (N_339,In_793,In_2047);
or U340 (N_340,In_1389,In_93);
and U341 (N_341,In_1899,In_2460);
and U342 (N_342,In_674,In_1350);
nor U343 (N_343,In_233,In_1516);
or U344 (N_344,In_2192,In_2572);
or U345 (N_345,In_227,In_2974);
nand U346 (N_346,In_1268,In_1964);
nor U347 (N_347,In_854,In_301);
xnor U348 (N_348,In_2972,In_1883);
nand U349 (N_349,In_1332,In_2609);
and U350 (N_350,In_2401,In_237);
nor U351 (N_351,In_2749,In_946);
or U352 (N_352,In_472,In_2379);
and U353 (N_353,In_2202,In_97);
nand U354 (N_354,In_18,In_15);
and U355 (N_355,In_1214,In_2207);
nand U356 (N_356,In_2005,In_2050);
nor U357 (N_357,In_2767,In_2658);
xnor U358 (N_358,In_2300,In_2993);
xnor U359 (N_359,In_337,In_1052);
xnor U360 (N_360,In_1460,In_952);
nor U361 (N_361,In_2825,In_575);
nand U362 (N_362,In_1971,In_326);
nor U363 (N_363,In_2169,In_1747);
nor U364 (N_364,In_612,In_2136);
xnor U365 (N_365,In_1082,In_1431);
and U366 (N_366,In_333,In_422);
nand U367 (N_367,In_1185,In_553);
and U368 (N_368,In_129,In_2683);
nor U369 (N_369,In_487,In_2435);
xor U370 (N_370,In_394,In_1667);
or U371 (N_371,In_245,In_1468);
xor U372 (N_372,In_1733,In_480);
or U373 (N_373,In_2008,In_1414);
and U374 (N_374,In_2088,In_1531);
nand U375 (N_375,In_837,In_983);
nor U376 (N_376,In_1051,In_2865);
nand U377 (N_377,In_2548,In_2696);
or U378 (N_378,In_53,In_628);
and U379 (N_379,In_1771,In_2318);
or U380 (N_380,In_849,In_2293);
and U381 (N_381,In_1535,In_2686);
nand U382 (N_382,In_2278,In_310);
nor U383 (N_383,In_2004,In_2492);
xor U384 (N_384,In_1782,In_1147);
xor U385 (N_385,In_2876,In_1068);
xor U386 (N_386,In_2553,In_357);
xor U387 (N_387,In_2628,In_1066);
or U388 (N_388,In_2180,In_2735);
or U389 (N_389,In_385,In_535);
nor U390 (N_390,In_706,In_2627);
xnor U391 (N_391,In_1811,In_1342);
xnor U392 (N_392,In_2531,In_531);
and U393 (N_393,In_2409,In_1303);
or U394 (N_394,In_1112,In_2604);
xnor U395 (N_395,In_2896,In_1402);
and U396 (N_396,In_416,In_2148);
and U397 (N_397,In_701,In_2644);
and U398 (N_398,In_2054,In_1862);
or U399 (N_399,In_1520,In_1840);
or U400 (N_400,In_2626,In_754);
and U401 (N_401,In_1114,In_151);
and U402 (N_402,In_2281,In_926);
xor U403 (N_403,In_388,In_2887);
xor U404 (N_404,In_1193,In_2712);
or U405 (N_405,In_1682,In_1908);
nor U406 (N_406,In_2776,In_2779);
nor U407 (N_407,In_2240,In_2692);
nand U408 (N_408,In_1334,In_1742);
or U409 (N_409,In_2590,In_2357);
and U410 (N_410,In_66,In_1007);
nor U411 (N_411,In_2105,In_1618);
or U412 (N_412,In_1948,In_580);
nand U413 (N_413,In_887,In_1756);
nor U414 (N_414,In_2470,In_699);
xor U415 (N_415,In_1596,In_2436);
or U416 (N_416,In_2542,In_705);
xnor U417 (N_417,In_2841,In_1670);
nor U418 (N_418,In_2491,In_2763);
nor U419 (N_419,In_1541,In_1829);
and U420 (N_420,In_1417,In_2322);
or U421 (N_421,In_975,In_1984);
or U422 (N_422,In_2049,In_2258);
or U423 (N_423,In_1049,In_454);
nor U424 (N_424,In_55,In_918);
nor U425 (N_425,In_2720,In_1127);
nor U426 (N_426,In_2107,In_3);
nand U427 (N_427,In_1955,In_1530);
nand U428 (N_428,In_1148,In_51);
xor U429 (N_429,In_902,In_1341);
or U430 (N_430,In_2945,In_1282);
or U431 (N_431,In_1732,In_2546);
nor U432 (N_432,In_2250,In_1188);
nand U433 (N_433,In_275,In_1063);
and U434 (N_434,In_1383,In_623);
or U435 (N_435,In_1824,In_2739);
and U436 (N_436,In_1124,In_1988);
nor U437 (N_437,In_1814,In_2495);
xnor U438 (N_438,In_1226,In_2171);
xor U439 (N_439,In_1416,In_2933);
nor U440 (N_440,In_2532,In_1040);
xor U441 (N_441,In_1967,In_1962);
xor U442 (N_442,In_1999,In_741);
xnor U443 (N_443,In_2196,In_846);
and U444 (N_444,In_2209,In_395);
nor U445 (N_445,In_1436,In_559);
or U446 (N_446,In_1797,In_2804);
nand U447 (N_447,In_2231,In_2963);
nor U448 (N_448,In_1177,In_2833);
xnor U449 (N_449,In_198,In_1691);
or U450 (N_450,In_2259,In_2279);
or U451 (N_451,In_2126,In_1842);
nand U452 (N_452,In_695,In_1222);
xnor U453 (N_453,In_2102,In_1609);
or U454 (N_454,In_569,In_2956);
and U455 (N_455,In_2390,In_1689);
nand U456 (N_456,In_1517,In_64);
or U457 (N_457,In_523,In_2501);
and U458 (N_458,In_1495,In_1493);
or U459 (N_459,In_2784,In_568);
or U460 (N_460,In_2806,In_2033);
and U461 (N_461,In_78,In_2596);
nor U462 (N_462,In_2404,In_1323);
and U463 (N_463,In_1773,In_638);
nor U464 (N_464,In_1805,In_401);
and U465 (N_465,In_438,In_1354);
or U466 (N_466,In_903,In_2271);
and U467 (N_467,In_479,In_723);
and U468 (N_468,In_691,In_50);
xor U469 (N_469,In_2367,In_370);
and U470 (N_470,In_2519,In_2566);
and U471 (N_471,In_2812,In_1504);
or U472 (N_472,In_2264,In_1053);
nor U473 (N_473,In_2997,In_1152);
nor U474 (N_474,In_953,In_497);
or U475 (N_475,In_2682,In_766);
or U476 (N_476,In_1026,In_2411);
xor U477 (N_477,In_2150,In_2465);
nand U478 (N_478,In_1308,In_1548);
nor U479 (N_479,In_1256,In_1046);
nand U480 (N_480,In_265,In_1084);
and U481 (N_481,In_1208,In_2425);
xnor U482 (N_482,In_2157,In_1074);
nand U483 (N_483,In_947,In_2472);
and U484 (N_484,In_720,In_2884);
nand U485 (N_485,In_899,In_971);
and U486 (N_486,In_400,In_1511);
nor U487 (N_487,In_2031,In_154);
nor U488 (N_488,In_1437,In_1358);
or U489 (N_489,In_1273,In_360);
nand U490 (N_490,In_2424,In_989);
nand U491 (N_491,In_1939,In_230);
xor U492 (N_492,In_1482,In_908);
and U493 (N_493,In_684,In_468);
and U494 (N_494,In_1477,In_736);
nand U495 (N_495,In_1380,In_1190);
nand U496 (N_496,In_2221,In_1015);
xnor U497 (N_497,In_41,In_307);
and U498 (N_498,In_1672,In_773);
xnor U499 (N_499,In_591,In_1674);
nand U500 (N_500,In_313,In_1987);
and U501 (N_501,In_2836,In_1715);
nand U502 (N_502,In_636,In_2719);
xor U503 (N_503,In_2166,In_919);
or U504 (N_504,In_403,In_2652);
and U505 (N_505,In_1794,In_325);
nor U506 (N_506,In_2257,In_2539);
or U507 (N_507,In_2455,In_2128);
xor U508 (N_508,In_2305,In_1762);
and U509 (N_509,In_2374,In_936);
xor U510 (N_510,In_1398,In_2790);
and U511 (N_511,In_2729,In_1599);
nand U512 (N_512,In_1928,In_2600);
and U513 (N_513,In_711,In_2311);
nor U514 (N_514,In_392,In_1901);
and U515 (N_515,In_2966,In_1631);
or U516 (N_516,In_2103,In_2170);
nor U517 (N_517,In_46,In_2267);
or U518 (N_518,In_2175,In_669);
xnor U519 (N_519,In_1311,In_1386);
xnor U520 (N_520,In_1832,In_1877);
or U521 (N_521,In_543,In_915);
nor U522 (N_522,In_537,In_456);
xnor U523 (N_523,In_692,In_506);
nor U524 (N_524,In_2560,In_323);
and U525 (N_525,In_2203,In_1036);
xor U526 (N_526,In_1692,In_1514);
xnor U527 (N_527,In_2282,In_1037);
nand U528 (N_528,In_1163,In_222);
nor U529 (N_529,In_1447,In_897);
or U530 (N_530,In_2019,In_1954);
and U531 (N_531,In_808,In_471);
or U532 (N_532,In_2955,In_2251);
xnor U533 (N_533,In_383,In_2718);
and U534 (N_534,In_1681,In_1157);
nor U535 (N_535,In_654,In_807);
nand U536 (N_536,In_2213,In_2289);
nand U537 (N_537,In_1079,In_302);
or U538 (N_538,In_475,In_9);
nand U539 (N_539,In_2372,In_1344);
nor U540 (N_540,In_2619,In_156);
and U541 (N_541,In_2707,In_2448);
nand U542 (N_542,In_1191,In_1166);
nor U543 (N_543,In_2383,In_2868);
or U544 (N_544,In_247,In_2517);
nand U545 (N_545,In_541,In_2867);
xor U546 (N_546,In_2642,In_611);
nor U547 (N_547,In_687,In_2303);
and U548 (N_548,In_1622,In_1047);
nor U549 (N_549,In_680,In_2829);
or U550 (N_550,In_1986,In_134);
nor U551 (N_551,In_2746,In_127);
nand U552 (N_552,In_2403,In_2028);
xnor U553 (N_553,In_817,In_2813);
or U554 (N_554,In_2866,In_1200);
xnor U555 (N_555,In_1428,In_1283);
nor U556 (N_556,In_1991,In_376);
nand U557 (N_557,In_2239,In_1331);
xnor U558 (N_558,In_82,In_2736);
xnor U559 (N_559,In_2743,In_2388);
or U560 (N_560,In_458,In_839);
nor U561 (N_561,In_2022,In_1553);
or U562 (N_562,In_1629,In_2768);
or U563 (N_563,In_1293,In_1287);
and U564 (N_564,In_1248,In_2371);
and U565 (N_565,In_2198,In_197);
or U566 (N_566,In_1789,In_2416);
or U567 (N_567,In_933,In_1255);
xor U568 (N_568,In_106,In_841);
and U569 (N_569,In_896,In_1977);
and U570 (N_570,In_882,In_1335);
or U571 (N_571,In_1748,In_2529);
or U572 (N_572,In_2087,In_140);
xnor U573 (N_573,In_524,In_789);
or U574 (N_574,In_1890,In_1641);
xor U575 (N_575,In_1932,In_2741);
and U576 (N_576,In_2557,In_2339);
xnor U577 (N_577,In_2893,In_1364);
and U578 (N_578,In_2242,In_1542);
nor U579 (N_579,In_1199,In_1846);
nor U580 (N_580,In_2344,In_2384);
or U581 (N_581,In_1173,In_273);
nand U582 (N_582,In_2562,In_1571);
and U583 (N_583,In_546,In_199);
nand U584 (N_584,In_2713,In_2935);
nor U585 (N_585,In_2861,In_116);
nor U586 (N_586,In_2063,In_1309);
nand U587 (N_587,In_1405,In_539);
or U588 (N_588,In_1777,In_2525);
and U589 (N_589,In_757,In_296);
nand U590 (N_590,In_2338,In_2431);
and U591 (N_591,In_1625,In_1325);
nand U592 (N_592,In_2832,In_2591);
xnor U593 (N_593,In_285,In_964);
and U594 (N_594,In_2838,In_1606);
and U595 (N_595,In_2944,In_725);
xor U596 (N_596,In_207,In_606);
nor U597 (N_597,In_144,In_604);
and U598 (N_598,In_1614,In_1101);
or U599 (N_599,In_1391,In_1552);
xor U600 (N_600,In_2574,In_1201);
nand U601 (N_601,In_594,In_1970);
or U602 (N_602,In_1607,In_2194);
and U603 (N_603,In_27,In_610);
nand U604 (N_604,In_372,In_1328);
nand U605 (N_605,In_123,In_2178);
nor U606 (N_606,In_719,In_928);
xnor U607 (N_607,In_1624,In_1589);
nor U608 (N_608,In_2670,In_921);
nand U609 (N_609,In_663,In_173);
or U610 (N_610,In_157,In_1837);
nor U611 (N_611,In_2449,In_2733);
nand U612 (N_612,In_1069,In_1766);
nand U613 (N_613,In_1903,In_1957);
or U614 (N_614,In_1770,In_2060);
xor U615 (N_615,In_1711,In_1247);
xor U616 (N_616,In_1969,In_2703);
xnor U617 (N_617,In_2316,In_1820);
nand U618 (N_618,In_2364,In_2852);
nand U619 (N_619,In_2726,In_2410);
and U620 (N_620,In_2466,In_1894);
nand U621 (N_621,In_1236,In_83);
nand U622 (N_622,In_661,In_2032);
or U623 (N_623,In_1515,In_1258);
or U624 (N_624,In_2285,In_1834);
nor U625 (N_625,In_2254,In_958);
nor U626 (N_626,In_2842,In_1088);
nor U627 (N_627,In_1243,In_1098);
nor U628 (N_628,In_1737,In_2874);
xor U629 (N_629,In_710,In_765);
nand U630 (N_630,In_821,In_1409);
xor U631 (N_631,In_1638,In_1149);
nand U632 (N_632,In_797,In_2860);
nor U633 (N_633,In_2352,In_405);
xor U634 (N_634,In_2846,In_354);
nand U635 (N_635,In_1103,In_865);
nor U636 (N_636,In_2853,In_2272);
nor U637 (N_637,In_2079,In_467);
xnor U638 (N_638,In_363,In_966);
nand U639 (N_639,In_1109,In_90);
and U640 (N_640,In_2205,In_1259);
nor U641 (N_641,In_1566,In_2369);
nand U642 (N_642,In_1319,In_823);
nand U643 (N_643,In_2487,In_934);
and U644 (N_644,In_2187,In_1288);
xor U645 (N_645,In_311,In_1872);
nand U646 (N_646,In_246,In_2688);
nand U647 (N_647,In_1724,In_1992);
nand U648 (N_648,In_1374,In_1312);
nand U649 (N_649,In_1313,In_2504);
xnor U650 (N_650,In_104,In_1701);
nand U651 (N_651,In_212,In_2734);
and U652 (N_652,In_427,In_2070);
and U653 (N_653,In_2922,In_2034);
or U654 (N_654,In_1677,In_662);
and U655 (N_655,In_182,In_2937);
nor U656 (N_656,In_2467,In_2914);
and U657 (N_657,In_526,In_1615);
nand U658 (N_658,In_1687,In_2775);
xnor U659 (N_659,In_2181,In_1743);
and U660 (N_660,In_1252,In_657);
and U661 (N_661,In_1584,In_1557);
nand U662 (N_662,In_2820,In_1406);
xor U663 (N_663,In_1630,In_1445);
and U664 (N_664,In_1097,In_2680);
nand U665 (N_665,In_1,In_124);
or U666 (N_666,In_2708,In_2351);
and U667 (N_667,In_2478,In_2040);
nand U668 (N_668,In_1180,In_1809);
xor U669 (N_669,In_419,In_2165);
or U670 (N_670,In_1534,In_2210);
nor U671 (N_671,In_1663,In_1787);
and U672 (N_672,In_595,In_1852);
nor U673 (N_673,In_2064,In_2214);
nor U674 (N_674,In_624,In_1175);
nor U675 (N_675,In_1642,In_1583);
nor U676 (N_676,In_1498,In_4);
xor U677 (N_677,In_549,In_1616);
or U678 (N_678,In_217,In_1561);
or U679 (N_679,In_498,In_813);
nor U680 (N_680,In_1806,In_601);
nand U681 (N_681,In_2398,In_1943);
nand U682 (N_682,In_2010,In_1716);
nor U683 (N_683,In_261,In_629);
and U684 (N_684,In_1608,In_453);
nor U685 (N_685,In_512,In_2052);
or U686 (N_686,In_170,In_959);
or U687 (N_687,In_1522,In_1904);
xnor U688 (N_688,In_1930,In_2023);
nor U689 (N_689,In_205,In_2009);
and U690 (N_690,In_2905,In_267);
nand U691 (N_691,In_1915,In_2894);
xnor U692 (N_692,In_532,In_2665);
nor U693 (N_693,In_132,In_2306);
or U694 (N_694,In_2057,In_819);
or U695 (N_695,In_378,In_1138);
and U696 (N_696,In_890,In_648);
or U697 (N_697,In_2855,In_1704);
xnor U698 (N_698,In_1435,In_1022);
or U699 (N_699,In_2946,In_1159);
or U700 (N_700,In_1627,In_1244);
or U701 (N_701,In_1178,In_2348);
and U702 (N_702,In_1595,In_1555);
xor U703 (N_703,In_2759,In_359);
and U704 (N_704,In_386,In_2412);
or U705 (N_705,In_2163,In_961);
and U706 (N_706,In_1951,In_2794);
or U707 (N_707,In_2066,In_228);
nor U708 (N_708,In_2457,In_2263);
and U709 (N_709,In_67,In_2236);
and U710 (N_710,In_1230,In_235);
and U711 (N_711,In_2603,In_1656);
or U712 (N_712,In_678,In_1018);
nor U713 (N_713,In_547,In_2452);
nor U714 (N_714,In_465,In_596);
nor U715 (N_715,In_1080,In_2578);
or U716 (N_716,In_1558,In_1772);
nor U717 (N_717,In_1666,In_898);
xnor U718 (N_718,In_2773,In_2260);
nand U719 (N_719,In_249,In_2002);
nand U720 (N_720,In_114,In_2536);
nand U721 (N_721,In_1918,In_2657);
and U722 (N_722,In_234,In_216);
xnor U723 (N_723,In_1947,In_1212);
nor U724 (N_724,In_2545,In_1831);
or U725 (N_725,In_1734,In_505);
xnor U726 (N_726,In_435,In_282);
nor U727 (N_727,In_113,In_2684);
nand U728 (N_728,In_1321,In_679);
or U729 (N_729,In_2901,In_2638);
xor U730 (N_730,In_1366,In_499);
and U731 (N_731,In_74,In_770);
nand U732 (N_732,In_822,In_1729);
nand U733 (N_733,In_633,In_344);
xnor U734 (N_734,In_2461,In_201);
nand U735 (N_735,In_20,In_2340);
and U736 (N_736,In_1705,In_870);
or U737 (N_737,In_1819,In_272);
xnor U738 (N_738,In_847,In_1119);
xor U739 (N_739,In_1337,In_1586);
nor U740 (N_740,In_2801,In_968);
xnor U741 (N_741,In_1480,In_1262);
nor U742 (N_742,In_1644,In_2715);
xor U743 (N_743,In_2858,In_1866);
nand U744 (N_744,In_1464,In_1001);
nor U745 (N_745,In_731,In_2942);
xor U746 (N_746,In_1478,In_2206);
nand U747 (N_747,In_2445,In_1916);
nor U748 (N_748,In_1512,In_484);
or U749 (N_749,In_166,In_799);
and U750 (N_750,In_162,In_294);
and U751 (N_751,In_1198,In_1499);
nor U752 (N_752,In_2570,In_2347);
nor U753 (N_753,In_109,In_2584);
and U754 (N_754,In_191,In_2463);
and U755 (N_755,In_1229,In_828);
and U756 (N_756,In_1696,In_2373);
or U757 (N_757,In_2249,In_2423);
nor U758 (N_758,In_963,In_1610);
or U759 (N_759,In_1953,In_30);
and U760 (N_760,In_984,In_794);
nor U761 (N_761,In_1736,In_2108);
xor U762 (N_762,In_1592,In_1298);
nor U763 (N_763,In_1290,In_2477);
or U764 (N_764,In_2230,In_298);
or U765 (N_765,In_1501,In_866);
nand U766 (N_766,In_1839,In_2931);
or U767 (N_767,In_2969,In_1502);
or U768 (N_768,In_627,In_675);
and U769 (N_769,In_1421,In_941);
or U770 (N_770,In_1204,In_321);
and U771 (N_771,In_779,In_1876);
and U772 (N_772,In_834,In_367);
xor U773 (N_773,In_1830,In_2748);
nor U774 (N_774,In_2149,In_1440);
xor U775 (N_775,In_2795,In_2991);
xnor U776 (N_776,In_21,In_1355);
nand U777 (N_777,In_2096,In_2247);
nand U778 (N_778,In_631,In_1161);
and U779 (N_779,In_1880,In_791);
nand U780 (N_780,In_2948,In_441);
nand U781 (N_781,In_567,In_503);
xnor U782 (N_782,In_258,In_862);
xnor U783 (N_783,In_555,In_2229);
xor U784 (N_784,In_1661,In_1574);
and U785 (N_785,In_1570,In_577);
nor U786 (N_786,In_1485,In_2599);
and U787 (N_787,In_2441,In_1043);
nor U788 (N_788,In_1024,In_163);
nor U789 (N_789,In_2244,In_96);
nor U790 (N_790,In_2189,In_2437);
and U791 (N_791,In_312,In_1154);
and U792 (N_792,In_1295,In_2907);
or U793 (N_793,In_1660,In_2920);
nor U794 (N_794,In_851,In_1639);
xnor U795 (N_795,In_2197,In_2006);
nand U796 (N_796,In_2800,In_2232);
xor U797 (N_797,In_2762,In_960);
xnor U798 (N_798,In_375,In_2336);
and U799 (N_799,In_211,In_974);
and U800 (N_800,In_2671,In_1042);
xnor U801 (N_801,In_1654,In_391);
xnor U802 (N_802,In_909,In_1441);
nor U803 (N_803,In_2863,In_576);
nor U804 (N_804,In_2827,In_1634);
nand U805 (N_805,In_1362,In_1551);
and U806 (N_806,In_995,In_1233);
nor U807 (N_807,In_2433,In_548);
or U808 (N_808,In_554,In_2426);
or U809 (N_809,In_1096,In_2377);
nor U810 (N_810,In_1220,In_2711);
nor U811 (N_811,In_972,In_1740);
xor U812 (N_812,In_1597,In_43);
or U813 (N_813,In_570,In_42);
xor U814 (N_814,In_1302,In_2450);
nand U815 (N_815,In_1678,In_1578);
xnor U816 (N_816,In_2056,In_262);
nor U817 (N_817,In_2702,In_1529);
xnor U818 (N_818,In_1184,In_2502);
xor U819 (N_819,In_2130,In_1452);
or U820 (N_820,In_2899,In_2454);
xnor U821 (N_821,In_1385,In_632);
xor U822 (N_822,In_2509,In_2622);
xnor U823 (N_823,In_1195,In_73);
nand U824 (N_824,In_2245,In_411);
and U825 (N_825,In_451,In_1750);
nand U826 (N_826,In_664,In_511);
xor U827 (N_827,In_2015,In_48);
nand U828 (N_828,In_2679,In_840);
and U829 (N_829,In_1532,In_2589);
nor U830 (N_830,In_1263,In_2625);
nand U831 (N_831,In_208,In_742);
nand U832 (N_832,In_1857,In_2757);
xor U833 (N_833,In_1454,In_192);
nor U834 (N_834,In_1296,In_744);
and U835 (N_835,In_1333,In_774);
or U836 (N_836,In_796,In_280);
and U837 (N_837,In_2610,In_110);
nor U838 (N_838,In_2824,In_478);
and U839 (N_839,In_1993,In_1058);
nand U840 (N_840,In_2071,In_329);
nor U841 (N_841,In_2669,In_2029);
nor U842 (N_842,In_149,In_1067);
nand U843 (N_843,In_1593,In_1708);
nor U844 (N_844,In_2508,In_1816);
or U845 (N_845,In_827,In_1881);
or U846 (N_846,In_2370,In_2990);
xnor U847 (N_847,In_1317,In_2730);
xor U848 (N_848,In_120,In_1061);
nand U849 (N_849,In_1340,In_1885);
nor U850 (N_850,In_2983,In_800);
nor U851 (N_851,In_1550,In_155);
and U852 (N_852,In_776,In_203);
nand U853 (N_853,In_2543,In_103);
and U854 (N_854,In_540,In_1848);
or U855 (N_855,In_1128,In_2518);
and U856 (N_856,In_826,In_815);
and U857 (N_857,In_0,In_260);
or U858 (N_858,In_1718,In_99);
nand U859 (N_859,In_2526,In_2592);
or U860 (N_860,In_269,In_2233);
nand U861 (N_861,In_426,In_160);
nor U862 (N_862,In_2550,In_1925);
nand U863 (N_863,In_1330,In_1849);
nor U864 (N_864,In_2782,In_2132);
and U865 (N_865,In_2139,In_656);
nand U866 (N_866,In_751,In_449);
or U867 (N_867,In_2319,In_2110);
nor U868 (N_868,In_2633,In_204);
xnor U869 (N_869,In_2101,In_1979);
or U870 (N_870,In_2885,In_2798);
nor U871 (N_871,In_990,In_696);
nand U872 (N_872,In_2078,In_1815);
nor U873 (N_873,In_2976,In_709);
nand U874 (N_874,In_1968,In_829);
nand U875 (N_875,In_1348,In_1151);
nand U876 (N_876,In_804,In_901);
nor U877 (N_877,In_2629,In_1792);
xor U878 (N_878,In_1463,In_469);
and U879 (N_879,In_398,In_1956);
nor U880 (N_880,In_1717,In_286);
nand U881 (N_881,In_11,In_1547);
and U882 (N_882,In_2880,In_1744);
and U883 (N_883,In_1013,In_1810);
nand U884 (N_884,In_8,In_1473);
nor U885 (N_885,In_407,In_1357);
nor U886 (N_886,In_1818,In_1073);
xor U887 (N_887,In_179,In_2770);
or U888 (N_888,In_514,In_1411);
or U889 (N_889,In_87,In_1778);
and U890 (N_890,In_2677,In_1310);
or U891 (N_891,In_752,In_1213);
xor U892 (N_892,In_1242,In_1653);
and U893 (N_893,In_1433,In_2396);
or U894 (N_894,In_161,In_948);
nor U895 (N_895,In_2443,In_743);
or U896 (N_896,In_1868,In_1741);
xor U897 (N_897,In_2632,In_1141);
nand U898 (N_898,In_1240,In_306);
nand U899 (N_899,In_579,In_1594);
nor U900 (N_900,In_685,In_2097);
nand U901 (N_901,In_973,In_2481);
or U902 (N_902,In_496,In_892);
nand U903 (N_903,In_1227,In_283);
nand U904 (N_904,In_988,In_1906);
nor U905 (N_905,In_707,In_787);
xnor U906 (N_906,In_2947,In_2881);
nor U907 (N_907,In_242,In_878);
and U908 (N_908,In_1423,In_1879);
or U909 (N_909,In_2067,In_450);
or U910 (N_910,In_374,In_2341);
xnor U911 (N_911,In_1192,In_2516);
and U912 (N_912,In_2637,In_1760);
xnor U913 (N_913,In_647,In_2299);
or U914 (N_914,In_171,In_1064);
xnor U915 (N_915,In_2402,In_1949);
xnor U916 (N_916,In_637,In_746);
nand U917 (N_917,In_2083,In_54);
xnor U918 (N_918,In_432,In_1169);
nor U919 (N_919,In_2482,In_578);
and U920 (N_920,In_447,In_2872);
nand U921 (N_921,In_1438,In_1425);
and U922 (N_922,In_474,In_2386);
xnor U923 (N_923,In_2320,In_52);
nor U924 (N_924,In_2915,In_445);
xnor U925 (N_925,In_1765,In_1965);
or U926 (N_926,In_343,In_2984);
and U927 (N_927,In_955,In_2823);
xor U928 (N_928,In_2480,In_121);
nor U929 (N_929,In_490,In_1390);
xnor U930 (N_930,In_1484,In_16);
nor U931 (N_931,In_443,In_2797);
nand U932 (N_932,In_2630,In_727);
xor U933 (N_933,In_1394,In_1339);
nor U934 (N_934,In_830,In_2113);
or U935 (N_935,In_979,In_1519);
or U936 (N_936,In_905,In_2895);
xor U937 (N_937,In_2647,In_715);
nor U938 (N_938,In_390,In_790);
or U939 (N_939,In_14,In_1853);
nor U940 (N_940,In_2791,In_1662);
nor U941 (N_941,In_2520,In_1057);
nor U942 (N_942,In_371,In_1981);
and U943 (N_943,In_2226,In_1160);
or U944 (N_944,In_2376,In_287);
nand U945 (N_945,In_2252,In_1071);
and U946 (N_946,In_1486,In_519);
and U947 (N_947,In_2659,In_186);
or U948 (N_948,In_2428,In_1933);
xor U949 (N_949,In_1845,In_1235);
and U950 (N_950,In_634,In_409);
and U951 (N_951,In_1415,In_895);
xor U952 (N_952,In_1521,In_352);
or U953 (N_953,In_1401,In_517);
nor U954 (N_954,In_2312,In_1926);
or U955 (N_955,In_745,In_1143);
nand U956 (N_956,In_1216,In_2810);
and U957 (N_957,In_768,In_704);
or U958 (N_958,In_1359,In_2856);
or U959 (N_959,In_605,In_1442);
nand U960 (N_960,In_1821,In_1779);
nand U961 (N_961,In_1215,In_906);
xor U962 (N_962,In_2690,In_1871);
and U963 (N_963,In_1983,In_1142);
and U964 (N_964,In_2142,In_1048);
nor U965 (N_965,In_1786,In_492);
or U966 (N_966,In_2605,In_1581);
nor U967 (N_967,In_1232,In_1767);
or U968 (N_968,In_2503,In_2224);
nor U969 (N_969,In_2131,In_232);
xnor U970 (N_970,In_1307,In_2286);
xor U971 (N_971,In_2065,In_1799);
nand U972 (N_972,In_1703,In_2307);
and U973 (N_973,In_729,In_1117);
xor U974 (N_974,In_2613,In_2154);
and U975 (N_975,In_681,In_274);
or U976 (N_976,In_2195,In_2000);
xnor U977 (N_977,In_2878,In_2522);
nor U978 (N_978,In_2897,In_221);
or U979 (N_979,In_1104,In_1370);
xnor U980 (N_980,In_2994,In_2636);
xor U981 (N_981,In_98,In_1785);
nor U982 (N_982,In_1898,In_2162);
and U983 (N_983,In_649,In_461);
and U984 (N_984,In_1399,In_2328);
nor U985 (N_985,In_2675,In_683);
xnor U986 (N_986,In_1759,In_92);
nor U987 (N_987,In_2965,In_29);
nor U988 (N_988,In_2464,In_1006);
nor U989 (N_989,In_2978,In_1719);
and U990 (N_990,In_187,In_126);
and U991 (N_991,In_85,In_2186);
nand U992 (N_992,In_476,In_1812);
and U993 (N_993,In_2588,In_1361);
or U994 (N_994,In_810,In_1960);
nor U995 (N_995,In_614,In_2406);
nand U996 (N_996,In_314,In_587);
or U997 (N_997,In_2201,In_2577);
nor U998 (N_998,In_130,In_2092);
and U999 (N_999,In_47,In_2510);
nor U1000 (N_1000,In_219,In_2998);
nor U1001 (N_1001,In_264,In_108);
or U1002 (N_1002,In_1062,In_1698);
nand U1003 (N_1003,In_2523,In_2104);
xor U1004 (N_1004,In_2953,In_781);
and U1005 (N_1005,In_34,In_5);
or U1006 (N_1006,In_342,In_893);
xor U1007 (N_1007,In_1913,In_382);
or U1008 (N_1008,In_2418,In_780);
xor U1009 (N_1009,In_1533,In_2988);
or U1010 (N_1010,In_2541,In_2814);
xor U1011 (N_1011,In_2200,In_788);
or U1012 (N_1012,In_618,In_1368);
and U1013 (N_1013,In_2615,In_1150);
nor U1014 (N_1014,In_1099,In_1572);
xor U1015 (N_1015,In_2046,In_2016);
nand U1016 (N_1016,In_2035,In_2919);
and U1017 (N_1017,In_172,In_1035);
and U1018 (N_1018,In_137,In_2961);
xnor U1019 (N_1019,In_2456,In_2704);
or U1020 (N_1020,In_65,In_2080);
xnor U1021 (N_1021,In_563,In_2044);
nor U1022 (N_1022,In_255,In_189);
or U1023 (N_1023,In_702,In_521);
xor U1024 (N_1024,In_2051,In_740);
and U1025 (N_1025,In_334,In_529);
nand U1026 (N_1026,In_2321,In_879);
xor U1027 (N_1027,In_168,In_809);
nand U1028 (N_1028,In_1320,In_2122);
and U1029 (N_1029,In_2662,In_2297);
nor U1030 (N_1030,In_40,In_2324);
or U1031 (N_1031,In_434,In_1585);
or U1032 (N_1032,In_802,In_2805);
or U1033 (N_1033,In_1855,In_1183);
and U1034 (N_1034,In_2616,In_2419);
xnor U1035 (N_1035,In_1944,In_2879);
xnor U1036 (N_1036,In_1269,In_957);
or U1037 (N_1037,In_184,In_1769);
and U1038 (N_1038,In_1727,In_138);
and U1039 (N_1039,In_19,In_1556);
nor U1040 (N_1040,In_1825,In_558);
and U1041 (N_1041,In_366,In_1375);
nand U1042 (N_1042,In_295,In_1804);
nand U1043 (N_1043,In_597,In_2177);
and U1044 (N_1044,In_2269,In_1537);
nor U1045 (N_1045,In_1775,In_2167);
xor U1046 (N_1046,In_1116,In_1923);
nor U1047 (N_1047,In_2222,In_297);
nor U1048 (N_1048,In_473,In_1754);
or U1049 (N_1049,In_2936,In_2650);
and U1050 (N_1050,In_2916,In_1446);
nor U1051 (N_1051,In_2118,In_2420);
and U1052 (N_1052,In_1250,In_2929);
nor U1053 (N_1053,In_987,In_231);
nand U1054 (N_1054,In_762,In_2660);
and U1055 (N_1055,In_84,In_2017);
xor U1056 (N_1056,In_2693,In_2185);
nor U1057 (N_1057,In_2834,In_2722);
or U1058 (N_1058,In_1582,In_1483);
nand U1059 (N_1059,In_916,In_1757);
nor U1060 (N_1060,In_2304,In_356);
and U1061 (N_1061,In_513,In_1279);
and U1062 (N_1062,In_2414,In_1137);
or U1063 (N_1063,In_644,In_1241);
or U1064 (N_1064,In_1503,In_2479);
and U1065 (N_1065,In_2077,In_1434);
nor U1066 (N_1066,In_1579,In_1587);
or U1067 (N_1067,In_2217,In_1917);
xor U1068 (N_1068,In_1559,In_1291);
nand U1069 (N_1069,In_1781,In_2141);
and U1070 (N_1070,In_566,In_728);
and U1071 (N_1071,In_682,In_2515);
and U1072 (N_1072,In_2215,In_1632);
nand U1073 (N_1073,In_1528,In_2011);
and U1074 (N_1074,In_2528,In_1121);
nor U1075 (N_1075,In_1253,In_1752);
nand U1076 (N_1076,In_2500,In_423);
nand U1077 (N_1077,In_2346,In_561);
or U1078 (N_1078,In_1731,In_2134);
nand U1079 (N_1079,In_341,In_1554);
xnor U1080 (N_1080,In_761,In_1017);
nand U1081 (N_1081,In_967,In_1412);
and U1082 (N_1082,In_500,In_2643);
xor U1083 (N_1083,In_2939,In_2921);
or U1084 (N_1084,In_206,In_489);
and U1085 (N_1085,In_2072,In_2646);
nand U1086 (N_1086,In_2999,In_1025);
and U1087 (N_1087,In_1974,In_2266);
xor U1088 (N_1088,In_2219,In_1620);
and U1089 (N_1089,In_429,In_1869);
xnor U1090 (N_1090,In_872,In_2568);
and U1091 (N_1091,In_2155,In_1424);
or U1092 (N_1092,In_2835,In_1299);
or U1093 (N_1093,In_1669,In_1467);
nand U1094 (N_1094,In_2290,In_1146);
or U1095 (N_1095,In_439,In_136);
and U1096 (N_1096,In_2446,In_102);
xnor U1097 (N_1097,In_2645,In_1936);
nand U1098 (N_1098,In_856,In_2821);
or U1099 (N_1099,In_1508,In_2569);
xor U1100 (N_1100,In_2787,In_1174);
and U1101 (N_1101,In_347,In_2624);
nand U1102 (N_1102,In_2453,In_71);
xor U1103 (N_1103,In_852,In_2840);
nand U1104 (N_1104,In_2772,In_2886);
and U1105 (N_1105,In_185,In_2294);
nor U1106 (N_1106,In_45,In_965);
nand U1107 (N_1107,In_38,In_1650);
nand U1108 (N_1108,In_1841,In_2287);
and U1109 (N_1109,In_111,In_969);
and U1110 (N_1110,In_2582,In_1649);
and U1111 (N_1111,In_2089,In_2549);
and U1112 (N_1112,In_753,In_408);
xor U1113 (N_1113,In_1249,In_2989);
or U1114 (N_1114,In_1790,In_2623);
xnor U1115 (N_1115,In_68,In_159);
and U1116 (N_1116,In_533,In_1838);
xor U1117 (N_1117,In_798,In_2191);
nand U1118 (N_1118,In_1491,In_1776);
nand U1119 (N_1119,In_931,In_1507);
xor U1120 (N_1120,In_835,In_2144);
and U1121 (N_1121,In_2173,In_2674);
or U1122 (N_1122,In_1912,In_2444);
nand U1123 (N_1123,In_266,In_1730);
and U1124 (N_1124,In_585,In_1472);
nor U1125 (N_1125,In_716,In_722);
and U1126 (N_1126,In_785,In_1034);
nand U1127 (N_1127,In_2750,In_236);
xnor U1128 (N_1128,In_956,In_1995);
and U1129 (N_1129,In_2617,In_690);
xnor U1130 (N_1130,In_2220,In_1605);
nor U1131 (N_1131,In_2486,In_760);
xnor U1132 (N_1132,In_1856,In_195);
or U1133 (N_1133,In_2497,In_1569);
nand U1134 (N_1134,In_322,In_23);
xor U1135 (N_1135,In_279,In_2327);
nor U1136 (N_1136,In_1365,In_1471);
or U1137 (N_1137,In_2038,In_738);
or U1138 (N_1138,In_152,In_1285);
or U1139 (N_1139,In_2385,In_2681);
nand U1140 (N_1140,In_2980,In_240);
xnor U1141 (N_1141,In_833,In_2378);
or U1142 (N_1142,In_1231,In_486);
nand U1143 (N_1143,In_2359,In_2218);
or U1144 (N_1144,In_1802,In_1874);
nand U1145 (N_1145,In_1897,In_993);
and U1146 (N_1146,In_874,In_2796);
or U1147 (N_1147,In_1381,In_2727);
and U1148 (N_1148,In_1565,In_2349);
or U1149 (N_1149,In_2193,In_2283);
nand U1150 (N_1150,In_2342,In_1963);
and U1151 (N_1151,In_1836,In_564);
nor U1152 (N_1152,In_299,In_795);
and U1153 (N_1153,In_552,In_1260);
nor U1154 (N_1154,In_868,In_2345);
nor U1155 (N_1155,In_697,In_2873);
xor U1156 (N_1156,In_1602,In_1780);
nand U1157 (N_1157,In_1694,In_2095);
and U1158 (N_1158,In_1106,In_1735);
or U1159 (N_1159,In_999,In_733);
or U1160 (N_1160,In_1573,In_1072);
xnor U1161 (N_1161,In_712,In_1864);
xor U1162 (N_1162,In_2527,In_838);
and U1163 (N_1163,In_884,In_671);
nand U1164 (N_1164,In_646,In_667);
nand U1165 (N_1165,In_2358,In_1027);
nor U1166 (N_1166,In_384,In_455);
nand U1167 (N_1167,In_2573,In_44);
or U1168 (N_1168,In_2731,In_2789);
and U1169 (N_1169,In_718,In_2586);
nand U1170 (N_1170,In_1945,In_263);
nor U1171 (N_1171,In_504,In_2728);
and U1172 (N_1172,In_590,In_1751);
nor U1173 (N_1173,In_2393,In_951);
nor U1174 (N_1174,In_2127,In_735);
nor U1175 (N_1175,In_330,In_56);
and U1176 (N_1176,In_2368,In_442);
nor U1177 (N_1177,In_891,In_1749);
and U1178 (N_1178,In_259,In_1959);
or U1179 (N_1179,In_2612,In_1426);
and U1180 (N_1180,In_2620,In_1455);
or U1181 (N_1181,In_404,In_2761);
nand U1182 (N_1182,In_2053,In_2803);
or U1183 (N_1183,In_2747,In_1929);
nor U1184 (N_1184,In_460,In_666);
nor U1185 (N_1185,In_803,In_368);
nor U1186 (N_1186,In_1827,In_1369);
nand U1187 (N_1187,In_1997,In_1021);
nor U1188 (N_1188,In_1012,In_912);
and U1189 (N_1189,In_1907,In_1577);
nor U1190 (N_1190,In_196,In_836);
xnor U1191 (N_1191,In_2639,In_1456);
nor U1192 (N_1192,In_145,In_939);
or U1193 (N_1193,In_1466,In_688);
or U1194 (N_1194,In_2476,In_1304);
or U1195 (N_1195,In_1580,In_1937);
nor U1196 (N_1196,In_508,In_786);
or U1197 (N_1197,In_1788,In_69);
nor U1198 (N_1198,In_2114,In_437);
nand U1199 (N_1199,In_1351,In_2745);
or U1200 (N_1200,In_2391,N_1100);
xnor U1201 (N_1201,In_858,N_268);
or U1202 (N_1202,N_32,In_527);
nand U1203 (N_1203,N_62,N_1191);
and U1204 (N_1204,N_543,N_301);
nand U1205 (N_1205,N_354,N_72);
xor U1206 (N_1206,N_259,In_2413);
nor U1207 (N_1207,N_997,N_1172);
or U1208 (N_1208,N_585,In_1713);
and U1209 (N_1209,In_2228,N_339);
xnor U1210 (N_1210,N_978,N_448);
or U1211 (N_1211,N_143,N_699);
nor U1212 (N_1212,In_1238,N_21);
nand U1213 (N_1213,N_563,In_2649);
nand U1214 (N_1214,N_815,N_390);
and U1215 (N_1215,In_209,In_1676);
and U1216 (N_1216,In_1941,N_1112);
or U1217 (N_1217,N_103,N_781);
nand U1218 (N_1218,N_411,In_1060);
nand U1219 (N_1219,N_635,N_518);
and U1220 (N_1220,N_787,In_860);
or U1221 (N_1221,In_2511,In_105);
nand U1222 (N_1222,In_2656,N_392);
xnor U1223 (N_1223,N_65,In_1706);
nand U1224 (N_1224,N_191,N_702);
or U1225 (N_1225,In_143,N_456);
nand U1226 (N_1226,In_2295,In_2698);
and U1227 (N_1227,In_2013,In_190);
xor U1228 (N_1228,In_58,N_1139);
or U1229 (N_1229,N_555,N_928);
and U1230 (N_1230,N_230,N_766);
and U1231 (N_1231,In_2954,In_2904);
and U1232 (N_1232,In_135,N_876);
and U1233 (N_1233,In_213,In_1408);
xnor U1234 (N_1234,N_93,N_1153);
nor U1235 (N_1235,N_600,N_811);
or U1236 (N_1236,In_2758,N_564);
nand U1237 (N_1237,N_1084,N_127);
or U1238 (N_1238,N_129,N_739);
nand U1239 (N_1239,In_2430,In_1055);
xor U1240 (N_1240,N_694,N_355);
nor U1241 (N_1241,In_1626,In_1755);
or U1242 (N_1242,N_803,In_355);
and U1243 (N_1243,N_653,N_688);
and U1244 (N_1244,N_490,N_409);
and U1245 (N_1245,N_3,N_288);
or U1246 (N_1246,In_1205,In_894);
nand U1247 (N_1247,N_910,N_179);
or U1248 (N_1248,In_147,N_350);
xor U1249 (N_1249,N_114,In_2653);
xnor U1250 (N_1250,In_1294,N_848);
nor U1251 (N_1251,N_971,In_2819);
or U1252 (N_1252,In_991,N_492);
and U1253 (N_1253,In_1686,N_300);
or U1254 (N_1254,N_960,N_894);
nand U1255 (N_1255,N_535,N_49);
or U1256 (N_1256,N_1098,N_1088);
nor U1257 (N_1257,In_2716,N_1134);
nor U1258 (N_1258,In_2594,N_623);
nand U1259 (N_1259,In_2802,In_2135);
nor U1260 (N_1260,In_1430,In_1345);
or U1261 (N_1261,N_839,N_202);
and U1262 (N_1262,In_1549,N_1045);
nand U1263 (N_1263,N_269,In_2576);
and U1264 (N_1264,N_712,N_472);
nor U1265 (N_1265,N_1011,N_613);
or U1266 (N_1266,In_717,N_571);
or U1267 (N_1267,N_576,N_184);
xor U1268 (N_1268,In_358,In_639);
nor U1269 (N_1269,In_985,N_1187);
or U1270 (N_1270,In_2766,N_1062);
and U1271 (N_1271,In_660,In_1315);
or U1272 (N_1272,N_598,N_888);
nor U1273 (N_1273,N_331,In_613);
nor U1274 (N_1274,N_692,In_1305);
or U1275 (N_1275,N_886,In_2179);
nand U1276 (N_1276,In_2962,N_484);
and U1277 (N_1277,N_356,In_462);
nor U1278 (N_1278,In_2208,N_588);
and U1279 (N_1279,N_667,N_324);
nor U1280 (N_1280,N_46,N_63);
nor U1281 (N_1281,N_1009,N_559);
nor U1282 (N_1282,In_1998,In_1950);
xnor U1283 (N_1283,N_295,N_728);
nand U1284 (N_1284,In_1217,N_539);
and U1285 (N_1285,In_501,N_551);
and U1286 (N_1286,N_890,In_645);
or U1287 (N_1287,In_2421,In_1086);
xnor U1288 (N_1288,In_2434,In_1568);
xor U1289 (N_1289,N_14,N_553);
nor U1290 (N_1290,N_181,N_1162);
xnor U1291 (N_1291,In_327,N_583);
xnor U1292 (N_1292,In_2362,N_109);
nand U1293 (N_1293,N_526,N_678);
xor U1294 (N_1294,In_2147,N_90);
and U1295 (N_1295,N_465,N_570);
or U1296 (N_1296,In_1546,N_774);
and U1297 (N_1297,N_206,N_167);
or U1298 (N_1298,In_1598,In_1567);
or U1299 (N_1299,In_1228,N_87);
nor U1300 (N_1300,In_79,N_603);
or U1301 (N_1301,In_976,N_340);
and U1302 (N_1302,N_926,N_681);
or U1303 (N_1303,N_1046,In_2268);
nand U1304 (N_1304,N_627,N_863);
nand U1305 (N_1305,N_517,In_238);
or U1306 (N_1306,N_901,N_1021);
nor U1307 (N_1307,N_174,N_446);
nand U1308 (N_1308,N_172,In_412);
or U1309 (N_1309,N_22,In_2212);
and U1310 (N_1310,N_56,In_2024);
or U1311 (N_1311,In_1000,N_383);
and U1312 (N_1312,In_59,N_393);
nor U1313 (N_1313,N_58,In_2400);
xnor U1314 (N_1314,N_791,In_431);
xnor U1315 (N_1315,In_572,In_1985);
or U1316 (N_1316,N_414,N_575);
xnor U1317 (N_1317,N_777,In_1544);
nor U1318 (N_1318,N_1087,In_2958);
and U1319 (N_1319,N_194,N_523);
nand U1320 (N_1320,N_1180,N_892);
xor U1321 (N_1321,In_749,In_1753);
and U1322 (N_1322,N_1176,N_469);
nor U1323 (N_1323,N_176,In_2857);
nor U1324 (N_1324,N_554,N_664);
and U1325 (N_1325,N_972,In_2654);
xnor U1326 (N_1326,N_332,N_483);
or U1327 (N_1327,In_1275,N_271);
xnor U1328 (N_1328,N_15,N_979);
nand U1329 (N_1329,In_1851,N_964);
or U1330 (N_1330,N_297,N_683);
xnor U1331 (N_1331,N_796,In_1379);
nor U1332 (N_1332,N_13,N_733);
nand U1333 (N_1333,N_887,N_691);
nand U1334 (N_1334,N_240,N_79);
xor U1335 (N_1335,N_474,N_990);
xor U1336 (N_1336,In_2337,N_146);
or U1337 (N_1337,N_77,N_333);
and U1338 (N_1338,In_1973,N_227);
nand U1339 (N_1339,N_567,N_1095);
and U1340 (N_1340,N_807,In_1489);
nor U1341 (N_1341,N_326,In_1224);
or U1342 (N_1342,In_176,N_632);
or U1343 (N_1343,N_716,N_629);
xnor U1344 (N_1344,N_258,N_151);
nor U1345 (N_1345,N_1174,In_1324);
and U1346 (N_1346,N_266,N_314);
nor U1347 (N_1347,N_207,N_342);
xor U1348 (N_1348,N_234,In_1010);
nor U1349 (N_1349,N_1074,N_372);
nor U1350 (N_1350,N_919,N_522);
and U1351 (N_1351,N_723,In_2732);
xor U1352 (N_1352,N_171,N_1189);
xnor U1353 (N_1353,N_75,In_2950);
or U1354 (N_1354,N_159,N_459);
nor U1355 (N_1355,N_64,N_854);
nand U1356 (N_1356,In_986,N_962);
or U1357 (N_1357,N_337,N_601);
nand U1358 (N_1358,N_1083,In_202);
nor U1359 (N_1359,In_1113,In_658);
nand U1360 (N_1360,In_1722,In_676);
nand U1361 (N_1361,N_1154,In_673);
or U1362 (N_1362,In_1878,In_2161);
nor U1363 (N_1363,N_514,N_581);
nor U1364 (N_1364,N_959,N_164);
and U1365 (N_1365,In_2086,In_1763);
or U1366 (N_1366,In_2640,N_1048);
and U1367 (N_1367,N_579,N_418);
nor U1368 (N_1368,In_215,In_1651);
or U1369 (N_1369,N_906,In_714);
or U1370 (N_1370,N_1033,N_647);
xnor U1371 (N_1371,N_1022,N_382);
nor U1372 (N_1372,N_663,N_403);
and U1373 (N_1373,N_91,N_873);
xnor U1374 (N_1374,N_361,N_408);
nand U1375 (N_1375,N_40,In_1056);
nand U1376 (N_1376,N_377,In_806);
and U1377 (N_1377,N_424,In_643);
and U1378 (N_1378,N_531,N_1096);
or U1379 (N_1379,In_482,N_558);
nor U1380 (N_1380,In_2512,N_609);
nor U1381 (N_1381,In_1545,In_818);
xnor U1382 (N_1382,N_1159,N_397);
or U1383 (N_1383,N_582,N_281);
nand U1384 (N_1384,N_987,N_1106);
and U1385 (N_1385,N_197,N_457);
nand U1386 (N_1386,N_55,In_2843);
xnor U1387 (N_1387,In_2552,In_1028);
or U1388 (N_1388,In_2085,In_2979);
and U1389 (N_1389,In_1209,N_1013);
nand U1390 (N_1390,In_2451,N_315);
or U1391 (N_1391,In_2673,N_78);
or U1392 (N_1392,N_123,N_20);
nor U1393 (N_1393,N_923,N_669);
xnor U1394 (N_1394,N_500,N_60);
xnor U1395 (N_1395,N_239,N_718);
and U1396 (N_1396,N_1026,N_52);
or U1397 (N_1397,N_441,In_616);
xor U1398 (N_1398,N_984,N_1185);
xor U1399 (N_1399,N_958,In_1604);
nand U1400 (N_1400,N_931,In_2898);
xnor U1401 (N_1401,In_252,N_1072);
and U1402 (N_1402,N_1165,N_318);
nor U1403 (N_1403,N_94,N_780);
nand U1404 (N_1404,N_875,In_1153);
or U1405 (N_1405,N_695,N_495);
nand U1406 (N_1406,N_1182,N_419);
or U1407 (N_1407,N_955,In_1077);
or U1408 (N_1408,N_957,N_726);
nor U1409 (N_1409,N_1117,N_652);
and U1410 (N_1410,N_161,N_360);
nand U1411 (N_1411,N_938,N_279);
or U1412 (N_1412,In_1922,N_686);
and U1413 (N_1413,In_651,In_277);
nand U1414 (N_1414,In_1693,In_239);
nand U1415 (N_1415,N_577,In_1536);
nand U1416 (N_1416,N_398,In_2783);
xor U1417 (N_1417,N_1144,N_1016);
nor U1418 (N_1418,In_582,In_1807);
nand U1419 (N_1419,N_1170,In_739);
nor U1420 (N_1420,N_918,N_454);
nor U1421 (N_1421,In_1527,N_814);
and U1422 (N_1422,N_643,N_306);
nand U1423 (N_1423,In_2387,N_250);
and U1424 (N_1424,N_144,In_2778);
or U1425 (N_1425,In_2971,N_1020);
nor U1426 (N_1426,In_1271,In_150);
or U1427 (N_1427,In_775,N_133);
xor U1428 (N_1428,N_710,N_816);
and U1429 (N_1429,N_110,N_1133);
nor U1430 (N_1430,N_199,N_1056);
or U1431 (N_1431,N_320,N_1094);
nand U1432 (N_1432,In_600,N_953);
xnor U1433 (N_1433,N_69,In_1496);
nand U1434 (N_1434,N_630,In_2940);
or U1435 (N_1435,In_397,N_602);
nand U1436 (N_1436,In_863,N_325);
or U1437 (N_1437,In_1210,N_826);
nand U1438 (N_1438,N_822,N_488);
or U1439 (N_1439,N_429,N_205);
or U1440 (N_1440,N_203,N_636);
xor U1441 (N_1441,In_2439,N_458);
or U1442 (N_1442,N_660,In_2190);
nand U1443 (N_1443,N_1086,N_335);
xor U1444 (N_1444,N_366,N_940);
or U1445 (N_1445,N_45,N_1038);
or U1446 (N_1446,N_169,N_658);
nand U1447 (N_1447,In_1494,In_2928);
or U1448 (N_1448,In_2808,N_675);
or U1449 (N_1449,N_1099,In_1801);
nor U1450 (N_1450,N_192,N_965);
nand U1451 (N_1451,N_120,N_1120);
nand U1452 (N_1452,N_437,N_925);
and U1453 (N_1453,N_274,N_608);
or U1454 (N_1454,N_348,In_60);
xor U1455 (N_1455,N_920,N_477);
xnor U1456 (N_1456,N_974,N_1060);
nand U1457 (N_1457,N_1066,In_598);
or U1458 (N_1458,N_713,In_194);
nand U1459 (N_1459,N_677,N_473);
or U1460 (N_1460,In_345,In_784);
xnor U1461 (N_1461,N_1090,N_497);
nand U1462 (N_1462,N_186,N_47);
nor U1463 (N_1463,In_1505,In_2407);
xor U1464 (N_1464,In_2484,In_2538);
and U1465 (N_1465,In_2117,N_772);
nor U1466 (N_1466,In_1360,N_1055);
and U1467 (N_1467,In_2555,In_1403);
xor U1468 (N_1468,N_177,In_349);
nor U1469 (N_1469,N_157,N_1156);
or U1470 (N_1470,N_769,N_891);
or U1471 (N_1471,N_445,N_696);
xnor U1472 (N_1472,In_932,N_349);
nor U1473 (N_1473,N_351,N_1105);
xnor U1474 (N_1474,In_292,N_435);
or U1475 (N_1475,N_1006,N_493);
nor U1476 (N_1476,In_1016,N_1044);
and U1477 (N_1477,In_2862,N_961);
xnor U1478 (N_1478,In_2815,In_2986);
and U1479 (N_1479,N_1183,N_933);
or U1480 (N_1480,N_638,In_2076);
xor U1481 (N_1481,N_294,In_1363);
xor U1482 (N_1482,In_1314,N_837);
nand U1483 (N_1483,In_2094,In_1870);
nor U1484 (N_1484,In_2262,N_307);
and U1485 (N_1485,In_1891,N_54);
and U1486 (N_1486,N_275,N_980);
nand U1487 (N_1487,In_2429,In_2143);
nor U1488 (N_1488,N_540,N_254);
or U1489 (N_1489,N_939,N_1168);
xnor U1490 (N_1490,N_927,N_670);
and U1491 (N_1491,N_420,N_1179);
and U1492 (N_1492,N_1115,N_756);
xor U1493 (N_1493,In_2635,N_977);
xnor U1494 (N_1494,N_140,In_2182);
nand U1495 (N_1495,In_1994,N_1075);
nor U1496 (N_1496,N_720,N_762);
nor U1497 (N_1497,In_2908,N_1129);
nand U1498 (N_1498,In_1921,In_2174);
nand U1499 (N_1499,N_736,N_806);
xor U1500 (N_1500,N_212,In_1931);
nand U1501 (N_1501,N_1097,N_819);
and U1502 (N_1502,N_804,N_634);
nand U1503 (N_1503,N_434,N_256);
and U1504 (N_1504,In_1091,In_1100);
nor U1505 (N_1505,N_820,N_124);
or U1506 (N_1506,N_1118,N_153);
xnor U1507 (N_1507,N_672,N_198);
nor U1508 (N_1508,N_359,N_166);
nand U1509 (N_1509,N_450,In_1817);
and U1510 (N_1510,N_840,N_412);
or U1511 (N_1511,N_1043,N_1093);
and U1512 (N_1512,N_520,N_183);
xnor U1513 (N_1513,N_1042,N_125);
nor U1514 (N_1514,In_767,In_2270);
nor U1515 (N_1515,N_797,In_2771);
and U1516 (N_1516,N_101,In_1695);
or U1517 (N_1517,N_385,N_673);
nor U1518 (N_1518,N_821,N_273);
or U1519 (N_1519,N_236,N_23);
nor U1520 (N_1520,N_462,In_2459);
and U1521 (N_1521,N_1190,In_1014);
nand U1522 (N_1522,In_1822,N_417);
and U1523 (N_1523,In_1978,N_903);
or U1524 (N_1524,In_2663,N_902);
nand U1525 (N_1525,N_433,N_651);
and U1526 (N_1526,N_1173,N_649);
and U1527 (N_1527,N_818,N_481);
and U1528 (N_1528,In_2483,N_415);
xor U1529 (N_1529,N_371,In_2571);
xnor U1530 (N_1530,In_290,N_914);
and U1531 (N_1531,N_1089,N_1135);
and U1532 (N_1532,N_1108,N_160);
nor U1533 (N_1533,N_966,N_869);
or U1534 (N_1534,N_232,In_686);
nor U1535 (N_1535,In_1600,In_1972);
nand U1536 (N_1536,In_2540,N_1037);
or U1537 (N_1537,N_389,N_499);
or U1538 (N_1538,In_528,N_995);
nand U1539 (N_1539,In_1338,N_685);
and U1540 (N_1540,N_621,N_374);
or U1541 (N_1541,In_1800,N_249);
nor U1542 (N_1542,N_264,N_530);
or U1543 (N_1543,N_352,N_1034);
nand U1544 (N_1544,N_1178,N_70);
xor U1545 (N_1545,N_864,N_771);
and U1546 (N_1546,In_100,In_1487);
or U1547 (N_1547,N_257,N_168);
xor U1548 (N_1548,In_2091,In_1265);
nor U1549 (N_1549,N_871,In_820);
and U1550 (N_1550,In_1892,In_2964);
and U1551 (N_1551,N_593,N_1155);
nor U1552 (N_1552,In_2754,N_36);
xnor U1553 (N_1553,N_568,N_730);
xor U1554 (N_1554,N_4,N_1010);
and U1555 (N_1555,N_790,N_237);
nor U1556 (N_1556,N_53,N_973);
or U1557 (N_1557,N_1110,In_88);
nor U1558 (N_1558,N_1057,In_2785);
and U1559 (N_1559,N_7,N_308);
xnor U1560 (N_1560,In_1251,N_883);
xor U1561 (N_1561,N_432,In_2415);
nand U1562 (N_1562,In_81,N_642);
nor U1563 (N_1563,N_1,N_480);
and U1564 (N_1564,N_89,In_2012);
or U1565 (N_1565,N_261,N_565);
and U1566 (N_1566,N_528,N_178);
xor U1567 (N_1567,N_1052,N_746);
nand U1568 (N_1568,N_607,N_687);
nand U1569 (N_1569,N_379,N_661);
nand U1570 (N_1570,N_1130,N_785);
nor U1571 (N_1571,N_1058,N_967);
nand U1572 (N_1572,In_1684,In_1444);
nand U1573 (N_1573,N_399,In_226);
xnor U1574 (N_1574,N_1177,N_130);
nor U1575 (N_1575,In_402,N_122);
and U1576 (N_1576,N_33,In_1683);
or U1577 (N_1577,N_421,N_700);
nor U1578 (N_1578,N_98,N_862);
xnor U1579 (N_1579,N_1123,N_721);
nor U1580 (N_1580,N_201,In_2717);
nor U1581 (N_1581,In_2280,In_2488);
nor U1582 (N_1582,N_2,In_2256);
xor U1583 (N_1583,In_2521,N_856);
nand U1584 (N_1584,N_589,In_2238);
nand U1585 (N_1585,N_1169,N_1141);
nor U1586 (N_1586,N_881,N_362);
xnor U1587 (N_1587,In_873,N_423);
nor U1588 (N_1588,N_646,N_665);
or U1589 (N_1589,N_674,N_668);
and U1590 (N_1590,N_711,In_31);
xor U1591 (N_1591,N_679,In_464);
and U1592 (N_1592,N_99,In_726);
and U1593 (N_1593,N_900,N_116);
or U1594 (N_1594,N_289,N_233);
or U1595 (N_1595,N_783,N_1003);
xor U1596 (N_1596,In_2471,In_2350);
nand U1597 (N_1597,In_1346,N_494);
nor U1598 (N_1598,In_1655,N_865);
xor U1599 (N_1599,N_624,N_1027);
or U1600 (N_1600,In_361,N_852);
xnor U1601 (N_1601,N_272,N_561);
and U1602 (N_1602,N_363,N_375);
xnor U1603 (N_1603,N_616,N_1029);
and U1604 (N_1604,N_843,In_117);
and U1605 (N_1605,In_339,In_1382);
nor U1606 (N_1606,N_948,N_440);
or U1607 (N_1607,N_989,In_253);
and U1608 (N_1608,N_968,N_615);
nor U1609 (N_1609,N_759,N_376);
and U1610 (N_1610,In_2125,N_1111);
nand U1611 (N_1611,N_1039,N_829);
xnor U1612 (N_1612,In_289,N_113);
xor U1613 (N_1613,In_2817,In_2830);
nor U1614 (N_1614,In_1833,N_929);
nor U1615 (N_1615,N_1079,N_1136);
nor U1616 (N_1616,N_1103,N_732);
or U1617 (N_1617,N_666,In_300);
nor U1618 (N_1618,N_1107,N_1121);
xnor U1619 (N_1619,N_801,N_943);
xor U1620 (N_1620,In_2,N_963);
and U1621 (N_1621,In_1905,N_365);
nor U1622 (N_1622,N_527,N_1124);
nand U1623 (N_1623,In_417,N_475);
and U1624 (N_1624,N_396,N_190);
nand U1625 (N_1625,In_1796,N_731);
nand U1626 (N_1626,In_536,N_30);
or U1627 (N_1627,N_38,N_825);
nor U1628 (N_1628,N_436,N_519);
and U1629 (N_1629,In_724,N_513);
nor U1630 (N_1630,In_315,In_1186);
and U1631 (N_1631,N_1114,N_1050);
nand U1632 (N_1632,In_1619,N_509);
and U1633 (N_1633,N_180,N_304);
nor U1634 (N_1634,N_631,N_126);
xnor U1635 (N_1635,N_283,N_976);
nand U1636 (N_1636,N_1030,N_388);
and U1637 (N_1637,In_2001,N_662);
and U1638 (N_1638,N_501,N_751);
or U1639 (N_1639,N_754,N_188);
nand U1640 (N_1640,In_2332,N_338);
nand U1641 (N_1641,In_1266,N_884);
and U1642 (N_1642,In_2847,N_66);
nor U1643 (N_1643,N_548,In_1488);
nand U1644 (N_1644,N_427,In_148);
nor U1645 (N_1645,N_846,N_132);
and U1646 (N_1646,N_932,In_923);
nor U1647 (N_1647,In_1090,In_2007);
xnor U1648 (N_1648,N_165,In_2888);
or U1649 (N_1649,N_701,N_1051);
and U1650 (N_1650,N_404,N_874);
nand U1651 (N_1651,In_1492,In_2355);
nor U1652 (N_1652,N_867,N_1049);
or U1653 (N_1653,N_1065,In_1844);
xor U1654 (N_1654,N_221,N_478);
and U1655 (N_1655,In_1791,In_584);
and U1656 (N_1656,In_1886,In_1418);
xnor U1657 (N_1657,In_76,N_1067);
xor U1658 (N_1658,In_1076,N_302);
nand U1659 (N_1659,N_1147,N_438);
nor U1660 (N_1660,N_245,In_2567);
or U1661 (N_1661,In_1164,N_1157);
xnor U1662 (N_1662,N_817,N_482);
xnor U1663 (N_1663,N_328,N_1005);
nand U1664 (N_1664,N_628,N_620);
or U1665 (N_1665,N_345,N_1140);
and U1666 (N_1666,N_1119,In_244);
nor U1667 (N_1667,N_1068,In_35);
nand U1668 (N_1668,In_2634,N_1025);
nor U1669 (N_1669,In_414,In_792);
nor U1670 (N_1670,N_861,N_850);
or U1671 (N_1671,In_2109,N_225);
xor U1672 (N_1672,In_2314,In_1388);
nand U1673 (N_1673,In_2353,N_722);
nor U1674 (N_1674,In_2828,N_135);
nor U1675 (N_1675,N_776,In_1318);
nand U1676 (N_1676,In_2799,In_2462);
xor U1677 (N_1677,N_842,N_511);
nor U1678 (N_1678,N_725,N_596);
nand U1679 (N_1679,N_341,N_34);
xor U1680 (N_1680,N_357,In_2151);
xor U1681 (N_1681,N_27,In_2301);
xor U1682 (N_1682,N_18,N_1143);
or U1683 (N_1683,N_562,N_805);
nand U1684 (N_1684,N_946,N_496);
nand U1685 (N_1685,In_2593,In_2037);
and U1686 (N_1686,In_1349,In_1707);
nand U1687 (N_1687,N_158,In_2943);
nand U1688 (N_1688,In_177,N_136);
and U1689 (N_1689,N_155,In_2172);
nor U1690 (N_1690,N_128,N_1145);
xor U1691 (N_1691,N_515,In_1461);
nand U1692 (N_1692,In_112,In_158);
and U1693 (N_1693,In_210,In_1085);
or U1694 (N_1694,In_1859,In_2335);
nand U1695 (N_1695,In_864,In_270);
xor U1696 (N_1696,N_908,In_2839);
nand U1697 (N_1697,N_213,In_2547);
nor U1698 (N_1698,N_1195,N_1019);
xor U1699 (N_1699,N_453,N_590);
or U1700 (N_1700,N_899,N_280);
xnor U1701 (N_1701,N_491,N_193);
xor U1702 (N_1702,N_449,N_868);
nor U1703 (N_1703,N_162,In_2291);
and U1704 (N_1704,N_758,N_1199);
nor U1705 (N_1705,In_1560,N_76);
nand U1706 (N_1706,N_706,N_877);
nor U1707 (N_1707,In_2235,In_516);
nor U1708 (N_1708,N_770,N_347);
xor U1709 (N_1709,In_2816,N_1102);
nand U1710 (N_1710,In_1835,N_464);
and U1711 (N_1711,In_75,N_8);
and U1712 (N_1712,N_83,In_369);
and U1713 (N_1713,N_97,N_106);
nor U1714 (N_1714,N_216,In_1372);
nor U1715 (N_1715,In_502,N_657);
nand U1716 (N_1716,N_285,N_43);
nor U1717 (N_1717,N_930,N_975);
nor U1718 (N_1718,N_611,N_296);
and U1719 (N_1719,N_541,In_2468);
nor U1720 (N_1720,N_1192,N_485);
nand U1721 (N_1721,In_164,In_950);
or U1722 (N_1722,In_2058,In_1092);
nand U1723 (N_1723,In_1621,N_671);
and U1724 (N_1724,In_119,N_578);
or U1725 (N_1725,N_11,N_1054);
xnor U1726 (N_1726,N_982,N_529);
nor U1727 (N_1727,In_2363,N_836);
nand U1728 (N_1728,N_690,N_154);
xor U1729 (N_1729,N_48,N_506);
or U1730 (N_1730,N_26,In_2248);
xor U1731 (N_1731,N_999,N_148);
nor U1732 (N_1732,N_784,In_1526);
or U1733 (N_1733,N_291,In_783);
nand U1734 (N_1734,N_1017,N_470);
xor U1735 (N_1735,N_752,In_1033);
or U1736 (N_1736,N_996,N_1161);
xnor U1737 (N_1737,In_1745,In_622);
nand U1738 (N_1738,N_747,N_619);
nand U1739 (N_1739,In_1657,N_329);
or U1740 (N_1740,In_2706,In_944);
xor U1741 (N_1741,N_945,N_265);
nor U1742 (N_1742,In_466,N_1032);
and U1743 (N_1743,In_318,In_2737);
or U1744 (N_1744,In_2043,N_391);
nand U1745 (N_1745,In_1506,N_895);
nor U1746 (N_1746,N_947,In_1257);
and U1747 (N_1747,N_163,N_533);
nor U1748 (N_1748,In_764,N_298);
nor U1749 (N_1749,N_1125,In_1671);
and U1750 (N_1750,N_556,In_278);
xnor U1751 (N_1751,In_1538,In_1378);
xnor U1752 (N_1752,N_1166,In_440);
xnor U1753 (N_1753,N_709,N_594);
xnor U1754 (N_1754,In_1952,In_1274);
nor U1755 (N_1755,In_694,In_1194);
xnor U1756 (N_1756,N_1001,N_364);
or U1757 (N_1757,N_400,N_1031);
nand U1758 (N_1758,N_952,In_340);
or U1759 (N_1759,N_170,N_743);
nand U1760 (N_1760,N_786,N_451);
nand U1761 (N_1761,N_909,N_231);
xor U1762 (N_1762,N_447,N_879);
and U1763 (N_1763,N_1171,In_399);
xnor U1764 (N_1764,N_546,In_1612);
or U1765 (N_1765,N_534,In_1685);
nor U1766 (N_1766,In_1680,N_878);
xor U1767 (N_1767,N_276,N_260);
and U1768 (N_1768,N_757,N_587);
or U1769 (N_1769,N_765,In_2273);
nand U1770 (N_1770,N_334,N_724);
nand U1771 (N_1771,N_416,N_387);
nand U1772 (N_1772,In_2970,In_2473);
nor U1773 (N_1773,N_956,N_460);
nand U1774 (N_1774,N_1002,In_2223);
nand U1775 (N_1775,In_1588,N_309);
or U1776 (N_1776,N_1035,N_800);
nor U1777 (N_1777,N_808,In_848);
nor U1778 (N_1778,N_386,N_644);
nand U1779 (N_1779,In_49,N_788);
or U1780 (N_1780,N_773,N_857);
and U1781 (N_1781,In_425,In_2499);
nand U1782 (N_1782,N_214,N_625);
nand U1783 (N_1783,N_405,N_704);
and U1784 (N_1784,N_431,N_941);
nand U1785 (N_1785,In_635,N_88);
or U1786 (N_1786,N_322,N_310);
nand U1787 (N_1787,In_1543,N_917);
or U1788 (N_1788,N_1078,N_1081);
or U1789 (N_1789,In_1958,N_1059);
or U1790 (N_1790,N_612,N_599);
nor U1791 (N_1791,N_1193,In_2275);
xor U1792 (N_1792,In_2026,In_2889);
xnor U1793 (N_1793,N_954,In_2422);
nand U1794 (N_1794,N_209,N_111);
and U1795 (N_1795,N_737,N_761);
nand U1796 (N_1796,In_2330,N_312);
xor U1797 (N_1797,In_2614,N_858);
and U1798 (N_1798,In_248,In_1875);
and U1799 (N_1799,In_2438,N_1138);
nor U1800 (N_1800,N_905,In_1353);
nor U1801 (N_1801,N_654,In_346);
xor U1802 (N_1802,In_2199,N_95);
nand U1803 (N_1803,In_904,In_2440);
and U1804 (N_1804,N_882,N_224);
or U1805 (N_1805,N_538,N_262);
xor U1806 (N_1806,N_860,N_218);
or U1807 (N_1807,N_467,N_698);
and U1808 (N_1808,In_1861,N_439);
nand U1809 (N_1809,N_911,N_915);
or U1810 (N_1810,N_617,In_1774);
xnor U1811 (N_1811,N_1018,N_604);
nor U1812 (N_1812,In_2308,N_693);
and U1813 (N_1813,In_620,N_986);
xor U1814 (N_1814,N_305,N_498);
nand U1815 (N_1815,N_1163,N_1070);
nand U1816 (N_1816,In_6,N_648);
nor U1817 (N_1817,N_131,In_2045);
and U1818 (N_1818,N_100,In_2906);
nand U1819 (N_1819,N_96,N_597);
or U1820 (N_1820,N_16,N_833);
or U1821 (N_1821,In_2216,N_220);
nand U1822 (N_1822,N_369,In_424);
nor U1823 (N_1823,N_1014,N_640);
and U1824 (N_1824,N_637,N_107);
and U1825 (N_1825,N_50,N_656);
nand U1826 (N_1826,N_645,In_1675);
and U1827 (N_1827,N_606,N_442);
and U1828 (N_1828,In_869,N_19);
and U1829 (N_1829,In_2329,N_557);
xor U1830 (N_1830,In_1469,N_219);
or U1831 (N_1831,N_738,N_247);
or U1832 (N_1832,N_1142,In_857);
and U1833 (N_1833,N_327,In_225);
or U1834 (N_1834,N_1082,N_394);
or U1835 (N_1835,N_1092,N_1085);
and U1836 (N_1836,N_150,N_80);
nand U1837 (N_1837,N_468,N_476);
nor U1838 (N_1838,In_2115,N_880);
and U1839 (N_1839,N_750,In_1393);
nand U1840 (N_1840,In_652,N_544);
and U1841 (N_1841,In_855,In_2537);
xor U1842 (N_1842,In_1725,N_838);
xnor U1843 (N_1843,N_748,N_745);
or U1844 (N_1844,N_373,N_1148);
and U1845 (N_1845,N_284,N_6);
and U1846 (N_1846,N_907,N_367);
xnor U1847 (N_1847,N_775,N_573);
or U1848 (N_1848,In_1659,N_512);
and U1849 (N_1849,N_277,N_729);
nand U1850 (N_1850,In_2039,N_552);
and U1851 (N_1851,N_73,N_487);
xnor U1852 (N_1852,In_2807,In_2458);
or U1853 (N_1853,N_727,In_1207);
nand U1854 (N_1854,N_242,N_626);
nor U1855 (N_1855,N_1061,N_536);
and U1856 (N_1856,In_2781,N_1181);
nor U1857 (N_1857,In_2788,In_36);
xnor U1858 (N_1858,In_2317,N_1008);
nor U1859 (N_1859,N_740,In_2152);
nor U1860 (N_1860,In_2607,In_2927);
xnor U1861 (N_1861,N_248,In_2809);
or U1862 (N_1862,N_137,N_985);
nor U1863 (N_1863,N_545,In_1316);
nor U1864 (N_1864,N_102,N_549);
xnor U1865 (N_1865,In_2891,N_828);
nand U1866 (N_1866,N_537,N_944);
and U1867 (N_1867,In_2469,N_1041);
xor U1868 (N_1868,N_115,In_2691);
xor U1869 (N_1869,N_35,N_370);
nor U1870 (N_1870,In_1911,In_328);
xor U1871 (N_1871,In_2912,N_278);
or U1872 (N_1872,N_1069,N_584);
or U1873 (N_1873,N_1028,N_368);
or U1874 (N_1874,N_9,N_639);
xnor U1875 (N_1875,N_1188,In_825);
nor U1876 (N_1876,In_2900,N_410);
nand U1877 (N_1877,In_542,N_1175);
xnor U1878 (N_1878,In_2709,N_145);
xor U1879 (N_1879,N_270,In_309);
nor U1880 (N_1880,N_108,N_1007);
or U1881 (N_1881,N_547,N_1158);
xor U1882 (N_1882,N_208,N_24);
or U1883 (N_1883,N_182,In_251);
xnor U1884 (N_1884,N_1132,In_2918);
xnor U1885 (N_1885,In_2288,N_204);
nand U1886 (N_1886,N_282,N_44);
and U1887 (N_1887,N_226,N_1150);
nand U1888 (N_1888,In_2563,N_897);
and U1889 (N_1889,N_793,N_443);
nand U1890 (N_1890,N_592,N_904);
nor U1891 (N_1891,In_2822,N_1076);
or U1892 (N_1892,N_574,In_2323);
or U1893 (N_1893,In_1059,In_1223);
or U1894 (N_1894,In_77,In_288);
and U1895 (N_1895,In_2111,In_747);
xor U1896 (N_1896,N_413,N_251);
xor U1897 (N_1897,In_1858,N_241);
or U1898 (N_1898,In_257,In_1462);
and U1899 (N_1899,N_719,In_2405);
nor U1900 (N_1900,N_25,In_2606);
and U1901 (N_1901,In_303,N_235);
xnor U1902 (N_1902,N_1012,N_17);
or U1903 (N_1903,N_152,N_841);
xor U1904 (N_1904,N_532,In_200);
or U1905 (N_1905,In_2648,N_228);
nor U1906 (N_1906,In_1002,N_353);
nand U1907 (N_1907,N_916,N_1196);
nor U1908 (N_1908,N_924,N_794);
xnor U1909 (N_1909,In_1900,In_619);
nor U1910 (N_1910,N_988,N_51);
nor U1911 (N_1911,N_1137,In_1044);
xor U1912 (N_1912,In_1927,N_149);
nor U1913 (N_1913,N_1071,N_1101);
nand U1914 (N_1914,N_849,In_2375);
xnor U1915 (N_1915,N_503,In_1564);
or U1916 (N_1916,N_981,N_622);
nand U1917 (N_1917,In_2493,In_2597);
or U1918 (N_1918,In_876,N_92);
xor U1919 (N_1919,In_2938,N_810);
and U1920 (N_1920,N_1164,In_1395);
xor U1921 (N_1921,N_605,In_1125);
xor U1922 (N_1922,In_1728,N_614);
or U1923 (N_1923,N_893,In_2977);
nand U1924 (N_1924,N_507,N_215);
nand U1925 (N_1925,N_1023,In_998);
and U1926 (N_1926,N_655,N_293);
nand U1927 (N_1927,In_2246,N_313);
nand U1928 (N_1928,N_1126,N_1131);
and U1929 (N_1929,N_789,N_697);
or U1930 (N_1930,N_229,N_799);
nand U1931 (N_1931,In_2932,N_141);
nor U1932 (N_1932,N_950,N_505);
nand U1933 (N_1933,N_994,In_1980);
or U1934 (N_1934,N_802,N_41);
xor U1935 (N_1935,N_767,N_336);
and U1936 (N_1936,In_2158,N_992);
xnor U1937 (N_1937,N_173,N_1184);
nor U1938 (N_1938,N_74,N_346);
or U1939 (N_1939,N_39,N_572);
and U1940 (N_1940,N_898,In_1518);
nor U1941 (N_1941,In_2723,N_211);
nor U1942 (N_1942,In_1029,In_1966);
or U1943 (N_1943,In_1457,N_489);
xnor U1944 (N_1944,N_749,In_1094);
nand U1945 (N_1945,N_401,In_193);
or U1946 (N_1946,In_2705,N_684);
xor U1947 (N_1947,N_253,N_117);
and U1948 (N_1948,N_112,In_698);
nand U1949 (N_1949,In_2740,N_1063);
xor U1950 (N_1950,N_121,In_428);
nor U1951 (N_1951,In_1221,N_983);
nor U1952 (N_1952,In_131,In_2274);
nand U1953 (N_1953,N_795,In_214);
nand U1954 (N_1954,In_396,N_1149);
xnor U1955 (N_1955,N_1109,In_1136);
nand U1956 (N_1956,N_1186,In_2744);
and U1957 (N_1957,N_1146,N_104);
xnor U1958 (N_1958,In_229,N_118);
or U1959 (N_1959,N_1000,In_1768);
nor U1960 (N_1960,In_881,N_896);
and U1961 (N_1961,N_384,In_2505);
nor U1962 (N_1962,N_455,In_1144);
xnor U1963 (N_1963,N_463,In_2631);
or U1964 (N_1964,In_935,N_1004);
and U1965 (N_1965,N_407,N_870);
nand U1966 (N_1966,N_866,N_1152);
nor U1967 (N_1967,N_61,N_969);
nand U1968 (N_1968,In_37,N_156);
xor U1969 (N_1969,N_189,N_735);
and U1970 (N_1970,In_2243,N_1116);
nor U1971 (N_1971,N_134,N_222);
and U1972 (N_1972,In_556,In_2742);
xnor U1973 (N_1973,N_851,N_566);
or U1974 (N_1974,N_10,N_844);
nand U1975 (N_1975,N_1040,In_2837);
nor U1976 (N_1976,N_428,N_591);
xor U1977 (N_1977,N_834,N_471);
nand U1978 (N_1978,In_2082,N_486);
nor U1979 (N_1979,N_1197,In_2697);
and U1980 (N_1980,In_2924,N_742);
or U1981 (N_1981,In_1850,N_659);
or U1982 (N_1982,N_452,In_494);
xor U1983 (N_1983,N_764,N_824);
or U1984 (N_1984,N_922,In_2959);
or U1985 (N_1985,In_2124,N_1047);
xor U1986 (N_1986,In_488,N_1036);
or U1987 (N_1987,N_105,N_760);
nor U1988 (N_1988,In_1714,N_610);
and U1989 (N_1989,N_406,N_316);
xnor U1990 (N_1990,N_82,N_422);
or U1991 (N_1991,N_586,N_937);
nand U1992 (N_1992,In_2844,N_524);
nand U1993 (N_1993,N_708,N_1080);
nor U1994 (N_1994,N_717,N_650);
nand U1995 (N_1995,N_217,N_936);
nand U1996 (N_1996,N_1024,N_921);
and U1997 (N_1997,N_778,N_823);
nor U1998 (N_1998,In_914,N_1194);
nand U1999 (N_1999,N_763,N_703);
or U2000 (N_2000,N_560,N_287);
nand U2001 (N_2001,In_1635,In_1292);
xnor U2002 (N_2002,N_1160,N_29);
xnor U2003 (N_2003,In_1197,N_319);
or U2004 (N_2004,N_299,N_768);
nor U2005 (N_2005,N_81,N_831);
or U2006 (N_2006,N_633,N_286);
or U2007 (N_2007,In_2554,N_267);
xnor U2008 (N_2008,N_714,N_1104);
nor U2009 (N_2009,N_138,In_1636);
nand U2010 (N_2010,In_1078,N_569);
xnor U2011 (N_2011,N_290,N_147);
or U2012 (N_2012,N_425,N_195);
nor U2013 (N_2013,In_389,In_276);
and U2014 (N_2014,N_395,N_37);
xor U2015 (N_2015,In_1336,N_1077);
nand U2016 (N_2016,N_913,N_508);
nor U2017 (N_2017,N_263,N_993);
and U2018 (N_2018,N_859,N_252);
nand U2019 (N_2019,N_28,In_885);
xnor U2020 (N_2020,N_755,N_303);
xor U2021 (N_2021,In_1276,N_246);
nand U2022 (N_2022,N_934,N_885);
nor U2023 (N_2023,N_142,In_250);
nand U2024 (N_2024,N_680,In_2204);
and U2025 (N_2025,N_991,N_461);
nor U2026 (N_2026,N_504,In_581);
or U2027 (N_2027,In_1031,N_516);
nand U2028 (N_2028,N_479,N_1113);
nand U2029 (N_2029,N_618,In_2397);
or U2030 (N_2030,N_744,N_185);
xnor U2031 (N_2031,In_977,N_1064);
or U2032 (N_2032,In_2475,N_381);
and U2033 (N_2033,In_1474,N_343);
nand U2034 (N_2034,N_187,N_935);
or U2035 (N_2035,N_855,In_57);
nand U2036 (N_2036,In_1746,N_57);
and U2037 (N_2037,N_792,N_330);
nor U2038 (N_2038,In_2417,N_42);
and U2039 (N_2039,N_317,N_809);
xnor U2040 (N_2040,In_1108,N_67);
xnor U2041 (N_2041,N_502,N_71);
xor U2042 (N_2042,N_430,In_1914);
xnor U2043 (N_2043,N_358,N_380);
nand U2044 (N_2044,N_889,N_139);
nand U2045 (N_2045,N_734,N_1091);
or U2046 (N_2046,In_1181,N_311);
nor U2047 (N_2047,N_845,In_1863);
nor U2048 (N_2048,N_676,In_2850);
nor U2049 (N_2049,N_426,N_85);
xor U2050 (N_2050,N_378,N_741);
nand U2051 (N_2051,N_12,In_1645);
and U2052 (N_2052,N_1127,N_1015);
nor U2053 (N_2053,N_86,N_550);
and U2054 (N_2054,N_238,N_1073);
and U2055 (N_2055,In_39,N_812);
and U2056 (N_2056,N_595,In_2027);
or U2057 (N_2057,In_883,In_2356);
nor U2058 (N_2058,N_1053,N_119);
nor U2059 (N_2059,N_753,N_689);
nor U2060 (N_2060,N_798,In_28);
xnor U2061 (N_2061,N_830,N_84);
xor U2062 (N_2062,N_949,In_2760);
and U2063 (N_2063,In_1167,In_1646);
or U2064 (N_2064,N_847,In_758);
and U2065 (N_2065,N_292,In_1910);
xnor U2066 (N_2066,N_402,N_31);
nand U2067 (N_2067,N_998,N_344);
and U2068 (N_2068,N_813,N_175);
nand U2069 (N_2069,N_827,N_210);
or U2070 (N_2070,N_912,N_510);
nor U2071 (N_2071,In_1371,N_0);
and U2072 (N_2072,N_323,N_682);
xor U2073 (N_2073,In_2380,In_2121);
and U2074 (N_2074,In_1459,N_5);
nor U2075 (N_2075,N_779,N_715);
nand U2076 (N_2076,N_832,In_609);
xnor U2077 (N_2077,N_59,N_223);
xnor U2078 (N_2078,N_444,N_466);
xor U2079 (N_2079,N_521,N_244);
or U2080 (N_2080,N_853,N_255);
or U2081 (N_2081,In_949,N_196);
or U2082 (N_2082,N_1122,N_782);
xnor U2083 (N_2083,N_321,N_835);
or U2084 (N_2084,In_1225,In_2967);
xor U2085 (N_2085,N_970,In_2685);
nor U2086 (N_2086,N_951,N_1167);
xnor U2087 (N_2087,N_243,In_1387);
and U2088 (N_2088,In_1140,N_542);
or U2089 (N_2089,N_1128,In_421);
nor U2090 (N_2090,N_705,In_1720);
and U2091 (N_2091,N_707,N_580);
nand U2092 (N_2092,N_641,N_1198);
or U2093 (N_2093,N_200,N_942);
and U2094 (N_2094,N_872,In_2561);
or U2095 (N_2095,N_68,In_1865);
or U2096 (N_2096,In_737,In_1087);
nor U2097 (N_2097,In_1976,N_1151);
nor U2098 (N_2098,In_1449,In_2183);
nor U2099 (N_2099,In_33,N_525);
and U2100 (N_2100,N_801,N_1151);
nand U2101 (N_2101,In_1345,N_956);
nor U2102 (N_2102,N_529,N_380);
xnor U2103 (N_2103,N_549,In_1973);
or U2104 (N_2104,In_303,In_2350);
and U2105 (N_2105,In_1316,In_1998);
xnor U2106 (N_2106,In_2521,In_739);
nor U2107 (N_2107,N_62,N_268);
nand U2108 (N_2108,N_670,N_342);
or U2109 (N_2109,In_1998,N_337);
nand U2110 (N_2110,N_256,N_500);
xor U2111 (N_2111,In_2742,N_690);
or U2112 (N_2112,N_881,N_1073);
xor U2113 (N_2113,In_2927,In_2547);
nor U2114 (N_2114,In_764,In_288);
xnor U2115 (N_2115,N_10,N_901);
and U2116 (N_2116,N_964,N_692);
or U2117 (N_2117,In_257,In_2538);
xor U2118 (N_2118,N_257,N_1076);
xor U2119 (N_2119,In_2421,N_825);
and U2120 (N_2120,N_133,N_566);
nand U2121 (N_2121,N_955,N_835);
or U2122 (N_2122,N_241,N_686);
nand U2123 (N_2123,In_2152,In_248);
and U2124 (N_2124,In_2323,In_57);
and U2125 (N_2125,In_1489,N_838);
nand U2126 (N_2126,In_673,N_477);
nor U2127 (N_2127,In_2117,In_289);
xnor U2128 (N_2128,In_2037,In_2817);
or U2129 (N_2129,N_1001,N_615);
or U2130 (N_2130,In_1878,N_363);
nand U2131 (N_2131,In_2594,N_613);
nor U2132 (N_2132,In_1657,N_837);
and U2133 (N_2133,N_48,N_159);
nor U2134 (N_2134,In_417,N_135);
xnor U2135 (N_2135,N_281,N_684);
nor U2136 (N_2136,In_2001,In_2417);
or U2137 (N_2137,In_1768,In_2499);
nand U2138 (N_2138,N_1018,N_340);
nand U2139 (N_2139,N_289,N_624);
or U2140 (N_2140,N_14,N_413);
xor U2141 (N_2141,N_535,N_1031);
xor U2142 (N_2142,N_596,N_24);
xnor U2143 (N_2143,N_1063,In_2183);
or U2144 (N_2144,In_2337,N_671);
nor U2145 (N_2145,N_1159,N_343);
or U2146 (N_2146,In_2537,In_1055);
and U2147 (N_2147,N_1147,N_455);
and U2148 (N_2148,In_425,In_2964);
and U2149 (N_2149,In_698,N_23);
xnor U2150 (N_2150,N_704,N_318);
nand U2151 (N_2151,N_1077,N_792);
xnor U2152 (N_2152,In_502,N_115);
nor U2153 (N_2153,In_1087,In_39);
xnor U2154 (N_2154,N_1033,N_360);
and U2155 (N_2155,N_42,N_1024);
nand U2156 (N_2156,N_188,In_1225);
nand U2157 (N_2157,In_425,In_2815);
nand U2158 (N_2158,In_389,N_689);
nor U2159 (N_2159,N_161,In_2246);
xor U2160 (N_2160,In_2235,N_461);
and U2161 (N_2161,N_1149,N_600);
or U2162 (N_2162,N_814,N_213);
nand U2163 (N_2163,N_391,N_403);
xor U2164 (N_2164,N_185,N_377);
nand U2165 (N_2165,In_2912,In_949);
xor U2166 (N_2166,In_2850,N_644);
xor U2167 (N_2167,N_78,N_138);
nor U2168 (N_2168,N_105,In_194);
nand U2169 (N_2169,In_1016,In_225);
and U2170 (N_2170,N_1106,N_809);
xor U2171 (N_2171,N_568,N_588);
xnor U2172 (N_2172,In_39,In_1276);
xnor U2173 (N_2173,N_654,N_933);
nand U2174 (N_2174,In_2691,N_492);
or U2175 (N_2175,N_319,N_637);
nand U2176 (N_2176,N_901,In_2656);
and U2177 (N_2177,N_508,N_1190);
nor U2178 (N_2178,In_1489,In_257);
xnor U2179 (N_2179,N_233,N_341);
and U2180 (N_2180,N_487,N_1198);
nand U2181 (N_2181,In_1459,N_170);
and U2182 (N_2182,In_2468,N_562);
and U2183 (N_2183,N_1100,N_342);
nand U2184 (N_2184,N_1151,N_250);
xor U2185 (N_2185,N_1113,N_34);
or U2186 (N_2186,N_96,In_277);
xnor U2187 (N_2187,N_1096,N_38);
nand U2188 (N_2188,In_1835,N_770);
nand U2189 (N_2189,N_261,N_1183);
or U2190 (N_2190,In_1010,N_392);
or U2191 (N_2191,N_1106,N_257);
xor U2192 (N_2192,N_1150,N_161);
nor U2193 (N_2193,In_2109,N_924);
nor U2194 (N_2194,In_349,N_166);
xor U2195 (N_2195,In_1921,In_2459);
and U2196 (N_2196,N_898,N_77);
or U2197 (N_2197,N_349,N_1062);
and U2198 (N_2198,N_937,N_379);
nand U2199 (N_2199,In_2906,N_74);
xnor U2200 (N_2200,N_900,In_1275);
or U2201 (N_2201,N_1191,In_1324);
nor U2202 (N_2202,In_1388,N_1165);
nand U2203 (N_2203,In_1353,In_1985);
nor U2204 (N_2204,N_1046,N_223);
nor U2205 (N_2205,N_567,N_753);
and U2206 (N_2206,N_659,N_870);
nor U2207 (N_2207,N_891,N_796);
xnor U2208 (N_2208,N_1070,N_91);
and U2209 (N_2209,N_251,N_65);
xnor U2210 (N_2210,N_567,In_494);
nor U2211 (N_2211,In_619,N_693);
xor U2212 (N_2212,N_1173,In_1619);
nand U2213 (N_2213,N_882,N_613);
or U2214 (N_2214,N_1199,In_2391);
nand U2215 (N_2215,N_938,N_1005);
xnor U2216 (N_2216,N_42,In_278);
xnor U2217 (N_2217,In_1635,In_2847);
nor U2218 (N_2218,In_2908,N_793);
nand U2219 (N_2219,N_1157,In_1225);
nor U2220 (N_2220,In_2977,N_666);
or U2221 (N_2221,In_369,N_365);
nand U2222 (N_2222,In_2363,N_305);
nor U2223 (N_2223,N_1187,N_543);
and U2224 (N_2224,In_1363,N_568);
and U2225 (N_2225,N_820,In_1746);
xor U2226 (N_2226,N_875,In_2135);
and U2227 (N_2227,N_1165,N_327);
or U2228 (N_2228,N_350,N_616);
nor U2229 (N_2229,N_830,In_1488);
and U2230 (N_2230,N_656,In_361);
and U2231 (N_2231,N_327,N_873);
and U2232 (N_2232,In_300,N_1106);
nor U2233 (N_2233,In_2469,N_571);
xor U2234 (N_2234,In_2434,N_571);
nand U2235 (N_2235,N_247,In_2391);
nand U2236 (N_2236,N_277,In_2977);
nand U2237 (N_2237,In_1378,In_658);
or U2238 (N_2238,N_383,In_2908);
or U2239 (N_2239,N_559,N_977);
and U2240 (N_2240,In_2808,In_464);
xnor U2241 (N_2241,N_224,In_651);
nor U2242 (N_2242,N_591,In_2027);
or U2243 (N_2243,In_2977,In_598);
nor U2244 (N_2244,N_57,N_1168);
and U2245 (N_2245,N_982,N_153);
xor U2246 (N_2246,N_515,N_338);
or U2247 (N_2247,N_455,N_626);
nand U2248 (N_2248,N_305,N_773);
nand U2249 (N_2249,In_2954,In_239);
and U2250 (N_2250,In_2332,N_19);
and U2251 (N_2251,N_397,N_966);
nand U2252 (N_2252,N_220,N_509);
nand U2253 (N_2253,N_944,N_4);
or U2254 (N_2254,N_313,N_194);
nor U2255 (N_2255,In_2228,N_711);
nor U2256 (N_2256,N_1145,N_911);
xnor U2257 (N_2257,N_668,In_2742);
nand U2258 (N_2258,N_43,N_762);
nand U2259 (N_2259,N_1003,N_874);
nand U2260 (N_2260,N_1123,N_257);
or U2261 (N_2261,In_440,In_200);
or U2262 (N_2262,N_329,In_1186);
and U2263 (N_2263,In_2499,N_910);
and U2264 (N_2264,N_201,In_784);
and U2265 (N_2265,N_84,N_661);
nand U2266 (N_2266,In_1905,N_1021);
or U2267 (N_2267,N_882,N_564);
nor U2268 (N_2268,N_313,N_58);
and U2269 (N_2269,N_554,N_1035);
and U2270 (N_2270,N_114,N_22);
or U2271 (N_2271,N_1087,In_1506);
or U2272 (N_2272,N_299,N_280);
xnor U2273 (N_2273,N_566,N_1127);
nand U2274 (N_2274,N_152,N_464);
and U2275 (N_2275,N_72,In_1100);
and U2276 (N_2276,N_906,N_49);
nand U2277 (N_2277,In_276,N_646);
and U2278 (N_2278,N_912,N_144);
xnor U2279 (N_2279,N_788,N_861);
nor U2280 (N_2280,In_1952,N_1143);
and U2281 (N_2281,In_1800,N_73);
and U2282 (N_2282,N_799,N_137);
nor U2283 (N_2283,N_524,N_94);
or U2284 (N_2284,In_767,N_1103);
nand U2285 (N_2285,N_620,In_1680);
nand U2286 (N_2286,N_569,In_462);
nor U2287 (N_2287,In_1224,N_327);
and U2288 (N_2288,N_231,N_709);
nor U2289 (N_2289,N_835,N_301);
and U2290 (N_2290,In_622,N_847);
nand U2291 (N_2291,N_293,In_214);
xnor U2292 (N_2292,In_1875,In_2723);
nand U2293 (N_2293,N_112,N_457);
nand U2294 (N_2294,In_2732,N_311);
xor U2295 (N_2295,N_305,N_1);
nand U2296 (N_2296,N_129,N_59);
and U2297 (N_2297,N_280,N_202);
nand U2298 (N_2298,In_1085,In_985);
or U2299 (N_2299,N_342,N_67);
or U2300 (N_2300,N_1193,In_2891);
nand U2301 (N_2301,In_1167,N_667);
nor U2302 (N_2302,N_221,In_2413);
nand U2303 (N_2303,In_2802,In_1294);
or U2304 (N_2304,In_1922,N_956);
nor U2305 (N_2305,N_406,In_873);
nor U2306 (N_2306,In_2744,N_658);
nand U2307 (N_2307,N_906,N_78);
xnor U2308 (N_2308,N_137,N_1133);
nor U2309 (N_2309,N_1068,In_277);
or U2310 (N_2310,In_1886,In_1745);
xor U2311 (N_2311,N_145,In_2238);
or U2312 (N_2312,N_1161,In_1318);
nor U2313 (N_2313,N_45,N_180);
nand U2314 (N_2314,In_2323,In_2649);
and U2315 (N_2315,N_122,N_769);
nand U2316 (N_2316,N_1035,N_969);
xnor U2317 (N_2317,N_438,N_532);
nand U2318 (N_2318,N_522,N_759);
nand U2319 (N_2319,In_2778,N_486);
nor U2320 (N_2320,N_1087,In_858);
and U2321 (N_2321,N_508,In_1077);
nor U2322 (N_2322,In_396,In_2158);
xnor U2323 (N_2323,N_409,N_398);
or U2324 (N_2324,N_488,N_1085);
nand U2325 (N_2325,N_629,N_875);
or U2326 (N_2326,In_1985,In_1911);
nor U2327 (N_2327,In_1087,N_1089);
xnor U2328 (N_2328,N_436,N_171);
or U2329 (N_2329,N_265,N_373);
or U2330 (N_2330,N_986,In_278);
or U2331 (N_2331,N_926,N_236);
xnor U2332 (N_2332,N_308,N_43);
xnor U2333 (N_2333,N_310,N_450);
or U2334 (N_2334,N_844,In_2649);
nor U2335 (N_2335,N_154,In_652);
xor U2336 (N_2336,N_423,In_1976);
xor U2337 (N_2337,In_1900,N_334);
nor U2338 (N_2338,N_558,N_749);
nand U2339 (N_2339,N_159,In_2888);
nor U2340 (N_2340,N_1115,In_1033);
nor U2341 (N_2341,N_761,N_931);
nor U2342 (N_2342,N_1184,N_521);
nand U2343 (N_2343,N_1073,N_738);
nor U2344 (N_2344,N_1009,In_2082);
nor U2345 (N_2345,N_123,In_1029);
xnor U2346 (N_2346,In_1536,In_2115);
nand U2347 (N_2347,N_191,In_315);
or U2348 (N_2348,N_618,N_231);
and U2349 (N_2349,N_578,N_426);
nand U2350 (N_2350,In_2124,N_699);
nand U2351 (N_2351,N_295,N_998);
nand U2352 (N_2352,N_388,N_458);
xnor U2353 (N_2353,N_945,N_949);
xnor U2354 (N_2354,N_1078,N_358);
xor U2355 (N_2355,N_904,In_1094);
nor U2356 (N_2356,N_707,N_1);
nand U2357 (N_2357,N_951,In_2026);
nor U2358 (N_2358,N_456,N_307);
or U2359 (N_2359,N_1078,In_1505);
nand U2360 (N_2360,N_29,In_2256);
or U2361 (N_2361,N_57,N_125);
or U2362 (N_2362,N_142,In_1016);
and U2363 (N_2363,N_1091,N_219);
xor U2364 (N_2364,In_1136,N_160);
and U2365 (N_2365,N_592,In_820);
or U2366 (N_2366,N_1115,N_1159);
nor U2367 (N_2367,N_263,In_414);
xnor U2368 (N_2368,N_309,In_784);
or U2369 (N_2369,N_781,N_732);
nor U2370 (N_2370,N_73,In_2950);
nand U2371 (N_2371,N_1160,N_578);
xor U2372 (N_2372,In_1604,N_141);
nand U2373 (N_2373,N_708,N_337);
or U2374 (N_2374,N_393,N_1048);
nor U2375 (N_2375,N_204,N_102);
and U2376 (N_2376,N_597,N_164);
and U2377 (N_2377,N_1148,N_1023);
nor U2378 (N_2378,In_2471,N_568);
nor U2379 (N_2379,N_576,N_1001);
xnor U2380 (N_2380,N_903,In_2043);
and U2381 (N_2381,N_37,N_17);
and U2382 (N_2382,N_1048,N_926);
xnor U2383 (N_2383,In_1560,N_320);
and U2384 (N_2384,N_157,N_916);
or U2385 (N_2385,N_56,N_894);
and U2386 (N_2386,N_570,In_2499);
nand U2387 (N_2387,In_2737,In_57);
or U2388 (N_2388,In_2172,N_1055);
nor U2389 (N_2389,In_2561,N_483);
nand U2390 (N_2390,N_138,In_1544);
nor U2391 (N_2391,N_1173,N_419);
or U2392 (N_2392,In_226,N_1052);
and U2393 (N_2393,N_451,In_210);
and U2394 (N_2394,N_343,N_279);
or U2395 (N_2395,N_629,N_295);
or U2396 (N_2396,N_419,N_424);
or U2397 (N_2397,N_407,In_1113);
nor U2398 (N_2398,N_807,In_355);
nand U2399 (N_2399,In_2451,In_1774);
or U2400 (N_2400,N_1714,N_1672);
or U2401 (N_2401,N_1543,N_1461);
and U2402 (N_2402,N_1772,N_2338);
or U2403 (N_2403,N_1715,N_1264);
xor U2404 (N_2404,N_2177,N_2081);
and U2405 (N_2405,N_1457,N_1420);
and U2406 (N_2406,N_1435,N_1650);
or U2407 (N_2407,N_1352,N_1547);
or U2408 (N_2408,N_2144,N_2072);
or U2409 (N_2409,N_1906,N_2077);
xnor U2410 (N_2410,N_1642,N_1580);
and U2411 (N_2411,N_1968,N_1503);
nand U2412 (N_2412,N_1934,N_1525);
xor U2413 (N_2413,N_1463,N_1896);
nand U2414 (N_2414,N_1568,N_1417);
or U2415 (N_2415,N_1982,N_1387);
and U2416 (N_2416,N_2108,N_1434);
or U2417 (N_2417,N_1647,N_1616);
nor U2418 (N_2418,N_1645,N_1830);
or U2419 (N_2419,N_1585,N_1865);
xor U2420 (N_2420,N_2176,N_1757);
and U2421 (N_2421,N_1952,N_1965);
nand U2422 (N_2422,N_1973,N_2193);
xor U2423 (N_2423,N_2245,N_2104);
nor U2424 (N_2424,N_2091,N_1839);
and U2425 (N_2425,N_2180,N_1700);
nor U2426 (N_2426,N_2271,N_1937);
nand U2427 (N_2427,N_1224,N_1786);
and U2428 (N_2428,N_2294,N_2254);
nor U2429 (N_2429,N_1891,N_1226);
or U2430 (N_2430,N_2341,N_1228);
nand U2431 (N_2431,N_2183,N_2034);
nor U2432 (N_2432,N_1671,N_1980);
nor U2433 (N_2433,N_2344,N_1563);
or U2434 (N_2434,N_1447,N_1635);
xor U2435 (N_2435,N_1901,N_1418);
and U2436 (N_2436,N_1837,N_1796);
nand U2437 (N_2437,N_2355,N_2178);
and U2438 (N_2438,N_1673,N_2367);
xnor U2439 (N_2439,N_1919,N_1595);
nor U2440 (N_2440,N_2377,N_2239);
nor U2441 (N_2441,N_1683,N_1974);
or U2442 (N_2442,N_1859,N_2241);
and U2443 (N_2443,N_1693,N_1208);
nor U2444 (N_2444,N_2036,N_2169);
nand U2445 (N_2445,N_1211,N_2114);
xor U2446 (N_2446,N_2362,N_1443);
or U2447 (N_2447,N_1343,N_1860);
or U2448 (N_2448,N_1766,N_1216);
or U2449 (N_2449,N_1354,N_1775);
nor U2450 (N_2450,N_2017,N_2150);
or U2451 (N_2451,N_1531,N_2010);
xor U2452 (N_2452,N_1994,N_1782);
nor U2453 (N_2453,N_1761,N_1357);
nor U2454 (N_2454,N_2262,N_1369);
and U2455 (N_2455,N_2272,N_2046);
and U2456 (N_2456,N_2020,N_1886);
xor U2457 (N_2457,N_1777,N_1899);
nand U2458 (N_2458,N_1695,N_2135);
and U2459 (N_2459,N_1458,N_1227);
and U2460 (N_2460,N_2352,N_1222);
nor U2461 (N_2461,N_1533,N_1736);
xnor U2462 (N_2462,N_1362,N_2249);
nor U2463 (N_2463,N_2201,N_1748);
nor U2464 (N_2464,N_1946,N_1963);
nand U2465 (N_2465,N_2029,N_2210);
nor U2466 (N_2466,N_2218,N_1419);
nand U2467 (N_2467,N_1338,N_1282);
xnor U2468 (N_2468,N_1425,N_1584);
and U2469 (N_2469,N_1862,N_1790);
and U2470 (N_2470,N_1769,N_1709);
nor U2471 (N_2471,N_1762,N_1827);
nor U2472 (N_2472,N_1691,N_2030);
xnor U2473 (N_2473,N_2267,N_2076);
nand U2474 (N_2474,N_1200,N_1852);
xnor U2475 (N_2475,N_1936,N_1781);
nand U2476 (N_2476,N_1276,N_2300);
or U2477 (N_2477,N_1460,N_1438);
and U2478 (N_2478,N_2000,N_1845);
and U2479 (N_2479,N_1634,N_1389);
or U2480 (N_2480,N_2316,N_1573);
xor U2481 (N_2481,N_1592,N_1971);
and U2482 (N_2482,N_1297,N_1487);
xor U2483 (N_2483,N_1491,N_2074);
and U2484 (N_2484,N_2379,N_1947);
xor U2485 (N_2485,N_1267,N_1725);
or U2486 (N_2486,N_1750,N_1524);
and U2487 (N_2487,N_1895,N_1552);
or U2488 (N_2488,N_2154,N_1307);
and U2489 (N_2489,N_1538,N_1667);
nand U2490 (N_2490,N_1441,N_1477);
xnor U2491 (N_2491,N_2045,N_1707);
and U2492 (N_2492,N_1578,N_1957);
nor U2493 (N_2493,N_2230,N_1739);
nor U2494 (N_2494,N_1253,N_1998);
and U2495 (N_2495,N_2202,N_1846);
and U2496 (N_2496,N_1215,N_2137);
nand U2497 (N_2497,N_2361,N_2158);
and U2498 (N_2498,N_1723,N_1334);
nor U2499 (N_2499,N_1662,N_2080);
nor U2500 (N_2500,N_2211,N_2263);
nand U2501 (N_2501,N_2208,N_1586);
and U2502 (N_2502,N_1666,N_1785);
and U2503 (N_2503,N_1887,N_1941);
xor U2504 (N_2504,N_1450,N_1989);
and U2505 (N_2505,N_1348,N_1238);
or U2506 (N_2506,N_2396,N_1841);
nor U2507 (N_2507,N_1356,N_1676);
and U2508 (N_2508,N_2198,N_2172);
nor U2509 (N_2509,N_2118,N_1631);
nand U2510 (N_2510,N_2206,N_1321);
and U2511 (N_2511,N_2179,N_1900);
nand U2512 (N_2512,N_2376,N_1892);
or U2513 (N_2513,N_1515,N_1923);
xnor U2514 (N_2514,N_2371,N_1655);
nand U2515 (N_2515,N_1521,N_2392);
nor U2516 (N_2516,N_1836,N_1591);
nor U2517 (N_2517,N_1445,N_2070);
xor U2518 (N_2518,N_1566,N_1350);
nand U2519 (N_2519,N_1905,N_2365);
nand U2520 (N_2520,N_1897,N_1269);
or U2521 (N_2521,N_2112,N_1867);
nor U2522 (N_2522,N_1411,N_2184);
or U2523 (N_2523,N_1404,N_1817);
nand U2524 (N_2524,N_1381,N_1997);
nor U2525 (N_2525,N_2311,N_1728);
nor U2526 (N_2526,N_1287,N_2251);
and U2527 (N_2527,N_1377,N_1665);
nor U2528 (N_2528,N_1623,N_1395);
or U2529 (N_2529,N_1880,N_1640);
and U2530 (N_2530,N_2105,N_2117);
xor U2531 (N_2531,N_1599,N_2028);
xnor U2532 (N_2532,N_1793,N_2012);
xor U2533 (N_2533,N_2189,N_1472);
nor U2534 (N_2534,N_2337,N_1606);
or U2535 (N_2535,N_2139,N_1433);
xnor U2536 (N_2536,N_2385,N_1383);
nand U2537 (N_2537,N_1696,N_2186);
nand U2538 (N_2538,N_2278,N_2102);
and U2539 (N_2539,N_1201,N_2242);
xor U2540 (N_2540,N_2357,N_1554);
and U2541 (N_2541,N_2207,N_1530);
and U2542 (N_2542,N_1265,N_1259);
and U2543 (N_2543,N_2369,N_1663);
xor U2544 (N_2544,N_1217,N_1614);
nor U2545 (N_2545,N_1581,N_2326);
and U2546 (N_2546,N_2312,N_1409);
nand U2547 (N_2547,N_2260,N_1468);
xnor U2548 (N_2548,N_1493,N_2063);
nor U2549 (N_2549,N_2225,N_1885);
and U2550 (N_2550,N_2044,N_2398);
and U2551 (N_2551,N_1382,N_1870);
nor U2552 (N_2552,N_1562,N_1660);
nand U2553 (N_2553,N_2234,N_2270);
or U2554 (N_2554,N_2097,N_2128);
nand U2555 (N_2555,N_2088,N_1558);
nor U2556 (N_2556,N_2136,N_2122);
and U2557 (N_2557,N_1909,N_1744);
xor U2558 (N_2558,N_2049,N_2228);
nand U2559 (N_2559,N_1626,N_2131);
nand U2560 (N_2560,N_1427,N_1235);
nand U2561 (N_2561,N_2191,N_1483);
or U2562 (N_2562,N_1708,N_2065);
and U2563 (N_2563,N_2366,N_2322);
xor U2564 (N_2564,N_2246,N_1355);
or U2565 (N_2565,N_1309,N_1609);
nor U2566 (N_2566,N_1551,N_1414);
or U2567 (N_2567,N_2282,N_1529);
or U2568 (N_2568,N_1312,N_2149);
nor U2569 (N_2569,N_2205,N_1453);
nand U2570 (N_2570,N_2343,N_2382);
nand U2571 (N_2571,N_2243,N_2190);
or U2572 (N_2572,N_1507,N_2353);
or U2573 (N_2573,N_2227,N_2025);
and U2574 (N_2574,N_2219,N_2006);
xor U2575 (N_2575,N_2059,N_1639);
or U2576 (N_2576,N_1432,N_1204);
or U2577 (N_2577,N_2022,N_1271);
nor U2578 (N_2578,N_1763,N_1540);
xor U2579 (N_2579,N_1467,N_1240);
nand U2580 (N_2580,N_2086,N_2297);
nor U2581 (N_2581,N_1603,N_1555);
and U2582 (N_2582,N_2129,N_1764);
xnor U2583 (N_2583,N_2364,N_2147);
nand U2584 (N_2584,N_1854,N_1485);
nor U2585 (N_2585,N_1661,N_1956);
xor U2586 (N_2586,N_1351,N_1832);
or U2587 (N_2587,N_1242,N_1788);
nor U2588 (N_2588,N_2220,N_1440);
nor U2589 (N_2589,N_1544,N_1303);
nor U2590 (N_2590,N_1986,N_1929);
or U2591 (N_2591,N_1394,N_2336);
xnor U2592 (N_2592,N_1679,N_2258);
nand U2593 (N_2593,N_1260,N_2142);
xor U2594 (N_2594,N_1430,N_1471);
or U2595 (N_2595,N_1340,N_1206);
and U2596 (N_2596,N_1392,N_1313);
nor U2597 (N_2597,N_2280,N_2141);
nor U2598 (N_2598,N_2281,N_2298);
nor U2599 (N_2599,N_1541,N_1977);
xnor U2600 (N_2600,N_1298,N_1539);
nand U2601 (N_2601,N_1278,N_1470);
and U2602 (N_2602,N_1735,N_1451);
nor U2603 (N_2603,N_1464,N_1942);
or U2604 (N_2604,N_1680,N_1806);
nor U2605 (N_2605,N_1992,N_1229);
and U2606 (N_2606,N_2162,N_1526);
nor U2607 (N_2607,N_1881,N_2052);
nand U2608 (N_2608,N_1528,N_2098);
or U2609 (N_2609,N_1294,N_2256);
nand U2610 (N_2610,N_1703,N_2055);
or U2611 (N_2611,N_1209,N_2389);
xnor U2612 (N_2612,N_1358,N_1500);
xnor U2613 (N_2613,N_1940,N_2164);
nand U2614 (N_2614,N_1508,N_1903);
and U2615 (N_2615,N_1424,N_2035);
and U2616 (N_2616,N_2330,N_1505);
or U2617 (N_2617,N_1494,N_1840);
and U2618 (N_2618,N_1615,N_1292);
or U2619 (N_2619,N_1426,N_1975);
xor U2620 (N_2620,N_1602,N_1345);
nand U2621 (N_2621,N_1911,N_1575);
or U2622 (N_2622,N_2069,N_1755);
or U2623 (N_2623,N_1306,N_1588);
or U2624 (N_2624,N_1834,N_1743);
nor U2625 (N_2625,N_1462,N_2231);
nand U2626 (N_2626,N_1318,N_2145);
xnor U2627 (N_2627,N_2004,N_2094);
or U2628 (N_2628,N_1564,N_1286);
nor U2629 (N_2629,N_2383,N_1720);
xor U2630 (N_2630,N_1368,N_1363);
nand U2631 (N_2631,N_2308,N_2229);
nor U2632 (N_2632,N_1455,N_1315);
nand U2633 (N_2633,N_2185,N_1499);
xor U2634 (N_2634,N_2333,N_1904);
and U2635 (N_2635,N_1617,N_1970);
nand U2636 (N_2636,N_1407,N_2244);
nor U2637 (N_2637,N_2323,N_2192);
or U2638 (N_2638,N_1324,N_2157);
xor U2639 (N_2639,N_1364,N_2339);
or U2640 (N_2640,N_2213,N_1810);
nor U2641 (N_2641,N_1613,N_1932);
xor U2642 (N_2642,N_1884,N_1958);
nand U2643 (N_2643,N_1285,N_1898);
nor U2644 (N_2644,N_1384,N_2286);
nand U2645 (N_2645,N_1469,N_1612);
nor U2646 (N_2646,N_1939,N_1331);
nand U2647 (N_2647,N_2127,N_2363);
nor U2648 (N_2648,N_2126,N_1439);
nand U2649 (N_2649,N_1776,N_1931);
or U2650 (N_2650,N_2130,N_1203);
or U2651 (N_2651,N_1789,N_2275);
xnor U2652 (N_2652,N_1847,N_2359);
or U2653 (N_2653,N_1593,N_2195);
nor U2654 (N_2654,N_2090,N_2288);
nor U2655 (N_2655,N_1516,N_2250);
nor U2656 (N_2656,N_2067,N_1636);
nor U2657 (N_2657,N_1628,N_2289);
nand U2658 (N_2658,N_1829,N_1648);
or U2659 (N_2659,N_2167,N_1824);
nor U2660 (N_2660,N_1681,N_1778);
and U2661 (N_2661,N_2050,N_1798);
nor U2662 (N_2662,N_1474,N_1621);
nand U2663 (N_2663,N_1589,N_1262);
and U2664 (N_2664,N_1912,N_1317);
nand U2665 (N_2665,N_2350,N_2273);
xnor U2666 (N_2666,N_1740,N_1787);
nand U2667 (N_2667,N_1657,N_2075);
xor U2668 (N_2668,N_1624,N_2007);
xnor U2669 (N_2669,N_2078,N_1237);
nor U2670 (N_2670,N_1448,N_2261);
xor U2671 (N_2671,N_1797,N_2236);
and U2672 (N_2672,N_2313,N_1514);
and U2673 (N_2673,N_1247,N_1984);
xnor U2674 (N_2674,N_2143,N_1288);
and U2675 (N_2675,N_2197,N_1746);
and U2676 (N_2676,N_1610,N_1482);
nand U2677 (N_2677,N_1938,N_1882);
xor U2678 (N_2678,N_1553,N_1257);
or U2679 (N_2679,N_1756,N_2039);
and U2680 (N_2680,N_1716,N_1379);
xor U2681 (N_2681,N_2238,N_1794);
xnor U2682 (N_2682,N_1370,N_1627);
nor U2683 (N_2683,N_1386,N_1868);
or U2684 (N_2684,N_2287,N_2093);
and U2685 (N_2685,N_2399,N_1976);
xor U2686 (N_2686,N_1652,N_1391);
xnor U2687 (N_2687,N_1773,N_1619);
nor U2688 (N_2688,N_1361,N_1783);
xor U2689 (N_2689,N_2394,N_1598);
nand U2690 (N_2690,N_1339,N_1653);
nand U2691 (N_2691,N_1221,N_1630);
xnor U2692 (N_2692,N_1502,N_2106);
nand U2693 (N_2693,N_1861,N_1871);
or U2694 (N_2694,N_1659,N_1643);
xor U2695 (N_2695,N_2222,N_1388);
and U2696 (N_2696,N_1918,N_2155);
xnor U2697 (N_2697,N_1536,N_1519);
and U2698 (N_2698,N_1765,N_1376);
xor U2699 (N_2699,N_2269,N_2368);
nand U2700 (N_2700,N_1944,N_1921);
nor U2701 (N_2701,N_1953,N_1452);
or U2702 (N_2702,N_1251,N_1727);
and U2703 (N_2703,N_2019,N_1858);
nor U2704 (N_2704,N_1724,N_1632);
nand U2705 (N_2705,N_1421,N_2274);
xnor U2706 (N_2706,N_2209,N_2056);
and U2707 (N_2707,N_1360,N_2014);
xnor U2708 (N_2708,N_2259,N_1478);
nor U2709 (N_2709,N_2332,N_1574);
nor U2710 (N_2710,N_2194,N_2087);
nand U2711 (N_2711,N_1995,N_1629);
xor U2712 (N_2712,N_1234,N_1583);
xnor U2713 (N_2713,N_1688,N_1760);
or U2714 (N_2714,N_1248,N_1279);
nand U2715 (N_2715,N_2174,N_1349);
or U2716 (N_2716,N_1875,N_2027);
and U2717 (N_2717,N_1926,N_2221);
and U2718 (N_2718,N_2224,N_2391);
nor U2719 (N_2719,N_2100,N_2299);
or U2720 (N_2720,N_1985,N_2134);
and U2721 (N_2721,N_2378,N_2089);
or U2722 (N_2722,N_1393,N_1816);
or U2723 (N_2723,N_1878,N_1560);
xor U2724 (N_2724,N_1908,N_2257);
xnor U2725 (N_2725,N_2223,N_1527);
or U2726 (N_2726,N_1523,N_1272);
nand U2727 (N_2727,N_1608,N_2043);
nand U2728 (N_2728,N_1729,N_2248);
and U2729 (N_2729,N_2133,N_1687);
or U2730 (N_2730,N_2292,N_1704);
nand U2731 (N_2731,N_1570,N_2226);
nand U2732 (N_2732,N_2021,N_1556);
or U2733 (N_2733,N_1396,N_1686);
and U2734 (N_2734,N_2016,N_1826);
and U2735 (N_2735,N_1668,N_1205);
nor U2736 (N_2736,N_2170,N_1813);
xor U2737 (N_2737,N_1930,N_1694);
nor U2738 (N_2738,N_2388,N_1987);
or U2739 (N_2739,N_2001,N_1273);
nand U2740 (N_2740,N_2342,N_2232);
xor U2741 (N_2741,N_1752,N_2051);
xor U2742 (N_2742,N_1751,N_2215);
or U2743 (N_2743,N_1734,N_2315);
or U2744 (N_2744,N_1481,N_1498);
nor U2745 (N_2745,N_1654,N_1576);
and U2746 (N_2746,N_1954,N_1917);
or U2747 (N_2747,N_1999,N_1844);
nor U2748 (N_2748,N_1803,N_1620);
or U2749 (N_2749,N_2032,N_1341);
nor U2750 (N_2750,N_1405,N_1415);
nor U2751 (N_2751,N_1480,N_1275);
nor U2752 (N_2752,N_2011,N_2096);
nand U2753 (N_2753,N_1722,N_1945);
xnor U2754 (N_2754,N_1506,N_1328);
or U2755 (N_2755,N_1822,N_1293);
nand U2756 (N_2756,N_1274,N_1733);
nand U2757 (N_2757,N_2182,N_1981);
nand U2758 (N_2758,N_2372,N_1828);
or U2759 (N_2759,N_1401,N_1767);
and U2760 (N_2760,N_1833,N_1486);
or U2761 (N_2761,N_2373,N_1838);
xor U2762 (N_2762,N_2058,N_1423);
nor U2763 (N_2763,N_1296,N_1289);
xnor U2764 (N_2764,N_2053,N_1325);
xnor U2765 (N_2765,N_1326,N_2121);
nor U2766 (N_2766,N_1484,N_1712);
nor U2767 (N_2767,N_1779,N_2293);
nand U2768 (N_2768,N_2203,N_1800);
or U2769 (N_2769,N_2387,N_1266);
nor U2770 (N_2770,N_1284,N_1823);
xnor U2771 (N_2771,N_1504,N_1398);
nand U2772 (N_2772,N_1295,N_1561);
xnor U2773 (N_2773,N_2370,N_2163);
nand U2774 (N_2774,N_1913,N_1644);
xnor U2775 (N_2775,N_2319,N_1802);
or U2776 (N_2776,N_2009,N_1928);
or U2777 (N_2777,N_1791,N_1475);
or U2778 (N_2778,N_1879,N_1815);
and U2779 (N_2779,N_1412,N_2068);
nand U2780 (N_2780,N_1705,N_1651);
or U2781 (N_2781,N_1428,N_1511);
or U2782 (N_2782,N_1397,N_1873);
nand U2783 (N_2783,N_2132,N_2165);
nor U2784 (N_2784,N_2037,N_2125);
nand U2785 (N_2785,N_1509,N_1459);
xor U2786 (N_2786,N_1549,N_2384);
or U2787 (N_2787,N_1322,N_1537);
nor U2788 (N_2788,N_1565,N_1812);
nor U2789 (N_2789,N_1571,N_2015);
or U2790 (N_2790,N_2374,N_1820);
and U2791 (N_2791,N_2151,N_2252);
nand U2792 (N_2792,N_1329,N_1730);
xnor U2793 (N_2793,N_1856,N_1801);
and U2794 (N_2794,N_1342,N_1545);
nand U2795 (N_2795,N_1255,N_1607);
or U2796 (N_2796,N_1416,N_2265);
nor U2797 (N_2797,N_1915,N_1559);
or U2798 (N_2798,N_1542,N_2013);
nand U2799 (N_2799,N_2095,N_2345);
and U2800 (N_2800,N_1969,N_2103);
and U2801 (N_2801,N_2255,N_1747);
nor U2802 (N_2802,N_1737,N_2119);
nor U2803 (N_2803,N_2302,N_1855);
or U2804 (N_2804,N_1336,N_2307);
nand U2805 (N_2805,N_1966,N_1770);
or U2806 (N_2806,N_1641,N_2283);
and U2807 (N_2807,N_1814,N_1674);
xnor U2808 (N_2808,N_1239,N_1596);
and U2809 (N_2809,N_1577,N_1916);
nor U2810 (N_2810,N_1490,N_2216);
xnor U2811 (N_2811,N_1380,N_2092);
or U2812 (N_2812,N_1925,N_1857);
nor U2813 (N_2813,N_1301,N_1572);
and U2814 (N_2814,N_1811,N_2187);
nor U2815 (N_2815,N_2101,N_1476);
xnor U2816 (N_2816,N_1220,N_1214);
xnor U2817 (N_2817,N_2356,N_1308);
nor U2818 (N_2818,N_2109,N_1567);
xor U2819 (N_2819,N_1496,N_1311);
nor U2820 (N_2820,N_1246,N_2181);
nor U2821 (N_2821,N_2306,N_1821);
xor U2822 (N_2822,N_1310,N_1371);
or U2823 (N_2823,N_1479,N_2296);
and U2824 (N_2824,N_1207,N_1698);
nand U2825 (N_2825,N_2214,N_2024);
nor U2826 (N_2826,N_1869,N_1988);
or U2827 (N_2827,N_1893,N_1579);
nand U2828 (N_2828,N_2393,N_1256);
and U2829 (N_2829,N_1850,N_2047);
nand U2830 (N_2830,N_1675,N_1232);
and U2831 (N_2831,N_1225,N_2124);
xor U2832 (N_2832,N_1670,N_2291);
nor U2833 (N_2833,N_1697,N_1978);
xnor U2834 (N_2834,N_1442,N_2386);
and U2835 (N_2835,N_2290,N_1601);
or U2836 (N_2836,N_1717,N_2375);
and U2837 (N_2837,N_2107,N_1236);
and U2838 (N_2838,N_2110,N_1245);
nand U2839 (N_2839,N_1263,N_2018);
xor U2840 (N_2840,N_2380,N_1637);
xnor U2841 (N_2841,N_1961,N_2175);
nand U2842 (N_2842,N_1202,N_1706);
and U2843 (N_2843,N_1692,N_2217);
nand U2844 (N_2844,N_1210,N_2354);
nand U2845 (N_2845,N_1557,N_2146);
or U2846 (N_2846,N_2123,N_1244);
xor U2847 (N_2847,N_1831,N_1283);
and U2848 (N_2848,N_1784,N_1753);
and U2849 (N_2849,N_1951,N_1849);
nor U2850 (N_2850,N_2054,N_1853);
xor U2851 (N_2851,N_1804,N_1243);
xor U2852 (N_2852,N_2060,N_2140);
and U2853 (N_2853,N_1254,N_1335);
nand U2854 (N_2854,N_1437,N_2204);
xnor U2855 (N_2855,N_1365,N_2279);
or U2856 (N_2856,N_2309,N_1792);
xor U2857 (N_2857,N_1732,N_1894);
xor U2858 (N_2858,N_1656,N_2304);
and U2859 (N_2859,N_2240,N_1550);
nand U2860 (N_2860,N_1213,N_1872);
xnor U2861 (N_2861,N_2188,N_1385);
nor U2862 (N_2862,N_1241,N_1972);
xnor U2863 (N_2863,N_2268,N_1611);
xor U2864 (N_2864,N_2066,N_1548);
nand U2865 (N_2865,N_1372,N_1413);
xor U2866 (N_2866,N_1600,N_1863);
nor U2867 (N_2867,N_1330,N_2284);
nand U2868 (N_2868,N_2253,N_1633);
nor U2869 (N_2869,N_1252,N_1488);
nor U2870 (N_2870,N_1902,N_1344);
nand U2871 (N_2871,N_2233,N_1809);
xor U2872 (N_2872,N_1406,N_2321);
xnor U2873 (N_2873,N_1299,N_1366);
or U2874 (N_2874,N_1738,N_1532);
and U2875 (N_2875,N_1390,N_1219);
or U2876 (N_2876,N_1333,N_1277);
and U2877 (N_2877,N_1690,N_2026);
and U2878 (N_2878,N_2073,N_1497);
or U2879 (N_2879,N_2325,N_1399);
nand U2880 (N_2880,N_1646,N_2264);
or U2881 (N_2881,N_2348,N_1701);
xnor U2882 (N_2882,N_2161,N_1268);
xnor U2883 (N_2883,N_2048,N_1304);
nand U2884 (N_2884,N_1501,N_1684);
nand U2885 (N_2885,N_2237,N_1771);
nand U2886 (N_2886,N_1281,N_1864);
nand U2887 (N_2887,N_2318,N_2395);
nand U2888 (N_2888,N_1669,N_2212);
and U2889 (N_2889,N_2346,N_2160);
nand U2890 (N_2890,N_2116,N_1745);
xor U2891 (N_2891,N_2038,N_1582);
and U2892 (N_2892,N_1517,N_1924);
and U2893 (N_2893,N_2040,N_1819);
xor U2894 (N_2894,N_1535,N_2320);
nor U2895 (N_2895,N_1590,N_1492);
and U2896 (N_2896,N_2235,N_1774);
nand U2897 (N_2897,N_1922,N_2071);
and U2898 (N_2898,N_2276,N_2023);
nor U2899 (N_2899,N_1795,N_1302);
and U2900 (N_2900,N_2062,N_1983);
and U2901 (N_2901,N_1754,N_1604);
or U2902 (N_2902,N_2247,N_1713);
nor U2903 (N_2903,N_2099,N_1638);
nand U2904 (N_2904,N_2340,N_2061);
or U2905 (N_2905,N_2196,N_2310);
and U2906 (N_2906,N_1710,N_1374);
nor U2907 (N_2907,N_2285,N_1726);
xor U2908 (N_2908,N_1231,N_1520);
and U2909 (N_2909,N_1682,N_2138);
and U2910 (N_2910,N_1948,N_1373);
or U2911 (N_2911,N_1258,N_1473);
or U2912 (N_2912,N_1848,N_1883);
or U2913 (N_2913,N_1910,N_1949);
nand U2914 (N_2914,N_1979,N_2349);
nor U2915 (N_2915,N_1843,N_2057);
and U2916 (N_2916,N_1907,N_1403);
nor U2917 (N_2917,N_2152,N_2082);
xor U2918 (N_2918,N_2334,N_1955);
xor U2919 (N_2919,N_1649,N_1605);
and U2920 (N_2920,N_2328,N_1920);
xnor U2921 (N_2921,N_1678,N_1962);
and U2922 (N_2922,N_2358,N_1518);
or U2923 (N_2923,N_1465,N_1410);
nand U2924 (N_2924,N_1943,N_2153);
nor U2925 (N_2925,N_2329,N_1664);
nand U2926 (N_2926,N_2173,N_1359);
nand U2927 (N_2927,N_1959,N_1622);
and U2928 (N_2928,N_1749,N_1316);
and U2929 (N_2929,N_1594,N_1291);
and U2930 (N_2930,N_2111,N_1250);
nor U2931 (N_2931,N_1993,N_2199);
or U2932 (N_2932,N_1489,N_2159);
xnor U2933 (N_2933,N_1935,N_2327);
and U2934 (N_2934,N_2360,N_1337);
or U2935 (N_2935,N_1569,N_1877);
and U2936 (N_2936,N_1718,N_1314);
nor U2937 (N_2937,N_1933,N_1991);
nor U2938 (N_2938,N_2083,N_1444);
nand U2939 (N_2939,N_1320,N_1449);
or U2940 (N_2940,N_1768,N_2148);
xor U2941 (N_2941,N_1851,N_1587);
nor U2942 (N_2942,N_2390,N_1346);
or U2943 (N_2943,N_1914,N_1597);
nor U2944 (N_2944,N_1731,N_1466);
xor U2945 (N_2945,N_2041,N_2079);
or U2946 (N_2946,N_2002,N_1780);
xor U2947 (N_2947,N_2031,N_1719);
nand U2948 (N_2948,N_1742,N_2171);
nand U2949 (N_2949,N_2115,N_1495);
nor U2950 (N_2950,N_1431,N_1512);
nor U2951 (N_2951,N_1741,N_1721);
nor U2952 (N_2952,N_2397,N_1402);
xor U2953 (N_2953,N_1805,N_1967);
or U2954 (N_2954,N_2277,N_1689);
or U2955 (N_2955,N_2033,N_2005);
or U2956 (N_2956,N_2295,N_2156);
and U2957 (N_2957,N_1964,N_1699);
or U2958 (N_2958,N_2113,N_1842);
or U2959 (N_2959,N_1327,N_1927);
xor U2960 (N_2960,N_1261,N_1876);
nor U2961 (N_2961,N_2317,N_2381);
nor U2962 (N_2962,N_1874,N_1888);
nor U2963 (N_2963,N_2166,N_2351);
nand U2964 (N_2964,N_1400,N_2064);
nand U2965 (N_2965,N_1218,N_1454);
nand U2966 (N_2966,N_1618,N_1702);
and U2967 (N_2967,N_1323,N_2324);
and U2968 (N_2968,N_1825,N_2347);
nand U2969 (N_2969,N_1990,N_2266);
or U2970 (N_2970,N_1429,N_1290);
or U2971 (N_2971,N_2200,N_2314);
nand U2972 (N_2972,N_1446,N_1249);
or U2973 (N_2973,N_1818,N_1332);
or U2974 (N_2974,N_1799,N_1300);
and U2975 (N_2975,N_2301,N_1677);
and U2976 (N_2976,N_1758,N_1889);
nand U2977 (N_2977,N_1212,N_1378);
and U2978 (N_2978,N_1950,N_1456);
and U2979 (N_2979,N_1513,N_2168);
nor U2980 (N_2980,N_1436,N_1367);
xnor U2981 (N_2981,N_1711,N_1534);
and U2982 (N_2982,N_2042,N_1422);
and U2983 (N_2983,N_1510,N_1658);
xor U2984 (N_2984,N_2331,N_1625);
nand U2985 (N_2985,N_1546,N_1347);
xor U2986 (N_2986,N_2305,N_1685);
nor U2987 (N_2987,N_1319,N_2085);
nor U2988 (N_2988,N_1408,N_1280);
or U2989 (N_2989,N_2003,N_1866);
nand U2990 (N_2990,N_1835,N_1759);
and U2991 (N_2991,N_1223,N_2335);
and U2992 (N_2992,N_1375,N_2008);
nor U2993 (N_2993,N_1305,N_1230);
or U2994 (N_2994,N_1890,N_1270);
nand U2995 (N_2995,N_1522,N_1353);
and U2996 (N_2996,N_1807,N_2303);
or U2997 (N_2997,N_2120,N_1233);
or U2998 (N_2998,N_1960,N_1996);
nand U2999 (N_2999,N_2084,N_1808);
or U3000 (N_3000,N_1465,N_1406);
or U3001 (N_3001,N_1776,N_1388);
xor U3002 (N_3002,N_2113,N_2261);
nand U3003 (N_3003,N_1977,N_1454);
nand U3004 (N_3004,N_2208,N_1280);
nand U3005 (N_3005,N_1758,N_1250);
xnor U3006 (N_3006,N_1994,N_1661);
xnor U3007 (N_3007,N_1400,N_2130);
nor U3008 (N_3008,N_1486,N_2363);
nand U3009 (N_3009,N_1271,N_1407);
nand U3010 (N_3010,N_1423,N_1784);
and U3011 (N_3011,N_1650,N_1734);
and U3012 (N_3012,N_2075,N_1727);
or U3013 (N_3013,N_1386,N_2327);
nor U3014 (N_3014,N_1659,N_1750);
nand U3015 (N_3015,N_2123,N_1422);
xnor U3016 (N_3016,N_1446,N_2316);
and U3017 (N_3017,N_2319,N_1673);
xnor U3018 (N_3018,N_1337,N_1809);
nor U3019 (N_3019,N_1225,N_1632);
and U3020 (N_3020,N_1244,N_1767);
xor U3021 (N_3021,N_2115,N_2355);
xor U3022 (N_3022,N_1308,N_1779);
or U3023 (N_3023,N_1327,N_1664);
nor U3024 (N_3024,N_1977,N_1457);
nand U3025 (N_3025,N_1475,N_1692);
or U3026 (N_3026,N_2356,N_1475);
and U3027 (N_3027,N_2031,N_2103);
or U3028 (N_3028,N_2296,N_2081);
and U3029 (N_3029,N_1809,N_1660);
nor U3030 (N_3030,N_2187,N_1320);
xor U3031 (N_3031,N_2322,N_1966);
xor U3032 (N_3032,N_1584,N_1393);
xor U3033 (N_3033,N_1947,N_1810);
xor U3034 (N_3034,N_1729,N_1785);
or U3035 (N_3035,N_1875,N_2272);
or U3036 (N_3036,N_2334,N_1259);
nor U3037 (N_3037,N_1301,N_1507);
or U3038 (N_3038,N_1502,N_2203);
nand U3039 (N_3039,N_1345,N_2049);
or U3040 (N_3040,N_1809,N_2333);
nand U3041 (N_3041,N_1314,N_1464);
xnor U3042 (N_3042,N_1987,N_1489);
nor U3043 (N_3043,N_1303,N_1317);
and U3044 (N_3044,N_1642,N_2276);
nor U3045 (N_3045,N_1850,N_1777);
or U3046 (N_3046,N_1472,N_1547);
nand U3047 (N_3047,N_1807,N_2384);
nand U3048 (N_3048,N_1830,N_1258);
nor U3049 (N_3049,N_2025,N_1769);
or U3050 (N_3050,N_1445,N_1661);
and U3051 (N_3051,N_2025,N_2271);
nor U3052 (N_3052,N_1562,N_1428);
xor U3053 (N_3053,N_2188,N_1361);
xnor U3054 (N_3054,N_2047,N_1820);
nand U3055 (N_3055,N_1322,N_1902);
and U3056 (N_3056,N_2221,N_1807);
nand U3057 (N_3057,N_1490,N_1593);
nand U3058 (N_3058,N_2207,N_1792);
and U3059 (N_3059,N_1251,N_2078);
nand U3060 (N_3060,N_1696,N_2101);
or U3061 (N_3061,N_1659,N_1512);
xor U3062 (N_3062,N_1305,N_1384);
or U3063 (N_3063,N_2338,N_1391);
and U3064 (N_3064,N_1263,N_2305);
and U3065 (N_3065,N_1698,N_1979);
nand U3066 (N_3066,N_1377,N_1643);
nand U3067 (N_3067,N_1590,N_1785);
and U3068 (N_3068,N_1740,N_1440);
nor U3069 (N_3069,N_2298,N_1726);
nor U3070 (N_3070,N_1683,N_1344);
and U3071 (N_3071,N_1605,N_2035);
xor U3072 (N_3072,N_1506,N_1319);
nor U3073 (N_3073,N_2326,N_1589);
xnor U3074 (N_3074,N_1438,N_1944);
xnor U3075 (N_3075,N_2383,N_1665);
or U3076 (N_3076,N_2029,N_2333);
and U3077 (N_3077,N_2099,N_1401);
nor U3078 (N_3078,N_2235,N_1981);
nand U3079 (N_3079,N_2093,N_1414);
and U3080 (N_3080,N_2161,N_1462);
and U3081 (N_3081,N_1737,N_1615);
nand U3082 (N_3082,N_1286,N_1561);
nand U3083 (N_3083,N_2005,N_1808);
and U3084 (N_3084,N_2177,N_1253);
nor U3085 (N_3085,N_2055,N_1839);
xnor U3086 (N_3086,N_1299,N_2076);
or U3087 (N_3087,N_2096,N_2345);
and U3088 (N_3088,N_1541,N_2322);
and U3089 (N_3089,N_1965,N_2145);
or U3090 (N_3090,N_1927,N_2141);
nand U3091 (N_3091,N_2160,N_1239);
or U3092 (N_3092,N_1803,N_1288);
nor U3093 (N_3093,N_1631,N_1382);
and U3094 (N_3094,N_2092,N_1559);
xor U3095 (N_3095,N_1416,N_2053);
xor U3096 (N_3096,N_1416,N_2233);
nor U3097 (N_3097,N_2124,N_1661);
and U3098 (N_3098,N_1867,N_2031);
or U3099 (N_3099,N_1848,N_1631);
and U3100 (N_3100,N_1867,N_1419);
xnor U3101 (N_3101,N_2026,N_1682);
nand U3102 (N_3102,N_2307,N_1214);
xor U3103 (N_3103,N_2015,N_1980);
or U3104 (N_3104,N_1539,N_2278);
and U3105 (N_3105,N_1257,N_2087);
and U3106 (N_3106,N_1962,N_2213);
nor U3107 (N_3107,N_1212,N_1955);
nand U3108 (N_3108,N_1932,N_2079);
or U3109 (N_3109,N_1355,N_1473);
nor U3110 (N_3110,N_1972,N_2155);
or U3111 (N_3111,N_1390,N_1689);
xor U3112 (N_3112,N_1441,N_1718);
xnor U3113 (N_3113,N_2161,N_1247);
nand U3114 (N_3114,N_2314,N_1517);
nand U3115 (N_3115,N_1304,N_2239);
nand U3116 (N_3116,N_2394,N_1498);
nand U3117 (N_3117,N_2164,N_2375);
nor U3118 (N_3118,N_1302,N_2280);
or U3119 (N_3119,N_1781,N_1818);
nand U3120 (N_3120,N_1461,N_2050);
and U3121 (N_3121,N_1646,N_1308);
and U3122 (N_3122,N_2273,N_1262);
nand U3123 (N_3123,N_1530,N_2015);
nor U3124 (N_3124,N_2103,N_1915);
and U3125 (N_3125,N_2289,N_1215);
xnor U3126 (N_3126,N_1979,N_1829);
or U3127 (N_3127,N_1715,N_1971);
nor U3128 (N_3128,N_1900,N_2357);
nor U3129 (N_3129,N_2129,N_2278);
or U3130 (N_3130,N_2250,N_1699);
xnor U3131 (N_3131,N_2255,N_1508);
xor U3132 (N_3132,N_1894,N_1914);
nor U3133 (N_3133,N_1487,N_1776);
and U3134 (N_3134,N_2027,N_1977);
and U3135 (N_3135,N_2067,N_1944);
nand U3136 (N_3136,N_1422,N_2010);
xor U3137 (N_3137,N_1724,N_1524);
nor U3138 (N_3138,N_1398,N_1618);
xor U3139 (N_3139,N_1260,N_1862);
xor U3140 (N_3140,N_1715,N_1388);
and U3141 (N_3141,N_1702,N_1310);
or U3142 (N_3142,N_1734,N_2226);
or U3143 (N_3143,N_2037,N_1786);
nor U3144 (N_3144,N_1675,N_1835);
xor U3145 (N_3145,N_2288,N_2141);
nand U3146 (N_3146,N_2168,N_1601);
and U3147 (N_3147,N_1827,N_2289);
nor U3148 (N_3148,N_1607,N_1793);
or U3149 (N_3149,N_1619,N_1256);
or U3150 (N_3150,N_1639,N_1430);
or U3151 (N_3151,N_1323,N_1832);
nand U3152 (N_3152,N_1668,N_1923);
nor U3153 (N_3153,N_2050,N_2058);
nand U3154 (N_3154,N_2379,N_1231);
and U3155 (N_3155,N_2122,N_1567);
nor U3156 (N_3156,N_1595,N_2067);
and U3157 (N_3157,N_1501,N_1384);
or U3158 (N_3158,N_1685,N_1255);
and U3159 (N_3159,N_1481,N_1637);
and U3160 (N_3160,N_1804,N_1689);
xnor U3161 (N_3161,N_1667,N_1438);
xnor U3162 (N_3162,N_1875,N_1363);
nand U3163 (N_3163,N_2234,N_2118);
or U3164 (N_3164,N_1223,N_1346);
nand U3165 (N_3165,N_2051,N_1924);
nor U3166 (N_3166,N_2079,N_2266);
nor U3167 (N_3167,N_1713,N_1894);
or U3168 (N_3168,N_2029,N_1508);
and U3169 (N_3169,N_1361,N_1566);
or U3170 (N_3170,N_1698,N_2161);
and U3171 (N_3171,N_1372,N_1272);
nor U3172 (N_3172,N_1615,N_2125);
nand U3173 (N_3173,N_1677,N_1671);
nand U3174 (N_3174,N_2363,N_1650);
and U3175 (N_3175,N_2200,N_2177);
and U3176 (N_3176,N_1672,N_1938);
or U3177 (N_3177,N_1893,N_1772);
nor U3178 (N_3178,N_1971,N_1217);
or U3179 (N_3179,N_2162,N_2307);
or U3180 (N_3180,N_1301,N_2012);
nand U3181 (N_3181,N_2011,N_1320);
nor U3182 (N_3182,N_2054,N_2105);
or U3183 (N_3183,N_1856,N_1958);
nor U3184 (N_3184,N_2236,N_1288);
nand U3185 (N_3185,N_1601,N_1957);
nand U3186 (N_3186,N_1807,N_1976);
nand U3187 (N_3187,N_2273,N_2302);
or U3188 (N_3188,N_1737,N_1273);
and U3189 (N_3189,N_2217,N_1355);
nor U3190 (N_3190,N_2286,N_1372);
nor U3191 (N_3191,N_1933,N_1870);
and U3192 (N_3192,N_1660,N_1520);
nand U3193 (N_3193,N_2363,N_1253);
xor U3194 (N_3194,N_1214,N_1784);
and U3195 (N_3195,N_1892,N_1556);
and U3196 (N_3196,N_1313,N_2114);
or U3197 (N_3197,N_2314,N_1275);
nor U3198 (N_3198,N_1748,N_2122);
or U3199 (N_3199,N_2113,N_2343);
nor U3200 (N_3200,N_2176,N_1961);
nand U3201 (N_3201,N_2086,N_2310);
or U3202 (N_3202,N_2110,N_2024);
xor U3203 (N_3203,N_2175,N_1605);
nor U3204 (N_3204,N_2346,N_1743);
and U3205 (N_3205,N_1692,N_1608);
or U3206 (N_3206,N_1297,N_1426);
and U3207 (N_3207,N_1995,N_1316);
nor U3208 (N_3208,N_1653,N_2178);
and U3209 (N_3209,N_2327,N_1929);
xnor U3210 (N_3210,N_2115,N_1561);
nor U3211 (N_3211,N_2333,N_2013);
xor U3212 (N_3212,N_2082,N_1623);
or U3213 (N_3213,N_2316,N_2376);
nand U3214 (N_3214,N_2170,N_1888);
nor U3215 (N_3215,N_1727,N_1877);
nor U3216 (N_3216,N_1702,N_2009);
xor U3217 (N_3217,N_1741,N_2386);
nand U3218 (N_3218,N_2238,N_1916);
and U3219 (N_3219,N_2238,N_1351);
xor U3220 (N_3220,N_1388,N_1851);
and U3221 (N_3221,N_2364,N_1228);
and U3222 (N_3222,N_1433,N_1657);
xor U3223 (N_3223,N_1714,N_1370);
nor U3224 (N_3224,N_1619,N_2009);
nor U3225 (N_3225,N_1588,N_1930);
and U3226 (N_3226,N_1274,N_1389);
nor U3227 (N_3227,N_1286,N_2325);
nor U3228 (N_3228,N_1659,N_1640);
xnor U3229 (N_3229,N_2256,N_1605);
nor U3230 (N_3230,N_1493,N_1715);
and U3231 (N_3231,N_1635,N_2098);
and U3232 (N_3232,N_1324,N_1634);
xnor U3233 (N_3233,N_1588,N_2164);
or U3234 (N_3234,N_1252,N_2204);
xor U3235 (N_3235,N_1383,N_2260);
and U3236 (N_3236,N_2142,N_2006);
or U3237 (N_3237,N_1799,N_2308);
or U3238 (N_3238,N_1664,N_1425);
nand U3239 (N_3239,N_1975,N_1296);
or U3240 (N_3240,N_2240,N_1989);
xor U3241 (N_3241,N_2161,N_2062);
or U3242 (N_3242,N_2378,N_1267);
and U3243 (N_3243,N_2213,N_1269);
or U3244 (N_3244,N_1477,N_1579);
nor U3245 (N_3245,N_1433,N_1310);
nand U3246 (N_3246,N_1472,N_1910);
and U3247 (N_3247,N_2322,N_1638);
or U3248 (N_3248,N_2231,N_1875);
nand U3249 (N_3249,N_1490,N_1220);
and U3250 (N_3250,N_1883,N_1725);
nor U3251 (N_3251,N_2090,N_1949);
nand U3252 (N_3252,N_1372,N_1769);
nand U3253 (N_3253,N_2313,N_1636);
and U3254 (N_3254,N_1363,N_2344);
nand U3255 (N_3255,N_1475,N_1956);
and U3256 (N_3256,N_2060,N_2309);
or U3257 (N_3257,N_1232,N_1890);
nor U3258 (N_3258,N_1244,N_2210);
xor U3259 (N_3259,N_1695,N_2128);
and U3260 (N_3260,N_1226,N_2080);
xor U3261 (N_3261,N_1605,N_1394);
nand U3262 (N_3262,N_1523,N_1927);
nand U3263 (N_3263,N_2308,N_1498);
nor U3264 (N_3264,N_1580,N_1538);
xnor U3265 (N_3265,N_1614,N_2152);
nor U3266 (N_3266,N_2189,N_1971);
nand U3267 (N_3267,N_1518,N_1394);
xnor U3268 (N_3268,N_1239,N_1662);
xnor U3269 (N_3269,N_2265,N_2337);
nand U3270 (N_3270,N_1999,N_1534);
nand U3271 (N_3271,N_2386,N_2299);
xor U3272 (N_3272,N_2263,N_1442);
nand U3273 (N_3273,N_1670,N_2347);
and U3274 (N_3274,N_1499,N_1887);
or U3275 (N_3275,N_1752,N_1662);
xnor U3276 (N_3276,N_1998,N_2271);
nand U3277 (N_3277,N_2198,N_1624);
nor U3278 (N_3278,N_1544,N_2094);
nand U3279 (N_3279,N_1665,N_2063);
nand U3280 (N_3280,N_2313,N_1895);
xor U3281 (N_3281,N_2384,N_2309);
or U3282 (N_3282,N_1560,N_2170);
and U3283 (N_3283,N_2203,N_2393);
xor U3284 (N_3284,N_1749,N_2242);
or U3285 (N_3285,N_2074,N_1397);
nor U3286 (N_3286,N_1359,N_1243);
xnor U3287 (N_3287,N_1851,N_1278);
or U3288 (N_3288,N_1224,N_1748);
nand U3289 (N_3289,N_1644,N_2328);
or U3290 (N_3290,N_1591,N_1952);
nand U3291 (N_3291,N_2047,N_1428);
nor U3292 (N_3292,N_2163,N_2051);
nand U3293 (N_3293,N_1313,N_2389);
nand U3294 (N_3294,N_1773,N_1636);
nand U3295 (N_3295,N_2015,N_1921);
and U3296 (N_3296,N_2153,N_1964);
or U3297 (N_3297,N_2153,N_1985);
xnor U3298 (N_3298,N_2223,N_1643);
nor U3299 (N_3299,N_1479,N_1718);
nand U3300 (N_3300,N_1970,N_2301);
or U3301 (N_3301,N_1255,N_1387);
or U3302 (N_3302,N_1688,N_2327);
xnor U3303 (N_3303,N_2046,N_1434);
nand U3304 (N_3304,N_1681,N_1216);
xnor U3305 (N_3305,N_1571,N_2055);
nor U3306 (N_3306,N_1546,N_2194);
or U3307 (N_3307,N_2321,N_1283);
nor U3308 (N_3308,N_2265,N_1790);
nor U3309 (N_3309,N_1287,N_2069);
and U3310 (N_3310,N_1410,N_1984);
xor U3311 (N_3311,N_1586,N_1977);
and U3312 (N_3312,N_2135,N_1560);
and U3313 (N_3313,N_1264,N_1433);
and U3314 (N_3314,N_1983,N_1388);
xor U3315 (N_3315,N_2144,N_2201);
and U3316 (N_3316,N_1760,N_2149);
or U3317 (N_3317,N_2168,N_2211);
and U3318 (N_3318,N_1648,N_2314);
nand U3319 (N_3319,N_1780,N_2200);
and U3320 (N_3320,N_2088,N_1308);
nor U3321 (N_3321,N_2039,N_1533);
xor U3322 (N_3322,N_1464,N_1543);
and U3323 (N_3323,N_2065,N_1948);
or U3324 (N_3324,N_1645,N_2033);
xnor U3325 (N_3325,N_2086,N_1993);
nor U3326 (N_3326,N_2217,N_2355);
or U3327 (N_3327,N_2125,N_2139);
xor U3328 (N_3328,N_1332,N_2090);
xor U3329 (N_3329,N_1744,N_2006);
nor U3330 (N_3330,N_1292,N_1309);
and U3331 (N_3331,N_2288,N_1661);
or U3332 (N_3332,N_1737,N_2105);
nor U3333 (N_3333,N_1707,N_1267);
or U3334 (N_3334,N_2123,N_1342);
or U3335 (N_3335,N_1832,N_2024);
nor U3336 (N_3336,N_1659,N_1333);
or U3337 (N_3337,N_2377,N_2396);
and U3338 (N_3338,N_2215,N_2336);
nor U3339 (N_3339,N_2094,N_1677);
and U3340 (N_3340,N_1552,N_1911);
and U3341 (N_3341,N_1679,N_1766);
or U3342 (N_3342,N_2120,N_1236);
xor U3343 (N_3343,N_2098,N_1963);
nor U3344 (N_3344,N_2303,N_2370);
xor U3345 (N_3345,N_1952,N_1595);
xor U3346 (N_3346,N_1393,N_1631);
or U3347 (N_3347,N_2308,N_2288);
xor U3348 (N_3348,N_2033,N_2103);
nand U3349 (N_3349,N_2214,N_1403);
and U3350 (N_3350,N_1690,N_1696);
nor U3351 (N_3351,N_2399,N_1231);
and U3352 (N_3352,N_2034,N_2255);
and U3353 (N_3353,N_1624,N_1524);
and U3354 (N_3354,N_2340,N_2375);
nand U3355 (N_3355,N_1432,N_2075);
nor U3356 (N_3356,N_1690,N_2254);
or U3357 (N_3357,N_1625,N_1321);
nor U3358 (N_3358,N_1291,N_2092);
xor U3359 (N_3359,N_2071,N_1935);
nand U3360 (N_3360,N_2019,N_2264);
and U3361 (N_3361,N_2346,N_1324);
nor U3362 (N_3362,N_1695,N_1347);
nand U3363 (N_3363,N_1256,N_1668);
or U3364 (N_3364,N_1254,N_1377);
or U3365 (N_3365,N_2276,N_1333);
nand U3366 (N_3366,N_1764,N_1526);
and U3367 (N_3367,N_2216,N_2242);
or U3368 (N_3368,N_1202,N_2115);
nor U3369 (N_3369,N_1903,N_1482);
nor U3370 (N_3370,N_1611,N_1573);
and U3371 (N_3371,N_2047,N_1426);
xnor U3372 (N_3372,N_1555,N_2399);
nand U3373 (N_3373,N_2063,N_1221);
or U3374 (N_3374,N_1999,N_1701);
or U3375 (N_3375,N_2356,N_1931);
nand U3376 (N_3376,N_1602,N_1498);
nor U3377 (N_3377,N_1496,N_2267);
xnor U3378 (N_3378,N_1925,N_1482);
nor U3379 (N_3379,N_1206,N_2368);
nand U3380 (N_3380,N_2143,N_1296);
or U3381 (N_3381,N_1381,N_2315);
and U3382 (N_3382,N_2302,N_2321);
or U3383 (N_3383,N_1517,N_2186);
nor U3384 (N_3384,N_1218,N_1854);
xor U3385 (N_3385,N_1200,N_2187);
xor U3386 (N_3386,N_1744,N_1610);
xor U3387 (N_3387,N_2153,N_1722);
or U3388 (N_3388,N_2383,N_1932);
or U3389 (N_3389,N_2071,N_2067);
and U3390 (N_3390,N_1725,N_2180);
nand U3391 (N_3391,N_2287,N_2077);
and U3392 (N_3392,N_2361,N_2076);
and U3393 (N_3393,N_1656,N_1734);
and U3394 (N_3394,N_2074,N_2280);
xor U3395 (N_3395,N_1464,N_1267);
nor U3396 (N_3396,N_1870,N_1629);
and U3397 (N_3397,N_1699,N_1375);
xor U3398 (N_3398,N_2388,N_2382);
xor U3399 (N_3399,N_2322,N_1771);
or U3400 (N_3400,N_1909,N_2265);
and U3401 (N_3401,N_2014,N_1281);
nand U3402 (N_3402,N_2313,N_1560);
nand U3403 (N_3403,N_1213,N_2033);
or U3404 (N_3404,N_2198,N_1529);
nand U3405 (N_3405,N_1948,N_1218);
xor U3406 (N_3406,N_2073,N_1276);
nor U3407 (N_3407,N_1802,N_1874);
nor U3408 (N_3408,N_1490,N_1252);
nor U3409 (N_3409,N_2207,N_1303);
nand U3410 (N_3410,N_2306,N_2395);
nor U3411 (N_3411,N_1246,N_1504);
xor U3412 (N_3412,N_1731,N_1630);
nor U3413 (N_3413,N_1889,N_2291);
xor U3414 (N_3414,N_1241,N_1208);
nor U3415 (N_3415,N_1420,N_1951);
nor U3416 (N_3416,N_1889,N_1454);
or U3417 (N_3417,N_2144,N_2310);
or U3418 (N_3418,N_1844,N_1413);
nand U3419 (N_3419,N_2021,N_1440);
or U3420 (N_3420,N_1705,N_1895);
xnor U3421 (N_3421,N_1417,N_1652);
nor U3422 (N_3422,N_2125,N_2070);
and U3423 (N_3423,N_1358,N_1961);
xor U3424 (N_3424,N_1487,N_1989);
or U3425 (N_3425,N_1729,N_1633);
nand U3426 (N_3426,N_1225,N_1784);
and U3427 (N_3427,N_1703,N_2136);
nand U3428 (N_3428,N_2346,N_1471);
nand U3429 (N_3429,N_2068,N_1752);
nand U3430 (N_3430,N_2354,N_1614);
or U3431 (N_3431,N_1346,N_2041);
xor U3432 (N_3432,N_1636,N_1574);
xnor U3433 (N_3433,N_1374,N_1260);
nand U3434 (N_3434,N_2094,N_1673);
nor U3435 (N_3435,N_1729,N_1678);
and U3436 (N_3436,N_1225,N_1744);
xor U3437 (N_3437,N_1703,N_1228);
and U3438 (N_3438,N_1709,N_1738);
nor U3439 (N_3439,N_1494,N_2012);
and U3440 (N_3440,N_1238,N_1399);
nand U3441 (N_3441,N_1275,N_2198);
xor U3442 (N_3442,N_1879,N_2361);
xor U3443 (N_3443,N_2357,N_2265);
nor U3444 (N_3444,N_1690,N_1577);
nor U3445 (N_3445,N_1380,N_2373);
and U3446 (N_3446,N_1578,N_1261);
or U3447 (N_3447,N_1585,N_1409);
or U3448 (N_3448,N_1671,N_1740);
xor U3449 (N_3449,N_1593,N_1635);
xnor U3450 (N_3450,N_2339,N_1974);
nand U3451 (N_3451,N_1757,N_2289);
and U3452 (N_3452,N_1938,N_1418);
or U3453 (N_3453,N_1292,N_1459);
xnor U3454 (N_3454,N_2291,N_1702);
nand U3455 (N_3455,N_1606,N_1210);
nor U3456 (N_3456,N_1247,N_1676);
xor U3457 (N_3457,N_1407,N_1272);
xnor U3458 (N_3458,N_2142,N_1946);
or U3459 (N_3459,N_2042,N_1747);
xnor U3460 (N_3460,N_1799,N_1436);
or U3461 (N_3461,N_1589,N_1259);
nor U3462 (N_3462,N_1335,N_2155);
or U3463 (N_3463,N_1507,N_1659);
nor U3464 (N_3464,N_1973,N_1645);
nor U3465 (N_3465,N_2297,N_1335);
xor U3466 (N_3466,N_1820,N_1288);
nor U3467 (N_3467,N_1678,N_1438);
nor U3468 (N_3468,N_1868,N_1846);
and U3469 (N_3469,N_2346,N_2099);
nand U3470 (N_3470,N_1211,N_2204);
nand U3471 (N_3471,N_1880,N_1851);
xnor U3472 (N_3472,N_2109,N_1303);
or U3473 (N_3473,N_2371,N_2397);
and U3474 (N_3474,N_1281,N_1608);
nand U3475 (N_3475,N_1665,N_2035);
xor U3476 (N_3476,N_1343,N_2254);
or U3477 (N_3477,N_1415,N_2114);
or U3478 (N_3478,N_1984,N_1355);
or U3479 (N_3479,N_1446,N_2364);
nor U3480 (N_3480,N_1249,N_1295);
nand U3481 (N_3481,N_1797,N_1431);
and U3482 (N_3482,N_2355,N_1576);
nor U3483 (N_3483,N_1252,N_1682);
and U3484 (N_3484,N_1300,N_2041);
xnor U3485 (N_3485,N_1832,N_1513);
and U3486 (N_3486,N_2024,N_1795);
nand U3487 (N_3487,N_1637,N_1693);
nor U3488 (N_3488,N_1506,N_1956);
nand U3489 (N_3489,N_1743,N_1241);
or U3490 (N_3490,N_2310,N_2246);
and U3491 (N_3491,N_1587,N_1224);
or U3492 (N_3492,N_2396,N_1393);
nor U3493 (N_3493,N_2386,N_2036);
and U3494 (N_3494,N_1427,N_2064);
or U3495 (N_3495,N_1868,N_1766);
or U3496 (N_3496,N_1913,N_2047);
or U3497 (N_3497,N_1842,N_1536);
nand U3498 (N_3498,N_2280,N_2321);
xnor U3499 (N_3499,N_1457,N_1883);
and U3500 (N_3500,N_1280,N_1438);
or U3501 (N_3501,N_1652,N_1480);
and U3502 (N_3502,N_1503,N_1502);
and U3503 (N_3503,N_1484,N_1303);
nand U3504 (N_3504,N_1633,N_2335);
or U3505 (N_3505,N_2229,N_1247);
or U3506 (N_3506,N_2324,N_1732);
xnor U3507 (N_3507,N_1693,N_2018);
or U3508 (N_3508,N_1383,N_2149);
and U3509 (N_3509,N_1723,N_2098);
nand U3510 (N_3510,N_2161,N_2116);
or U3511 (N_3511,N_2116,N_2393);
or U3512 (N_3512,N_2300,N_1877);
and U3513 (N_3513,N_1833,N_1261);
nand U3514 (N_3514,N_1411,N_2088);
xnor U3515 (N_3515,N_1834,N_1914);
and U3516 (N_3516,N_1639,N_2162);
nand U3517 (N_3517,N_2126,N_1320);
xnor U3518 (N_3518,N_1543,N_1203);
nor U3519 (N_3519,N_2164,N_1582);
xnor U3520 (N_3520,N_1478,N_1354);
xnor U3521 (N_3521,N_1414,N_1663);
or U3522 (N_3522,N_1365,N_1208);
and U3523 (N_3523,N_1416,N_2225);
xnor U3524 (N_3524,N_2236,N_1996);
nor U3525 (N_3525,N_1512,N_1471);
xor U3526 (N_3526,N_1876,N_2202);
or U3527 (N_3527,N_1436,N_2043);
or U3528 (N_3528,N_1885,N_1964);
nor U3529 (N_3529,N_1314,N_1201);
and U3530 (N_3530,N_2274,N_2224);
and U3531 (N_3531,N_1285,N_1934);
xnor U3532 (N_3532,N_2232,N_1310);
nand U3533 (N_3533,N_1906,N_1247);
or U3534 (N_3534,N_1396,N_1299);
nand U3535 (N_3535,N_1209,N_1366);
or U3536 (N_3536,N_2278,N_1356);
nor U3537 (N_3537,N_1203,N_1846);
or U3538 (N_3538,N_2036,N_1813);
and U3539 (N_3539,N_1644,N_1780);
or U3540 (N_3540,N_1575,N_1758);
xnor U3541 (N_3541,N_1818,N_1899);
nor U3542 (N_3542,N_1522,N_1282);
or U3543 (N_3543,N_1582,N_1836);
or U3544 (N_3544,N_1950,N_1522);
and U3545 (N_3545,N_2131,N_1737);
nor U3546 (N_3546,N_1696,N_1323);
nand U3547 (N_3547,N_1968,N_1539);
nor U3548 (N_3548,N_1367,N_1828);
or U3549 (N_3549,N_1570,N_1579);
nand U3550 (N_3550,N_1506,N_2370);
nand U3551 (N_3551,N_1582,N_1546);
xnor U3552 (N_3552,N_2230,N_1579);
and U3553 (N_3553,N_1396,N_2217);
xor U3554 (N_3554,N_1507,N_2154);
nand U3555 (N_3555,N_2370,N_1530);
or U3556 (N_3556,N_1653,N_1512);
nand U3557 (N_3557,N_2368,N_1761);
nand U3558 (N_3558,N_2036,N_1638);
or U3559 (N_3559,N_1969,N_1231);
nor U3560 (N_3560,N_2340,N_1847);
xnor U3561 (N_3561,N_1765,N_1371);
nor U3562 (N_3562,N_1552,N_1441);
or U3563 (N_3563,N_2204,N_1430);
or U3564 (N_3564,N_1574,N_1552);
nor U3565 (N_3565,N_1775,N_1962);
nor U3566 (N_3566,N_2289,N_2234);
and U3567 (N_3567,N_2055,N_1353);
xnor U3568 (N_3568,N_1348,N_1706);
xnor U3569 (N_3569,N_1253,N_1918);
or U3570 (N_3570,N_1877,N_2108);
nor U3571 (N_3571,N_2226,N_1319);
and U3572 (N_3572,N_1894,N_2052);
xnor U3573 (N_3573,N_1819,N_1226);
nor U3574 (N_3574,N_2350,N_1662);
and U3575 (N_3575,N_2146,N_1746);
or U3576 (N_3576,N_2226,N_2285);
or U3577 (N_3577,N_1732,N_2221);
xor U3578 (N_3578,N_2194,N_2141);
and U3579 (N_3579,N_1283,N_2043);
or U3580 (N_3580,N_1994,N_1312);
and U3581 (N_3581,N_1227,N_1614);
nand U3582 (N_3582,N_1610,N_2102);
xnor U3583 (N_3583,N_1609,N_1836);
nand U3584 (N_3584,N_1803,N_1227);
xor U3585 (N_3585,N_1500,N_1258);
nand U3586 (N_3586,N_1664,N_1378);
and U3587 (N_3587,N_1683,N_1266);
and U3588 (N_3588,N_2358,N_1834);
nand U3589 (N_3589,N_2353,N_2069);
xnor U3590 (N_3590,N_1320,N_1671);
nand U3591 (N_3591,N_2274,N_1474);
nand U3592 (N_3592,N_2128,N_2135);
or U3593 (N_3593,N_2027,N_2121);
xnor U3594 (N_3594,N_2310,N_1336);
or U3595 (N_3595,N_2120,N_1435);
or U3596 (N_3596,N_1642,N_2189);
and U3597 (N_3597,N_2080,N_2208);
nand U3598 (N_3598,N_2253,N_2139);
nand U3599 (N_3599,N_1272,N_1325);
and U3600 (N_3600,N_3109,N_3160);
nand U3601 (N_3601,N_2508,N_2941);
nor U3602 (N_3602,N_3499,N_2713);
or U3603 (N_3603,N_3113,N_3529);
and U3604 (N_3604,N_2815,N_3398);
or U3605 (N_3605,N_3395,N_3356);
and U3606 (N_3606,N_2425,N_3584);
nand U3607 (N_3607,N_3348,N_2765);
nand U3608 (N_3608,N_3086,N_3040);
xor U3609 (N_3609,N_3097,N_2449);
xnor U3610 (N_3610,N_3433,N_2457);
and U3611 (N_3611,N_2939,N_3256);
nor U3612 (N_3612,N_3462,N_2679);
and U3613 (N_3613,N_3202,N_2977);
nand U3614 (N_3614,N_2572,N_3077);
xnor U3615 (N_3615,N_3385,N_2946);
xor U3616 (N_3616,N_3224,N_3142);
xnor U3617 (N_3617,N_2924,N_3330);
or U3618 (N_3618,N_2988,N_3134);
xor U3619 (N_3619,N_3360,N_3203);
or U3620 (N_3620,N_3414,N_2829);
nor U3621 (N_3621,N_2538,N_2813);
nor U3622 (N_3622,N_2549,N_3285);
and U3623 (N_3623,N_3260,N_2424);
nor U3624 (N_3624,N_2524,N_3429);
nand U3625 (N_3625,N_2413,N_3280);
nor U3626 (N_3626,N_2608,N_2741);
nand U3627 (N_3627,N_2727,N_2915);
nor U3628 (N_3628,N_3310,N_3112);
xor U3629 (N_3629,N_2701,N_2827);
and U3630 (N_3630,N_2806,N_2786);
nor U3631 (N_3631,N_2913,N_2753);
nand U3632 (N_3632,N_3015,N_3172);
or U3633 (N_3633,N_3495,N_3471);
nor U3634 (N_3634,N_3527,N_3507);
and U3635 (N_3635,N_3235,N_2527);
nor U3636 (N_3636,N_3177,N_3592);
nor U3637 (N_3637,N_3323,N_2867);
xor U3638 (N_3638,N_2529,N_3315);
nand U3639 (N_3639,N_2636,N_3291);
and U3640 (N_3640,N_2522,N_3476);
or U3641 (N_3641,N_2699,N_3418);
or U3642 (N_3642,N_2430,N_2991);
nor U3643 (N_3643,N_2757,N_2691);
nand U3644 (N_3644,N_2626,N_3312);
xnor U3645 (N_3645,N_3426,N_2485);
xnor U3646 (N_3646,N_2803,N_3123);
or U3647 (N_3647,N_2534,N_2483);
xor U3648 (N_3648,N_2982,N_2631);
nand U3649 (N_3649,N_3251,N_2942);
and U3650 (N_3650,N_3490,N_2853);
nand U3651 (N_3651,N_3294,N_3333);
xnor U3652 (N_3652,N_2825,N_2561);
xor U3653 (N_3653,N_3214,N_3493);
nor U3654 (N_3654,N_2515,N_3195);
xor U3655 (N_3655,N_3267,N_2726);
nor U3656 (N_3656,N_3271,N_3481);
xnor U3657 (N_3657,N_3517,N_3149);
nand U3658 (N_3658,N_3552,N_2749);
and U3659 (N_3659,N_3536,N_2956);
nand U3660 (N_3660,N_3340,N_3037);
and U3661 (N_3661,N_2676,N_3187);
nor U3662 (N_3662,N_2970,N_3232);
xnor U3663 (N_3663,N_2783,N_2670);
nor U3664 (N_3664,N_3266,N_2730);
xor U3665 (N_3665,N_2432,N_2934);
or U3666 (N_3666,N_2586,N_3531);
and U3667 (N_3667,N_3023,N_3598);
or U3668 (N_3668,N_3108,N_2710);
and U3669 (N_3669,N_3181,N_3401);
or U3670 (N_3670,N_3443,N_3081);
and U3671 (N_3671,N_2408,N_3168);
or U3672 (N_3672,N_3128,N_3198);
and U3673 (N_3673,N_2580,N_2844);
or U3674 (N_3674,N_2778,N_3072);
and U3675 (N_3675,N_2505,N_2474);
nor U3676 (N_3676,N_3163,N_3487);
and U3677 (N_3677,N_2969,N_2482);
or U3678 (N_3678,N_3156,N_3287);
or U3679 (N_3679,N_2661,N_2568);
or U3680 (N_3680,N_3464,N_3259);
nor U3681 (N_3681,N_3332,N_2569);
or U3682 (N_3682,N_2948,N_3103);
nor U3683 (N_3683,N_2651,N_2625);
and U3684 (N_3684,N_3222,N_2677);
or U3685 (N_3685,N_3295,N_3009);
nand U3686 (N_3686,N_3573,N_2921);
or U3687 (N_3687,N_3211,N_2732);
xor U3688 (N_3688,N_3049,N_3125);
nor U3689 (N_3689,N_3245,N_3590);
xnor U3690 (N_3690,N_3229,N_3197);
xor U3691 (N_3691,N_3297,N_2884);
nor U3692 (N_3692,N_2704,N_3524);
nor U3693 (N_3693,N_3199,N_3051);
nor U3694 (N_3694,N_3533,N_3270);
xnor U3695 (N_3695,N_3269,N_2781);
nor U3696 (N_3696,N_2849,N_3078);
xnor U3697 (N_3697,N_2464,N_3130);
or U3698 (N_3698,N_2875,N_3405);
nor U3699 (N_3699,N_3550,N_3132);
nor U3700 (N_3700,N_3062,N_3007);
nand U3701 (N_3701,N_2775,N_2647);
or U3702 (N_3702,N_3553,N_2675);
and U3703 (N_3703,N_2512,N_3101);
nand U3704 (N_3704,N_3389,N_3338);
or U3705 (N_3705,N_3148,N_3070);
xnor U3706 (N_3706,N_2936,N_2405);
and U3707 (N_3707,N_3560,N_3377);
nand U3708 (N_3708,N_2695,N_3154);
nor U3709 (N_3709,N_3191,N_3067);
xor U3710 (N_3710,N_3447,N_2664);
and U3711 (N_3711,N_2724,N_3206);
nand U3712 (N_3712,N_2693,N_2901);
and U3713 (N_3713,N_3435,N_2949);
and U3714 (N_3714,N_2862,N_3423);
and U3715 (N_3715,N_2443,N_2617);
or U3716 (N_3716,N_2850,N_2622);
and U3717 (N_3717,N_3557,N_3327);
xnor U3718 (N_3718,N_2518,N_3308);
xor U3719 (N_3719,N_2492,N_2876);
and U3720 (N_3720,N_2609,N_3298);
nand U3721 (N_3721,N_2770,N_2983);
nor U3722 (N_3722,N_3428,N_2869);
nand U3723 (N_3723,N_2491,N_2906);
xor U3724 (N_3724,N_2634,N_3463);
and U3725 (N_3725,N_2782,N_3339);
xor U3726 (N_3726,N_2541,N_2579);
and U3727 (N_3727,N_3140,N_3151);
and U3728 (N_3728,N_3209,N_3219);
nor U3729 (N_3729,N_3087,N_2873);
nand U3730 (N_3730,N_2531,N_3545);
nor U3731 (N_3731,N_2771,N_2723);
and U3732 (N_3732,N_2514,N_3478);
or U3733 (N_3733,N_2826,N_2814);
xnor U3734 (N_3734,N_2592,N_3155);
nand U3735 (N_3735,N_3014,N_2865);
or U3736 (N_3736,N_3193,N_2932);
and U3737 (N_3737,N_3376,N_2583);
xnor U3738 (N_3738,N_3508,N_3434);
nor U3739 (N_3739,N_2907,N_2828);
xnor U3740 (N_3740,N_3064,N_2461);
xor U3741 (N_3741,N_2658,N_2400);
xnor U3742 (N_3742,N_2410,N_3003);
xor U3743 (N_3743,N_2859,N_3074);
nand U3744 (N_3744,N_2629,N_2415);
or U3745 (N_3745,N_2767,N_2451);
xor U3746 (N_3746,N_2893,N_2804);
nand U3747 (N_3747,N_3406,N_2516);
and U3748 (N_3748,N_3368,N_2950);
nor U3749 (N_3749,N_3196,N_3561);
or U3750 (N_3750,N_3413,N_3419);
or U3751 (N_3751,N_2802,N_2858);
nand U3752 (N_3752,N_3358,N_3501);
or U3753 (N_3753,N_3397,N_3523);
xnor U3754 (N_3754,N_2823,N_2868);
and U3755 (N_3755,N_2750,N_3516);
or U3756 (N_3756,N_2896,N_2821);
or U3757 (N_3757,N_3546,N_2479);
and U3758 (N_3758,N_3379,N_2480);
nor U3759 (N_3759,N_2470,N_3482);
xnor U3760 (N_3760,N_3026,N_3165);
nor U3761 (N_3761,N_2458,N_2532);
or U3762 (N_3762,N_3359,N_2957);
nand U3763 (N_3763,N_2905,N_2509);
and U3764 (N_3764,N_2818,N_2728);
and U3765 (N_3765,N_2967,N_3188);
nor U3766 (N_3766,N_2902,N_3141);
nor U3767 (N_3767,N_3100,N_2718);
or U3768 (N_3768,N_3486,N_2431);
nor U3769 (N_3769,N_3567,N_3432);
nor U3770 (N_3770,N_2848,N_2928);
xnor U3771 (N_3771,N_2879,N_2558);
or U3772 (N_3772,N_3378,N_3104);
and U3773 (N_3773,N_2841,N_2955);
nand U3774 (N_3774,N_3004,N_2553);
and U3775 (N_3775,N_2454,N_2605);
and U3776 (N_3776,N_2570,N_3460);
and U3777 (N_3777,N_2460,N_2698);
and U3778 (N_3778,N_3056,N_2819);
or U3779 (N_3779,N_2528,N_2809);
xor U3780 (N_3780,N_3370,N_2715);
and U3781 (N_3781,N_3253,N_2504);
and U3782 (N_3782,N_2618,N_2922);
nand U3783 (N_3783,N_2787,N_3542);
and U3784 (N_3784,N_3325,N_2542);
nand U3785 (N_3785,N_3238,N_2581);
nor U3786 (N_3786,N_2801,N_3381);
and U3787 (N_3787,N_3183,N_2736);
nor U3788 (N_3788,N_2852,N_3489);
and U3789 (N_3789,N_3512,N_3411);
or U3790 (N_3790,N_3083,N_2564);
or U3791 (N_3791,N_2401,N_2519);
xor U3792 (N_3792,N_3532,N_2523);
or U3793 (N_3793,N_2591,N_3029);
and U3794 (N_3794,N_3446,N_3479);
and U3795 (N_3795,N_2900,N_3458);
and U3796 (N_3796,N_3288,N_2799);
xor U3797 (N_3797,N_2638,N_2697);
nand U3798 (N_3798,N_2978,N_2652);
xor U3799 (N_3799,N_3293,N_2412);
nor U3800 (N_3800,N_3440,N_3513);
nand U3801 (N_3801,N_3137,N_2448);
and U3802 (N_3802,N_2627,N_3357);
nand U3803 (N_3803,N_3541,N_2436);
xnor U3804 (N_3804,N_3350,N_3492);
or U3805 (N_3805,N_3236,N_3170);
and U3806 (N_3806,N_2838,N_2597);
and U3807 (N_3807,N_2992,N_2798);
or U3808 (N_3808,N_2551,N_3371);
and U3809 (N_3809,N_3472,N_3052);
or U3810 (N_3810,N_2857,N_2986);
xor U3811 (N_3811,N_2899,N_3581);
nand U3812 (N_3812,N_2477,N_3000);
nor U3813 (N_3813,N_3534,N_2686);
nand U3814 (N_3814,N_3485,N_2433);
nor U3815 (N_3815,N_2927,N_3555);
nand U3816 (N_3816,N_3496,N_3331);
nand U3817 (N_3817,N_3242,N_3393);
nand U3818 (N_3818,N_2716,N_3564);
nor U3819 (N_3819,N_3093,N_2587);
xnor U3820 (N_3820,N_2925,N_2807);
xor U3821 (N_3821,N_3351,N_2878);
nand U3822 (N_3822,N_2834,N_2759);
nand U3823 (N_3823,N_3153,N_2565);
nor U3824 (N_3824,N_2473,N_2860);
or U3825 (N_3825,N_2830,N_2785);
nor U3826 (N_3826,N_2935,N_3574);
or U3827 (N_3827,N_3402,N_2667);
nand U3828 (N_3828,N_2720,N_2422);
and U3829 (N_3829,N_3572,N_3240);
nand U3830 (N_3830,N_3283,N_3504);
xor U3831 (N_3831,N_2447,N_3438);
nor U3832 (N_3832,N_2507,N_3178);
xor U3833 (N_3833,N_2998,N_3380);
and U3834 (N_3834,N_3257,N_3115);
or U3835 (N_3835,N_2526,N_2874);
and U3836 (N_3836,N_3556,N_2758);
and U3837 (N_3837,N_3076,N_2835);
nor U3838 (N_3838,N_2703,N_3234);
xnor U3839 (N_3839,N_3537,N_3018);
xor U3840 (N_3840,N_3246,N_2620);
nor U3841 (N_3841,N_2793,N_2499);
and U3842 (N_3842,N_2673,N_2854);
and U3843 (N_3843,N_2498,N_2926);
and U3844 (N_3844,N_3272,N_2440);
nor U3845 (N_3845,N_2914,N_2689);
nor U3846 (N_3846,N_2891,N_3275);
nor U3847 (N_3847,N_3375,N_2734);
nand U3848 (N_3848,N_2560,N_2623);
nor U3849 (N_3849,N_3075,N_3346);
or U3850 (N_3850,N_3215,N_2712);
and U3851 (N_3851,N_2585,N_2747);
and U3852 (N_3852,N_2863,N_3047);
nor U3853 (N_3853,N_2450,N_2488);
or U3854 (N_3854,N_3248,N_2903);
xor U3855 (N_3855,N_3261,N_3528);
xnor U3856 (N_3856,N_2660,N_2714);
or U3857 (N_3857,N_3596,N_3036);
nor U3858 (N_3858,N_3551,N_2556);
xor U3859 (N_3859,N_2656,N_2981);
xnor U3860 (N_3860,N_2886,N_3563);
nand U3861 (N_3861,N_3582,N_2657);
nand U3862 (N_3862,N_2536,N_2404);
nand U3863 (N_3863,N_3210,N_2446);
nand U3864 (N_3864,N_3013,N_3186);
nor U3865 (N_3865,N_2453,N_3373);
and U3866 (N_3866,N_2769,N_3354);
nor U3867 (N_3867,N_3129,N_3417);
and U3868 (N_3868,N_3300,N_2511);
nor U3869 (N_3869,N_3502,N_2641);
nor U3870 (N_3870,N_3326,N_3290);
nor U3871 (N_3871,N_3353,N_3090);
xor U3872 (N_3872,N_3344,N_3363);
and U3873 (N_3873,N_2615,N_2607);
xor U3874 (N_3874,N_3028,N_3519);
nor U3875 (N_3875,N_3032,N_3425);
xor U3876 (N_3876,N_3289,N_2952);
or U3877 (N_3877,N_2577,N_3583);
nor U3878 (N_3878,N_3558,N_3320);
nor U3879 (N_3879,N_2495,N_2500);
and U3880 (N_3880,N_3535,N_3525);
xor U3881 (N_3881,N_3152,N_3150);
and U3882 (N_3882,N_3343,N_2467);
nand U3883 (N_3883,N_3088,N_3466);
and U3884 (N_3884,N_3473,N_3207);
nor U3885 (N_3885,N_3030,N_2434);
and U3886 (N_3886,N_3459,N_3063);
nand U3887 (N_3887,N_2537,N_2764);
or U3888 (N_3888,N_2871,N_3164);
xnor U3889 (N_3889,N_2895,N_3017);
nor U3890 (N_3890,N_3384,N_3355);
and U3891 (N_3891,N_3410,N_3050);
and U3892 (N_3892,N_2610,N_3475);
nand U3893 (N_3893,N_3409,N_3252);
and U3894 (N_3894,N_3135,N_3571);
and U3895 (N_3895,N_3306,N_2420);
and U3896 (N_3896,N_3352,N_3589);
and U3897 (N_3897,N_2472,N_2910);
xnor U3898 (N_3898,N_3102,N_2960);
nor U3899 (N_3899,N_3569,N_2795);
or U3900 (N_3900,N_2582,N_2469);
nand U3901 (N_3901,N_2546,N_3190);
or U3902 (N_3902,N_3230,N_3329);
nand U3903 (N_3903,N_3530,N_3205);
nand U3904 (N_3904,N_2465,N_2822);
xnor U3905 (N_3905,N_3099,N_2547);
xnor U3906 (N_3906,N_2776,N_3361);
xnor U3907 (N_3907,N_3092,N_3105);
or U3908 (N_3908,N_3302,N_3503);
nand U3909 (N_3909,N_2678,N_3282);
nand U3910 (N_3910,N_2904,N_2725);
xor U3911 (N_3911,N_3314,N_2911);
or U3912 (N_3912,N_2442,N_2683);
and U3913 (N_3913,N_3345,N_2722);
nand U3914 (N_3914,N_2655,N_2428);
nor U3915 (N_3915,N_2444,N_3279);
or U3916 (N_3916,N_3176,N_3587);
nor U3917 (N_3917,N_3391,N_3416);
and U3918 (N_3918,N_2437,N_2774);
nand U3919 (N_3919,N_2554,N_2740);
nand U3920 (N_3920,N_2402,N_3046);
nand U3921 (N_3921,N_2598,N_3568);
or U3922 (N_3922,N_3388,N_3538);
or U3923 (N_3923,N_2919,N_2595);
nand U3924 (N_3924,N_3500,N_2692);
nand U3925 (N_3925,N_2997,N_3467);
or U3926 (N_3926,N_3147,N_3237);
and U3927 (N_3927,N_2590,N_2816);
nand U3928 (N_3928,N_2411,N_3126);
nand U3929 (N_3929,N_2681,N_2810);
nor U3930 (N_3930,N_3559,N_3316);
nand U3931 (N_3931,N_2567,N_2520);
xor U3932 (N_3932,N_2671,N_3578);
and U3933 (N_3933,N_3031,N_2885);
nand U3934 (N_3934,N_2755,N_3119);
nand U3935 (N_3935,N_2796,N_2435);
nand U3936 (N_3936,N_3362,N_2763);
and U3937 (N_3937,N_3208,N_2650);
or U3938 (N_3938,N_2596,N_2709);
and U3939 (N_3939,N_2694,N_3184);
or U3940 (N_3940,N_3167,N_3011);
or U3941 (N_3941,N_2975,N_3107);
nand U3942 (N_3942,N_3212,N_2912);
or U3943 (N_3943,N_2880,N_2929);
xnor U3944 (N_3944,N_3437,N_3055);
nor U3945 (N_3945,N_2632,N_3044);
xnor U3946 (N_3946,N_2672,N_2773);
or U3947 (N_3947,N_3595,N_2502);
and U3948 (N_3948,N_2644,N_2780);
and U3949 (N_3949,N_2653,N_2481);
nand U3950 (N_3950,N_2584,N_3313);
or U3951 (N_3951,N_2888,N_2619);
or U3952 (N_3952,N_2945,N_3057);
and U3953 (N_3953,N_2972,N_3022);
and U3954 (N_3954,N_3182,N_2861);
or U3955 (N_3955,N_2812,N_2628);
nor U3956 (N_3956,N_3158,N_2604);
nor U3957 (N_3957,N_3042,N_2930);
xor U3958 (N_3958,N_3328,N_3421);
or U3959 (N_3959,N_3024,N_3053);
nor U3960 (N_3960,N_2702,N_2974);
nand U3961 (N_3961,N_3204,N_3069);
nor U3962 (N_3962,N_2687,N_3318);
nand U3963 (N_3963,N_3580,N_3514);
nand U3964 (N_3964,N_2471,N_2484);
nand U3965 (N_3965,N_3250,N_2792);
or U3966 (N_3966,N_2883,N_3258);
and U3967 (N_3967,N_2958,N_2616);
and U3968 (N_3968,N_2940,N_3497);
or U3969 (N_3969,N_2497,N_3082);
nand U3970 (N_3970,N_3073,N_3133);
xnor U3971 (N_3971,N_3365,N_3008);
or U3972 (N_3972,N_2937,N_3274);
nand U3973 (N_3973,N_2866,N_3562);
and U3974 (N_3974,N_3012,N_2872);
or U3975 (N_3975,N_2521,N_3591);
nand U3976 (N_3976,N_2719,N_3465);
and U3977 (N_3977,N_3400,N_3217);
nor U3978 (N_3978,N_3094,N_3444);
and U3979 (N_3979,N_3139,N_3146);
nor U3980 (N_3980,N_2831,N_3278);
and U3981 (N_3981,N_2820,N_3526);
or U3982 (N_3982,N_2779,N_3060);
or U3983 (N_3983,N_3570,N_3065);
or U3984 (N_3984,N_3021,N_3403);
nor U3985 (N_3985,N_2639,N_3450);
and U3986 (N_3986,N_2426,N_2462);
and U3987 (N_3987,N_3436,N_2962);
nor U3988 (N_3988,N_2762,N_3392);
and U3989 (N_3989,N_3220,N_3445);
nor U3990 (N_3990,N_3520,N_2744);
nor U3991 (N_3991,N_2643,N_2976);
xor U3992 (N_3992,N_2494,N_2964);
or U3993 (N_3993,N_3084,N_3175);
or U3994 (N_3994,N_3366,N_3002);
nor U3995 (N_3995,N_3068,N_3264);
or U3996 (N_3996,N_2766,N_2419);
xnor U3997 (N_3997,N_2407,N_3456);
nand U3998 (N_3998,N_2984,N_2555);
nand U3999 (N_3999,N_3543,N_3241);
nor U4000 (N_4000,N_3189,N_3544);
nand U4001 (N_4001,N_3001,N_3061);
and U4002 (N_4002,N_2543,N_3399);
or U4003 (N_4003,N_2920,N_2705);
or U4004 (N_4004,N_2682,N_2513);
or U4005 (N_4005,N_3268,N_2635);
xnor U4006 (N_4006,N_2665,N_2909);
nor U4007 (N_4007,N_3225,N_3045);
nor U4008 (N_4008,N_3455,N_2761);
and U4009 (N_4009,N_2421,N_3174);
nor U4010 (N_4010,N_2993,N_2995);
and U4011 (N_4011,N_2559,N_3054);
or U4012 (N_4012,N_3127,N_3226);
nand U4013 (N_4013,N_3079,N_3511);
xnor U4014 (N_4014,N_3593,N_3342);
or U4015 (N_4015,N_3390,N_3281);
and U4016 (N_4016,N_3424,N_3249);
or U4017 (N_4017,N_3066,N_2668);
nor U4018 (N_4018,N_2892,N_2735);
and U4019 (N_4019,N_2539,N_2423);
or U4020 (N_4020,N_2600,N_3304);
or U4021 (N_4021,N_3506,N_2696);
nand U4022 (N_4022,N_2847,N_3451);
nor U4023 (N_4023,N_2601,N_3071);
and U4024 (N_4024,N_3138,N_2666);
nand U4025 (N_4025,N_2708,N_3038);
and U4026 (N_4026,N_2800,N_3265);
or U4027 (N_4027,N_2545,N_2923);
nand U4028 (N_4028,N_2637,N_2602);
or U4029 (N_4029,N_2966,N_2706);
nand U4030 (N_4030,N_2550,N_2409);
xor U4031 (N_4031,N_3020,N_3309);
or U4032 (N_4032,N_3349,N_2890);
xnor U4033 (N_4033,N_3035,N_3468);
xnor U4034 (N_4034,N_3303,N_3159);
xor U4035 (N_4035,N_2938,N_2788);
nor U4036 (N_4036,N_2478,N_2576);
nand U4037 (N_4037,N_2754,N_3470);
xor U4038 (N_4038,N_3586,N_3145);
xnor U4039 (N_4039,N_3491,N_2717);
and U4040 (N_4040,N_2989,N_3454);
nand U4041 (N_4041,N_3483,N_3301);
or U4042 (N_4042,N_2700,N_3161);
nand U4043 (N_4043,N_3407,N_2490);
nand U4044 (N_4044,N_3453,N_3311);
nand U4045 (N_4045,N_2990,N_2662);
and U4046 (N_4046,N_2496,N_2599);
or U4047 (N_4047,N_3422,N_3484);
nand U4048 (N_4048,N_3273,N_2603);
or U4049 (N_4049,N_3307,N_2768);
and U4050 (N_4050,N_2760,N_2611);
nor U4051 (N_4051,N_2455,N_2917);
or U4052 (N_4052,N_2416,N_2908);
xor U4053 (N_4053,N_3548,N_3043);
nor U4054 (N_4054,N_3091,N_3157);
and U4055 (N_4055,N_2731,N_2613);
xor U4056 (N_4056,N_2951,N_2737);
xor U4057 (N_4057,N_2417,N_2742);
or U4058 (N_4058,N_2851,N_2503);
nor U4059 (N_4059,N_3059,N_3469);
and U4060 (N_4060,N_3085,N_3080);
nor U4061 (N_4061,N_3131,N_2646);
nand U4062 (N_4062,N_2832,N_2606);
xor U4063 (N_4063,N_2535,N_2663);
xor U4064 (N_4064,N_3034,N_3039);
nand U4065 (N_4065,N_2540,N_3201);
xor U4066 (N_4066,N_3317,N_3041);
nand U4067 (N_4067,N_3120,N_3341);
nor U4068 (N_4068,N_3382,N_2640);
nand U4069 (N_4069,N_3239,N_2877);
nor U4070 (N_4070,N_3025,N_2476);
or U4071 (N_4071,N_3367,N_2965);
and U4072 (N_4072,N_2797,N_3539);
and U4073 (N_4073,N_2648,N_3033);
nor U4074 (N_4074,N_3277,N_3494);
xnor U4075 (N_4075,N_2685,N_2979);
nand U4076 (N_4076,N_3337,N_2808);
nor U4077 (N_4077,N_3319,N_3200);
and U4078 (N_4078,N_3404,N_2475);
or U4079 (N_4079,N_3566,N_3394);
nand U4080 (N_4080,N_2711,N_3565);
xnor U4081 (N_4081,N_2566,N_3515);
nand U4082 (N_4082,N_2743,N_2506);
nor U4083 (N_4083,N_3477,N_2466);
or U4084 (N_4084,N_2563,N_2486);
nor U4085 (N_4085,N_2968,N_3431);
and U4086 (N_4086,N_2777,N_2882);
nand U4087 (N_4087,N_3585,N_2578);
and U4088 (N_4088,N_2530,N_2842);
xnor U4089 (N_4089,N_2756,N_2552);
or U4090 (N_4090,N_2973,N_2414);
xor U4091 (N_4091,N_3114,N_2918);
and U4092 (N_4092,N_2573,N_3442);
xor U4093 (N_4093,N_3118,N_2575);
xnor U4094 (N_4094,N_3106,N_3096);
nand U4095 (N_4095,N_3457,N_2748);
xor U4096 (N_4096,N_3439,N_2489);
and U4097 (N_4097,N_3322,N_2954);
nor U4098 (N_4098,N_3488,N_3347);
and U4099 (N_4099,N_3016,N_2953);
nand U4100 (N_4100,N_3192,N_2688);
nand U4101 (N_4101,N_3218,N_2784);
nor U4102 (N_4102,N_3336,N_3521);
or U4103 (N_4103,N_3180,N_3334);
or U4104 (N_4104,N_2947,N_3427);
xnor U4105 (N_4105,N_2994,N_2746);
nand U4106 (N_4106,N_2721,N_3110);
or U4107 (N_4107,N_2733,N_3296);
xnor U4108 (N_4108,N_2855,N_3213);
nand U4109 (N_4109,N_3474,N_2898);
xor U4110 (N_4110,N_2963,N_2811);
or U4111 (N_4111,N_2438,N_3324);
and U4112 (N_4112,N_2739,N_2614);
nor U4113 (N_4113,N_2593,N_3522);
xor U4114 (N_4114,N_3597,N_2642);
nand U4115 (N_4115,N_2791,N_2654);
xnor U4116 (N_4116,N_3374,N_3171);
and U4117 (N_4117,N_3594,N_3048);
nor U4118 (N_4118,N_3441,N_2824);
or U4119 (N_4119,N_3448,N_2621);
nand U4120 (N_4120,N_2589,N_2790);
nand U4121 (N_4121,N_3305,N_2897);
xor U4122 (N_4122,N_3010,N_2501);
nand U4123 (N_4123,N_3223,N_3227);
nor U4124 (N_4124,N_2463,N_3518);
nor U4125 (N_4125,N_2840,N_2889);
nor U4126 (N_4126,N_2944,N_2959);
nand U4127 (N_4127,N_3098,N_3122);
or U4128 (N_4128,N_3185,N_3372);
xor U4129 (N_4129,N_2630,N_2680);
or U4130 (N_4130,N_3169,N_3547);
or U4131 (N_4131,N_2833,N_2837);
xnor U4132 (N_4132,N_2943,N_2817);
xnor U4133 (N_4133,N_2441,N_2772);
or U4134 (N_4134,N_2427,N_2894);
and U4135 (N_4135,N_2439,N_2805);
nor U4136 (N_4136,N_3505,N_3412);
and U4137 (N_4137,N_3244,N_3576);
nor U4138 (N_4138,N_3228,N_2406);
xor U4139 (N_4139,N_2931,N_2403);
and U4140 (N_4140,N_3233,N_3540);
or U4141 (N_4141,N_2794,N_3579);
xor U4142 (N_4142,N_2659,N_3284);
and U4143 (N_4143,N_3599,N_3089);
or U4144 (N_4144,N_2612,N_2445);
nor U4145 (N_4145,N_2971,N_3173);
and U4146 (N_4146,N_2864,N_2845);
nand U4147 (N_4147,N_3449,N_2510);
nor U4148 (N_4148,N_2839,N_3117);
or U4149 (N_4149,N_3292,N_2562);
and U4150 (N_4150,N_2487,N_2870);
nand U4151 (N_4151,N_2525,N_3276);
or U4152 (N_4152,N_3095,N_2669);
xnor U4153 (N_4153,N_2633,N_2980);
or U4154 (N_4154,N_3286,N_2836);
nor U4155 (N_4155,N_3577,N_3243);
nor U4156 (N_4156,N_3162,N_3263);
nand U4157 (N_4157,N_2588,N_3321);
and U4158 (N_4158,N_2881,N_3058);
xnor U4159 (N_4159,N_3498,N_2846);
nand U4160 (N_4160,N_2933,N_2985);
nor U4161 (N_4161,N_2887,N_3111);
xor U4162 (N_4162,N_2533,N_2987);
or U4163 (N_4163,N_3415,N_2517);
or U4164 (N_4164,N_3124,N_3247);
xnor U4165 (N_4165,N_3369,N_2751);
xnor U4166 (N_4166,N_3005,N_3510);
xnor U4167 (N_4167,N_3386,N_2459);
and U4168 (N_4168,N_2557,N_3255);
nand U4169 (N_4169,N_2684,N_3136);
nand U4170 (N_4170,N_2624,N_2544);
xnor U4171 (N_4171,N_2752,N_3194);
and U4172 (N_4172,N_2856,N_3116);
nand U4173 (N_4173,N_3299,N_2843);
nor U4174 (N_4174,N_3254,N_3509);
and U4175 (N_4175,N_2674,N_3452);
nand U4176 (N_4176,N_3461,N_3480);
nor U4177 (N_4177,N_3383,N_3262);
nand U4178 (N_4178,N_3166,N_2418);
or U4179 (N_4179,N_3027,N_3221);
or U4180 (N_4180,N_3143,N_3575);
and U4181 (N_4181,N_3121,N_2690);
and U4182 (N_4182,N_2707,N_3179);
nor U4183 (N_4183,N_2493,N_2452);
xnor U4184 (N_4184,N_2729,N_3430);
and U4185 (N_4185,N_2738,N_2745);
nor U4186 (N_4186,N_3408,N_3216);
and U4187 (N_4187,N_2789,N_2649);
or U4188 (N_4188,N_2429,N_2996);
nand U4189 (N_4189,N_2468,N_2574);
nor U4190 (N_4190,N_2999,N_3420);
nor U4191 (N_4191,N_2548,N_3006);
nor U4192 (N_4192,N_2456,N_2645);
and U4193 (N_4193,N_2571,N_2916);
and U4194 (N_4194,N_3554,N_3588);
xnor U4195 (N_4195,N_3019,N_3335);
and U4196 (N_4196,N_3396,N_3549);
nand U4197 (N_4197,N_3231,N_3387);
and U4198 (N_4198,N_2961,N_3364);
nand U4199 (N_4199,N_2594,N_3144);
and U4200 (N_4200,N_2550,N_3226);
nand U4201 (N_4201,N_3181,N_2716);
and U4202 (N_4202,N_2572,N_2431);
xor U4203 (N_4203,N_3411,N_3023);
or U4204 (N_4204,N_2875,N_3460);
nand U4205 (N_4205,N_2805,N_3172);
or U4206 (N_4206,N_2598,N_2647);
nor U4207 (N_4207,N_2689,N_2458);
or U4208 (N_4208,N_2729,N_2707);
nand U4209 (N_4209,N_3243,N_3149);
or U4210 (N_4210,N_2570,N_2775);
or U4211 (N_4211,N_2836,N_3261);
nor U4212 (N_4212,N_3018,N_3576);
or U4213 (N_4213,N_3025,N_2896);
nor U4214 (N_4214,N_3358,N_2972);
and U4215 (N_4215,N_3259,N_2569);
nand U4216 (N_4216,N_3331,N_3111);
nor U4217 (N_4217,N_2761,N_3250);
and U4218 (N_4218,N_2663,N_2482);
and U4219 (N_4219,N_2954,N_3025);
or U4220 (N_4220,N_2468,N_2680);
or U4221 (N_4221,N_3227,N_2485);
or U4222 (N_4222,N_3562,N_3325);
xnor U4223 (N_4223,N_2863,N_2646);
xnor U4224 (N_4224,N_3006,N_2408);
xor U4225 (N_4225,N_3347,N_3261);
nand U4226 (N_4226,N_2672,N_2531);
nor U4227 (N_4227,N_2644,N_2577);
xor U4228 (N_4228,N_2505,N_3028);
nor U4229 (N_4229,N_3256,N_3288);
nor U4230 (N_4230,N_2913,N_3102);
or U4231 (N_4231,N_3102,N_2515);
nor U4232 (N_4232,N_2467,N_2533);
or U4233 (N_4233,N_3038,N_2844);
nand U4234 (N_4234,N_2876,N_3120);
and U4235 (N_4235,N_2979,N_2690);
nor U4236 (N_4236,N_3315,N_2624);
or U4237 (N_4237,N_3376,N_2658);
nand U4238 (N_4238,N_2433,N_2766);
xor U4239 (N_4239,N_2829,N_2566);
nand U4240 (N_4240,N_2568,N_2541);
or U4241 (N_4241,N_2887,N_2715);
or U4242 (N_4242,N_3524,N_3113);
xnor U4243 (N_4243,N_3572,N_2810);
nand U4244 (N_4244,N_2638,N_2931);
and U4245 (N_4245,N_3037,N_3380);
and U4246 (N_4246,N_3196,N_2861);
nor U4247 (N_4247,N_2558,N_2896);
or U4248 (N_4248,N_2478,N_2797);
and U4249 (N_4249,N_3416,N_2652);
and U4250 (N_4250,N_2752,N_2452);
xnor U4251 (N_4251,N_3281,N_3379);
or U4252 (N_4252,N_3126,N_3451);
or U4253 (N_4253,N_3240,N_3471);
xnor U4254 (N_4254,N_2875,N_2721);
nand U4255 (N_4255,N_3267,N_2408);
nor U4256 (N_4256,N_3402,N_2897);
nand U4257 (N_4257,N_2744,N_3487);
and U4258 (N_4258,N_2702,N_3135);
xor U4259 (N_4259,N_2463,N_3147);
nand U4260 (N_4260,N_3224,N_3153);
nand U4261 (N_4261,N_3558,N_3475);
or U4262 (N_4262,N_2840,N_3106);
nand U4263 (N_4263,N_2865,N_3175);
nand U4264 (N_4264,N_2970,N_2559);
or U4265 (N_4265,N_3476,N_2644);
or U4266 (N_4266,N_2809,N_3229);
nand U4267 (N_4267,N_3436,N_3278);
and U4268 (N_4268,N_2664,N_3415);
nand U4269 (N_4269,N_3482,N_3402);
nor U4270 (N_4270,N_2767,N_3370);
nor U4271 (N_4271,N_3185,N_2684);
and U4272 (N_4272,N_3094,N_3414);
or U4273 (N_4273,N_2467,N_3454);
nor U4274 (N_4274,N_2608,N_3380);
nor U4275 (N_4275,N_3169,N_2426);
nand U4276 (N_4276,N_2513,N_3070);
xor U4277 (N_4277,N_3018,N_2877);
xor U4278 (N_4278,N_2849,N_2588);
nor U4279 (N_4279,N_3371,N_3528);
xor U4280 (N_4280,N_2940,N_2982);
nor U4281 (N_4281,N_3349,N_3452);
nand U4282 (N_4282,N_3281,N_3409);
nand U4283 (N_4283,N_2540,N_2919);
nor U4284 (N_4284,N_3505,N_3263);
xnor U4285 (N_4285,N_3370,N_3369);
nand U4286 (N_4286,N_2481,N_3595);
and U4287 (N_4287,N_3471,N_2763);
or U4288 (N_4288,N_2816,N_2428);
xnor U4289 (N_4289,N_3000,N_3371);
and U4290 (N_4290,N_3491,N_3356);
nor U4291 (N_4291,N_3384,N_2501);
nor U4292 (N_4292,N_3438,N_2500);
and U4293 (N_4293,N_3391,N_2565);
and U4294 (N_4294,N_2824,N_3454);
nor U4295 (N_4295,N_3512,N_3486);
and U4296 (N_4296,N_2620,N_2595);
or U4297 (N_4297,N_3136,N_2419);
nor U4298 (N_4298,N_2762,N_3451);
or U4299 (N_4299,N_2426,N_3545);
nand U4300 (N_4300,N_3112,N_2757);
or U4301 (N_4301,N_2705,N_2421);
nor U4302 (N_4302,N_3544,N_2532);
nand U4303 (N_4303,N_2566,N_3247);
xnor U4304 (N_4304,N_3496,N_3088);
nor U4305 (N_4305,N_3256,N_3221);
or U4306 (N_4306,N_3064,N_3576);
or U4307 (N_4307,N_3260,N_2754);
or U4308 (N_4308,N_2976,N_2631);
xor U4309 (N_4309,N_3250,N_2476);
or U4310 (N_4310,N_2562,N_3290);
or U4311 (N_4311,N_2442,N_3033);
or U4312 (N_4312,N_2626,N_2661);
nand U4313 (N_4313,N_3239,N_3232);
or U4314 (N_4314,N_3389,N_3023);
and U4315 (N_4315,N_3096,N_3298);
and U4316 (N_4316,N_2755,N_3034);
nand U4317 (N_4317,N_3462,N_2729);
xnor U4318 (N_4318,N_3250,N_3552);
nand U4319 (N_4319,N_3512,N_3383);
nor U4320 (N_4320,N_3123,N_2495);
and U4321 (N_4321,N_3261,N_2857);
or U4322 (N_4322,N_2645,N_2750);
xnor U4323 (N_4323,N_2812,N_2516);
or U4324 (N_4324,N_3438,N_3234);
xor U4325 (N_4325,N_2951,N_3091);
or U4326 (N_4326,N_2797,N_3061);
xor U4327 (N_4327,N_2791,N_3567);
or U4328 (N_4328,N_3172,N_3344);
or U4329 (N_4329,N_3544,N_2597);
xor U4330 (N_4330,N_2693,N_3129);
xnor U4331 (N_4331,N_3265,N_2563);
and U4332 (N_4332,N_3372,N_2818);
xnor U4333 (N_4333,N_3318,N_3269);
nor U4334 (N_4334,N_3568,N_2423);
and U4335 (N_4335,N_2887,N_2418);
or U4336 (N_4336,N_3332,N_3286);
or U4337 (N_4337,N_2884,N_3163);
xor U4338 (N_4338,N_2709,N_3462);
and U4339 (N_4339,N_2423,N_3405);
and U4340 (N_4340,N_3192,N_2406);
or U4341 (N_4341,N_2735,N_2686);
and U4342 (N_4342,N_3529,N_2469);
nor U4343 (N_4343,N_2558,N_2572);
xor U4344 (N_4344,N_2415,N_3352);
or U4345 (N_4345,N_2626,N_3101);
nand U4346 (N_4346,N_2906,N_2951);
or U4347 (N_4347,N_3461,N_3152);
nand U4348 (N_4348,N_3177,N_3524);
nand U4349 (N_4349,N_3545,N_2882);
or U4350 (N_4350,N_2787,N_3431);
xnor U4351 (N_4351,N_2997,N_2509);
or U4352 (N_4352,N_3306,N_2977);
nand U4353 (N_4353,N_3406,N_2441);
nor U4354 (N_4354,N_2451,N_3176);
or U4355 (N_4355,N_2918,N_2791);
xor U4356 (N_4356,N_3475,N_3349);
and U4357 (N_4357,N_3396,N_3397);
and U4358 (N_4358,N_2902,N_2424);
nand U4359 (N_4359,N_3398,N_2493);
nor U4360 (N_4360,N_3109,N_3003);
and U4361 (N_4361,N_3156,N_3387);
or U4362 (N_4362,N_2418,N_3006);
nand U4363 (N_4363,N_3599,N_3330);
xnor U4364 (N_4364,N_2539,N_3352);
or U4365 (N_4365,N_3161,N_2576);
nor U4366 (N_4366,N_3347,N_2460);
and U4367 (N_4367,N_2911,N_2553);
xor U4368 (N_4368,N_2833,N_2960);
nor U4369 (N_4369,N_2818,N_3148);
xnor U4370 (N_4370,N_3501,N_3516);
nor U4371 (N_4371,N_2906,N_3225);
xor U4372 (N_4372,N_3562,N_3277);
nor U4373 (N_4373,N_3211,N_3332);
xnor U4374 (N_4374,N_2724,N_3466);
or U4375 (N_4375,N_2637,N_3281);
nand U4376 (N_4376,N_3237,N_3063);
and U4377 (N_4377,N_2406,N_2512);
nor U4378 (N_4378,N_2561,N_3353);
and U4379 (N_4379,N_2402,N_3284);
and U4380 (N_4380,N_2772,N_2455);
nor U4381 (N_4381,N_2888,N_3593);
xnor U4382 (N_4382,N_2725,N_3509);
nor U4383 (N_4383,N_2432,N_3376);
and U4384 (N_4384,N_2430,N_3413);
and U4385 (N_4385,N_3516,N_3204);
nand U4386 (N_4386,N_2549,N_3322);
and U4387 (N_4387,N_2493,N_3590);
nor U4388 (N_4388,N_3128,N_3007);
nand U4389 (N_4389,N_2523,N_2532);
nor U4390 (N_4390,N_2947,N_3150);
and U4391 (N_4391,N_3014,N_2612);
and U4392 (N_4392,N_2934,N_3132);
nor U4393 (N_4393,N_3394,N_3286);
xnor U4394 (N_4394,N_3191,N_3585);
nand U4395 (N_4395,N_2628,N_2514);
or U4396 (N_4396,N_3141,N_2579);
and U4397 (N_4397,N_3170,N_3075);
nand U4398 (N_4398,N_2851,N_3301);
xor U4399 (N_4399,N_3038,N_3419);
xor U4400 (N_4400,N_3207,N_3388);
or U4401 (N_4401,N_3212,N_3168);
nand U4402 (N_4402,N_2650,N_3331);
and U4403 (N_4403,N_2819,N_2712);
nand U4404 (N_4404,N_3328,N_3506);
nor U4405 (N_4405,N_3379,N_3477);
nor U4406 (N_4406,N_3518,N_2596);
nor U4407 (N_4407,N_2601,N_3400);
xor U4408 (N_4408,N_2782,N_2827);
or U4409 (N_4409,N_2626,N_3495);
and U4410 (N_4410,N_2406,N_2888);
xnor U4411 (N_4411,N_2551,N_2827);
and U4412 (N_4412,N_2642,N_2912);
nand U4413 (N_4413,N_2447,N_3305);
and U4414 (N_4414,N_3077,N_2571);
xor U4415 (N_4415,N_2948,N_3475);
xor U4416 (N_4416,N_2433,N_2787);
nand U4417 (N_4417,N_2498,N_2430);
nand U4418 (N_4418,N_3090,N_3340);
xor U4419 (N_4419,N_3101,N_3277);
or U4420 (N_4420,N_3514,N_3340);
nor U4421 (N_4421,N_3336,N_2965);
or U4422 (N_4422,N_3323,N_3332);
and U4423 (N_4423,N_2547,N_3322);
and U4424 (N_4424,N_3599,N_3562);
xor U4425 (N_4425,N_2792,N_3374);
or U4426 (N_4426,N_3579,N_3287);
nand U4427 (N_4427,N_2750,N_3045);
and U4428 (N_4428,N_2793,N_3540);
and U4429 (N_4429,N_2914,N_2783);
or U4430 (N_4430,N_2671,N_2574);
nor U4431 (N_4431,N_2857,N_3086);
nand U4432 (N_4432,N_2451,N_2429);
or U4433 (N_4433,N_2701,N_2731);
or U4434 (N_4434,N_3321,N_3178);
nand U4435 (N_4435,N_2604,N_2763);
nand U4436 (N_4436,N_3072,N_2409);
nand U4437 (N_4437,N_2500,N_3372);
nor U4438 (N_4438,N_3072,N_2876);
nor U4439 (N_4439,N_2715,N_2459);
nand U4440 (N_4440,N_3008,N_3304);
nand U4441 (N_4441,N_2470,N_2456);
or U4442 (N_4442,N_3013,N_2490);
or U4443 (N_4443,N_2654,N_2923);
and U4444 (N_4444,N_3060,N_2913);
and U4445 (N_4445,N_3341,N_3504);
and U4446 (N_4446,N_3348,N_2797);
xnor U4447 (N_4447,N_2540,N_3058);
and U4448 (N_4448,N_3230,N_2677);
xor U4449 (N_4449,N_3185,N_2828);
and U4450 (N_4450,N_3332,N_2667);
or U4451 (N_4451,N_3462,N_3091);
nand U4452 (N_4452,N_2411,N_3518);
nor U4453 (N_4453,N_3048,N_2495);
and U4454 (N_4454,N_3005,N_3125);
xor U4455 (N_4455,N_2749,N_2733);
xor U4456 (N_4456,N_2764,N_2559);
or U4457 (N_4457,N_2476,N_3051);
and U4458 (N_4458,N_3507,N_2425);
xor U4459 (N_4459,N_3510,N_2688);
nand U4460 (N_4460,N_2489,N_2675);
or U4461 (N_4461,N_2628,N_3147);
nand U4462 (N_4462,N_3087,N_3193);
and U4463 (N_4463,N_2970,N_2706);
and U4464 (N_4464,N_3549,N_3513);
or U4465 (N_4465,N_2936,N_3429);
or U4466 (N_4466,N_3025,N_2982);
nand U4467 (N_4467,N_2819,N_3542);
and U4468 (N_4468,N_3555,N_2736);
and U4469 (N_4469,N_3067,N_3555);
nor U4470 (N_4470,N_3145,N_3495);
or U4471 (N_4471,N_3396,N_2674);
nor U4472 (N_4472,N_2854,N_3046);
nand U4473 (N_4473,N_3039,N_2503);
nor U4474 (N_4474,N_2514,N_3323);
nor U4475 (N_4475,N_2778,N_3540);
xor U4476 (N_4476,N_3275,N_2443);
nand U4477 (N_4477,N_3431,N_3298);
nand U4478 (N_4478,N_3194,N_2501);
nand U4479 (N_4479,N_3015,N_2852);
nand U4480 (N_4480,N_3554,N_2926);
nor U4481 (N_4481,N_3524,N_3254);
or U4482 (N_4482,N_2940,N_2515);
xnor U4483 (N_4483,N_2560,N_2586);
xnor U4484 (N_4484,N_2760,N_3428);
nor U4485 (N_4485,N_2875,N_3346);
and U4486 (N_4486,N_3210,N_2989);
or U4487 (N_4487,N_2870,N_3060);
or U4488 (N_4488,N_3397,N_3466);
nor U4489 (N_4489,N_3558,N_2431);
nand U4490 (N_4490,N_2652,N_3593);
xnor U4491 (N_4491,N_2975,N_2540);
and U4492 (N_4492,N_3369,N_2572);
xor U4493 (N_4493,N_2431,N_3168);
nand U4494 (N_4494,N_3105,N_3365);
nor U4495 (N_4495,N_3317,N_3138);
xor U4496 (N_4496,N_3284,N_2951);
and U4497 (N_4497,N_2497,N_2792);
nand U4498 (N_4498,N_2991,N_3504);
nand U4499 (N_4499,N_2936,N_2928);
or U4500 (N_4500,N_3362,N_3023);
and U4501 (N_4501,N_2596,N_2774);
and U4502 (N_4502,N_2687,N_3506);
nor U4503 (N_4503,N_3421,N_2570);
nor U4504 (N_4504,N_3082,N_2630);
or U4505 (N_4505,N_2748,N_3172);
or U4506 (N_4506,N_3216,N_2797);
or U4507 (N_4507,N_3469,N_2523);
and U4508 (N_4508,N_2661,N_3434);
xnor U4509 (N_4509,N_3510,N_3468);
and U4510 (N_4510,N_2425,N_3030);
and U4511 (N_4511,N_2897,N_2554);
or U4512 (N_4512,N_3174,N_2850);
nor U4513 (N_4513,N_3436,N_2904);
nor U4514 (N_4514,N_2720,N_2760);
xor U4515 (N_4515,N_2645,N_3511);
or U4516 (N_4516,N_3107,N_2505);
nor U4517 (N_4517,N_2519,N_3046);
nor U4518 (N_4518,N_3188,N_3409);
xor U4519 (N_4519,N_2520,N_2835);
and U4520 (N_4520,N_2506,N_3125);
xnor U4521 (N_4521,N_2770,N_2866);
or U4522 (N_4522,N_2927,N_2872);
nor U4523 (N_4523,N_2885,N_2546);
nand U4524 (N_4524,N_2897,N_3289);
and U4525 (N_4525,N_2439,N_2843);
and U4526 (N_4526,N_3465,N_2744);
and U4527 (N_4527,N_2943,N_2611);
or U4528 (N_4528,N_3426,N_3163);
xor U4529 (N_4529,N_2414,N_3381);
xor U4530 (N_4530,N_3122,N_3239);
xor U4531 (N_4531,N_2988,N_2753);
and U4532 (N_4532,N_3379,N_3214);
and U4533 (N_4533,N_3093,N_2533);
xor U4534 (N_4534,N_3507,N_2504);
nand U4535 (N_4535,N_3251,N_3158);
nand U4536 (N_4536,N_3378,N_3366);
xor U4537 (N_4537,N_2783,N_3235);
nor U4538 (N_4538,N_2497,N_2875);
nand U4539 (N_4539,N_3490,N_3371);
xnor U4540 (N_4540,N_3511,N_2649);
or U4541 (N_4541,N_3157,N_2624);
or U4542 (N_4542,N_3421,N_2517);
or U4543 (N_4543,N_2916,N_3495);
or U4544 (N_4544,N_3466,N_2813);
or U4545 (N_4545,N_3421,N_2581);
and U4546 (N_4546,N_2579,N_2775);
or U4547 (N_4547,N_3426,N_2526);
or U4548 (N_4548,N_2656,N_3150);
and U4549 (N_4549,N_2408,N_2784);
or U4550 (N_4550,N_3375,N_2454);
xor U4551 (N_4551,N_3402,N_3171);
nand U4552 (N_4552,N_3403,N_3335);
xor U4553 (N_4553,N_3482,N_3383);
xor U4554 (N_4554,N_3058,N_3073);
xnor U4555 (N_4555,N_2860,N_3088);
nor U4556 (N_4556,N_3294,N_3468);
nand U4557 (N_4557,N_3467,N_3080);
nor U4558 (N_4558,N_2684,N_3249);
xor U4559 (N_4559,N_2825,N_3088);
nand U4560 (N_4560,N_3153,N_3068);
or U4561 (N_4561,N_2562,N_2853);
and U4562 (N_4562,N_3049,N_3405);
or U4563 (N_4563,N_2632,N_2982);
and U4564 (N_4564,N_2472,N_3087);
and U4565 (N_4565,N_2941,N_3276);
and U4566 (N_4566,N_3574,N_3390);
or U4567 (N_4567,N_2926,N_3423);
or U4568 (N_4568,N_3123,N_3157);
xor U4569 (N_4569,N_3523,N_3518);
nor U4570 (N_4570,N_2914,N_2664);
nand U4571 (N_4571,N_3363,N_2576);
or U4572 (N_4572,N_3183,N_3195);
nor U4573 (N_4573,N_3515,N_2692);
or U4574 (N_4574,N_2706,N_3576);
nand U4575 (N_4575,N_2468,N_2611);
nor U4576 (N_4576,N_2815,N_3476);
or U4577 (N_4577,N_3251,N_3152);
xor U4578 (N_4578,N_3005,N_2532);
xnor U4579 (N_4579,N_2665,N_2997);
xnor U4580 (N_4580,N_3421,N_2776);
and U4581 (N_4581,N_2487,N_2416);
or U4582 (N_4582,N_3169,N_3118);
or U4583 (N_4583,N_3150,N_3577);
xor U4584 (N_4584,N_3360,N_2502);
xor U4585 (N_4585,N_2844,N_2749);
nand U4586 (N_4586,N_3532,N_3267);
or U4587 (N_4587,N_2467,N_2712);
and U4588 (N_4588,N_3029,N_2741);
and U4589 (N_4589,N_3040,N_3104);
or U4590 (N_4590,N_2942,N_3200);
and U4591 (N_4591,N_3057,N_2558);
xor U4592 (N_4592,N_3424,N_2490);
xnor U4593 (N_4593,N_2566,N_2968);
xor U4594 (N_4594,N_3167,N_3077);
nand U4595 (N_4595,N_3362,N_3388);
or U4596 (N_4596,N_2964,N_3161);
or U4597 (N_4597,N_3176,N_2411);
and U4598 (N_4598,N_2551,N_3327);
or U4599 (N_4599,N_2478,N_2528);
and U4600 (N_4600,N_2407,N_3085);
or U4601 (N_4601,N_3241,N_3343);
nand U4602 (N_4602,N_3128,N_2418);
xor U4603 (N_4603,N_3557,N_3085);
and U4604 (N_4604,N_2716,N_2553);
nor U4605 (N_4605,N_3477,N_2836);
or U4606 (N_4606,N_2906,N_2755);
xnor U4607 (N_4607,N_3323,N_3535);
nor U4608 (N_4608,N_3303,N_3362);
nor U4609 (N_4609,N_2687,N_3143);
and U4610 (N_4610,N_2670,N_2790);
or U4611 (N_4611,N_3495,N_2702);
and U4612 (N_4612,N_2959,N_2641);
and U4613 (N_4613,N_2731,N_3407);
xnor U4614 (N_4614,N_3171,N_2738);
nand U4615 (N_4615,N_2618,N_2520);
nand U4616 (N_4616,N_3435,N_2529);
nor U4617 (N_4617,N_2698,N_3561);
xnor U4618 (N_4618,N_2612,N_3065);
or U4619 (N_4619,N_3044,N_3407);
nor U4620 (N_4620,N_2502,N_3418);
and U4621 (N_4621,N_2847,N_3239);
nand U4622 (N_4622,N_3460,N_3129);
xnor U4623 (N_4623,N_3259,N_2674);
nor U4624 (N_4624,N_3465,N_2692);
nor U4625 (N_4625,N_2993,N_2474);
xor U4626 (N_4626,N_3223,N_3511);
and U4627 (N_4627,N_2702,N_2774);
nor U4628 (N_4628,N_3551,N_3198);
xor U4629 (N_4629,N_2710,N_2615);
or U4630 (N_4630,N_2424,N_3476);
and U4631 (N_4631,N_3027,N_2618);
nand U4632 (N_4632,N_3152,N_3208);
xor U4633 (N_4633,N_3324,N_2504);
and U4634 (N_4634,N_3478,N_3480);
or U4635 (N_4635,N_3583,N_2936);
nand U4636 (N_4636,N_2916,N_2745);
nor U4637 (N_4637,N_2781,N_3426);
xor U4638 (N_4638,N_2508,N_3231);
or U4639 (N_4639,N_2653,N_3340);
nand U4640 (N_4640,N_3164,N_3298);
nor U4641 (N_4641,N_2591,N_3247);
and U4642 (N_4642,N_2733,N_3468);
or U4643 (N_4643,N_3072,N_3248);
xor U4644 (N_4644,N_2612,N_2472);
nor U4645 (N_4645,N_3442,N_3185);
and U4646 (N_4646,N_2711,N_3588);
xor U4647 (N_4647,N_2992,N_3156);
nand U4648 (N_4648,N_3478,N_3441);
or U4649 (N_4649,N_2796,N_2893);
nand U4650 (N_4650,N_2759,N_2816);
xnor U4651 (N_4651,N_3076,N_2710);
nand U4652 (N_4652,N_3370,N_2737);
nor U4653 (N_4653,N_2496,N_3013);
nand U4654 (N_4654,N_2749,N_2983);
or U4655 (N_4655,N_2507,N_3195);
or U4656 (N_4656,N_3265,N_3080);
nor U4657 (N_4657,N_3297,N_3296);
or U4658 (N_4658,N_2762,N_2412);
and U4659 (N_4659,N_2461,N_3265);
nand U4660 (N_4660,N_3071,N_3512);
nor U4661 (N_4661,N_3522,N_3480);
and U4662 (N_4662,N_2697,N_2520);
and U4663 (N_4663,N_3351,N_3258);
xor U4664 (N_4664,N_3056,N_3206);
nor U4665 (N_4665,N_3052,N_3528);
or U4666 (N_4666,N_3251,N_3359);
or U4667 (N_4667,N_2881,N_3021);
and U4668 (N_4668,N_3420,N_3094);
nand U4669 (N_4669,N_2964,N_2555);
or U4670 (N_4670,N_2624,N_3413);
xor U4671 (N_4671,N_2464,N_2836);
nand U4672 (N_4672,N_2728,N_3391);
nand U4673 (N_4673,N_2754,N_3049);
and U4674 (N_4674,N_3076,N_2933);
nor U4675 (N_4675,N_2552,N_3409);
or U4676 (N_4676,N_3268,N_3440);
or U4677 (N_4677,N_3290,N_2583);
nand U4678 (N_4678,N_2488,N_3558);
and U4679 (N_4679,N_3092,N_3473);
and U4680 (N_4680,N_3024,N_3466);
or U4681 (N_4681,N_2932,N_3568);
nor U4682 (N_4682,N_3548,N_2569);
or U4683 (N_4683,N_2420,N_2474);
xor U4684 (N_4684,N_3385,N_3353);
or U4685 (N_4685,N_3375,N_3516);
nand U4686 (N_4686,N_2860,N_2973);
xnor U4687 (N_4687,N_3528,N_2464);
and U4688 (N_4688,N_2788,N_2898);
and U4689 (N_4689,N_3150,N_2858);
nand U4690 (N_4690,N_2716,N_3419);
nand U4691 (N_4691,N_2536,N_3377);
and U4692 (N_4692,N_2553,N_3272);
xnor U4693 (N_4693,N_2604,N_3031);
nand U4694 (N_4694,N_3459,N_3386);
and U4695 (N_4695,N_2527,N_2842);
nand U4696 (N_4696,N_2532,N_3373);
xor U4697 (N_4697,N_2524,N_2792);
or U4698 (N_4698,N_2974,N_2890);
nor U4699 (N_4699,N_2614,N_3328);
nand U4700 (N_4700,N_2443,N_2411);
or U4701 (N_4701,N_3421,N_3068);
nor U4702 (N_4702,N_3027,N_3482);
or U4703 (N_4703,N_3541,N_3559);
xor U4704 (N_4704,N_2605,N_2486);
nor U4705 (N_4705,N_3269,N_3172);
nand U4706 (N_4706,N_3055,N_2442);
xor U4707 (N_4707,N_2553,N_2825);
or U4708 (N_4708,N_2659,N_2444);
and U4709 (N_4709,N_2609,N_3100);
nor U4710 (N_4710,N_3344,N_3590);
and U4711 (N_4711,N_3125,N_2420);
or U4712 (N_4712,N_2427,N_3260);
or U4713 (N_4713,N_2579,N_2811);
and U4714 (N_4714,N_3006,N_3483);
xor U4715 (N_4715,N_2815,N_2645);
nor U4716 (N_4716,N_2605,N_2624);
and U4717 (N_4717,N_3413,N_3500);
nand U4718 (N_4718,N_2845,N_2783);
xor U4719 (N_4719,N_2419,N_2810);
nor U4720 (N_4720,N_2443,N_3193);
and U4721 (N_4721,N_3158,N_3422);
and U4722 (N_4722,N_3051,N_2876);
xnor U4723 (N_4723,N_2552,N_3497);
or U4724 (N_4724,N_3121,N_3162);
or U4725 (N_4725,N_2905,N_3163);
xor U4726 (N_4726,N_2752,N_2575);
nand U4727 (N_4727,N_2698,N_3440);
or U4728 (N_4728,N_2711,N_2656);
nand U4729 (N_4729,N_3485,N_2628);
nor U4730 (N_4730,N_3562,N_2503);
xor U4731 (N_4731,N_2450,N_2940);
or U4732 (N_4732,N_3074,N_3269);
or U4733 (N_4733,N_3000,N_3410);
and U4734 (N_4734,N_2550,N_2586);
or U4735 (N_4735,N_3232,N_2465);
and U4736 (N_4736,N_3274,N_2436);
nand U4737 (N_4737,N_2884,N_3434);
and U4738 (N_4738,N_2959,N_2649);
and U4739 (N_4739,N_3401,N_3502);
and U4740 (N_4740,N_3102,N_2796);
and U4741 (N_4741,N_2929,N_2651);
or U4742 (N_4742,N_2824,N_2459);
and U4743 (N_4743,N_3008,N_3139);
nor U4744 (N_4744,N_3192,N_3555);
or U4745 (N_4745,N_3143,N_3265);
or U4746 (N_4746,N_2940,N_3356);
or U4747 (N_4747,N_3176,N_3270);
nor U4748 (N_4748,N_3099,N_3389);
nor U4749 (N_4749,N_2582,N_2797);
nor U4750 (N_4750,N_3231,N_2792);
nand U4751 (N_4751,N_2639,N_2899);
and U4752 (N_4752,N_3495,N_3228);
and U4753 (N_4753,N_2448,N_3085);
xor U4754 (N_4754,N_3352,N_2721);
nor U4755 (N_4755,N_3303,N_2752);
nand U4756 (N_4756,N_3423,N_3580);
xor U4757 (N_4757,N_2851,N_2577);
and U4758 (N_4758,N_2706,N_2433);
or U4759 (N_4759,N_3159,N_3273);
nand U4760 (N_4760,N_3590,N_3066);
or U4761 (N_4761,N_2440,N_3133);
xor U4762 (N_4762,N_3453,N_3381);
nor U4763 (N_4763,N_3060,N_3284);
nand U4764 (N_4764,N_2409,N_2800);
and U4765 (N_4765,N_3347,N_2441);
xor U4766 (N_4766,N_2604,N_3294);
and U4767 (N_4767,N_3035,N_2428);
xnor U4768 (N_4768,N_2635,N_2658);
nand U4769 (N_4769,N_2751,N_2566);
xor U4770 (N_4770,N_3030,N_2461);
or U4771 (N_4771,N_2820,N_2490);
nand U4772 (N_4772,N_2703,N_3289);
and U4773 (N_4773,N_3105,N_2622);
nor U4774 (N_4774,N_3083,N_2631);
xnor U4775 (N_4775,N_2646,N_2589);
xor U4776 (N_4776,N_3556,N_2633);
xor U4777 (N_4777,N_3532,N_2987);
or U4778 (N_4778,N_3535,N_3070);
nand U4779 (N_4779,N_3524,N_2980);
nor U4780 (N_4780,N_3586,N_3340);
nand U4781 (N_4781,N_2922,N_3547);
nor U4782 (N_4782,N_2865,N_3162);
and U4783 (N_4783,N_3224,N_2542);
nand U4784 (N_4784,N_2886,N_3531);
nand U4785 (N_4785,N_3502,N_2792);
xnor U4786 (N_4786,N_2978,N_2726);
and U4787 (N_4787,N_3194,N_2800);
nand U4788 (N_4788,N_3034,N_2490);
or U4789 (N_4789,N_2999,N_3265);
or U4790 (N_4790,N_3525,N_3519);
and U4791 (N_4791,N_2658,N_2517);
nand U4792 (N_4792,N_3290,N_2578);
nand U4793 (N_4793,N_3509,N_3494);
nor U4794 (N_4794,N_2968,N_3475);
nand U4795 (N_4795,N_2860,N_2534);
xor U4796 (N_4796,N_2519,N_2403);
or U4797 (N_4797,N_3279,N_3177);
xor U4798 (N_4798,N_2710,N_3433);
xnor U4799 (N_4799,N_3308,N_2920);
or U4800 (N_4800,N_4706,N_4143);
nand U4801 (N_4801,N_3888,N_3683);
xnor U4802 (N_4802,N_4236,N_3899);
nand U4803 (N_4803,N_3853,N_4131);
xnor U4804 (N_4804,N_3749,N_4391);
nand U4805 (N_4805,N_3696,N_4051);
nor U4806 (N_4806,N_4402,N_4770);
xnor U4807 (N_4807,N_4323,N_4485);
nor U4808 (N_4808,N_4258,N_3827);
and U4809 (N_4809,N_3699,N_4431);
or U4810 (N_4810,N_3919,N_4118);
and U4811 (N_4811,N_4022,N_3859);
nor U4812 (N_4812,N_4496,N_4309);
nor U4813 (N_4813,N_3755,N_4082);
or U4814 (N_4814,N_4384,N_4318);
nand U4815 (N_4815,N_4441,N_4169);
or U4816 (N_4816,N_3608,N_4013);
and U4817 (N_4817,N_4634,N_4540);
or U4818 (N_4818,N_4733,N_4599);
nor U4819 (N_4819,N_3780,N_4716);
nand U4820 (N_4820,N_4667,N_4685);
nor U4821 (N_4821,N_4604,N_4561);
xnor U4822 (N_4822,N_3718,N_4306);
or U4823 (N_4823,N_4030,N_3657);
and U4824 (N_4824,N_4150,N_3975);
nor U4825 (N_4825,N_4272,N_4301);
and U4826 (N_4826,N_4074,N_4750);
and U4827 (N_4827,N_4524,N_3843);
or U4828 (N_4828,N_3627,N_4167);
nor U4829 (N_4829,N_4268,N_4397);
xor U4830 (N_4830,N_4584,N_4459);
xnor U4831 (N_4831,N_3961,N_4601);
nor U4832 (N_4832,N_3765,N_4193);
or U4833 (N_4833,N_4758,N_4152);
nand U4834 (N_4834,N_3973,N_3686);
and U4835 (N_4835,N_4092,N_3828);
nand U4836 (N_4836,N_4280,N_4279);
or U4837 (N_4837,N_4113,N_3785);
and U4838 (N_4838,N_4620,N_3882);
and U4839 (N_4839,N_4385,N_4104);
xnor U4840 (N_4840,N_3790,N_4029);
nand U4841 (N_4841,N_3792,N_4626);
xor U4842 (N_4842,N_4573,N_3869);
nor U4843 (N_4843,N_4180,N_3668);
xor U4844 (N_4844,N_4375,N_4224);
nand U4845 (N_4845,N_3670,N_3730);
nand U4846 (N_4846,N_4125,N_3639);
nand U4847 (N_4847,N_3705,N_3922);
xnor U4848 (N_4848,N_4221,N_3737);
nor U4849 (N_4849,N_4010,N_4738);
xor U4850 (N_4850,N_4068,N_4484);
nand U4851 (N_4851,N_4035,N_4126);
nor U4852 (N_4852,N_3773,N_4265);
nand U4853 (N_4853,N_4712,N_4646);
and U4854 (N_4854,N_4614,N_3753);
and U4855 (N_4855,N_4465,N_4781);
and U4856 (N_4856,N_3767,N_4392);
or U4857 (N_4857,N_4471,N_4290);
nor U4858 (N_4858,N_4046,N_3962);
xnor U4859 (N_4859,N_4040,N_3816);
xor U4860 (N_4860,N_4166,N_4789);
nor U4861 (N_4861,N_4711,N_4110);
nand U4862 (N_4862,N_4671,N_4625);
and U4863 (N_4863,N_3815,N_4579);
xnor U4864 (N_4864,N_4755,N_4346);
nand U4865 (N_4865,N_4648,N_4090);
nor U4866 (N_4866,N_4203,N_3929);
or U4867 (N_4867,N_3793,N_4562);
and U4868 (N_4868,N_4731,N_4592);
nor U4869 (N_4869,N_4565,N_4713);
xor U4870 (N_4870,N_4421,N_4552);
nand U4871 (N_4871,N_4136,N_3864);
nor U4872 (N_4872,N_3720,N_3889);
nand U4873 (N_4873,N_4657,N_3948);
and U4874 (N_4874,N_3867,N_4762);
or U4875 (N_4875,N_3750,N_3873);
nor U4876 (N_4876,N_4264,N_4518);
nand U4877 (N_4877,N_4137,N_4525);
nand U4878 (N_4878,N_4386,N_4133);
nor U4879 (N_4879,N_4448,N_4075);
and U4880 (N_4880,N_4768,N_3930);
and U4881 (N_4881,N_4393,N_3703);
or U4882 (N_4882,N_4239,N_3745);
and U4883 (N_4883,N_4588,N_4432);
nor U4884 (N_4884,N_4747,N_3808);
nor U4885 (N_4885,N_4057,N_4653);
nand U4886 (N_4886,N_4778,N_3974);
nand U4887 (N_4887,N_4248,N_3671);
nor U4888 (N_4888,N_4242,N_3878);
nor U4889 (N_4889,N_3817,N_4662);
and U4890 (N_4890,N_3908,N_4553);
nand U4891 (N_4891,N_4455,N_4718);
or U4892 (N_4892,N_4590,N_4005);
or U4893 (N_4893,N_4099,N_3661);
and U4894 (N_4894,N_4313,N_4497);
nand U4895 (N_4895,N_3868,N_4660);
nand U4896 (N_4896,N_4335,N_4668);
nor U4897 (N_4897,N_3850,N_3890);
and U4898 (N_4898,N_3998,N_4149);
nand U4899 (N_4899,N_4535,N_4440);
xnor U4900 (N_4900,N_4021,N_3698);
nand U4901 (N_4901,N_3824,N_3652);
xnor U4902 (N_4902,N_3723,N_4098);
nor U4903 (N_4903,N_3732,N_3846);
and U4904 (N_4904,N_3988,N_4558);
nor U4905 (N_4905,N_4454,N_4189);
nand U4906 (N_4906,N_4516,N_4447);
nor U4907 (N_4907,N_4434,N_4340);
nor U4908 (N_4908,N_3777,N_4076);
nand U4909 (N_4909,N_3641,N_3976);
and U4910 (N_4910,N_4526,N_4492);
nor U4911 (N_4911,N_3746,N_3787);
xnor U4912 (N_4912,N_4539,N_4387);
xor U4913 (N_4913,N_3937,N_4453);
or U4914 (N_4914,N_3701,N_3783);
xnor U4915 (N_4915,N_3757,N_3968);
or U4916 (N_4916,N_4311,N_4019);
or U4917 (N_4917,N_4720,N_3965);
or U4918 (N_4918,N_3942,N_4106);
and U4919 (N_4919,N_3761,N_3616);
nand U4920 (N_4920,N_4055,N_3642);
and U4921 (N_4921,N_3996,N_4709);
and U4922 (N_4922,N_3969,N_4664);
nand U4923 (N_4923,N_4025,N_4223);
nand U4924 (N_4924,N_4594,N_4237);
and U4925 (N_4925,N_4372,N_4756);
xor U4926 (N_4926,N_4480,N_4319);
xnor U4927 (N_4927,N_4532,N_4370);
nand U4928 (N_4928,N_3911,N_4343);
or U4929 (N_4929,N_4038,N_4546);
xnor U4930 (N_4930,N_4690,N_4211);
nor U4931 (N_4931,N_4663,N_3833);
nand U4932 (N_4932,N_4234,N_4452);
or U4933 (N_4933,N_4586,N_4139);
xnor U4934 (N_4934,N_4080,N_3883);
and U4935 (N_4935,N_3904,N_3759);
nand U4936 (N_4936,N_3631,N_4537);
nand U4937 (N_4937,N_4328,N_4503);
and U4938 (N_4938,N_4761,N_4643);
and U4939 (N_4939,N_3622,N_4276);
and U4940 (N_4940,N_4534,N_4305);
or U4941 (N_4941,N_4517,N_4398);
nand U4942 (N_4942,N_4331,N_4570);
nor U4943 (N_4943,N_4753,N_4209);
xnor U4944 (N_4944,N_4141,N_4155);
and U4945 (N_4945,N_4593,N_4316);
or U4946 (N_4946,N_4487,N_4184);
and U4947 (N_4947,N_4160,N_4514);
xnor U4948 (N_4948,N_4597,N_4219);
nor U4949 (N_4949,N_4702,N_4363);
nor U4950 (N_4950,N_3966,N_4610);
nor U4951 (N_4951,N_4495,N_4191);
or U4952 (N_4952,N_4270,N_3636);
and U4953 (N_4953,N_4481,N_3805);
nor U4954 (N_4954,N_4457,N_4719);
and U4955 (N_4955,N_3741,N_3902);
nand U4956 (N_4956,N_3635,N_4108);
and U4957 (N_4957,N_3721,N_4689);
or U4958 (N_4958,N_4122,N_4489);
nor U4959 (N_4959,N_3964,N_3949);
or U4960 (N_4960,N_4053,N_4119);
or U4961 (N_4961,N_4228,N_4470);
or U4962 (N_4962,N_3821,N_4024);
or U4963 (N_4963,N_3852,N_4230);
xnor U4964 (N_4964,N_4674,N_4249);
nand U4965 (N_4965,N_3934,N_4679);
xnor U4966 (N_4966,N_3989,N_3624);
or U4967 (N_4967,N_4142,N_4416);
xor U4968 (N_4968,N_3943,N_4278);
and U4969 (N_4969,N_3865,N_4582);
or U4970 (N_4970,N_3754,N_4430);
nor U4971 (N_4971,N_4530,N_3825);
and U4972 (N_4972,N_3945,N_4446);
or U4973 (N_4973,N_4473,N_3611);
xor U4974 (N_4974,N_4369,N_4501);
xnor U4975 (N_4975,N_4255,N_4275);
nand U4976 (N_4976,N_3630,N_4563);
and U4977 (N_4977,N_4476,N_3664);
or U4978 (N_4978,N_4418,N_4377);
and U4979 (N_4979,N_3604,N_3665);
nand U4980 (N_4980,N_4292,N_4608);
and U4981 (N_4981,N_4066,N_3912);
or U4982 (N_4982,N_3806,N_3713);
xor U4983 (N_4983,N_4672,N_4031);
nand U4984 (N_4984,N_3885,N_4782);
xnor U4985 (N_4985,N_4569,N_4611);
and U4986 (N_4986,N_3690,N_3687);
nand U4987 (N_4987,N_3724,N_4609);
and U4988 (N_4988,N_3860,N_4656);
xnor U4989 (N_4989,N_3650,N_3640);
xor U4990 (N_4990,N_4566,N_4645);
xor U4991 (N_4991,N_4324,N_3870);
xnor U4992 (N_4992,N_4794,N_3752);
xor U4993 (N_4993,N_4329,N_4683);
or U4994 (N_4994,N_3798,N_4721);
or U4995 (N_4995,N_3857,N_4124);
xor U4996 (N_4996,N_4135,N_3736);
and U4997 (N_4997,N_3907,N_4214);
xnor U4998 (N_4998,N_4355,N_3967);
nor U4999 (N_4999,N_4103,N_4414);
nor U5000 (N_5000,N_3840,N_4380);
or U5001 (N_5001,N_3638,N_4572);
nand U5002 (N_5002,N_4680,N_4542);
xor U5003 (N_5003,N_3880,N_4776);
nor U5004 (N_5004,N_4458,N_4638);
nor U5005 (N_5005,N_3841,N_4262);
nand U5006 (N_5006,N_3995,N_4735);
or U5007 (N_5007,N_3771,N_3971);
xor U5008 (N_5008,N_3905,N_4771);
and U5009 (N_5009,N_3603,N_4274);
nand U5010 (N_5010,N_4208,N_4033);
nor U5011 (N_5011,N_4088,N_4682);
xor U5012 (N_5012,N_4741,N_3855);
nand U5013 (N_5013,N_3960,N_4337);
xnor U5014 (N_5014,N_3688,N_4576);
xnor U5015 (N_5015,N_4308,N_3692);
xnor U5016 (N_5016,N_4232,N_4161);
xnor U5017 (N_5017,N_4206,N_3914);
and U5018 (N_5018,N_3726,N_4006);
xor U5019 (N_5019,N_4783,N_4354);
or U5020 (N_5020,N_4358,N_4326);
nand U5021 (N_5021,N_3795,N_4395);
and U5022 (N_5022,N_4288,N_3913);
xnor U5023 (N_5023,N_3784,N_4538);
nand U5024 (N_5024,N_3715,N_4202);
nand U5025 (N_5025,N_4406,N_3836);
and U5026 (N_5026,N_4687,N_4240);
and U5027 (N_5027,N_4763,N_3881);
nand U5028 (N_5028,N_4298,N_4460);
xnor U5029 (N_5029,N_3766,N_3666);
nor U5030 (N_5030,N_4708,N_4294);
or U5031 (N_5031,N_3660,N_3756);
nor U5032 (N_5032,N_4500,N_4423);
nor U5033 (N_5033,N_4543,N_4574);
and U5034 (N_5034,N_4407,N_3981);
xnor U5035 (N_5035,N_3619,N_4533);
xnor U5036 (N_5036,N_4351,N_3844);
xnor U5037 (N_5037,N_4474,N_4304);
nand U5038 (N_5038,N_4449,N_4164);
nand U5039 (N_5039,N_4284,N_3993);
xor U5040 (N_5040,N_3662,N_3955);
and U5041 (N_5041,N_3658,N_4580);
nor U5042 (N_5042,N_4462,N_4725);
xnor U5043 (N_5043,N_3957,N_4757);
and U5044 (N_5044,N_3609,N_4047);
nand U5045 (N_5045,N_3801,N_4394);
nand U5046 (N_5046,N_4784,N_4371);
nor U5047 (N_5047,N_3891,N_3782);
nor U5048 (N_5048,N_4165,N_4256);
and U5049 (N_5049,N_3941,N_3606);
or U5050 (N_5050,N_4201,N_4606);
xnor U5051 (N_5051,N_3977,N_4127);
or U5052 (N_5052,N_4178,N_4691);
and U5053 (N_5053,N_4085,N_3927);
nor U5054 (N_5054,N_4128,N_4595);
or U5055 (N_5055,N_4365,N_4396);
or U5056 (N_5056,N_3959,N_3926);
and U5057 (N_5057,N_4041,N_3681);
or U5058 (N_5058,N_4271,N_4486);
xor U5059 (N_5059,N_3663,N_3747);
and U5060 (N_5060,N_4204,N_3731);
nand U5061 (N_5061,N_4154,N_4764);
xor U5062 (N_5062,N_4095,N_3739);
and U5063 (N_5063,N_3951,N_4225);
nor U5064 (N_5064,N_4056,N_3924);
xor U5065 (N_5065,N_4008,N_3980);
xor U5066 (N_5066,N_4176,N_4675);
or U5067 (N_5067,N_4623,N_4069);
xnor U5068 (N_5068,N_3762,N_4244);
or U5069 (N_5069,N_4527,N_4296);
nand U5070 (N_5070,N_4723,N_4109);
or U5071 (N_5071,N_4303,N_4145);
nand U5072 (N_5072,N_4320,N_4064);
nand U5073 (N_5073,N_4216,N_4312);
xor U5074 (N_5074,N_4378,N_4138);
and U5075 (N_5075,N_3637,N_4529);
nand U5076 (N_5076,N_3990,N_4357);
xnor U5077 (N_5077,N_3875,N_4531);
xor U5078 (N_5078,N_3618,N_3615);
or U5079 (N_5079,N_4661,N_4374);
nor U5080 (N_5080,N_4267,N_4630);
nand U5081 (N_5081,N_4699,N_4456);
and U5082 (N_5082,N_3823,N_4425);
nand U5083 (N_5083,N_4600,N_4156);
or U5084 (N_5084,N_4436,N_4192);
and U5085 (N_5085,N_4468,N_4724);
xor U5086 (N_5086,N_3653,N_4696);
and U5087 (N_5087,N_3778,N_4445);
and U5088 (N_5088,N_3605,N_4307);
and U5089 (N_5089,N_3693,N_4635);
or U5090 (N_5090,N_4213,N_4334);
nand U5091 (N_5091,N_3886,N_4737);
nor U5092 (N_5092,N_4246,N_4442);
nand U5093 (N_5093,N_4793,N_4121);
xnor U5094 (N_5094,N_4642,N_4508);
or U5095 (N_5095,N_4097,N_3751);
nor U5096 (N_5096,N_4359,N_3839);
and U5097 (N_5097,N_3710,N_4297);
nand U5098 (N_5098,N_3626,N_4100);
nand U5099 (N_5099,N_3917,N_4190);
and U5100 (N_5100,N_4676,N_4637);
xor U5101 (N_5101,N_3614,N_3818);
nand U5102 (N_5102,N_3940,N_4158);
nor U5103 (N_5103,N_3684,N_4507);
xnor U5104 (N_5104,N_4017,N_4797);
nand U5105 (N_5105,N_3896,N_4235);
xor U5106 (N_5106,N_4171,N_3620);
nor U5107 (N_5107,N_3717,N_4791);
and U5108 (N_5108,N_4144,N_4252);
nand U5109 (N_5109,N_3901,N_3772);
and U5110 (N_5110,N_4727,N_3769);
nor U5111 (N_5111,N_4515,N_3863);
nor U5112 (N_5112,N_4159,N_3768);
xnor U5113 (N_5113,N_4077,N_4697);
and U5114 (N_5114,N_4198,N_3809);
xor U5115 (N_5115,N_4506,N_4027);
nand U5116 (N_5116,N_4379,N_4622);
and U5117 (N_5117,N_4020,N_4767);
nand U5118 (N_5118,N_4603,N_3939);
nor U5119 (N_5119,N_4651,N_4598);
and U5120 (N_5120,N_4116,N_4577);
nor U5121 (N_5121,N_3845,N_4678);
nand U5122 (N_5122,N_4405,N_3725);
or U5123 (N_5123,N_4799,N_3842);
and U5124 (N_5124,N_4388,N_3789);
or U5125 (N_5125,N_4695,N_4205);
and U5126 (N_5126,N_4123,N_3689);
or U5127 (N_5127,N_4752,N_4479);
or U5128 (N_5128,N_4681,N_4117);
nand U5129 (N_5129,N_4686,N_4222);
or U5130 (N_5130,N_4581,N_4281);
nand U5131 (N_5131,N_3879,N_3800);
xnor U5132 (N_5132,N_4728,N_4439);
or U5133 (N_5133,N_3675,N_3849);
or U5134 (N_5134,N_4684,N_3740);
or U5135 (N_5135,N_4015,N_4605);
xor U5136 (N_5136,N_3695,N_4583);
or U5137 (N_5137,N_4490,N_4000);
xor U5138 (N_5138,N_4383,N_4641);
nand U5139 (N_5139,N_4036,N_3837);
nor U5140 (N_5140,N_3925,N_4437);
xor U5141 (N_5141,N_3970,N_4701);
nand U5142 (N_5142,N_4382,N_4785);
nand U5143 (N_5143,N_4499,N_3621);
nor U5144 (N_5144,N_4060,N_4322);
nand U5145 (N_5145,N_3685,N_4536);
xor U5146 (N_5146,N_3794,N_3947);
or U5147 (N_5147,N_4049,N_3994);
nand U5148 (N_5148,N_3956,N_4283);
or U5149 (N_5149,N_4617,N_4067);
nor U5150 (N_5150,N_4618,N_4101);
or U5151 (N_5151,N_4408,N_4426);
and U5152 (N_5152,N_4774,N_3654);
nand U5153 (N_5153,N_4420,N_3810);
nand U5154 (N_5154,N_4512,N_3972);
and U5155 (N_5155,N_4707,N_3735);
nand U5156 (N_5156,N_4004,N_3952);
or U5157 (N_5157,N_4792,N_4636);
xor U5158 (N_5158,N_3678,N_3682);
xnor U5159 (N_5159,N_4177,N_4482);
nor U5160 (N_5160,N_4415,N_4710);
nor U5161 (N_5161,N_3733,N_4148);
or U5162 (N_5162,N_4287,N_4293);
xor U5163 (N_5163,N_4245,N_3851);
or U5164 (N_5164,N_3822,N_4559);
nand U5165 (N_5165,N_4591,N_4528);
nor U5166 (N_5166,N_4016,N_3950);
xnor U5167 (N_5167,N_4666,N_4732);
and U5168 (N_5168,N_4520,N_4647);
xor U5169 (N_5169,N_4018,N_3655);
nor U5170 (N_5170,N_4743,N_4568);
nand U5171 (N_5171,N_4417,N_4014);
xnor U5172 (N_5172,N_4295,N_3763);
nand U5173 (N_5173,N_4772,N_4780);
nor U5174 (N_5174,N_4325,N_4475);
nand U5175 (N_5175,N_3708,N_4194);
nor U5176 (N_5176,N_4607,N_3674);
nand U5177 (N_5177,N_4717,N_4009);
or U5178 (N_5178,N_4350,N_4612);
xor U5179 (N_5179,N_3673,N_3838);
and U5180 (N_5180,N_3744,N_3656);
nor U5181 (N_5181,N_4112,N_4332);
or U5182 (N_5182,N_4111,N_3986);
nand U5183 (N_5183,N_4070,N_4129);
xor U5184 (N_5184,N_4333,N_4032);
or U5185 (N_5185,N_3804,N_4409);
nor U5186 (N_5186,N_4341,N_4649);
xor U5187 (N_5187,N_3877,N_4045);
xnor U5188 (N_5188,N_4162,N_4754);
nor U5189 (N_5189,N_4362,N_3711);
xor U5190 (N_5190,N_4745,N_3812);
and U5191 (N_5191,N_3649,N_4629);
nand U5192 (N_5192,N_4314,N_4050);
or U5193 (N_5193,N_4188,N_4083);
xor U5194 (N_5194,N_3788,N_4483);
xor U5195 (N_5195,N_4548,N_4217);
or U5196 (N_5196,N_3920,N_4419);
nand U5197 (N_5197,N_3909,N_3617);
xor U5198 (N_5198,N_4179,N_4115);
nand U5199 (N_5199,N_3832,N_3694);
nor U5200 (N_5200,N_3643,N_4744);
xor U5201 (N_5201,N_4114,N_4187);
nand U5202 (N_5202,N_4786,N_4510);
xor U5203 (N_5203,N_3979,N_4412);
or U5204 (N_5204,N_4102,N_4659);
and U5205 (N_5205,N_4063,N_3985);
or U5206 (N_5206,N_4344,N_3647);
nor U5207 (N_5207,N_3835,N_4389);
nand U5208 (N_5208,N_4748,N_3910);
or U5209 (N_5209,N_4410,N_3781);
or U5210 (N_5210,N_4795,N_4310);
nand U5211 (N_5211,N_4700,N_4093);
xor U5212 (N_5212,N_3704,N_4621);
nor U5213 (N_5213,N_4196,N_4183);
nand U5214 (N_5214,N_4511,N_4215);
and U5215 (N_5215,N_4413,N_4360);
nand U5216 (N_5216,N_4153,N_4229);
nand U5217 (N_5217,N_3774,N_3872);
nand U5218 (N_5218,N_4749,N_4551);
or U5219 (N_5219,N_4729,N_4522);
xnor U5220 (N_5220,N_4073,N_4130);
and U5221 (N_5221,N_3677,N_3814);
nand U5222 (N_5222,N_4347,N_3680);
nor U5223 (N_5223,N_4567,N_4627);
nor U5224 (N_5224,N_4173,N_4502);
or U5225 (N_5225,N_4317,N_3978);
and U5226 (N_5226,N_4348,N_3871);
xnor U5227 (N_5227,N_3729,N_4266);
nor U5228 (N_5228,N_3770,N_4596);
nor U5229 (N_5229,N_4012,N_4564);
and U5230 (N_5230,N_4488,N_4059);
nand U5231 (N_5231,N_3811,N_4521);
nor U5232 (N_5232,N_4698,N_3628);
and U5233 (N_5233,N_4401,N_3983);
nand U5234 (N_5234,N_4058,N_3779);
and U5235 (N_5235,N_4644,N_3602);
nand U5236 (N_5236,N_3894,N_3932);
and U5237 (N_5237,N_4556,N_3764);
and U5238 (N_5238,N_4472,N_4422);
nand U5239 (N_5239,N_4003,N_4739);
nand U5240 (N_5240,N_3936,N_4545);
or U5241 (N_5241,N_4790,N_4231);
nand U5242 (N_5242,N_3676,N_4054);
or U5243 (N_5243,N_4619,N_4218);
xor U5244 (N_5244,N_4151,N_3672);
xor U5245 (N_5245,N_3820,N_4321);
or U5246 (N_5246,N_4091,N_3796);
xor U5247 (N_5247,N_4438,N_4544);
and U5248 (N_5248,N_3892,N_4477);
nor U5249 (N_5249,N_3776,N_4376);
and U5250 (N_5250,N_3797,N_4011);
nand U5251 (N_5251,N_4726,N_4238);
nand U5252 (N_5252,N_4742,N_4157);
nor U5253 (N_5253,N_4286,N_4775);
nor U5254 (N_5254,N_4094,N_4443);
or U5255 (N_5255,N_3707,N_4463);
nand U5256 (N_5256,N_4260,N_4736);
nand U5257 (N_5257,N_4693,N_4107);
nand U5258 (N_5258,N_3897,N_3858);
nor U5259 (N_5259,N_4704,N_4769);
or U5260 (N_5260,N_4105,N_4478);
nand U5261 (N_5261,N_3997,N_4613);
nor U5262 (N_5262,N_4199,N_4163);
xnor U5263 (N_5263,N_3760,N_3610);
nand U5264 (N_5264,N_3900,N_4361);
or U5265 (N_5265,N_3876,N_4373);
nor U5266 (N_5266,N_4028,N_3791);
nor U5267 (N_5267,N_4336,N_3982);
xor U5268 (N_5268,N_4220,N_4247);
and U5269 (N_5269,N_4773,N_4513);
and U5270 (N_5270,N_4044,N_3953);
nand U5271 (N_5271,N_4081,N_4428);
xnor U5272 (N_5272,N_4364,N_3963);
xnor U5273 (N_5273,N_4182,N_4034);
xnor U5274 (N_5274,N_4450,N_3923);
xnor U5275 (N_5275,N_4705,N_3775);
xnor U5276 (N_5276,N_4779,N_4547);
or U5277 (N_5277,N_3854,N_4146);
xor U5278 (N_5278,N_3629,N_3758);
or U5279 (N_5279,N_3743,N_4259);
and U5280 (N_5280,N_3944,N_3691);
or U5281 (N_5281,N_4241,N_4504);
and U5282 (N_5282,N_4078,N_4043);
xor U5283 (N_5283,N_3916,N_4451);
xnor U5284 (N_5284,N_4291,N_4427);
nand U5285 (N_5285,N_4253,N_4692);
nor U5286 (N_5286,N_4652,N_4352);
and U5287 (N_5287,N_3634,N_3722);
nor U5288 (N_5288,N_3623,N_4381);
nor U5289 (N_5289,N_4195,N_3700);
xor U5290 (N_5290,N_4461,N_4147);
or U5291 (N_5291,N_4251,N_4519);
or U5292 (N_5292,N_4185,N_4086);
and U5293 (N_5293,N_4368,N_4665);
and U5294 (N_5294,N_4120,N_4403);
and U5295 (N_5295,N_4424,N_4655);
nor U5296 (N_5296,N_3632,N_4065);
nand U5297 (N_5297,N_4227,N_4134);
or U5298 (N_5298,N_4339,N_4345);
nand U5299 (N_5299,N_3697,N_4688);
nand U5300 (N_5300,N_4226,N_3893);
xor U5301 (N_5301,N_4039,N_4541);
and U5302 (N_5302,N_4494,N_4263);
nor U5303 (N_5303,N_3931,N_3915);
or U5304 (N_5304,N_4315,N_4498);
nor U5305 (N_5305,N_4285,N_3861);
and U5306 (N_5306,N_3874,N_3728);
and U5307 (N_5307,N_4677,N_4788);
nor U5308 (N_5308,N_3625,N_3935);
xor U5309 (N_5309,N_4289,N_3706);
and U5310 (N_5310,N_4585,N_4523);
and U5311 (N_5311,N_4273,N_4589);
or U5312 (N_5312,N_3709,N_4673);
nor U5313 (N_5313,N_3601,N_3847);
xnor U5314 (N_5314,N_3807,N_3786);
nand U5315 (N_5315,N_4175,N_4411);
and U5316 (N_5316,N_3648,N_4404);
nor U5317 (N_5317,N_4624,N_3799);
xor U5318 (N_5318,N_4026,N_3612);
xnor U5319 (N_5319,N_4639,N_3613);
and U5320 (N_5320,N_4299,N_4282);
or U5321 (N_5321,N_3830,N_4560);
xnor U5322 (N_5322,N_4250,N_3887);
and U5323 (N_5323,N_4342,N_4766);
xor U5324 (N_5324,N_4796,N_4089);
xor U5325 (N_5325,N_3742,N_3644);
and U5326 (N_5326,N_3895,N_4444);
nand U5327 (N_5327,N_4257,N_4658);
nor U5328 (N_5328,N_4730,N_4399);
xor U5329 (N_5329,N_4079,N_4042);
and U5330 (N_5330,N_4174,N_4670);
xnor U5331 (N_5331,N_3918,N_4277);
or U5332 (N_5332,N_3600,N_4466);
nor U5333 (N_5333,N_4367,N_4715);
and U5334 (N_5334,N_4181,N_4650);
xnor U5335 (N_5335,N_4703,N_4084);
xor U5336 (N_5336,N_4002,N_4615);
nor U5337 (N_5337,N_4760,N_3903);
and U5338 (N_5338,N_4338,N_4571);
xor U5339 (N_5339,N_4746,N_3702);
nand U5340 (N_5340,N_3714,N_3679);
nor U5341 (N_5341,N_4493,N_4096);
nand U5342 (N_5342,N_4554,N_4631);
or U5343 (N_5343,N_4212,N_4327);
and U5344 (N_5344,N_4654,N_4616);
and U5345 (N_5345,N_4429,N_3954);
and U5346 (N_5346,N_4798,N_3803);
nand U5347 (N_5347,N_4550,N_3958);
and U5348 (N_5348,N_3802,N_3884);
nor U5349 (N_5349,N_4669,N_3834);
nand U5350 (N_5350,N_4200,N_4602);
and U5351 (N_5351,N_4072,N_3813);
nand U5352 (N_5352,N_4210,N_3719);
nor U5353 (N_5353,N_4062,N_4491);
and U5354 (N_5354,N_4464,N_3999);
or U5355 (N_5355,N_3938,N_4435);
xnor U5356 (N_5356,N_3738,N_4694);
or U5357 (N_5357,N_3633,N_3991);
xor U5358 (N_5358,N_4140,N_4587);
nand U5359 (N_5359,N_4400,N_4037);
or U5360 (N_5360,N_4302,N_3856);
and U5361 (N_5361,N_4001,N_4557);
xor U5362 (N_5362,N_3646,N_3659);
and U5363 (N_5363,N_4640,N_4765);
and U5364 (N_5364,N_4632,N_4061);
and U5365 (N_5365,N_4555,N_4300);
nor U5366 (N_5366,N_3669,N_4170);
nor U5367 (N_5367,N_4087,N_4207);
nor U5368 (N_5368,N_4722,N_4172);
nand U5369 (N_5369,N_3727,N_4366);
xor U5370 (N_5370,N_3829,N_4007);
and U5371 (N_5371,N_3946,N_4048);
xnor U5372 (N_5372,N_3748,N_4353);
nor U5373 (N_5373,N_3645,N_4261);
and U5374 (N_5374,N_4740,N_4132);
nand U5375 (N_5375,N_3928,N_4186);
or U5376 (N_5376,N_3734,N_4349);
or U5377 (N_5377,N_4071,N_4390);
nand U5378 (N_5378,N_4243,N_3651);
xor U5379 (N_5379,N_3933,N_4549);
and U5380 (N_5380,N_4254,N_4633);
or U5381 (N_5381,N_4330,N_3898);
and U5382 (N_5382,N_4233,N_3819);
xnor U5383 (N_5383,N_4787,N_4052);
and U5384 (N_5384,N_4168,N_4578);
nor U5385 (N_5385,N_3866,N_4356);
nand U5386 (N_5386,N_3984,N_4269);
nand U5387 (N_5387,N_3607,N_4759);
and U5388 (N_5388,N_3831,N_4714);
or U5389 (N_5389,N_4433,N_4777);
xnor U5390 (N_5390,N_3862,N_3848);
nor U5391 (N_5391,N_3667,N_3826);
or U5392 (N_5392,N_4751,N_4469);
nand U5393 (N_5393,N_4505,N_4575);
and U5394 (N_5394,N_4734,N_3992);
xnor U5395 (N_5395,N_3906,N_3921);
nor U5396 (N_5396,N_4628,N_3987);
or U5397 (N_5397,N_4023,N_4467);
xor U5398 (N_5398,N_4509,N_4197);
or U5399 (N_5399,N_3712,N_3716);
xor U5400 (N_5400,N_4020,N_3922);
or U5401 (N_5401,N_4408,N_4107);
nand U5402 (N_5402,N_4126,N_3795);
or U5403 (N_5403,N_3900,N_4445);
or U5404 (N_5404,N_3615,N_4079);
and U5405 (N_5405,N_4165,N_3782);
nor U5406 (N_5406,N_4535,N_3909);
xnor U5407 (N_5407,N_4721,N_4163);
and U5408 (N_5408,N_4006,N_4200);
and U5409 (N_5409,N_4529,N_4248);
and U5410 (N_5410,N_3916,N_3996);
nand U5411 (N_5411,N_4394,N_3704);
nand U5412 (N_5412,N_4499,N_3917);
xnor U5413 (N_5413,N_4607,N_3865);
and U5414 (N_5414,N_3715,N_4479);
xnor U5415 (N_5415,N_3839,N_4109);
xor U5416 (N_5416,N_3612,N_4000);
nor U5417 (N_5417,N_4406,N_4020);
or U5418 (N_5418,N_4578,N_4245);
or U5419 (N_5419,N_4739,N_4683);
nand U5420 (N_5420,N_3752,N_3653);
or U5421 (N_5421,N_4016,N_4066);
or U5422 (N_5422,N_4581,N_4130);
nand U5423 (N_5423,N_4756,N_3884);
or U5424 (N_5424,N_4772,N_4678);
or U5425 (N_5425,N_4601,N_4471);
or U5426 (N_5426,N_3730,N_4783);
xor U5427 (N_5427,N_3910,N_4674);
and U5428 (N_5428,N_3647,N_4580);
nand U5429 (N_5429,N_4432,N_3750);
nor U5430 (N_5430,N_4485,N_4439);
or U5431 (N_5431,N_4058,N_4449);
or U5432 (N_5432,N_4386,N_4752);
and U5433 (N_5433,N_4041,N_3721);
and U5434 (N_5434,N_4004,N_4126);
xor U5435 (N_5435,N_4466,N_4241);
nor U5436 (N_5436,N_4241,N_4085);
or U5437 (N_5437,N_4698,N_3759);
and U5438 (N_5438,N_4204,N_4641);
or U5439 (N_5439,N_3676,N_4253);
or U5440 (N_5440,N_4787,N_4589);
xnor U5441 (N_5441,N_4719,N_4518);
nor U5442 (N_5442,N_4263,N_3694);
nor U5443 (N_5443,N_4611,N_4550);
xor U5444 (N_5444,N_4278,N_4166);
xnor U5445 (N_5445,N_4476,N_4651);
xnor U5446 (N_5446,N_4363,N_4490);
xor U5447 (N_5447,N_4393,N_4404);
nand U5448 (N_5448,N_4269,N_4010);
and U5449 (N_5449,N_4196,N_3874);
xnor U5450 (N_5450,N_4452,N_4329);
xnor U5451 (N_5451,N_3641,N_4728);
or U5452 (N_5452,N_4365,N_4437);
nor U5453 (N_5453,N_3857,N_4784);
nand U5454 (N_5454,N_4502,N_4686);
and U5455 (N_5455,N_4499,N_4321);
nand U5456 (N_5456,N_4707,N_4659);
or U5457 (N_5457,N_4035,N_4075);
and U5458 (N_5458,N_3674,N_4698);
xnor U5459 (N_5459,N_4095,N_4400);
nand U5460 (N_5460,N_3971,N_4269);
xnor U5461 (N_5461,N_4369,N_3821);
nand U5462 (N_5462,N_4746,N_4235);
or U5463 (N_5463,N_3827,N_3801);
nor U5464 (N_5464,N_3902,N_4347);
nand U5465 (N_5465,N_3665,N_4735);
or U5466 (N_5466,N_3736,N_4532);
nand U5467 (N_5467,N_3970,N_4051);
nor U5468 (N_5468,N_4071,N_4202);
and U5469 (N_5469,N_4318,N_4789);
nor U5470 (N_5470,N_3762,N_3905);
and U5471 (N_5471,N_3918,N_3828);
xnor U5472 (N_5472,N_3706,N_4261);
nor U5473 (N_5473,N_4524,N_3995);
and U5474 (N_5474,N_3685,N_4232);
nand U5475 (N_5475,N_3779,N_3686);
or U5476 (N_5476,N_3825,N_4192);
or U5477 (N_5477,N_3958,N_4505);
nor U5478 (N_5478,N_4023,N_4130);
xnor U5479 (N_5479,N_4791,N_3860);
xnor U5480 (N_5480,N_3938,N_4652);
and U5481 (N_5481,N_3756,N_4478);
nor U5482 (N_5482,N_4023,N_4190);
or U5483 (N_5483,N_4661,N_4729);
and U5484 (N_5484,N_4795,N_4778);
nand U5485 (N_5485,N_4586,N_4037);
xor U5486 (N_5486,N_3799,N_3997);
xor U5487 (N_5487,N_3752,N_4209);
or U5488 (N_5488,N_4168,N_4128);
xnor U5489 (N_5489,N_4615,N_3991);
nor U5490 (N_5490,N_4113,N_3841);
or U5491 (N_5491,N_4132,N_4379);
xor U5492 (N_5492,N_4787,N_4180);
nand U5493 (N_5493,N_3840,N_4493);
xor U5494 (N_5494,N_4511,N_3901);
and U5495 (N_5495,N_4310,N_3620);
nor U5496 (N_5496,N_4185,N_4174);
and U5497 (N_5497,N_3860,N_4067);
or U5498 (N_5498,N_4689,N_4125);
nand U5499 (N_5499,N_4467,N_3799);
xor U5500 (N_5500,N_4200,N_3716);
nand U5501 (N_5501,N_3639,N_4373);
xor U5502 (N_5502,N_3657,N_3844);
or U5503 (N_5503,N_4045,N_3871);
nor U5504 (N_5504,N_4229,N_4471);
xor U5505 (N_5505,N_4540,N_3922);
xnor U5506 (N_5506,N_4041,N_4541);
xor U5507 (N_5507,N_3661,N_4608);
nor U5508 (N_5508,N_4373,N_4736);
nor U5509 (N_5509,N_4334,N_4703);
and U5510 (N_5510,N_3823,N_4053);
nand U5511 (N_5511,N_4099,N_3651);
xnor U5512 (N_5512,N_4446,N_3683);
nor U5513 (N_5513,N_3623,N_4051);
xnor U5514 (N_5514,N_4760,N_4016);
xor U5515 (N_5515,N_4587,N_3632);
and U5516 (N_5516,N_4406,N_3963);
xnor U5517 (N_5517,N_3834,N_3979);
xnor U5518 (N_5518,N_4531,N_4066);
and U5519 (N_5519,N_4123,N_4224);
and U5520 (N_5520,N_4418,N_4287);
nand U5521 (N_5521,N_4297,N_4054);
or U5522 (N_5522,N_4568,N_4190);
and U5523 (N_5523,N_4239,N_3967);
nor U5524 (N_5524,N_4718,N_4341);
and U5525 (N_5525,N_4433,N_3972);
and U5526 (N_5526,N_4194,N_4145);
nand U5527 (N_5527,N_4016,N_4488);
xnor U5528 (N_5528,N_4382,N_3604);
xnor U5529 (N_5529,N_4654,N_3909);
nand U5530 (N_5530,N_3603,N_4719);
nor U5531 (N_5531,N_3839,N_4576);
nor U5532 (N_5532,N_4428,N_4450);
or U5533 (N_5533,N_4784,N_3678);
nor U5534 (N_5534,N_3667,N_3946);
nor U5535 (N_5535,N_4705,N_4303);
or U5536 (N_5536,N_4565,N_3970);
nor U5537 (N_5537,N_4768,N_4624);
xnor U5538 (N_5538,N_4737,N_4069);
nand U5539 (N_5539,N_4129,N_4187);
and U5540 (N_5540,N_3887,N_4793);
xor U5541 (N_5541,N_4777,N_4633);
nor U5542 (N_5542,N_4506,N_3642);
nand U5543 (N_5543,N_4753,N_4463);
xnor U5544 (N_5544,N_3764,N_4066);
nor U5545 (N_5545,N_4643,N_4595);
or U5546 (N_5546,N_3637,N_4314);
xor U5547 (N_5547,N_3963,N_3834);
xnor U5548 (N_5548,N_4495,N_4519);
nand U5549 (N_5549,N_3742,N_3717);
and U5550 (N_5550,N_3828,N_4406);
nor U5551 (N_5551,N_3724,N_4581);
and U5552 (N_5552,N_3864,N_3768);
nor U5553 (N_5553,N_3825,N_4273);
xor U5554 (N_5554,N_4311,N_3804);
xor U5555 (N_5555,N_4651,N_3885);
or U5556 (N_5556,N_3760,N_4639);
nand U5557 (N_5557,N_4309,N_4711);
and U5558 (N_5558,N_4746,N_3749);
nand U5559 (N_5559,N_4259,N_4229);
or U5560 (N_5560,N_4382,N_4305);
nor U5561 (N_5561,N_4386,N_4439);
xor U5562 (N_5562,N_3688,N_4720);
or U5563 (N_5563,N_4107,N_4177);
or U5564 (N_5564,N_3622,N_4015);
nand U5565 (N_5565,N_3988,N_4583);
nand U5566 (N_5566,N_4506,N_4014);
nor U5567 (N_5567,N_4322,N_3872);
xor U5568 (N_5568,N_4542,N_3746);
xor U5569 (N_5569,N_4422,N_4311);
or U5570 (N_5570,N_3900,N_3910);
and U5571 (N_5571,N_4498,N_4161);
xor U5572 (N_5572,N_4262,N_4779);
xnor U5573 (N_5573,N_4345,N_4288);
and U5574 (N_5574,N_3667,N_4131);
xor U5575 (N_5575,N_4622,N_3687);
nand U5576 (N_5576,N_4391,N_4515);
nor U5577 (N_5577,N_3658,N_3917);
xor U5578 (N_5578,N_4592,N_3931);
xor U5579 (N_5579,N_4075,N_4106);
or U5580 (N_5580,N_3683,N_3748);
and U5581 (N_5581,N_3619,N_4330);
and U5582 (N_5582,N_3657,N_3726);
or U5583 (N_5583,N_3961,N_3902);
and U5584 (N_5584,N_4100,N_4511);
nor U5585 (N_5585,N_4217,N_4235);
xnor U5586 (N_5586,N_4216,N_4157);
and U5587 (N_5587,N_4336,N_3807);
nor U5588 (N_5588,N_4453,N_4423);
and U5589 (N_5589,N_3896,N_4471);
nor U5590 (N_5590,N_4478,N_4243);
or U5591 (N_5591,N_4789,N_3618);
and U5592 (N_5592,N_4097,N_3746);
or U5593 (N_5593,N_4700,N_3651);
nand U5594 (N_5594,N_4197,N_4739);
or U5595 (N_5595,N_4053,N_4374);
or U5596 (N_5596,N_4041,N_3639);
nor U5597 (N_5597,N_4606,N_3972);
or U5598 (N_5598,N_4743,N_3601);
nand U5599 (N_5599,N_4009,N_3929);
or U5600 (N_5600,N_4432,N_4357);
nand U5601 (N_5601,N_4292,N_4319);
and U5602 (N_5602,N_3622,N_3908);
xor U5603 (N_5603,N_4088,N_3994);
nor U5604 (N_5604,N_4691,N_3635);
and U5605 (N_5605,N_4765,N_3954);
nor U5606 (N_5606,N_4078,N_4118);
nand U5607 (N_5607,N_4199,N_3750);
nor U5608 (N_5608,N_3915,N_4558);
nor U5609 (N_5609,N_4433,N_4151);
nor U5610 (N_5610,N_3677,N_4613);
nand U5611 (N_5611,N_3788,N_3754);
nand U5612 (N_5612,N_4405,N_4392);
nor U5613 (N_5613,N_4610,N_3681);
xnor U5614 (N_5614,N_4227,N_4116);
nor U5615 (N_5615,N_4705,N_3911);
nand U5616 (N_5616,N_3858,N_4688);
or U5617 (N_5617,N_3938,N_3939);
nand U5618 (N_5618,N_3625,N_4587);
xnor U5619 (N_5619,N_4188,N_4388);
and U5620 (N_5620,N_3992,N_4157);
xnor U5621 (N_5621,N_4176,N_3735);
nor U5622 (N_5622,N_4702,N_4340);
nor U5623 (N_5623,N_3650,N_3662);
and U5624 (N_5624,N_3833,N_3925);
nand U5625 (N_5625,N_3952,N_3873);
xnor U5626 (N_5626,N_4764,N_3885);
or U5627 (N_5627,N_3799,N_3830);
and U5628 (N_5628,N_4478,N_4163);
xnor U5629 (N_5629,N_4509,N_3906);
nor U5630 (N_5630,N_4008,N_4665);
xor U5631 (N_5631,N_3804,N_4623);
nor U5632 (N_5632,N_3646,N_4620);
and U5633 (N_5633,N_3810,N_4313);
nand U5634 (N_5634,N_3944,N_4681);
or U5635 (N_5635,N_4385,N_4241);
or U5636 (N_5636,N_4582,N_4040);
xor U5637 (N_5637,N_3600,N_3780);
xor U5638 (N_5638,N_3988,N_3717);
nand U5639 (N_5639,N_4251,N_3978);
nand U5640 (N_5640,N_4205,N_3957);
and U5641 (N_5641,N_4115,N_4474);
or U5642 (N_5642,N_4616,N_4773);
nand U5643 (N_5643,N_4694,N_4279);
and U5644 (N_5644,N_4240,N_4231);
and U5645 (N_5645,N_4169,N_4157);
xnor U5646 (N_5646,N_3629,N_3740);
nor U5647 (N_5647,N_3700,N_4518);
nor U5648 (N_5648,N_4204,N_3639);
or U5649 (N_5649,N_4521,N_4571);
nand U5650 (N_5650,N_4291,N_4724);
nand U5651 (N_5651,N_3856,N_3642);
or U5652 (N_5652,N_3759,N_3873);
xor U5653 (N_5653,N_4061,N_4747);
xor U5654 (N_5654,N_4283,N_4799);
xor U5655 (N_5655,N_4065,N_4145);
nor U5656 (N_5656,N_3778,N_4709);
nor U5657 (N_5657,N_4564,N_4721);
and U5658 (N_5658,N_4623,N_4177);
xor U5659 (N_5659,N_4516,N_4498);
xnor U5660 (N_5660,N_4316,N_4447);
and U5661 (N_5661,N_3970,N_3975);
xor U5662 (N_5662,N_4551,N_4601);
and U5663 (N_5663,N_3672,N_4049);
nor U5664 (N_5664,N_4148,N_4465);
or U5665 (N_5665,N_4703,N_4501);
or U5666 (N_5666,N_4176,N_4146);
xnor U5667 (N_5667,N_4361,N_4657);
and U5668 (N_5668,N_4371,N_3804);
and U5669 (N_5669,N_4167,N_4197);
or U5670 (N_5670,N_3651,N_3998);
nor U5671 (N_5671,N_4754,N_4545);
nand U5672 (N_5672,N_4746,N_4451);
nor U5673 (N_5673,N_4637,N_4653);
nor U5674 (N_5674,N_3641,N_3705);
nor U5675 (N_5675,N_3654,N_4241);
or U5676 (N_5676,N_4172,N_3862);
or U5677 (N_5677,N_3642,N_4320);
nor U5678 (N_5678,N_4653,N_4747);
and U5679 (N_5679,N_4394,N_4269);
or U5680 (N_5680,N_4423,N_4374);
and U5681 (N_5681,N_4209,N_3974);
or U5682 (N_5682,N_4264,N_3999);
or U5683 (N_5683,N_4196,N_4016);
and U5684 (N_5684,N_3727,N_4357);
nor U5685 (N_5685,N_4077,N_4184);
or U5686 (N_5686,N_4168,N_3896);
nand U5687 (N_5687,N_4691,N_4771);
xor U5688 (N_5688,N_4744,N_4336);
or U5689 (N_5689,N_4737,N_4156);
and U5690 (N_5690,N_4525,N_4501);
or U5691 (N_5691,N_4652,N_4026);
and U5692 (N_5692,N_4518,N_3892);
nor U5693 (N_5693,N_3921,N_4443);
xnor U5694 (N_5694,N_3997,N_3941);
and U5695 (N_5695,N_3755,N_4045);
xor U5696 (N_5696,N_4774,N_4739);
xor U5697 (N_5697,N_4063,N_3821);
xnor U5698 (N_5698,N_4122,N_4786);
xor U5699 (N_5699,N_3703,N_4124);
xor U5700 (N_5700,N_4342,N_4587);
or U5701 (N_5701,N_3910,N_4020);
nor U5702 (N_5702,N_4139,N_3787);
or U5703 (N_5703,N_4004,N_4275);
or U5704 (N_5704,N_3712,N_3727);
nand U5705 (N_5705,N_4235,N_3749);
and U5706 (N_5706,N_4402,N_4766);
or U5707 (N_5707,N_4645,N_4459);
nand U5708 (N_5708,N_4290,N_4243);
nand U5709 (N_5709,N_4118,N_3874);
and U5710 (N_5710,N_3929,N_4194);
or U5711 (N_5711,N_4239,N_4619);
and U5712 (N_5712,N_4389,N_4477);
nand U5713 (N_5713,N_4346,N_4710);
nand U5714 (N_5714,N_4629,N_3702);
nor U5715 (N_5715,N_4286,N_4549);
nand U5716 (N_5716,N_4281,N_4509);
xnor U5717 (N_5717,N_4150,N_4435);
nor U5718 (N_5718,N_4679,N_4534);
or U5719 (N_5719,N_4324,N_4103);
xnor U5720 (N_5720,N_4739,N_3904);
nor U5721 (N_5721,N_3797,N_4798);
and U5722 (N_5722,N_4447,N_4205);
nand U5723 (N_5723,N_3712,N_4455);
xor U5724 (N_5724,N_4262,N_4093);
xnor U5725 (N_5725,N_4797,N_3665);
nand U5726 (N_5726,N_3987,N_4338);
xor U5727 (N_5727,N_4714,N_4265);
and U5728 (N_5728,N_4127,N_4191);
and U5729 (N_5729,N_4005,N_4766);
nor U5730 (N_5730,N_4153,N_4532);
nor U5731 (N_5731,N_4737,N_4453);
nor U5732 (N_5732,N_4215,N_4008);
xor U5733 (N_5733,N_3754,N_4077);
nor U5734 (N_5734,N_4626,N_4357);
nor U5735 (N_5735,N_4259,N_4385);
nor U5736 (N_5736,N_4237,N_4684);
or U5737 (N_5737,N_3891,N_3616);
nor U5738 (N_5738,N_4626,N_4038);
nor U5739 (N_5739,N_4444,N_3617);
nand U5740 (N_5740,N_4248,N_4104);
and U5741 (N_5741,N_4419,N_4723);
nand U5742 (N_5742,N_4204,N_4485);
nor U5743 (N_5743,N_3695,N_4092);
and U5744 (N_5744,N_3622,N_4099);
xnor U5745 (N_5745,N_4277,N_3862);
or U5746 (N_5746,N_4260,N_4437);
nor U5747 (N_5747,N_4343,N_3889);
and U5748 (N_5748,N_4039,N_4278);
or U5749 (N_5749,N_4032,N_4518);
nand U5750 (N_5750,N_4729,N_3642);
or U5751 (N_5751,N_3662,N_4282);
xor U5752 (N_5752,N_4439,N_3683);
xor U5753 (N_5753,N_4359,N_4314);
xnor U5754 (N_5754,N_4563,N_4252);
xnor U5755 (N_5755,N_4644,N_3641);
xor U5756 (N_5756,N_3999,N_4215);
nand U5757 (N_5757,N_4281,N_4499);
nand U5758 (N_5758,N_3918,N_3891);
or U5759 (N_5759,N_4627,N_4144);
and U5760 (N_5760,N_4533,N_4398);
nand U5761 (N_5761,N_4050,N_3747);
and U5762 (N_5762,N_4485,N_3833);
nor U5763 (N_5763,N_4792,N_4274);
and U5764 (N_5764,N_4750,N_3855);
and U5765 (N_5765,N_3880,N_3896);
and U5766 (N_5766,N_3867,N_3689);
or U5767 (N_5767,N_4359,N_3613);
xnor U5768 (N_5768,N_4747,N_4518);
nor U5769 (N_5769,N_3864,N_4382);
nor U5770 (N_5770,N_4277,N_4414);
nor U5771 (N_5771,N_4688,N_4108);
nor U5772 (N_5772,N_3872,N_3780);
or U5773 (N_5773,N_3944,N_4744);
or U5774 (N_5774,N_4641,N_4407);
nor U5775 (N_5775,N_3872,N_3841);
and U5776 (N_5776,N_4095,N_4232);
nor U5777 (N_5777,N_4382,N_4622);
nand U5778 (N_5778,N_4650,N_4124);
xnor U5779 (N_5779,N_3838,N_4442);
or U5780 (N_5780,N_4680,N_4605);
xor U5781 (N_5781,N_4604,N_3986);
xnor U5782 (N_5782,N_4269,N_4609);
and U5783 (N_5783,N_3706,N_3816);
and U5784 (N_5784,N_4413,N_4268);
and U5785 (N_5785,N_3922,N_3666);
nand U5786 (N_5786,N_4458,N_3838);
or U5787 (N_5787,N_3946,N_4441);
xnor U5788 (N_5788,N_3621,N_4434);
nand U5789 (N_5789,N_4711,N_4290);
nor U5790 (N_5790,N_4472,N_3947);
xor U5791 (N_5791,N_4572,N_4792);
or U5792 (N_5792,N_4096,N_3625);
or U5793 (N_5793,N_4128,N_4339);
and U5794 (N_5794,N_4722,N_3862);
and U5795 (N_5795,N_4436,N_4590);
nand U5796 (N_5796,N_4043,N_3660);
and U5797 (N_5797,N_4274,N_4606);
nand U5798 (N_5798,N_3678,N_3815);
xor U5799 (N_5799,N_4672,N_4259);
xnor U5800 (N_5800,N_4412,N_4524);
nand U5801 (N_5801,N_4065,N_4706);
xor U5802 (N_5802,N_4099,N_3844);
nor U5803 (N_5803,N_3932,N_3789);
and U5804 (N_5804,N_4290,N_4416);
nand U5805 (N_5805,N_4300,N_4549);
and U5806 (N_5806,N_3708,N_4691);
xnor U5807 (N_5807,N_4368,N_4453);
and U5808 (N_5808,N_4587,N_3681);
and U5809 (N_5809,N_4585,N_4578);
nand U5810 (N_5810,N_4504,N_4618);
or U5811 (N_5811,N_4243,N_4127);
xnor U5812 (N_5812,N_3814,N_3939);
nand U5813 (N_5813,N_4317,N_4673);
and U5814 (N_5814,N_4630,N_4358);
and U5815 (N_5815,N_4011,N_4100);
nor U5816 (N_5816,N_4160,N_4487);
nand U5817 (N_5817,N_4044,N_4158);
or U5818 (N_5818,N_4599,N_4696);
or U5819 (N_5819,N_4305,N_4120);
and U5820 (N_5820,N_4160,N_3822);
or U5821 (N_5821,N_4527,N_3857);
or U5822 (N_5822,N_4746,N_4782);
or U5823 (N_5823,N_3706,N_4183);
nand U5824 (N_5824,N_4333,N_4547);
nor U5825 (N_5825,N_4341,N_3654);
nand U5826 (N_5826,N_4126,N_3827);
or U5827 (N_5827,N_4061,N_4116);
or U5828 (N_5828,N_3605,N_4315);
and U5829 (N_5829,N_4237,N_4758);
xor U5830 (N_5830,N_3993,N_4227);
xor U5831 (N_5831,N_4034,N_3760);
or U5832 (N_5832,N_4775,N_4396);
xnor U5833 (N_5833,N_3644,N_4759);
xor U5834 (N_5834,N_4565,N_3982);
and U5835 (N_5835,N_4096,N_4404);
and U5836 (N_5836,N_4475,N_3882);
nand U5837 (N_5837,N_3722,N_3977);
nor U5838 (N_5838,N_4350,N_4725);
nand U5839 (N_5839,N_3752,N_4581);
or U5840 (N_5840,N_4108,N_4335);
xor U5841 (N_5841,N_4172,N_4557);
or U5842 (N_5842,N_4131,N_4397);
xor U5843 (N_5843,N_4194,N_3887);
and U5844 (N_5844,N_4749,N_4527);
nor U5845 (N_5845,N_4074,N_3920);
and U5846 (N_5846,N_4288,N_4264);
nand U5847 (N_5847,N_3790,N_3729);
nand U5848 (N_5848,N_4336,N_4223);
xor U5849 (N_5849,N_4772,N_3679);
nor U5850 (N_5850,N_4380,N_4609);
xnor U5851 (N_5851,N_4301,N_3671);
nand U5852 (N_5852,N_4079,N_3874);
or U5853 (N_5853,N_3632,N_3839);
and U5854 (N_5854,N_3942,N_4180);
and U5855 (N_5855,N_4229,N_4731);
nand U5856 (N_5856,N_4014,N_3649);
or U5857 (N_5857,N_3763,N_4407);
or U5858 (N_5858,N_4527,N_4609);
and U5859 (N_5859,N_4327,N_4688);
xnor U5860 (N_5860,N_4477,N_3713);
xnor U5861 (N_5861,N_4145,N_4504);
or U5862 (N_5862,N_4391,N_4629);
and U5863 (N_5863,N_4501,N_4546);
or U5864 (N_5864,N_4202,N_4355);
xor U5865 (N_5865,N_3678,N_4459);
xnor U5866 (N_5866,N_4461,N_4605);
nor U5867 (N_5867,N_4232,N_3919);
and U5868 (N_5868,N_3737,N_4333);
and U5869 (N_5869,N_3710,N_3980);
and U5870 (N_5870,N_4706,N_4046);
xor U5871 (N_5871,N_4621,N_4547);
xor U5872 (N_5872,N_4645,N_4314);
or U5873 (N_5873,N_4118,N_3926);
or U5874 (N_5874,N_3848,N_4199);
or U5875 (N_5875,N_3693,N_3726);
xor U5876 (N_5876,N_4020,N_3889);
xnor U5877 (N_5877,N_4761,N_3679);
and U5878 (N_5878,N_4503,N_3863);
nand U5879 (N_5879,N_3946,N_4271);
or U5880 (N_5880,N_3825,N_4477);
and U5881 (N_5881,N_3864,N_4437);
or U5882 (N_5882,N_3977,N_4700);
nor U5883 (N_5883,N_3776,N_3902);
and U5884 (N_5884,N_3782,N_4788);
nand U5885 (N_5885,N_4524,N_4238);
nand U5886 (N_5886,N_4508,N_4428);
or U5887 (N_5887,N_4059,N_4166);
or U5888 (N_5888,N_3954,N_3910);
and U5889 (N_5889,N_4421,N_4643);
nor U5890 (N_5890,N_4286,N_3835);
and U5891 (N_5891,N_3791,N_3897);
xnor U5892 (N_5892,N_4084,N_3834);
or U5893 (N_5893,N_3727,N_3753);
nor U5894 (N_5894,N_3618,N_4159);
nand U5895 (N_5895,N_4607,N_4338);
nor U5896 (N_5896,N_4514,N_3997);
or U5897 (N_5897,N_4790,N_3928);
or U5898 (N_5898,N_3993,N_3721);
nand U5899 (N_5899,N_3843,N_3862);
nor U5900 (N_5900,N_4541,N_3669);
nor U5901 (N_5901,N_3864,N_3813);
xnor U5902 (N_5902,N_3778,N_4163);
nor U5903 (N_5903,N_4768,N_4568);
nor U5904 (N_5904,N_4693,N_3613);
nand U5905 (N_5905,N_3740,N_4435);
nand U5906 (N_5906,N_4671,N_4330);
or U5907 (N_5907,N_4238,N_4402);
xor U5908 (N_5908,N_3782,N_4084);
or U5909 (N_5909,N_4757,N_4308);
nand U5910 (N_5910,N_4351,N_4099);
or U5911 (N_5911,N_4518,N_4328);
nand U5912 (N_5912,N_4547,N_4376);
nor U5913 (N_5913,N_4086,N_4795);
nand U5914 (N_5914,N_4502,N_4270);
nor U5915 (N_5915,N_4196,N_4082);
nor U5916 (N_5916,N_4051,N_4584);
nand U5917 (N_5917,N_3779,N_3646);
nor U5918 (N_5918,N_3972,N_4077);
nor U5919 (N_5919,N_3627,N_4122);
or U5920 (N_5920,N_4264,N_4083);
nor U5921 (N_5921,N_3840,N_4128);
nand U5922 (N_5922,N_3826,N_4073);
nor U5923 (N_5923,N_4363,N_4113);
and U5924 (N_5924,N_4450,N_4382);
nand U5925 (N_5925,N_4518,N_3773);
nor U5926 (N_5926,N_4665,N_3684);
nand U5927 (N_5927,N_4179,N_3701);
nor U5928 (N_5928,N_4547,N_3997);
nand U5929 (N_5929,N_4063,N_4396);
nor U5930 (N_5930,N_4121,N_4071);
xor U5931 (N_5931,N_4791,N_4417);
and U5932 (N_5932,N_3869,N_4568);
nor U5933 (N_5933,N_4233,N_4733);
or U5934 (N_5934,N_4506,N_4199);
or U5935 (N_5935,N_3714,N_4508);
and U5936 (N_5936,N_4251,N_4620);
nor U5937 (N_5937,N_3841,N_3820);
and U5938 (N_5938,N_4718,N_4218);
and U5939 (N_5939,N_3951,N_4349);
xnor U5940 (N_5940,N_4605,N_4476);
or U5941 (N_5941,N_4614,N_3967);
or U5942 (N_5942,N_3686,N_3650);
and U5943 (N_5943,N_3931,N_3700);
or U5944 (N_5944,N_4652,N_4297);
or U5945 (N_5945,N_3839,N_4139);
or U5946 (N_5946,N_4044,N_3810);
nand U5947 (N_5947,N_4509,N_3913);
or U5948 (N_5948,N_3857,N_4652);
xor U5949 (N_5949,N_4424,N_4527);
or U5950 (N_5950,N_4212,N_3623);
xnor U5951 (N_5951,N_3621,N_3783);
xnor U5952 (N_5952,N_4144,N_4168);
nor U5953 (N_5953,N_4363,N_4771);
xnor U5954 (N_5954,N_3935,N_3608);
nor U5955 (N_5955,N_3851,N_3864);
nor U5956 (N_5956,N_4213,N_4627);
nand U5957 (N_5957,N_3701,N_4707);
nand U5958 (N_5958,N_4787,N_4702);
nor U5959 (N_5959,N_4216,N_4489);
nor U5960 (N_5960,N_3608,N_3965);
nor U5961 (N_5961,N_4514,N_4631);
nor U5962 (N_5962,N_3964,N_4552);
and U5963 (N_5963,N_4623,N_4152);
or U5964 (N_5964,N_4741,N_4681);
or U5965 (N_5965,N_4478,N_4680);
nor U5966 (N_5966,N_4113,N_4007);
or U5967 (N_5967,N_4282,N_4119);
and U5968 (N_5968,N_3601,N_3998);
nor U5969 (N_5969,N_4264,N_4216);
xnor U5970 (N_5970,N_4467,N_4675);
or U5971 (N_5971,N_4021,N_4033);
or U5972 (N_5972,N_3766,N_4782);
nand U5973 (N_5973,N_3832,N_4526);
or U5974 (N_5974,N_4165,N_4781);
and U5975 (N_5975,N_4444,N_4055);
and U5976 (N_5976,N_3955,N_4669);
nand U5977 (N_5977,N_3660,N_4260);
and U5978 (N_5978,N_4052,N_3967);
or U5979 (N_5979,N_4366,N_4050);
or U5980 (N_5980,N_4749,N_4626);
nand U5981 (N_5981,N_4018,N_4567);
nor U5982 (N_5982,N_3845,N_3939);
or U5983 (N_5983,N_4152,N_4670);
or U5984 (N_5984,N_4372,N_4517);
or U5985 (N_5985,N_3628,N_4073);
xor U5986 (N_5986,N_3752,N_3618);
xnor U5987 (N_5987,N_4730,N_4439);
or U5988 (N_5988,N_4279,N_3684);
or U5989 (N_5989,N_3988,N_4073);
and U5990 (N_5990,N_4596,N_4326);
and U5991 (N_5991,N_3968,N_3635);
xor U5992 (N_5992,N_3651,N_4434);
or U5993 (N_5993,N_4649,N_4030);
and U5994 (N_5994,N_4189,N_3681);
nand U5995 (N_5995,N_3959,N_3963);
nand U5996 (N_5996,N_3702,N_4241);
or U5997 (N_5997,N_3691,N_4302);
nand U5998 (N_5998,N_3728,N_4491);
and U5999 (N_5999,N_4187,N_4494);
xor U6000 (N_6000,N_5454,N_4848);
and U6001 (N_6001,N_5089,N_5813);
xor U6002 (N_6002,N_5963,N_5024);
nor U6003 (N_6003,N_5838,N_5561);
nor U6004 (N_6004,N_5753,N_5055);
and U6005 (N_6005,N_5956,N_5589);
xnor U6006 (N_6006,N_5400,N_5286);
and U6007 (N_6007,N_5904,N_5695);
xnor U6008 (N_6008,N_5258,N_4939);
and U6009 (N_6009,N_5134,N_5525);
or U6010 (N_6010,N_5802,N_5394);
or U6011 (N_6011,N_5976,N_4978);
nand U6012 (N_6012,N_5713,N_5957);
and U6013 (N_6013,N_5169,N_5056);
nor U6014 (N_6014,N_4871,N_5836);
nor U6015 (N_6015,N_4995,N_5047);
nand U6016 (N_6016,N_4919,N_5913);
or U6017 (N_6017,N_5881,N_4974);
xor U6018 (N_6018,N_4957,N_5717);
xnor U6019 (N_6019,N_5935,N_5609);
nand U6020 (N_6020,N_5355,N_4849);
nor U6021 (N_6021,N_5853,N_5673);
nor U6022 (N_6022,N_5545,N_5923);
xnor U6023 (N_6023,N_5390,N_5057);
nor U6024 (N_6024,N_5697,N_5041);
nand U6025 (N_6025,N_4963,N_5008);
or U6026 (N_6026,N_5073,N_4899);
and U6027 (N_6027,N_5377,N_5527);
or U6028 (N_6028,N_4851,N_5109);
and U6029 (N_6029,N_4937,N_5485);
nor U6030 (N_6030,N_5029,N_4825);
and U6031 (N_6031,N_5875,N_5971);
nor U6032 (N_6032,N_5471,N_5841);
and U6033 (N_6033,N_5920,N_5859);
and U6034 (N_6034,N_5621,N_4840);
nand U6035 (N_6035,N_5322,N_4812);
nor U6036 (N_6036,N_4852,N_4805);
and U6037 (N_6037,N_5227,N_5314);
and U6038 (N_6038,N_5529,N_5608);
xor U6039 (N_6039,N_5229,N_5603);
and U6040 (N_6040,N_5431,N_5679);
and U6041 (N_6041,N_5358,N_5764);
nand U6042 (N_6042,N_5905,N_5741);
or U6043 (N_6043,N_5184,N_5715);
nor U6044 (N_6044,N_5505,N_4846);
xor U6045 (N_6045,N_5486,N_5567);
nand U6046 (N_6046,N_5309,N_5623);
nor U6047 (N_6047,N_5224,N_4810);
xor U6048 (N_6048,N_5844,N_4920);
nor U6049 (N_6049,N_5404,N_5150);
nand U6050 (N_6050,N_5834,N_5676);
xor U6051 (N_6051,N_5968,N_5949);
nor U6052 (N_6052,N_4924,N_4865);
nand U6053 (N_6053,N_5279,N_5724);
and U6054 (N_6054,N_5398,N_5362);
xor U6055 (N_6055,N_5438,N_5332);
xor U6056 (N_6056,N_5062,N_5661);
nor U6057 (N_6057,N_4996,N_5852);
nand U6058 (N_6058,N_5862,N_5918);
or U6059 (N_6059,N_5705,N_5240);
nand U6060 (N_6060,N_5165,N_5936);
and U6061 (N_6061,N_5563,N_5141);
xnor U6062 (N_6062,N_5129,N_5425);
or U6063 (N_6063,N_5909,N_5696);
xnor U6064 (N_6064,N_5074,N_4886);
and U6065 (N_6065,N_5759,N_5995);
nand U6066 (N_6066,N_5095,N_5625);
nand U6067 (N_6067,N_5974,N_5843);
or U6068 (N_6068,N_5714,N_5718);
nand U6069 (N_6069,N_5234,N_5353);
or U6070 (N_6070,N_5452,N_5096);
and U6071 (N_6071,N_4972,N_4965);
and U6072 (N_6072,N_5618,N_5858);
and U6073 (N_6073,N_5285,N_5414);
nor U6074 (N_6074,N_4959,N_5916);
or U6075 (N_6075,N_5065,N_5448);
or U6076 (N_6076,N_5765,N_5778);
nor U6077 (N_6077,N_5372,N_5958);
nor U6078 (N_6078,N_5253,N_4925);
xnor U6079 (N_6079,N_5139,N_4949);
or U6080 (N_6080,N_5610,N_4822);
and U6081 (N_6081,N_5620,N_5921);
nor U6082 (N_6082,N_5788,N_5287);
nand U6083 (N_6083,N_5578,N_5756);
and U6084 (N_6084,N_5748,N_5536);
and U6085 (N_6085,N_5386,N_5543);
nand U6086 (N_6086,N_5116,N_5941);
nand U6087 (N_6087,N_4998,N_5829);
xor U6088 (N_6088,N_4975,N_5099);
xor U6089 (N_6089,N_5461,N_5734);
nand U6090 (N_6090,N_4904,N_5035);
and U6091 (N_6091,N_4860,N_5602);
and U6092 (N_6092,N_5180,N_5861);
nor U6093 (N_6093,N_4879,N_5146);
xnor U6094 (N_6094,N_5364,N_5653);
nor U6095 (N_6095,N_5850,N_5729);
xnor U6096 (N_6096,N_5367,N_5186);
nand U6097 (N_6097,N_4801,N_5190);
nor U6098 (N_6098,N_5984,N_5927);
and U6099 (N_6099,N_4945,N_5886);
nand U6100 (N_6100,N_4976,N_5412);
or U6101 (N_6101,N_5239,N_5635);
or U6102 (N_6102,N_5628,N_5710);
nand U6103 (N_6103,N_4930,N_5342);
and U6104 (N_6104,N_5330,N_5014);
or U6105 (N_6105,N_5061,N_5381);
nand U6106 (N_6106,N_5467,N_5245);
xor U6107 (N_6107,N_5553,N_5703);
or U6108 (N_6108,N_5954,N_5745);
and U6109 (N_6109,N_5274,N_5269);
or U6110 (N_6110,N_5551,N_4864);
xnor U6111 (N_6111,N_5535,N_5985);
or U6112 (N_6112,N_4923,N_5945);
nor U6113 (N_6113,N_5106,N_5893);
and U6114 (N_6114,N_5664,N_5280);
xor U6115 (N_6115,N_5012,N_5604);
or U6116 (N_6116,N_5097,N_5117);
and U6117 (N_6117,N_5494,N_5375);
xor U6118 (N_6118,N_5233,N_5906);
xor U6119 (N_6119,N_5864,N_4917);
xor U6120 (N_6120,N_5627,N_5063);
nor U6121 (N_6121,N_5994,N_4802);
nor U6122 (N_6122,N_4897,N_5633);
nor U6123 (N_6123,N_5907,N_5672);
xnor U6124 (N_6124,N_5164,N_5617);
and U6125 (N_6125,N_5052,N_5104);
nand U6126 (N_6126,N_5823,N_5284);
xor U6127 (N_6127,N_5112,N_4824);
and U6128 (N_6128,N_5903,N_4944);
nor U6129 (N_6129,N_5481,N_5201);
nand U6130 (N_6130,N_5771,N_5382);
xor U6131 (N_6131,N_5100,N_5579);
nor U6132 (N_6132,N_5347,N_5520);
and U6133 (N_6133,N_5468,N_5747);
or U6134 (N_6134,N_5365,N_4988);
nand U6135 (N_6135,N_5017,N_5986);
and U6136 (N_6136,N_5098,N_5491);
nor U6137 (N_6137,N_4818,N_5113);
nand U6138 (N_6138,N_5870,N_5121);
nand U6139 (N_6139,N_5736,N_5631);
or U6140 (N_6140,N_5781,N_5878);
xor U6141 (N_6141,N_4815,N_5163);
nor U6142 (N_6142,N_5825,N_5938);
and U6143 (N_6143,N_4985,N_5510);
and U6144 (N_6144,N_5716,N_4882);
nor U6145 (N_6145,N_5143,N_4809);
nand U6146 (N_6146,N_5289,N_5222);
nand U6147 (N_6147,N_5212,N_5706);
nand U6148 (N_6148,N_5622,N_5526);
or U6149 (N_6149,N_5389,N_4915);
xnor U6150 (N_6150,N_5880,N_5599);
or U6151 (N_6151,N_5115,N_5148);
or U6152 (N_6152,N_5203,N_4887);
or U6153 (N_6153,N_5969,N_5187);
nor U6154 (N_6154,N_5891,N_5384);
nor U6155 (N_6155,N_5130,N_4829);
and U6156 (N_6156,N_5763,N_5084);
nor U6157 (N_6157,N_5369,N_5982);
xnor U6158 (N_6158,N_4991,N_5872);
nand U6159 (N_6159,N_5449,N_5987);
nand U6160 (N_6160,N_5254,N_5940);
nor U6161 (N_6161,N_5789,N_5256);
or U6162 (N_6162,N_5442,N_5223);
and U6163 (N_6163,N_5154,N_5569);
xnor U6164 (N_6164,N_5170,N_5827);
xnor U6165 (N_6165,N_5726,N_5410);
and U6166 (N_6166,N_5686,N_5639);
nor U6167 (N_6167,N_4950,N_5460);
nand U6168 (N_6168,N_5477,N_5315);
nand U6169 (N_6169,N_5168,N_5898);
nor U6170 (N_6170,N_5496,N_5430);
or U6171 (N_6171,N_4987,N_5319);
or U6172 (N_6172,N_5721,N_4908);
nor U6173 (N_6173,N_5316,N_5798);
and U6174 (N_6174,N_5380,N_5867);
nand U6175 (N_6175,N_4940,N_5119);
or U6176 (N_6176,N_5826,N_5429);
nand U6177 (N_6177,N_5135,N_5495);
nand U6178 (N_6178,N_5027,N_5970);
nand U6179 (N_6179,N_5324,N_5281);
nand U6180 (N_6180,N_5632,N_5517);
and U6181 (N_6181,N_4916,N_5732);
nand U6182 (N_6182,N_4979,N_5470);
or U6183 (N_6183,N_5659,N_5774);
and U6184 (N_6184,N_5352,N_5719);
or U6185 (N_6185,N_5444,N_5007);
or U6186 (N_6186,N_5871,N_4835);
or U6187 (N_6187,N_5782,N_5492);
or U6188 (N_6188,N_5767,N_4855);
nor U6189 (N_6189,N_5638,N_5819);
nand U6190 (N_6190,N_5848,N_5990);
xor U6191 (N_6191,N_5205,N_5926);
and U6192 (N_6192,N_5426,N_5594);
nand U6193 (N_6193,N_5243,N_5405);
and U6194 (N_6194,N_5040,N_5683);
and U6195 (N_6195,N_5787,N_5513);
nor U6196 (N_6196,N_5651,N_4977);
nor U6197 (N_6197,N_5327,N_5952);
xnor U6198 (N_6198,N_5411,N_5593);
nor U6199 (N_6199,N_5402,N_5271);
nand U6200 (N_6200,N_5965,N_5038);
and U6201 (N_6201,N_5574,N_5733);
nor U6202 (N_6202,N_5195,N_5225);
and U6203 (N_6203,N_5354,N_5743);
nor U6204 (N_6204,N_5383,N_5152);
xnor U6205 (N_6205,N_5601,N_5300);
nand U6206 (N_6206,N_5036,N_5303);
nand U6207 (N_6207,N_5246,N_5801);
xor U6208 (N_6208,N_5413,N_4967);
nand U6209 (N_6209,N_5434,N_5919);
and U6210 (N_6210,N_4837,N_5208);
nand U6211 (N_6211,N_5888,N_4942);
nand U6212 (N_6212,N_5908,N_5291);
or U6213 (N_6213,N_5803,N_5396);
and U6214 (N_6214,N_5323,N_5453);
xor U6215 (N_6215,N_5842,N_5820);
nand U6216 (N_6216,N_5302,N_5348);
or U6217 (N_6217,N_5979,N_4956);
or U6218 (N_6218,N_5528,N_5626);
xnor U6219 (N_6219,N_4958,N_5101);
or U6220 (N_6220,N_5128,N_5232);
xnor U6221 (N_6221,N_5216,N_4885);
and U6222 (N_6222,N_5740,N_5977);
nor U6223 (N_6223,N_5972,N_5497);
or U6224 (N_6224,N_5544,N_5590);
nor U6225 (N_6225,N_5293,N_5072);
nor U6226 (N_6226,N_5147,N_5175);
xnor U6227 (N_6227,N_5435,N_4907);
or U6228 (N_6228,N_5176,N_5018);
or U6229 (N_6229,N_5554,N_5882);
xor U6230 (N_6230,N_5643,N_5215);
nor U6231 (N_6231,N_5863,N_5159);
nand U6232 (N_6232,N_5772,N_5149);
nor U6233 (N_6233,N_5070,N_5607);
and U6234 (N_6234,N_5179,N_5701);
and U6235 (N_6235,N_5276,N_5649);
and U6236 (N_6236,N_5731,N_5500);
nor U6237 (N_6237,N_5722,N_5125);
or U6238 (N_6238,N_4867,N_5524);
xor U6239 (N_6239,N_5845,N_5019);
xor U6240 (N_6240,N_4936,N_5711);
and U6241 (N_6241,N_5688,N_5983);
nor U6242 (N_6242,N_5564,N_4935);
and U6243 (N_6243,N_5887,N_5451);
or U6244 (N_6244,N_5665,N_5156);
xnor U6245 (N_6245,N_5652,N_5251);
nor U6246 (N_6246,N_5334,N_5899);
xnor U6247 (N_6247,N_5779,N_5515);
xnor U6248 (N_6248,N_4832,N_5988);
or U6249 (N_6249,N_4821,N_4933);
or U6250 (N_6250,N_5081,N_5720);
nand U6251 (N_6251,N_5847,N_5039);
nor U6252 (N_6252,N_5502,N_5546);
nor U6253 (N_6253,N_4913,N_5445);
or U6254 (N_6254,N_5944,N_5463);
or U6255 (N_6255,N_5370,N_5521);
or U6256 (N_6256,N_5091,N_5851);
nand U6257 (N_6257,N_5523,N_4961);
nand U6258 (N_6258,N_4847,N_5612);
nand U6259 (N_6259,N_5948,N_5387);
nand U6260 (N_6260,N_5237,N_5700);
nand U6261 (N_6261,N_5754,N_5160);
nor U6262 (N_6262,N_5346,N_5751);
xor U6263 (N_6263,N_5450,N_5489);
nor U6264 (N_6264,N_5548,N_5484);
nand U6265 (N_6265,N_5896,N_5832);
or U6266 (N_6266,N_5436,N_5522);
or U6267 (N_6267,N_5849,N_5951);
nor U6268 (N_6268,N_5480,N_4827);
xor U6269 (N_6269,N_4863,N_4866);
or U6270 (N_6270,N_5457,N_5110);
xnor U6271 (N_6271,N_5640,N_4836);
nor U6272 (N_6272,N_5378,N_5499);
nor U6273 (N_6273,N_5374,N_5268);
xnor U6274 (N_6274,N_5614,N_5991);
nor U6275 (N_6275,N_5576,N_5616);
or U6276 (N_6276,N_5531,N_5242);
or U6277 (N_6277,N_5644,N_5928);
nor U6278 (N_6278,N_5708,N_4898);
xnor U6279 (N_6279,N_5199,N_5808);
xnor U6280 (N_6280,N_4909,N_5955);
nor U6281 (N_6281,N_5595,N_5458);
nand U6282 (N_6282,N_5973,N_5306);
and U6283 (N_6283,N_5860,N_5959);
nand U6284 (N_6284,N_5762,N_5534);
or U6285 (N_6285,N_5680,N_5816);
xor U6286 (N_6286,N_5937,N_5547);
xor U6287 (N_6287,N_5385,N_5770);
nor U6288 (N_6288,N_5037,N_5189);
and U6289 (N_6289,N_4853,N_5768);
or U6290 (N_6290,N_4808,N_5540);
or U6291 (N_6291,N_4931,N_5158);
nand U6292 (N_6292,N_4932,N_5839);
or U6293 (N_6293,N_5259,N_5343);
nor U6294 (N_6294,N_5999,N_5173);
or U6295 (N_6295,N_5194,N_4841);
xnor U6296 (N_6296,N_5549,N_4946);
xor U6297 (N_6297,N_5992,N_5698);
nand U6298 (N_6298,N_5821,N_5566);
nor U6299 (N_6299,N_5325,N_5464);
nand U6300 (N_6300,N_4947,N_5191);
nand U6301 (N_6301,N_4928,N_5421);
xnor U6302 (N_6302,N_5138,N_5577);
xor U6303 (N_6303,N_5079,N_5118);
nand U6304 (N_6304,N_5478,N_4929);
nand U6305 (N_6305,N_5304,N_5255);
and U6306 (N_6306,N_5479,N_5877);
xnor U6307 (N_6307,N_5641,N_4970);
or U6308 (N_6308,N_5932,N_5423);
nand U6309 (N_6309,N_5294,N_5723);
nor U6310 (N_6310,N_5068,N_5010);
xor U6311 (N_6311,N_5217,N_5111);
nor U6312 (N_6312,N_4893,N_5586);
nor U6313 (N_6313,N_5766,N_5320);
xnor U6314 (N_6314,N_5911,N_5211);
or U6315 (N_6315,N_5066,N_5917);
nor U6316 (N_6316,N_4884,N_4895);
nand U6317 (N_6317,N_5830,N_5854);
xor U6318 (N_6318,N_5783,N_5814);
and U6319 (N_6319,N_4870,N_5171);
nand U6320 (N_6320,N_5933,N_5780);
or U6321 (N_6321,N_5359,N_5668);
xor U6322 (N_6322,N_4969,N_5746);
xor U6323 (N_6323,N_5312,N_5401);
nor U6324 (N_6324,N_4952,N_5082);
nor U6325 (N_6325,N_5025,N_5824);
nand U6326 (N_6326,N_5835,N_4894);
nand U6327 (N_6327,N_5086,N_5220);
xnor U6328 (N_6328,N_5556,N_5562);
and U6329 (N_6329,N_5691,N_4997);
and U6330 (N_6330,N_5376,N_5034);
or U6331 (N_6331,N_5584,N_5794);
or U6332 (N_6332,N_5596,N_5501);
nor U6333 (N_6333,N_5307,N_5178);
nand U6334 (N_6334,N_4823,N_5427);
or U6335 (N_6335,N_5252,N_5656);
or U6336 (N_6336,N_5516,N_5559);
or U6337 (N_6337,N_5388,N_5784);
or U6338 (N_6338,N_5934,N_5206);
xnor U6339 (N_6339,N_5519,N_5026);
xor U6340 (N_6340,N_5837,N_5122);
and U6341 (N_6341,N_5455,N_5810);
nor U6342 (N_6342,N_5929,N_5424);
nor U6343 (N_6343,N_5094,N_5108);
nor U6344 (N_6344,N_5157,N_5235);
nand U6345 (N_6345,N_4910,N_5188);
or U6346 (N_6346,N_5582,N_5667);
nor U6347 (N_6347,N_5231,N_4984);
or U6348 (N_6348,N_5465,N_5333);
xor U6349 (N_6349,N_5321,N_5588);
xor U6350 (N_6350,N_5060,N_5339);
nand U6351 (N_6351,N_5702,N_5511);
or U6352 (N_6352,N_5273,N_5571);
and U6353 (N_6353,N_4869,N_5092);
or U6354 (N_6354,N_5296,N_5075);
and U6355 (N_6355,N_5699,N_5264);
xor U6356 (N_6356,N_5407,N_5833);
nand U6357 (N_6357,N_5238,N_5758);
nor U6358 (N_6358,N_5730,N_5869);
or U6359 (N_6359,N_5792,N_5349);
xor U6360 (N_6360,N_5960,N_5800);
nand U6361 (N_6361,N_5504,N_5537);
xnor U6362 (N_6362,N_5379,N_5634);
nor U6363 (N_6363,N_5214,N_5822);
nor U6364 (N_6364,N_5775,N_5681);
nor U6365 (N_6365,N_4964,N_4989);
xnor U6366 (N_6366,N_4968,N_5466);
nor U6367 (N_6367,N_5914,N_5670);
xor U6368 (N_6368,N_5636,N_5755);
and U6369 (N_6369,N_5474,N_5883);
nand U6370 (N_6370,N_5915,N_5687);
or U6371 (N_6371,N_5675,N_5140);
nand U6372 (N_6372,N_5953,N_5288);
or U6373 (N_6373,N_5087,N_4814);
xor U6374 (N_6374,N_5183,N_5738);
xnor U6375 (N_6375,N_5692,N_5344);
or U6376 (N_6376,N_5704,N_5587);
and U6377 (N_6377,N_5226,N_5042);
nand U6378 (N_6378,N_5689,N_4888);
nand U6379 (N_6379,N_5200,N_4900);
xor U6380 (N_6380,N_4982,N_5488);
or U6381 (N_6381,N_5674,N_5361);
or U6382 (N_6382,N_5897,N_4838);
nor U6383 (N_6383,N_5298,N_5777);
nor U6384 (N_6384,N_4816,N_5317);
nor U6385 (N_6385,N_5210,N_5533);
and U6386 (N_6386,N_5900,N_5076);
nor U6387 (N_6387,N_5518,N_5657);
and U6388 (N_6388,N_5895,N_5003);
xor U6389 (N_6389,N_5155,N_5290);
nand U6390 (N_6390,N_5998,N_5669);
or U6391 (N_6391,N_5428,N_5126);
nor U6392 (N_6392,N_5310,N_5080);
nor U6393 (N_6393,N_5085,N_5337);
xnor U6394 (N_6394,N_5508,N_4859);
nand U6395 (N_6395,N_4806,N_5363);
xnor U6396 (N_6396,N_4912,N_5313);
and U6397 (N_6397,N_5804,N_4902);
nand U6398 (N_6398,N_5305,N_5270);
nand U6399 (N_6399,N_5114,N_5403);
nor U6400 (N_6400,N_5942,N_4800);
and U6401 (N_6401,N_5446,N_5866);
and U6402 (N_6402,N_4861,N_5542);
nor U6403 (N_6403,N_5630,N_5493);
or U6404 (N_6404,N_5760,N_5966);
xor U6405 (N_6405,N_4819,N_4872);
or U6406 (N_6406,N_5202,N_5067);
xor U6407 (N_6407,N_5658,N_4901);
and U6408 (N_6408,N_5725,N_5555);
xor U6409 (N_6409,N_5440,N_4891);
or U6410 (N_6410,N_5776,N_5439);
nand U6411 (N_6411,N_5831,N_5473);
nor U6412 (N_6412,N_5815,N_5120);
or U6413 (N_6413,N_5417,N_5006);
and U6414 (N_6414,N_5432,N_5624);
or U6415 (N_6415,N_5295,N_5786);
or U6416 (N_6416,N_5193,N_4842);
or U6417 (N_6417,N_5020,N_5811);
nor U6418 (N_6418,N_5637,N_5077);
and U6419 (N_6419,N_5030,N_5013);
nor U6420 (N_6420,N_4896,N_4986);
xor U6421 (N_6421,N_5196,N_5884);
or U6422 (N_6422,N_5694,N_5873);
nor U6423 (N_6423,N_5336,N_5538);
nor U6424 (N_6424,N_4843,N_5509);
nand U6425 (N_6425,N_4811,N_5591);
xnor U6426 (N_6426,N_5447,N_5818);
xor U6427 (N_6427,N_5943,N_4966);
nand U6428 (N_6428,N_5185,N_5650);
or U6429 (N_6429,N_5560,N_5441);
xnor U6430 (N_6430,N_5581,N_5048);
xor U6431 (N_6431,N_5498,N_5791);
nand U6432 (N_6432,N_5053,N_4889);
xnor U6433 (N_6433,N_5228,N_5373);
or U6434 (N_6434,N_5476,N_4941);
or U6435 (N_6435,N_5964,N_5272);
or U6436 (N_6436,N_4877,N_5598);
nand U6437 (N_6437,N_5318,N_4934);
nor U6438 (N_6438,N_5058,N_4954);
nand U6439 (N_6439,N_5805,N_5123);
nand U6440 (N_6440,N_5172,N_5503);
xnor U6441 (N_6441,N_5350,N_5204);
nand U6442 (N_6442,N_5459,N_5663);
or U6443 (N_6443,N_5666,N_5419);
xnor U6444 (N_6444,N_5236,N_5311);
nor U6445 (N_6445,N_5045,N_5487);
nor U6446 (N_6446,N_5677,N_5894);
and U6447 (N_6447,N_4905,N_4830);
xor U6448 (N_6448,N_4834,N_5059);
xnor U6449 (N_6449,N_5016,N_5512);
or U6450 (N_6450,N_5023,N_5865);
nor U6451 (N_6451,N_5433,N_5000);
or U6452 (N_6452,N_5795,N_5366);
and U6453 (N_6453,N_5785,N_5422);
or U6454 (N_6454,N_5153,N_5391);
nand U6455 (N_6455,N_5331,N_5064);
nand U6456 (N_6456,N_5613,N_5876);
xnor U6457 (N_6457,N_4955,N_5541);
xnor U6458 (N_6458,N_5277,N_5090);
nor U6459 (N_6459,N_5054,N_5221);
or U6460 (N_6460,N_5744,N_5292);
and U6461 (N_6461,N_5249,N_5757);
nand U6462 (N_6462,N_5338,N_4820);
and U6463 (N_6463,N_5244,N_4906);
xor U6464 (N_6464,N_5137,N_5532);
xnor U6465 (N_6465,N_4831,N_5278);
nor U6466 (N_6466,N_5167,N_4858);
nor U6467 (N_6467,N_5558,N_5133);
and U6468 (N_6468,N_4813,N_5855);
nor U6469 (N_6469,N_4857,N_4962);
nor U6470 (N_6470,N_5088,N_4807);
and U6471 (N_6471,N_5345,N_5671);
nor U6472 (N_6472,N_4953,N_5901);
and U6473 (N_6473,N_5335,N_5793);
nand U6474 (N_6474,N_4903,N_5539);
nor U6475 (N_6475,N_4868,N_5218);
and U6476 (N_6476,N_4826,N_4983);
nor U6477 (N_6477,N_5572,N_5475);
or U6478 (N_6478,N_5739,N_5326);
nor U6479 (N_6479,N_4839,N_4918);
nor U6480 (N_6480,N_5482,N_5606);
nor U6481 (N_6481,N_5071,N_4990);
nor U6482 (N_6482,N_5182,N_5127);
nand U6483 (N_6483,N_5028,N_5550);
nand U6484 (N_6484,N_5015,N_4883);
nor U6485 (N_6485,N_5409,N_4890);
nand U6486 (N_6486,N_5806,N_5997);
nor U6487 (N_6487,N_4881,N_5151);
nor U6488 (N_6488,N_5297,N_5874);
nor U6489 (N_6489,N_5809,N_5145);
and U6490 (N_6490,N_4844,N_5946);
nand U6491 (N_6491,N_5565,N_5248);
or U6492 (N_6492,N_5885,N_5207);
and U6493 (N_6493,N_5742,N_5654);
nor U6494 (N_6494,N_5962,N_5629);
xor U6495 (N_6495,N_5856,N_5769);
or U6496 (N_6496,N_5043,N_5456);
and U6497 (N_6497,N_5685,N_5910);
nand U6498 (N_6498,N_5605,N_5592);
xnor U6499 (N_6499,N_5177,N_5727);
nand U6500 (N_6500,N_5712,N_5728);
or U6501 (N_6501,N_5469,N_5230);
nand U6502 (N_6502,N_5507,N_5462);
nand U6503 (N_6503,N_5001,N_5198);
xor U6504 (N_6504,N_5597,N_4938);
xor U6505 (N_6505,N_5570,N_5580);
and U6506 (N_6506,N_5392,N_5690);
nand U6507 (N_6507,N_5993,N_5472);
and U6508 (N_6508,N_5132,N_4876);
and U6509 (N_6509,N_5046,N_5619);
nor U6510 (N_6510,N_5735,N_5161);
nor U6511 (N_6511,N_5032,N_5328);
or U6512 (N_6512,N_4845,N_5418);
or U6513 (N_6513,N_5393,N_5261);
xor U6514 (N_6514,N_5357,N_5981);
xor U6515 (N_6515,N_5051,N_5371);
xnor U6516 (N_6516,N_5351,N_4960);
or U6517 (N_6517,N_5749,N_4951);
or U6518 (N_6518,N_4828,N_5980);
nor U6519 (N_6519,N_5103,N_5506);
nor U6520 (N_6520,N_5299,N_5266);
and U6521 (N_6521,N_5005,N_5752);
or U6522 (N_6522,N_5707,N_4873);
nand U6523 (N_6523,N_5124,N_4922);
or U6524 (N_6524,N_5890,N_4803);
nor U6525 (N_6525,N_5102,N_4892);
or U6526 (N_6526,N_5583,N_5490);
and U6527 (N_6527,N_4875,N_5930);
xnor U6528 (N_6528,N_4943,N_5002);
nand U6529 (N_6529,N_5420,N_5912);
nor U6530 (N_6530,N_5049,N_5807);
and U6531 (N_6531,N_5950,N_5750);
and U6532 (N_6532,N_5166,N_5267);
xor U6533 (N_6533,N_5961,N_5967);
nor U6534 (N_6534,N_5648,N_4992);
nor U6535 (N_6535,N_4874,N_5530);
or U6536 (N_6536,N_5136,N_5615);
or U6537 (N_6537,N_4980,N_4804);
nand U6538 (N_6538,N_5263,N_5611);
and U6539 (N_6539,N_5069,N_5213);
xor U6540 (N_6540,N_4948,N_4999);
or U6541 (N_6541,N_5416,N_5131);
xnor U6542 (N_6542,N_4880,N_5209);
xnor U6543 (N_6543,N_5761,N_5879);
xnor U6544 (N_6544,N_5892,N_5360);
xnor U6545 (N_6545,N_5642,N_5797);
nand U6546 (N_6546,N_5857,N_4993);
or U6547 (N_6547,N_5265,N_5600);
nand U6548 (N_6548,N_5031,N_5368);
or U6549 (N_6549,N_5585,N_5356);
or U6550 (N_6550,N_5250,N_5573);
nor U6551 (N_6551,N_5796,N_5975);
and U6552 (N_6552,N_5406,N_5682);
nand U6553 (N_6553,N_5282,N_5437);
nor U6554 (N_6554,N_5011,N_5902);
xor U6555 (N_6555,N_5678,N_5192);
xnor U6556 (N_6556,N_5107,N_5397);
or U6557 (N_6557,N_5399,N_5050);
nor U6558 (N_6558,N_5308,N_5078);
or U6559 (N_6559,N_5799,N_5568);
and U6560 (N_6560,N_4878,N_5105);
and U6561 (N_6561,N_5925,N_5162);
and U6562 (N_6562,N_4854,N_5989);
or U6563 (N_6563,N_4973,N_4981);
and U6564 (N_6564,N_5329,N_4926);
nor U6565 (N_6565,N_5083,N_5408);
and U6566 (N_6566,N_4971,N_5033);
or U6567 (N_6567,N_4927,N_5247);
or U6568 (N_6568,N_5840,N_4850);
xnor U6569 (N_6569,N_5812,N_5645);
nor U6570 (N_6570,N_5889,N_5340);
or U6571 (N_6571,N_4994,N_5647);
and U6572 (N_6572,N_5093,N_5004);
xnor U6573 (N_6573,N_5931,N_5301);
and U6574 (N_6574,N_5939,N_5773);
xor U6575 (N_6575,N_5737,N_5197);
and U6576 (N_6576,N_4911,N_5655);
nor U6577 (N_6577,N_5846,N_5144);
and U6578 (N_6578,N_5241,N_5662);
xnor U6579 (N_6579,N_5947,N_5924);
and U6580 (N_6580,N_5817,N_5575);
xor U6581 (N_6581,N_5415,N_5022);
and U6582 (N_6582,N_5443,N_5868);
xor U6583 (N_6583,N_4856,N_5552);
and U6584 (N_6584,N_5275,N_5262);
or U6585 (N_6585,N_4914,N_5978);
nand U6586 (N_6586,N_5996,N_5009);
nand U6587 (N_6587,N_5514,N_5174);
nor U6588 (N_6588,N_5181,N_5219);
or U6589 (N_6589,N_5828,N_5021);
or U6590 (N_6590,N_5260,N_5922);
and U6591 (N_6591,N_4833,N_5557);
xnor U6592 (N_6592,N_4817,N_5684);
or U6593 (N_6593,N_5693,N_5790);
xnor U6594 (N_6594,N_5395,N_5341);
nor U6595 (N_6595,N_5709,N_5646);
nand U6596 (N_6596,N_5142,N_5044);
or U6597 (N_6597,N_5483,N_5257);
and U6598 (N_6598,N_5283,N_5660);
and U6599 (N_6599,N_4862,N_4921);
xor U6600 (N_6600,N_4807,N_5372);
xor U6601 (N_6601,N_5624,N_5108);
nor U6602 (N_6602,N_5717,N_5143);
nand U6603 (N_6603,N_5208,N_5704);
nor U6604 (N_6604,N_4926,N_5879);
nand U6605 (N_6605,N_5011,N_5695);
xnor U6606 (N_6606,N_5947,N_5080);
nor U6607 (N_6607,N_5872,N_4869);
and U6608 (N_6608,N_5751,N_5816);
nand U6609 (N_6609,N_5671,N_5153);
nand U6610 (N_6610,N_5632,N_5280);
xnor U6611 (N_6611,N_5056,N_5585);
nand U6612 (N_6612,N_5221,N_4882);
nor U6613 (N_6613,N_5588,N_4828);
nor U6614 (N_6614,N_5984,N_5811);
or U6615 (N_6615,N_4819,N_5283);
nor U6616 (N_6616,N_4862,N_5716);
nand U6617 (N_6617,N_4846,N_5420);
nand U6618 (N_6618,N_4801,N_5403);
nor U6619 (N_6619,N_4850,N_5268);
xnor U6620 (N_6620,N_5557,N_5620);
nand U6621 (N_6621,N_4940,N_5901);
xor U6622 (N_6622,N_5499,N_5690);
nand U6623 (N_6623,N_5936,N_5959);
and U6624 (N_6624,N_5969,N_5363);
xnor U6625 (N_6625,N_5938,N_5164);
or U6626 (N_6626,N_5390,N_5185);
nor U6627 (N_6627,N_5770,N_5509);
nand U6628 (N_6628,N_5700,N_4969);
nor U6629 (N_6629,N_5256,N_5486);
xor U6630 (N_6630,N_5354,N_5316);
and U6631 (N_6631,N_4892,N_4997);
and U6632 (N_6632,N_5176,N_5897);
nor U6633 (N_6633,N_4976,N_5226);
nand U6634 (N_6634,N_5145,N_5372);
and U6635 (N_6635,N_5279,N_4987);
and U6636 (N_6636,N_5120,N_5330);
and U6637 (N_6637,N_5057,N_5922);
and U6638 (N_6638,N_5078,N_5920);
xnor U6639 (N_6639,N_5667,N_4885);
or U6640 (N_6640,N_5072,N_5541);
and U6641 (N_6641,N_5469,N_5560);
nand U6642 (N_6642,N_4995,N_5099);
or U6643 (N_6643,N_5042,N_4904);
or U6644 (N_6644,N_5844,N_4955);
xnor U6645 (N_6645,N_5153,N_5296);
or U6646 (N_6646,N_5576,N_5288);
or U6647 (N_6647,N_5851,N_5611);
nor U6648 (N_6648,N_5650,N_5434);
xor U6649 (N_6649,N_4830,N_5663);
xnor U6650 (N_6650,N_5815,N_5830);
and U6651 (N_6651,N_5074,N_4855);
or U6652 (N_6652,N_5920,N_5139);
nor U6653 (N_6653,N_4984,N_5920);
xor U6654 (N_6654,N_5173,N_5188);
nand U6655 (N_6655,N_5200,N_5553);
or U6656 (N_6656,N_5064,N_5070);
and U6657 (N_6657,N_5105,N_5259);
and U6658 (N_6658,N_4812,N_4966);
or U6659 (N_6659,N_4936,N_5935);
and U6660 (N_6660,N_5797,N_5223);
or U6661 (N_6661,N_5245,N_5980);
and U6662 (N_6662,N_5384,N_5667);
xnor U6663 (N_6663,N_4981,N_5206);
xnor U6664 (N_6664,N_5238,N_5202);
xor U6665 (N_6665,N_5145,N_5576);
xor U6666 (N_6666,N_5136,N_5768);
nor U6667 (N_6667,N_5349,N_4998);
nand U6668 (N_6668,N_4871,N_5184);
nor U6669 (N_6669,N_5723,N_5504);
nand U6670 (N_6670,N_5269,N_4879);
nor U6671 (N_6671,N_5708,N_5393);
and U6672 (N_6672,N_5705,N_5305);
nor U6673 (N_6673,N_5070,N_5271);
or U6674 (N_6674,N_5692,N_5473);
nand U6675 (N_6675,N_5080,N_4869);
nor U6676 (N_6676,N_5152,N_4919);
nor U6677 (N_6677,N_5839,N_5688);
nor U6678 (N_6678,N_5674,N_5222);
xnor U6679 (N_6679,N_5661,N_4938);
or U6680 (N_6680,N_5286,N_5665);
or U6681 (N_6681,N_4986,N_5260);
nand U6682 (N_6682,N_5163,N_5402);
and U6683 (N_6683,N_5005,N_4927);
or U6684 (N_6684,N_5769,N_5478);
xor U6685 (N_6685,N_4947,N_5600);
and U6686 (N_6686,N_5864,N_5729);
nor U6687 (N_6687,N_5216,N_5531);
xor U6688 (N_6688,N_5802,N_5576);
nand U6689 (N_6689,N_5087,N_5079);
nor U6690 (N_6690,N_4981,N_5445);
xor U6691 (N_6691,N_5803,N_5698);
nand U6692 (N_6692,N_4885,N_5804);
nand U6693 (N_6693,N_4836,N_5162);
xor U6694 (N_6694,N_5406,N_5423);
xor U6695 (N_6695,N_4994,N_5988);
nor U6696 (N_6696,N_5724,N_4999);
and U6697 (N_6697,N_5635,N_5154);
nor U6698 (N_6698,N_4918,N_5352);
or U6699 (N_6699,N_5450,N_5340);
and U6700 (N_6700,N_5258,N_5140);
and U6701 (N_6701,N_5890,N_5674);
nand U6702 (N_6702,N_5136,N_5821);
nor U6703 (N_6703,N_5917,N_5474);
nand U6704 (N_6704,N_4975,N_5354);
nand U6705 (N_6705,N_4888,N_5513);
xnor U6706 (N_6706,N_5728,N_5904);
nand U6707 (N_6707,N_5282,N_4962);
and U6708 (N_6708,N_5815,N_5115);
xnor U6709 (N_6709,N_5769,N_5848);
and U6710 (N_6710,N_5175,N_5722);
nor U6711 (N_6711,N_5093,N_5868);
or U6712 (N_6712,N_5438,N_5831);
nand U6713 (N_6713,N_5790,N_4962);
and U6714 (N_6714,N_5412,N_4889);
or U6715 (N_6715,N_5400,N_5080);
nor U6716 (N_6716,N_5443,N_5016);
nand U6717 (N_6717,N_5199,N_5646);
nand U6718 (N_6718,N_4841,N_5730);
xnor U6719 (N_6719,N_5318,N_5531);
nand U6720 (N_6720,N_4975,N_5701);
and U6721 (N_6721,N_5136,N_5511);
nor U6722 (N_6722,N_5476,N_5736);
nor U6723 (N_6723,N_5359,N_5093);
nand U6724 (N_6724,N_4919,N_5789);
nor U6725 (N_6725,N_5821,N_5129);
nor U6726 (N_6726,N_5911,N_5171);
nor U6727 (N_6727,N_5245,N_5428);
nor U6728 (N_6728,N_5155,N_5568);
xor U6729 (N_6729,N_5940,N_5436);
nor U6730 (N_6730,N_5682,N_5839);
xnor U6731 (N_6731,N_4819,N_5213);
nand U6732 (N_6732,N_5271,N_5182);
nand U6733 (N_6733,N_4886,N_4852);
nor U6734 (N_6734,N_5581,N_5363);
xor U6735 (N_6735,N_5316,N_5497);
and U6736 (N_6736,N_5838,N_5872);
nand U6737 (N_6737,N_5759,N_5723);
or U6738 (N_6738,N_5562,N_5406);
and U6739 (N_6739,N_5548,N_5423);
and U6740 (N_6740,N_5795,N_5809);
and U6741 (N_6741,N_5977,N_5545);
xnor U6742 (N_6742,N_5885,N_5170);
xor U6743 (N_6743,N_5922,N_4997);
nand U6744 (N_6744,N_5505,N_5897);
nor U6745 (N_6745,N_5433,N_5110);
and U6746 (N_6746,N_5064,N_5674);
and U6747 (N_6747,N_5524,N_5174);
or U6748 (N_6748,N_5619,N_5875);
and U6749 (N_6749,N_5527,N_5267);
and U6750 (N_6750,N_5694,N_5029);
and U6751 (N_6751,N_5520,N_5677);
nor U6752 (N_6752,N_4894,N_5830);
or U6753 (N_6753,N_5895,N_4892);
nor U6754 (N_6754,N_5027,N_5296);
xor U6755 (N_6755,N_5147,N_5223);
nor U6756 (N_6756,N_5927,N_5782);
xnor U6757 (N_6757,N_4992,N_4851);
nand U6758 (N_6758,N_5491,N_5898);
nor U6759 (N_6759,N_5925,N_5745);
xnor U6760 (N_6760,N_5942,N_5954);
nand U6761 (N_6761,N_5574,N_4961);
and U6762 (N_6762,N_5553,N_5424);
xor U6763 (N_6763,N_5001,N_5171);
nand U6764 (N_6764,N_4839,N_5377);
nand U6765 (N_6765,N_5238,N_4976);
nand U6766 (N_6766,N_4822,N_4898);
or U6767 (N_6767,N_5920,N_5828);
nand U6768 (N_6768,N_5312,N_5777);
and U6769 (N_6769,N_5016,N_4967);
xor U6770 (N_6770,N_5941,N_4969);
or U6771 (N_6771,N_5106,N_5015);
nand U6772 (N_6772,N_4992,N_4954);
xor U6773 (N_6773,N_4911,N_4927);
xnor U6774 (N_6774,N_5562,N_4918);
or U6775 (N_6775,N_5146,N_5492);
nand U6776 (N_6776,N_5537,N_5617);
nor U6777 (N_6777,N_4858,N_5410);
or U6778 (N_6778,N_5992,N_5032);
nor U6779 (N_6779,N_4829,N_5791);
xor U6780 (N_6780,N_5604,N_5967);
xor U6781 (N_6781,N_5741,N_5420);
nor U6782 (N_6782,N_4846,N_5356);
nor U6783 (N_6783,N_5001,N_5084);
xor U6784 (N_6784,N_5929,N_4992);
nand U6785 (N_6785,N_4902,N_5906);
or U6786 (N_6786,N_5729,N_5005);
and U6787 (N_6787,N_5327,N_5446);
xor U6788 (N_6788,N_5542,N_5851);
xnor U6789 (N_6789,N_5122,N_4921);
xor U6790 (N_6790,N_5591,N_5137);
xor U6791 (N_6791,N_5166,N_5384);
or U6792 (N_6792,N_4913,N_5735);
nor U6793 (N_6793,N_5952,N_4948);
xnor U6794 (N_6794,N_5597,N_5948);
or U6795 (N_6795,N_5961,N_5182);
nor U6796 (N_6796,N_5730,N_4802);
xor U6797 (N_6797,N_5772,N_5839);
nand U6798 (N_6798,N_5508,N_5999);
nor U6799 (N_6799,N_5332,N_5281);
nand U6800 (N_6800,N_5498,N_4977);
nor U6801 (N_6801,N_5141,N_4924);
xnor U6802 (N_6802,N_5673,N_4964);
or U6803 (N_6803,N_5052,N_5512);
nor U6804 (N_6804,N_5325,N_5202);
nor U6805 (N_6805,N_5911,N_5529);
nor U6806 (N_6806,N_5000,N_5378);
xnor U6807 (N_6807,N_4986,N_5141);
nand U6808 (N_6808,N_5391,N_4948);
nor U6809 (N_6809,N_5783,N_5670);
nor U6810 (N_6810,N_5659,N_4824);
and U6811 (N_6811,N_5554,N_5889);
nor U6812 (N_6812,N_5978,N_5878);
nor U6813 (N_6813,N_4985,N_5690);
nor U6814 (N_6814,N_5103,N_5788);
nor U6815 (N_6815,N_5801,N_5028);
and U6816 (N_6816,N_5102,N_5599);
nand U6817 (N_6817,N_5623,N_5124);
nor U6818 (N_6818,N_5737,N_4908);
xor U6819 (N_6819,N_5518,N_5894);
or U6820 (N_6820,N_5126,N_5001);
nor U6821 (N_6821,N_5225,N_5075);
and U6822 (N_6822,N_5963,N_5306);
nand U6823 (N_6823,N_4962,N_5348);
nor U6824 (N_6824,N_5309,N_5036);
xnor U6825 (N_6825,N_5048,N_5221);
nand U6826 (N_6826,N_4920,N_5424);
and U6827 (N_6827,N_4944,N_4857);
or U6828 (N_6828,N_5565,N_5990);
nand U6829 (N_6829,N_4913,N_5606);
nor U6830 (N_6830,N_4937,N_5205);
nand U6831 (N_6831,N_5974,N_5849);
or U6832 (N_6832,N_4830,N_5167);
xnor U6833 (N_6833,N_4886,N_5282);
or U6834 (N_6834,N_5275,N_5273);
nand U6835 (N_6835,N_5694,N_4974);
or U6836 (N_6836,N_4990,N_5939);
or U6837 (N_6837,N_5324,N_5516);
xnor U6838 (N_6838,N_5093,N_5765);
nand U6839 (N_6839,N_4895,N_5599);
nand U6840 (N_6840,N_5326,N_5430);
xor U6841 (N_6841,N_5260,N_5059);
nand U6842 (N_6842,N_5800,N_5763);
nor U6843 (N_6843,N_5528,N_5676);
nor U6844 (N_6844,N_4860,N_5417);
or U6845 (N_6845,N_5793,N_5685);
or U6846 (N_6846,N_5673,N_5216);
and U6847 (N_6847,N_5530,N_5271);
nand U6848 (N_6848,N_5161,N_5455);
xor U6849 (N_6849,N_5328,N_5949);
xor U6850 (N_6850,N_4807,N_5470);
or U6851 (N_6851,N_5622,N_5951);
xnor U6852 (N_6852,N_4992,N_5486);
or U6853 (N_6853,N_5987,N_5589);
xnor U6854 (N_6854,N_4831,N_5867);
nand U6855 (N_6855,N_5295,N_5261);
nor U6856 (N_6856,N_5527,N_5866);
or U6857 (N_6857,N_5785,N_5925);
nand U6858 (N_6858,N_5247,N_5295);
and U6859 (N_6859,N_4927,N_5053);
nand U6860 (N_6860,N_5085,N_5599);
nand U6861 (N_6861,N_5837,N_5200);
nor U6862 (N_6862,N_5818,N_5443);
xor U6863 (N_6863,N_5973,N_5115);
nand U6864 (N_6864,N_5204,N_5908);
or U6865 (N_6865,N_5949,N_5908);
nor U6866 (N_6866,N_5440,N_5321);
nand U6867 (N_6867,N_5127,N_4867);
and U6868 (N_6868,N_5845,N_5224);
nor U6869 (N_6869,N_5506,N_5455);
or U6870 (N_6870,N_5667,N_5897);
and U6871 (N_6871,N_5244,N_5785);
or U6872 (N_6872,N_4821,N_5273);
nand U6873 (N_6873,N_5141,N_5917);
xnor U6874 (N_6874,N_5086,N_5950);
nand U6875 (N_6875,N_5770,N_5372);
nand U6876 (N_6876,N_5507,N_5533);
and U6877 (N_6877,N_5208,N_5799);
or U6878 (N_6878,N_5688,N_5004);
or U6879 (N_6879,N_5338,N_5467);
nor U6880 (N_6880,N_5378,N_5761);
nor U6881 (N_6881,N_5200,N_5801);
and U6882 (N_6882,N_5573,N_5102);
and U6883 (N_6883,N_5047,N_5583);
or U6884 (N_6884,N_5853,N_5680);
nand U6885 (N_6885,N_5262,N_4858);
nor U6886 (N_6886,N_5689,N_5057);
or U6887 (N_6887,N_5312,N_5682);
or U6888 (N_6888,N_5705,N_5278);
and U6889 (N_6889,N_4931,N_5090);
or U6890 (N_6890,N_5059,N_5035);
nor U6891 (N_6891,N_5354,N_4941);
xnor U6892 (N_6892,N_5274,N_5702);
or U6893 (N_6893,N_5160,N_5459);
nor U6894 (N_6894,N_5470,N_5935);
or U6895 (N_6895,N_5163,N_5184);
and U6896 (N_6896,N_5853,N_5295);
or U6897 (N_6897,N_5654,N_5390);
nor U6898 (N_6898,N_4850,N_5803);
nor U6899 (N_6899,N_5800,N_5479);
and U6900 (N_6900,N_5098,N_5873);
xnor U6901 (N_6901,N_4909,N_5246);
or U6902 (N_6902,N_4922,N_5385);
and U6903 (N_6903,N_5682,N_5344);
xor U6904 (N_6904,N_5771,N_4965);
or U6905 (N_6905,N_5353,N_5847);
or U6906 (N_6906,N_5443,N_5682);
and U6907 (N_6907,N_5793,N_5313);
and U6908 (N_6908,N_4989,N_5946);
or U6909 (N_6909,N_5662,N_5307);
or U6910 (N_6910,N_5572,N_5101);
nor U6911 (N_6911,N_4911,N_5931);
or U6912 (N_6912,N_5741,N_5097);
nand U6913 (N_6913,N_5212,N_5112);
nand U6914 (N_6914,N_5142,N_5362);
nand U6915 (N_6915,N_5324,N_5316);
or U6916 (N_6916,N_5992,N_5035);
xor U6917 (N_6917,N_5518,N_5233);
and U6918 (N_6918,N_4810,N_5418);
nand U6919 (N_6919,N_5857,N_5070);
or U6920 (N_6920,N_5647,N_5040);
or U6921 (N_6921,N_4890,N_5887);
nand U6922 (N_6922,N_5377,N_5462);
nand U6923 (N_6923,N_5862,N_5509);
or U6924 (N_6924,N_5008,N_5851);
or U6925 (N_6925,N_5228,N_4953);
and U6926 (N_6926,N_4835,N_4993);
or U6927 (N_6927,N_5589,N_5629);
nor U6928 (N_6928,N_5836,N_5338);
and U6929 (N_6929,N_5553,N_5505);
nor U6930 (N_6930,N_5503,N_4808);
and U6931 (N_6931,N_5507,N_5276);
or U6932 (N_6932,N_5238,N_5104);
or U6933 (N_6933,N_5653,N_5032);
nor U6934 (N_6934,N_5286,N_4818);
nor U6935 (N_6935,N_5246,N_5406);
xnor U6936 (N_6936,N_5167,N_5113);
nor U6937 (N_6937,N_4926,N_5406);
or U6938 (N_6938,N_5113,N_5768);
nor U6939 (N_6939,N_5338,N_5295);
nand U6940 (N_6940,N_5266,N_5432);
xor U6941 (N_6941,N_5562,N_5292);
or U6942 (N_6942,N_5417,N_5239);
or U6943 (N_6943,N_5732,N_4942);
xor U6944 (N_6944,N_5642,N_5112);
nand U6945 (N_6945,N_5491,N_5962);
nand U6946 (N_6946,N_5686,N_5261);
nor U6947 (N_6947,N_5300,N_5773);
and U6948 (N_6948,N_5856,N_5116);
xor U6949 (N_6949,N_5242,N_4969);
or U6950 (N_6950,N_5004,N_5932);
nor U6951 (N_6951,N_5625,N_5958);
or U6952 (N_6952,N_5138,N_5845);
or U6953 (N_6953,N_5006,N_5316);
or U6954 (N_6954,N_5989,N_5856);
nor U6955 (N_6955,N_4833,N_5693);
xor U6956 (N_6956,N_5135,N_5891);
and U6957 (N_6957,N_5508,N_4970);
or U6958 (N_6958,N_5157,N_5163);
and U6959 (N_6959,N_5359,N_5734);
nor U6960 (N_6960,N_4852,N_5623);
xnor U6961 (N_6961,N_5973,N_5998);
xnor U6962 (N_6962,N_5944,N_5559);
or U6963 (N_6963,N_5638,N_5549);
xnor U6964 (N_6964,N_5613,N_5768);
or U6965 (N_6965,N_5717,N_5660);
nor U6966 (N_6966,N_5369,N_5154);
nor U6967 (N_6967,N_5584,N_5171);
nor U6968 (N_6968,N_5226,N_5197);
and U6969 (N_6969,N_4870,N_5472);
nor U6970 (N_6970,N_5080,N_5361);
xor U6971 (N_6971,N_5721,N_4934);
or U6972 (N_6972,N_5422,N_5893);
nor U6973 (N_6973,N_5657,N_5700);
or U6974 (N_6974,N_5771,N_5403);
or U6975 (N_6975,N_5217,N_5228);
and U6976 (N_6976,N_5568,N_5153);
or U6977 (N_6977,N_4880,N_4884);
nor U6978 (N_6978,N_5773,N_5492);
or U6979 (N_6979,N_5999,N_5000);
nor U6980 (N_6980,N_5573,N_5593);
xnor U6981 (N_6981,N_5494,N_4990);
xnor U6982 (N_6982,N_5376,N_5719);
nand U6983 (N_6983,N_5783,N_4901);
and U6984 (N_6984,N_5330,N_5043);
or U6985 (N_6985,N_4906,N_4817);
xor U6986 (N_6986,N_5446,N_4856);
xnor U6987 (N_6987,N_5571,N_5583);
and U6988 (N_6988,N_5639,N_5910);
and U6989 (N_6989,N_5228,N_5019);
nand U6990 (N_6990,N_5935,N_5593);
xor U6991 (N_6991,N_4993,N_4812);
nor U6992 (N_6992,N_5670,N_5785);
nand U6993 (N_6993,N_4855,N_5956);
nand U6994 (N_6994,N_4913,N_5477);
nand U6995 (N_6995,N_4867,N_5479);
or U6996 (N_6996,N_5960,N_5105);
nor U6997 (N_6997,N_5867,N_5572);
nor U6998 (N_6998,N_5672,N_5408);
or U6999 (N_6999,N_4977,N_5810);
nor U7000 (N_7000,N_5093,N_5138);
xnor U7001 (N_7001,N_5243,N_5679);
and U7002 (N_7002,N_5615,N_4998);
and U7003 (N_7003,N_5343,N_4962);
nand U7004 (N_7004,N_5471,N_5207);
and U7005 (N_7005,N_5692,N_5678);
or U7006 (N_7006,N_5668,N_5317);
or U7007 (N_7007,N_5694,N_5560);
or U7008 (N_7008,N_5830,N_5784);
nor U7009 (N_7009,N_5469,N_4968);
nor U7010 (N_7010,N_5070,N_5292);
or U7011 (N_7011,N_5546,N_5586);
or U7012 (N_7012,N_5969,N_4957);
xnor U7013 (N_7013,N_5490,N_5926);
nand U7014 (N_7014,N_5078,N_5828);
or U7015 (N_7015,N_4889,N_5694);
or U7016 (N_7016,N_5289,N_5337);
nand U7017 (N_7017,N_5450,N_5599);
xor U7018 (N_7018,N_5410,N_5535);
nor U7019 (N_7019,N_5756,N_5970);
nor U7020 (N_7020,N_4867,N_5300);
nor U7021 (N_7021,N_5578,N_5713);
or U7022 (N_7022,N_5466,N_5272);
nor U7023 (N_7023,N_5113,N_5376);
nor U7024 (N_7024,N_4828,N_5294);
and U7025 (N_7025,N_5719,N_5245);
nand U7026 (N_7026,N_5719,N_5828);
nor U7027 (N_7027,N_5842,N_5074);
or U7028 (N_7028,N_4936,N_5948);
nor U7029 (N_7029,N_5487,N_5083);
nand U7030 (N_7030,N_5153,N_5362);
or U7031 (N_7031,N_5999,N_4945);
nor U7032 (N_7032,N_5447,N_5827);
nand U7033 (N_7033,N_4983,N_5316);
xnor U7034 (N_7034,N_4847,N_5691);
xnor U7035 (N_7035,N_5622,N_5446);
nor U7036 (N_7036,N_5114,N_5151);
xnor U7037 (N_7037,N_5146,N_5935);
xor U7038 (N_7038,N_5453,N_5898);
xor U7039 (N_7039,N_5981,N_5095);
nor U7040 (N_7040,N_5968,N_4948);
nand U7041 (N_7041,N_4800,N_5130);
xor U7042 (N_7042,N_5419,N_5559);
and U7043 (N_7043,N_5524,N_5762);
nor U7044 (N_7044,N_5733,N_5644);
nor U7045 (N_7045,N_5627,N_5755);
and U7046 (N_7046,N_4970,N_5110);
nand U7047 (N_7047,N_5944,N_5143);
nand U7048 (N_7048,N_4892,N_5708);
xnor U7049 (N_7049,N_5305,N_5844);
and U7050 (N_7050,N_5133,N_5168);
nand U7051 (N_7051,N_5643,N_5315);
or U7052 (N_7052,N_5234,N_4976);
and U7053 (N_7053,N_5925,N_5618);
or U7054 (N_7054,N_5604,N_5726);
nand U7055 (N_7055,N_5380,N_4997);
nor U7056 (N_7056,N_4830,N_5744);
and U7057 (N_7057,N_5885,N_5173);
and U7058 (N_7058,N_5418,N_4873);
nor U7059 (N_7059,N_4814,N_5150);
and U7060 (N_7060,N_5220,N_5659);
or U7061 (N_7061,N_5499,N_5432);
nor U7062 (N_7062,N_5384,N_5360);
and U7063 (N_7063,N_5067,N_4935);
nand U7064 (N_7064,N_5671,N_4944);
nand U7065 (N_7065,N_5431,N_5017);
nor U7066 (N_7066,N_4822,N_5748);
or U7067 (N_7067,N_4964,N_5290);
nand U7068 (N_7068,N_5620,N_5889);
nor U7069 (N_7069,N_5427,N_5795);
or U7070 (N_7070,N_4852,N_4870);
nand U7071 (N_7071,N_5544,N_5188);
or U7072 (N_7072,N_5511,N_5357);
nor U7073 (N_7073,N_5947,N_5172);
and U7074 (N_7074,N_5936,N_5483);
nand U7075 (N_7075,N_5365,N_5224);
nand U7076 (N_7076,N_4988,N_5754);
xor U7077 (N_7077,N_5015,N_5393);
xnor U7078 (N_7078,N_5589,N_5900);
or U7079 (N_7079,N_4970,N_5933);
or U7080 (N_7080,N_5424,N_5648);
xnor U7081 (N_7081,N_5422,N_5688);
nor U7082 (N_7082,N_5487,N_5425);
and U7083 (N_7083,N_5392,N_5822);
and U7084 (N_7084,N_5896,N_5494);
and U7085 (N_7085,N_5259,N_5861);
and U7086 (N_7086,N_5094,N_4872);
and U7087 (N_7087,N_4981,N_5033);
and U7088 (N_7088,N_5141,N_5153);
nor U7089 (N_7089,N_5177,N_5000);
and U7090 (N_7090,N_5740,N_5942);
and U7091 (N_7091,N_5115,N_5446);
nor U7092 (N_7092,N_4979,N_5976);
xor U7093 (N_7093,N_5293,N_5893);
or U7094 (N_7094,N_5074,N_5095);
xnor U7095 (N_7095,N_5415,N_5844);
nand U7096 (N_7096,N_4901,N_4908);
and U7097 (N_7097,N_4926,N_5702);
nand U7098 (N_7098,N_5006,N_5376);
nor U7099 (N_7099,N_5267,N_5886);
nand U7100 (N_7100,N_5671,N_5542);
xnor U7101 (N_7101,N_5199,N_5968);
or U7102 (N_7102,N_5013,N_4906);
or U7103 (N_7103,N_5666,N_5186);
nor U7104 (N_7104,N_5375,N_5251);
or U7105 (N_7105,N_5086,N_4909);
xor U7106 (N_7106,N_5191,N_5680);
or U7107 (N_7107,N_5602,N_5568);
and U7108 (N_7108,N_5401,N_5394);
xnor U7109 (N_7109,N_5311,N_5487);
xnor U7110 (N_7110,N_5575,N_4882);
xor U7111 (N_7111,N_5691,N_4801);
and U7112 (N_7112,N_4995,N_5384);
nand U7113 (N_7113,N_4843,N_5120);
nor U7114 (N_7114,N_4997,N_5158);
xnor U7115 (N_7115,N_5984,N_4967);
and U7116 (N_7116,N_5692,N_4997);
nor U7117 (N_7117,N_5447,N_5351);
nor U7118 (N_7118,N_5722,N_5758);
and U7119 (N_7119,N_5563,N_5835);
and U7120 (N_7120,N_4811,N_5953);
nor U7121 (N_7121,N_5712,N_5348);
nor U7122 (N_7122,N_5701,N_5484);
and U7123 (N_7123,N_5738,N_5072);
and U7124 (N_7124,N_4855,N_5187);
nor U7125 (N_7125,N_5897,N_5691);
and U7126 (N_7126,N_5850,N_4812);
and U7127 (N_7127,N_4830,N_5193);
nand U7128 (N_7128,N_5754,N_5456);
nor U7129 (N_7129,N_5000,N_5625);
and U7130 (N_7130,N_5783,N_4859);
xor U7131 (N_7131,N_5826,N_5671);
nor U7132 (N_7132,N_4807,N_5778);
xor U7133 (N_7133,N_5397,N_4988);
xor U7134 (N_7134,N_5841,N_5185);
nor U7135 (N_7135,N_5591,N_5797);
and U7136 (N_7136,N_5579,N_5795);
nor U7137 (N_7137,N_4904,N_4871);
nand U7138 (N_7138,N_5204,N_5890);
xnor U7139 (N_7139,N_5239,N_5789);
nand U7140 (N_7140,N_5070,N_4921);
or U7141 (N_7141,N_5672,N_5130);
or U7142 (N_7142,N_5976,N_5712);
or U7143 (N_7143,N_5671,N_5509);
nand U7144 (N_7144,N_4843,N_5549);
xnor U7145 (N_7145,N_5791,N_5927);
nand U7146 (N_7146,N_5413,N_5974);
nor U7147 (N_7147,N_5958,N_5459);
nor U7148 (N_7148,N_4883,N_4898);
or U7149 (N_7149,N_5319,N_5444);
or U7150 (N_7150,N_5168,N_5495);
and U7151 (N_7151,N_5971,N_5779);
nor U7152 (N_7152,N_4996,N_5043);
xnor U7153 (N_7153,N_5708,N_5691);
or U7154 (N_7154,N_5693,N_5470);
nor U7155 (N_7155,N_4991,N_5562);
nor U7156 (N_7156,N_5181,N_5000);
xnor U7157 (N_7157,N_5025,N_5595);
xnor U7158 (N_7158,N_5451,N_5848);
and U7159 (N_7159,N_5575,N_5856);
nand U7160 (N_7160,N_5964,N_5776);
and U7161 (N_7161,N_5847,N_5585);
xor U7162 (N_7162,N_5206,N_5381);
nand U7163 (N_7163,N_5833,N_5032);
and U7164 (N_7164,N_5632,N_4939);
nand U7165 (N_7165,N_5366,N_4912);
nand U7166 (N_7166,N_5910,N_5773);
nor U7167 (N_7167,N_5355,N_5545);
nand U7168 (N_7168,N_5397,N_4836);
or U7169 (N_7169,N_5528,N_4958);
nor U7170 (N_7170,N_5469,N_5799);
nor U7171 (N_7171,N_5919,N_5230);
and U7172 (N_7172,N_5912,N_5324);
or U7173 (N_7173,N_5544,N_5652);
or U7174 (N_7174,N_4996,N_5925);
nor U7175 (N_7175,N_4894,N_5847);
xnor U7176 (N_7176,N_5257,N_5985);
xnor U7177 (N_7177,N_5450,N_4977);
and U7178 (N_7178,N_4887,N_5803);
nor U7179 (N_7179,N_5378,N_5889);
nor U7180 (N_7180,N_5611,N_5243);
and U7181 (N_7181,N_4961,N_5733);
nand U7182 (N_7182,N_5416,N_5232);
and U7183 (N_7183,N_4882,N_5825);
and U7184 (N_7184,N_5232,N_5181);
or U7185 (N_7185,N_5970,N_5457);
or U7186 (N_7186,N_5700,N_5728);
or U7187 (N_7187,N_5172,N_5517);
xor U7188 (N_7188,N_5375,N_5439);
nor U7189 (N_7189,N_5504,N_5333);
and U7190 (N_7190,N_4872,N_5622);
nor U7191 (N_7191,N_5475,N_5039);
and U7192 (N_7192,N_5074,N_5576);
or U7193 (N_7193,N_4850,N_4978);
and U7194 (N_7194,N_5661,N_5304);
nand U7195 (N_7195,N_4854,N_4884);
nand U7196 (N_7196,N_5150,N_5736);
nand U7197 (N_7197,N_4872,N_5979);
nor U7198 (N_7198,N_5474,N_5826);
nor U7199 (N_7199,N_4825,N_5248);
or U7200 (N_7200,N_6644,N_6654);
nand U7201 (N_7201,N_6300,N_6801);
nor U7202 (N_7202,N_6894,N_6501);
and U7203 (N_7203,N_6678,N_6960);
xnor U7204 (N_7204,N_6477,N_7033);
nor U7205 (N_7205,N_6151,N_7168);
nand U7206 (N_7206,N_6819,N_6861);
nand U7207 (N_7207,N_6561,N_7175);
xor U7208 (N_7208,N_6294,N_6718);
nand U7209 (N_7209,N_6295,N_7012);
nor U7210 (N_7210,N_6145,N_6345);
or U7211 (N_7211,N_6549,N_6122);
nor U7212 (N_7212,N_6408,N_6733);
and U7213 (N_7213,N_6053,N_6916);
nand U7214 (N_7214,N_6160,N_6860);
nor U7215 (N_7215,N_6218,N_7190);
nand U7216 (N_7216,N_7112,N_6926);
nor U7217 (N_7217,N_6986,N_6072);
or U7218 (N_7218,N_6080,N_7151);
nand U7219 (N_7219,N_6128,N_6040);
nand U7220 (N_7220,N_6256,N_6748);
and U7221 (N_7221,N_6852,N_6132);
nand U7222 (N_7222,N_7071,N_6747);
nor U7223 (N_7223,N_6090,N_6514);
nand U7224 (N_7224,N_6872,N_6778);
nor U7225 (N_7225,N_6254,N_7008);
nor U7226 (N_7226,N_6486,N_7022);
nor U7227 (N_7227,N_6194,N_6837);
and U7228 (N_7228,N_6634,N_6683);
nand U7229 (N_7229,N_6669,N_6436);
or U7230 (N_7230,N_6279,N_6878);
and U7231 (N_7231,N_6223,N_6662);
nor U7232 (N_7232,N_6923,N_6035);
xor U7233 (N_7233,N_6133,N_6949);
or U7234 (N_7234,N_7040,N_6285);
xor U7235 (N_7235,N_7171,N_6025);
or U7236 (N_7236,N_6731,N_6277);
and U7237 (N_7237,N_6399,N_6234);
nor U7238 (N_7238,N_6444,N_6425);
xnor U7239 (N_7239,N_6435,N_6512);
and U7240 (N_7240,N_6934,N_6608);
and U7241 (N_7241,N_7153,N_6150);
and U7242 (N_7242,N_7166,N_6557);
and U7243 (N_7243,N_6970,N_6955);
and U7244 (N_7244,N_6163,N_6572);
nor U7245 (N_7245,N_6773,N_7149);
xnor U7246 (N_7246,N_6362,N_7034);
and U7247 (N_7247,N_6258,N_6140);
xor U7248 (N_7248,N_6148,N_6830);
nor U7249 (N_7249,N_6244,N_6762);
xnor U7250 (N_7250,N_7030,N_7066);
and U7251 (N_7251,N_6403,N_6288);
and U7252 (N_7252,N_6152,N_6793);
and U7253 (N_7253,N_6219,N_6702);
and U7254 (N_7254,N_7142,N_6430);
nand U7255 (N_7255,N_6344,N_7067);
and U7256 (N_7256,N_6456,N_6680);
nor U7257 (N_7257,N_6143,N_7000);
or U7258 (N_7258,N_6776,N_6112);
nand U7259 (N_7259,N_6202,N_6497);
xor U7260 (N_7260,N_6114,N_6358);
nor U7261 (N_7261,N_7177,N_7176);
and U7262 (N_7262,N_6742,N_6336);
and U7263 (N_7263,N_6893,N_6653);
or U7264 (N_7264,N_6078,N_6792);
xor U7265 (N_7265,N_6469,N_6439);
xor U7266 (N_7266,N_6799,N_6382);
and U7267 (N_7267,N_6073,N_6999);
or U7268 (N_7268,N_6730,N_6782);
and U7269 (N_7269,N_6790,N_6154);
or U7270 (N_7270,N_7156,N_6343);
nand U7271 (N_7271,N_6593,N_6672);
or U7272 (N_7272,N_6282,N_7100);
xor U7273 (N_7273,N_7121,N_6175);
nor U7274 (N_7274,N_6475,N_6856);
nand U7275 (N_7275,N_6009,N_7003);
and U7276 (N_7276,N_6900,N_6927);
nor U7277 (N_7277,N_6650,N_6239);
nand U7278 (N_7278,N_7126,N_6104);
xnor U7279 (N_7279,N_6166,N_7078);
xnor U7280 (N_7280,N_6183,N_7089);
nor U7281 (N_7281,N_6178,N_6798);
or U7282 (N_7282,N_6576,N_6979);
nand U7283 (N_7283,N_7140,N_6422);
xnor U7284 (N_7284,N_6041,N_6481);
nor U7285 (N_7285,N_6310,N_6100);
or U7286 (N_7286,N_6741,N_6325);
xnor U7287 (N_7287,N_6626,N_6119);
nor U7288 (N_7288,N_6751,N_6535);
nand U7289 (N_7289,N_6800,N_6048);
nor U7290 (N_7290,N_6779,N_6752);
and U7291 (N_7291,N_6516,N_6489);
xor U7292 (N_7292,N_6677,N_7026);
xor U7293 (N_7293,N_6618,N_7104);
xnor U7294 (N_7294,N_7145,N_6997);
nor U7295 (N_7295,N_6468,N_6607);
nor U7296 (N_7296,N_6319,N_6524);
xor U7297 (N_7297,N_7125,N_6307);
nor U7298 (N_7298,N_6598,N_6404);
nand U7299 (N_7299,N_6391,N_6571);
or U7300 (N_7300,N_6587,N_6933);
or U7301 (N_7301,N_6974,N_7063);
nor U7302 (N_7302,N_6724,N_7198);
nor U7303 (N_7303,N_6236,N_7082);
xnor U7304 (N_7304,N_7095,N_7130);
or U7305 (N_7305,N_6763,N_6428);
xnor U7306 (N_7306,N_6116,N_6541);
xnor U7307 (N_7307,N_6186,N_6588);
or U7308 (N_7308,N_6983,N_6103);
and U7309 (N_7309,N_6780,N_6994);
and U7310 (N_7310,N_6595,N_6210);
nor U7311 (N_7311,N_6612,N_6509);
xnor U7312 (N_7312,N_6251,N_6919);
nand U7313 (N_7313,N_6450,N_7194);
and U7314 (N_7314,N_6111,N_6328);
xor U7315 (N_7315,N_6392,N_6615);
or U7316 (N_7316,N_6975,N_6357);
or U7317 (N_7317,N_6250,N_6705);
and U7318 (N_7318,N_6135,N_6338);
nand U7319 (N_7319,N_6658,N_6764);
nand U7320 (N_7320,N_6364,N_6014);
xnor U7321 (N_7321,N_6192,N_6268);
xnor U7322 (N_7322,N_6701,N_6846);
xor U7323 (N_7323,N_6023,N_6094);
nor U7324 (N_7324,N_6857,N_6998);
and U7325 (N_7325,N_6959,N_6036);
xnor U7326 (N_7326,N_6670,N_7010);
nand U7327 (N_7327,N_6520,N_6305);
or U7328 (N_7328,N_6432,N_6273);
and U7329 (N_7329,N_6840,N_6944);
or U7330 (N_7330,N_6452,N_6329);
and U7331 (N_7331,N_6229,N_6322);
or U7332 (N_7332,N_6067,N_7132);
xnor U7333 (N_7333,N_6573,N_6704);
and U7334 (N_7334,N_6353,N_6636);
or U7335 (N_7335,N_6815,N_6579);
xnor U7336 (N_7336,N_6113,N_6264);
nor U7337 (N_7337,N_6333,N_6966);
xor U7338 (N_7338,N_6605,N_6191);
nor U7339 (N_7339,N_6496,N_7119);
and U7340 (N_7340,N_6597,N_7094);
nor U7341 (N_7341,N_6941,N_6086);
or U7342 (N_7342,N_6845,N_6739);
and U7343 (N_7343,N_6811,N_6942);
nand U7344 (N_7344,N_6007,N_7160);
or U7345 (N_7345,N_7157,N_6045);
and U7346 (N_7346,N_6199,N_6249);
xor U7347 (N_7347,N_6577,N_6813);
and U7348 (N_7348,N_6320,N_6686);
or U7349 (N_7349,N_6352,N_7128);
nand U7350 (N_7350,N_6386,N_6698);
nor U7351 (N_7351,N_7009,N_6914);
nand U7352 (N_7352,N_7045,N_6717);
or U7353 (N_7353,N_6296,N_6483);
or U7354 (N_7354,N_6374,N_7088);
and U7355 (N_7355,N_6185,N_6238);
nor U7356 (N_7356,N_7187,N_6476);
xnor U7357 (N_7357,N_6370,N_7133);
nand U7358 (N_7358,N_6899,N_7056);
and U7359 (N_7359,N_7087,N_6534);
nand U7360 (N_7360,N_6141,N_6548);
and U7361 (N_7361,N_7159,N_6714);
or U7362 (N_7362,N_6648,N_6440);
and U7363 (N_7363,N_6095,N_6075);
nand U7364 (N_7364,N_7037,N_6537);
and U7365 (N_7365,N_6695,N_6463);
xor U7366 (N_7366,N_7058,N_6129);
or U7367 (N_7367,N_6335,N_7189);
or U7368 (N_7368,N_6225,N_6963);
and U7369 (N_7369,N_6233,N_7025);
and U7370 (N_7370,N_6580,N_6124);
nor U7371 (N_7371,N_6954,N_7069);
or U7372 (N_7372,N_6976,N_6876);
nand U7373 (N_7373,N_6110,N_6118);
xor U7374 (N_7374,N_6874,N_6720);
nand U7375 (N_7375,N_6130,N_6749);
nand U7376 (N_7376,N_6995,N_6126);
nor U7377 (N_7377,N_6044,N_6624);
nor U7378 (N_7378,N_6049,N_6804);
xor U7379 (N_7379,N_6550,N_6885);
xor U7380 (N_7380,N_6667,N_6409);
nor U7381 (N_7381,N_7174,N_7050);
nand U7382 (N_7382,N_7154,N_7091);
and U7383 (N_7383,N_6865,N_6292);
and U7384 (N_7384,N_6841,N_6488);
or U7385 (N_7385,N_6434,N_7110);
or U7386 (N_7386,N_6581,N_6827);
nand U7387 (N_7387,N_6613,N_6478);
and U7388 (N_7388,N_6886,N_6082);
nand U7389 (N_7389,N_6659,N_6835);
or U7390 (N_7390,N_6671,N_6473);
nor U7391 (N_7391,N_6787,N_6125);
and U7392 (N_7392,N_6931,N_6538);
nand U7393 (N_7393,N_7021,N_6155);
xor U7394 (N_7394,N_7074,N_6853);
nor U7395 (N_7395,N_6190,N_6508);
or U7396 (N_7396,N_6068,N_6136);
xnor U7397 (N_7397,N_6372,N_6586);
nor U7398 (N_7398,N_6661,N_6204);
xnor U7399 (N_7399,N_6105,N_6065);
xor U7400 (N_7400,N_6891,N_6467);
nand U7401 (N_7401,N_6389,N_7014);
and U7402 (N_7402,N_6500,N_6039);
or U7403 (N_7403,N_6551,N_6211);
or U7404 (N_7404,N_6308,N_6716);
and U7405 (N_7405,N_6755,N_6699);
or U7406 (N_7406,N_6521,N_6957);
nand U7407 (N_7407,N_6474,N_7013);
nor U7408 (N_7408,N_6775,N_7053);
nor U7409 (N_7409,N_6879,N_6276);
nand U7410 (N_7410,N_6750,N_6123);
and U7411 (N_7411,N_6361,N_7134);
or U7412 (N_7412,N_6611,N_6760);
or U7413 (N_7413,N_7081,N_6664);
nand U7414 (N_7414,N_6226,N_6363);
xor U7415 (N_7415,N_6688,N_6585);
or U7416 (N_7416,N_6419,N_6317);
nand U7417 (N_7417,N_7120,N_7020);
nand U7418 (N_7418,N_6070,N_6703);
xnor U7419 (N_7419,N_6943,N_6263);
nor U7420 (N_7420,N_7011,N_6937);
xnor U7421 (N_7421,N_6138,N_7167);
xnor U7422 (N_7422,N_6584,N_7105);
and U7423 (N_7423,N_6545,N_6058);
nand U7424 (N_7424,N_6795,N_6806);
and U7425 (N_7425,N_6540,N_7085);
xnor U7426 (N_7426,N_7035,N_6640);
nor U7427 (N_7427,N_6553,N_6245);
and U7428 (N_7428,N_6694,N_6884);
or U7429 (N_7429,N_6479,N_6085);
and U7430 (N_7430,N_6283,N_6224);
nand U7431 (N_7431,N_6794,N_6988);
and U7432 (N_7432,N_6518,N_6629);
xnor U7433 (N_7433,N_7129,N_6134);
nand U7434 (N_7434,N_6930,N_6565);
nor U7435 (N_7435,N_6797,N_7170);
and U7436 (N_7436,N_6301,N_6863);
and U7437 (N_7437,N_6708,N_6610);
or U7438 (N_7438,N_6940,N_6924);
and U7439 (N_7439,N_6334,N_6599);
or U7440 (N_7440,N_6167,N_6395);
or U7441 (N_7441,N_6341,N_6063);
or U7442 (N_7442,N_6563,N_6472);
or U7443 (N_7443,N_6713,N_6982);
and U7444 (N_7444,N_6120,N_6482);
or U7445 (N_7445,N_7072,N_6438);
and U7446 (N_7446,N_6836,N_7183);
nor U7447 (N_7447,N_6866,N_6616);
xnor U7448 (N_7448,N_6366,N_6875);
and U7449 (N_7449,N_6981,N_6139);
or U7450 (N_7450,N_6871,N_6069);
or U7451 (N_7451,N_6102,N_6589);
or U7452 (N_7452,N_6614,N_6423);
and U7453 (N_7453,N_6715,N_6992);
and U7454 (N_7454,N_6619,N_6868);
and U7455 (N_7455,N_6003,N_6777);
or U7456 (N_7456,N_6099,N_6850);
nand U7457 (N_7457,N_7131,N_6071);
or U7458 (N_7458,N_6195,N_7114);
xnor U7459 (N_7459,N_6212,N_6280);
and U7460 (N_7460,N_6769,N_6359);
xnor U7461 (N_7461,N_6485,N_6274);
xor U7462 (N_7462,N_6842,N_6735);
and U7463 (N_7463,N_6643,N_6889);
and U7464 (N_7464,N_6744,N_6625);
or U7465 (N_7465,N_6617,N_6037);
nor U7466 (N_7466,N_7028,N_6847);
xor U7467 (N_7467,N_6767,N_6913);
xnor U7468 (N_7468,N_6005,N_6843);
xnor U7469 (N_7469,N_7073,N_6869);
xnor U7470 (N_7470,N_6887,N_6367);
nand U7471 (N_7471,N_6832,N_6791);
xor U7472 (N_7472,N_7099,N_6505);
and U7473 (N_7473,N_6969,N_7164);
nand U7474 (N_7474,N_6691,N_7017);
nor U7475 (N_7475,N_7179,N_6552);
nor U7476 (N_7476,N_6302,N_6405);
or U7477 (N_7477,N_6412,N_6407);
nand U7478 (N_7478,N_6024,N_6312);
nand U7479 (N_7479,N_6905,N_6948);
or U7480 (N_7480,N_6493,N_7075);
and U7481 (N_7481,N_6162,N_6465);
xor U7482 (N_7482,N_6001,N_6360);
and U7483 (N_7483,N_6029,N_6645);
or U7484 (N_7484,N_6569,N_6725);
nand U7485 (N_7485,N_7143,N_7098);
and U7486 (N_7486,N_6161,N_6578);
or U7487 (N_7487,N_6838,N_6093);
xor U7488 (N_7488,N_6401,N_6179);
xor U7489 (N_7489,N_6098,N_6622);
and U7490 (N_7490,N_6621,N_6968);
nand U7491 (N_7491,N_6303,N_6384);
or U7492 (N_7492,N_6796,N_6503);
and U7493 (N_7493,N_7158,N_6042);
and U7494 (N_7494,N_6700,N_7042);
nand U7495 (N_7495,N_6892,N_6453);
xor U7496 (N_7496,N_6530,N_6906);
nand U7497 (N_7497,N_7006,N_6709);
or U7498 (N_7498,N_6925,N_6809);
nor U7499 (N_7499,N_6375,N_6376);
and U7500 (N_7500,N_6117,N_7047);
xnor U7501 (N_7501,N_6396,N_6447);
xor U7502 (N_7502,N_7004,N_6682);
nand U7503 (N_7503,N_7052,N_6693);
xnor U7504 (N_7504,N_6373,N_7064);
and U7505 (N_7505,N_6696,N_6187);
nor U7506 (N_7506,N_7137,N_6921);
nand U7507 (N_7507,N_6985,N_6172);
nor U7508 (N_7508,N_6337,N_6737);
and U7509 (N_7509,N_6026,N_6910);
nor U7510 (N_7510,N_6281,N_6196);
and U7511 (N_7511,N_6785,N_6759);
xnor U7512 (N_7512,N_6817,N_6385);
nand U7513 (N_7513,N_6083,N_6928);
nor U7514 (N_7514,N_6631,N_6461);
nand U7515 (N_7515,N_6091,N_6306);
or U7516 (N_7516,N_6079,N_7127);
nand U7517 (N_7517,N_6637,N_7188);
nor U7518 (N_7518,N_6265,N_6560);
nand U7519 (N_7519,N_6402,N_6649);
or U7520 (N_7520,N_6786,N_6665);
or U7521 (N_7521,N_6416,N_6200);
or U7522 (N_7522,N_6076,N_6464);
or U7523 (N_7523,N_6674,N_6594);
xnor U7524 (N_7524,N_6030,N_7079);
nor U7525 (N_7525,N_6290,N_6170);
nor U7526 (N_7526,N_6547,N_6298);
and U7527 (N_7527,N_6570,N_6829);
nand U7528 (N_7528,N_7061,N_6908);
nor U7529 (N_7529,N_6896,N_6146);
or U7530 (N_7530,N_6177,N_6858);
nand U7531 (N_7531,N_6340,N_6575);
nand U7532 (N_7532,N_6673,N_6772);
and U7533 (N_7533,N_7117,N_7049);
and U7534 (N_7534,N_6774,N_7031);
and U7535 (N_7535,N_7147,N_6922);
and U7536 (N_7536,N_6807,N_6215);
or U7537 (N_7537,N_6088,N_6938);
nor U7538 (N_7538,N_6816,N_6690);
nor U7539 (N_7539,N_6046,N_6502);
nand U7540 (N_7540,N_7138,N_6583);
nor U7541 (N_7541,N_6297,N_6657);
and U7542 (N_7542,N_6346,N_6993);
nand U7543 (N_7543,N_7155,N_6904);
nand U7544 (N_7544,N_6164,N_6433);
or U7545 (N_7545,N_6964,N_7005);
nand U7546 (N_7546,N_6021,N_6859);
nor U7547 (N_7547,N_6655,N_7116);
xnor U7548 (N_7548,N_7015,N_7165);
nand U7549 (N_7549,N_6084,N_6266);
xnor U7550 (N_7550,N_6912,N_6834);
xnor U7551 (N_7551,N_6457,N_6542);
xnor U7552 (N_7552,N_6443,N_6324);
nand U7553 (N_7553,N_6828,N_7054);
nor U7554 (N_7554,N_6158,N_7135);
nor U7555 (N_7555,N_6973,N_6867);
or U7556 (N_7556,N_6387,N_6380);
and U7557 (N_7557,N_6946,N_6877);
nand U7558 (N_7558,N_7195,N_6564);
nor U7559 (N_7559,N_7106,N_6627);
nand U7560 (N_7560,N_6153,N_6812);
and U7561 (N_7561,N_6721,N_6052);
nand U7562 (N_7562,N_6729,N_6349);
nor U7563 (N_7563,N_6459,N_7123);
or U7564 (N_7564,N_7111,N_6064);
xnor U7565 (N_7565,N_6855,N_7083);
nand U7566 (N_7566,N_6454,N_6159);
xor U7567 (N_7567,N_6765,N_6028);
and U7568 (N_7568,N_6754,N_6059);
and U7569 (N_7569,N_6209,N_6424);
nor U7570 (N_7570,N_6544,N_6907);
nor U7571 (N_7571,N_6227,N_6499);
or U7572 (N_7572,N_6201,N_6470);
nand U7573 (N_7573,N_6293,N_6442);
or U7574 (N_7574,N_6350,N_6991);
nand U7575 (N_7575,N_6490,N_6554);
xor U7576 (N_7576,N_7180,N_6808);
xnor U7577 (N_7577,N_6451,N_6216);
xnor U7578 (N_7578,N_6883,N_6533);
and U7579 (N_7579,N_7080,N_6417);
nand U7580 (N_7580,N_6971,N_6318);
xnor U7581 (N_7581,N_6050,N_7191);
nand U7582 (N_7582,N_6556,N_7001);
xor U7583 (N_7583,N_6066,N_6781);
and U7584 (N_7584,N_6719,N_6525);
nor U7585 (N_7585,N_7051,N_6675);
and U7586 (N_7586,N_6017,N_6397);
nor U7587 (N_7587,N_6685,N_6789);
xor U7588 (N_7588,N_6558,N_6471);
xnor U7589 (N_7589,N_6019,N_6681);
or U7590 (N_7590,N_6936,N_7048);
nor U7591 (N_7591,N_6331,N_6668);
and U7592 (N_7592,N_7108,N_6873);
and U7593 (N_7593,N_6016,N_6348);
and U7594 (N_7594,N_6057,N_6379);
and U7595 (N_7595,N_6047,N_7019);
or U7596 (N_7596,N_6722,N_6531);
and U7597 (N_7597,N_6413,N_7115);
xnor U7598 (N_7598,N_6184,N_6639);
xor U7599 (N_7599,N_7181,N_6020);
or U7600 (N_7600,N_6137,N_7161);
nand U7601 (N_7601,N_7185,N_6393);
nand U7602 (N_7602,N_6429,N_6510);
or U7603 (N_7603,N_7118,N_6445);
or U7604 (N_7604,N_7062,N_6043);
or U7605 (N_7605,N_6222,N_6909);
and U7606 (N_7606,N_6723,N_6820);
nand U7607 (N_7607,N_6519,N_6054);
nand U7608 (N_7608,N_6299,N_6513);
and U7609 (N_7609,N_6032,N_7182);
and U7610 (N_7610,N_6289,N_6523);
xor U7611 (N_7611,N_6903,N_6568);
nand U7612 (N_7612,N_6844,N_6487);
nor U7613 (N_7613,N_6205,N_6314);
xnor U7614 (N_7614,N_7097,N_6498);
nand U7615 (N_7615,N_6018,N_6426);
and U7616 (N_7616,N_6783,N_6526);
nand U7617 (N_7617,N_6240,N_6822);
nor U7618 (N_7618,N_6606,N_6339);
and U7619 (N_7619,N_6246,N_6269);
and U7620 (N_7620,N_6562,N_6010);
nand U7621 (N_7621,N_7046,N_6491);
xor U7622 (N_7622,N_6270,N_7192);
xor U7623 (N_7623,N_7136,N_7007);
or U7624 (N_7624,N_6932,N_6630);
nor U7625 (N_7625,N_6652,N_6740);
xnor U7626 (N_7626,N_6448,N_7096);
and U7627 (N_7627,N_6803,N_6351);
nor U7628 (N_7628,N_7059,N_7065);
nand U7629 (N_7629,N_6398,N_6539);
xnor U7630 (N_7630,N_6207,N_7018);
xnor U7631 (N_7631,N_6628,N_6458);
nand U7632 (N_7632,N_6378,N_6736);
nor U7633 (N_7633,N_7102,N_6623);
xnor U7634 (N_7634,N_6732,N_6347);
and U7635 (N_7635,N_6635,N_7173);
and U7636 (N_7636,N_6824,N_6825);
xnor U7637 (N_7637,N_6734,N_6743);
nand U7638 (N_7638,N_6275,N_6646);
xnor U7639 (N_7639,N_6590,N_6947);
or U7640 (N_7640,N_6862,N_6849);
or U7641 (N_7641,N_6831,N_6697);
and U7642 (N_7642,N_6950,N_7197);
xnor U7643 (N_7643,N_6230,N_6420);
nor U7644 (N_7644,N_6601,N_6323);
or U7645 (N_7645,N_7092,N_6818);
nand U7646 (N_7646,N_6480,N_6977);
and U7647 (N_7647,N_6257,N_6745);
xnor U7648 (N_7648,N_6770,N_6157);
nor U7649 (N_7649,N_6761,N_6410);
nand U7650 (N_7650,N_6121,N_6559);
and U7651 (N_7651,N_6984,N_6006);
and U7652 (N_7652,N_6097,N_7101);
nand U7653 (N_7653,N_6437,N_7055);
nand U7654 (N_7654,N_6990,N_6706);
nand U7655 (N_7655,N_7113,N_6660);
and U7656 (N_7656,N_6414,N_6371);
or U7657 (N_7657,N_6566,N_6898);
or U7658 (N_7658,N_6171,N_7178);
or U7659 (N_7659,N_6929,N_6259);
nand U7660 (N_7660,N_7043,N_7057);
or U7661 (N_7661,N_7084,N_6707);
and U7662 (N_7662,N_6144,N_6272);
or U7663 (N_7663,N_6768,N_6766);
nor U7664 (N_7664,N_6089,N_6142);
nand U7665 (N_7665,N_6206,N_6355);
nand U7666 (N_7666,N_6961,N_6895);
nor U7667 (N_7667,N_6823,N_6107);
xnor U7668 (N_7668,N_6427,N_6055);
or U7669 (N_7669,N_7044,N_6165);
and U7670 (N_7670,N_6945,N_6332);
xnor U7671 (N_7671,N_7038,N_6851);
or U7672 (N_7672,N_6788,N_6309);
nor U7673 (N_7673,N_6077,N_6492);
and U7674 (N_7674,N_6756,N_6253);
nand U7675 (N_7675,N_6168,N_6935);
nand U7676 (N_7676,N_6038,N_6529);
or U7677 (N_7677,N_6002,N_6753);
nor U7678 (N_7678,N_7199,N_7186);
nand U7679 (N_7679,N_6096,N_6180);
or U7680 (N_7680,N_6242,N_6684);
and U7681 (N_7681,N_7109,N_6802);
xor U7682 (N_7682,N_7148,N_6814);
xnor U7683 (N_7683,N_6011,N_6365);
and U7684 (N_7684,N_6555,N_6746);
nor U7685 (N_7685,N_6711,N_6647);
or U7686 (N_7686,N_7162,N_7070);
or U7687 (N_7687,N_6663,N_6321);
or U7688 (N_7688,N_6390,N_6261);
and U7689 (N_7689,N_6517,N_6784);
nor U7690 (N_7690,N_6953,N_6666);
or U7691 (N_7691,N_6679,N_6870);
nor U7692 (N_7692,N_6342,N_6208);
nand U7693 (N_7693,N_6839,N_7122);
nand U7694 (N_7694,N_6854,N_6805);
nand U7695 (N_7695,N_6915,N_6013);
nand U7696 (N_7696,N_6147,N_6400);
nor U7697 (N_7697,N_6821,N_6441);
or U7698 (N_7698,N_7193,N_6446);
or U7699 (N_7699,N_6888,N_6081);
xnor U7700 (N_7700,N_6462,N_6603);
xnor U7701 (N_7701,N_6591,N_6848);
and U7702 (N_7702,N_6727,N_6656);
xnor U7703 (N_7703,N_7041,N_6235);
nor U7704 (N_7704,N_7141,N_6494);
nand U7705 (N_7705,N_6217,N_6710);
and U7706 (N_7706,N_6056,N_6012);
and U7707 (N_7707,N_6176,N_6356);
nor U7708 (N_7708,N_6074,N_6431);
nor U7709 (N_7709,N_7024,N_6231);
nand U7710 (N_7710,N_7124,N_7029);
xor U7711 (N_7711,N_6728,N_6291);
or U7712 (N_7712,N_7032,N_6101);
and U7713 (N_7713,N_7036,N_6149);
and U7714 (N_7714,N_6304,N_6543);
or U7715 (N_7715,N_6109,N_6316);
or U7716 (N_7716,N_6255,N_6506);
and U7717 (N_7717,N_6546,N_6383);
or U7718 (N_7718,N_6956,N_6632);
and U7719 (N_7719,N_6582,N_6826);
or U7720 (N_7720,N_7076,N_6388);
nand U7721 (N_7721,N_6127,N_6466);
nand U7722 (N_7722,N_7139,N_6965);
nor U7723 (N_7723,N_6061,N_6574);
and U7724 (N_7724,N_6193,N_7107);
nand U7725 (N_7725,N_6864,N_6108);
or U7726 (N_7726,N_6511,N_6411);
and U7727 (N_7727,N_6368,N_6189);
nor U7728 (N_7728,N_6641,N_6182);
nand U7729 (N_7729,N_6455,N_6771);
nor U7730 (N_7730,N_6214,N_6567);
nand U7731 (N_7731,N_7086,N_6972);
xnor U7732 (N_7732,N_6504,N_6004);
nor U7733 (N_7733,N_7163,N_6284);
and U7734 (N_7734,N_6330,N_6008);
nor U7735 (N_7735,N_6484,N_7016);
nand U7736 (N_7736,N_6980,N_6228);
and U7737 (N_7737,N_6592,N_6156);
nor U7738 (N_7738,N_7146,N_6460);
xor U7739 (N_7739,N_6022,N_6087);
and U7740 (N_7740,N_6687,N_6248);
or U7741 (N_7741,N_6951,N_6911);
nor U7742 (N_7742,N_7169,N_6092);
nor U7743 (N_7743,N_6033,N_6958);
or U7744 (N_7744,N_6181,N_7077);
xor U7745 (N_7745,N_6369,N_6527);
nand U7746 (N_7746,N_6738,N_6051);
nand U7747 (N_7747,N_6689,N_6833);
xnor U7748 (N_7748,N_6880,N_6326);
nand U7749 (N_7749,N_7068,N_6354);
or U7750 (N_7750,N_6757,N_7172);
nand U7751 (N_7751,N_6188,N_6247);
and U7752 (N_7752,N_6174,N_6377);
xnor U7753 (N_7753,N_6421,N_6620);
nor U7754 (N_7754,N_6692,N_6651);
nand U7755 (N_7755,N_6267,N_6882);
or U7756 (N_7756,N_6169,N_7027);
or U7757 (N_7757,N_7152,N_6602);
nor U7758 (N_7758,N_6712,N_6027);
or U7759 (N_7759,N_6060,N_6203);
xor U7760 (N_7760,N_6600,N_6115);
and U7761 (N_7761,N_6758,N_7023);
and U7762 (N_7762,N_7060,N_6902);
nand U7763 (N_7763,N_6262,N_7002);
nor U7764 (N_7764,N_6287,N_6890);
xor U7765 (N_7765,N_6197,N_6726);
nor U7766 (N_7766,N_6031,N_6418);
nor U7767 (N_7767,N_6604,N_6939);
or U7768 (N_7768,N_6920,N_6015);
and U7769 (N_7769,N_6260,N_6313);
nor U7770 (N_7770,N_7144,N_6173);
nor U7771 (N_7771,N_6286,N_6406);
nand U7772 (N_7772,N_6241,N_6633);
nor U7773 (N_7773,N_7090,N_6220);
xnor U7774 (N_7774,N_6106,N_6962);
xor U7775 (N_7775,N_6522,N_6243);
xor U7776 (N_7776,N_6327,N_6881);
nor U7777 (N_7777,N_6252,N_6918);
nand U7778 (N_7778,N_6062,N_6989);
or U7779 (N_7779,N_6897,N_6676);
and U7780 (N_7780,N_6449,N_7184);
or U7781 (N_7781,N_6000,N_6638);
nor U7782 (N_7782,N_7150,N_6642);
and U7783 (N_7783,N_6131,N_6394);
nand U7784 (N_7784,N_6917,N_6810);
nand U7785 (N_7785,N_7196,N_6415);
nand U7786 (N_7786,N_6315,N_6237);
xor U7787 (N_7787,N_7039,N_6232);
and U7788 (N_7788,N_6901,N_6987);
nor U7789 (N_7789,N_6996,N_6609);
nand U7790 (N_7790,N_6213,N_6532);
nor U7791 (N_7791,N_6311,N_6596);
nor U7792 (N_7792,N_6536,N_6952);
xnor U7793 (N_7793,N_6507,N_6198);
or U7794 (N_7794,N_6978,N_7093);
and U7795 (N_7795,N_6271,N_6278);
or U7796 (N_7796,N_6528,N_6034);
xor U7797 (N_7797,N_7103,N_6967);
xnor U7798 (N_7798,N_6495,N_6221);
nand U7799 (N_7799,N_6515,N_6381);
or U7800 (N_7800,N_6829,N_6449);
nand U7801 (N_7801,N_6824,N_6331);
xor U7802 (N_7802,N_6772,N_6459);
or U7803 (N_7803,N_6048,N_6532);
or U7804 (N_7804,N_6001,N_6089);
nor U7805 (N_7805,N_6690,N_6870);
xor U7806 (N_7806,N_6810,N_6538);
or U7807 (N_7807,N_6488,N_7182);
and U7808 (N_7808,N_6319,N_7146);
and U7809 (N_7809,N_6925,N_6746);
xnor U7810 (N_7810,N_6693,N_6633);
nor U7811 (N_7811,N_6975,N_6115);
nor U7812 (N_7812,N_6024,N_6341);
xor U7813 (N_7813,N_6963,N_6281);
nand U7814 (N_7814,N_6344,N_6934);
nand U7815 (N_7815,N_6254,N_6751);
nand U7816 (N_7816,N_6202,N_6702);
and U7817 (N_7817,N_6226,N_6584);
nor U7818 (N_7818,N_7167,N_6777);
or U7819 (N_7819,N_6801,N_6099);
xor U7820 (N_7820,N_6428,N_6536);
and U7821 (N_7821,N_6248,N_6775);
or U7822 (N_7822,N_6700,N_6569);
and U7823 (N_7823,N_6676,N_6918);
or U7824 (N_7824,N_6485,N_6494);
and U7825 (N_7825,N_6386,N_7081);
nor U7826 (N_7826,N_6456,N_6991);
xnor U7827 (N_7827,N_6158,N_6751);
nand U7828 (N_7828,N_6355,N_6724);
and U7829 (N_7829,N_6890,N_6594);
nor U7830 (N_7830,N_7112,N_6737);
xnor U7831 (N_7831,N_6474,N_6591);
and U7832 (N_7832,N_6633,N_6991);
nand U7833 (N_7833,N_6046,N_7072);
nor U7834 (N_7834,N_6122,N_6425);
xnor U7835 (N_7835,N_6728,N_6065);
nand U7836 (N_7836,N_6964,N_6050);
xor U7837 (N_7837,N_6071,N_6997);
nand U7838 (N_7838,N_7004,N_7008);
nor U7839 (N_7839,N_6675,N_6471);
or U7840 (N_7840,N_7068,N_7199);
or U7841 (N_7841,N_6293,N_7083);
or U7842 (N_7842,N_6292,N_6763);
or U7843 (N_7843,N_7169,N_6392);
and U7844 (N_7844,N_6002,N_6817);
nor U7845 (N_7845,N_7006,N_6776);
nor U7846 (N_7846,N_6764,N_7072);
and U7847 (N_7847,N_6184,N_6263);
nor U7848 (N_7848,N_6417,N_6895);
and U7849 (N_7849,N_7063,N_6169);
and U7850 (N_7850,N_6018,N_6162);
or U7851 (N_7851,N_6252,N_6186);
and U7852 (N_7852,N_6693,N_7039);
or U7853 (N_7853,N_6352,N_6827);
nand U7854 (N_7854,N_6188,N_6422);
and U7855 (N_7855,N_6155,N_6814);
xor U7856 (N_7856,N_6984,N_6315);
xnor U7857 (N_7857,N_6727,N_6068);
nor U7858 (N_7858,N_6690,N_6101);
and U7859 (N_7859,N_7093,N_6605);
nor U7860 (N_7860,N_6321,N_6757);
nand U7861 (N_7861,N_7147,N_7153);
or U7862 (N_7862,N_7163,N_6799);
xnor U7863 (N_7863,N_6451,N_6655);
nor U7864 (N_7864,N_6782,N_6896);
nor U7865 (N_7865,N_6491,N_6587);
and U7866 (N_7866,N_6439,N_6567);
or U7867 (N_7867,N_6815,N_6994);
nand U7868 (N_7868,N_6497,N_6115);
or U7869 (N_7869,N_6227,N_6645);
or U7870 (N_7870,N_6990,N_6118);
or U7871 (N_7871,N_6131,N_6823);
and U7872 (N_7872,N_6916,N_6045);
nor U7873 (N_7873,N_6800,N_7087);
or U7874 (N_7874,N_7090,N_6991);
xnor U7875 (N_7875,N_7064,N_7117);
xor U7876 (N_7876,N_6394,N_7113);
xor U7877 (N_7877,N_6036,N_7160);
and U7878 (N_7878,N_6972,N_6040);
xor U7879 (N_7879,N_6305,N_6445);
xnor U7880 (N_7880,N_6299,N_7084);
xnor U7881 (N_7881,N_7060,N_6822);
nand U7882 (N_7882,N_6830,N_6899);
nor U7883 (N_7883,N_7047,N_7097);
nand U7884 (N_7884,N_6472,N_6703);
xor U7885 (N_7885,N_7000,N_7183);
nor U7886 (N_7886,N_6620,N_6653);
or U7887 (N_7887,N_6499,N_6004);
nand U7888 (N_7888,N_6300,N_6374);
nand U7889 (N_7889,N_7070,N_6087);
nand U7890 (N_7890,N_6440,N_6942);
or U7891 (N_7891,N_6603,N_6449);
or U7892 (N_7892,N_6532,N_6999);
or U7893 (N_7893,N_6695,N_6377);
or U7894 (N_7894,N_6883,N_6632);
and U7895 (N_7895,N_6627,N_6073);
or U7896 (N_7896,N_6523,N_7122);
or U7897 (N_7897,N_6230,N_6441);
and U7898 (N_7898,N_6316,N_6599);
xor U7899 (N_7899,N_6038,N_7102);
nand U7900 (N_7900,N_7159,N_6938);
and U7901 (N_7901,N_7117,N_6989);
and U7902 (N_7902,N_6921,N_6496);
nand U7903 (N_7903,N_6385,N_6697);
xnor U7904 (N_7904,N_6318,N_6005);
nor U7905 (N_7905,N_6939,N_6242);
or U7906 (N_7906,N_7025,N_6646);
and U7907 (N_7907,N_6344,N_6512);
and U7908 (N_7908,N_6495,N_6583);
and U7909 (N_7909,N_6715,N_6175);
and U7910 (N_7910,N_6318,N_6648);
nand U7911 (N_7911,N_7161,N_6706);
and U7912 (N_7912,N_7106,N_6360);
or U7913 (N_7913,N_6673,N_6549);
or U7914 (N_7914,N_6353,N_6890);
nand U7915 (N_7915,N_6461,N_6746);
and U7916 (N_7916,N_6730,N_6560);
or U7917 (N_7917,N_6375,N_7094);
nor U7918 (N_7918,N_7103,N_6365);
nand U7919 (N_7919,N_6316,N_6290);
xor U7920 (N_7920,N_6152,N_6048);
nand U7921 (N_7921,N_6060,N_7168);
nor U7922 (N_7922,N_6388,N_6189);
or U7923 (N_7923,N_6148,N_6782);
nor U7924 (N_7924,N_6446,N_6148);
or U7925 (N_7925,N_6021,N_6754);
nor U7926 (N_7926,N_6703,N_6576);
or U7927 (N_7927,N_7062,N_6636);
or U7928 (N_7928,N_6366,N_6955);
nand U7929 (N_7929,N_6872,N_6648);
and U7930 (N_7930,N_7057,N_6689);
xnor U7931 (N_7931,N_6698,N_6227);
or U7932 (N_7932,N_6183,N_6389);
and U7933 (N_7933,N_6131,N_6596);
or U7934 (N_7934,N_6445,N_6783);
or U7935 (N_7935,N_6624,N_6830);
xor U7936 (N_7936,N_6267,N_6839);
nor U7937 (N_7937,N_7196,N_6447);
and U7938 (N_7938,N_6314,N_7103);
nand U7939 (N_7939,N_6663,N_6212);
nand U7940 (N_7940,N_7012,N_6208);
nor U7941 (N_7941,N_6803,N_6279);
xnor U7942 (N_7942,N_6143,N_6993);
nor U7943 (N_7943,N_7178,N_7054);
nor U7944 (N_7944,N_6760,N_6232);
and U7945 (N_7945,N_6215,N_6727);
nor U7946 (N_7946,N_6280,N_6372);
and U7947 (N_7947,N_6422,N_6133);
nand U7948 (N_7948,N_6646,N_7072);
xor U7949 (N_7949,N_6388,N_7031);
nand U7950 (N_7950,N_7002,N_6309);
nand U7951 (N_7951,N_6878,N_6717);
nor U7952 (N_7952,N_6517,N_6566);
and U7953 (N_7953,N_7197,N_6172);
and U7954 (N_7954,N_6661,N_6647);
nand U7955 (N_7955,N_6471,N_6588);
nor U7956 (N_7956,N_7007,N_6585);
nand U7957 (N_7957,N_7077,N_6937);
nand U7958 (N_7958,N_6215,N_6024);
xnor U7959 (N_7959,N_6135,N_6076);
or U7960 (N_7960,N_6436,N_6777);
or U7961 (N_7961,N_6354,N_6644);
nor U7962 (N_7962,N_6541,N_6221);
nor U7963 (N_7963,N_6384,N_6236);
nor U7964 (N_7964,N_6616,N_6515);
nor U7965 (N_7965,N_7105,N_6447);
and U7966 (N_7966,N_6445,N_6397);
or U7967 (N_7967,N_6825,N_6873);
nand U7968 (N_7968,N_6244,N_6526);
nand U7969 (N_7969,N_7119,N_6961);
nand U7970 (N_7970,N_6669,N_6082);
and U7971 (N_7971,N_6027,N_6011);
nor U7972 (N_7972,N_6043,N_6138);
xor U7973 (N_7973,N_6797,N_6595);
xor U7974 (N_7974,N_6724,N_6653);
xor U7975 (N_7975,N_6756,N_6684);
nand U7976 (N_7976,N_6512,N_6026);
xnor U7977 (N_7977,N_6319,N_6045);
or U7978 (N_7978,N_6023,N_6304);
xnor U7979 (N_7979,N_6700,N_6742);
xor U7980 (N_7980,N_6670,N_6072);
xor U7981 (N_7981,N_6687,N_6464);
and U7982 (N_7982,N_7126,N_6997);
or U7983 (N_7983,N_6691,N_6287);
xor U7984 (N_7984,N_6175,N_6258);
nand U7985 (N_7985,N_6652,N_7152);
xor U7986 (N_7986,N_6508,N_6563);
nand U7987 (N_7987,N_6652,N_6165);
xnor U7988 (N_7988,N_6314,N_6384);
or U7989 (N_7989,N_6424,N_6579);
nor U7990 (N_7990,N_6934,N_6360);
nand U7991 (N_7991,N_6302,N_6724);
and U7992 (N_7992,N_6646,N_6013);
and U7993 (N_7993,N_6457,N_7198);
xor U7994 (N_7994,N_6746,N_6634);
xnor U7995 (N_7995,N_6693,N_6097);
xor U7996 (N_7996,N_6081,N_6499);
nor U7997 (N_7997,N_7079,N_7057);
xor U7998 (N_7998,N_7061,N_6218);
nand U7999 (N_7999,N_7095,N_6135);
nor U8000 (N_8000,N_6949,N_7115);
nand U8001 (N_8001,N_6795,N_6588);
nand U8002 (N_8002,N_6294,N_6827);
nand U8003 (N_8003,N_6678,N_7180);
or U8004 (N_8004,N_6599,N_6378);
or U8005 (N_8005,N_6466,N_6727);
nor U8006 (N_8006,N_6380,N_7031);
or U8007 (N_8007,N_6200,N_6410);
xor U8008 (N_8008,N_6245,N_6513);
and U8009 (N_8009,N_6808,N_6315);
or U8010 (N_8010,N_6735,N_6670);
nand U8011 (N_8011,N_7027,N_6545);
xor U8012 (N_8012,N_6612,N_6802);
nand U8013 (N_8013,N_6850,N_6857);
or U8014 (N_8014,N_6617,N_7076);
xor U8015 (N_8015,N_6488,N_7135);
nor U8016 (N_8016,N_6032,N_6224);
nand U8017 (N_8017,N_6571,N_6887);
nand U8018 (N_8018,N_6907,N_6441);
or U8019 (N_8019,N_6178,N_6427);
or U8020 (N_8020,N_6663,N_6449);
or U8021 (N_8021,N_6542,N_7096);
or U8022 (N_8022,N_6966,N_7189);
xor U8023 (N_8023,N_6786,N_6094);
and U8024 (N_8024,N_6395,N_6662);
or U8025 (N_8025,N_6102,N_6326);
and U8026 (N_8026,N_6555,N_6161);
nand U8027 (N_8027,N_6645,N_6408);
xnor U8028 (N_8028,N_6262,N_6086);
nand U8029 (N_8029,N_7158,N_6628);
or U8030 (N_8030,N_6733,N_6710);
and U8031 (N_8031,N_6177,N_6212);
nand U8032 (N_8032,N_6491,N_6046);
nand U8033 (N_8033,N_6112,N_6146);
xor U8034 (N_8034,N_6511,N_6728);
nor U8035 (N_8035,N_6361,N_6271);
nand U8036 (N_8036,N_6974,N_6756);
xnor U8037 (N_8037,N_7087,N_6593);
nor U8038 (N_8038,N_6527,N_6107);
or U8039 (N_8039,N_6622,N_7175);
xnor U8040 (N_8040,N_6491,N_6771);
or U8041 (N_8041,N_6525,N_6240);
nor U8042 (N_8042,N_6298,N_6728);
xor U8043 (N_8043,N_6344,N_7162);
nand U8044 (N_8044,N_6488,N_6761);
and U8045 (N_8045,N_6433,N_6306);
xor U8046 (N_8046,N_6293,N_7184);
nand U8047 (N_8047,N_6529,N_6081);
nor U8048 (N_8048,N_6879,N_6146);
and U8049 (N_8049,N_7154,N_6003);
xor U8050 (N_8050,N_6404,N_6809);
nand U8051 (N_8051,N_7129,N_6852);
or U8052 (N_8052,N_6185,N_6437);
nor U8053 (N_8053,N_6691,N_6701);
nand U8054 (N_8054,N_6099,N_6906);
nor U8055 (N_8055,N_6308,N_6751);
or U8056 (N_8056,N_7163,N_7023);
and U8057 (N_8057,N_6229,N_6376);
nor U8058 (N_8058,N_6443,N_6823);
nor U8059 (N_8059,N_6452,N_6477);
and U8060 (N_8060,N_6679,N_6451);
xnor U8061 (N_8061,N_6527,N_6472);
xnor U8062 (N_8062,N_6437,N_6984);
or U8063 (N_8063,N_6693,N_6474);
and U8064 (N_8064,N_6293,N_6324);
nand U8065 (N_8065,N_6083,N_7182);
and U8066 (N_8066,N_6298,N_6327);
or U8067 (N_8067,N_6512,N_6575);
nor U8068 (N_8068,N_6730,N_6281);
nor U8069 (N_8069,N_6001,N_6529);
xor U8070 (N_8070,N_6213,N_7168);
or U8071 (N_8071,N_6402,N_6250);
xor U8072 (N_8072,N_6476,N_6892);
or U8073 (N_8073,N_7154,N_6883);
and U8074 (N_8074,N_6080,N_6853);
xnor U8075 (N_8075,N_6017,N_6209);
nor U8076 (N_8076,N_7082,N_6165);
nand U8077 (N_8077,N_7106,N_6460);
nor U8078 (N_8078,N_6477,N_6618);
nor U8079 (N_8079,N_6499,N_6412);
xnor U8080 (N_8080,N_6379,N_6735);
xor U8081 (N_8081,N_6834,N_6007);
xor U8082 (N_8082,N_6587,N_6200);
xnor U8083 (N_8083,N_6821,N_6203);
xor U8084 (N_8084,N_6357,N_7105);
or U8085 (N_8085,N_6500,N_6501);
nor U8086 (N_8086,N_6589,N_6367);
nand U8087 (N_8087,N_6836,N_6043);
and U8088 (N_8088,N_6410,N_7154);
nand U8089 (N_8089,N_6618,N_6144);
nor U8090 (N_8090,N_7072,N_6047);
nor U8091 (N_8091,N_6419,N_7190);
and U8092 (N_8092,N_6786,N_6670);
or U8093 (N_8093,N_6015,N_6445);
and U8094 (N_8094,N_6484,N_7060);
nand U8095 (N_8095,N_6152,N_6309);
or U8096 (N_8096,N_6926,N_6100);
xnor U8097 (N_8097,N_6129,N_6507);
or U8098 (N_8098,N_6612,N_6933);
xor U8099 (N_8099,N_6120,N_6660);
nand U8100 (N_8100,N_6651,N_6549);
xor U8101 (N_8101,N_6238,N_6027);
and U8102 (N_8102,N_6944,N_6827);
xor U8103 (N_8103,N_6617,N_6830);
nand U8104 (N_8104,N_6501,N_6958);
xnor U8105 (N_8105,N_6226,N_6402);
nor U8106 (N_8106,N_6347,N_6730);
or U8107 (N_8107,N_6851,N_6978);
xor U8108 (N_8108,N_7058,N_6073);
or U8109 (N_8109,N_6299,N_6212);
nand U8110 (N_8110,N_6131,N_7016);
or U8111 (N_8111,N_7104,N_6913);
and U8112 (N_8112,N_6409,N_6255);
xor U8113 (N_8113,N_6757,N_6750);
xor U8114 (N_8114,N_6695,N_6223);
nor U8115 (N_8115,N_6034,N_6986);
nand U8116 (N_8116,N_6671,N_6351);
xnor U8117 (N_8117,N_7036,N_6616);
or U8118 (N_8118,N_6144,N_7175);
and U8119 (N_8119,N_6726,N_7028);
nand U8120 (N_8120,N_7012,N_6346);
xor U8121 (N_8121,N_6395,N_7163);
nor U8122 (N_8122,N_6315,N_6032);
or U8123 (N_8123,N_7046,N_6125);
or U8124 (N_8124,N_6992,N_7077);
xnor U8125 (N_8125,N_7143,N_6988);
nand U8126 (N_8126,N_6136,N_6473);
or U8127 (N_8127,N_6262,N_6574);
xnor U8128 (N_8128,N_7151,N_6203);
nand U8129 (N_8129,N_7115,N_6323);
and U8130 (N_8130,N_6439,N_6642);
xor U8131 (N_8131,N_6785,N_6386);
nor U8132 (N_8132,N_6306,N_7039);
or U8133 (N_8133,N_7191,N_7067);
and U8134 (N_8134,N_7019,N_7084);
and U8135 (N_8135,N_6767,N_6303);
xnor U8136 (N_8136,N_6128,N_6648);
and U8137 (N_8137,N_6717,N_6933);
or U8138 (N_8138,N_7056,N_6930);
or U8139 (N_8139,N_6869,N_6633);
xor U8140 (N_8140,N_6895,N_6322);
and U8141 (N_8141,N_6482,N_6770);
or U8142 (N_8142,N_6857,N_6189);
nor U8143 (N_8143,N_7001,N_6630);
nor U8144 (N_8144,N_6996,N_6075);
nand U8145 (N_8145,N_7175,N_6278);
nor U8146 (N_8146,N_6757,N_6985);
and U8147 (N_8147,N_6408,N_6804);
nor U8148 (N_8148,N_6063,N_6023);
xor U8149 (N_8149,N_6203,N_6377);
or U8150 (N_8150,N_7083,N_6845);
nor U8151 (N_8151,N_7081,N_7108);
nand U8152 (N_8152,N_6528,N_6683);
nand U8153 (N_8153,N_7099,N_6666);
or U8154 (N_8154,N_6658,N_6363);
xor U8155 (N_8155,N_6784,N_6629);
nand U8156 (N_8156,N_6072,N_6293);
nor U8157 (N_8157,N_7147,N_6109);
and U8158 (N_8158,N_6926,N_6467);
nor U8159 (N_8159,N_6141,N_6639);
or U8160 (N_8160,N_6631,N_6811);
nor U8161 (N_8161,N_6706,N_6487);
and U8162 (N_8162,N_6024,N_6711);
and U8163 (N_8163,N_6572,N_6791);
nor U8164 (N_8164,N_6984,N_6754);
or U8165 (N_8165,N_6628,N_7133);
or U8166 (N_8166,N_6610,N_6780);
nor U8167 (N_8167,N_6358,N_6307);
nand U8168 (N_8168,N_7025,N_6502);
nand U8169 (N_8169,N_6930,N_6960);
nor U8170 (N_8170,N_7044,N_6802);
or U8171 (N_8171,N_6001,N_6079);
or U8172 (N_8172,N_7160,N_6942);
xnor U8173 (N_8173,N_6309,N_6219);
xnor U8174 (N_8174,N_6416,N_6981);
and U8175 (N_8175,N_6583,N_6392);
and U8176 (N_8176,N_6250,N_6827);
nor U8177 (N_8177,N_6656,N_6730);
nand U8178 (N_8178,N_6641,N_6738);
nor U8179 (N_8179,N_6247,N_6797);
or U8180 (N_8180,N_6831,N_6158);
nor U8181 (N_8181,N_6824,N_6298);
or U8182 (N_8182,N_6998,N_6638);
xor U8183 (N_8183,N_6592,N_6568);
and U8184 (N_8184,N_6097,N_6202);
nand U8185 (N_8185,N_6131,N_6589);
nor U8186 (N_8186,N_7106,N_6006);
nand U8187 (N_8187,N_6388,N_6351);
and U8188 (N_8188,N_6917,N_6048);
or U8189 (N_8189,N_6093,N_6026);
nor U8190 (N_8190,N_6623,N_6163);
or U8191 (N_8191,N_6814,N_6870);
and U8192 (N_8192,N_6569,N_6315);
nand U8193 (N_8193,N_7054,N_6203);
and U8194 (N_8194,N_6200,N_7064);
and U8195 (N_8195,N_7194,N_6991);
or U8196 (N_8196,N_6677,N_6633);
or U8197 (N_8197,N_6695,N_6770);
or U8198 (N_8198,N_6062,N_7049);
or U8199 (N_8199,N_6987,N_6120);
and U8200 (N_8200,N_7157,N_6856);
nand U8201 (N_8201,N_6348,N_7164);
nand U8202 (N_8202,N_6668,N_6008);
nor U8203 (N_8203,N_6105,N_6604);
nand U8204 (N_8204,N_6843,N_6907);
nand U8205 (N_8205,N_6184,N_6947);
xnor U8206 (N_8206,N_6951,N_7182);
and U8207 (N_8207,N_6879,N_6575);
xnor U8208 (N_8208,N_6317,N_6308);
nand U8209 (N_8209,N_6158,N_6081);
or U8210 (N_8210,N_6386,N_6802);
or U8211 (N_8211,N_6749,N_6783);
and U8212 (N_8212,N_6789,N_6737);
or U8213 (N_8213,N_6128,N_6092);
xnor U8214 (N_8214,N_6681,N_6900);
and U8215 (N_8215,N_6615,N_7163);
xor U8216 (N_8216,N_6275,N_6360);
nor U8217 (N_8217,N_6947,N_7081);
nand U8218 (N_8218,N_6454,N_7050);
and U8219 (N_8219,N_6683,N_7180);
xnor U8220 (N_8220,N_6516,N_6267);
and U8221 (N_8221,N_7159,N_7087);
nor U8222 (N_8222,N_6723,N_6199);
xor U8223 (N_8223,N_6919,N_7103);
or U8224 (N_8224,N_7177,N_6617);
xnor U8225 (N_8225,N_6776,N_7147);
nor U8226 (N_8226,N_6221,N_6320);
nand U8227 (N_8227,N_6912,N_7171);
or U8228 (N_8228,N_6013,N_6412);
nand U8229 (N_8229,N_6354,N_6844);
nand U8230 (N_8230,N_6432,N_6476);
or U8231 (N_8231,N_6667,N_6549);
and U8232 (N_8232,N_7187,N_6904);
xnor U8233 (N_8233,N_6782,N_7137);
or U8234 (N_8234,N_6884,N_6622);
nand U8235 (N_8235,N_7154,N_6206);
nand U8236 (N_8236,N_7157,N_6863);
nor U8237 (N_8237,N_6834,N_6034);
and U8238 (N_8238,N_6498,N_6146);
and U8239 (N_8239,N_6152,N_6325);
nor U8240 (N_8240,N_7158,N_7008);
or U8241 (N_8241,N_6468,N_6795);
nor U8242 (N_8242,N_6443,N_6427);
xor U8243 (N_8243,N_6441,N_6687);
nor U8244 (N_8244,N_6023,N_7119);
nand U8245 (N_8245,N_6546,N_6766);
or U8246 (N_8246,N_7048,N_6175);
nor U8247 (N_8247,N_6124,N_6269);
and U8248 (N_8248,N_6764,N_6724);
xnor U8249 (N_8249,N_6982,N_6296);
or U8250 (N_8250,N_7179,N_6760);
and U8251 (N_8251,N_6697,N_6315);
nor U8252 (N_8252,N_6642,N_6132);
nor U8253 (N_8253,N_6836,N_6014);
or U8254 (N_8254,N_7056,N_6520);
or U8255 (N_8255,N_6716,N_6052);
nor U8256 (N_8256,N_6319,N_6558);
nor U8257 (N_8257,N_6854,N_6320);
or U8258 (N_8258,N_6383,N_6527);
or U8259 (N_8259,N_6441,N_6967);
and U8260 (N_8260,N_6111,N_6503);
and U8261 (N_8261,N_6440,N_6853);
nor U8262 (N_8262,N_6977,N_6165);
and U8263 (N_8263,N_6214,N_6270);
nor U8264 (N_8264,N_7023,N_6213);
or U8265 (N_8265,N_6881,N_6364);
nor U8266 (N_8266,N_7105,N_6049);
and U8267 (N_8267,N_6934,N_6849);
and U8268 (N_8268,N_6257,N_6688);
nand U8269 (N_8269,N_6651,N_7152);
nand U8270 (N_8270,N_7080,N_6151);
or U8271 (N_8271,N_6599,N_6213);
and U8272 (N_8272,N_6933,N_7057);
or U8273 (N_8273,N_6044,N_6185);
nand U8274 (N_8274,N_6416,N_6605);
nand U8275 (N_8275,N_6598,N_6335);
or U8276 (N_8276,N_6592,N_6967);
nor U8277 (N_8277,N_6202,N_6491);
or U8278 (N_8278,N_6697,N_6024);
or U8279 (N_8279,N_7096,N_6464);
and U8280 (N_8280,N_7034,N_6601);
nand U8281 (N_8281,N_6366,N_6229);
nand U8282 (N_8282,N_6975,N_7105);
nand U8283 (N_8283,N_6894,N_6937);
nor U8284 (N_8284,N_6985,N_6134);
and U8285 (N_8285,N_6270,N_7182);
nand U8286 (N_8286,N_7102,N_6406);
or U8287 (N_8287,N_6626,N_6351);
and U8288 (N_8288,N_7124,N_6471);
nor U8289 (N_8289,N_6630,N_6048);
nor U8290 (N_8290,N_7164,N_6160);
nand U8291 (N_8291,N_6067,N_6024);
nor U8292 (N_8292,N_6298,N_6702);
and U8293 (N_8293,N_6948,N_7013);
or U8294 (N_8294,N_6826,N_6078);
nand U8295 (N_8295,N_7082,N_6564);
and U8296 (N_8296,N_6060,N_6378);
xnor U8297 (N_8297,N_6853,N_6028);
nand U8298 (N_8298,N_6189,N_7064);
and U8299 (N_8299,N_6626,N_7197);
or U8300 (N_8300,N_6681,N_6767);
and U8301 (N_8301,N_7112,N_6076);
xnor U8302 (N_8302,N_6737,N_6933);
or U8303 (N_8303,N_6936,N_6381);
nand U8304 (N_8304,N_7158,N_6218);
or U8305 (N_8305,N_6686,N_7180);
nand U8306 (N_8306,N_6011,N_6807);
nand U8307 (N_8307,N_6503,N_6263);
and U8308 (N_8308,N_6880,N_6439);
nor U8309 (N_8309,N_6705,N_6142);
nand U8310 (N_8310,N_6945,N_7175);
nor U8311 (N_8311,N_6770,N_6947);
xor U8312 (N_8312,N_7111,N_6267);
nor U8313 (N_8313,N_6015,N_6155);
xor U8314 (N_8314,N_6957,N_6197);
or U8315 (N_8315,N_6658,N_6841);
nand U8316 (N_8316,N_6848,N_6821);
or U8317 (N_8317,N_6181,N_6951);
nand U8318 (N_8318,N_6375,N_6280);
nor U8319 (N_8319,N_6241,N_6700);
xor U8320 (N_8320,N_6958,N_6305);
xor U8321 (N_8321,N_7032,N_6444);
or U8322 (N_8322,N_6603,N_7087);
nor U8323 (N_8323,N_6094,N_6772);
nand U8324 (N_8324,N_6798,N_6579);
and U8325 (N_8325,N_6020,N_6627);
nor U8326 (N_8326,N_6327,N_6585);
or U8327 (N_8327,N_7137,N_6024);
or U8328 (N_8328,N_6810,N_6749);
nand U8329 (N_8329,N_6839,N_7044);
xor U8330 (N_8330,N_6284,N_6997);
nand U8331 (N_8331,N_6448,N_6237);
nor U8332 (N_8332,N_6249,N_7126);
or U8333 (N_8333,N_6703,N_6223);
nand U8334 (N_8334,N_6919,N_6940);
or U8335 (N_8335,N_6712,N_6362);
and U8336 (N_8336,N_6044,N_6293);
and U8337 (N_8337,N_6792,N_6410);
nand U8338 (N_8338,N_6834,N_6801);
xnor U8339 (N_8339,N_6699,N_6892);
nand U8340 (N_8340,N_6518,N_7040);
or U8341 (N_8341,N_6486,N_6053);
or U8342 (N_8342,N_7052,N_7120);
xnor U8343 (N_8343,N_6911,N_6662);
xor U8344 (N_8344,N_6317,N_6380);
xor U8345 (N_8345,N_6254,N_6683);
nand U8346 (N_8346,N_6820,N_6088);
xnor U8347 (N_8347,N_6301,N_6289);
or U8348 (N_8348,N_7136,N_6880);
xnor U8349 (N_8349,N_6526,N_6648);
nor U8350 (N_8350,N_6148,N_6759);
nor U8351 (N_8351,N_6257,N_6770);
nand U8352 (N_8352,N_6367,N_6097);
or U8353 (N_8353,N_6020,N_6788);
nor U8354 (N_8354,N_7134,N_6961);
nor U8355 (N_8355,N_7129,N_7085);
xor U8356 (N_8356,N_6853,N_6284);
xor U8357 (N_8357,N_6264,N_7071);
and U8358 (N_8358,N_7021,N_6452);
nand U8359 (N_8359,N_6790,N_6455);
or U8360 (N_8360,N_6782,N_6295);
nand U8361 (N_8361,N_6640,N_6271);
and U8362 (N_8362,N_6592,N_6395);
or U8363 (N_8363,N_7137,N_6769);
or U8364 (N_8364,N_6359,N_7089);
xor U8365 (N_8365,N_6558,N_6967);
xor U8366 (N_8366,N_6698,N_6773);
nor U8367 (N_8367,N_6113,N_6890);
or U8368 (N_8368,N_6223,N_7171);
and U8369 (N_8369,N_6860,N_7154);
nor U8370 (N_8370,N_6262,N_6385);
or U8371 (N_8371,N_6569,N_6316);
and U8372 (N_8372,N_6789,N_6181);
nand U8373 (N_8373,N_6305,N_6703);
or U8374 (N_8374,N_7142,N_6852);
and U8375 (N_8375,N_6872,N_6736);
and U8376 (N_8376,N_6743,N_6566);
and U8377 (N_8377,N_7062,N_6454);
xor U8378 (N_8378,N_7086,N_6788);
and U8379 (N_8379,N_6944,N_6357);
and U8380 (N_8380,N_7051,N_6849);
or U8381 (N_8381,N_6940,N_6011);
nor U8382 (N_8382,N_7194,N_7119);
nand U8383 (N_8383,N_6552,N_6412);
and U8384 (N_8384,N_6106,N_6644);
or U8385 (N_8385,N_7158,N_6116);
xor U8386 (N_8386,N_6298,N_6224);
and U8387 (N_8387,N_6698,N_6703);
nand U8388 (N_8388,N_6932,N_6283);
nor U8389 (N_8389,N_7140,N_6198);
or U8390 (N_8390,N_6089,N_6230);
nand U8391 (N_8391,N_7020,N_6614);
and U8392 (N_8392,N_6223,N_6430);
nor U8393 (N_8393,N_6898,N_6525);
and U8394 (N_8394,N_7134,N_6613);
nor U8395 (N_8395,N_6996,N_6946);
nand U8396 (N_8396,N_6113,N_6334);
nor U8397 (N_8397,N_7052,N_6334);
or U8398 (N_8398,N_6302,N_6360);
nor U8399 (N_8399,N_6917,N_7022);
nand U8400 (N_8400,N_7464,N_7586);
xor U8401 (N_8401,N_7515,N_7739);
nand U8402 (N_8402,N_8055,N_7822);
nor U8403 (N_8403,N_7745,N_8237);
nand U8404 (N_8404,N_7936,N_8296);
nand U8405 (N_8405,N_7396,N_7317);
and U8406 (N_8406,N_8252,N_7664);
nor U8407 (N_8407,N_7200,N_7565);
xnor U8408 (N_8408,N_8398,N_7212);
nand U8409 (N_8409,N_7452,N_7905);
nor U8410 (N_8410,N_8391,N_7696);
xnor U8411 (N_8411,N_8286,N_7342);
and U8412 (N_8412,N_7730,N_8281);
nand U8413 (N_8413,N_8021,N_8336);
or U8414 (N_8414,N_7714,N_8335);
nand U8415 (N_8415,N_8146,N_7559);
and U8416 (N_8416,N_7793,N_7271);
and U8417 (N_8417,N_7891,N_7475);
or U8418 (N_8418,N_7695,N_7362);
or U8419 (N_8419,N_7201,N_8151);
xor U8420 (N_8420,N_7859,N_7879);
and U8421 (N_8421,N_7647,N_8191);
and U8422 (N_8422,N_8388,N_7335);
nand U8423 (N_8423,N_7848,N_8042);
or U8424 (N_8424,N_8187,N_8179);
nand U8425 (N_8425,N_7389,N_7371);
and U8426 (N_8426,N_7492,N_7959);
xnor U8427 (N_8427,N_7281,N_7689);
and U8428 (N_8428,N_7743,N_8135);
nor U8429 (N_8429,N_7736,N_8376);
nor U8430 (N_8430,N_7645,N_7336);
and U8431 (N_8431,N_7938,N_7811);
and U8432 (N_8432,N_7868,N_7272);
or U8433 (N_8433,N_7843,N_8069);
and U8434 (N_8434,N_7478,N_8190);
nor U8435 (N_8435,N_8166,N_8355);
or U8436 (N_8436,N_7309,N_7930);
and U8437 (N_8437,N_7680,N_7874);
and U8438 (N_8438,N_7289,N_8087);
or U8439 (N_8439,N_7704,N_7882);
or U8440 (N_8440,N_7635,N_7778);
xor U8441 (N_8441,N_7679,N_7451);
nand U8442 (N_8442,N_8383,N_8071);
nor U8443 (N_8443,N_7410,N_7668);
nand U8444 (N_8444,N_8368,N_7246);
or U8445 (N_8445,N_7324,N_8299);
nand U8446 (N_8446,N_7477,N_7249);
xnor U8447 (N_8447,N_8082,N_7998);
xnor U8448 (N_8448,N_7211,N_7983);
or U8449 (N_8449,N_7278,N_8291);
or U8450 (N_8450,N_8352,N_7250);
nand U8451 (N_8451,N_8210,N_7306);
and U8452 (N_8452,N_8140,N_8269);
and U8453 (N_8453,N_8095,N_8310);
xor U8454 (N_8454,N_7571,N_7513);
nor U8455 (N_8455,N_7481,N_8288);
and U8456 (N_8456,N_8364,N_7840);
or U8457 (N_8457,N_7919,N_7523);
or U8458 (N_8458,N_7528,N_7267);
and U8459 (N_8459,N_7213,N_7230);
xor U8460 (N_8460,N_7671,N_7996);
nor U8461 (N_8461,N_7821,N_8350);
and U8462 (N_8462,N_7673,N_7297);
nor U8463 (N_8463,N_7881,N_7514);
xnor U8464 (N_8464,N_7439,N_7404);
or U8465 (N_8465,N_7277,N_7502);
and U8466 (N_8466,N_8211,N_7982);
or U8467 (N_8467,N_7588,N_7912);
and U8468 (N_8468,N_8092,N_7691);
nand U8469 (N_8469,N_8287,N_7248);
nor U8470 (N_8470,N_8363,N_7659);
nor U8471 (N_8471,N_7901,N_7628);
nand U8472 (N_8472,N_7416,N_7710);
nor U8473 (N_8473,N_7366,N_7665);
or U8474 (N_8474,N_7796,N_7622);
and U8475 (N_8475,N_7214,N_7290);
or U8476 (N_8476,N_7826,N_7794);
xor U8477 (N_8477,N_8107,N_8349);
nand U8478 (N_8478,N_7705,N_7786);
xor U8479 (N_8479,N_8038,N_7910);
and U8480 (N_8480,N_8386,N_7238);
xnor U8481 (N_8481,N_7991,N_7471);
xnor U8482 (N_8482,N_7886,N_7259);
nor U8483 (N_8483,N_7470,N_7841);
nand U8484 (N_8484,N_7803,N_8147);
nor U8485 (N_8485,N_7862,N_7429);
or U8486 (N_8486,N_7880,N_7781);
and U8487 (N_8487,N_7694,N_7724);
xor U8488 (N_8488,N_7600,N_8058);
nor U8489 (N_8489,N_7906,N_7999);
and U8490 (N_8490,N_7964,N_7631);
or U8491 (N_8491,N_7707,N_8195);
nor U8492 (N_8492,N_7712,N_8235);
nor U8493 (N_8493,N_8198,N_7591);
xor U8494 (N_8494,N_8102,N_7207);
or U8495 (N_8495,N_7677,N_7374);
nand U8496 (N_8496,N_8158,N_7800);
nand U8497 (N_8497,N_8157,N_7735);
nand U8498 (N_8498,N_7785,N_7792);
nand U8499 (N_8499,N_8262,N_8257);
and U8500 (N_8500,N_7825,N_7334);
nand U8501 (N_8501,N_8313,N_7675);
xor U8502 (N_8502,N_8277,N_7723);
xor U8503 (N_8503,N_7969,N_7392);
xor U8504 (N_8504,N_7526,N_7564);
xor U8505 (N_8505,N_8337,N_8251);
xnor U8506 (N_8506,N_7529,N_7256);
nand U8507 (N_8507,N_7618,N_8346);
and U8508 (N_8508,N_8233,N_8026);
and U8509 (N_8509,N_7986,N_8358);
nand U8510 (N_8510,N_7340,N_7884);
xor U8511 (N_8511,N_7940,N_7836);
or U8512 (N_8512,N_7908,N_7764);
or U8513 (N_8513,N_7889,N_7266);
and U8514 (N_8514,N_7239,N_8183);
xnor U8515 (N_8515,N_7369,N_7810);
and U8516 (N_8516,N_8327,N_7789);
nand U8517 (N_8517,N_7976,N_7890);
nor U8518 (N_8518,N_7417,N_8070);
xnor U8519 (N_8519,N_7364,N_7546);
xor U8520 (N_8520,N_7900,N_7717);
nor U8521 (N_8521,N_7592,N_7467);
xor U8522 (N_8522,N_8155,N_7233);
nor U8523 (N_8523,N_7399,N_7867);
or U8524 (N_8524,N_7657,N_7970);
and U8525 (N_8525,N_7473,N_7483);
and U8526 (N_8526,N_7832,N_7395);
or U8527 (N_8527,N_7954,N_7298);
nor U8528 (N_8528,N_8315,N_7258);
nor U8529 (N_8529,N_8282,N_7204);
nand U8530 (N_8530,N_7388,N_8320);
nand U8531 (N_8531,N_7567,N_7227);
or U8532 (N_8532,N_7509,N_7241);
or U8533 (N_8533,N_8115,N_7563);
nand U8534 (N_8534,N_7621,N_8113);
or U8535 (N_8535,N_8098,N_7994);
xor U8536 (N_8536,N_7343,N_7533);
nor U8537 (N_8537,N_7779,N_8278);
nor U8538 (N_8538,N_7965,N_8172);
xnor U8539 (N_8539,N_8075,N_7354);
or U8540 (N_8540,N_7402,N_7819);
nand U8541 (N_8541,N_7275,N_8127);
nor U8542 (N_8542,N_7927,N_8019);
and U8543 (N_8543,N_7686,N_8354);
nor U8544 (N_8544,N_7975,N_7658);
xnor U8545 (N_8545,N_7548,N_7302);
or U8546 (N_8546,N_7368,N_8043);
xnor U8547 (N_8547,N_8230,N_7944);
or U8548 (N_8548,N_7350,N_8074);
nor U8549 (N_8549,N_8049,N_7961);
nor U8550 (N_8550,N_7605,N_8143);
nor U8551 (N_8551,N_7359,N_7461);
and U8552 (N_8552,N_8004,N_7687);
or U8553 (N_8553,N_8148,N_8256);
xnor U8554 (N_8554,N_7597,N_7418);
nor U8555 (N_8555,N_7721,N_7812);
or U8556 (N_8556,N_7842,N_7445);
xnor U8557 (N_8557,N_7957,N_7762);
or U8558 (N_8558,N_7333,N_8059);
nor U8559 (N_8559,N_8046,N_8351);
or U8560 (N_8560,N_7243,N_7305);
or U8561 (N_8561,N_8361,N_7503);
nor U8562 (N_8562,N_8062,N_8311);
nor U8563 (N_8563,N_8253,N_7419);
and U8564 (N_8564,N_8142,N_8040);
xor U8565 (N_8565,N_7878,N_8054);
nor U8566 (N_8566,N_7413,N_7873);
or U8567 (N_8567,N_8118,N_7282);
or U8568 (N_8568,N_7920,N_8395);
and U8569 (N_8569,N_7479,N_7960);
nor U8570 (N_8570,N_7829,N_8194);
xnor U8571 (N_8571,N_7459,N_7987);
nor U8572 (N_8572,N_7897,N_8290);
nor U8573 (N_8573,N_7728,N_7294);
nor U8574 (N_8574,N_7663,N_8080);
nand U8575 (N_8575,N_7255,N_7845);
and U8576 (N_8576,N_7457,N_7620);
nand U8577 (N_8577,N_7922,N_8159);
and U8578 (N_8578,N_7491,N_8356);
xnor U8579 (N_8579,N_7780,N_8226);
and U8580 (N_8580,N_7405,N_7538);
nor U8581 (N_8581,N_7817,N_8340);
or U8582 (N_8582,N_8052,N_8264);
nand U8583 (N_8583,N_8061,N_8228);
nand U8584 (N_8584,N_7766,N_7426);
or U8585 (N_8585,N_8248,N_8242);
nor U8586 (N_8586,N_7641,N_7234);
and U8587 (N_8587,N_7430,N_8099);
and U8588 (N_8588,N_7440,N_7504);
xnor U8589 (N_8589,N_7387,N_8073);
and U8590 (N_8590,N_7776,N_7593);
and U8591 (N_8591,N_7231,N_7236);
xor U8592 (N_8592,N_7301,N_7676);
nor U8593 (N_8593,N_7844,N_7557);
nand U8594 (N_8594,N_7929,N_8295);
nor U8595 (N_8595,N_8161,N_7685);
xor U8596 (N_8596,N_8379,N_8084);
or U8597 (N_8597,N_8217,N_7487);
xnor U8598 (N_8598,N_7412,N_8163);
xnor U8599 (N_8599,N_8177,N_8318);
and U8600 (N_8600,N_7537,N_7383);
nand U8601 (N_8601,N_7913,N_7403);
nand U8602 (N_8602,N_7835,N_8342);
nor U8603 (N_8603,N_7536,N_8063);
and U8604 (N_8604,N_7318,N_7332);
nor U8605 (N_8605,N_7669,N_7299);
nor U8606 (N_8606,N_7784,N_8182);
or U8607 (N_8607,N_8220,N_8067);
and U8608 (N_8608,N_8189,N_8185);
or U8609 (N_8609,N_7903,N_7887);
nand U8610 (N_8610,N_8112,N_8018);
nand U8611 (N_8611,N_7254,N_8109);
or U8612 (N_8612,N_8164,N_8271);
xnor U8613 (N_8613,N_7818,N_7208);
or U8614 (N_8614,N_7224,N_7598);
nand U8615 (N_8615,N_7656,N_8083);
xnor U8616 (N_8616,N_7352,N_7494);
xnor U8617 (N_8617,N_7923,N_7542);
or U8618 (N_8618,N_7460,N_7797);
or U8619 (N_8619,N_7619,N_8044);
and U8620 (N_8620,N_8333,N_8072);
or U8621 (N_8621,N_8394,N_7360);
and U8622 (N_8622,N_7367,N_7636);
xnor U8623 (N_8623,N_7361,N_8249);
nor U8624 (N_8624,N_8330,N_7414);
nand U8625 (N_8625,N_7666,N_7490);
xnor U8626 (N_8626,N_7222,N_8197);
nand U8627 (N_8627,N_7376,N_7303);
nor U8628 (N_8628,N_7719,N_8254);
nor U8629 (N_8629,N_7265,N_7761);
and U8630 (N_8630,N_8234,N_8300);
and U8631 (N_8631,N_7612,N_7759);
xor U8632 (N_8632,N_8276,N_8348);
and U8633 (N_8633,N_7338,N_7217);
xor U8634 (N_8634,N_7575,N_8374);
nand U8635 (N_8635,N_8137,N_7511);
or U8636 (N_8636,N_8227,N_8028);
and U8637 (N_8637,N_7941,N_8384);
nand U8638 (N_8638,N_7942,N_7715);
or U8639 (N_8639,N_7323,N_7604);
or U8640 (N_8640,N_8312,N_7462);
nor U8641 (N_8641,N_8365,N_7824);
nor U8642 (N_8642,N_7599,N_7623);
and U8643 (N_8643,N_7770,N_7499);
xor U8644 (N_8644,N_8317,N_7322);
and U8645 (N_8645,N_7311,N_7220);
nand U8646 (N_8646,N_8002,N_8274);
and U8647 (N_8647,N_7654,N_7949);
xnor U8648 (N_8648,N_8293,N_8218);
xor U8649 (N_8649,N_7876,N_7894);
nand U8650 (N_8650,N_8231,N_8273);
and U8651 (N_8651,N_7978,N_7314);
nand U8652 (N_8652,N_7948,N_7951);
xnor U8653 (N_8653,N_7837,N_7611);
and U8654 (N_8654,N_8008,N_8360);
nand U8655 (N_8655,N_7740,N_7773);
or U8656 (N_8656,N_7209,N_8141);
xor U8657 (N_8657,N_8206,N_7437);
nand U8658 (N_8658,N_8272,N_8285);
nand U8659 (N_8659,N_7329,N_8123);
xnor U8660 (N_8660,N_7261,N_7391);
and U8661 (N_8661,N_7603,N_7650);
and U8662 (N_8662,N_7447,N_7915);
or U8663 (N_8663,N_7857,N_7992);
xnor U8664 (N_8664,N_8309,N_7775);
and U8665 (N_8665,N_7203,N_7956);
or U8666 (N_8666,N_7966,N_7210);
nor U8667 (N_8667,N_8378,N_7221);
or U8668 (N_8668,N_7828,N_8027);
and U8669 (N_8669,N_8266,N_7555);
nand U8670 (N_8670,N_7560,N_7484);
or U8671 (N_8671,N_7614,N_7974);
xnor U8672 (N_8672,N_8292,N_7624);
and U8673 (N_8673,N_7807,N_7415);
xor U8674 (N_8674,N_7649,N_7458);
nand U8675 (N_8675,N_7284,N_7240);
xnor U8676 (N_8676,N_7286,N_7547);
nor U8677 (N_8677,N_8304,N_7813);
nand U8678 (N_8678,N_8000,N_7720);
nand U8679 (N_8679,N_7485,N_7427);
nor U8680 (N_8680,N_7864,N_8184);
or U8681 (N_8681,N_8088,N_7292);
nand U8682 (N_8682,N_8250,N_8319);
xnor U8683 (N_8683,N_8385,N_7771);
xnor U8684 (N_8684,N_8196,N_7896);
and U8685 (N_8685,N_7544,N_7726);
and U8686 (N_8686,N_7521,N_7269);
or U8687 (N_8687,N_7595,N_7823);
xor U8688 (N_8688,N_7506,N_7850);
nor U8689 (N_8689,N_8090,N_7655);
nor U8690 (N_8690,N_7809,N_7997);
and U8691 (N_8691,N_7285,N_7320);
nor U8692 (N_8692,N_7651,N_7979);
nand U8693 (N_8693,N_7273,N_8245);
nor U8694 (N_8694,N_7508,N_7788);
nor U8695 (N_8695,N_7288,N_8007);
or U8696 (N_8696,N_7804,N_7748);
or U8697 (N_8697,N_7875,N_7328);
xor U8698 (N_8698,N_7407,N_7205);
xnor U8699 (N_8699,N_7510,N_7590);
nand U8700 (N_8700,N_7851,N_7709);
xor U8701 (N_8701,N_7385,N_7488);
xnor U8702 (N_8702,N_7355,N_7384);
nor U8703 (N_8703,N_7370,N_8302);
or U8704 (N_8704,N_7398,N_7926);
and U8705 (N_8705,N_7225,N_7993);
xor U8706 (N_8706,N_8322,N_8373);
or U8707 (N_8707,N_7394,N_7519);
or U8708 (N_8708,N_7257,N_8057);
or U8709 (N_8709,N_7815,N_7463);
or U8710 (N_8710,N_7252,N_7319);
nor U8711 (N_8711,N_7373,N_7917);
nor U8712 (N_8712,N_8301,N_8205);
and U8713 (N_8713,N_7283,N_8047);
and U8714 (N_8714,N_7379,N_7895);
and U8715 (N_8715,N_8013,N_7223);
xnor U8716 (N_8716,N_8387,N_7262);
and U8717 (N_8717,N_7228,N_7950);
nand U8718 (N_8718,N_8041,N_8036);
xor U8719 (N_8719,N_7550,N_8174);
nor U8720 (N_8720,N_7237,N_8323);
xor U8721 (N_8721,N_7545,N_7420);
or U8722 (N_8722,N_8341,N_7424);
xor U8723 (N_8723,N_7711,N_8023);
or U8724 (N_8724,N_7708,N_8066);
and U8725 (N_8725,N_8160,N_8369);
or U8726 (N_8726,N_7629,N_7375);
xnor U8727 (N_8727,N_8357,N_7968);
nor U8728 (N_8728,N_7648,N_7280);
and U8729 (N_8729,N_7313,N_8329);
nand U8730 (N_8730,N_7742,N_8175);
and U8731 (N_8731,N_7465,N_7852);
and U8732 (N_8732,N_7907,N_7307);
xnor U8733 (N_8733,N_8265,N_8039);
and U8734 (N_8734,N_7667,N_8168);
nand U8735 (N_8735,N_8106,N_7752);
xnor U8736 (N_8736,N_7357,N_7562);
and U8737 (N_8737,N_7493,N_7646);
and U8738 (N_8738,N_7767,N_7914);
nand U8739 (N_8739,N_7806,N_7798);
nor U8740 (N_8740,N_7469,N_7849);
or U8741 (N_8741,N_7566,N_7753);
or U8742 (N_8742,N_7263,N_7718);
and U8743 (N_8743,N_7633,N_7870);
nand U8744 (N_8744,N_7855,N_8035);
or U8745 (N_8745,N_7931,N_8068);
xor U8746 (N_8746,N_8119,N_7963);
and U8747 (N_8747,N_8201,N_7400);
xnor U8748 (N_8748,N_7955,N_8239);
nor U8749 (N_8749,N_7749,N_7935);
nand U8750 (N_8750,N_8136,N_7757);
xor U8751 (N_8751,N_8307,N_7741);
nand U8752 (N_8752,N_8077,N_7251);
nor U8753 (N_8753,N_8014,N_7732);
nand U8754 (N_8754,N_7422,N_8316);
nor U8755 (N_8755,N_8104,N_8133);
nand U8756 (N_8756,N_8126,N_8381);
and U8757 (N_8757,N_7702,N_7758);
and U8758 (N_8758,N_7672,N_7684);
xnor U8759 (N_8759,N_7530,N_7703);
xnor U8760 (N_8760,N_8339,N_7326);
nor U8761 (N_8761,N_8096,N_7872);
and U8762 (N_8762,N_7561,N_8324);
nor U8763 (N_8763,N_7638,N_7406);
and U8764 (N_8764,N_7507,N_7834);
nand U8765 (N_8765,N_7751,N_7808);
nor U8766 (N_8766,N_7674,N_7518);
xnor U8767 (N_8767,N_8297,N_8371);
or U8768 (N_8768,N_7939,N_7909);
or U8769 (N_8769,N_8236,N_8048);
xor U8770 (N_8770,N_8162,N_8353);
xor U8771 (N_8771,N_7962,N_7589);
nand U8772 (N_8772,N_7833,N_7434);
nor U8773 (N_8773,N_7584,N_7443);
nor U8774 (N_8774,N_7682,N_8382);
and U8775 (N_8775,N_8214,N_7330);
nand U8776 (N_8776,N_7421,N_8392);
or U8777 (N_8777,N_8122,N_7693);
or U8778 (N_8778,N_8085,N_8076);
and U8779 (N_8779,N_7791,N_7928);
and U8780 (N_8780,N_8125,N_7308);
and U8781 (N_8781,N_7782,N_7229);
nor U8782 (N_8782,N_8243,N_7517);
nor U8783 (N_8783,N_7777,N_7380);
or U8784 (N_8784,N_7501,N_7552);
nor U8785 (N_8785,N_7356,N_7270);
nand U8786 (N_8786,N_8093,N_7856);
nor U8787 (N_8787,N_7643,N_7769);
xor U8788 (N_8788,N_8212,N_7683);
nor U8789 (N_8789,N_8009,N_7678);
xor U8790 (N_8790,N_8241,N_8006);
nand U8791 (N_8791,N_7206,N_7937);
and U8792 (N_8792,N_7670,N_7454);
and U8793 (N_8793,N_8114,N_7347);
or U8794 (N_8794,N_7339,N_7432);
and U8795 (N_8795,N_7731,N_7660);
nand U8796 (N_8796,N_8131,N_7397);
xnor U8797 (N_8797,N_7495,N_8110);
nor U8798 (N_8798,N_7553,N_7594);
xnor U8799 (N_8799,N_7390,N_8219);
nand U8800 (N_8800,N_8130,N_7497);
xnor U8801 (N_8801,N_7408,N_8200);
or U8802 (N_8802,N_7893,N_7918);
nand U8803 (N_8803,N_7747,N_7582);
nand U8804 (N_8804,N_7932,N_7304);
or U8805 (N_8805,N_7353,N_8389);
or U8806 (N_8806,N_7315,N_7482);
and U8807 (N_8807,N_8005,N_8033);
and U8808 (N_8808,N_7428,N_7756);
xnor U8809 (N_8809,N_8144,N_8030);
or U8810 (N_8810,N_7701,N_8138);
nand U8811 (N_8811,N_8390,N_7573);
nand U8812 (N_8812,N_7988,N_7316);
and U8813 (N_8813,N_8305,N_7378);
nor U8814 (N_8814,N_8064,N_8208);
or U8815 (N_8815,N_8176,N_8065);
nand U8816 (N_8816,N_7877,N_7698);
xor U8817 (N_8817,N_7568,N_7312);
nand U8818 (N_8818,N_8334,N_8079);
and U8819 (N_8819,N_8025,N_8268);
or U8820 (N_8820,N_7274,N_7232);
and U8821 (N_8821,N_7442,N_7578);
xnor U8822 (N_8822,N_7688,N_7476);
nor U8823 (N_8823,N_7898,N_7737);
or U8824 (N_8824,N_7455,N_8367);
and U8825 (N_8825,N_7435,N_8258);
xor U8826 (N_8826,N_8359,N_7549);
or U8827 (N_8827,N_7321,N_7535);
nand U8828 (N_8828,N_7543,N_8022);
nand U8829 (N_8829,N_8154,N_8259);
or U8830 (N_8830,N_7838,N_7990);
or U8831 (N_8831,N_7574,N_7943);
or U8832 (N_8832,N_7692,N_8193);
nor U8833 (N_8833,N_8267,N_7722);
nand U8834 (N_8834,N_7661,N_7456);
nand U8835 (N_8835,N_7706,N_7995);
and U8836 (N_8836,N_7522,N_8202);
nor U8837 (N_8837,N_7587,N_7626);
xor U8838 (N_8838,N_7602,N_7934);
xor U8839 (N_8839,N_8139,N_7699);
and U8840 (N_8840,N_8101,N_7358);
nor U8841 (N_8841,N_7480,N_8186);
nand U8842 (N_8842,N_7579,N_7754);
nand U8843 (N_8843,N_7377,N_7958);
and U8844 (N_8844,N_8100,N_7431);
xor U8845 (N_8845,N_8171,N_7554);
nand U8846 (N_8846,N_7760,N_7520);
and U8847 (N_8847,N_7662,N_8016);
xor U8848 (N_8848,N_8129,N_7831);
xnor U8849 (N_8849,N_7973,N_7570);
nor U8850 (N_8850,N_7733,N_7690);
or U8851 (N_8851,N_8229,N_7532);
xor U8852 (N_8852,N_8001,N_7489);
nand U8853 (N_8853,N_7977,N_8017);
xor U8854 (N_8854,N_8050,N_7746);
nand U8855 (N_8855,N_7637,N_8314);
and U8856 (N_8856,N_7606,N_8037);
nor U8857 (N_8857,N_7541,N_7772);
nor U8858 (N_8858,N_8366,N_8051);
nand U8859 (N_8859,N_7863,N_8108);
or U8860 (N_8860,N_7524,N_7734);
nor U8861 (N_8861,N_8280,N_7534);
nand U8862 (N_8862,N_7630,N_8167);
nand U8863 (N_8863,N_7866,N_7531);
or U8864 (N_8864,N_7348,N_7827);
xnor U8865 (N_8865,N_8283,N_7765);
or U8866 (N_8866,N_7946,N_8153);
xor U8867 (N_8867,N_8263,N_7858);
xor U8868 (N_8868,N_8308,N_7438);
and U8869 (N_8869,N_7902,N_7972);
xnor U8870 (N_8870,N_7805,N_8180);
xnor U8871 (N_8871,N_7583,N_8173);
and U8872 (N_8872,N_7681,N_7981);
nor U8873 (N_8873,N_7925,N_8343);
nor U8874 (N_8874,N_7245,N_7409);
nor U8875 (N_8875,N_8192,N_7615);
and U8876 (N_8876,N_7854,N_8362);
and U8877 (N_8877,N_8199,N_7572);
nor U8878 (N_8878,N_7401,N_7755);
nand U8879 (N_8879,N_7892,N_7512);
nand U8880 (N_8880,N_8255,N_8223);
or U8881 (N_8881,N_7953,N_7924);
or U8882 (N_8882,N_7750,N_8103);
nor U8883 (N_8883,N_7505,N_7446);
nand U8884 (N_8884,N_8156,N_7774);
or U8885 (N_8885,N_7300,N_8105);
nand U8886 (N_8886,N_7453,N_7349);
nand U8887 (N_8887,N_7883,N_8240);
xor U8888 (N_8888,N_7727,N_7653);
nor U8889 (N_8889,N_8116,N_7363);
nand U8890 (N_8890,N_7260,N_7644);
or U8891 (N_8891,N_7382,N_8326);
xnor U8892 (N_8892,N_7985,N_7527);
nand U8893 (N_8893,N_7569,N_8120);
and U8894 (N_8894,N_7853,N_8011);
or U8895 (N_8895,N_7799,N_8306);
or U8896 (N_8896,N_7423,N_7474);
xnor U8897 (N_8897,N_8117,N_7632);
nor U8898 (N_8898,N_7839,N_7816);
or U8899 (N_8899,N_7264,N_7642);
nor U8900 (N_8900,N_7716,N_8344);
nor U8901 (N_8901,N_7744,N_7441);
or U8902 (N_8902,N_8020,N_7971);
nand U8903 (N_8903,N_8056,N_7634);
or U8904 (N_8904,N_8380,N_7616);
or U8905 (N_8905,N_8209,N_8224);
nor U8906 (N_8906,N_8284,N_7617);
nand U8907 (N_8907,N_7888,N_7989);
xor U8908 (N_8908,N_8347,N_7219);
and U8909 (N_8909,N_7607,N_7551);
and U8910 (N_8910,N_7345,N_7911);
and U8911 (N_8911,N_8279,N_8328);
or U8912 (N_8912,N_7293,N_8332);
xnor U8913 (N_8913,N_7202,N_8338);
nand U8914 (N_8914,N_8331,N_7581);
nor U8915 (N_8915,N_7331,N_7865);
or U8916 (N_8916,N_7768,N_8260);
and U8917 (N_8917,N_8010,N_7861);
nand U8918 (N_8918,N_7393,N_7627);
nand U8919 (N_8919,N_8149,N_8024);
xnor U8920 (N_8920,N_8375,N_7291);
and U8921 (N_8921,N_7860,N_7904);
nor U8922 (N_8922,N_8399,N_7433);
nor U8923 (N_8923,N_7967,N_7577);
nor U8924 (N_8924,N_7444,N_8213);
nor U8925 (N_8925,N_8170,N_8060);
nor U8926 (N_8926,N_7372,N_7386);
nand U8927 (N_8927,N_8370,N_7729);
nor U8928 (N_8928,N_7610,N_7247);
or U8929 (N_8929,N_7576,N_8089);
xor U8930 (N_8930,N_7500,N_8222);
xor U8931 (N_8931,N_7486,N_8145);
nand U8932 (N_8932,N_8003,N_8015);
or U8933 (N_8933,N_7885,N_7327);
or U8934 (N_8934,N_7425,N_7235);
nand U8935 (N_8935,N_7787,N_8289);
and U8936 (N_8936,N_8078,N_7287);
and U8937 (N_8937,N_8094,N_7801);
and U8938 (N_8938,N_7795,N_8393);
and U8939 (N_8939,N_7449,N_7763);
nor U8940 (N_8940,N_7279,N_8165);
and U8941 (N_8941,N_8261,N_7596);
and U8942 (N_8942,N_7916,N_7613);
or U8943 (N_8943,N_7242,N_8372);
or U8944 (N_8944,N_7700,N_8207);
nand U8945 (N_8945,N_7608,N_7448);
xor U8946 (N_8946,N_8377,N_7346);
or U8947 (N_8947,N_7947,N_7411);
or U8948 (N_8948,N_7790,N_8128);
nand U8949 (N_8949,N_7847,N_8124);
xor U8950 (N_8950,N_7899,N_8325);
xor U8951 (N_8951,N_7738,N_8396);
xor U8952 (N_8952,N_7498,N_8294);
or U8953 (N_8953,N_8247,N_8303);
and U8954 (N_8954,N_8178,N_8150);
or U8955 (N_8955,N_7830,N_7496);
nor U8956 (N_8956,N_7337,N_7871);
nand U8957 (N_8957,N_8097,N_7381);
or U8958 (N_8958,N_8298,N_8012);
nand U8959 (N_8959,N_8270,N_7365);
xor U8960 (N_8960,N_7226,N_7341);
nor U8961 (N_8961,N_7933,N_7472);
xnor U8962 (N_8962,N_8111,N_8045);
nand U8963 (N_8963,N_7869,N_7639);
nand U8964 (N_8964,N_8188,N_8132);
or U8965 (N_8965,N_7697,N_7601);
nor U8966 (N_8966,N_7325,N_8181);
or U8967 (N_8967,N_8086,N_8031);
nand U8968 (N_8968,N_8029,N_8321);
or U8969 (N_8969,N_8345,N_7516);
or U8970 (N_8970,N_8232,N_7984);
and U8971 (N_8971,N_7725,N_7295);
and U8972 (N_8972,N_8244,N_8203);
nand U8973 (N_8973,N_8134,N_7802);
xor U8974 (N_8974,N_7625,N_8246);
nand U8975 (N_8975,N_8053,N_7820);
and U8976 (N_8976,N_8221,N_7539);
or U8977 (N_8977,N_7980,N_7945);
and U8978 (N_8978,N_7814,N_8034);
xnor U8979 (N_8979,N_7466,N_7952);
or U8980 (N_8980,N_7580,N_8225);
and U8981 (N_8981,N_7216,N_7846);
nand U8982 (N_8982,N_8169,N_7296);
nand U8983 (N_8983,N_7436,N_8081);
or U8984 (N_8984,N_7713,N_8215);
and U8985 (N_8985,N_8238,N_8216);
or U8986 (N_8986,N_7351,N_8121);
and U8987 (N_8987,N_7344,N_8397);
nor U8988 (N_8988,N_8204,N_7218);
and U8989 (N_8989,N_7253,N_7556);
nand U8990 (N_8990,N_7640,N_7558);
xnor U8991 (N_8991,N_7276,N_7609);
nand U8992 (N_8992,N_8152,N_7585);
nor U8993 (N_8993,N_7215,N_8032);
xor U8994 (N_8994,N_7783,N_8091);
nor U8995 (N_8995,N_7652,N_7310);
nand U8996 (N_8996,N_7468,N_7268);
nor U8997 (N_8997,N_7525,N_8275);
nor U8998 (N_8998,N_7450,N_7540);
or U8999 (N_8999,N_7921,N_7244);
xor U9000 (N_9000,N_7687,N_7540);
nor U9001 (N_9001,N_8269,N_7785);
nand U9002 (N_9002,N_7685,N_7323);
xor U9003 (N_9003,N_8307,N_8174);
and U9004 (N_9004,N_7712,N_7440);
or U9005 (N_9005,N_7204,N_7988);
nor U9006 (N_9006,N_7289,N_7537);
nor U9007 (N_9007,N_7873,N_7226);
and U9008 (N_9008,N_8308,N_7930);
or U9009 (N_9009,N_8104,N_7921);
nor U9010 (N_9010,N_8373,N_8255);
xor U9011 (N_9011,N_7678,N_7556);
or U9012 (N_9012,N_7882,N_8063);
nor U9013 (N_9013,N_7932,N_7643);
nor U9014 (N_9014,N_7765,N_7461);
nor U9015 (N_9015,N_7470,N_7535);
nand U9016 (N_9016,N_7370,N_7913);
and U9017 (N_9017,N_8014,N_8292);
nor U9018 (N_9018,N_8169,N_8304);
xnor U9019 (N_9019,N_7570,N_7758);
xor U9020 (N_9020,N_8216,N_8086);
nor U9021 (N_9021,N_7977,N_7992);
or U9022 (N_9022,N_7862,N_7796);
or U9023 (N_9023,N_8288,N_7413);
nor U9024 (N_9024,N_7576,N_8213);
nor U9025 (N_9025,N_7531,N_7420);
and U9026 (N_9026,N_7546,N_7248);
nand U9027 (N_9027,N_8142,N_7723);
or U9028 (N_9028,N_7938,N_7466);
xor U9029 (N_9029,N_8178,N_8065);
and U9030 (N_9030,N_7417,N_7964);
nand U9031 (N_9031,N_7632,N_7978);
xor U9032 (N_9032,N_8087,N_7383);
nor U9033 (N_9033,N_8163,N_7927);
xnor U9034 (N_9034,N_8147,N_7259);
xor U9035 (N_9035,N_7525,N_7443);
xnor U9036 (N_9036,N_7368,N_7916);
nand U9037 (N_9037,N_7508,N_7684);
xnor U9038 (N_9038,N_7293,N_7723);
nor U9039 (N_9039,N_8376,N_7617);
nor U9040 (N_9040,N_8182,N_7333);
or U9041 (N_9041,N_7795,N_7402);
nor U9042 (N_9042,N_7519,N_7290);
xnor U9043 (N_9043,N_7376,N_7972);
or U9044 (N_9044,N_7574,N_8042);
nor U9045 (N_9045,N_7714,N_8204);
and U9046 (N_9046,N_7226,N_7841);
or U9047 (N_9047,N_7789,N_7567);
or U9048 (N_9048,N_7991,N_7824);
xnor U9049 (N_9049,N_7540,N_8342);
and U9050 (N_9050,N_7914,N_7833);
nor U9051 (N_9051,N_7861,N_8148);
nor U9052 (N_9052,N_7324,N_7595);
nor U9053 (N_9053,N_7475,N_8055);
nand U9054 (N_9054,N_7547,N_7302);
and U9055 (N_9055,N_8298,N_7294);
and U9056 (N_9056,N_7623,N_7995);
nand U9057 (N_9057,N_7415,N_7779);
or U9058 (N_9058,N_7644,N_8283);
nor U9059 (N_9059,N_7342,N_8214);
xnor U9060 (N_9060,N_8068,N_8099);
and U9061 (N_9061,N_7201,N_7221);
nand U9062 (N_9062,N_7387,N_8294);
and U9063 (N_9063,N_7419,N_7338);
nand U9064 (N_9064,N_8072,N_7899);
and U9065 (N_9065,N_7919,N_7968);
and U9066 (N_9066,N_8142,N_8360);
xnor U9067 (N_9067,N_7450,N_7726);
or U9068 (N_9068,N_7761,N_7626);
or U9069 (N_9069,N_8385,N_7586);
or U9070 (N_9070,N_7281,N_8246);
xnor U9071 (N_9071,N_7462,N_8000);
or U9072 (N_9072,N_8092,N_8233);
nor U9073 (N_9073,N_7464,N_7357);
or U9074 (N_9074,N_8167,N_7378);
nand U9075 (N_9075,N_8344,N_7757);
nor U9076 (N_9076,N_8113,N_7561);
or U9077 (N_9077,N_8175,N_7460);
nor U9078 (N_9078,N_7497,N_8047);
xnor U9079 (N_9079,N_8355,N_8392);
or U9080 (N_9080,N_7614,N_7394);
or U9081 (N_9081,N_8151,N_7663);
nand U9082 (N_9082,N_7307,N_8375);
nor U9083 (N_9083,N_7611,N_7380);
xnor U9084 (N_9084,N_7909,N_7385);
or U9085 (N_9085,N_7656,N_7568);
nand U9086 (N_9086,N_7822,N_7695);
nand U9087 (N_9087,N_7433,N_7386);
xor U9088 (N_9088,N_7242,N_7863);
and U9089 (N_9089,N_7508,N_7200);
and U9090 (N_9090,N_8063,N_7825);
and U9091 (N_9091,N_7771,N_7247);
or U9092 (N_9092,N_8290,N_7766);
xor U9093 (N_9093,N_7390,N_7964);
nor U9094 (N_9094,N_7707,N_8347);
or U9095 (N_9095,N_7428,N_7217);
nor U9096 (N_9096,N_7339,N_7541);
nand U9097 (N_9097,N_8202,N_7295);
nor U9098 (N_9098,N_7370,N_8358);
and U9099 (N_9099,N_7789,N_7674);
nor U9100 (N_9100,N_7774,N_7723);
nand U9101 (N_9101,N_7262,N_7415);
and U9102 (N_9102,N_8281,N_7323);
and U9103 (N_9103,N_7823,N_7316);
nor U9104 (N_9104,N_7927,N_7834);
or U9105 (N_9105,N_8205,N_7247);
or U9106 (N_9106,N_8088,N_8156);
nor U9107 (N_9107,N_7904,N_7300);
or U9108 (N_9108,N_7202,N_7604);
nand U9109 (N_9109,N_7432,N_7921);
xnor U9110 (N_9110,N_7415,N_8356);
nand U9111 (N_9111,N_8154,N_8371);
nand U9112 (N_9112,N_8369,N_7333);
nand U9113 (N_9113,N_8202,N_8024);
and U9114 (N_9114,N_7288,N_7854);
xnor U9115 (N_9115,N_8379,N_8388);
xnor U9116 (N_9116,N_7658,N_8341);
and U9117 (N_9117,N_8013,N_7986);
nand U9118 (N_9118,N_7814,N_8069);
nor U9119 (N_9119,N_8163,N_7315);
or U9120 (N_9120,N_8058,N_7557);
nor U9121 (N_9121,N_8193,N_7822);
or U9122 (N_9122,N_7732,N_8051);
nor U9123 (N_9123,N_8095,N_7729);
xnor U9124 (N_9124,N_7565,N_8217);
or U9125 (N_9125,N_7603,N_7288);
and U9126 (N_9126,N_7974,N_7885);
nand U9127 (N_9127,N_7823,N_8212);
or U9128 (N_9128,N_7824,N_7814);
or U9129 (N_9129,N_7276,N_8002);
xor U9130 (N_9130,N_7692,N_7378);
xor U9131 (N_9131,N_7768,N_7957);
and U9132 (N_9132,N_7576,N_7923);
xor U9133 (N_9133,N_7569,N_7713);
nand U9134 (N_9134,N_7723,N_8149);
and U9135 (N_9135,N_7444,N_7613);
and U9136 (N_9136,N_8357,N_8307);
or U9137 (N_9137,N_7661,N_7849);
and U9138 (N_9138,N_8390,N_7709);
nand U9139 (N_9139,N_8393,N_8043);
or U9140 (N_9140,N_7807,N_8282);
nor U9141 (N_9141,N_7253,N_7672);
or U9142 (N_9142,N_7777,N_7950);
nand U9143 (N_9143,N_8258,N_8357);
and U9144 (N_9144,N_7202,N_7843);
nand U9145 (N_9145,N_7993,N_7478);
nor U9146 (N_9146,N_8273,N_7201);
xor U9147 (N_9147,N_8361,N_7963);
nand U9148 (N_9148,N_7803,N_7471);
or U9149 (N_9149,N_8290,N_8091);
and U9150 (N_9150,N_7616,N_7249);
or U9151 (N_9151,N_7399,N_7492);
nand U9152 (N_9152,N_7295,N_7788);
and U9153 (N_9153,N_7932,N_7428);
nor U9154 (N_9154,N_7527,N_7886);
xnor U9155 (N_9155,N_8317,N_7370);
nor U9156 (N_9156,N_8149,N_7713);
or U9157 (N_9157,N_8209,N_8313);
xnor U9158 (N_9158,N_8124,N_7401);
nor U9159 (N_9159,N_7652,N_7840);
xor U9160 (N_9160,N_8063,N_8081);
xnor U9161 (N_9161,N_8110,N_7990);
or U9162 (N_9162,N_7494,N_7245);
or U9163 (N_9163,N_7344,N_8232);
nand U9164 (N_9164,N_7846,N_7650);
nand U9165 (N_9165,N_8158,N_7853);
and U9166 (N_9166,N_8143,N_8345);
or U9167 (N_9167,N_7250,N_7889);
and U9168 (N_9168,N_7641,N_8311);
nand U9169 (N_9169,N_8008,N_7412);
and U9170 (N_9170,N_8176,N_7241);
nand U9171 (N_9171,N_7450,N_7967);
nand U9172 (N_9172,N_7461,N_7539);
or U9173 (N_9173,N_7219,N_7929);
nand U9174 (N_9174,N_7424,N_7867);
nand U9175 (N_9175,N_7740,N_7475);
and U9176 (N_9176,N_7237,N_8073);
and U9177 (N_9177,N_7911,N_8356);
xor U9178 (N_9178,N_8063,N_8002);
nand U9179 (N_9179,N_7281,N_7919);
or U9180 (N_9180,N_8115,N_8197);
nand U9181 (N_9181,N_7549,N_7796);
xnor U9182 (N_9182,N_7934,N_8040);
and U9183 (N_9183,N_7353,N_7939);
nand U9184 (N_9184,N_8145,N_7979);
or U9185 (N_9185,N_7815,N_7408);
nand U9186 (N_9186,N_8270,N_7649);
or U9187 (N_9187,N_7366,N_8066);
and U9188 (N_9188,N_7611,N_7819);
nand U9189 (N_9189,N_7831,N_7694);
or U9190 (N_9190,N_8191,N_7579);
or U9191 (N_9191,N_8277,N_7911);
xnor U9192 (N_9192,N_7386,N_7900);
or U9193 (N_9193,N_7953,N_8270);
nand U9194 (N_9194,N_8079,N_7622);
xor U9195 (N_9195,N_8324,N_7550);
nand U9196 (N_9196,N_7963,N_7625);
nand U9197 (N_9197,N_7758,N_7998);
nor U9198 (N_9198,N_7773,N_8371);
and U9199 (N_9199,N_7660,N_7738);
nand U9200 (N_9200,N_7661,N_7643);
or U9201 (N_9201,N_8030,N_8028);
xor U9202 (N_9202,N_7636,N_8363);
nor U9203 (N_9203,N_7474,N_7997);
nor U9204 (N_9204,N_8185,N_8068);
nand U9205 (N_9205,N_8340,N_7399);
nand U9206 (N_9206,N_7550,N_7250);
nand U9207 (N_9207,N_7538,N_7215);
or U9208 (N_9208,N_7315,N_7828);
or U9209 (N_9209,N_8335,N_8176);
and U9210 (N_9210,N_7319,N_7468);
nand U9211 (N_9211,N_7233,N_8349);
or U9212 (N_9212,N_8145,N_8195);
nor U9213 (N_9213,N_8227,N_7426);
nand U9214 (N_9214,N_8117,N_7409);
xnor U9215 (N_9215,N_7783,N_7515);
and U9216 (N_9216,N_8031,N_8116);
nor U9217 (N_9217,N_8109,N_8229);
and U9218 (N_9218,N_7448,N_8054);
or U9219 (N_9219,N_7359,N_8134);
xor U9220 (N_9220,N_7332,N_7246);
nand U9221 (N_9221,N_7813,N_8022);
and U9222 (N_9222,N_7896,N_8061);
nand U9223 (N_9223,N_8235,N_7203);
nand U9224 (N_9224,N_7927,N_8247);
and U9225 (N_9225,N_7668,N_7216);
and U9226 (N_9226,N_8344,N_7504);
xnor U9227 (N_9227,N_7541,N_8382);
and U9228 (N_9228,N_7462,N_7343);
nand U9229 (N_9229,N_7575,N_7415);
nor U9230 (N_9230,N_7230,N_8014);
nand U9231 (N_9231,N_7964,N_8056);
and U9232 (N_9232,N_7248,N_7223);
and U9233 (N_9233,N_8314,N_7374);
and U9234 (N_9234,N_8399,N_7969);
or U9235 (N_9235,N_8332,N_7590);
or U9236 (N_9236,N_7402,N_8382);
nor U9237 (N_9237,N_8244,N_7822);
nand U9238 (N_9238,N_7396,N_8283);
or U9239 (N_9239,N_7279,N_8168);
or U9240 (N_9240,N_7627,N_7817);
nand U9241 (N_9241,N_7272,N_8181);
and U9242 (N_9242,N_8172,N_7373);
xor U9243 (N_9243,N_7793,N_8245);
and U9244 (N_9244,N_7865,N_7406);
nand U9245 (N_9245,N_7983,N_7483);
or U9246 (N_9246,N_7241,N_7979);
nand U9247 (N_9247,N_7601,N_8348);
xnor U9248 (N_9248,N_7607,N_7527);
nor U9249 (N_9249,N_8087,N_7852);
nand U9250 (N_9250,N_7851,N_7975);
nand U9251 (N_9251,N_8246,N_7357);
xnor U9252 (N_9252,N_7436,N_7250);
nor U9253 (N_9253,N_8353,N_7490);
or U9254 (N_9254,N_8114,N_7550);
or U9255 (N_9255,N_7919,N_7756);
or U9256 (N_9256,N_8223,N_7637);
and U9257 (N_9257,N_7376,N_7280);
and U9258 (N_9258,N_7551,N_8049);
nand U9259 (N_9259,N_8379,N_7846);
nor U9260 (N_9260,N_7799,N_8088);
xor U9261 (N_9261,N_8082,N_7698);
nand U9262 (N_9262,N_7266,N_7840);
and U9263 (N_9263,N_8038,N_8088);
nand U9264 (N_9264,N_7870,N_7829);
nand U9265 (N_9265,N_7907,N_8051);
nand U9266 (N_9266,N_8390,N_8154);
and U9267 (N_9267,N_7530,N_7747);
nand U9268 (N_9268,N_7289,N_7638);
nand U9269 (N_9269,N_7449,N_8238);
and U9270 (N_9270,N_7463,N_7414);
and U9271 (N_9271,N_7921,N_7292);
nand U9272 (N_9272,N_8185,N_8237);
or U9273 (N_9273,N_7241,N_8059);
xnor U9274 (N_9274,N_7263,N_7913);
nor U9275 (N_9275,N_7910,N_7254);
and U9276 (N_9276,N_7804,N_7718);
or U9277 (N_9277,N_7585,N_7923);
and U9278 (N_9278,N_8172,N_7989);
and U9279 (N_9279,N_8091,N_7355);
xnor U9280 (N_9280,N_7512,N_7608);
and U9281 (N_9281,N_7961,N_7795);
and U9282 (N_9282,N_7758,N_7803);
nor U9283 (N_9283,N_7588,N_7800);
and U9284 (N_9284,N_7656,N_8347);
and U9285 (N_9285,N_7525,N_7869);
or U9286 (N_9286,N_7468,N_8375);
nor U9287 (N_9287,N_7899,N_7665);
nand U9288 (N_9288,N_7998,N_7380);
nand U9289 (N_9289,N_7647,N_8134);
xor U9290 (N_9290,N_8152,N_7391);
xnor U9291 (N_9291,N_7722,N_8041);
or U9292 (N_9292,N_7267,N_8394);
and U9293 (N_9293,N_7462,N_7463);
nand U9294 (N_9294,N_7777,N_7626);
xnor U9295 (N_9295,N_7477,N_8058);
and U9296 (N_9296,N_8220,N_8336);
nor U9297 (N_9297,N_7377,N_8199);
xnor U9298 (N_9298,N_8226,N_7584);
and U9299 (N_9299,N_7265,N_8152);
and U9300 (N_9300,N_8064,N_7774);
or U9301 (N_9301,N_7800,N_7884);
and U9302 (N_9302,N_7761,N_7774);
and U9303 (N_9303,N_8337,N_7428);
nor U9304 (N_9304,N_7866,N_8193);
or U9305 (N_9305,N_7501,N_8316);
and U9306 (N_9306,N_7730,N_7771);
nor U9307 (N_9307,N_7345,N_8279);
and U9308 (N_9308,N_8098,N_7748);
nor U9309 (N_9309,N_7856,N_7282);
xor U9310 (N_9310,N_8088,N_8289);
xnor U9311 (N_9311,N_8075,N_7683);
and U9312 (N_9312,N_7274,N_8018);
nor U9313 (N_9313,N_7437,N_7200);
xor U9314 (N_9314,N_7470,N_8190);
xnor U9315 (N_9315,N_7262,N_7277);
and U9316 (N_9316,N_7358,N_7758);
and U9317 (N_9317,N_7307,N_8203);
xor U9318 (N_9318,N_8157,N_8243);
xor U9319 (N_9319,N_7391,N_8367);
nor U9320 (N_9320,N_7320,N_7510);
xnor U9321 (N_9321,N_7532,N_8065);
nand U9322 (N_9322,N_8012,N_7669);
and U9323 (N_9323,N_7435,N_7967);
or U9324 (N_9324,N_7793,N_7480);
nand U9325 (N_9325,N_8317,N_7974);
nor U9326 (N_9326,N_7760,N_8379);
and U9327 (N_9327,N_7660,N_7874);
nand U9328 (N_9328,N_8063,N_7573);
or U9329 (N_9329,N_8188,N_8335);
and U9330 (N_9330,N_7878,N_7450);
nor U9331 (N_9331,N_8237,N_7371);
nor U9332 (N_9332,N_7512,N_7679);
nor U9333 (N_9333,N_7572,N_7702);
and U9334 (N_9334,N_7440,N_8281);
or U9335 (N_9335,N_7920,N_8226);
nor U9336 (N_9336,N_7301,N_8068);
and U9337 (N_9337,N_7747,N_7214);
nor U9338 (N_9338,N_7553,N_7538);
and U9339 (N_9339,N_7470,N_7965);
and U9340 (N_9340,N_8014,N_7520);
nor U9341 (N_9341,N_7510,N_7983);
nand U9342 (N_9342,N_8115,N_7475);
or U9343 (N_9343,N_7582,N_8187);
nand U9344 (N_9344,N_7212,N_7820);
nor U9345 (N_9345,N_8335,N_8251);
nor U9346 (N_9346,N_7624,N_7413);
nand U9347 (N_9347,N_7473,N_7736);
xnor U9348 (N_9348,N_8344,N_8298);
nor U9349 (N_9349,N_7331,N_7486);
or U9350 (N_9350,N_7893,N_8222);
xnor U9351 (N_9351,N_7898,N_7206);
and U9352 (N_9352,N_8045,N_7685);
nand U9353 (N_9353,N_8183,N_7242);
or U9354 (N_9354,N_8253,N_7629);
nor U9355 (N_9355,N_7291,N_8391);
nand U9356 (N_9356,N_7660,N_7907);
nand U9357 (N_9357,N_7270,N_7218);
nor U9358 (N_9358,N_7981,N_8112);
and U9359 (N_9359,N_7495,N_7318);
xor U9360 (N_9360,N_7394,N_8148);
nand U9361 (N_9361,N_7975,N_7451);
and U9362 (N_9362,N_8074,N_8080);
and U9363 (N_9363,N_8211,N_7544);
xor U9364 (N_9364,N_8270,N_8243);
and U9365 (N_9365,N_7867,N_7300);
and U9366 (N_9366,N_8380,N_8054);
nand U9367 (N_9367,N_7382,N_8243);
or U9368 (N_9368,N_7495,N_8254);
nor U9369 (N_9369,N_7437,N_8175);
nand U9370 (N_9370,N_7830,N_7915);
nor U9371 (N_9371,N_8025,N_7627);
nand U9372 (N_9372,N_7410,N_8185);
or U9373 (N_9373,N_7806,N_8119);
and U9374 (N_9374,N_8093,N_8289);
and U9375 (N_9375,N_7547,N_8343);
xor U9376 (N_9376,N_7516,N_7318);
nor U9377 (N_9377,N_7513,N_8113);
and U9378 (N_9378,N_7511,N_7823);
and U9379 (N_9379,N_8134,N_8372);
and U9380 (N_9380,N_7789,N_7424);
nor U9381 (N_9381,N_7546,N_7940);
and U9382 (N_9382,N_7946,N_8046);
and U9383 (N_9383,N_8352,N_7478);
xnor U9384 (N_9384,N_7402,N_7287);
or U9385 (N_9385,N_7378,N_7593);
or U9386 (N_9386,N_8107,N_7606);
nand U9387 (N_9387,N_7607,N_7938);
and U9388 (N_9388,N_7261,N_8250);
nor U9389 (N_9389,N_7833,N_8351);
nor U9390 (N_9390,N_8323,N_8107);
nor U9391 (N_9391,N_8195,N_8162);
nor U9392 (N_9392,N_7568,N_7967);
or U9393 (N_9393,N_8218,N_7832);
nor U9394 (N_9394,N_7382,N_7654);
nand U9395 (N_9395,N_8319,N_8115);
nor U9396 (N_9396,N_7930,N_7706);
and U9397 (N_9397,N_7707,N_7871);
or U9398 (N_9398,N_7532,N_7606);
xnor U9399 (N_9399,N_8336,N_7708);
nand U9400 (N_9400,N_7427,N_7389);
nor U9401 (N_9401,N_7629,N_8358);
xnor U9402 (N_9402,N_7478,N_8216);
or U9403 (N_9403,N_7968,N_8305);
xor U9404 (N_9404,N_7382,N_7855);
or U9405 (N_9405,N_8064,N_8135);
xor U9406 (N_9406,N_8169,N_7455);
nand U9407 (N_9407,N_8131,N_7792);
nor U9408 (N_9408,N_7498,N_8088);
and U9409 (N_9409,N_8241,N_7667);
nor U9410 (N_9410,N_7600,N_7854);
and U9411 (N_9411,N_8042,N_8374);
nand U9412 (N_9412,N_7618,N_8307);
xor U9413 (N_9413,N_7725,N_7224);
nor U9414 (N_9414,N_8199,N_7531);
and U9415 (N_9415,N_8371,N_8157);
xor U9416 (N_9416,N_7865,N_8362);
nand U9417 (N_9417,N_8312,N_7725);
or U9418 (N_9418,N_8095,N_7376);
nor U9419 (N_9419,N_8338,N_8010);
or U9420 (N_9420,N_7638,N_7562);
nand U9421 (N_9421,N_8327,N_8126);
nand U9422 (N_9422,N_8316,N_7204);
and U9423 (N_9423,N_7555,N_8041);
xor U9424 (N_9424,N_8077,N_7570);
and U9425 (N_9425,N_7517,N_7295);
nand U9426 (N_9426,N_8002,N_8219);
or U9427 (N_9427,N_7708,N_8124);
and U9428 (N_9428,N_8268,N_7691);
and U9429 (N_9429,N_7824,N_8070);
or U9430 (N_9430,N_7374,N_7651);
xnor U9431 (N_9431,N_7644,N_7983);
nor U9432 (N_9432,N_7829,N_7722);
nand U9433 (N_9433,N_7960,N_8216);
or U9434 (N_9434,N_8373,N_8307);
xor U9435 (N_9435,N_7436,N_7351);
nand U9436 (N_9436,N_8360,N_7557);
and U9437 (N_9437,N_7245,N_8269);
xor U9438 (N_9438,N_8023,N_7201);
nand U9439 (N_9439,N_7946,N_8313);
xor U9440 (N_9440,N_7438,N_7509);
xor U9441 (N_9441,N_7961,N_7375);
and U9442 (N_9442,N_7856,N_7629);
nand U9443 (N_9443,N_8111,N_7421);
nand U9444 (N_9444,N_8236,N_7762);
nand U9445 (N_9445,N_7555,N_7357);
xor U9446 (N_9446,N_7223,N_8213);
xnor U9447 (N_9447,N_7272,N_7729);
nor U9448 (N_9448,N_7429,N_7952);
xnor U9449 (N_9449,N_8154,N_7312);
nand U9450 (N_9450,N_7724,N_8059);
and U9451 (N_9451,N_8343,N_7574);
nand U9452 (N_9452,N_7913,N_8235);
nand U9453 (N_9453,N_8367,N_8154);
and U9454 (N_9454,N_7656,N_8173);
nor U9455 (N_9455,N_7411,N_8366);
or U9456 (N_9456,N_7419,N_8278);
nor U9457 (N_9457,N_7347,N_7628);
nor U9458 (N_9458,N_7671,N_7450);
xnor U9459 (N_9459,N_7519,N_7352);
nor U9460 (N_9460,N_7909,N_7581);
xnor U9461 (N_9461,N_7798,N_7241);
or U9462 (N_9462,N_7229,N_7681);
and U9463 (N_9463,N_7556,N_7696);
nor U9464 (N_9464,N_7997,N_7914);
and U9465 (N_9465,N_8014,N_8248);
or U9466 (N_9466,N_7519,N_8270);
xor U9467 (N_9467,N_7661,N_7262);
nand U9468 (N_9468,N_7785,N_8047);
or U9469 (N_9469,N_8273,N_7905);
nor U9470 (N_9470,N_8397,N_7384);
nor U9471 (N_9471,N_8376,N_7953);
and U9472 (N_9472,N_7935,N_7361);
nor U9473 (N_9473,N_7990,N_7564);
nor U9474 (N_9474,N_7563,N_8124);
nand U9475 (N_9475,N_7951,N_7692);
or U9476 (N_9476,N_7432,N_8377);
or U9477 (N_9477,N_8155,N_8123);
and U9478 (N_9478,N_8270,N_8351);
and U9479 (N_9479,N_7637,N_7972);
or U9480 (N_9480,N_8247,N_8182);
nand U9481 (N_9481,N_8035,N_7214);
nor U9482 (N_9482,N_8387,N_7345);
and U9483 (N_9483,N_7768,N_7530);
or U9484 (N_9484,N_8086,N_7669);
or U9485 (N_9485,N_7663,N_8284);
nand U9486 (N_9486,N_7545,N_7698);
and U9487 (N_9487,N_7701,N_7611);
and U9488 (N_9488,N_7527,N_7231);
nand U9489 (N_9489,N_7978,N_7968);
or U9490 (N_9490,N_8230,N_7614);
nand U9491 (N_9491,N_8378,N_8343);
or U9492 (N_9492,N_7362,N_7499);
or U9493 (N_9493,N_7913,N_7585);
and U9494 (N_9494,N_7988,N_7789);
nor U9495 (N_9495,N_8109,N_7283);
nor U9496 (N_9496,N_7478,N_7391);
nand U9497 (N_9497,N_7999,N_7293);
nand U9498 (N_9498,N_7817,N_7546);
xor U9499 (N_9499,N_7354,N_7901);
or U9500 (N_9500,N_7512,N_8048);
or U9501 (N_9501,N_8282,N_7779);
or U9502 (N_9502,N_7402,N_8357);
nand U9503 (N_9503,N_8243,N_7252);
and U9504 (N_9504,N_7754,N_8274);
nand U9505 (N_9505,N_7931,N_7724);
and U9506 (N_9506,N_7947,N_7261);
xnor U9507 (N_9507,N_7853,N_8198);
nand U9508 (N_9508,N_7713,N_7732);
or U9509 (N_9509,N_8097,N_8347);
nor U9510 (N_9510,N_7821,N_7605);
nand U9511 (N_9511,N_8326,N_7978);
nand U9512 (N_9512,N_7617,N_7513);
xor U9513 (N_9513,N_7389,N_7891);
and U9514 (N_9514,N_8239,N_7874);
nand U9515 (N_9515,N_8368,N_8105);
or U9516 (N_9516,N_7383,N_7938);
and U9517 (N_9517,N_8253,N_7790);
nand U9518 (N_9518,N_7626,N_7877);
nor U9519 (N_9519,N_8000,N_7557);
or U9520 (N_9520,N_8242,N_7743);
nor U9521 (N_9521,N_7827,N_7381);
nand U9522 (N_9522,N_7452,N_8034);
xor U9523 (N_9523,N_7491,N_7642);
and U9524 (N_9524,N_7847,N_7508);
nor U9525 (N_9525,N_8353,N_7404);
nand U9526 (N_9526,N_8306,N_8086);
and U9527 (N_9527,N_8190,N_8103);
or U9528 (N_9528,N_7391,N_7630);
xnor U9529 (N_9529,N_7654,N_7519);
nor U9530 (N_9530,N_8050,N_8126);
or U9531 (N_9531,N_7855,N_8288);
and U9532 (N_9532,N_8227,N_7859);
or U9533 (N_9533,N_8086,N_8273);
nor U9534 (N_9534,N_7726,N_8199);
or U9535 (N_9535,N_8272,N_8189);
or U9536 (N_9536,N_8161,N_7723);
and U9537 (N_9537,N_7761,N_8122);
nand U9538 (N_9538,N_7873,N_7848);
xor U9539 (N_9539,N_7688,N_8222);
xor U9540 (N_9540,N_7607,N_7479);
nor U9541 (N_9541,N_7287,N_7668);
nand U9542 (N_9542,N_8012,N_7963);
xor U9543 (N_9543,N_8234,N_8260);
and U9544 (N_9544,N_8155,N_8020);
and U9545 (N_9545,N_7391,N_7225);
or U9546 (N_9546,N_7223,N_8161);
nor U9547 (N_9547,N_7665,N_8099);
xor U9548 (N_9548,N_7383,N_8325);
nor U9549 (N_9549,N_7393,N_7792);
nor U9550 (N_9550,N_7401,N_8394);
nand U9551 (N_9551,N_7514,N_7217);
nor U9552 (N_9552,N_7825,N_7291);
or U9553 (N_9553,N_8082,N_7535);
nor U9554 (N_9554,N_7805,N_7985);
nor U9555 (N_9555,N_7725,N_7870);
nand U9556 (N_9556,N_8191,N_8080);
and U9557 (N_9557,N_8123,N_8220);
or U9558 (N_9558,N_7762,N_7577);
xor U9559 (N_9559,N_7764,N_8134);
xnor U9560 (N_9560,N_7982,N_8291);
and U9561 (N_9561,N_7421,N_8223);
nand U9562 (N_9562,N_7223,N_7750);
xor U9563 (N_9563,N_7989,N_7328);
nor U9564 (N_9564,N_7269,N_7431);
and U9565 (N_9565,N_7311,N_7825);
and U9566 (N_9566,N_7342,N_8058);
nor U9567 (N_9567,N_8267,N_8040);
xor U9568 (N_9568,N_7883,N_7778);
nor U9569 (N_9569,N_7699,N_7435);
xnor U9570 (N_9570,N_7521,N_8205);
nand U9571 (N_9571,N_7916,N_7804);
nand U9572 (N_9572,N_8342,N_7605);
or U9573 (N_9573,N_7917,N_7524);
xnor U9574 (N_9574,N_7833,N_8180);
nor U9575 (N_9575,N_8326,N_7815);
and U9576 (N_9576,N_7235,N_8370);
nand U9577 (N_9577,N_7345,N_7238);
or U9578 (N_9578,N_7286,N_8104);
nor U9579 (N_9579,N_8089,N_7567);
nor U9580 (N_9580,N_7721,N_7468);
or U9581 (N_9581,N_8342,N_7531);
xnor U9582 (N_9582,N_7265,N_7397);
nand U9583 (N_9583,N_7466,N_7945);
xor U9584 (N_9584,N_7811,N_7696);
or U9585 (N_9585,N_7210,N_8311);
nor U9586 (N_9586,N_7802,N_7595);
or U9587 (N_9587,N_7909,N_7730);
and U9588 (N_9588,N_8139,N_7292);
nand U9589 (N_9589,N_7997,N_7705);
nand U9590 (N_9590,N_7474,N_7386);
and U9591 (N_9591,N_8276,N_7230);
xnor U9592 (N_9592,N_7787,N_7210);
or U9593 (N_9593,N_7319,N_8066);
xnor U9594 (N_9594,N_7716,N_8345);
nor U9595 (N_9595,N_8391,N_7299);
nor U9596 (N_9596,N_7528,N_7631);
or U9597 (N_9597,N_8040,N_7737);
or U9598 (N_9598,N_8021,N_8193);
or U9599 (N_9599,N_8208,N_7334);
nor U9600 (N_9600,N_9240,N_8806);
or U9601 (N_9601,N_8487,N_9068);
nor U9602 (N_9602,N_9464,N_9223);
or U9603 (N_9603,N_9165,N_9413);
xnor U9604 (N_9604,N_8883,N_8637);
and U9605 (N_9605,N_8524,N_9439);
nand U9606 (N_9606,N_8607,N_8915);
nand U9607 (N_9607,N_8832,N_9216);
nor U9608 (N_9608,N_8685,N_8467);
nand U9609 (N_9609,N_8454,N_8777);
or U9610 (N_9610,N_9561,N_8711);
or U9611 (N_9611,N_9486,N_9229);
xor U9612 (N_9612,N_8845,N_9198);
and U9613 (N_9613,N_9112,N_9237);
and U9614 (N_9614,N_8407,N_9014);
nand U9615 (N_9615,N_9347,N_9479);
xor U9616 (N_9616,N_8597,N_9009);
nand U9617 (N_9617,N_8472,N_9061);
and U9618 (N_9618,N_9300,N_9338);
nor U9619 (N_9619,N_8692,N_8439);
nor U9620 (N_9620,N_8464,N_8859);
and U9621 (N_9621,N_9493,N_9100);
nand U9622 (N_9622,N_9277,N_8408);
nor U9623 (N_9623,N_9353,N_8432);
and U9624 (N_9624,N_9513,N_9386);
nand U9625 (N_9625,N_8961,N_8780);
and U9626 (N_9626,N_9005,N_8446);
or U9627 (N_9627,N_9156,N_8947);
xnor U9628 (N_9628,N_9304,N_9458);
xor U9629 (N_9629,N_8652,N_9474);
or U9630 (N_9630,N_8774,N_8686);
or U9631 (N_9631,N_8745,N_9242);
nand U9632 (N_9632,N_8940,N_8691);
or U9633 (N_9633,N_9398,N_9451);
nand U9634 (N_9634,N_9220,N_8603);
or U9635 (N_9635,N_8536,N_9105);
xor U9636 (N_9636,N_8715,N_8929);
and U9637 (N_9637,N_9440,N_9149);
nand U9638 (N_9638,N_9247,N_9031);
nand U9639 (N_9639,N_9143,N_9426);
nand U9640 (N_9640,N_8834,N_8746);
nor U9641 (N_9641,N_8705,N_8583);
or U9642 (N_9642,N_8800,N_8694);
or U9643 (N_9643,N_8903,N_9555);
xnor U9644 (N_9644,N_9423,N_8846);
or U9645 (N_9645,N_8957,N_8612);
and U9646 (N_9646,N_9572,N_9401);
and U9647 (N_9647,N_9550,N_8619);
nor U9648 (N_9648,N_9408,N_8604);
and U9649 (N_9649,N_8457,N_9511);
or U9650 (N_9650,N_9375,N_9567);
nand U9651 (N_9651,N_9089,N_9383);
xor U9652 (N_9652,N_8435,N_8789);
or U9653 (N_9653,N_9271,N_9318);
nand U9654 (N_9654,N_8977,N_9209);
and U9655 (N_9655,N_9202,N_8966);
and U9656 (N_9656,N_9453,N_8754);
nand U9657 (N_9657,N_8868,N_9121);
nor U9658 (N_9658,N_8700,N_8649);
nand U9659 (N_9659,N_8493,N_8932);
xnor U9660 (N_9660,N_8647,N_9134);
xor U9661 (N_9661,N_9399,N_8816);
nor U9662 (N_9662,N_8635,N_8999);
and U9663 (N_9663,N_8993,N_8554);
nor U9664 (N_9664,N_9189,N_9183);
or U9665 (N_9665,N_8858,N_9234);
nor U9666 (N_9666,N_8904,N_8876);
or U9667 (N_9667,N_9448,N_9050);
nand U9668 (N_9668,N_8786,N_8570);
or U9669 (N_9669,N_8781,N_8920);
nand U9670 (N_9670,N_9460,N_8519);
nand U9671 (N_9671,N_8926,N_9226);
or U9672 (N_9672,N_9060,N_8443);
and U9673 (N_9673,N_9406,N_9133);
xor U9674 (N_9674,N_8899,N_8797);
or U9675 (N_9675,N_8425,N_8989);
nor U9676 (N_9676,N_8974,N_9163);
nand U9677 (N_9677,N_8739,N_9580);
nor U9678 (N_9678,N_9267,N_9321);
and U9679 (N_9679,N_8831,N_8508);
xor U9680 (N_9680,N_9475,N_9340);
and U9681 (N_9681,N_9040,N_9144);
or U9682 (N_9682,N_9161,N_8605);
nand U9683 (N_9683,N_8488,N_8861);
xor U9684 (N_9684,N_8665,N_9431);
nor U9685 (N_9685,N_9319,N_8535);
nand U9686 (N_9686,N_9503,N_9492);
xor U9687 (N_9687,N_8849,N_9549);
and U9688 (N_9688,N_8482,N_8547);
xor U9689 (N_9689,N_9192,N_8842);
or U9690 (N_9690,N_8474,N_9313);
nand U9691 (N_9691,N_8577,N_9369);
nor U9692 (N_9692,N_8623,N_9544);
or U9693 (N_9693,N_9489,N_8772);
nor U9694 (N_9694,N_8550,N_9568);
nor U9695 (N_9695,N_8882,N_8941);
nor U9696 (N_9696,N_9291,N_9096);
nand U9697 (N_9697,N_8848,N_9152);
nand U9698 (N_9698,N_8783,N_9562);
and U9699 (N_9699,N_8466,N_9598);
or U9700 (N_9700,N_8891,N_9188);
and U9701 (N_9701,N_8960,N_8709);
or U9702 (N_9702,N_8679,N_8981);
or U9703 (N_9703,N_9368,N_8927);
nand U9704 (N_9704,N_9181,N_8541);
nand U9705 (N_9705,N_8833,N_8617);
nor U9706 (N_9706,N_9290,N_8835);
nand U9707 (N_9707,N_8996,N_9029);
nand U9708 (N_9708,N_8862,N_9552);
or U9709 (N_9709,N_9557,N_9257);
xor U9710 (N_9710,N_9113,N_8756);
nor U9711 (N_9711,N_8706,N_9403);
or U9712 (N_9712,N_8499,N_8656);
xnor U9713 (N_9713,N_9442,N_9505);
xnor U9714 (N_9714,N_8664,N_9421);
xor U9715 (N_9715,N_9323,N_8825);
xnor U9716 (N_9716,N_8818,N_9091);
nor U9717 (N_9717,N_9485,N_8463);
and U9718 (N_9718,N_8870,N_8813);
nand U9719 (N_9719,N_9055,N_8836);
and U9720 (N_9720,N_8651,N_8838);
or U9721 (N_9721,N_9044,N_9255);
xor U9722 (N_9722,N_8515,N_8918);
or U9723 (N_9723,N_9200,N_9024);
xnor U9724 (N_9724,N_9296,N_9175);
or U9725 (N_9725,N_8479,N_8791);
and U9726 (N_9726,N_8802,N_9350);
and U9727 (N_9727,N_8532,N_8520);
xnor U9728 (N_9728,N_9582,N_9452);
xnor U9729 (N_9729,N_9302,N_9420);
and U9730 (N_9730,N_9190,N_8478);
and U9731 (N_9731,N_8555,N_8695);
nand U9732 (N_9732,N_8452,N_9073);
or U9733 (N_9733,N_8702,N_9488);
or U9734 (N_9734,N_9483,N_9095);
and U9735 (N_9735,N_9027,N_8648);
or U9736 (N_9736,N_8863,N_9397);
and U9737 (N_9737,N_8782,N_9404);
nand U9738 (N_9738,N_8629,N_9494);
or U9739 (N_9739,N_9245,N_9136);
nand U9740 (N_9740,N_8733,N_9554);
nand U9741 (N_9741,N_8608,N_9160);
or U9742 (N_9742,N_9534,N_8423);
and U9743 (N_9743,N_8563,N_8560);
xor U9744 (N_9744,N_8809,N_8442);
or U9745 (N_9745,N_8760,N_9219);
nand U9746 (N_9746,N_8917,N_9306);
xor U9747 (N_9747,N_8406,N_8880);
or U9748 (N_9748,N_9239,N_9177);
nand U9749 (N_9749,N_8798,N_8494);
nor U9750 (N_9750,N_8765,N_8919);
and U9751 (N_9751,N_8663,N_8624);
or U9752 (N_9752,N_8573,N_8860);
nor U9753 (N_9753,N_9221,N_9123);
nand U9754 (N_9754,N_9496,N_9354);
nor U9755 (N_9755,N_8865,N_8755);
and U9756 (N_9756,N_8998,N_9543);
nor U9757 (N_9757,N_8699,N_8935);
xnor U9758 (N_9758,N_9072,N_9070);
and U9759 (N_9759,N_9418,N_8529);
and U9760 (N_9760,N_9179,N_9141);
nand U9761 (N_9761,N_9301,N_8574);
nor U9762 (N_9762,N_8805,N_9059);
xor U9763 (N_9763,N_8567,N_9305);
nor U9764 (N_9764,N_8548,N_9480);
nand U9765 (N_9765,N_8726,N_9395);
nor U9766 (N_9766,N_8586,N_9329);
nand U9767 (N_9767,N_9436,N_9583);
nand U9768 (N_9768,N_8588,N_8748);
xnor U9769 (N_9769,N_9108,N_9530);
nor U9770 (N_9770,N_9589,N_8698);
nand U9771 (N_9771,N_8433,N_9343);
and U9772 (N_9772,N_9570,N_8579);
xnor U9773 (N_9773,N_9285,N_8538);
or U9774 (N_9774,N_9118,N_8819);
or U9775 (N_9775,N_9541,N_9062);
and U9776 (N_9776,N_9414,N_8502);
or U9777 (N_9777,N_8662,N_9011);
or U9778 (N_9778,N_8741,N_8844);
nand U9779 (N_9779,N_8984,N_9129);
nand U9780 (N_9780,N_8730,N_9218);
or U9781 (N_9781,N_9187,N_9115);
or U9782 (N_9782,N_8785,N_8728);
and U9783 (N_9783,N_8717,N_8930);
xnor U9784 (N_9784,N_9125,N_9571);
or U9785 (N_9785,N_8719,N_9235);
nor U9786 (N_9786,N_9127,N_9457);
xor U9787 (N_9787,N_9046,N_9253);
nor U9788 (N_9788,N_8486,N_9191);
nand U9789 (N_9789,N_8767,N_9331);
nand U9790 (N_9790,N_8622,N_8757);
nand U9791 (N_9791,N_9010,N_9284);
nor U9792 (N_9792,N_8814,N_8743);
nand U9793 (N_9793,N_8507,N_9204);
or U9794 (N_9794,N_8952,N_9279);
or U9795 (N_9795,N_9384,N_8751);
or U9796 (N_9796,N_9491,N_9522);
nand U9797 (N_9797,N_8584,N_9259);
xor U9798 (N_9798,N_8992,N_9325);
nor U9799 (N_9799,N_8410,N_9154);
nand U9800 (N_9800,N_8804,N_8533);
xnor U9801 (N_9801,N_8946,N_9392);
nor U9802 (N_9802,N_9022,N_8485);
nand U9803 (N_9803,N_9114,N_8815);
or U9804 (N_9804,N_9506,N_9456);
or U9805 (N_9805,N_8986,N_8944);
or U9806 (N_9806,N_9167,N_9214);
nand U9807 (N_9807,N_8411,N_9248);
nor U9808 (N_9808,N_8824,N_8762);
or U9809 (N_9809,N_8596,N_9264);
nor U9810 (N_9810,N_9090,N_9415);
or U9811 (N_9811,N_9574,N_9539);
or U9812 (N_9812,N_8690,N_9042);
and U9813 (N_9813,N_8747,N_8997);
nor U9814 (N_9814,N_9232,N_8572);
nor U9815 (N_9815,N_9287,N_9314);
nand U9816 (N_9816,N_8630,N_8578);
and U9817 (N_9817,N_8907,N_9435);
nand U9818 (N_9818,N_8530,N_9510);
xnor U9819 (N_9819,N_8978,N_9047);
nor U9820 (N_9820,N_9288,N_9416);
or U9821 (N_9821,N_9071,N_8484);
and U9822 (N_9822,N_9504,N_8793);
nand U9823 (N_9823,N_9332,N_9577);
xnor U9824 (N_9824,N_8820,N_9205);
xnor U9825 (N_9825,N_8516,N_9518);
and U9826 (N_9826,N_9286,N_8811);
or U9827 (N_9827,N_8483,N_8489);
xnor U9828 (N_9828,N_9551,N_8626);
xnor U9829 (N_9829,N_8437,N_8826);
xnor U9830 (N_9830,N_8985,N_8459);
nand U9831 (N_9831,N_8497,N_8585);
or U9832 (N_9832,N_9131,N_9429);
nand U9833 (N_9833,N_9213,N_9462);
xor U9834 (N_9834,N_9361,N_9039);
nor U9835 (N_9835,N_9564,N_8720);
nor U9836 (N_9836,N_8616,N_8713);
or U9837 (N_9837,N_9434,N_9527);
nand U9838 (N_9838,N_9281,N_9363);
or U9839 (N_9839,N_8953,N_9256);
nand U9840 (N_9840,N_8436,N_9251);
nor U9841 (N_9841,N_9120,N_8632);
xor U9842 (N_9842,N_8921,N_8776);
nor U9843 (N_9843,N_9147,N_9182);
nor U9844 (N_9844,N_9591,N_9324);
nand U9845 (N_9845,N_9389,N_9124);
nor U9846 (N_9846,N_9393,N_9007);
and U9847 (N_9847,N_8803,N_8693);
xor U9848 (N_9848,N_9227,N_8556);
xnor U9849 (N_9849,N_8796,N_9473);
xnor U9850 (N_9850,N_9030,N_8707);
or U9851 (N_9851,N_9390,N_8643);
xnor U9852 (N_9852,N_9079,N_9508);
or U9853 (N_9853,N_9269,N_9316);
or U9854 (N_9854,N_8523,N_9579);
or U9855 (N_9855,N_9026,N_9367);
nand U9856 (N_9856,N_9352,N_8988);
xnor U9857 (N_9857,N_9588,N_9203);
xnor U9858 (N_9858,N_9412,N_8594);
nor U9859 (N_9859,N_9596,N_9020);
and U9860 (N_9860,N_8606,N_8902);
nor U9861 (N_9861,N_9049,N_8634);
nand U9862 (N_9862,N_9312,N_9166);
or U9863 (N_9863,N_8898,N_8644);
or U9864 (N_9864,N_9322,N_9444);
nor U9865 (N_9865,N_8905,N_9584);
and U9866 (N_9866,N_8874,N_8794);
nor U9867 (N_9867,N_9428,N_8956);
or U9868 (N_9868,N_9171,N_8681);
nor U9869 (N_9869,N_8689,N_9015);
xnor U9870 (N_9870,N_9465,N_9560);
and U9871 (N_9871,N_9116,N_9535);
or U9872 (N_9872,N_8799,N_8448);
xor U9873 (N_9873,N_8792,N_9587);
or U9874 (N_9874,N_9258,N_9034);
xor U9875 (N_9875,N_8668,N_8429);
and U9876 (N_9876,N_9529,N_9419);
or U9877 (N_9877,N_8673,N_8414);
and U9878 (N_9878,N_9374,N_8945);
or U9879 (N_9879,N_8795,N_8601);
nand U9880 (N_9880,N_8642,N_8853);
and U9881 (N_9881,N_8683,N_8742);
nand U9882 (N_9882,N_8650,N_8591);
nor U9883 (N_9883,N_9487,N_9507);
or U9884 (N_9884,N_9110,N_8473);
nand U9885 (N_9885,N_8812,N_9087);
xor U9886 (N_9886,N_9307,N_9335);
nor U9887 (N_9887,N_8959,N_8864);
xnor U9888 (N_9888,N_9337,N_9446);
and U9889 (N_9889,N_9599,N_9359);
xnor U9890 (N_9890,N_8503,N_8766);
or U9891 (N_9891,N_9278,N_8923);
nor U9892 (N_9892,N_9586,N_9012);
or U9893 (N_9893,N_8655,N_8498);
nor U9894 (N_9894,N_8771,N_8504);
nor U9895 (N_9895,N_9417,N_8893);
and U9896 (N_9896,N_8722,N_9159);
or U9897 (N_9897,N_9001,N_9261);
and U9898 (N_9898,N_9477,N_9490);
nand U9899 (N_9899,N_8445,N_9447);
and U9900 (N_9900,N_9400,N_9525);
nand U9901 (N_9901,N_8469,N_9233);
xnor U9902 (N_9902,N_8744,N_9468);
nand U9903 (N_9903,N_9531,N_8913);
and U9904 (N_9904,N_8735,N_8491);
nor U9905 (N_9905,N_9153,N_9019);
nor U9906 (N_9906,N_8906,N_9275);
nor U9907 (N_9907,N_9260,N_9138);
xor U9908 (N_9908,N_8732,N_9208);
xor U9909 (N_9909,N_8564,N_8495);
and U9910 (N_9910,N_9249,N_9481);
or U9911 (N_9911,N_9002,N_8708);
nand U9912 (N_9912,N_9008,N_9524);
xor U9913 (N_9913,N_8640,N_9088);
nor U9914 (N_9914,N_8413,N_8506);
and U9915 (N_9915,N_8723,N_8928);
or U9916 (N_9916,N_8509,N_8416);
xnor U9917 (N_9917,N_8545,N_9333);
xnor U9918 (N_9918,N_8587,N_9471);
and U9919 (N_9919,N_9207,N_9372);
nor U9920 (N_9920,N_8511,N_8561);
nand U9921 (N_9921,N_8675,N_9262);
or U9922 (N_9922,N_9362,N_9597);
xor U9923 (N_9923,N_8962,N_9268);
nor U9924 (N_9924,N_9553,N_9000);
xnor U9925 (N_9925,N_9168,N_8696);
and U9926 (N_9926,N_8636,N_9132);
nor U9927 (N_9927,N_9065,N_9520);
or U9928 (N_9928,N_9142,N_8847);
and U9929 (N_9929,N_9578,N_8740);
nand U9930 (N_9930,N_8595,N_9193);
nor U9931 (N_9931,N_9309,N_9157);
xor U9932 (N_9932,N_9536,N_9075);
nand U9933 (N_9933,N_8867,N_8759);
nor U9934 (N_9934,N_8419,N_8540);
xnor U9935 (N_9935,N_8866,N_9130);
and U9936 (N_9936,N_8678,N_9533);
xnor U9937 (N_9937,N_9320,N_8975);
nor U9938 (N_9938,N_8614,N_9150);
nand U9939 (N_9939,N_9559,N_9495);
and U9940 (N_9940,N_8982,N_8857);
and U9941 (N_9941,N_9484,N_9443);
nor U9942 (N_9942,N_8991,N_9581);
or U9943 (N_9943,N_8551,N_9348);
or U9944 (N_9944,N_8639,N_8557);
and U9945 (N_9945,N_8426,N_8476);
and U9946 (N_9946,N_9151,N_9140);
nand U9947 (N_9947,N_9006,N_9174);
nand U9948 (N_9948,N_9206,N_9173);
nor U9949 (N_9949,N_9217,N_9357);
or U9950 (N_9950,N_9407,N_8697);
xnor U9951 (N_9951,N_9212,N_9074);
xor U9952 (N_9952,N_8534,N_9238);
and U9953 (N_9953,N_9424,N_8471);
or U9954 (N_9954,N_8477,N_9425);
or U9955 (N_9955,N_8440,N_8527);
nand U9956 (N_9956,N_9328,N_8949);
and U9957 (N_9957,N_8618,N_8787);
or U9958 (N_9958,N_8518,N_9101);
nand U9959 (N_9959,N_8566,N_8676);
xnor U9960 (N_9960,N_8894,N_9083);
nor U9961 (N_9961,N_8914,N_9365);
nand U9962 (N_9962,N_8731,N_8613);
nor U9963 (N_9963,N_8768,N_8987);
and U9964 (N_9964,N_9199,N_9308);
xnor U9965 (N_9965,N_8670,N_9461);
nor U9966 (N_9966,N_8521,N_9515);
xor U9967 (N_9967,N_8828,N_8703);
or U9968 (N_9968,N_8610,N_9294);
nor U9969 (N_9969,N_8910,N_8990);
nor U9970 (N_9970,N_8531,N_9122);
and U9971 (N_9971,N_8434,N_9438);
xnor U9972 (N_9972,N_9405,N_8421);
or U9973 (N_9973,N_9241,N_8528);
nand U9974 (N_9974,N_9195,N_9593);
nor U9975 (N_9975,N_9086,N_9469);
nor U9976 (N_9976,N_9119,N_8983);
and U9977 (N_9977,N_8881,N_9080);
xor U9978 (N_9978,N_9117,N_8770);
or U9979 (N_9979,N_9076,N_8450);
nand U9980 (N_9980,N_9111,N_8729);
nand U9981 (N_9981,N_9037,N_9585);
and U9982 (N_9982,N_8465,N_9592);
xnor U9983 (N_9983,N_8453,N_9519);
xor U9984 (N_9984,N_9211,N_9215);
nand U9985 (N_9985,N_8852,N_8537);
or U9986 (N_9986,N_9162,N_9317);
nand U9987 (N_9987,N_8934,N_9021);
nand U9988 (N_9988,N_9243,N_8680);
nor U9989 (N_9989,N_8837,N_8925);
nor U9990 (N_9990,N_8420,N_9292);
or U9991 (N_9991,N_8775,N_9499);
xnor U9992 (N_9992,N_8973,N_9067);
nand U9993 (N_9993,N_9103,N_9053);
nand U9994 (N_9994,N_9128,N_8955);
or U9995 (N_9995,N_9376,N_8539);
nand U9996 (N_9996,N_9180,N_8628);
or U9997 (N_9997,N_8427,N_9422);
nand U9998 (N_9998,N_9263,N_9274);
nand U9999 (N_9999,N_8887,N_8638);
or U10000 (N_10000,N_8688,N_8401);
nand U10001 (N_10001,N_9538,N_9498);
and U10002 (N_10002,N_8549,N_8758);
xor U10003 (N_10003,N_8950,N_9194);
nand U10004 (N_10004,N_9135,N_9532);
and U10005 (N_10005,N_8620,N_9228);
or U10006 (N_10006,N_9360,N_8712);
xnor U10007 (N_10007,N_9336,N_9409);
or U10008 (N_10008,N_8951,N_8942);
or U10009 (N_10009,N_9058,N_8937);
nand U10010 (N_10010,N_8417,N_8470);
and U10011 (N_10011,N_9084,N_8451);
or U10012 (N_10012,N_8969,N_9517);
nand U10013 (N_10013,N_9590,N_9373);
or U10014 (N_10014,N_9097,N_8734);
and U10015 (N_10015,N_8823,N_8994);
nor U10016 (N_10016,N_9379,N_9197);
nor U10017 (N_10017,N_9236,N_9502);
or U10018 (N_10018,N_9225,N_9545);
xor U10019 (N_10019,N_8895,N_8682);
or U10020 (N_10020,N_9158,N_9003);
or U10021 (N_10021,N_8954,N_8590);
and U10022 (N_10022,N_9282,N_9346);
and U10023 (N_10023,N_9546,N_8856);
and U10024 (N_10024,N_9043,N_9509);
nor U10025 (N_10025,N_9077,N_8764);
and U10026 (N_10026,N_8901,N_9482);
xor U10027 (N_10027,N_9371,N_8995);
or U10028 (N_10028,N_9041,N_8580);
or U10029 (N_10029,N_9516,N_8840);
and U10030 (N_10030,N_9547,N_9164);
nor U10031 (N_10031,N_9558,N_9450);
nor U10032 (N_10032,N_8611,N_9295);
or U10033 (N_10033,N_8873,N_9437);
or U10034 (N_10034,N_9230,N_8412);
or U10035 (N_10035,N_8843,N_9540);
and U10036 (N_10036,N_8447,N_8671);
nand U10037 (N_10037,N_8615,N_8589);
nand U10038 (N_10038,N_9273,N_9170);
xor U10039 (N_10039,N_9478,N_9430);
xor U10040 (N_10040,N_9311,N_8911);
nor U10041 (N_10041,N_9345,N_9283);
or U10042 (N_10042,N_8460,N_9575);
nand U10043 (N_10043,N_9381,N_9201);
xnor U10044 (N_10044,N_9459,N_8641);
nand U10045 (N_10045,N_8542,N_9250);
or U10046 (N_10046,N_9016,N_9254);
and U10047 (N_10047,N_8916,N_9394);
nor U10048 (N_10048,N_9342,N_9548);
and U10049 (N_10049,N_8943,N_9056);
xnor U10050 (N_10050,N_8431,N_8822);
nor U10051 (N_10051,N_8877,N_8889);
nor U10052 (N_10052,N_8514,N_8871);
nand U10053 (N_10053,N_8778,N_8571);
xnor U10054 (N_10054,N_8609,N_8592);
and U10055 (N_10055,N_8409,N_9449);
xnor U10056 (N_10056,N_8599,N_8582);
nand U10057 (N_10057,N_9013,N_8888);
xnor U10058 (N_10058,N_8963,N_8627);
xnor U10059 (N_10059,N_8562,N_8908);
nor U10060 (N_10060,N_8854,N_8875);
nand U10061 (N_10061,N_8544,N_8701);
and U10062 (N_10062,N_8677,N_8481);
or U10063 (N_10063,N_8672,N_9210);
nand U10064 (N_10064,N_9036,N_9104);
xnor U10065 (N_10065,N_9265,N_9472);
and U10066 (N_10066,N_9402,N_9266);
or U10067 (N_10067,N_8968,N_9576);
nand U10068 (N_10068,N_8438,N_8621);
xor U10069 (N_10069,N_9396,N_8922);
xor U10070 (N_10070,N_9093,N_9387);
or U10071 (N_10071,N_9556,N_8807);
and U10072 (N_10072,N_8501,N_9512);
xnor U10073 (N_10073,N_8939,N_8565);
and U10074 (N_10074,N_8801,N_8879);
or U10075 (N_10075,N_8492,N_9356);
nor U10076 (N_10076,N_9280,N_8496);
xor U10077 (N_10077,N_8553,N_9018);
nor U10078 (N_10078,N_8851,N_8725);
xor U10079 (N_10079,N_8512,N_9391);
and U10080 (N_10080,N_9476,N_8449);
or U10081 (N_10081,N_8724,N_9364);
and U10082 (N_10082,N_9094,N_8552);
nor U10083 (N_10083,N_9004,N_9098);
nor U10084 (N_10084,N_8654,N_8422);
and U10085 (N_10085,N_9045,N_8896);
or U10086 (N_10086,N_8885,N_8829);
xor U10087 (N_10087,N_9303,N_8788);
nor U10088 (N_10088,N_8575,N_9382);
nor U10089 (N_10089,N_9048,N_9410);
or U10090 (N_10090,N_9052,N_8892);
or U10091 (N_10091,N_8827,N_8710);
nand U10092 (N_10092,N_8727,N_9246);
nand U10093 (N_10093,N_8721,N_8890);
nor U10094 (N_10094,N_9565,N_8458);
nor U10095 (N_10095,N_9032,N_9537);
xor U10096 (N_10096,N_9102,N_8657);
xor U10097 (N_10097,N_9563,N_8884);
and U10098 (N_10098,N_8653,N_8666);
nand U10099 (N_10099,N_9573,N_8704);
or U10100 (N_10100,N_8808,N_8581);
nand U10101 (N_10101,N_8569,N_8602);
nor U10102 (N_10102,N_8970,N_9099);
xor U10103 (N_10103,N_9252,N_9566);
nor U10104 (N_10104,N_8716,N_9595);
nor U10105 (N_10105,N_9388,N_9038);
or U10106 (N_10106,N_8424,N_8980);
and U10107 (N_10107,N_8749,N_8522);
nand U10108 (N_10108,N_8645,N_9289);
and U10109 (N_10109,N_8773,N_8912);
nand U10110 (N_10110,N_9231,N_8684);
and U10111 (N_10111,N_8964,N_8475);
nand U10112 (N_10112,N_8455,N_9569);
xnor U10113 (N_10113,N_8461,N_8405);
xnor U10114 (N_10114,N_8718,N_9334);
nand U10115 (N_10115,N_8568,N_9501);
xnor U10116 (N_10116,N_9351,N_8872);
and U10117 (N_10117,N_9139,N_9349);
xnor U10118 (N_10118,N_9092,N_8687);
or U10119 (N_10119,N_9054,N_8855);
nor U10120 (N_10120,N_8971,N_8821);
or U10121 (N_10121,N_9222,N_9355);
and U10122 (N_10122,N_8593,N_8546);
nand U10123 (N_10123,N_8886,N_9023);
or U10124 (N_10124,N_9064,N_9178);
and U10125 (N_10125,N_8979,N_8415);
nor U10126 (N_10126,N_8878,N_8661);
nand U10127 (N_10127,N_9297,N_9521);
nor U10128 (N_10128,N_9145,N_8738);
nand U10129 (N_10129,N_9148,N_8633);
nand U10130 (N_10130,N_9315,N_8525);
nand U10131 (N_10131,N_8714,N_9035);
nand U10132 (N_10132,N_8938,N_9186);
or U10133 (N_10133,N_8936,N_9299);
or U10134 (N_10134,N_9184,N_8736);
xor U10135 (N_10135,N_9378,N_8403);
nand U10136 (N_10136,N_8933,N_9081);
xnor U10137 (N_10137,N_8784,N_9172);
or U10138 (N_10138,N_9126,N_9528);
nor U10139 (N_10139,N_9497,N_9017);
or U10140 (N_10140,N_8817,N_9244);
nor U10141 (N_10141,N_8598,N_9293);
or U10142 (N_10142,N_9445,N_8790);
xor U10143 (N_10143,N_9327,N_9339);
and U10144 (N_10144,N_8669,N_8428);
nor U10145 (N_10145,N_8965,N_9082);
or U10146 (N_10146,N_8404,N_9514);
or U10147 (N_10147,N_9500,N_9033);
or U10148 (N_10148,N_9377,N_9594);
nand U10149 (N_10149,N_9542,N_9066);
and U10150 (N_10150,N_8869,N_8924);
and U10151 (N_10151,N_9411,N_8625);
nor U10152 (N_10152,N_9427,N_9137);
or U10153 (N_10153,N_9107,N_9466);
and U10154 (N_10154,N_8958,N_8444);
nand U10155 (N_10155,N_8753,N_8559);
xor U10156 (N_10156,N_9069,N_9270);
and U10157 (N_10157,N_8558,N_9063);
nor U10158 (N_10158,N_9385,N_9433);
xor U10159 (N_10159,N_9272,N_9463);
nor U10160 (N_10160,N_8660,N_8658);
and U10161 (N_10161,N_8976,N_8897);
or U10162 (N_10162,N_8505,N_8462);
nand U10163 (N_10163,N_8830,N_8646);
nor U10164 (N_10164,N_9344,N_8576);
or U10165 (N_10165,N_8850,N_9155);
and U10166 (N_10166,N_8402,N_8441);
nand U10167 (N_10167,N_8948,N_9298);
nand U10168 (N_10168,N_9196,N_9455);
nor U10169 (N_10169,N_8631,N_9441);
or U10170 (N_10170,N_9106,N_9051);
or U10171 (N_10171,N_8909,N_9276);
nand U10172 (N_10172,N_9523,N_9176);
nor U10173 (N_10173,N_9057,N_8839);
or U10174 (N_10174,N_9078,N_8972);
nor U10175 (N_10175,N_8667,N_8931);
xor U10176 (N_10176,N_9330,N_8967);
nor U10177 (N_10177,N_8500,N_8418);
xnor U10178 (N_10178,N_8468,N_8490);
nand U10179 (N_10179,N_9224,N_9370);
nor U10180 (N_10180,N_8430,N_9109);
xor U10181 (N_10181,N_9085,N_8517);
and U10182 (N_10182,N_9526,N_9146);
and U10183 (N_10183,N_8750,N_8841);
xnor U10184 (N_10184,N_9025,N_9380);
nand U10185 (N_10185,N_9169,N_9326);
xnor U10186 (N_10186,N_9028,N_8659);
nor U10187 (N_10187,N_9470,N_8763);
xnor U10188 (N_10188,N_8900,N_8513);
xnor U10189 (N_10189,N_8769,N_8480);
nand U10190 (N_10190,N_9366,N_9358);
xor U10191 (N_10191,N_9467,N_9454);
nand U10192 (N_10192,N_8779,N_8761);
nand U10193 (N_10193,N_8752,N_8510);
xor U10194 (N_10194,N_8526,N_8674);
or U10195 (N_10195,N_9185,N_8737);
nor U10196 (N_10196,N_9341,N_8543);
or U10197 (N_10197,N_9432,N_8810);
nand U10198 (N_10198,N_8456,N_8400);
xor U10199 (N_10199,N_8600,N_9310);
xor U10200 (N_10200,N_9009,N_8576);
nor U10201 (N_10201,N_8925,N_8618);
nor U10202 (N_10202,N_8979,N_8407);
nand U10203 (N_10203,N_8660,N_8749);
nor U10204 (N_10204,N_8540,N_8686);
nand U10205 (N_10205,N_8666,N_9040);
nor U10206 (N_10206,N_9536,N_9170);
and U10207 (N_10207,N_9207,N_8578);
or U10208 (N_10208,N_8517,N_8904);
nor U10209 (N_10209,N_8589,N_9322);
nor U10210 (N_10210,N_8874,N_9403);
or U10211 (N_10211,N_8486,N_9245);
nor U10212 (N_10212,N_8927,N_9070);
or U10213 (N_10213,N_8694,N_9092);
nand U10214 (N_10214,N_9427,N_9192);
xor U10215 (N_10215,N_9413,N_9422);
or U10216 (N_10216,N_9592,N_8848);
nor U10217 (N_10217,N_9380,N_8572);
nand U10218 (N_10218,N_9200,N_9525);
or U10219 (N_10219,N_8408,N_9038);
nand U10220 (N_10220,N_8503,N_9404);
nor U10221 (N_10221,N_9026,N_9268);
nand U10222 (N_10222,N_8539,N_9451);
or U10223 (N_10223,N_8798,N_9145);
xnor U10224 (N_10224,N_9349,N_8991);
xor U10225 (N_10225,N_8707,N_9144);
nor U10226 (N_10226,N_9123,N_8501);
nor U10227 (N_10227,N_8433,N_9158);
nor U10228 (N_10228,N_8599,N_9498);
or U10229 (N_10229,N_8408,N_9538);
nor U10230 (N_10230,N_9270,N_8906);
nand U10231 (N_10231,N_9219,N_9427);
nand U10232 (N_10232,N_9033,N_9190);
xnor U10233 (N_10233,N_9375,N_8704);
xor U10234 (N_10234,N_9072,N_8591);
nand U10235 (N_10235,N_9115,N_8667);
and U10236 (N_10236,N_9495,N_9460);
nand U10237 (N_10237,N_9588,N_8510);
or U10238 (N_10238,N_9046,N_9538);
nand U10239 (N_10239,N_9519,N_9351);
xor U10240 (N_10240,N_9132,N_8878);
nor U10241 (N_10241,N_9508,N_9001);
nor U10242 (N_10242,N_8731,N_9312);
and U10243 (N_10243,N_8842,N_8851);
nand U10244 (N_10244,N_8657,N_8492);
or U10245 (N_10245,N_8736,N_9202);
xor U10246 (N_10246,N_9466,N_9300);
nand U10247 (N_10247,N_8675,N_9274);
and U10248 (N_10248,N_8875,N_8446);
nor U10249 (N_10249,N_8650,N_9563);
and U10250 (N_10250,N_9015,N_9262);
and U10251 (N_10251,N_8551,N_8800);
xor U10252 (N_10252,N_9017,N_8599);
and U10253 (N_10253,N_8658,N_9252);
nor U10254 (N_10254,N_8502,N_9003);
and U10255 (N_10255,N_9388,N_8557);
nand U10256 (N_10256,N_8867,N_8663);
nor U10257 (N_10257,N_8875,N_8988);
nand U10258 (N_10258,N_9236,N_9199);
or U10259 (N_10259,N_9487,N_9363);
or U10260 (N_10260,N_9273,N_8633);
nand U10261 (N_10261,N_8648,N_8916);
or U10262 (N_10262,N_9455,N_8864);
nor U10263 (N_10263,N_9471,N_9596);
and U10264 (N_10264,N_9119,N_9276);
or U10265 (N_10265,N_9235,N_8725);
xnor U10266 (N_10266,N_9584,N_9169);
xnor U10267 (N_10267,N_9339,N_9441);
xor U10268 (N_10268,N_9574,N_8580);
or U10269 (N_10269,N_8627,N_9436);
nand U10270 (N_10270,N_9526,N_8525);
xnor U10271 (N_10271,N_9040,N_8844);
nor U10272 (N_10272,N_8407,N_9379);
or U10273 (N_10273,N_9155,N_8713);
nand U10274 (N_10274,N_9462,N_8480);
nor U10275 (N_10275,N_9427,N_9420);
and U10276 (N_10276,N_8719,N_8978);
and U10277 (N_10277,N_8895,N_8950);
and U10278 (N_10278,N_8774,N_8863);
xnor U10279 (N_10279,N_8737,N_8839);
or U10280 (N_10280,N_9433,N_8496);
or U10281 (N_10281,N_8811,N_8891);
or U10282 (N_10282,N_9351,N_8760);
and U10283 (N_10283,N_9127,N_9351);
nand U10284 (N_10284,N_8721,N_8416);
xor U10285 (N_10285,N_8728,N_8896);
nor U10286 (N_10286,N_9525,N_9570);
xor U10287 (N_10287,N_8889,N_9295);
and U10288 (N_10288,N_8820,N_8962);
nand U10289 (N_10289,N_8795,N_8722);
xnor U10290 (N_10290,N_8734,N_9178);
nand U10291 (N_10291,N_8400,N_8793);
nand U10292 (N_10292,N_9574,N_8819);
and U10293 (N_10293,N_9412,N_9520);
nor U10294 (N_10294,N_9222,N_8696);
or U10295 (N_10295,N_9147,N_9133);
nor U10296 (N_10296,N_8708,N_9542);
or U10297 (N_10297,N_9570,N_9127);
or U10298 (N_10298,N_8444,N_9353);
and U10299 (N_10299,N_8451,N_9586);
nor U10300 (N_10300,N_8757,N_8407);
xor U10301 (N_10301,N_9434,N_8883);
xnor U10302 (N_10302,N_9532,N_9133);
nand U10303 (N_10303,N_9465,N_8800);
xnor U10304 (N_10304,N_8943,N_8613);
and U10305 (N_10305,N_9307,N_9258);
nor U10306 (N_10306,N_9459,N_9592);
nor U10307 (N_10307,N_8564,N_8511);
and U10308 (N_10308,N_9321,N_9166);
or U10309 (N_10309,N_9043,N_8411);
and U10310 (N_10310,N_9327,N_9137);
or U10311 (N_10311,N_8963,N_9427);
nor U10312 (N_10312,N_8908,N_9252);
nor U10313 (N_10313,N_8843,N_9571);
and U10314 (N_10314,N_9295,N_9134);
nand U10315 (N_10315,N_8498,N_9015);
and U10316 (N_10316,N_8439,N_9456);
nand U10317 (N_10317,N_8569,N_8845);
and U10318 (N_10318,N_8896,N_8964);
and U10319 (N_10319,N_9367,N_8757);
nor U10320 (N_10320,N_9492,N_9106);
or U10321 (N_10321,N_8706,N_9486);
and U10322 (N_10322,N_9250,N_9517);
and U10323 (N_10323,N_9340,N_9341);
xnor U10324 (N_10324,N_9541,N_9514);
xor U10325 (N_10325,N_8662,N_9299);
and U10326 (N_10326,N_8468,N_9195);
or U10327 (N_10327,N_9407,N_8880);
and U10328 (N_10328,N_8609,N_8710);
xnor U10329 (N_10329,N_8634,N_8621);
and U10330 (N_10330,N_8872,N_9284);
nand U10331 (N_10331,N_8909,N_8602);
xor U10332 (N_10332,N_8500,N_9114);
nor U10333 (N_10333,N_8675,N_8812);
xor U10334 (N_10334,N_8828,N_8977);
and U10335 (N_10335,N_8692,N_9583);
nand U10336 (N_10336,N_9014,N_9171);
nand U10337 (N_10337,N_8526,N_8872);
or U10338 (N_10338,N_9561,N_8692);
xor U10339 (N_10339,N_9039,N_8554);
xor U10340 (N_10340,N_8765,N_9556);
nand U10341 (N_10341,N_8585,N_8857);
nor U10342 (N_10342,N_9226,N_8859);
xnor U10343 (N_10343,N_9060,N_9245);
xor U10344 (N_10344,N_8477,N_9059);
xor U10345 (N_10345,N_9193,N_8923);
xor U10346 (N_10346,N_9305,N_8691);
xor U10347 (N_10347,N_9442,N_9424);
nand U10348 (N_10348,N_8918,N_9381);
nand U10349 (N_10349,N_9020,N_9373);
nand U10350 (N_10350,N_9054,N_8920);
xnor U10351 (N_10351,N_9577,N_8488);
nor U10352 (N_10352,N_8898,N_8533);
and U10353 (N_10353,N_8891,N_8990);
xnor U10354 (N_10354,N_8766,N_8838);
or U10355 (N_10355,N_9543,N_9185);
nand U10356 (N_10356,N_8545,N_9036);
and U10357 (N_10357,N_9268,N_8969);
and U10358 (N_10358,N_8452,N_8555);
nor U10359 (N_10359,N_9278,N_8843);
nand U10360 (N_10360,N_9472,N_8545);
and U10361 (N_10361,N_9027,N_9280);
nor U10362 (N_10362,N_8797,N_8513);
nand U10363 (N_10363,N_8773,N_9459);
xor U10364 (N_10364,N_8500,N_9298);
xor U10365 (N_10365,N_8462,N_9217);
nor U10366 (N_10366,N_8476,N_8573);
xnor U10367 (N_10367,N_9247,N_9193);
xor U10368 (N_10368,N_9071,N_8603);
nor U10369 (N_10369,N_9436,N_8738);
nand U10370 (N_10370,N_8665,N_9351);
nand U10371 (N_10371,N_8895,N_8636);
or U10372 (N_10372,N_9320,N_8559);
nand U10373 (N_10373,N_8989,N_8571);
nor U10374 (N_10374,N_8915,N_8464);
nor U10375 (N_10375,N_9029,N_8713);
xor U10376 (N_10376,N_8966,N_8663);
or U10377 (N_10377,N_8937,N_8868);
or U10378 (N_10378,N_8981,N_9109);
nand U10379 (N_10379,N_9512,N_8958);
or U10380 (N_10380,N_8969,N_8989);
or U10381 (N_10381,N_8780,N_9420);
nor U10382 (N_10382,N_9220,N_8708);
or U10383 (N_10383,N_9393,N_8447);
xor U10384 (N_10384,N_8778,N_9385);
xor U10385 (N_10385,N_8443,N_8583);
xnor U10386 (N_10386,N_9008,N_9067);
xnor U10387 (N_10387,N_8793,N_9508);
or U10388 (N_10388,N_9089,N_9473);
xnor U10389 (N_10389,N_9097,N_9334);
nor U10390 (N_10390,N_8419,N_8576);
xor U10391 (N_10391,N_9137,N_8861);
or U10392 (N_10392,N_8869,N_8446);
nor U10393 (N_10393,N_9547,N_8855);
xor U10394 (N_10394,N_9145,N_8792);
xnor U10395 (N_10395,N_8509,N_9588);
xor U10396 (N_10396,N_9411,N_8956);
and U10397 (N_10397,N_9496,N_9228);
or U10398 (N_10398,N_8607,N_9441);
nand U10399 (N_10399,N_8569,N_9454);
nand U10400 (N_10400,N_8888,N_9399);
and U10401 (N_10401,N_9579,N_9095);
and U10402 (N_10402,N_8511,N_8759);
and U10403 (N_10403,N_8981,N_8984);
xor U10404 (N_10404,N_9325,N_9025);
nor U10405 (N_10405,N_9563,N_9456);
nor U10406 (N_10406,N_9080,N_8857);
and U10407 (N_10407,N_9101,N_8737);
and U10408 (N_10408,N_8504,N_9423);
or U10409 (N_10409,N_9390,N_8672);
nor U10410 (N_10410,N_9050,N_9523);
nor U10411 (N_10411,N_8687,N_9333);
or U10412 (N_10412,N_9059,N_9173);
xnor U10413 (N_10413,N_9450,N_9037);
and U10414 (N_10414,N_8686,N_8773);
nor U10415 (N_10415,N_9390,N_8984);
nand U10416 (N_10416,N_9166,N_9196);
and U10417 (N_10417,N_8809,N_8661);
or U10418 (N_10418,N_8432,N_9094);
nor U10419 (N_10419,N_8719,N_8950);
nor U10420 (N_10420,N_8552,N_9092);
and U10421 (N_10421,N_8732,N_9160);
or U10422 (N_10422,N_9054,N_9444);
or U10423 (N_10423,N_8871,N_9088);
xor U10424 (N_10424,N_9519,N_9330);
xor U10425 (N_10425,N_8966,N_8812);
and U10426 (N_10426,N_8604,N_9336);
nand U10427 (N_10427,N_8465,N_8791);
and U10428 (N_10428,N_9177,N_9163);
xnor U10429 (N_10429,N_8770,N_8738);
and U10430 (N_10430,N_9019,N_8780);
nor U10431 (N_10431,N_8808,N_8635);
nand U10432 (N_10432,N_9286,N_9481);
xnor U10433 (N_10433,N_8708,N_9036);
nand U10434 (N_10434,N_9151,N_9032);
and U10435 (N_10435,N_9554,N_8679);
nor U10436 (N_10436,N_9455,N_8763);
xnor U10437 (N_10437,N_9493,N_9541);
nand U10438 (N_10438,N_9398,N_8603);
nand U10439 (N_10439,N_9436,N_9453);
xor U10440 (N_10440,N_8735,N_9148);
nand U10441 (N_10441,N_9489,N_8831);
or U10442 (N_10442,N_8816,N_8625);
nand U10443 (N_10443,N_8943,N_9274);
and U10444 (N_10444,N_9569,N_9528);
or U10445 (N_10445,N_9413,N_8470);
xnor U10446 (N_10446,N_9134,N_8557);
xor U10447 (N_10447,N_9123,N_8995);
or U10448 (N_10448,N_9296,N_8427);
and U10449 (N_10449,N_9597,N_9499);
nor U10450 (N_10450,N_9576,N_8971);
xnor U10451 (N_10451,N_8417,N_9244);
nand U10452 (N_10452,N_8819,N_9056);
and U10453 (N_10453,N_9302,N_8564);
or U10454 (N_10454,N_8797,N_9462);
nand U10455 (N_10455,N_9481,N_9023);
or U10456 (N_10456,N_9398,N_8978);
or U10457 (N_10457,N_8728,N_9566);
or U10458 (N_10458,N_8538,N_8550);
nor U10459 (N_10459,N_9057,N_8560);
nor U10460 (N_10460,N_9486,N_9002);
and U10461 (N_10461,N_9502,N_8558);
and U10462 (N_10462,N_9378,N_8604);
nor U10463 (N_10463,N_8568,N_8825);
and U10464 (N_10464,N_8490,N_8549);
nor U10465 (N_10465,N_8923,N_8848);
xor U10466 (N_10466,N_9397,N_8968);
xor U10467 (N_10467,N_9377,N_9346);
nor U10468 (N_10468,N_9201,N_9014);
nand U10469 (N_10469,N_8925,N_8794);
or U10470 (N_10470,N_9151,N_9079);
nor U10471 (N_10471,N_9082,N_9103);
or U10472 (N_10472,N_8494,N_8552);
and U10473 (N_10473,N_8815,N_8788);
nand U10474 (N_10474,N_9418,N_9114);
nand U10475 (N_10475,N_9344,N_8873);
nand U10476 (N_10476,N_8598,N_9526);
and U10477 (N_10477,N_9545,N_8936);
or U10478 (N_10478,N_8528,N_9198);
xor U10479 (N_10479,N_9443,N_9174);
and U10480 (N_10480,N_9240,N_9147);
nor U10481 (N_10481,N_8836,N_9327);
or U10482 (N_10482,N_8747,N_9158);
and U10483 (N_10483,N_8648,N_8685);
nor U10484 (N_10484,N_9321,N_8745);
and U10485 (N_10485,N_8937,N_8802);
nand U10486 (N_10486,N_9287,N_8759);
nand U10487 (N_10487,N_9580,N_8929);
nand U10488 (N_10488,N_9597,N_8753);
or U10489 (N_10489,N_9320,N_8684);
nand U10490 (N_10490,N_9189,N_8578);
nand U10491 (N_10491,N_8631,N_8833);
and U10492 (N_10492,N_8539,N_8680);
nand U10493 (N_10493,N_9146,N_9103);
xnor U10494 (N_10494,N_9414,N_9197);
nand U10495 (N_10495,N_9362,N_8754);
xnor U10496 (N_10496,N_8419,N_9086);
and U10497 (N_10497,N_9132,N_9464);
and U10498 (N_10498,N_8940,N_9052);
xor U10499 (N_10499,N_8603,N_8610);
and U10500 (N_10500,N_9141,N_8813);
or U10501 (N_10501,N_9529,N_9385);
xnor U10502 (N_10502,N_8734,N_8710);
or U10503 (N_10503,N_8768,N_8412);
nand U10504 (N_10504,N_9313,N_9378);
nor U10505 (N_10505,N_9597,N_8807);
or U10506 (N_10506,N_9586,N_9022);
or U10507 (N_10507,N_9045,N_9241);
nor U10508 (N_10508,N_8796,N_8818);
nand U10509 (N_10509,N_8831,N_9364);
xnor U10510 (N_10510,N_8466,N_9119);
nand U10511 (N_10511,N_9024,N_9139);
nand U10512 (N_10512,N_8881,N_8506);
or U10513 (N_10513,N_9310,N_9271);
and U10514 (N_10514,N_9167,N_9163);
nor U10515 (N_10515,N_8528,N_8894);
nor U10516 (N_10516,N_8455,N_9119);
nand U10517 (N_10517,N_9421,N_9168);
and U10518 (N_10518,N_8469,N_9083);
nand U10519 (N_10519,N_9016,N_8929);
nand U10520 (N_10520,N_8780,N_9228);
xor U10521 (N_10521,N_9409,N_9203);
nor U10522 (N_10522,N_9123,N_8570);
and U10523 (N_10523,N_9220,N_9570);
nor U10524 (N_10524,N_9156,N_9472);
xor U10525 (N_10525,N_8481,N_8417);
and U10526 (N_10526,N_9190,N_9237);
nor U10527 (N_10527,N_8968,N_9471);
nand U10528 (N_10528,N_9379,N_8999);
nand U10529 (N_10529,N_8643,N_8844);
and U10530 (N_10530,N_8938,N_8467);
nor U10531 (N_10531,N_8869,N_9334);
and U10532 (N_10532,N_9400,N_9143);
nand U10533 (N_10533,N_9198,N_9147);
and U10534 (N_10534,N_8965,N_9404);
nor U10535 (N_10535,N_8499,N_8850);
and U10536 (N_10536,N_9043,N_8868);
nor U10537 (N_10537,N_8977,N_8903);
nand U10538 (N_10538,N_8758,N_8451);
nor U10539 (N_10539,N_9385,N_8409);
nor U10540 (N_10540,N_8615,N_8602);
xor U10541 (N_10541,N_9164,N_9309);
nor U10542 (N_10542,N_8542,N_8647);
xor U10543 (N_10543,N_9508,N_8652);
nor U10544 (N_10544,N_9423,N_9441);
and U10545 (N_10545,N_9134,N_8653);
and U10546 (N_10546,N_8417,N_8941);
xnor U10547 (N_10547,N_9363,N_9116);
xnor U10548 (N_10548,N_9251,N_9182);
and U10549 (N_10549,N_8606,N_8583);
nor U10550 (N_10550,N_9420,N_8982);
nand U10551 (N_10551,N_9361,N_8777);
nand U10552 (N_10552,N_8902,N_8712);
and U10553 (N_10553,N_8918,N_9525);
xnor U10554 (N_10554,N_8858,N_8556);
and U10555 (N_10555,N_8979,N_9065);
or U10556 (N_10556,N_9505,N_8653);
xor U10557 (N_10557,N_8530,N_8835);
and U10558 (N_10558,N_8640,N_8466);
nand U10559 (N_10559,N_9372,N_9438);
and U10560 (N_10560,N_8957,N_9067);
xnor U10561 (N_10561,N_8689,N_8819);
and U10562 (N_10562,N_8631,N_9549);
or U10563 (N_10563,N_8938,N_8781);
or U10564 (N_10564,N_8646,N_8451);
xnor U10565 (N_10565,N_8817,N_8781);
nand U10566 (N_10566,N_9197,N_8546);
or U10567 (N_10567,N_9434,N_8434);
or U10568 (N_10568,N_9389,N_8981);
and U10569 (N_10569,N_9353,N_9252);
or U10570 (N_10570,N_8744,N_8825);
xnor U10571 (N_10571,N_9408,N_9041);
nand U10572 (N_10572,N_8608,N_9211);
and U10573 (N_10573,N_8786,N_9185);
nor U10574 (N_10574,N_8466,N_8464);
and U10575 (N_10575,N_9490,N_8598);
xor U10576 (N_10576,N_8945,N_9568);
and U10577 (N_10577,N_8794,N_8440);
and U10578 (N_10578,N_9296,N_9422);
xor U10579 (N_10579,N_8777,N_9585);
or U10580 (N_10580,N_8597,N_8543);
or U10581 (N_10581,N_8693,N_9579);
nand U10582 (N_10582,N_9547,N_8415);
nand U10583 (N_10583,N_9143,N_9024);
or U10584 (N_10584,N_9249,N_8617);
xor U10585 (N_10585,N_8440,N_8682);
nand U10586 (N_10586,N_9072,N_9009);
nor U10587 (N_10587,N_8779,N_9227);
and U10588 (N_10588,N_8424,N_8404);
nand U10589 (N_10589,N_9141,N_9076);
or U10590 (N_10590,N_8673,N_9373);
or U10591 (N_10591,N_9160,N_8958);
nor U10592 (N_10592,N_8525,N_9220);
and U10593 (N_10593,N_8512,N_8681);
and U10594 (N_10594,N_9059,N_9230);
nand U10595 (N_10595,N_9462,N_8862);
and U10596 (N_10596,N_9481,N_9445);
xnor U10597 (N_10597,N_9417,N_9442);
nand U10598 (N_10598,N_9368,N_8637);
and U10599 (N_10599,N_8589,N_9421);
nand U10600 (N_10600,N_9010,N_9362);
xor U10601 (N_10601,N_9081,N_9533);
and U10602 (N_10602,N_9145,N_8771);
or U10603 (N_10603,N_8654,N_8551);
xor U10604 (N_10604,N_8740,N_9507);
xor U10605 (N_10605,N_9082,N_8685);
xnor U10606 (N_10606,N_8575,N_9208);
nand U10607 (N_10607,N_9520,N_8708);
or U10608 (N_10608,N_8808,N_9267);
nand U10609 (N_10609,N_9165,N_8409);
nor U10610 (N_10610,N_8650,N_8560);
xnor U10611 (N_10611,N_8760,N_9348);
or U10612 (N_10612,N_9031,N_9069);
xor U10613 (N_10613,N_9347,N_9386);
and U10614 (N_10614,N_9250,N_9305);
nor U10615 (N_10615,N_9460,N_9274);
and U10616 (N_10616,N_8664,N_9055);
and U10617 (N_10617,N_9578,N_8643);
nor U10618 (N_10618,N_8506,N_8801);
xnor U10619 (N_10619,N_9086,N_8955);
and U10620 (N_10620,N_8502,N_9025);
nor U10621 (N_10621,N_9265,N_8438);
nand U10622 (N_10622,N_9434,N_8583);
nor U10623 (N_10623,N_9341,N_8691);
nand U10624 (N_10624,N_8732,N_8685);
and U10625 (N_10625,N_9476,N_9211);
xor U10626 (N_10626,N_9156,N_9432);
nand U10627 (N_10627,N_8882,N_8809);
or U10628 (N_10628,N_8938,N_8995);
or U10629 (N_10629,N_9271,N_8872);
and U10630 (N_10630,N_8445,N_9527);
nand U10631 (N_10631,N_8507,N_9268);
nand U10632 (N_10632,N_8743,N_8672);
nor U10633 (N_10633,N_8841,N_9301);
xnor U10634 (N_10634,N_9592,N_9413);
and U10635 (N_10635,N_9419,N_8573);
nor U10636 (N_10636,N_8575,N_9244);
xnor U10637 (N_10637,N_9408,N_8633);
nor U10638 (N_10638,N_9407,N_9380);
and U10639 (N_10639,N_8929,N_9545);
or U10640 (N_10640,N_8733,N_8538);
and U10641 (N_10641,N_8864,N_9348);
or U10642 (N_10642,N_9186,N_9040);
nor U10643 (N_10643,N_9321,N_9470);
and U10644 (N_10644,N_8448,N_9397);
nor U10645 (N_10645,N_9040,N_8870);
xor U10646 (N_10646,N_8660,N_9300);
xor U10647 (N_10647,N_9057,N_8786);
and U10648 (N_10648,N_8714,N_8583);
xnor U10649 (N_10649,N_9439,N_9365);
or U10650 (N_10650,N_9592,N_9432);
nand U10651 (N_10651,N_9202,N_9341);
nand U10652 (N_10652,N_8475,N_8470);
nand U10653 (N_10653,N_9462,N_9253);
xnor U10654 (N_10654,N_8831,N_8881);
nand U10655 (N_10655,N_9473,N_8760);
nand U10656 (N_10656,N_9103,N_9153);
or U10657 (N_10657,N_9198,N_9061);
nor U10658 (N_10658,N_9076,N_8804);
xor U10659 (N_10659,N_8788,N_8464);
xnor U10660 (N_10660,N_9046,N_8816);
nand U10661 (N_10661,N_9269,N_8598);
nand U10662 (N_10662,N_8477,N_8488);
nand U10663 (N_10663,N_8887,N_8574);
nor U10664 (N_10664,N_9567,N_9069);
nand U10665 (N_10665,N_8582,N_9384);
nand U10666 (N_10666,N_9103,N_9489);
or U10667 (N_10667,N_9556,N_9457);
xnor U10668 (N_10668,N_8830,N_9461);
nor U10669 (N_10669,N_9149,N_9561);
xor U10670 (N_10670,N_8847,N_8447);
nor U10671 (N_10671,N_8976,N_8674);
nor U10672 (N_10672,N_8429,N_9551);
nand U10673 (N_10673,N_8686,N_8427);
nand U10674 (N_10674,N_9252,N_9304);
nand U10675 (N_10675,N_8832,N_8735);
or U10676 (N_10676,N_9437,N_8867);
and U10677 (N_10677,N_8453,N_8929);
xnor U10678 (N_10678,N_8779,N_9453);
nand U10679 (N_10679,N_8625,N_9484);
and U10680 (N_10680,N_8881,N_8500);
or U10681 (N_10681,N_9417,N_8875);
nand U10682 (N_10682,N_9387,N_9038);
nand U10683 (N_10683,N_9087,N_8714);
and U10684 (N_10684,N_8549,N_9357);
and U10685 (N_10685,N_9306,N_8537);
nor U10686 (N_10686,N_9123,N_8580);
nor U10687 (N_10687,N_9048,N_8913);
xor U10688 (N_10688,N_9556,N_8449);
nand U10689 (N_10689,N_8871,N_8454);
nor U10690 (N_10690,N_9518,N_9199);
or U10691 (N_10691,N_8422,N_9338);
nand U10692 (N_10692,N_9052,N_9395);
nand U10693 (N_10693,N_8678,N_8934);
nor U10694 (N_10694,N_9120,N_8531);
and U10695 (N_10695,N_9539,N_8447);
or U10696 (N_10696,N_8413,N_9261);
or U10697 (N_10697,N_9256,N_9513);
and U10698 (N_10698,N_8567,N_8707);
nand U10699 (N_10699,N_9275,N_9145);
xnor U10700 (N_10700,N_8923,N_8858);
or U10701 (N_10701,N_9246,N_8810);
and U10702 (N_10702,N_9135,N_9478);
nor U10703 (N_10703,N_9432,N_8820);
xor U10704 (N_10704,N_8705,N_9125);
nand U10705 (N_10705,N_8933,N_9277);
nand U10706 (N_10706,N_9486,N_9302);
and U10707 (N_10707,N_9312,N_8596);
nand U10708 (N_10708,N_8456,N_8580);
and U10709 (N_10709,N_8641,N_9499);
xnor U10710 (N_10710,N_9420,N_9443);
nand U10711 (N_10711,N_8912,N_9187);
or U10712 (N_10712,N_8725,N_9244);
nand U10713 (N_10713,N_9405,N_8755);
or U10714 (N_10714,N_8531,N_8853);
nand U10715 (N_10715,N_8931,N_9434);
xor U10716 (N_10716,N_8880,N_8426);
nor U10717 (N_10717,N_8792,N_9599);
and U10718 (N_10718,N_8866,N_9336);
and U10719 (N_10719,N_8820,N_8716);
nor U10720 (N_10720,N_8953,N_9325);
nor U10721 (N_10721,N_8508,N_8541);
or U10722 (N_10722,N_8518,N_8960);
nor U10723 (N_10723,N_8996,N_9400);
nor U10724 (N_10724,N_9585,N_8737);
nor U10725 (N_10725,N_9132,N_9444);
nor U10726 (N_10726,N_9404,N_9122);
or U10727 (N_10727,N_9284,N_8480);
nor U10728 (N_10728,N_8435,N_9222);
nand U10729 (N_10729,N_8810,N_9206);
nor U10730 (N_10730,N_8833,N_8494);
or U10731 (N_10731,N_9005,N_9109);
xnor U10732 (N_10732,N_8731,N_8431);
or U10733 (N_10733,N_9003,N_9294);
or U10734 (N_10734,N_8551,N_9336);
nand U10735 (N_10735,N_9428,N_8984);
or U10736 (N_10736,N_8788,N_8501);
xor U10737 (N_10737,N_8952,N_9232);
nor U10738 (N_10738,N_9371,N_8432);
and U10739 (N_10739,N_9080,N_8494);
xor U10740 (N_10740,N_9369,N_8709);
or U10741 (N_10741,N_8744,N_9351);
nand U10742 (N_10742,N_9389,N_8824);
xnor U10743 (N_10743,N_9039,N_8766);
nor U10744 (N_10744,N_9366,N_9064);
nor U10745 (N_10745,N_9416,N_8732);
xor U10746 (N_10746,N_9168,N_8516);
xor U10747 (N_10747,N_8936,N_9352);
or U10748 (N_10748,N_8905,N_9576);
nand U10749 (N_10749,N_9313,N_8872);
and U10750 (N_10750,N_9035,N_9287);
nand U10751 (N_10751,N_8515,N_9435);
nand U10752 (N_10752,N_9376,N_9562);
and U10753 (N_10753,N_8605,N_9593);
nand U10754 (N_10754,N_9222,N_9108);
nand U10755 (N_10755,N_9358,N_9229);
xor U10756 (N_10756,N_9575,N_8446);
nor U10757 (N_10757,N_9369,N_9255);
or U10758 (N_10758,N_9393,N_9515);
nand U10759 (N_10759,N_9043,N_8598);
xnor U10760 (N_10760,N_8587,N_9340);
nand U10761 (N_10761,N_8784,N_8842);
xnor U10762 (N_10762,N_9189,N_8986);
or U10763 (N_10763,N_8722,N_8433);
or U10764 (N_10764,N_9541,N_8870);
xor U10765 (N_10765,N_8506,N_9068);
or U10766 (N_10766,N_8584,N_9268);
or U10767 (N_10767,N_9231,N_8775);
nor U10768 (N_10768,N_8517,N_9285);
nor U10769 (N_10769,N_9538,N_8959);
nand U10770 (N_10770,N_8846,N_9153);
nand U10771 (N_10771,N_9411,N_9208);
nand U10772 (N_10772,N_8461,N_9199);
or U10773 (N_10773,N_8487,N_8626);
and U10774 (N_10774,N_8695,N_8592);
and U10775 (N_10775,N_9386,N_9352);
nor U10776 (N_10776,N_9189,N_9597);
nor U10777 (N_10777,N_8627,N_9218);
nand U10778 (N_10778,N_9560,N_8658);
or U10779 (N_10779,N_9258,N_9025);
nand U10780 (N_10780,N_8585,N_9176);
and U10781 (N_10781,N_8868,N_8582);
nand U10782 (N_10782,N_9519,N_9064);
xnor U10783 (N_10783,N_8541,N_8992);
and U10784 (N_10784,N_9168,N_8694);
xor U10785 (N_10785,N_8768,N_9584);
xnor U10786 (N_10786,N_9482,N_8495);
nor U10787 (N_10787,N_9012,N_9429);
or U10788 (N_10788,N_9263,N_8642);
xnor U10789 (N_10789,N_9124,N_8977);
and U10790 (N_10790,N_8731,N_9556);
nand U10791 (N_10791,N_9344,N_8727);
and U10792 (N_10792,N_8505,N_8875);
or U10793 (N_10793,N_9507,N_8927);
or U10794 (N_10794,N_9321,N_9506);
or U10795 (N_10795,N_9126,N_8758);
xor U10796 (N_10796,N_8835,N_9269);
nor U10797 (N_10797,N_8776,N_8503);
nand U10798 (N_10798,N_8562,N_8816);
or U10799 (N_10799,N_8507,N_9198);
xor U10800 (N_10800,N_9879,N_9704);
nand U10801 (N_10801,N_10402,N_9712);
and U10802 (N_10802,N_9745,N_10584);
or U10803 (N_10803,N_10091,N_9648);
and U10804 (N_10804,N_10775,N_9770);
xnor U10805 (N_10805,N_9881,N_9794);
nand U10806 (N_10806,N_9996,N_9692);
and U10807 (N_10807,N_10772,N_10532);
nand U10808 (N_10808,N_9743,N_10347);
xnor U10809 (N_10809,N_10266,N_10469);
xnor U10810 (N_10810,N_10499,N_10278);
and U10811 (N_10811,N_10738,N_10484);
xor U10812 (N_10812,N_10729,N_9840);
xor U10813 (N_10813,N_10442,N_10130);
xnor U10814 (N_10814,N_10166,N_10217);
or U10815 (N_10815,N_10700,N_9889);
nor U10816 (N_10816,N_10142,N_10722);
and U10817 (N_10817,N_10099,N_9867);
nor U10818 (N_10818,N_9786,N_9863);
xnor U10819 (N_10819,N_10560,N_10631);
nor U10820 (N_10820,N_10026,N_9857);
or U10821 (N_10821,N_9781,N_10332);
xnor U10822 (N_10822,N_10602,N_10762);
nand U10823 (N_10823,N_10500,N_10032);
or U10824 (N_10824,N_9731,N_9732);
nand U10825 (N_10825,N_10765,N_10301);
nand U10826 (N_10826,N_10497,N_10521);
xor U10827 (N_10827,N_10557,N_9640);
nand U10828 (N_10828,N_9870,N_10368);
nor U10829 (N_10829,N_9662,N_10465);
or U10830 (N_10830,N_9850,N_10637);
or U10831 (N_10831,N_10248,N_10022);
xor U10832 (N_10832,N_9896,N_10378);
and U10833 (N_10833,N_10669,N_9807);
and U10834 (N_10834,N_10671,N_10651);
xnor U10835 (N_10835,N_10229,N_10744);
xnor U10836 (N_10836,N_9902,N_10286);
nand U10837 (N_10837,N_10512,N_10116);
nand U10838 (N_10838,N_9943,N_9631);
or U10839 (N_10839,N_9971,N_9792);
nand U10840 (N_10840,N_10698,N_9940);
or U10841 (N_10841,N_9643,N_10231);
nand U10842 (N_10842,N_9811,N_10134);
nor U10843 (N_10843,N_10063,N_10333);
nand U10844 (N_10844,N_9929,N_10405);
xor U10845 (N_10845,N_10413,N_9769);
or U10846 (N_10846,N_10783,N_9819);
nand U10847 (N_10847,N_10473,N_10764);
xnor U10848 (N_10848,N_10177,N_10420);
xnor U10849 (N_10849,N_10639,N_10244);
xnor U10850 (N_10850,N_10159,N_9644);
nor U10851 (N_10851,N_10003,N_10119);
nor U10852 (N_10852,N_10542,N_10553);
nand U10853 (N_10853,N_10054,N_10516);
nand U10854 (N_10854,N_10567,N_10001);
xor U10855 (N_10855,N_10184,N_10580);
xor U10856 (N_10856,N_10093,N_9854);
or U10857 (N_10857,N_9734,N_10665);
nor U10858 (N_10858,N_9744,N_10260);
xnor U10859 (N_10859,N_10436,N_10150);
and U10860 (N_10860,N_10431,N_10559);
or U10861 (N_10861,N_10742,N_10658);
and U10862 (N_10862,N_10132,N_10704);
xor U10863 (N_10863,N_9768,N_10523);
nor U10864 (N_10864,N_9754,N_9873);
xnor U10865 (N_10865,N_10741,N_10520);
or U10866 (N_10866,N_10797,N_10190);
and U10867 (N_10867,N_10207,N_10642);
and U10868 (N_10868,N_9829,N_10398);
nor U10869 (N_10869,N_10292,N_10196);
or U10870 (N_10870,N_10392,N_10691);
xor U10871 (N_10871,N_9703,N_10287);
xnor U10872 (N_10872,N_9671,N_10007);
or U10873 (N_10873,N_10156,N_10135);
nor U10874 (N_10874,N_9755,N_9664);
or U10875 (N_10875,N_10182,N_9893);
xor U10876 (N_10876,N_10483,N_10787);
or U10877 (N_10877,N_10176,N_9606);
and U10878 (N_10878,N_10302,N_10218);
nor U10879 (N_10879,N_10367,N_10450);
or U10880 (N_10880,N_10443,N_10318);
or U10881 (N_10881,N_10048,N_9605);
and U10882 (N_10882,N_9942,N_9908);
xor U10883 (N_10883,N_10137,N_10654);
xor U10884 (N_10884,N_10299,N_10566);
nand U10885 (N_10885,N_9735,N_10718);
xor U10886 (N_10886,N_10033,N_10234);
and U10887 (N_10887,N_10608,N_9696);
nand U10888 (N_10888,N_9956,N_10065);
or U10889 (N_10889,N_9772,N_9787);
and U10890 (N_10890,N_10322,N_10243);
and U10891 (N_10891,N_10617,N_9953);
and U10892 (N_10892,N_10627,N_10240);
xnor U10893 (N_10893,N_10501,N_10437);
nor U10894 (N_10894,N_10111,N_10004);
nor U10895 (N_10895,N_10423,N_9773);
and U10896 (N_10896,N_10364,N_10352);
and U10897 (N_10897,N_9615,N_9777);
or U10898 (N_10898,N_10650,N_9888);
or U10899 (N_10899,N_10416,N_10538);
nor U10900 (N_10900,N_9668,N_10160);
and U10901 (N_10901,N_10222,N_10289);
or U10902 (N_10902,N_9721,N_9900);
xor U10903 (N_10903,N_10399,N_10635);
nor U10904 (N_10904,N_9834,N_10548);
xor U10905 (N_10905,N_10746,N_10038);
or U10906 (N_10906,N_10327,N_9730);
or U10907 (N_10907,N_9860,N_9844);
nor U10908 (N_10908,N_9613,N_9812);
or U10909 (N_10909,N_9765,N_9973);
nor U10910 (N_10910,N_10268,N_10601);
nand U10911 (N_10911,N_10773,N_10097);
nand U10912 (N_10912,N_10027,N_10664);
or U10913 (N_10913,N_9915,N_10355);
or U10914 (N_10914,N_10334,N_10254);
and U10915 (N_10915,N_10146,N_10149);
nand U10916 (N_10916,N_9992,N_10165);
or U10917 (N_10917,N_10181,N_9793);
nor U10918 (N_10918,N_9959,N_10070);
or U10919 (N_10919,N_10689,N_10776);
xor U10920 (N_10920,N_9666,N_10264);
and U10921 (N_10921,N_10466,N_9716);
and U10922 (N_10922,N_10171,N_9823);
nand U10923 (N_10923,N_10707,N_9747);
and U10924 (N_10924,N_10572,N_10319);
xnor U10925 (N_10925,N_10373,N_10793);
nand U10926 (N_10926,N_9691,N_10767);
xnor U10927 (N_10927,N_10585,N_9837);
nand U10928 (N_10928,N_10663,N_10481);
xnor U10929 (N_10929,N_10730,N_10646);
and U10930 (N_10930,N_9861,N_10710);
xor U10931 (N_10931,N_9993,N_9830);
nor U10932 (N_10932,N_10056,N_9906);
xnor U10933 (N_10933,N_9872,N_9907);
nand U10934 (N_10934,N_9767,N_10300);
and U10935 (N_10935,N_10779,N_9763);
nand U10936 (N_10936,N_9986,N_9928);
xor U10937 (N_10937,N_10147,N_10396);
or U10938 (N_10938,N_9707,N_10652);
xnor U10939 (N_10939,N_10647,N_10385);
nand U10940 (N_10940,N_9690,N_10514);
nor U10941 (N_10941,N_9706,N_10384);
nor U10942 (N_10942,N_9980,N_10183);
or U10943 (N_10943,N_10628,N_10692);
nand U10944 (N_10944,N_9880,N_9693);
and U10945 (N_10945,N_9848,N_9816);
nand U10946 (N_10946,N_10439,N_9877);
nor U10947 (N_10947,N_10587,N_10502);
or U10948 (N_10948,N_10204,N_10331);
or U10949 (N_10949,N_10417,N_10382);
or U10950 (N_10950,N_10645,N_10276);
and U10951 (N_10951,N_10239,N_9783);
nor U10952 (N_10952,N_10518,N_10238);
nor U10953 (N_10953,N_10379,N_10510);
xor U10954 (N_10954,N_10257,N_10008);
and U10955 (N_10955,N_9627,N_10386);
xor U10956 (N_10956,N_9689,N_10073);
xnor U10957 (N_10957,N_9701,N_9798);
nand U10958 (N_10958,N_10100,N_10269);
xor U10959 (N_10959,N_9874,N_10090);
nor U10960 (N_10960,N_10479,N_10085);
xor U10961 (N_10961,N_10412,N_9602);
xor U10962 (N_10962,N_10154,N_10258);
nor U10963 (N_10963,N_9795,N_10640);
or U10964 (N_10964,N_9739,N_9868);
nor U10965 (N_10965,N_9626,N_10155);
or U10966 (N_10966,N_10297,N_9717);
nand U10967 (N_10967,N_9601,N_9875);
nor U10968 (N_10968,N_10788,N_10072);
xnor U10969 (N_10969,N_9898,N_10380);
or U10970 (N_10970,N_10115,N_9618);
xnor U10971 (N_10971,N_10720,N_10095);
or U10972 (N_10972,N_10068,N_10513);
or U10973 (N_10973,N_10603,N_9727);
and U10974 (N_10974,N_10066,N_10002);
xnor U10975 (N_10975,N_10325,N_9709);
nand U10976 (N_10976,N_10113,N_10360);
nor U10977 (N_10977,N_9964,N_9923);
nor U10978 (N_10978,N_9612,N_9651);
xnor U10979 (N_10979,N_9858,N_10748);
and U10980 (N_10980,N_9920,N_9610);
nand U10981 (N_10981,N_10010,N_10271);
nor U10982 (N_10982,N_10487,N_10724);
nor U10983 (N_10983,N_10711,N_10426);
nand U10984 (N_10984,N_9890,N_10476);
or U10985 (N_10985,N_9634,N_10213);
or U10986 (N_10986,N_10285,N_9660);
or U10987 (N_10987,N_10141,N_9657);
or U10988 (N_10988,N_10547,N_10434);
and U10989 (N_10989,N_10583,N_9912);
or U10990 (N_10990,N_9820,N_10697);
nor U10991 (N_10991,N_10610,N_9977);
or U10992 (N_10992,N_9897,N_10064);
nor U10993 (N_10993,N_10577,N_9698);
nor U10994 (N_10994,N_9839,N_9815);
nor U10995 (N_10995,N_10662,N_9936);
or U10996 (N_10996,N_10158,N_9825);
nand U10997 (N_10997,N_9608,N_9913);
or U10998 (N_10998,N_10758,N_9904);
xor U10999 (N_10999,N_9683,N_10098);
xnor U11000 (N_11000,N_9699,N_9742);
or U11001 (N_11001,N_10388,N_10112);
nor U11002 (N_11002,N_9617,N_10754);
nor U11003 (N_11003,N_9632,N_10133);
or U11004 (N_11004,N_9686,N_9728);
or U11005 (N_11005,N_9740,N_10556);
and U11006 (N_11006,N_10723,N_10528);
xor U11007 (N_11007,N_10127,N_10312);
xor U11008 (N_11008,N_9984,N_10125);
or U11009 (N_11009,N_9982,N_10050);
xor U11010 (N_11010,N_10363,N_9841);
xnor U11011 (N_11011,N_10202,N_9822);
nand U11012 (N_11012,N_10798,N_10452);
nor U11013 (N_11013,N_10415,N_10470);
xor U11014 (N_11014,N_9905,N_10592);
or U11015 (N_11015,N_9925,N_10667);
xor U11016 (N_11016,N_10209,N_10504);
or U11017 (N_11017,N_9719,N_9779);
or U11018 (N_11018,N_10590,N_10612);
and U11019 (N_11019,N_10283,N_9711);
or U11020 (N_11020,N_10794,N_9609);
nand U11021 (N_11021,N_10699,N_10259);
or U11022 (N_11022,N_10023,N_9994);
nor U11023 (N_11023,N_10406,N_9974);
or U11024 (N_11024,N_9970,N_10565);
or U11025 (N_11025,N_10727,N_9921);
nor U11026 (N_11026,N_10421,N_10461);
and U11027 (N_11027,N_10533,N_10227);
xnor U11028 (N_11028,N_10422,N_10435);
and U11029 (N_11029,N_10397,N_10079);
xnor U11030 (N_11030,N_10551,N_10344);
xor U11031 (N_11031,N_10638,N_10526);
xor U11032 (N_11032,N_10685,N_10371);
and U11033 (N_11033,N_10148,N_10449);
xnor U11034 (N_11034,N_9780,N_9814);
or U11035 (N_11035,N_10366,N_10770);
nand U11036 (N_11036,N_10161,N_10145);
xor U11037 (N_11037,N_9673,N_9737);
nand U11038 (N_11038,N_10677,N_10404);
and U11039 (N_11039,N_10537,N_10763);
or U11040 (N_11040,N_10107,N_9990);
nand U11041 (N_11041,N_10686,N_10725);
nor U11042 (N_11042,N_9797,N_10527);
xnor U11043 (N_11043,N_9947,N_9979);
and U11044 (N_11044,N_10361,N_10558);
and U11045 (N_11045,N_10530,N_10769);
xor U11046 (N_11046,N_9941,N_9883);
xnor U11047 (N_11047,N_10309,N_10236);
nand U11048 (N_11048,N_9991,N_10524);
nor U11049 (N_11049,N_10562,N_9955);
and U11050 (N_11050,N_10294,N_9661);
xnor U11051 (N_11051,N_10784,N_10430);
nor U11052 (N_11052,N_10569,N_9778);
nand U11053 (N_11053,N_10338,N_10489);
or U11054 (N_11054,N_10792,N_10340);
and U11055 (N_11055,N_10216,N_10785);
xor U11056 (N_11056,N_9948,N_10045);
xnor U11057 (N_11057,N_10401,N_9914);
nand U11058 (N_11058,N_10534,N_9946);
xor U11059 (N_11059,N_9876,N_10307);
xnor U11060 (N_11060,N_10205,N_10478);
xor U11061 (N_11061,N_10136,N_10349);
nand U11062 (N_11062,N_9639,N_10211);
or U11063 (N_11063,N_9659,N_10057);
xor U11064 (N_11064,N_10101,N_10543);
or U11065 (N_11065,N_10621,N_10120);
xor U11066 (N_11066,N_10224,N_10721);
nand U11067 (N_11067,N_10626,N_9957);
nand U11068 (N_11068,N_10105,N_9852);
nand U11069 (N_11069,N_10212,N_10680);
xor U11070 (N_11070,N_10082,N_10611);
nor U11071 (N_11071,N_10242,N_10458);
and U11072 (N_11072,N_10108,N_9909);
nand U11073 (N_11073,N_10365,N_9865);
and U11074 (N_11074,N_10317,N_10006);
nor U11075 (N_11075,N_10314,N_10357);
or U11076 (N_11076,N_9851,N_10594);
and U11077 (N_11077,N_9855,N_10353);
nand U11078 (N_11078,N_10372,N_9718);
xor U11079 (N_11079,N_10732,N_9759);
or U11080 (N_11080,N_10529,N_9903);
and U11081 (N_11081,N_10702,N_10606);
nand U11082 (N_11082,N_10480,N_10288);
nor U11083 (N_11083,N_10624,N_10106);
and U11084 (N_11084,N_10076,N_10376);
nand U11085 (N_11085,N_9654,N_10246);
or U11086 (N_11086,N_10153,N_10736);
nand U11087 (N_11087,N_9918,N_9931);
and U11088 (N_11088,N_10522,N_9636);
nand U11089 (N_11089,N_9824,N_9945);
or U11090 (N_11090,N_10012,N_10315);
and U11091 (N_11091,N_9887,N_10778);
xnor U11092 (N_11092,N_10273,N_10109);
nor U11093 (N_11093,N_10467,N_10745);
or U11094 (N_11094,N_10274,N_10561);
xnor U11095 (N_11095,N_9746,N_10102);
nand U11096 (N_11096,N_9658,N_9997);
nand U11097 (N_11097,N_9916,N_10028);
nand U11098 (N_11098,N_10495,N_10221);
nand U11099 (N_11099,N_9622,N_9968);
xnor U11100 (N_11100,N_10061,N_9620);
nand U11101 (N_11101,N_9776,N_9619);
xor U11102 (N_11102,N_10418,N_10016);
xor U11103 (N_11103,N_9607,N_10320);
or U11104 (N_11104,N_10630,N_10117);
nand U11105 (N_11105,N_10174,N_10080);
and U11106 (N_11106,N_10053,N_10672);
and U11107 (N_11107,N_10474,N_9761);
or U11108 (N_11108,N_10345,N_10199);
and U11109 (N_11109,N_10343,N_10506);
and U11110 (N_11110,N_10081,N_9714);
and U11111 (N_11111,N_9774,N_10069);
nor U11112 (N_11112,N_10613,N_10539);
and U11113 (N_11113,N_9821,N_10573);
nor U11114 (N_11114,N_10241,N_9645);
or U11115 (N_11115,N_9641,N_9702);
and U11116 (N_11116,N_10280,N_10498);
nand U11117 (N_11117,N_10040,N_10129);
nor U11118 (N_11118,N_9764,N_10261);
nor U11119 (N_11119,N_9987,N_9842);
nand U11120 (N_11120,N_10164,N_10716);
nor U11121 (N_11121,N_10042,N_10578);
or U11122 (N_11122,N_10409,N_10037);
and U11123 (N_11123,N_9804,N_10550);
and U11124 (N_11124,N_10508,N_10139);
xor U11125 (N_11125,N_10535,N_10089);
xnor U11126 (N_11126,N_10179,N_9625);
or U11127 (N_11127,N_10735,N_10428);
nand U11128 (N_11128,N_9911,N_10673);
or U11129 (N_11129,N_10708,N_10296);
xor U11130 (N_11130,N_10503,N_10679);
or U11131 (N_11131,N_10761,N_10600);
nand U11132 (N_11132,N_10214,N_10751);
nand U11133 (N_11133,N_10641,N_10362);
xnor U11134 (N_11134,N_9813,N_10219);
nor U11135 (N_11135,N_9655,N_10486);
and U11136 (N_11136,N_10438,N_9782);
xnor U11137 (N_11137,N_10634,N_10310);
and U11138 (N_11138,N_9801,N_10393);
xnor U11139 (N_11139,N_10693,N_10541);
or U11140 (N_11140,N_10247,N_9790);
nor U11141 (N_11141,N_10615,N_10011);
and U11142 (N_11142,N_10563,N_10387);
or U11143 (N_11143,N_9808,N_10144);
xnor U11144 (N_11144,N_9800,N_9736);
nor U11145 (N_11145,N_10575,N_10305);
xnor U11146 (N_11146,N_10041,N_9802);
nand U11147 (N_11147,N_10690,N_9669);
or U11148 (N_11148,N_9628,N_10643);
xor U11149 (N_11149,N_9674,N_10737);
and U11150 (N_11150,N_10351,N_10451);
nand U11151 (N_11151,N_10370,N_10195);
nor U11152 (N_11152,N_9845,N_10756);
and U11153 (N_11153,N_10021,N_10311);
or U11154 (N_11154,N_10703,N_10786);
or U11155 (N_11155,N_10123,N_10509);
nor U11156 (N_11156,N_9952,N_10799);
nor U11157 (N_11157,N_9944,N_9679);
nor U11158 (N_11158,N_10014,N_10705);
nor U11159 (N_11159,N_10168,N_10715);
nor U11160 (N_11160,N_10570,N_9999);
nand U11161 (N_11161,N_10607,N_10094);
and U11162 (N_11162,N_9705,N_9653);
nor U11163 (N_11163,N_10574,N_9843);
nor U11164 (N_11164,N_9919,N_10471);
xnor U11165 (N_11165,N_10281,N_10517);
nor U11166 (N_11166,N_10226,N_10675);
xor U11167 (N_11167,N_10688,N_10230);
nand U11168 (N_11168,N_10713,N_10448);
or U11169 (N_11169,N_9624,N_10284);
xnor U11170 (N_11170,N_9775,N_10348);
or U11171 (N_11171,N_10381,N_9884);
xor U11172 (N_11172,N_9939,N_10411);
nor U11173 (N_11173,N_10337,N_9616);
and U11174 (N_11174,N_10389,N_9937);
and U11175 (N_11175,N_10649,N_10103);
or U11176 (N_11176,N_10187,N_10395);
and U11177 (N_11177,N_10425,N_10734);
nand U11178 (N_11178,N_10043,N_9809);
or U11179 (N_11179,N_9985,N_9961);
nand U11180 (N_11180,N_9603,N_9988);
nor U11181 (N_11181,N_9933,N_10225);
xnor U11182 (N_11182,N_10203,N_10644);
nand U11183 (N_11183,N_9962,N_10193);
or U11184 (N_11184,N_10316,N_10118);
nor U11185 (N_11185,N_9965,N_10684);
or U11186 (N_11186,N_9832,N_10687);
xnor U11187 (N_11187,N_10121,N_9638);
and U11188 (N_11188,N_10157,N_10676);
or U11189 (N_11189,N_10131,N_10408);
nor U11190 (N_11190,N_9785,N_9859);
nand U11191 (N_11191,N_10752,N_10346);
xnor U11192 (N_11192,N_10733,N_10579);
xnor U11193 (N_11193,N_10067,N_10463);
nor U11194 (N_11194,N_10666,N_10163);
nand U11195 (N_11195,N_9927,N_10493);
nor U11196 (N_11196,N_10092,N_10329);
nand U11197 (N_11197,N_10005,N_10429);
or U11198 (N_11198,N_10394,N_10681);
or U11199 (N_11199,N_10682,N_10013);
nand U11200 (N_11200,N_10536,N_9922);
nor U11201 (N_11201,N_10249,N_10052);
nor U11202 (N_11202,N_9878,N_10326);
nor U11203 (N_11203,N_10782,N_10024);
nor U11204 (N_11204,N_10321,N_10588);
xor U11205 (N_11205,N_10075,N_9642);
nor U11206 (N_11206,N_10694,N_10668);
nor U11207 (N_11207,N_10304,N_9688);
or U11208 (N_11208,N_10445,N_9614);
xnor U11209 (N_11209,N_10460,N_9885);
and U11210 (N_11210,N_10616,N_9604);
and U11211 (N_11211,N_10128,N_9756);
xnor U11212 (N_11212,N_9685,N_9960);
or U11213 (N_11213,N_9932,N_10410);
xor U11214 (N_11214,N_9715,N_10220);
and U11215 (N_11215,N_10757,N_10743);
and U11216 (N_11216,N_10777,N_10341);
nand U11217 (N_11217,N_10455,N_10462);
nand U11218 (N_11218,N_10564,N_10477);
xor U11219 (N_11219,N_9750,N_9924);
xnor U11220 (N_11220,N_10414,N_10739);
xnor U11221 (N_11221,N_9670,N_9621);
xor U11222 (N_11222,N_10457,N_10747);
xnor U11223 (N_11223,N_9676,N_9725);
and U11224 (N_11224,N_10060,N_10152);
nand U11225 (N_11225,N_9694,N_9895);
nor U11226 (N_11226,N_10126,N_10740);
or U11227 (N_11227,N_9871,N_10055);
nor U11228 (N_11228,N_10019,N_9665);
or U11229 (N_11229,N_10440,N_9749);
and U11230 (N_11230,N_9853,N_9771);
or U11231 (N_11231,N_10768,N_9752);
or U11232 (N_11232,N_10604,N_10760);
nor U11233 (N_11233,N_10655,N_9647);
nor U11234 (N_11234,N_10492,N_9784);
and U11235 (N_11235,N_10358,N_10308);
and U11236 (N_11236,N_10554,N_10036);
nand U11237 (N_11237,N_10104,N_10192);
xor U11238 (N_11238,N_9796,N_10235);
and U11239 (N_11239,N_10009,N_10597);
and U11240 (N_11240,N_9869,N_10545);
and U11241 (N_11241,N_9726,N_10251);
nor U11242 (N_11242,N_10593,N_10263);
nor U11243 (N_11243,N_10726,N_10661);
nor U11244 (N_11244,N_10619,N_10277);
xnor U11245 (N_11245,N_10058,N_9677);
nand U11246 (N_11246,N_10790,N_10374);
or U11247 (N_11247,N_10456,N_10335);
xor U11248 (N_11248,N_9762,N_9864);
and U11249 (N_11249,N_9681,N_9910);
nand U11250 (N_11250,N_10110,N_10596);
nand U11251 (N_11251,N_10712,N_10755);
and U11252 (N_11252,N_9799,N_10488);
or U11253 (N_11253,N_9649,N_10206);
or U11254 (N_11254,N_10201,N_10375);
and U11255 (N_11255,N_10208,N_9810);
nor U11256 (N_11256,N_10444,N_10197);
or U11257 (N_11257,N_10490,N_10482);
or U11258 (N_11258,N_10369,N_10599);
or U11259 (N_11259,N_10178,N_10122);
nor U11260 (N_11260,N_10622,N_9926);
or U11261 (N_11261,N_9803,N_9733);
nor U11262 (N_11262,N_10256,N_10015);
xor U11263 (N_11263,N_10419,N_10706);
nand U11264 (N_11264,N_10245,N_10485);
nand U11265 (N_11265,N_10568,N_10447);
and U11266 (N_11266,N_10459,N_10046);
or U11267 (N_11267,N_10390,N_10051);
nand U11268 (N_11268,N_10047,N_10062);
nor U11269 (N_11269,N_9697,N_9788);
or U11270 (N_11270,N_10591,N_10771);
or U11271 (N_11271,N_9847,N_10795);
or U11272 (N_11272,N_10781,N_9656);
and U11273 (N_11273,N_9967,N_9751);
or U11274 (N_11274,N_10549,N_10586);
nor U11275 (N_11275,N_9989,N_10709);
nor U11276 (N_11276,N_9766,N_10552);
and U11277 (N_11277,N_10546,N_10427);
nand U11278 (N_11278,N_10540,N_9826);
nor U11279 (N_11279,N_10198,N_10432);
nor U11280 (N_11280,N_9635,N_10265);
or U11281 (N_11281,N_10791,N_10670);
nor U11282 (N_11282,N_9846,N_9856);
nand U11283 (N_11283,N_9680,N_9667);
and U11284 (N_11284,N_9831,N_9713);
nand U11285 (N_11285,N_9866,N_9724);
or U11286 (N_11286,N_10728,N_10620);
nand U11287 (N_11287,N_9805,N_10291);
nor U11288 (N_11288,N_10170,N_10083);
and U11289 (N_11289,N_10223,N_10789);
nand U11290 (N_11290,N_9998,N_10034);
nand U11291 (N_11291,N_10185,N_10629);
or U11292 (N_11292,N_10491,N_10044);
nor U11293 (N_11293,N_10515,N_10189);
xor U11294 (N_11294,N_10074,N_10678);
or U11295 (N_11295,N_9708,N_10519);
nor U11296 (N_11296,N_10632,N_9828);
nor U11297 (N_11297,N_10753,N_9710);
nand U11298 (N_11298,N_10200,N_10270);
nor U11299 (N_11299,N_10749,N_10544);
nor U11300 (N_11300,N_9949,N_10433);
nor U11301 (N_11301,N_9950,N_10636);
nor U11302 (N_11302,N_10173,N_10759);
and U11303 (N_11303,N_10210,N_10138);
nor U11304 (N_11304,N_9748,N_10228);
and U11305 (N_11305,N_10354,N_10186);
xor U11306 (N_11306,N_10303,N_10330);
nand U11307 (N_11307,N_10525,N_9975);
and U11308 (N_11308,N_9817,N_9981);
nor U11309 (N_11309,N_9741,N_10169);
and U11310 (N_11310,N_9862,N_9723);
or U11311 (N_11311,N_10030,N_10581);
and U11312 (N_11312,N_9672,N_10000);
and U11313 (N_11313,N_10233,N_9650);
or U11314 (N_11314,N_10336,N_10162);
nand U11315 (N_11315,N_9894,N_10696);
xor U11316 (N_11316,N_10496,N_9827);
and U11317 (N_11317,N_10143,N_10172);
or U11318 (N_11318,N_10407,N_9682);
xnor U11319 (N_11319,N_9934,N_10188);
nand U11320 (N_11320,N_10029,N_10290);
or U11321 (N_11321,N_10494,N_10657);
or U11322 (N_11322,N_10719,N_9978);
xor U11323 (N_11323,N_9684,N_9891);
or U11324 (N_11324,N_10267,N_9882);
nor U11325 (N_11325,N_10383,N_9722);
nand U11326 (N_11326,N_10059,N_9833);
nand U11327 (N_11327,N_10774,N_10731);
and U11328 (N_11328,N_9935,N_9849);
or U11329 (N_11329,N_10191,N_9838);
nor U11330 (N_11330,N_9835,N_10031);
nand U11331 (N_11331,N_10614,N_10275);
xnor U11332 (N_11332,N_10531,N_9629);
nand U11333 (N_11333,N_10582,N_10253);
xnor U11334 (N_11334,N_9646,N_10589);
nand U11335 (N_11335,N_10424,N_10648);
or U11336 (N_11336,N_9983,N_9652);
nand U11337 (N_11337,N_10324,N_10250);
and U11338 (N_11338,N_10262,N_10025);
nor U11339 (N_11339,N_9818,N_10167);
xor U11340 (N_11340,N_10215,N_10237);
nand U11341 (N_11341,N_10077,N_10605);
nor U11342 (N_11342,N_9901,N_10454);
or U11343 (N_11343,N_9623,N_10511);
nor U11344 (N_11344,N_9637,N_10293);
xor U11345 (N_11345,N_9806,N_9687);
xnor U11346 (N_11346,N_10780,N_10279);
nor U11347 (N_11347,N_9836,N_10020);
xnor U11348 (N_11348,N_9678,N_10656);
xnor U11349 (N_11349,N_10683,N_9930);
xnor U11350 (N_11350,N_10356,N_10086);
nand U11351 (N_11351,N_10295,N_10660);
xnor U11352 (N_11352,N_10282,N_10571);
nand U11353 (N_11353,N_10576,N_10087);
or U11354 (N_11354,N_9757,N_10633);
xor U11355 (N_11355,N_10766,N_10674);
nor U11356 (N_11356,N_10609,N_10350);
or U11357 (N_11357,N_9791,N_10391);
nand U11358 (N_11358,N_9966,N_9954);
xor U11359 (N_11359,N_10049,N_9633);
or U11360 (N_11360,N_10403,N_10328);
xnor U11361 (N_11361,N_10232,N_10323);
nand U11362 (N_11362,N_9969,N_9951);
nor U11363 (N_11363,N_10313,N_10359);
nand U11364 (N_11364,N_10507,N_9700);
nand U11365 (N_11365,N_10717,N_9789);
and U11366 (N_11366,N_9630,N_9600);
or U11367 (N_11367,N_10598,N_10078);
and U11368 (N_11368,N_10255,N_10475);
xor U11369 (N_11369,N_9760,N_10441);
nor U11370 (N_11370,N_10595,N_10453);
xor U11371 (N_11371,N_10194,N_9663);
or U11372 (N_11372,N_9892,N_10377);
or U11373 (N_11373,N_9976,N_10175);
and U11374 (N_11374,N_10035,N_9899);
and U11375 (N_11375,N_10750,N_9753);
nand U11376 (N_11376,N_10472,N_9972);
nand U11377 (N_11377,N_10088,N_10446);
nor U11378 (N_11378,N_10555,N_10252);
xnor U11379 (N_11379,N_9611,N_10180);
xor U11380 (N_11380,N_10017,N_10114);
and U11381 (N_11381,N_10084,N_9675);
and U11382 (N_11382,N_10124,N_9938);
xnor U11383 (N_11383,N_9886,N_9720);
xor U11384 (N_11384,N_10618,N_9958);
and U11385 (N_11385,N_10701,N_9758);
or U11386 (N_11386,N_10298,N_10796);
and U11387 (N_11387,N_10400,N_9917);
or U11388 (N_11388,N_10140,N_9738);
xor U11389 (N_11389,N_10505,N_10071);
and U11390 (N_11390,N_10468,N_10039);
or U11391 (N_11391,N_10018,N_10695);
nand U11392 (N_11392,N_9729,N_9963);
nor U11393 (N_11393,N_10653,N_10623);
and U11394 (N_11394,N_10625,N_10339);
or U11395 (N_11395,N_9995,N_10342);
nand U11396 (N_11396,N_10272,N_9695);
nand U11397 (N_11397,N_10151,N_10659);
xor U11398 (N_11398,N_10464,N_10714);
xnor U11399 (N_11399,N_10096,N_10306);
or U11400 (N_11400,N_10242,N_10722);
nand U11401 (N_11401,N_9907,N_10397);
or U11402 (N_11402,N_10684,N_10009);
or U11403 (N_11403,N_10269,N_10730);
and U11404 (N_11404,N_9757,N_10577);
nor U11405 (N_11405,N_9793,N_9841);
or U11406 (N_11406,N_10630,N_10050);
nand U11407 (N_11407,N_10787,N_10485);
nor U11408 (N_11408,N_10741,N_10292);
nand U11409 (N_11409,N_9928,N_10107);
nand U11410 (N_11410,N_9962,N_10436);
xnor U11411 (N_11411,N_10209,N_10689);
xor U11412 (N_11412,N_9705,N_10236);
xor U11413 (N_11413,N_10138,N_9724);
nand U11414 (N_11414,N_10084,N_10087);
or U11415 (N_11415,N_10009,N_9981);
or U11416 (N_11416,N_9648,N_9795);
nor U11417 (N_11417,N_9606,N_10523);
and U11418 (N_11418,N_10369,N_10108);
xor U11419 (N_11419,N_10007,N_10688);
nand U11420 (N_11420,N_10584,N_10528);
xor U11421 (N_11421,N_10733,N_10532);
or U11422 (N_11422,N_9707,N_10155);
and U11423 (N_11423,N_10113,N_9808);
or U11424 (N_11424,N_9610,N_10536);
or U11425 (N_11425,N_10108,N_9648);
nor U11426 (N_11426,N_10474,N_10309);
and U11427 (N_11427,N_9850,N_9967);
xnor U11428 (N_11428,N_10733,N_10174);
and U11429 (N_11429,N_10718,N_10501);
nor U11430 (N_11430,N_9624,N_9895);
xnor U11431 (N_11431,N_9912,N_10135);
and U11432 (N_11432,N_10552,N_10182);
xnor U11433 (N_11433,N_10176,N_10364);
or U11434 (N_11434,N_10523,N_10463);
nand U11435 (N_11435,N_10793,N_10365);
or U11436 (N_11436,N_10549,N_10739);
and U11437 (N_11437,N_9630,N_9669);
and U11438 (N_11438,N_10065,N_10753);
nor U11439 (N_11439,N_9765,N_10449);
xnor U11440 (N_11440,N_9602,N_9636);
and U11441 (N_11441,N_10367,N_9693);
xor U11442 (N_11442,N_10091,N_9771);
and U11443 (N_11443,N_9602,N_9938);
nor U11444 (N_11444,N_10795,N_10680);
nand U11445 (N_11445,N_10701,N_10333);
xnor U11446 (N_11446,N_9869,N_10171);
nand U11447 (N_11447,N_10296,N_10453);
nor U11448 (N_11448,N_9608,N_10782);
nor U11449 (N_11449,N_10042,N_10331);
xor U11450 (N_11450,N_10569,N_10355);
nand U11451 (N_11451,N_9946,N_9840);
xor U11452 (N_11452,N_9909,N_10411);
or U11453 (N_11453,N_10049,N_9982);
or U11454 (N_11454,N_9806,N_9779);
or U11455 (N_11455,N_10457,N_9617);
and U11456 (N_11456,N_10093,N_10391);
nor U11457 (N_11457,N_9817,N_10627);
xnor U11458 (N_11458,N_10622,N_9778);
or U11459 (N_11459,N_9633,N_9729);
nor U11460 (N_11460,N_10110,N_10330);
nand U11461 (N_11461,N_10647,N_10643);
and U11462 (N_11462,N_9966,N_9987);
or U11463 (N_11463,N_10513,N_10572);
nor U11464 (N_11464,N_9616,N_10322);
xor U11465 (N_11465,N_10413,N_9742);
and U11466 (N_11466,N_10305,N_10126);
xor U11467 (N_11467,N_10300,N_9669);
or U11468 (N_11468,N_9833,N_10418);
and U11469 (N_11469,N_10077,N_9798);
and U11470 (N_11470,N_10086,N_10475);
or U11471 (N_11471,N_10292,N_10479);
xnor U11472 (N_11472,N_10483,N_10435);
and U11473 (N_11473,N_9770,N_9626);
and U11474 (N_11474,N_10256,N_10355);
nand U11475 (N_11475,N_9857,N_10453);
or U11476 (N_11476,N_9866,N_10519);
nand U11477 (N_11477,N_10326,N_9626);
xnor U11478 (N_11478,N_10328,N_10427);
xor U11479 (N_11479,N_10353,N_10705);
nand U11480 (N_11480,N_9997,N_10044);
or U11481 (N_11481,N_10435,N_9993);
and U11482 (N_11482,N_9738,N_9783);
xor U11483 (N_11483,N_10207,N_10357);
and U11484 (N_11484,N_10555,N_9640);
and U11485 (N_11485,N_10301,N_10797);
or U11486 (N_11486,N_10188,N_10688);
xnor U11487 (N_11487,N_10640,N_9943);
nand U11488 (N_11488,N_10714,N_10108);
and U11489 (N_11489,N_10117,N_10165);
and U11490 (N_11490,N_10713,N_10124);
and U11491 (N_11491,N_10189,N_10479);
xnor U11492 (N_11492,N_10139,N_9633);
xor U11493 (N_11493,N_10002,N_10475);
nor U11494 (N_11494,N_9912,N_10589);
and U11495 (N_11495,N_10128,N_10234);
xnor U11496 (N_11496,N_10747,N_9756);
nor U11497 (N_11497,N_10657,N_9714);
or U11498 (N_11498,N_9681,N_10538);
xnor U11499 (N_11499,N_10785,N_9704);
nand U11500 (N_11500,N_9855,N_10705);
nand U11501 (N_11501,N_10554,N_9908);
nand U11502 (N_11502,N_9707,N_10404);
xnor U11503 (N_11503,N_10463,N_10702);
nand U11504 (N_11504,N_10377,N_10174);
and U11505 (N_11505,N_10652,N_10634);
or U11506 (N_11506,N_10383,N_10426);
or U11507 (N_11507,N_10087,N_10518);
xnor U11508 (N_11508,N_10612,N_9993);
nand U11509 (N_11509,N_10178,N_9794);
xnor U11510 (N_11510,N_10724,N_9790);
xnor U11511 (N_11511,N_10064,N_10617);
or U11512 (N_11512,N_10684,N_9864);
xnor U11513 (N_11513,N_9681,N_10749);
nor U11514 (N_11514,N_10634,N_9751);
or U11515 (N_11515,N_10401,N_10142);
nand U11516 (N_11516,N_9732,N_10495);
xnor U11517 (N_11517,N_9652,N_10431);
nand U11518 (N_11518,N_9979,N_10766);
xor U11519 (N_11519,N_10518,N_9703);
or U11520 (N_11520,N_10097,N_9991);
xnor U11521 (N_11521,N_9854,N_9910);
nor U11522 (N_11522,N_10245,N_10357);
xor U11523 (N_11523,N_9644,N_10365);
xnor U11524 (N_11524,N_10313,N_9699);
nand U11525 (N_11525,N_10769,N_9956);
xor U11526 (N_11526,N_10382,N_10599);
and U11527 (N_11527,N_9639,N_10706);
or U11528 (N_11528,N_9763,N_10203);
or U11529 (N_11529,N_10088,N_10076);
nor U11530 (N_11530,N_10513,N_9789);
nand U11531 (N_11531,N_9645,N_9633);
or U11532 (N_11532,N_10576,N_10124);
and U11533 (N_11533,N_10467,N_9641);
nor U11534 (N_11534,N_9929,N_9612);
xor U11535 (N_11535,N_10087,N_10566);
or U11536 (N_11536,N_9725,N_10709);
and U11537 (N_11537,N_9607,N_9933);
or U11538 (N_11538,N_9812,N_10018);
nor U11539 (N_11539,N_10613,N_10338);
nor U11540 (N_11540,N_9868,N_10353);
nor U11541 (N_11541,N_10260,N_9628);
nor U11542 (N_11542,N_9804,N_10251);
nor U11543 (N_11543,N_10572,N_10735);
and U11544 (N_11544,N_9794,N_10050);
nor U11545 (N_11545,N_10372,N_10695);
nor U11546 (N_11546,N_9692,N_10297);
or U11547 (N_11547,N_10713,N_9944);
and U11548 (N_11548,N_10597,N_10645);
xnor U11549 (N_11549,N_9746,N_9748);
or U11550 (N_11550,N_10561,N_10616);
xor U11551 (N_11551,N_10248,N_10433);
and U11552 (N_11552,N_10167,N_10118);
or U11553 (N_11553,N_10006,N_9899);
nor U11554 (N_11554,N_9782,N_9829);
and U11555 (N_11555,N_10658,N_9940);
xnor U11556 (N_11556,N_9801,N_10150);
xor U11557 (N_11557,N_10510,N_10013);
xnor U11558 (N_11558,N_10261,N_10193);
nor U11559 (N_11559,N_10655,N_10590);
nand U11560 (N_11560,N_9603,N_9894);
or U11561 (N_11561,N_9620,N_9739);
nand U11562 (N_11562,N_10202,N_10325);
nor U11563 (N_11563,N_10418,N_10513);
xnor U11564 (N_11564,N_10150,N_10021);
and U11565 (N_11565,N_10386,N_10144);
nand U11566 (N_11566,N_10718,N_9754);
or U11567 (N_11567,N_9848,N_10509);
nor U11568 (N_11568,N_10477,N_10582);
or U11569 (N_11569,N_10696,N_10704);
nor U11570 (N_11570,N_10648,N_9698);
or U11571 (N_11571,N_9919,N_9852);
xnor U11572 (N_11572,N_10272,N_10189);
nand U11573 (N_11573,N_9844,N_10386);
xor U11574 (N_11574,N_10771,N_10633);
nand U11575 (N_11575,N_10372,N_10177);
or U11576 (N_11576,N_10551,N_10436);
nor U11577 (N_11577,N_10679,N_10413);
and U11578 (N_11578,N_9748,N_10193);
and U11579 (N_11579,N_10087,N_9933);
xor U11580 (N_11580,N_10653,N_10047);
nand U11581 (N_11581,N_9702,N_9688);
and U11582 (N_11582,N_10134,N_10441);
xor U11583 (N_11583,N_10389,N_9801);
nor U11584 (N_11584,N_9618,N_9832);
nand U11585 (N_11585,N_9961,N_10191);
nor U11586 (N_11586,N_9840,N_10343);
nand U11587 (N_11587,N_10769,N_9885);
or U11588 (N_11588,N_10067,N_10757);
nor U11589 (N_11589,N_10756,N_10322);
xor U11590 (N_11590,N_10747,N_10417);
and U11591 (N_11591,N_10612,N_10755);
and U11592 (N_11592,N_10089,N_10100);
and U11593 (N_11593,N_10071,N_10465);
and U11594 (N_11594,N_10586,N_10645);
nand U11595 (N_11595,N_9637,N_10723);
nand U11596 (N_11596,N_10744,N_10226);
nor U11597 (N_11597,N_9838,N_10374);
xor U11598 (N_11598,N_9731,N_10775);
and U11599 (N_11599,N_9642,N_10012);
or U11600 (N_11600,N_9966,N_10050);
nand U11601 (N_11601,N_10373,N_10789);
or U11602 (N_11602,N_9887,N_10747);
xor U11603 (N_11603,N_10693,N_9739);
xnor U11604 (N_11604,N_10271,N_10676);
xor U11605 (N_11605,N_9628,N_10689);
nor U11606 (N_11606,N_10037,N_9690);
nand U11607 (N_11607,N_9878,N_9872);
or U11608 (N_11608,N_9900,N_10197);
and U11609 (N_11609,N_10212,N_10624);
nor U11610 (N_11610,N_10152,N_10432);
xnor U11611 (N_11611,N_10206,N_10194);
or U11612 (N_11612,N_10016,N_10405);
nand U11613 (N_11613,N_9773,N_10168);
xnor U11614 (N_11614,N_10028,N_10293);
nand U11615 (N_11615,N_10088,N_10113);
nor U11616 (N_11616,N_10145,N_10535);
nand U11617 (N_11617,N_10112,N_9758);
and U11618 (N_11618,N_10690,N_10165);
nand U11619 (N_11619,N_9620,N_10306);
xnor U11620 (N_11620,N_10480,N_9782);
or U11621 (N_11621,N_10151,N_10188);
and U11622 (N_11622,N_9759,N_9629);
nor U11623 (N_11623,N_10061,N_10175);
xnor U11624 (N_11624,N_10421,N_10184);
nor U11625 (N_11625,N_10531,N_10274);
and U11626 (N_11626,N_10014,N_9822);
and U11627 (N_11627,N_10300,N_10450);
nand U11628 (N_11628,N_10718,N_9610);
and U11629 (N_11629,N_10653,N_10585);
nand U11630 (N_11630,N_9867,N_10597);
or U11631 (N_11631,N_10117,N_9690);
and U11632 (N_11632,N_10289,N_9866);
xnor U11633 (N_11633,N_10779,N_10663);
and U11634 (N_11634,N_9649,N_9705);
nor U11635 (N_11635,N_10080,N_10181);
nand U11636 (N_11636,N_10105,N_10352);
nor U11637 (N_11637,N_10736,N_10628);
or U11638 (N_11638,N_10255,N_10390);
nand U11639 (N_11639,N_10165,N_10126);
or U11640 (N_11640,N_10790,N_10741);
nor U11641 (N_11641,N_9724,N_10668);
nor U11642 (N_11642,N_10321,N_9695);
and U11643 (N_11643,N_10463,N_10157);
nor U11644 (N_11644,N_9910,N_10532);
xor U11645 (N_11645,N_9662,N_9983);
nor U11646 (N_11646,N_10136,N_9776);
nand U11647 (N_11647,N_10351,N_9822);
or U11648 (N_11648,N_9773,N_10784);
and U11649 (N_11649,N_10568,N_10672);
and U11650 (N_11650,N_10558,N_9914);
and U11651 (N_11651,N_10321,N_10296);
nand U11652 (N_11652,N_10283,N_9657);
xor U11653 (N_11653,N_10118,N_10591);
or U11654 (N_11654,N_9826,N_9882);
nor U11655 (N_11655,N_9755,N_10501);
and U11656 (N_11656,N_10054,N_10102);
nor U11657 (N_11657,N_9919,N_9695);
nand U11658 (N_11658,N_9895,N_9848);
and U11659 (N_11659,N_10375,N_9811);
nand U11660 (N_11660,N_10735,N_9646);
and U11661 (N_11661,N_10198,N_9972);
xnor U11662 (N_11662,N_10545,N_9931);
or U11663 (N_11663,N_10466,N_10195);
or U11664 (N_11664,N_10542,N_10238);
nor U11665 (N_11665,N_10538,N_10549);
or U11666 (N_11666,N_10377,N_10417);
xor U11667 (N_11667,N_9966,N_10507);
or U11668 (N_11668,N_10779,N_10351);
xnor U11669 (N_11669,N_10232,N_9871);
nor U11670 (N_11670,N_10595,N_9879);
and U11671 (N_11671,N_10598,N_10084);
and U11672 (N_11672,N_10084,N_10687);
xnor U11673 (N_11673,N_9904,N_10354);
and U11674 (N_11674,N_10427,N_9937);
or U11675 (N_11675,N_10252,N_9669);
nand U11676 (N_11676,N_9653,N_9739);
and U11677 (N_11677,N_10083,N_10155);
nor U11678 (N_11678,N_9978,N_9744);
and U11679 (N_11679,N_10356,N_10427);
nor U11680 (N_11680,N_10198,N_10550);
nand U11681 (N_11681,N_10722,N_9987);
xor U11682 (N_11682,N_10077,N_10602);
and U11683 (N_11683,N_10257,N_10070);
xor U11684 (N_11684,N_10704,N_10509);
nor U11685 (N_11685,N_10157,N_9846);
nor U11686 (N_11686,N_10526,N_9871);
or U11687 (N_11687,N_10046,N_9863);
nor U11688 (N_11688,N_9905,N_9867);
xnor U11689 (N_11689,N_10102,N_10076);
nor U11690 (N_11690,N_10342,N_10773);
xnor U11691 (N_11691,N_10436,N_10571);
or U11692 (N_11692,N_10725,N_10782);
xor U11693 (N_11693,N_10563,N_9996);
and U11694 (N_11694,N_9671,N_9779);
nor U11695 (N_11695,N_10728,N_10457);
and U11696 (N_11696,N_10798,N_10263);
or U11697 (N_11697,N_9766,N_9707);
nor U11698 (N_11698,N_10388,N_10536);
and U11699 (N_11699,N_9924,N_10304);
and U11700 (N_11700,N_10493,N_9660);
xor U11701 (N_11701,N_10751,N_9979);
and U11702 (N_11702,N_10339,N_10301);
and U11703 (N_11703,N_10579,N_10681);
nor U11704 (N_11704,N_10539,N_10018);
nand U11705 (N_11705,N_10320,N_10151);
xnor U11706 (N_11706,N_10348,N_10791);
or U11707 (N_11707,N_9726,N_9952);
xnor U11708 (N_11708,N_9750,N_10204);
nor U11709 (N_11709,N_10101,N_9723);
nand U11710 (N_11710,N_9814,N_9614);
xnor U11711 (N_11711,N_10757,N_10731);
and U11712 (N_11712,N_10602,N_10295);
or U11713 (N_11713,N_10377,N_10783);
and U11714 (N_11714,N_10699,N_10336);
xor U11715 (N_11715,N_10420,N_9872);
xnor U11716 (N_11716,N_10008,N_10414);
nand U11717 (N_11717,N_10699,N_10657);
and U11718 (N_11718,N_9951,N_10356);
nand U11719 (N_11719,N_10626,N_9835);
nand U11720 (N_11720,N_10434,N_10610);
nor U11721 (N_11721,N_10005,N_10309);
nand U11722 (N_11722,N_9799,N_10057);
and U11723 (N_11723,N_10182,N_9676);
nand U11724 (N_11724,N_9837,N_9651);
and U11725 (N_11725,N_10125,N_10770);
or U11726 (N_11726,N_10018,N_9620);
xnor U11727 (N_11727,N_10040,N_9799);
xnor U11728 (N_11728,N_10677,N_10495);
and U11729 (N_11729,N_10112,N_10781);
xor U11730 (N_11730,N_10717,N_10666);
or U11731 (N_11731,N_10456,N_10671);
nor U11732 (N_11732,N_9670,N_10684);
xor U11733 (N_11733,N_10089,N_10134);
or U11734 (N_11734,N_10484,N_9963);
nand U11735 (N_11735,N_9867,N_9728);
xnor U11736 (N_11736,N_9717,N_9926);
xnor U11737 (N_11737,N_10455,N_9983);
nor U11738 (N_11738,N_10008,N_10663);
or U11739 (N_11739,N_10392,N_10775);
or U11740 (N_11740,N_10784,N_9931);
nor U11741 (N_11741,N_10516,N_9992);
xor U11742 (N_11742,N_10465,N_10049);
or U11743 (N_11743,N_10478,N_10065);
nor U11744 (N_11744,N_10212,N_10208);
xor U11745 (N_11745,N_10634,N_10108);
nor U11746 (N_11746,N_9761,N_10511);
nand U11747 (N_11747,N_10701,N_9609);
xnor U11748 (N_11748,N_9975,N_10274);
and U11749 (N_11749,N_9602,N_10260);
and U11750 (N_11750,N_10363,N_10360);
or U11751 (N_11751,N_9602,N_9706);
nand U11752 (N_11752,N_10637,N_10517);
xor U11753 (N_11753,N_9942,N_10263);
nor U11754 (N_11754,N_10369,N_9849);
nand U11755 (N_11755,N_10066,N_10142);
and U11756 (N_11756,N_10438,N_10090);
and U11757 (N_11757,N_10464,N_9815);
or U11758 (N_11758,N_10407,N_10333);
nand U11759 (N_11759,N_10026,N_10643);
and U11760 (N_11760,N_10620,N_9748);
and U11761 (N_11761,N_9871,N_10073);
xnor U11762 (N_11762,N_10302,N_10053);
or U11763 (N_11763,N_10425,N_9789);
nand U11764 (N_11764,N_10386,N_9606);
nor U11765 (N_11765,N_9781,N_10509);
or U11766 (N_11766,N_10508,N_10517);
nand U11767 (N_11767,N_9921,N_10203);
nor U11768 (N_11768,N_10620,N_10271);
xnor U11769 (N_11769,N_9650,N_10216);
or U11770 (N_11770,N_10397,N_10123);
nand U11771 (N_11771,N_10633,N_9605);
xnor U11772 (N_11772,N_9769,N_10582);
nand U11773 (N_11773,N_10027,N_10777);
xor U11774 (N_11774,N_10124,N_9976);
nand U11775 (N_11775,N_9839,N_10652);
nor U11776 (N_11776,N_10383,N_10442);
xnor U11777 (N_11777,N_10684,N_10775);
xor U11778 (N_11778,N_10172,N_10480);
and U11779 (N_11779,N_10426,N_10776);
nor U11780 (N_11780,N_10053,N_10079);
nand U11781 (N_11781,N_10421,N_10396);
nor U11782 (N_11782,N_9677,N_9719);
nand U11783 (N_11783,N_10386,N_9989);
xnor U11784 (N_11784,N_9957,N_10256);
nor U11785 (N_11785,N_10276,N_10388);
and U11786 (N_11786,N_10321,N_10005);
xnor U11787 (N_11787,N_10023,N_10436);
nand U11788 (N_11788,N_10587,N_10684);
xor U11789 (N_11789,N_10043,N_9877);
nand U11790 (N_11790,N_9769,N_10326);
nor U11791 (N_11791,N_10470,N_9968);
and U11792 (N_11792,N_10300,N_10202);
xnor U11793 (N_11793,N_10569,N_10457);
nand U11794 (N_11794,N_9923,N_10494);
nand U11795 (N_11795,N_10076,N_10455);
and U11796 (N_11796,N_9846,N_10513);
or U11797 (N_11797,N_9647,N_10787);
nor U11798 (N_11798,N_10103,N_10205);
or U11799 (N_11799,N_10677,N_10115);
nand U11800 (N_11800,N_9623,N_10429);
or U11801 (N_11801,N_10413,N_10124);
nand U11802 (N_11802,N_10154,N_10189);
nand U11803 (N_11803,N_10549,N_9676);
and U11804 (N_11804,N_10465,N_10102);
xor U11805 (N_11805,N_10626,N_10554);
and U11806 (N_11806,N_10051,N_10395);
and U11807 (N_11807,N_10017,N_9698);
and U11808 (N_11808,N_10248,N_10375);
and U11809 (N_11809,N_10686,N_9843);
xnor U11810 (N_11810,N_10784,N_10737);
nor U11811 (N_11811,N_9988,N_9660);
xor U11812 (N_11812,N_9602,N_10553);
and U11813 (N_11813,N_10152,N_9915);
and U11814 (N_11814,N_9689,N_10676);
and U11815 (N_11815,N_9878,N_10402);
nand U11816 (N_11816,N_10681,N_10364);
xor U11817 (N_11817,N_9704,N_10657);
nor U11818 (N_11818,N_10015,N_10348);
nand U11819 (N_11819,N_9787,N_10722);
nand U11820 (N_11820,N_9822,N_10796);
and U11821 (N_11821,N_10585,N_10214);
xor U11822 (N_11822,N_9699,N_9625);
nand U11823 (N_11823,N_9845,N_9943);
nand U11824 (N_11824,N_10785,N_10617);
xor U11825 (N_11825,N_9813,N_10756);
xor U11826 (N_11826,N_9997,N_9649);
nand U11827 (N_11827,N_10386,N_10678);
xnor U11828 (N_11828,N_10200,N_9725);
nor U11829 (N_11829,N_10569,N_10052);
and U11830 (N_11830,N_9687,N_10466);
nor U11831 (N_11831,N_10142,N_10666);
nand U11832 (N_11832,N_10380,N_10319);
xor U11833 (N_11833,N_9912,N_10131);
nand U11834 (N_11834,N_9885,N_9854);
xnor U11835 (N_11835,N_10333,N_9746);
nand U11836 (N_11836,N_10215,N_10689);
nand U11837 (N_11837,N_10202,N_9739);
xor U11838 (N_11838,N_9892,N_10204);
or U11839 (N_11839,N_10346,N_10047);
xor U11840 (N_11840,N_10518,N_9794);
xor U11841 (N_11841,N_10616,N_10492);
nor U11842 (N_11842,N_9978,N_10257);
xor U11843 (N_11843,N_10662,N_9662);
xnor U11844 (N_11844,N_10468,N_9698);
nand U11845 (N_11845,N_10188,N_9956);
and U11846 (N_11846,N_10462,N_9762);
xnor U11847 (N_11847,N_9784,N_9608);
nor U11848 (N_11848,N_10779,N_9964);
nor U11849 (N_11849,N_10731,N_9646);
or U11850 (N_11850,N_10222,N_9928);
or U11851 (N_11851,N_9888,N_10663);
xor U11852 (N_11852,N_9993,N_9939);
or U11853 (N_11853,N_10030,N_10212);
or U11854 (N_11854,N_10165,N_10101);
or U11855 (N_11855,N_10515,N_10473);
or U11856 (N_11856,N_10797,N_10653);
and U11857 (N_11857,N_9745,N_10786);
or U11858 (N_11858,N_10246,N_10212);
nor U11859 (N_11859,N_9927,N_10067);
and U11860 (N_11860,N_10399,N_10385);
nor U11861 (N_11861,N_10398,N_10666);
xnor U11862 (N_11862,N_9978,N_9957);
or U11863 (N_11863,N_9791,N_9991);
nand U11864 (N_11864,N_9988,N_9664);
or U11865 (N_11865,N_9941,N_10036);
xor U11866 (N_11866,N_10384,N_10641);
nor U11867 (N_11867,N_9769,N_10741);
nor U11868 (N_11868,N_9835,N_10586);
nor U11869 (N_11869,N_10785,N_9713);
or U11870 (N_11870,N_10473,N_9812);
or U11871 (N_11871,N_10668,N_10341);
or U11872 (N_11872,N_10259,N_10556);
and U11873 (N_11873,N_9686,N_9644);
nor U11874 (N_11874,N_10395,N_10217);
nor U11875 (N_11875,N_10185,N_10679);
xnor U11876 (N_11876,N_10740,N_10251);
and U11877 (N_11877,N_9912,N_10174);
or U11878 (N_11878,N_9605,N_10069);
nor U11879 (N_11879,N_10671,N_10275);
nand U11880 (N_11880,N_10672,N_10691);
nor U11881 (N_11881,N_10323,N_10491);
and U11882 (N_11882,N_9918,N_10371);
nand U11883 (N_11883,N_10103,N_10001);
and U11884 (N_11884,N_10362,N_10517);
xor U11885 (N_11885,N_10003,N_10642);
nand U11886 (N_11886,N_10211,N_10761);
nor U11887 (N_11887,N_10146,N_10033);
nand U11888 (N_11888,N_9844,N_10197);
xor U11889 (N_11889,N_10234,N_10112);
xor U11890 (N_11890,N_10038,N_10168);
and U11891 (N_11891,N_10036,N_10462);
nand U11892 (N_11892,N_9616,N_10188);
nand U11893 (N_11893,N_9993,N_10255);
xor U11894 (N_11894,N_10728,N_9801);
or U11895 (N_11895,N_10436,N_9878);
nor U11896 (N_11896,N_10571,N_9898);
and U11897 (N_11897,N_10007,N_10446);
nor U11898 (N_11898,N_10435,N_10404);
nand U11899 (N_11899,N_9706,N_10798);
xor U11900 (N_11900,N_9858,N_9932);
nand U11901 (N_11901,N_10164,N_9699);
nor U11902 (N_11902,N_10238,N_10391);
xor U11903 (N_11903,N_9734,N_10098);
xor U11904 (N_11904,N_10276,N_10037);
or U11905 (N_11905,N_10234,N_9767);
nor U11906 (N_11906,N_10531,N_10637);
xor U11907 (N_11907,N_9923,N_9857);
xnor U11908 (N_11908,N_9711,N_10290);
nand U11909 (N_11909,N_10553,N_10250);
and U11910 (N_11910,N_10433,N_10782);
xor U11911 (N_11911,N_9771,N_10003);
xor U11912 (N_11912,N_10387,N_9869);
xnor U11913 (N_11913,N_9801,N_10715);
xor U11914 (N_11914,N_10366,N_10197);
xnor U11915 (N_11915,N_10485,N_10194);
or U11916 (N_11916,N_9703,N_10180);
nor U11917 (N_11917,N_9821,N_10504);
nor U11918 (N_11918,N_10623,N_10461);
or U11919 (N_11919,N_9966,N_10112);
xor U11920 (N_11920,N_10492,N_9670);
and U11921 (N_11921,N_10145,N_9679);
and U11922 (N_11922,N_9736,N_10449);
nand U11923 (N_11923,N_10075,N_10067);
and U11924 (N_11924,N_9964,N_10745);
nor U11925 (N_11925,N_9602,N_9940);
nor U11926 (N_11926,N_9672,N_10251);
xnor U11927 (N_11927,N_10587,N_10779);
nor U11928 (N_11928,N_9859,N_10191);
xor U11929 (N_11929,N_9934,N_9748);
nand U11930 (N_11930,N_10040,N_9631);
nand U11931 (N_11931,N_9917,N_10203);
and U11932 (N_11932,N_10335,N_10085);
or U11933 (N_11933,N_10691,N_10688);
and U11934 (N_11934,N_10412,N_10166);
xor U11935 (N_11935,N_10244,N_10538);
or U11936 (N_11936,N_10615,N_9920);
and U11937 (N_11937,N_9678,N_9868);
or U11938 (N_11938,N_9977,N_10771);
or U11939 (N_11939,N_10325,N_10001);
and U11940 (N_11940,N_10782,N_10783);
or U11941 (N_11941,N_10103,N_10724);
or U11942 (N_11942,N_10719,N_9982);
and U11943 (N_11943,N_9600,N_10433);
and U11944 (N_11944,N_9666,N_10611);
xor U11945 (N_11945,N_10126,N_10070);
nor U11946 (N_11946,N_10442,N_9740);
and U11947 (N_11947,N_9615,N_10400);
or U11948 (N_11948,N_9767,N_9789);
nor U11949 (N_11949,N_9957,N_9876);
or U11950 (N_11950,N_9967,N_10439);
xnor U11951 (N_11951,N_9861,N_10025);
xor U11952 (N_11952,N_10663,N_10394);
nand U11953 (N_11953,N_10639,N_10059);
or U11954 (N_11954,N_10531,N_10712);
or U11955 (N_11955,N_9977,N_9755);
and U11956 (N_11956,N_10134,N_10021);
xnor U11957 (N_11957,N_9927,N_9796);
or U11958 (N_11958,N_10193,N_10581);
nand U11959 (N_11959,N_10483,N_10086);
xor U11960 (N_11960,N_10115,N_10426);
and U11961 (N_11961,N_10257,N_9812);
xnor U11962 (N_11962,N_9901,N_10065);
nor U11963 (N_11963,N_9704,N_10452);
xor U11964 (N_11964,N_10472,N_9667);
or U11965 (N_11965,N_10776,N_10220);
and U11966 (N_11966,N_9992,N_10166);
and U11967 (N_11967,N_10548,N_10633);
nand U11968 (N_11968,N_10576,N_10165);
nor U11969 (N_11969,N_10548,N_10257);
nand U11970 (N_11970,N_10361,N_9819);
nor U11971 (N_11971,N_10746,N_10074);
and U11972 (N_11972,N_9771,N_9856);
nor U11973 (N_11973,N_10561,N_10597);
and U11974 (N_11974,N_9692,N_9897);
xor U11975 (N_11975,N_9601,N_10598);
or U11976 (N_11976,N_10760,N_9871);
xor U11977 (N_11977,N_10032,N_10295);
and U11978 (N_11978,N_9888,N_10729);
xnor U11979 (N_11979,N_9822,N_10734);
xor U11980 (N_11980,N_9894,N_10693);
or U11981 (N_11981,N_10136,N_10362);
nor U11982 (N_11982,N_10082,N_9983);
nand U11983 (N_11983,N_9945,N_10438);
nor U11984 (N_11984,N_10759,N_10339);
xor U11985 (N_11985,N_9949,N_10256);
nand U11986 (N_11986,N_9749,N_10586);
nor U11987 (N_11987,N_10378,N_10321);
xnor U11988 (N_11988,N_10696,N_9719);
nor U11989 (N_11989,N_10287,N_9672);
or U11990 (N_11990,N_9919,N_10066);
nor U11991 (N_11991,N_10727,N_10168);
nand U11992 (N_11992,N_10237,N_10253);
and U11993 (N_11993,N_10074,N_10426);
and U11994 (N_11994,N_10613,N_9971);
nand U11995 (N_11995,N_10483,N_10068);
and U11996 (N_11996,N_10748,N_10762);
or U11997 (N_11997,N_10143,N_10106);
nor U11998 (N_11998,N_9888,N_10527);
and U11999 (N_11999,N_10401,N_10757);
nor U12000 (N_12000,N_11527,N_11987);
nor U12001 (N_12001,N_11631,N_11869);
nor U12002 (N_12002,N_11881,N_11727);
or U12003 (N_12003,N_11338,N_10965);
nor U12004 (N_12004,N_11788,N_10907);
or U12005 (N_12005,N_11503,N_11502);
and U12006 (N_12006,N_11893,N_11783);
nand U12007 (N_12007,N_11237,N_11029);
or U12008 (N_12008,N_10958,N_10826);
and U12009 (N_12009,N_11397,N_11958);
xnor U12010 (N_12010,N_11887,N_11567);
nor U12011 (N_12011,N_11110,N_11256);
or U12012 (N_12012,N_11196,N_11455);
nor U12013 (N_12013,N_11461,N_11773);
xnor U12014 (N_12014,N_11889,N_11373);
nor U12015 (N_12015,N_11506,N_11806);
nand U12016 (N_12016,N_11711,N_10909);
xnor U12017 (N_12017,N_10819,N_11764);
and U12018 (N_12018,N_11908,N_11482);
and U12019 (N_12019,N_11756,N_11736);
or U12020 (N_12020,N_11609,N_10840);
nand U12021 (N_12021,N_11653,N_11369);
or U12022 (N_12022,N_11524,N_11480);
xnor U12023 (N_12023,N_11345,N_11552);
nor U12024 (N_12024,N_10821,N_11048);
nor U12025 (N_12025,N_11374,N_11819);
and U12026 (N_12026,N_11250,N_11953);
or U12027 (N_12027,N_10946,N_11423);
xnor U12028 (N_12028,N_11106,N_10857);
and U12029 (N_12029,N_11745,N_11422);
nor U12030 (N_12030,N_10845,N_11620);
nand U12031 (N_12031,N_11675,N_11429);
and U12032 (N_12032,N_11521,N_11238);
xor U12033 (N_12033,N_11608,N_11544);
nand U12034 (N_12034,N_11467,N_11769);
or U12035 (N_12035,N_10871,N_11353);
xor U12036 (N_12036,N_10829,N_11744);
nor U12037 (N_12037,N_10966,N_11504);
xnor U12038 (N_12038,N_10942,N_11817);
xor U12039 (N_12039,N_11629,N_10868);
nand U12040 (N_12040,N_11842,N_11257);
and U12041 (N_12041,N_11963,N_11207);
or U12042 (N_12042,N_11417,N_11137);
and U12043 (N_12043,N_11335,N_10924);
or U12044 (N_12044,N_11976,N_11796);
nand U12045 (N_12045,N_11245,N_11244);
nor U12046 (N_12046,N_11367,N_11154);
nor U12047 (N_12047,N_11886,N_11160);
nand U12048 (N_12048,N_10832,N_11410);
nor U12049 (N_12049,N_10849,N_11197);
and U12050 (N_12050,N_11464,N_11743);
and U12051 (N_12051,N_11329,N_11688);
or U12052 (N_12052,N_10866,N_11265);
nand U12053 (N_12053,N_11651,N_11258);
xnor U12054 (N_12054,N_11680,N_11710);
nand U12055 (N_12055,N_10985,N_11451);
or U12056 (N_12056,N_11514,N_11066);
xnor U12057 (N_12057,N_11926,N_11771);
or U12058 (N_12058,N_11898,N_11900);
nand U12059 (N_12059,N_11937,N_11253);
or U12060 (N_12060,N_10861,N_11087);
nor U12061 (N_12061,N_11610,N_11492);
xor U12062 (N_12062,N_11316,N_11565);
nor U12063 (N_12063,N_11936,N_11600);
nand U12064 (N_12064,N_11861,N_10839);
or U12065 (N_12065,N_11479,N_11089);
nand U12066 (N_12066,N_11208,N_11008);
or U12067 (N_12067,N_11985,N_11759);
and U12068 (N_12068,N_11334,N_10919);
nor U12069 (N_12069,N_11853,N_10895);
and U12070 (N_12070,N_11722,N_11115);
and U12071 (N_12071,N_11645,N_10921);
nand U12072 (N_12072,N_10859,N_11992);
and U12073 (N_12073,N_11101,N_11165);
xnor U12074 (N_12074,N_11532,N_11302);
nor U12075 (N_12075,N_11324,N_10976);
nand U12076 (N_12076,N_11077,N_10908);
xnor U12077 (N_12077,N_11203,N_10830);
nand U12078 (N_12078,N_11844,N_11589);
nand U12079 (N_12079,N_11116,N_11109);
nand U12080 (N_12080,N_11179,N_11959);
nor U12081 (N_12081,N_10884,N_11857);
nand U12082 (N_12082,N_10864,N_11108);
nand U12083 (N_12083,N_11990,N_11453);
nor U12084 (N_12084,N_10936,N_11734);
nand U12085 (N_12085,N_11498,N_10929);
nor U12086 (N_12086,N_11950,N_11342);
xor U12087 (N_12087,N_11080,N_11475);
nor U12088 (N_12088,N_11272,N_11728);
xor U12089 (N_12089,N_10996,N_11884);
xnor U12090 (N_12090,N_11988,N_11548);
xnor U12091 (N_12091,N_11776,N_11571);
nor U12092 (N_12092,N_11222,N_11432);
and U12093 (N_12093,N_11828,N_11568);
or U12094 (N_12094,N_11639,N_10964);
and U12095 (N_12095,N_11454,N_11184);
xnor U12096 (N_12096,N_11533,N_11906);
xor U12097 (N_12097,N_11189,N_11173);
nand U12098 (N_12098,N_10860,N_11669);
or U12099 (N_12099,N_10945,N_11279);
nor U12100 (N_12100,N_11810,N_10977);
nor U12101 (N_12101,N_11216,N_10865);
and U12102 (N_12102,N_11843,N_11136);
xnor U12103 (N_12103,N_11779,N_11124);
xor U12104 (N_12104,N_11932,N_11473);
and U12105 (N_12105,N_11726,N_11161);
or U12106 (N_12106,N_11882,N_11677);
nor U12107 (N_12107,N_11462,N_10954);
xor U12108 (N_12108,N_10960,N_11888);
xor U12109 (N_12109,N_11581,N_10915);
nand U12110 (N_12110,N_11712,N_11666);
xnor U12111 (N_12111,N_10975,N_11540);
or U12112 (N_12112,N_11385,N_11646);
xor U12113 (N_12113,N_11403,N_11640);
or U12114 (N_12114,N_11939,N_11399);
nand U12115 (N_12115,N_11508,N_10880);
and U12116 (N_12116,N_10938,N_11699);
xor U12117 (N_12117,N_11672,N_10898);
and U12118 (N_12118,N_11217,N_11448);
or U12119 (N_12119,N_10984,N_10978);
or U12120 (N_12120,N_11255,N_11580);
or U12121 (N_12121,N_11472,N_11126);
nor U12122 (N_12122,N_11167,N_10824);
and U12123 (N_12123,N_11248,N_11660);
nor U12124 (N_12124,N_11971,N_11595);
and U12125 (N_12125,N_10961,N_11519);
and U12126 (N_12126,N_10883,N_11206);
nand U12127 (N_12127,N_11445,N_11079);
and U12128 (N_12128,N_11793,N_11935);
xnor U12129 (N_12129,N_11435,N_10801);
nand U12130 (N_12130,N_11328,N_11026);
nor U12131 (N_12131,N_11363,N_11618);
or U12132 (N_12132,N_11713,N_11017);
and U12133 (N_12133,N_11121,N_10931);
and U12134 (N_12134,N_11310,N_11763);
or U12135 (N_12135,N_11528,N_11516);
xor U12136 (N_12136,N_11686,N_11298);
xor U12137 (N_12137,N_11187,N_11915);
and U12138 (N_12138,N_11043,N_11252);
or U12139 (N_12139,N_11947,N_11729);
nor U12140 (N_12140,N_10935,N_11558);
or U12141 (N_12141,N_11049,N_11998);
xor U12142 (N_12142,N_11180,N_11259);
or U12143 (N_12143,N_11765,N_11406);
and U12144 (N_12144,N_10843,N_11068);
nor U12145 (N_12145,N_10879,N_11930);
nor U12146 (N_12146,N_11344,N_10998);
nand U12147 (N_12147,N_11053,N_11182);
nor U12148 (N_12148,N_11957,N_11780);
xnor U12149 (N_12149,N_10948,N_11896);
xor U12150 (N_12150,N_11254,N_11185);
nor U12151 (N_12151,N_11201,N_11829);
or U12152 (N_12152,N_11323,N_10856);
nand U12153 (N_12153,N_11837,N_11892);
nor U12154 (N_12154,N_11671,N_11211);
xnor U12155 (N_12155,N_10885,N_11082);
and U12156 (N_12156,N_11487,N_10897);
or U12157 (N_12157,N_11670,N_11542);
nor U12158 (N_12158,N_11941,N_11718);
and U12159 (N_12159,N_11058,N_11750);
nor U12160 (N_12160,N_11860,N_10991);
nand U12161 (N_12161,N_11280,N_11365);
or U12162 (N_12162,N_11442,N_11952);
xor U12163 (N_12163,N_11227,N_11940);
nor U12164 (N_12164,N_10927,N_11883);
nor U12165 (N_12165,N_11798,N_11929);
nand U12166 (N_12166,N_11264,N_11288);
xor U12167 (N_12167,N_11046,N_11863);
and U12168 (N_12168,N_10983,N_11458);
nand U12169 (N_12169,N_11865,N_11911);
nor U12170 (N_12170,N_11358,N_11530);
nor U12171 (N_12171,N_10850,N_11578);
xor U12172 (N_12172,N_11716,N_11212);
nor U12173 (N_12173,N_11691,N_11613);
nor U12174 (N_12174,N_10882,N_11577);
nor U12175 (N_12175,N_11683,N_11536);
nor U12176 (N_12176,N_11014,N_11286);
and U12177 (N_12177,N_10980,N_11975);
nor U12178 (N_12178,N_11013,N_11384);
nor U12179 (N_12179,N_10893,N_11515);
xnor U12180 (N_12180,N_11658,N_11456);
or U12181 (N_12181,N_11372,N_11551);
nand U12182 (N_12182,N_11692,N_11795);
or U12183 (N_12183,N_10876,N_11166);
xnor U12184 (N_12184,N_11493,N_11431);
and U12185 (N_12185,N_11282,N_11107);
nor U12186 (N_12186,N_11420,N_11546);
xnor U12187 (N_12187,N_11918,N_11535);
xor U12188 (N_12188,N_11181,N_11590);
and U12189 (N_12189,N_10838,N_11785);
xor U12190 (N_12190,N_11060,N_11539);
and U12191 (N_12191,N_11875,N_11510);
xor U12192 (N_12192,N_11877,N_11944);
nand U12193 (N_12193,N_11447,N_11740);
and U12194 (N_12194,N_11574,N_11809);
and U12195 (N_12195,N_11025,N_11300);
xor U12196 (N_12196,N_11015,N_11566);
and U12197 (N_12197,N_11522,N_11619);
nand U12198 (N_12198,N_11348,N_10806);
xor U12199 (N_12199,N_11923,N_10877);
and U12200 (N_12200,N_11802,N_11767);
nand U12201 (N_12201,N_11127,N_10926);
or U12202 (N_12202,N_11063,N_10917);
nand U12203 (N_12203,N_11925,N_11113);
and U12204 (N_12204,N_11949,N_11512);
and U12205 (N_12205,N_11204,N_11317);
xor U12206 (N_12206,N_11656,N_11313);
and U12207 (N_12207,N_11596,N_11159);
or U12208 (N_12208,N_11021,N_11123);
or U12209 (N_12209,N_10911,N_11390);
nor U12210 (N_12210,N_11325,N_10950);
xnor U12211 (N_12211,N_11553,N_11102);
nand U12212 (N_12212,N_11138,N_11964);
nand U12213 (N_12213,N_11847,N_11851);
nand U12214 (N_12214,N_11093,N_11823);
or U12215 (N_12215,N_11638,N_11174);
or U12216 (N_12216,N_11615,N_11766);
xor U12217 (N_12217,N_11215,N_11150);
or U12218 (N_12218,N_11018,N_11205);
nand U12219 (N_12219,N_11848,N_10842);
or U12220 (N_12220,N_11426,N_11523);
or U12221 (N_12221,N_10818,N_11130);
or U12222 (N_12222,N_11684,N_11748);
nand U12223 (N_12223,N_11057,N_11826);
nand U12224 (N_12224,N_11491,N_11168);
and U12225 (N_12225,N_11091,N_11706);
nand U12226 (N_12226,N_10982,N_11597);
nor U12227 (N_12227,N_11778,N_11122);
xor U12228 (N_12228,N_11913,N_11634);
and U12229 (N_12229,N_11956,N_11903);
nand U12230 (N_12230,N_11312,N_11813);
and U12231 (N_12231,N_10862,N_11866);
and U12232 (N_12232,N_11904,N_11315);
and U12233 (N_12233,N_11376,N_11999);
nor U12234 (N_12234,N_11128,N_10802);
nor U12235 (N_12235,N_11816,N_10881);
xor U12236 (N_12236,N_11924,N_11855);
nor U12237 (N_12237,N_11019,N_10928);
nor U12238 (N_12238,N_11318,N_11583);
nor U12239 (N_12239,N_11867,N_11352);
nand U12240 (N_12240,N_11507,N_10994);
nand U12241 (N_12241,N_11649,N_11398);
nand U12242 (N_12242,N_11233,N_11346);
or U12243 (N_12243,N_11220,N_11709);
nand U12244 (N_12244,N_11362,N_11997);
nand U12245 (N_12245,N_10890,N_11062);
and U12246 (N_12246,N_11685,N_11486);
nand U12247 (N_12247,N_11152,N_10989);
or U12248 (N_12248,N_11995,N_10906);
nor U12249 (N_12249,N_10835,N_11236);
nand U12250 (N_12250,N_11452,N_11188);
or U12251 (N_12251,N_11591,N_11274);
nand U12252 (N_12252,N_10831,N_10803);
nand U12253 (N_12253,N_10834,N_11096);
and U12254 (N_12254,N_10956,N_11902);
xnor U12255 (N_12255,N_11234,N_11219);
nand U12256 (N_12256,N_10968,N_11322);
and U12257 (N_12257,N_11920,N_11614);
or U12258 (N_12258,N_11587,N_11977);
xnor U12259 (N_12259,N_11477,N_11223);
or U12260 (N_12260,N_11243,N_11917);
and U12261 (N_12261,N_10999,N_11643);
or U12262 (N_12262,N_11293,N_11210);
nand U12263 (N_12263,N_11478,N_11720);
nor U12264 (N_12264,N_10969,N_10937);
xnor U12265 (N_12265,N_11267,N_11351);
xor U12266 (N_12266,N_11876,N_10943);
nand U12267 (N_12267,N_11287,N_11022);
and U12268 (N_12268,N_11943,N_11945);
nand U12269 (N_12269,N_11177,N_11617);
xor U12270 (N_12270,N_11249,N_11679);
nor U12271 (N_12271,N_10833,N_11226);
xnor U12272 (N_12272,N_11045,N_11554);
nor U12273 (N_12273,N_10955,N_11421);
nand U12274 (N_12274,N_11011,N_11576);
or U12275 (N_12275,N_11291,N_11572);
nor U12276 (N_12276,N_11144,N_11443);
and U12277 (N_12277,N_11466,N_11509);
xnor U12278 (N_12278,N_11919,N_11163);
xnor U12279 (N_12279,N_11602,N_11735);
and U12280 (N_12280,N_11601,N_11537);
nand U12281 (N_12281,N_11702,N_11784);
or U12282 (N_12282,N_11616,N_11933);
or U12283 (N_12283,N_11714,N_11650);
or U12284 (N_12284,N_11490,N_11132);
and U12285 (N_12285,N_11307,N_11178);
or U12286 (N_12286,N_11419,N_11834);
xor U12287 (N_12287,N_11885,N_11072);
nand U12288 (N_12288,N_11209,N_10808);
and U12289 (N_12289,N_10963,N_10992);
and U12290 (N_12290,N_11550,N_11786);
xor U12291 (N_12291,N_10837,N_11797);
and U12292 (N_12292,N_10986,N_11849);
nand U12293 (N_12293,N_11588,N_11818);
xnor U12294 (N_12294,N_11457,N_11946);
xnor U12295 (N_12295,N_11474,N_11719);
nor U12296 (N_12296,N_11016,N_11967);
nand U12297 (N_12297,N_11791,N_10940);
and U12298 (N_12298,N_11761,N_11934);
xor U12299 (N_12299,N_11682,N_11199);
xor U12300 (N_12300,N_11739,N_11299);
xnor U12301 (N_12301,N_11175,N_11931);
nor U12302 (N_12302,N_11864,N_11067);
or U12303 (N_12303,N_11982,N_11703);
xnor U12304 (N_12304,N_11721,N_11119);
nor U12305 (N_12305,N_11341,N_11158);
or U12306 (N_12306,N_11357,N_11760);
or U12307 (N_12307,N_10804,N_11141);
and U12308 (N_12308,N_11434,N_11270);
nand U12309 (N_12309,N_10853,N_11470);
or U12310 (N_12310,N_11733,N_10995);
nor U12311 (N_12311,N_11153,N_11526);
and U12312 (N_12312,N_11371,N_11051);
and U12313 (N_12313,N_11584,N_11561);
or U12314 (N_12314,N_11586,N_11543);
or U12315 (N_12315,N_11593,N_11505);
or U12316 (N_12316,N_10889,N_11225);
nor U12317 (N_12317,N_11961,N_11641);
or U12318 (N_12318,N_11483,N_11061);
nand U12319 (N_12319,N_11890,N_11003);
nor U12320 (N_12320,N_10887,N_11803);
xor U12321 (N_12321,N_11356,N_11143);
and U12322 (N_12322,N_11501,N_11753);
xor U12323 (N_12323,N_10809,N_11044);
nor U12324 (N_12324,N_11134,N_11039);
nor U12325 (N_12325,N_11002,N_11630);
xnor U12326 (N_12326,N_10971,N_11573);
and U12327 (N_12327,N_11488,N_11380);
and U12328 (N_12328,N_11984,N_11069);
and U12329 (N_12329,N_11195,N_11081);
and U12330 (N_12330,N_11497,N_11500);
nor U12331 (N_12331,N_11559,N_11052);
nand U12332 (N_12332,N_11870,N_11155);
or U12333 (N_12333,N_11331,N_11375);
nand U12334 (N_12334,N_11804,N_11912);
xor U12335 (N_12335,N_11781,N_11742);
and U12336 (N_12336,N_11789,N_11606);
xnor U12337 (N_12337,N_11241,N_11190);
or U12338 (N_12338,N_11268,N_11942);
nand U12339 (N_12339,N_11193,N_11731);
nand U12340 (N_12340,N_10930,N_11907);
nand U12341 (N_12341,N_11273,N_11036);
xor U12342 (N_12342,N_11030,N_11084);
and U12343 (N_12343,N_11973,N_11518);
and U12344 (N_12344,N_10970,N_11401);
and U12345 (N_12345,N_10910,N_11825);
and U12346 (N_12346,N_11050,N_11446);
nor U12347 (N_12347,N_11404,N_11556);
xor U12348 (N_12348,N_11347,N_11135);
or U12349 (N_12349,N_11575,N_11221);
nor U12350 (N_12350,N_11103,N_11476);
nor U12351 (N_12351,N_11970,N_11749);
nor U12352 (N_12352,N_10813,N_11192);
and U12353 (N_12353,N_10867,N_11652);
nand U12354 (N_12354,N_11308,N_11545);
xor U12355 (N_12355,N_11437,N_11996);
and U12356 (N_12356,N_11297,N_11836);
or U12357 (N_12357,N_11910,N_10959);
and U12358 (N_12358,N_11805,N_11838);
xor U12359 (N_12359,N_11582,N_11668);
nor U12360 (N_12360,N_11071,N_11520);
xnor U12361 (N_12361,N_11757,N_11485);
xor U12362 (N_12362,N_11856,N_11162);
or U12363 (N_12363,N_11858,N_11275);
xnor U12364 (N_12364,N_11407,N_11659);
nor U12365 (N_12365,N_11674,N_10851);
or U12366 (N_12366,N_11146,N_11151);
nor U12367 (N_12367,N_11624,N_11415);
nand U12368 (N_12368,N_11306,N_11411);
nand U12369 (N_12369,N_11854,N_11276);
and U12370 (N_12370,N_11962,N_10817);
nor U12371 (N_12371,N_10952,N_11343);
or U12372 (N_12372,N_10878,N_11794);
and U12373 (N_12373,N_11040,N_11625);
xor U12374 (N_12374,N_11400,N_11833);
nor U12375 (N_12375,N_11261,N_11320);
or U12376 (N_12376,N_10918,N_11628);
and U12377 (N_12377,N_11598,N_11468);
xor U12378 (N_12378,N_11230,N_11042);
or U12379 (N_12379,N_11263,N_11056);
nor U12380 (N_12380,N_11831,N_10903);
nor U12381 (N_12381,N_11690,N_11301);
nand U12382 (N_12382,N_11768,N_11644);
nor U12383 (N_12383,N_11463,N_10870);
nor U12384 (N_12384,N_11820,N_11339);
or U12385 (N_12385,N_11547,N_11228);
nor U12386 (N_12386,N_11633,N_11555);
nor U12387 (N_12387,N_11772,N_11960);
nand U12388 (N_12388,N_11186,N_11862);
xnor U12389 (N_12389,N_11413,N_11094);
and U12390 (N_12390,N_11777,N_11387);
xor U12391 (N_12391,N_11388,N_10847);
nor U12392 (N_12392,N_11133,N_11078);
nor U12393 (N_12393,N_11292,N_11028);
or U12394 (N_12394,N_11808,N_10822);
or U12395 (N_12395,N_11746,N_10951);
xnor U12396 (N_12396,N_11840,N_10913);
and U12397 (N_12397,N_11835,N_10823);
xnor U12398 (N_12398,N_11213,N_11266);
and U12399 (N_12399,N_11986,N_11755);
or U12400 (N_12400,N_11235,N_11076);
nor U12401 (N_12401,N_11383,N_11354);
nor U12402 (N_12402,N_11024,N_11707);
xor U12403 (N_12403,N_11489,N_11377);
nand U12404 (N_12404,N_11156,N_11147);
nand U12405 (N_12405,N_11815,N_11741);
or U12406 (N_12406,N_11438,N_11529);
nand U12407 (N_12407,N_11111,N_11277);
or U12408 (N_12408,N_10899,N_11708);
nand U12409 (N_12409,N_11654,N_11097);
and U12410 (N_12410,N_11965,N_11176);
or U12411 (N_12411,N_11449,N_11285);
nand U12412 (N_12412,N_10934,N_11894);
nand U12413 (N_12413,N_11499,N_10947);
nand U12414 (N_12414,N_10891,N_11305);
or U12415 (N_12415,N_11364,N_11775);
and U12416 (N_12416,N_10912,N_10925);
and U12417 (N_12417,N_11993,N_11031);
nor U12418 (N_12418,N_11416,N_11607);
nand U12419 (N_12419,N_11541,N_11065);
xor U12420 (N_12420,N_10923,N_11402);
and U12421 (N_12421,N_11004,N_11635);
and U12422 (N_12422,N_11758,N_11661);
xor U12423 (N_12423,N_11260,N_10836);
nand U12424 (N_12424,N_11782,N_10973);
nand U12425 (N_12425,N_10896,N_11336);
or U12426 (N_12426,N_11202,N_11909);
or U12427 (N_12427,N_11859,N_11418);
or U12428 (N_12428,N_11099,N_11296);
nor U12429 (N_12429,N_11172,N_11622);
and U12430 (N_12430,N_11513,N_11140);
nor U12431 (N_12431,N_11118,N_10920);
or U12432 (N_12432,N_11754,N_11811);
or U12433 (N_12433,N_11396,N_11319);
nor U12434 (N_12434,N_11484,N_10990);
nand U12435 (N_12435,N_11899,N_11000);
or U12436 (N_12436,N_11284,N_11368);
nor U12437 (N_12437,N_11564,N_11966);
or U12438 (N_12438,N_11878,N_11007);
and U12439 (N_12439,N_11157,N_10993);
and U12440 (N_12440,N_10800,N_11605);
nor U12441 (N_12441,N_10810,N_11075);
or U12442 (N_12442,N_11494,N_11662);
nand U12443 (N_12443,N_11278,N_11450);
and U12444 (N_12444,N_11409,N_11969);
xnor U12445 (N_12445,N_11511,N_10872);
or U12446 (N_12446,N_10841,N_11839);
nand U12447 (N_12447,N_11538,N_11465);
and U12448 (N_12448,N_11637,N_11392);
or U12449 (N_12449,N_11311,N_11035);
and U12450 (N_12450,N_11240,N_11393);
or U12451 (N_12451,N_11408,N_11897);
and U12452 (N_12452,N_11585,N_11955);
and U12453 (N_12453,N_11246,N_11251);
nor U12454 (N_12454,N_11557,N_11092);
and U12455 (N_12455,N_10852,N_11295);
or U12456 (N_12456,N_11980,N_10820);
and U12457 (N_12457,N_11164,N_11531);
and U12458 (N_12458,N_10949,N_11852);
and U12459 (N_12459,N_11822,N_10812);
nor U12460 (N_12460,N_10827,N_11112);
nor U12461 (N_12461,N_11978,N_11821);
or U12462 (N_12462,N_11350,N_10815);
nand U12463 (N_12463,N_10933,N_11830);
or U12464 (N_12464,N_11579,N_11626);
or U12465 (N_12465,N_10869,N_11436);
or U12466 (N_12466,N_11738,N_11090);
nor U12467 (N_12467,N_11337,N_10854);
or U12468 (N_12468,N_10888,N_11697);
and U12469 (N_12469,N_11701,N_10848);
or U12470 (N_12470,N_11023,N_11366);
xnor U12471 (N_12471,N_11262,N_11200);
or U12472 (N_12472,N_10902,N_11938);
xnor U12473 (N_12473,N_11972,N_11694);
nor U12474 (N_12474,N_11762,N_11954);
and U12475 (N_12475,N_11349,N_11665);
nand U12476 (N_12476,N_10825,N_11979);
and U12477 (N_12477,N_11927,N_11807);
or U12478 (N_12478,N_10814,N_11621);
and U12479 (N_12479,N_10807,N_11715);
nor U12480 (N_12480,N_11647,N_10987);
or U12481 (N_12481,N_11717,N_10957);
and U12482 (N_12482,N_10974,N_11054);
xor U12483 (N_12483,N_11229,N_10932);
xnor U12484 (N_12484,N_11994,N_11370);
or U12485 (N_12485,N_11460,N_11774);
and U12486 (N_12486,N_11034,N_11827);
xor U12487 (N_12487,N_11379,N_11242);
nand U12488 (N_12488,N_11790,N_11664);
xor U12489 (N_12489,N_11632,N_10863);
xor U12490 (N_12490,N_11657,N_11841);
or U12491 (N_12491,N_10944,N_11098);
xor U12492 (N_12492,N_10844,N_11636);
and U12493 (N_12493,N_11439,N_11327);
xor U12494 (N_12494,N_11309,N_11145);
xor U12495 (N_12495,N_11868,N_11283);
and U12496 (N_12496,N_11012,N_11874);
xnor U12497 (N_12497,N_11517,N_11330);
and U12498 (N_12498,N_11395,N_11604);
nor U12499 (N_12499,N_11332,N_10901);
xor U12500 (N_12500,N_11020,N_11290);
xnor U12501 (N_12501,N_11627,N_11611);
nor U12502 (N_12502,N_11723,N_11386);
nor U12503 (N_12503,N_11623,N_11333);
or U12504 (N_12504,N_11381,N_10904);
or U12505 (N_12505,N_11901,N_11032);
nor U12506 (N_12506,N_11047,N_11495);
xor U12507 (N_12507,N_11394,N_11673);
nor U12508 (N_12508,N_10886,N_11704);
xor U12509 (N_12509,N_11006,N_11027);
xnor U12510 (N_12510,N_11191,N_11951);
and U12511 (N_12511,N_11360,N_11444);
nand U12512 (N_12512,N_11599,N_11412);
nand U12513 (N_12513,N_11139,N_11983);
nor U12514 (N_12514,N_10816,N_11695);
or U12515 (N_12515,N_11800,N_11441);
xor U12516 (N_12516,N_10874,N_11525);
or U12517 (N_12517,N_11799,N_11705);
nand U12518 (N_12518,N_11428,N_11104);
or U12519 (N_12519,N_11059,N_11981);
nand U12520 (N_12520,N_11751,N_11010);
nand U12521 (N_12521,N_11724,N_11037);
and U12522 (N_12522,N_11005,N_11814);
or U12523 (N_12523,N_11321,N_11073);
and U12524 (N_12524,N_11114,N_11787);
nor U12525 (N_12525,N_11088,N_11991);
nand U12526 (N_12526,N_11471,N_11382);
or U12527 (N_12527,N_11824,N_11129);
nor U12528 (N_12528,N_11569,N_11871);
nor U12529 (N_12529,N_11214,N_10916);
nand U12530 (N_12530,N_11916,N_11770);
nor U12531 (N_12531,N_11033,N_11359);
xnor U12532 (N_12532,N_11534,N_11170);
or U12533 (N_12533,N_11698,N_11038);
or U12534 (N_12534,N_11663,N_11271);
nand U12535 (N_12535,N_11687,N_11120);
nor U12536 (N_12536,N_11001,N_11433);
and U12537 (N_12537,N_11880,N_10828);
nand U12538 (N_12538,N_11725,N_11730);
nand U12539 (N_12539,N_10805,N_11563);
nor U12540 (N_12540,N_11678,N_11086);
nand U12541 (N_12541,N_10972,N_10979);
or U12542 (N_12542,N_11231,N_11218);
nor U12543 (N_12543,N_11696,N_11125);
nand U12544 (N_12544,N_11430,N_11667);
nand U12545 (N_12545,N_11747,N_11648);
xor U12546 (N_12546,N_11655,N_11459);
or U12547 (N_12547,N_11224,N_10962);
xor U12548 (N_12548,N_11303,N_11198);
nand U12549 (N_12549,N_11732,N_11879);
nor U12550 (N_12550,N_11440,N_11100);
or U12551 (N_12551,N_11592,N_11414);
nand U12552 (N_12552,N_11737,N_11921);
nand U12553 (N_12553,N_11425,N_11832);
nor U12554 (N_12554,N_11281,N_10811);
xor U12555 (N_12555,N_11922,N_10988);
nor U12556 (N_12556,N_11391,N_11183);
and U12557 (N_12557,N_11105,N_11239);
or U12558 (N_12558,N_11232,N_11594);
nand U12559 (N_12559,N_11681,N_11070);
or U12560 (N_12560,N_11496,N_10922);
xnor U12561 (N_12561,N_11171,N_10939);
nand U12562 (N_12562,N_11948,N_11928);
or U12563 (N_12563,N_11314,N_11792);
and U12564 (N_12564,N_11845,N_11469);
or U12565 (N_12565,N_11304,N_11294);
nand U12566 (N_12566,N_11693,N_11612);
and U12567 (N_12567,N_11149,N_11169);
and U12568 (N_12568,N_11914,N_11872);
nor U12569 (N_12569,N_11676,N_11549);
and U12570 (N_12570,N_11974,N_11055);
or U12571 (N_12571,N_11895,N_11700);
or U12572 (N_12572,N_10953,N_11846);
or U12573 (N_12573,N_10981,N_11427);
nor U12574 (N_12574,N_11142,N_11269);
nor U12575 (N_12575,N_11562,N_11405);
nand U12576 (N_12576,N_11642,N_11689);
or U12577 (N_12577,N_11095,N_11481);
or U12578 (N_12578,N_11117,N_11968);
nor U12579 (N_12579,N_11326,N_11812);
nor U12580 (N_12580,N_11361,N_11083);
or U12581 (N_12581,N_10858,N_11850);
xnor U12582 (N_12582,N_11148,N_10967);
and U12583 (N_12583,N_10894,N_10846);
nand U12584 (N_12584,N_11801,N_11560);
xnor U12585 (N_12585,N_11989,N_11194);
nand U12586 (N_12586,N_11873,N_11752);
xnor U12587 (N_12587,N_11009,N_11905);
and U12588 (N_12588,N_11891,N_11247);
and U12589 (N_12589,N_10905,N_11389);
and U12590 (N_12590,N_10900,N_11603);
nand U12591 (N_12591,N_11424,N_10914);
nand U12592 (N_12592,N_11074,N_11289);
or U12593 (N_12593,N_10941,N_10892);
and U12594 (N_12594,N_11570,N_11340);
nand U12595 (N_12595,N_10875,N_11355);
xnor U12596 (N_12596,N_11131,N_11378);
nor U12597 (N_12597,N_11085,N_10855);
xnor U12598 (N_12598,N_10873,N_11041);
nand U12599 (N_12599,N_11064,N_10997);
and U12600 (N_12600,N_11784,N_10935);
or U12601 (N_12601,N_10889,N_11647);
and U12602 (N_12602,N_11789,N_11489);
nor U12603 (N_12603,N_11766,N_11919);
nand U12604 (N_12604,N_11726,N_11673);
or U12605 (N_12605,N_10901,N_11824);
or U12606 (N_12606,N_11376,N_11685);
or U12607 (N_12607,N_11954,N_11939);
nor U12608 (N_12608,N_11861,N_11031);
and U12609 (N_12609,N_10910,N_11279);
and U12610 (N_12610,N_11527,N_10948);
nand U12611 (N_12611,N_11739,N_11435);
and U12612 (N_12612,N_11902,N_11569);
or U12613 (N_12613,N_11647,N_11792);
or U12614 (N_12614,N_11866,N_10917);
xor U12615 (N_12615,N_11360,N_11431);
or U12616 (N_12616,N_11529,N_11857);
and U12617 (N_12617,N_11727,N_11589);
xor U12618 (N_12618,N_10855,N_11401);
and U12619 (N_12619,N_11088,N_11828);
nor U12620 (N_12620,N_10847,N_11660);
or U12621 (N_12621,N_10853,N_10949);
nor U12622 (N_12622,N_11755,N_11849);
nor U12623 (N_12623,N_11077,N_11669);
and U12624 (N_12624,N_10928,N_11520);
nand U12625 (N_12625,N_10905,N_11401);
xor U12626 (N_12626,N_11656,N_11104);
or U12627 (N_12627,N_11151,N_11284);
and U12628 (N_12628,N_10820,N_11426);
xor U12629 (N_12629,N_11538,N_11198);
nand U12630 (N_12630,N_11281,N_11160);
xnor U12631 (N_12631,N_10948,N_11327);
or U12632 (N_12632,N_11946,N_10848);
xor U12633 (N_12633,N_11398,N_11548);
nor U12634 (N_12634,N_11390,N_11175);
xnor U12635 (N_12635,N_11665,N_11241);
xor U12636 (N_12636,N_11733,N_10991);
or U12637 (N_12637,N_11036,N_11025);
nand U12638 (N_12638,N_11077,N_11795);
nand U12639 (N_12639,N_11778,N_11982);
xnor U12640 (N_12640,N_11098,N_11449);
nor U12641 (N_12641,N_11243,N_11847);
xnor U12642 (N_12642,N_11704,N_11273);
nand U12643 (N_12643,N_11746,N_11372);
and U12644 (N_12644,N_11447,N_11756);
nor U12645 (N_12645,N_11906,N_11698);
xnor U12646 (N_12646,N_11552,N_11944);
xnor U12647 (N_12647,N_11991,N_10911);
nand U12648 (N_12648,N_10842,N_11207);
nor U12649 (N_12649,N_11611,N_10999);
xnor U12650 (N_12650,N_11965,N_11461);
or U12651 (N_12651,N_11033,N_11994);
xor U12652 (N_12652,N_11444,N_11159);
nor U12653 (N_12653,N_11325,N_11505);
nor U12654 (N_12654,N_11462,N_11673);
and U12655 (N_12655,N_11876,N_11880);
and U12656 (N_12656,N_11792,N_11065);
and U12657 (N_12657,N_11321,N_10909);
nor U12658 (N_12658,N_11263,N_11222);
or U12659 (N_12659,N_11536,N_11099);
or U12660 (N_12660,N_11865,N_11907);
nand U12661 (N_12661,N_11201,N_11780);
and U12662 (N_12662,N_11456,N_11902);
nand U12663 (N_12663,N_11515,N_11475);
and U12664 (N_12664,N_11478,N_11460);
and U12665 (N_12665,N_11092,N_11837);
nor U12666 (N_12666,N_11067,N_11830);
xor U12667 (N_12667,N_11045,N_11314);
and U12668 (N_12668,N_11539,N_11651);
nor U12669 (N_12669,N_10864,N_11127);
and U12670 (N_12670,N_11784,N_11275);
and U12671 (N_12671,N_11690,N_11046);
nand U12672 (N_12672,N_11950,N_11312);
nand U12673 (N_12673,N_11202,N_11860);
nand U12674 (N_12674,N_11043,N_10844);
xnor U12675 (N_12675,N_11947,N_11759);
nor U12676 (N_12676,N_11952,N_11193);
and U12677 (N_12677,N_11111,N_11579);
or U12678 (N_12678,N_10966,N_11141);
xor U12679 (N_12679,N_11351,N_10871);
or U12680 (N_12680,N_11743,N_11828);
nor U12681 (N_12681,N_11983,N_11198);
xnor U12682 (N_12682,N_10920,N_10814);
and U12683 (N_12683,N_11223,N_11979);
nor U12684 (N_12684,N_11535,N_11739);
xor U12685 (N_12685,N_11388,N_11891);
nor U12686 (N_12686,N_11358,N_11894);
nand U12687 (N_12687,N_10921,N_11304);
nor U12688 (N_12688,N_11769,N_11498);
nand U12689 (N_12689,N_11650,N_10978);
or U12690 (N_12690,N_11614,N_10907);
and U12691 (N_12691,N_11717,N_11517);
or U12692 (N_12692,N_11494,N_10922);
or U12693 (N_12693,N_11654,N_11478);
or U12694 (N_12694,N_10846,N_11902);
nand U12695 (N_12695,N_11861,N_11769);
and U12696 (N_12696,N_11185,N_11480);
or U12697 (N_12697,N_11933,N_11637);
nor U12698 (N_12698,N_11903,N_11101);
nand U12699 (N_12699,N_11767,N_10968);
nor U12700 (N_12700,N_11423,N_11997);
or U12701 (N_12701,N_11323,N_11425);
and U12702 (N_12702,N_11747,N_11673);
nand U12703 (N_12703,N_11368,N_11233);
or U12704 (N_12704,N_10991,N_11507);
or U12705 (N_12705,N_11441,N_11093);
nand U12706 (N_12706,N_11462,N_10875);
nor U12707 (N_12707,N_11640,N_11490);
nand U12708 (N_12708,N_11078,N_11496);
nor U12709 (N_12709,N_10957,N_11737);
nor U12710 (N_12710,N_11720,N_11304);
nor U12711 (N_12711,N_11892,N_10888);
or U12712 (N_12712,N_11300,N_11046);
nor U12713 (N_12713,N_10842,N_11248);
and U12714 (N_12714,N_11798,N_11048);
nor U12715 (N_12715,N_11513,N_11894);
nor U12716 (N_12716,N_11385,N_11248);
nand U12717 (N_12717,N_11285,N_10957);
nor U12718 (N_12718,N_11084,N_11367);
or U12719 (N_12719,N_11963,N_11957);
nand U12720 (N_12720,N_11935,N_11509);
or U12721 (N_12721,N_11983,N_11289);
and U12722 (N_12722,N_11036,N_11739);
nand U12723 (N_12723,N_11006,N_11524);
and U12724 (N_12724,N_11195,N_10912);
xor U12725 (N_12725,N_11570,N_11575);
xnor U12726 (N_12726,N_11595,N_10828);
or U12727 (N_12727,N_11705,N_11715);
xnor U12728 (N_12728,N_11017,N_11213);
and U12729 (N_12729,N_10804,N_11236);
xnor U12730 (N_12730,N_11841,N_11392);
xnor U12731 (N_12731,N_11116,N_11247);
nor U12732 (N_12732,N_11255,N_11755);
and U12733 (N_12733,N_11065,N_11306);
or U12734 (N_12734,N_11072,N_11597);
and U12735 (N_12735,N_11360,N_11369);
and U12736 (N_12736,N_11612,N_10961);
or U12737 (N_12737,N_11115,N_11062);
nor U12738 (N_12738,N_11920,N_11165);
or U12739 (N_12739,N_10802,N_11107);
and U12740 (N_12740,N_11170,N_11369);
and U12741 (N_12741,N_11536,N_11934);
and U12742 (N_12742,N_11017,N_11284);
nand U12743 (N_12743,N_10957,N_11101);
xnor U12744 (N_12744,N_11965,N_11082);
nand U12745 (N_12745,N_11207,N_11513);
or U12746 (N_12746,N_10911,N_11446);
nand U12747 (N_12747,N_10861,N_10956);
and U12748 (N_12748,N_11135,N_11821);
nand U12749 (N_12749,N_11554,N_11097);
xor U12750 (N_12750,N_11871,N_11894);
or U12751 (N_12751,N_10988,N_11074);
and U12752 (N_12752,N_11559,N_11981);
nand U12753 (N_12753,N_11290,N_11823);
xnor U12754 (N_12754,N_11968,N_11155);
nor U12755 (N_12755,N_11857,N_11304);
xnor U12756 (N_12756,N_11156,N_11744);
and U12757 (N_12757,N_10844,N_10816);
or U12758 (N_12758,N_10962,N_10855);
nor U12759 (N_12759,N_11157,N_11003);
or U12760 (N_12760,N_11182,N_11586);
and U12761 (N_12761,N_10889,N_11049);
or U12762 (N_12762,N_11519,N_11898);
nor U12763 (N_12763,N_11952,N_11213);
xnor U12764 (N_12764,N_10971,N_11987);
nand U12765 (N_12765,N_11342,N_11651);
xnor U12766 (N_12766,N_11273,N_10888);
nand U12767 (N_12767,N_11890,N_11500);
nand U12768 (N_12768,N_11487,N_11407);
xnor U12769 (N_12769,N_11787,N_11347);
nand U12770 (N_12770,N_11768,N_10854);
nand U12771 (N_12771,N_11681,N_10921);
or U12772 (N_12772,N_11466,N_11870);
xnor U12773 (N_12773,N_11638,N_11218);
nor U12774 (N_12774,N_11654,N_11483);
nor U12775 (N_12775,N_11124,N_11805);
nor U12776 (N_12776,N_11712,N_10858);
and U12777 (N_12777,N_11749,N_11099);
xnor U12778 (N_12778,N_11622,N_11839);
xor U12779 (N_12779,N_10999,N_11023);
nor U12780 (N_12780,N_10974,N_10817);
nand U12781 (N_12781,N_11415,N_10837);
nor U12782 (N_12782,N_11536,N_11056);
and U12783 (N_12783,N_11084,N_11960);
nor U12784 (N_12784,N_11972,N_11628);
nand U12785 (N_12785,N_11925,N_11417);
xor U12786 (N_12786,N_11023,N_11320);
nand U12787 (N_12787,N_11468,N_11193);
nand U12788 (N_12788,N_11181,N_10836);
and U12789 (N_12789,N_11555,N_10931);
nor U12790 (N_12790,N_11067,N_11302);
nand U12791 (N_12791,N_10906,N_11354);
xor U12792 (N_12792,N_10989,N_10877);
xnor U12793 (N_12793,N_11416,N_11496);
or U12794 (N_12794,N_11820,N_11261);
nor U12795 (N_12795,N_11141,N_11860);
nand U12796 (N_12796,N_11079,N_11973);
nand U12797 (N_12797,N_11154,N_11312);
nand U12798 (N_12798,N_11036,N_11623);
or U12799 (N_12799,N_11128,N_10998);
or U12800 (N_12800,N_11207,N_11573);
nand U12801 (N_12801,N_10836,N_11230);
nor U12802 (N_12802,N_11800,N_11701);
nand U12803 (N_12803,N_11156,N_11586);
or U12804 (N_12804,N_11099,N_11178);
nand U12805 (N_12805,N_11179,N_11167);
and U12806 (N_12806,N_11986,N_11677);
and U12807 (N_12807,N_11030,N_11963);
or U12808 (N_12808,N_11628,N_10859);
and U12809 (N_12809,N_11610,N_11112);
nand U12810 (N_12810,N_11996,N_10920);
nand U12811 (N_12811,N_11835,N_11150);
or U12812 (N_12812,N_11282,N_11268);
xnor U12813 (N_12813,N_11194,N_11431);
or U12814 (N_12814,N_11472,N_10993);
nor U12815 (N_12815,N_11181,N_11051);
nor U12816 (N_12816,N_11181,N_10908);
and U12817 (N_12817,N_11940,N_11996);
nor U12818 (N_12818,N_11503,N_11062);
or U12819 (N_12819,N_11412,N_11489);
and U12820 (N_12820,N_11367,N_11148);
or U12821 (N_12821,N_11736,N_10963);
nor U12822 (N_12822,N_11531,N_11342);
nor U12823 (N_12823,N_11159,N_11287);
nand U12824 (N_12824,N_11295,N_11240);
or U12825 (N_12825,N_11806,N_11847);
nand U12826 (N_12826,N_11270,N_11290);
xnor U12827 (N_12827,N_11694,N_11380);
or U12828 (N_12828,N_11095,N_10893);
nor U12829 (N_12829,N_10805,N_11938);
or U12830 (N_12830,N_11978,N_11774);
and U12831 (N_12831,N_11038,N_10875);
nand U12832 (N_12832,N_11533,N_11192);
nor U12833 (N_12833,N_11226,N_10869);
nand U12834 (N_12834,N_10954,N_11689);
or U12835 (N_12835,N_11245,N_11412);
nor U12836 (N_12836,N_11479,N_11505);
nand U12837 (N_12837,N_11506,N_10841);
and U12838 (N_12838,N_11918,N_11444);
or U12839 (N_12839,N_10992,N_11429);
xor U12840 (N_12840,N_11326,N_10951);
xnor U12841 (N_12841,N_11964,N_11175);
nand U12842 (N_12842,N_10838,N_11752);
or U12843 (N_12843,N_11547,N_11733);
or U12844 (N_12844,N_11546,N_11586);
nand U12845 (N_12845,N_11591,N_11512);
nand U12846 (N_12846,N_11743,N_11621);
xor U12847 (N_12847,N_11944,N_10813);
nor U12848 (N_12848,N_10894,N_11732);
and U12849 (N_12849,N_10990,N_11843);
nor U12850 (N_12850,N_11414,N_11670);
nor U12851 (N_12851,N_10936,N_11074);
nor U12852 (N_12852,N_11777,N_11318);
or U12853 (N_12853,N_11066,N_11758);
nand U12854 (N_12854,N_11536,N_11250);
or U12855 (N_12855,N_10822,N_10858);
nand U12856 (N_12856,N_11116,N_10863);
or U12857 (N_12857,N_11505,N_11128);
or U12858 (N_12858,N_11423,N_10928);
nor U12859 (N_12859,N_11439,N_11869);
nand U12860 (N_12860,N_11352,N_11860);
and U12861 (N_12861,N_10912,N_11650);
nor U12862 (N_12862,N_11486,N_10962);
nand U12863 (N_12863,N_10892,N_11078);
and U12864 (N_12864,N_11948,N_11192);
and U12865 (N_12865,N_11099,N_11339);
nand U12866 (N_12866,N_11079,N_11297);
or U12867 (N_12867,N_10951,N_11915);
xnor U12868 (N_12868,N_11881,N_11557);
xor U12869 (N_12869,N_11670,N_11882);
nor U12870 (N_12870,N_11332,N_11006);
nor U12871 (N_12871,N_10950,N_11239);
nand U12872 (N_12872,N_10978,N_11445);
xor U12873 (N_12873,N_11165,N_11750);
or U12874 (N_12874,N_11401,N_11883);
nor U12875 (N_12875,N_11670,N_10922);
nand U12876 (N_12876,N_11269,N_10878);
nand U12877 (N_12877,N_11965,N_11181);
and U12878 (N_12878,N_10891,N_11622);
xnor U12879 (N_12879,N_11627,N_11936);
and U12880 (N_12880,N_11885,N_11787);
or U12881 (N_12881,N_11320,N_11260);
and U12882 (N_12882,N_11576,N_11431);
or U12883 (N_12883,N_11583,N_11090);
xor U12884 (N_12884,N_11806,N_11300);
or U12885 (N_12885,N_11817,N_11862);
or U12886 (N_12886,N_11939,N_11890);
nor U12887 (N_12887,N_11058,N_11460);
or U12888 (N_12888,N_11311,N_11501);
or U12889 (N_12889,N_11903,N_11614);
xnor U12890 (N_12890,N_11858,N_11482);
and U12891 (N_12891,N_11602,N_11375);
or U12892 (N_12892,N_11556,N_11958);
nor U12893 (N_12893,N_11965,N_10813);
nand U12894 (N_12894,N_10868,N_11177);
and U12895 (N_12895,N_11359,N_11689);
nor U12896 (N_12896,N_11636,N_11841);
or U12897 (N_12897,N_11648,N_11231);
and U12898 (N_12898,N_11065,N_11548);
nor U12899 (N_12899,N_11083,N_11542);
nor U12900 (N_12900,N_11033,N_10886);
nor U12901 (N_12901,N_11897,N_10872);
or U12902 (N_12902,N_10979,N_11844);
xnor U12903 (N_12903,N_11829,N_11749);
nor U12904 (N_12904,N_11245,N_10899);
xnor U12905 (N_12905,N_11285,N_11806);
nor U12906 (N_12906,N_11694,N_11171);
xnor U12907 (N_12907,N_11018,N_11173);
xor U12908 (N_12908,N_11142,N_11186);
nand U12909 (N_12909,N_11931,N_11148);
or U12910 (N_12910,N_10800,N_11885);
or U12911 (N_12911,N_11676,N_11074);
xnor U12912 (N_12912,N_11927,N_11583);
xnor U12913 (N_12913,N_11493,N_11162);
nand U12914 (N_12914,N_11667,N_11575);
xor U12915 (N_12915,N_11791,N_11883);
xor U12916 (N_12916,N_11531,N_11385);
nand U12917 (N_12917,N_11850,N_11105);
nor U12918 (N_12918,N_11236,N_11367);
nor U12919 (N_12919,N_11875,N_11661);
nand U12920 (N_12920,N_11050,N_11838);
nor U12921 (N_12921,N_11090,N_11089);
xor U12922 (N_12922,N_10849,N_11878);
or U12923 (N_12923,N_11527,N_11666);
nand U12924 (N_12924,N_11239,N_11017);
nand U12925 (N_12925,N_10882,N_11454);
nor U12926 (N_12926,N_11858,N_11496);
xor U12927 (N_12927,N_11918,N_11825);
nor U12928 (N_12928,N_11330,N_10911);
or U12929 (N_12929,N_11690,N_11390);
xnor U12930 (N_12930,N_10944,N_11596);
nor U12931 (N_12931,N_11938,N_10859);
xnor U12932 (N_12932,N_11413,N_10979);
and U12933 (N_12933,N_11169,N_11268);
xor U12934 (N_12934,N_11980,N_11491);
and U12935 (N_12935,N_11034,N_10916);
xnor U12936 (N_12936,N_11494,N_10903);
and U12937 (N_12937,N_11015,N_10906);
and U12938 (N_12938,N_11350,N_10989);
nor U12939 (N_12939,N_11019,N_11076);
xor U12940 (N_12940,N_11871,N_11714);
nor U12941 (N_12941,N_11915,N_10868);
nor U12942 (N_12942,N_11002,N_11700);
and U12943 (N_12943,N_11086,N_11063);
nand U12944 (N_12944,N_11017,N_10810);
or U12945 (N_12945,N_11948,N_11111);
or U12946 (N_12946,N_11300,N_11618);
nor U12947 (N_12947,N_11761,N_11884);
nor U12948 (N_12948,N_11110,N_11897);
and U12949 (N_12949,N_10884,N_11882);
nor U12950 (N_12950,N_11794,N_11484);
xor U12951 (N_12951,N_10929,N_11532);
and U12952 (N_12952,N_10951,N_10957);
and U12953 (N_12953,N_11280,N_11432);
and U12954 (N_12954,N_11196,N_11036);
and U12955 (N_12955,N_11377,N_11702);
or U12956 (N_12956,N_11357,N_11827);
xor U12957 (N_12957,N_11892,N_11962);
and U12958 (N_12958,N_11673,N_11408);
and U12959 (N_12959,N_11498,N_11651);
or U12960 (N_12960,N_11617,N_11705);
nand U12961 (N_12961,N_10947,N_11291);
and U12962 (N_12962,N_11984,N_11974);
nand U12963 (N_12963,N_11375,N_11045);
nor U12964 (N_12964,N_10860,N_11472);
xor U12965 (N_12965,N_11014,N_11114);
nand U12966 (N_12966,N_11775,N_11905);
and U12967 (N_12967,N_11174,N_11034);
xor U12968 (N_12968,N_10888,N_11181);
xor U12969 (N_12969,N_10970,N_11632);
or U12970 (N_12970,N_11619,N_11555);
nor U12971 (N_12971,N_11079,N_11584);
nor U12972 (N_12972,N_10819,N_11134);
nand U12973 (N_12973,N_11797,N_11387);
nand U12974 (N_12974,N_10873,N_11990);
or U12975 (N_12975,N_11243,N_11866);
nor U12976 (N_12976,N_10925,N_11682);
xor U12977 (N_12977,N_11040,N_11120);
nand U12978 (N_12978,N_11423,N_11719);
and U12979 (N_12979,N_11957,N_11532);
xor U12980 (N_12980,N_11698,N_11445);
nor U12981 (N_12981,N_10925,N_11393);
nor U12982 (N_12982,N_11754,N_11265);
nand U12983 (N_12983,N_11363,N_11423);
nand U12984 (N_12984,N_10907,N_11581);
nor U12985 (N_12985,N_11086,N_10988);
nor U12986 (N_12986,N_10950,N_11760);
xor U12987 (N_12987,N_11916,N_10951);
nor U12988 (N_12988,N_11309,N_11952);
or U12989 (N_12989,N_11217,N_11869);
or U12990 (N_12990,N_11988,N_11671);
nand U12991 (N_12991,N_10952,N_10922);
xor U12992 (N_12992,N_10970,N_11081);
nand U12993 (N_12993,N_11178,N_11354);
xnor U12994 (N_12994,N_11420,N_11834);
xor U12995 (N_12995,N_11509,N_11347);
nand U12996 (N_12996,N_11198,N_11141);
and U12997 (N_12997,N_11440,N_11992);
or U12998 (N_12998,N_11337,N_11930);
xor U12999 (N_12999,N_11225,N_11982);
xnor U13000 (N_13000,N_10885,N_10913);
xor U13001 (N_13001,N_11992,N_10942);
nand U13002 (N_13002,N_10840,N_10975);
xnor U13003 (N_13003,N_11334,N_11053);
nand U13004 (N_13004,N_11261,N_11905);
nor U13005 (N_13005,N_11633,N_11752);
or U13006 (N_13006,N_11147,N_11390);
xnor U13007 (N_13007,N_11074,N_11341);
nand U13008 (N_13008,N_11282,N_11362);
nor U13009 (N_13009,N_10910,N_11170);
nand U13010 (N_13010,N_10904,N_11084);
nor U13011 (N_13011,N_10947,N_11787);
xnor U13012 (N_13012,N_10865,N_10804);
nor U13013 (N_13013,N_11838,N_11128);
or U13014 (N_13014,N_11513,N_11344);
or U13015 (N_13015,N_10804,N_11022);
xnor U13016 (N_13016,N_11279,N_11251);
nand U13017 (N_13017,N_10984,N_11594);
xor U13018 (N_13018,N_10984,N_11561);
xnor U13019 (N_13019,N_11034,N_11620);
and U13020 (N_13020,N_11802,N_10993);
or U13021 (N_13021,N_11521,N_11476);
nand U13022 (N_13022,N_11725,N_11796);
and U13023 (N_13023,N_11430,N_11009);
xor U13024 (N_13024,N_11499,N_11632);
nand U13025 (N_13025,N_11286,N_11151);
nand U13026 (N_13026,N_11569,N_11472);
and U13027 (N_13027,N_11460,N_11323);
nand U13028 (N_13028,N_11872,N_10882);
and U13029 (N_13029,N_11769,N_11385);
or U13030 (N_13030,N_11191,N_11755);
xor U13031 (N_13031,N_11408,N_11850);
nor U13032 (N_13032,N_11084,N_11515);
xor U13033 (N_13033,N_11209,N_11454);
or U13034 (N_13034,N_10974,N_11343);
and U13035 (N_13035,N_11112,N_11234);
xor U13036 (N_13036,N_11767,N_11663);
or U13037 (N_13037,N_11508,N_11848);
nand U13038 (N_13038,N_11286,N_10881);
xor U13039 (N_13039,N_11728,N_11430);
nand U13040 (N_13040,N_11912,N_11299);
nor U13041 (N_13041,N_11377,N_11432);
nand U13042 (N_13042,N_11901,N_11108);
nand U13043 (N_13043,N_10961,N_11385);
or U13044 (N_13044,N_11017,N_10947);
and U13045 (N_13045,N_11960,N_11757);
nor U13046 (N_13046,N_11947,N_11932);
xor U13047 (N_13047,N_11704,N_11558);
nand U13048 (N_13048,N_11353,N_11889);
nor U13049 (N_13049,N_11330,N_11153);
nor U13050 (N_13050,N_10976,N_11928);
nor U13051 (N_13051,N_11939,N_11547);
or U13052 (N_13052,N_11535,N_11812);
nor U13053 (N_13053,N_11968,N_10892);
xor U13054 (N_13054,N_11383,N_10887);
nand U13055 (N_13055,N_11564,N_11842);
xnor U13056 (N_13056,N_10847,N_10954);
nand U13057 (N_13057,N_10806,N_11905);
nor U13058 (N_13058,N_11879,N_11490);
and U13059 (N_13059,N_11095,N_10839);
nor U13060 (N_13060,N_11850,N_11964);
nor U13061 (N_13061,N_10980,N_11313);
xnor U13062 (N_13062,N_11231,N_11116);
nor U13063 (N_13063,N_11043,N_11357);
or U13064 (N_13064,N_10939,N_10926);
nor U13065 (N_13065,N_11201,N_11499);
xor U13066 (N_13066,N_11254,N_11707);
or U13067 (N_13067,N_11244,N_10974);
nand U13068 (N_13068,N_11512,N_11088);
xnor U13069 (N_13069,N_11551,N_11059);
nor U13070 (N_13070,N_11660,N_11024);
nor U13071 (N_13071,N_11979,N_11383);
nor U13072 (N_13072,N_11759,N_11427);
or U13073 (N_13073,N_11930,N_11170);
or U13074 (N_13074,N_10858,N_10948);
or U13075 (N_13075,N_11110,N_10813);
or U13076 (N_13076,N_10915,N_11938);
and U13077 (N_13077,N_10944,N_11440);
xor U13078 (N_13078,N_11077,N_11133);
xor U13079 (N_13079,N_11838,N_11732);
or U13080 (N_13080,N_11158,N_11687);
nor U13081 (N_13081,N_11195,N_11828);
nand U13082 (N_13082,N_11270,N_11069);
nand U13083 (N_13083,N_11481,N_11655);
xor U13084 (N_13084,N_10917,N_11009);
nor U13085 (N_13085,N_11703,N_11590);
xor U13086 (N_13086,N_11827,N_11027);
nand U13087 (N_13087,N_11886,N_11530);
nand U13088 (N_13088,N_11553,N_11126);
nand U13089 (N_13089,N_11624,N_11104);
xnor U13090 (N_13090,N_11478,N_11841);
xnor U13091 (N_13091,N_11978,N_10856);
nor U13092 (N_13092,N_11154,N_11134);
or U13093 (N_13093,N_11788,N_11437);
nand U13094 (N_13094,N_11797,N_11338);
or U13095 (N_13095,N_11548,N_11674);
nor U13096 (N_13096,N_11341,N_11574);
xnor U13097 (N_13097,N_11330,N_11688);
nand U13098 (N_13098,N_11619,N_10810);
xor U13099 (N_13099,N_11013,N_11335);
and U13100 (N_13100,N_10905,N_11962);
or U13101 (N_13101,N_11619,N_11909);
and U13102 (N_13102,N_11996,N_11224);
or U13103 (N_13103,N_11064,N_11208);
nor U13104 (N_13104,N_11819,N_11556);
xor U13105 (N_13105,N_11663,N_11712);
nand U13106 (N_13106,N_11424,N_11046);
nor U13107 (N_13107,N_11097,N_11600);
nand U13108 (N_13108,N_11924,N_11922);
or U13109 (N_13109,N_11648,N_11167);
and U13110 (N_13110,N_11766,N_11550);
or U13111 (N_13111,N_11610,N_10956);
nand U13112 (N_13112,N_11953,N_10907);
nor U13113 (N_13113,N_11854,N_11076);
nand U13114 (N_13114,N_11410,N_10806);
or U13115 (N_13115,N_10851,N_11865);
xor U13116 (N_13116,N_11715,N_11389);
nand U13117 (N_13117,N_10838,N_11262);
and U13118 (N_13118,N_10962,N_10940);
xnor U13119 (N_13119,N_11633,N_11772);
xnor U13120 (N_13120,N_11993,N_11648);
and U13121 (N_13121,N_11940,N_11435);
nand U13122 (N_13122,N_11684,N_11033);
nor U13123 (N_13123,N_10861,N_11315);
and U13124 (N_13124,N_10810,N_11440);
and U13125 (N_13125,N_11248,N_11824);
nand U13126 (N_13126,N_11230,N_10976);
nand U13127 (N_13127,N_11771,N_11369);
and U13128 (N_13128,N_11856,N_11587);
or U13129 (N_13129,N_11848,N_11516);
or U13130 (N_13130,N_11152,N_11229);
nand U13131 (N_13131,N_10972,N_11372);
nand U13132 (N_13132,N_11355,N_11759);
nor U13133 (N_13133,N_11721,N_11291);
and U13134 (N_13134,N_11795,N_11406);
nand U13135 (N_13135,N_11380,N_11132);
and U13136 (N_13136,N_11868,N_11947);
nor U13137 (N_13137,N_11980,N_11794);
xnor U13138 (N_13138,N_11692,N_11935);
nor U13139 (N_13139,N_10915,N_11104);
or U13140 (N_13140,N_11404,N_11089);
nand U13141 (N_13141,N_11759,N_10999);
xor U13142 (N_13142,N_11091,N_11813);
nor U13143 (N_13143,N_11201,N_10928);
or U13144 (N_13144,N_11377,N_11404);
and U13145 (N_13145,N_10892,N_10901);
or U13146 (N_13146,N_11277,N_11842);
or U13147 (N_13147,N_11278,N_11267);
nand U13148 (N_13148,N_11355,N_10844);
or U13149 (N_13149,N_10931,N_10908);
and U13150 (N_13150,N_11198,N_11949);
or U13151 (N_13151,N_11998,N_11833);
and U13152 (N_13152,N_11967,N_11272);
and U13153 (N_13153,N_10970,N_11362);
and U13154 (N_13154,N_10804,N_11667);
nor U13155 (N_13155,N_11891,N_11887);
nor U13156 (N_13156,N_11600,N_11872);
xnor U13157 (N_13157,N_11303,N_11257);
nand U13158 (N_13158,N_11630,N_10825);
nand U13159 (N_13159,N_11828,N_11922);
xnor U13160 (N_13160,N_11458,N_11514);
nand U13161 (N_13161,N_11369,N_11448);
nand U13162 (N_13162,N_10946,N_11847);
nand U13163 (N_13163,N_11854,N_11534);
nand U13164 (N_13164,N_11880,N_11760);
xnor U13165 (N_13165,N_11448,N_11972);
or U13166 (N_13166,N_11334,N_10818);
nand U13167 (N_13167,N_11090,N_11402);
and U13168 (N_13168,N_11351,N_11926);
nor U13169 (N_13169,N_11181,N_10880);
and U13170 (N_13170,N_11934,N_10848);
nor U13171 (N_13171,N_11383,N_10935);
or U13172 (N_13172,N_11173,N_11424);
and U13173 (N_13173,N_11349,N_11294);
xor U13174 (N_13174,N_11222,N_11230);
xnor U13175 (N_13175,N_10841,N_11899);
nand U13176 (N_13176,N_11711,N_10831);
xnor U13177 (N_13177,N_11064,N_11234);
xor U13178 (N_13178,N_11896,N_11877);
nor U13179 (N_13179,N_11420,N_11169);
nand U13180 (N_13180,N_11573,N_10879);
nor U13181 (N_13181,N_11918,N_11355);
nand U13182 (N_13182,N_10944,N_11739);
nor U13183 (N_13183,N_11228,N_11125);
or U13184 (N_13184,N_11015,N_11595);
and U13185 (N_13185,N_11281,N_10836);
xor U13186 (N_13186,N_11296,N_11098);
nand U13187 (N_13187,N_11974,N_11203);
or U13188 (N_13188,N_11525,N_11458);
and U13189 (N_13189,N_11584,N_11422);
and U13190 (N_13190,N_11335,N_11940);
or U13191 (N_13191,N_10916,N_10854);
nand U13192 (N_13192,N_10904,N_11380);
nor U13193 (N_13193,N_11254,N_11657);
and U13194 (N_13194,N_10924,N_11008);
xor U13195 (N_13195,N_11553,N_11825);
or U13196 (N_13196,N_10983,N_11607);
nor U13197 (N_13197,N_11805,N_11581);
xor U13198 (N_13198,N_11837,N_11999);
nand U13199 (N_13199,N_10968,N_11559);
nand U13200 (N_13200,N_12498,N_12574);
nand U13201 (N_13201,N_12112,N_12292);
or U13202 (N_13202,N_12225,N_12944);
nand U13203 (N_13203,N_12061,N_12911);
and U13204 (N_13204,N_12862,N_12737);
nor U13205 (N_13205,N_12321,N_12833);
or U13206 (N_13206,N_12961,N_12098);
or U13207 (N_13207,N_12805,N_12053);
nand U13208 (N_13208,N_12883,N_12204);
xor U13209 (N_13209,N_12629,N_12210);
and U13210 (N_13210,N_12764,N_12712);
or U13211 (N_13211,N_12155,N_12298);
nand U13212 (N_13212,N_12234,N_13171);
nand U13213 (N_13213,N_12845,N_12886);
or U13214 (N_13214,N_12227,N_12280);
and U13215 (N_13215,N_12624,N_13183);
nor U13216 (N_13216,N_12897,N_13056);
nor U13217 (N_13217,N_12362,N_13094);
nor U13218 (N_13218,N_12487,N_12311);
xor U13219 (N_13219,N_12054,N_12882);
nor U13220 (N_13220,N_12465,N_12668);
and U13221 (N_13221,N_12790,N_12052);
and U13222 (N_13222,N_12994,N_13083);
and U13223 (N_13223,N_12593,N_12476);
xor U13224 (N_13224,N_12508,N_12929);
nand U13225 (N_13225,N_12426,N_12720);
nand U13226 (N_13226,N_12735,N_13103);
or U13227 (N_13227,N_12938,N_12050);
nand U13228 (N_13228,N_13159,N_12137);
nand U13229 (N_13229,N_12603,N_12524);
and U13230 (N_13230,N_12519,N_12307);
nor U13231 (N_13231,N_12041,N_12209);
nor U13232 (N_13232,N_12653,N_13121);
and U13233 (N_13233,N_12374,N_12043);
and U13234 (N_13234,N_12654,N_12433);
and U13235 (N_13235,N_12088,N_12934);
nor U13236 (N_13236,N_12305,N_12147);
or U13237 (N_13237,N_12384,N_12449);
or U13238 (N_13238,N_12471,N_12100);
and U13239 (N_13239,N_12528,N_12446);
or U13240 (N_13240,N_12847,N_12564);
and U13241 (N_13241,N_12985,N_13130);
and U13242 (N_13242,N_12729,N_12756);
nand U13243 (N_13243,N_12804,N_12576);
or U13244 (N_13244,N_12551,N_12191);
nor U13245 (N_13245,N_12345,N_12690);
xor U13246 (N_13246,N_12027,N_12327);
nor U13247 (N_13247,N_12024,N_12424);
nor U13248 (N_13248,N_12419,N_12830);
nor U13249 (N_13249,N_12232,N_12279);
nor U13250 (N_13250,N_13093,N_12349);
xnor U13251 (N_13251,N_12208,N_13075);
or U13252 (N_13252,N_12365,N_12778);
or U13253 (N_13253,N_12352,N_12417);
and U13254 (N_13254,N_13125,N_12219);
xnor U13255 (N_13255,N_12565,N_12109);
nand U13256 (N_13256,N_12619,N_13179);
xor U13257 (N_13257,N_12108,N_12107);
or U13258 (N_13258,N_12399,N_12910);
and U13259 (N_13259,N_12990,N_12829);
and U13260 (N_13260,N_13185,N_12730);
xnor U13261 (N_13261,N_12843,N_12427);
nor U13262 (N_13262,N_12788,N_12135);
and U13263 (N_13263,N_13018,N_12379);
xnor U13264 (N_13264,N_13011,N_12009);
nand U13265 (N_13265,N_12981,N_12706);
and U13266 (N_13266,N_12699,N_12505);
or U13267 (N_13267,N_13104,N_12748);
or U13268 (N_13268,N_13062,N_12262);
xor U13269 (N_13269,N_12033,N_13143);
or U13270 (N_13270,N_12917,N_12357);
nor U13271 (N_13271,N_13055,N_12794);
nor U13272 (N_13272,N_13016,N_12765);
and U13273 (N_13273,N_12138,N_12688);
nand U13274 (N_13274,N_12675,N_12148);
and U13275 (N_13275,N_12233,N_12317);
and U13276 (N_13276,N_12569,N_12587);
nand U13277 (N_13277,N_12451,N_12080);
and U13278 (N_13278,N_12001,N_13110);
nor U13279 (N_13279,N_12895,N_12295);
nand U13280 (N_13280,N_12669,N_12622);
and U13281 (N_13281,N_12247,N_12383);
nand U13282 (N_13282,N_12769,N_12812);
or U13283 (N_13283,N_12177,N_12557);
and U13284 (N_13284,N_13137,N_12570);
nor U13285 (N_13285,N_12343,N_12057);
xnor U13286 (N_13286,N_12309,N_12051);
nand U13287 (N_13287,N_12468,N_12578);
or U13288 (N_13288,N_12407,N_12436);
or U13289 (N_13289,N_13024,N_12742);
xor U13290 (N_13290,N_12430,N_12858);
xor U13291 (N_13291,N_12205,N_12531);
and U13292 (N_13292,N_12185,N_12809);
nand U13293 (N_13293,N_12456,N_12122);
or U13294 (N_13294,N_13022,N_13132);
and U13295 (N_13295,N_12579,N_12891);
or U13296 (N_13296,N_13058,N_12650);
nand U13297 (N_13297,N_12784,N_12827);
xor U13298 (N_13298,N_12179,N_12418);
nor U13299 (N_13299,N_12077,N_12752);
and U13300 (N_13300,N_12447,N_12710);
xnor U13301 (N_13301,N_12940,N_13178);
nand U13302 (N_13302,N_12455,N_12034);
and U13303 (N_13303,N_12491,N_12662);
or U13304 (N_13304,N_12063,N_12144);
or U13305 (N_13305,N_12055,N_12517);
nor U13306 (N_13306,N_13184,N_12953);
nand U13307 (N_13307,N_12502,N_12119);
or U13308 (N_13308,N_13161,N_13014);
and U13309 (N_13309,N_13105,N_12873);
nor U13310 (N_13310,N_12242,N_12060);
nand U13311 (N_13311,N_12036,N_12150);
and U13312 (N_13312,N_12116,N_12149);
or U13313 (N_13313,N_12723,N_12416);
and U13314 (N_13314,N_12610,N_12902);
nor U13315 (N_13315,N_13048,N_12297);
nand U13316 (N_13316,N_12585,N_12442);
nand U13317 (N_13317,N_12963,N_12620);
or U13318 (N_13318,N_12773,N_12454);
nand U13319 (N_13319,N_12463,N_13051);
nand U13320 (N_13320,N_12874,N_12967);
nand U13321 (N_13321,N_12721,N_12299);
and U13322 (N_13322,N_12012,N_12350);
nand U13323 (N_13323,N_12779,N_12277);
or U13324 (N_13324,N_12700,N_12923);
or U13325 (N_13325,N_12597,N_13151);
nor U13326 (N_13326,N_12334,N_13067);
xor U13327 (N_13327,N_12615,N_12482);
xor U13328 (N_13328,N_12607,N_12255);
or U13329 (N_13329,N_12397,N_12010);
and U13330 (N_13330,N_12927,N_12583);
xor U13331 (N_13331,N_12022,N_12113);
xnor U13332 (N_13332,N_12821,N_12747);
nand U13333 (N_13333,N_12089,N_12452);
nor U13334 (N_13334,N_13095,N_12134);
xor U13335 (N_13335,N_12448,N_13060);
nand U13336 (N_13336,N_12474,N_12217);
nor U13337 (N_13337,N_12887,N_12393);
nand U13338 (N_13338,N_12796,N_12924);
and U13339 (N_13339,N_12888,N_13124);
xnor U13340 (N_13340,N_13158,N_12868);
xor U13341 (N_13341,N_13101,N_12017);
nor U13342 (N_13342,N_12450,N_12807);
xnor U13343 (N_13343,N_12271,N_12000);
xnor U13344 (N_13344,N_13091,N_12332);
nor U13345 (N_13345,N_13135,N_12102);
and U13346 (N_13346,N_13152,N_12997);
nand U13347 (N_13347,N_13173,N_12406);
nand U13348 (N_13348,N_13133,N_12682);
nand U13349 (N_13349,N_12038,N_13042);
nor U13350 (N_13350,N_12640,N_12328);
nor U13351 (N_13351,N_12029,N_12396);
xnor U13352 (N_13352,N_12866,N_12259);
or U13353 (N_13353,N_12946,N_12340);
nor U13354 (N_13354,N_12475,N_12582);
nand U13355 (N_13355,N_12818,N_12118);
nand U13356 (N_13356,N_12800,N_13144);
or U13357 (N_13357,N_12381,N_12049);
nor U13358 (N_13358,N_13082,N_12839);
nor U13359 (N_13359,N_12440,N_12342);
xor U13360 (N_13360,N_13057,N_12300);
and U13361 (N_13361,N_12285,N_12513);
and U13362 (N_13362,N_12799,N_12670);
xor U13363 (N_13363,N_12453,N_12457);
and U13364 (N_13364,N_12971,N_12376);
and U13365 (N_13365,N_12999,N_12750);
nor U13366 (N_13366,N_12308,N_12534);
and U13367 (N_13367,N_12731,N_13096);
and U13368 (N_13368,N_13072,N_12439);
nor U13369 (N_13369,N_12405,N_12264);
nor U13370 (N_13370,N_12479,N_12473);
or U13371 (N_13371,N_12266,N_12002);
xnor U13372 (N_13372,N_12877,N_12065);
and U13373 (N_13373,N_12364,N_12058);
xor U13374 (N_13374,N_12973,N_12630);
xnor U13375 (N_13375,N_12694,N_12717);
xor U13376 (N_13376,N_13070,N_13197);
nand U13377 (N_13377,N_13068,N_12972);
and U13378 (N_13378,N_12312,N_12951);
and U13379 (N_13379,N_12485,N_12962);
xor U13380 (N_13380,N_12533,N_12166);
nand U13381 (N_13381,N_13112,N_12884);
nor U13382 (N_13382,N_12656,N_12811);
and U13383 (N_13383,N_12532,N_12422);
nand U13384 (N_13384,N_12757,N_12193);
and U13385 (N_13385,N_12443,N_12616);
or U13386 (N_13386,N_12195,N_12703);
nor U13387 (N_13387,N_12728,N_13054);
xor U13388 (N_13388,N_12510,N_12156);
nor U13389 (N_13389,N_12718,N_12361);
nand U13390 (N_13390,N_12636,N_12272);
and U13391 (N_13391,N_12905,N_12339);
xor U13392 (N_13392,N_12791,N_13028);
nand U13393 (N_13393,N_12380,N_12503);
xor U13394 (N_13394,N_12167,N_12127);
nor U13395 (N_13395,N_12499,N_12173);
nor U13396 (N_13396,N_12368,N_13165);
or U13397 (N_13397,N_12254,N_12639);
and U13398 (N_13398,N_13063,N_12207);
and U13399 (N_13399,N_12248,N_12943);
and U13400 (N_13400,N_12310,N_12019);
and U13401 (N_13401,N_12337,N_12995);
nand U13402 (N_13402,N_13041,N_12132);
xor U13403 (N_13403,N_12542,N_12732);
nor U13404 (N_13404,N_12081,N_12320);
and U13405 (N_13405,N_12637,N_12575);
and U13406 (N_13406,N_13079,N_13084);
xnor U13407 (N_13407,N_12992,N_12462);
and U13408 (N_13408,N_12856,N_12664);
nand U13409 (N_13409,N_12850,N_12228);
xnor U13410 (N_13410,N_12875,N_13120);
and U13411 (N_13411,N_12007,N_12776);
nand U13412 (N_13412,N_12025,N_12743);
nor U13413 (N_13413,N_13193,N_13150);
or U13414 (N_13414,N_13102,N_12263);
xor U13415 (N_13415,N_12898,N_12387);
xnor U13416 (N_13416,N_12901,N_13123);
or U13417 (N_13417,N_12908,N_12042);
or U13418 (N_13418,N_12047,N_12226);
or U13419 (N_13419,N_12032,N_12329);
and U13420 (N_13420,N_12993,N_12145);
or U13421 (N_13421,N_12082,N_12642);
xor U13422 (N_13422,N_13186,N_12142);
and U13423 (N_13423,N_12326,N_13046);
xor U13424 (N_13424,N_12618,N_12835);
nor U13425 (N_13425,N_12389,N_12704);
nor U13426 (N_13426,N_12235,N_12644);
nand U13427 (N_13427,N_12168,N_12781);
or U13428 (N_13428,N_12016,N_12023);
xor U13429 (N_13429,N_12527,N_12104);
xnor U13430 (N_13430,N_12558,N_13090);
nor U13431 (N_13431,N_12537,N_12536);
and U13432 (N_13432,N_12628,N_12400);
and U13433 (N_13433,N_12239,N_12657);
xor U13434 (N_13434,N_12880,N_12673);
nor U13435 (N_13435,N_12655,N_13050);
nor U13436 (N_13436,N_12478,N_12702);
nand U13437 (N_13437,N_12870,N_12031);
or U13438 (N_13438,N_12614,N_12714);
nor U13439 (N_13439,N_12562,N_12554);
xnor U13440 (N_13440,N_12079,N_12988);
or U13441 (N_13441,N_12356,N_12170);
nor U13442 (N_13442,N_13169,N_12851);
and U13443 (N_13443,N_12878,N_12236);
and U13444 (N_13444,N_12011,N_12801);
and U13445 (N_13445,N_12813,N_12472);
nor U13446 (N_13446,N_12716,N_13030);
nor U13447 (N_13447,N_12401,N_12955);
or U13448 (N_13448,N_12709,N_12281);
nand U13449 (N_13449,N_13164,N_12826);
xor U13450 (N_13450,N_12093,N_12483);
and U13451 (N_13451,N_12677,N_13032);
nand U13452 (N_13452,N_12005,N_12651);
nand U13453 (N_13453,N_12645,N_12832);
nor U13454 (N_13454,N_13116,N_12896);
or U13455 (N_13455,N_12547,N_12486);
xor U13456 (N_13456,N_13162,N_12529);
and U13457 (N_13457,N_13113,N_12461);
nand U13458 (N_13458,N_12899,N_12931);
nor U13459 (N_13459,N_12283,N_12560);
nor U13460 (N_13460,N_12746,N_13080);
and U13461 (N_13461,N_12488,N_12783);
xor U13462 (N_13462,N_12984,N_12164);
or U13463 (N_13463,N_12759,N_12391);
nor U13464 (N_13464,N_12261,N_13040);
nand U13465 (N_13465,N_12840,N_12431);
xnor U13466 (N_13466,N_12404,N_12838);
nand U13467 (N_13467,N_12187,N_12289);
xnor U13468 (N_13468,N_12606,N_12392);
xor U13469 (N_13469,N_12303,N_12663);
xnor U13470 (N_13470,N_13174,N_12514);
nor U13471 (N_13471,N_12815,N_12493);
nand U13472 (N_13472,N_12692,N_12341);
and U13473 (N_13473,N_12154,N_12083);
and U13474 (N_13474,N_12375,N_12220);
nand U13475 (N_13475,N_12998,N_12871);
and U13476 (N_13476,N_12763,N_13004);
or U13477 (N_13477,N_12111,N_12026);
nor U13478 (N_13478,N_12828,N_12947);
xor U13479 (N_13479,N_12741,N_12608);
nor U13480 (N_13480,N_12561,N_12189);
and U13481 (N_13481,N_12852,N_12385);
or U13482 (N_13482,N_12857,N_12413);
nor U13483 (N_13483,N_13008,N_12894);
nand U13484 (N_13484,N_12099,N_12954);
nand U13485 (N_13485,N_12591,N_13140);
xnor U13486 (N_13486,N_13195,N_12789);
nand U13487 (N_13487,N_12133,N_12192);
or U13488 (N_13488,N_12612,N_13047);
or U13489 (N_13489,N_12398,N_12293);
or U13490 (N_13490,N_12194,N_12035);
and U13491 (N_13491,N_12577,N_12546);
and U13492 (N_13492,N_12360,N_12588);
nand U13493 (N_13493,N_13027,N_12378);
or U13494 (N_13494,N_12056,N_12964);
nand U13495 (N_13495,N_12105,N_12094);
and U13496 (N_13496,N_12495,N_12768);
xnor U13497 (N_13497,N_12627,N_12045);
nor U13498 (N_13498,N_13035,N_12631);
nor U13499 (N_13499,N_12581,N_13023);
or U13500 (N_13500,N_12257,N_12370);
nand U13501 (N_13501,N_12806,N_12250);
nand U13502 (N_13502,N_12315,N_12141);
nand U13503 (N_13503,N_12820,N_12719);
xor U13504 (N_13504,N_12090,N_13122);
nor U13505 (N_13505,N_12872,N_12020);
and U13506 (N_13506,N_12435,N_12237);
nor U13507 (N_13507,N_12190,N_13038);
xnor U13508 (N_13508,N_13196,N_12745);
and U13509 (N_13509,N_12355,N_12124);
nor U13510 (N_13510,N_12958,N_12184);
or U13511 (N_13511,N_12139,N_12975);
or U13512 (N_13512,N_12621,N_12548);
nand U13513 (N_13513,N_13108,N_12904);
nor U13514 (N_13514,N_12296,N_12539);
nand U13515 (N_13515,N_12960,N_12390);
and U13516 (N_13516,N_12733,N_12867);
xnor U13517 (N_13517,N_12347,N_12408);
xor U13518 (N_13518,N_12161,N_12635);
or U13519 (N_13519,N_12460,N_12241);
and U13520 (N_13520,N_12555,N_13085);
or U13521 (N_13521,N_12594,N_12824);
nand U13522 (N_13522,N_12087,N_12649);
and U13523 (N_13523,N_12445,N_12202);
or U13524 (N_13524,N_12331,N_12306);
xor U13525 (N_13525,N_12335,N_12402);
or U13526 (N_13526,N_12535,N_12046);
xor U13527 (N_13527,N_12346,N_12777);
or U13528 (N_13528,N_12101,N_12919);
and U13529 (N_13529,N_12200,N_13087);
or U13530 (N_13530,N_13100,N_12726);
xor U13531 (N_13531,N_12792,N_12921);
nand U13532 (N_13532,N_13044,N_12085);
nand U13533 (N_13533,N_12437,N_12130);
or U13534 (N_13534,N_13025,N_12749);
and U13535 (N_13535,N_12040,N_12751);
xnor U13536 (N_13536,N_12980,N_12667);
and U13537 (N_13537,N_12403,N_13157);
nor U13538 (N_13538,N_12203,N_13010);
nand U13539 (N_13539,N_13129,N_13190);
xnor U13540 (N_13540,N_13127,N_12216);
nor U13541 (N_13541,N_12782,N_12643);
nor U13542 (N_13542,N_13136,N_12222);
and U13543 (N_13543,N_12253,N_12925);
or U13544 (N_13544,N_12013,N_12157);
xnor U13545 (N_13545,N_12808,N_12367);
nand U13546 (N_13546,N_12996,N_13053);
and U13547 (N_13547,N_13145,N_12991);
and U13548 (N_13548,N_12853,N_12595);
or U13549 (N_13549,N_12568,N_12441);
and U13550 (N_13550,N_12836,N_12918);
and U13551 (N_13551,N_12267,N_12125);
nand U13552 (N_13552,N_12273,N_12844);
nand U13553 (N_13553,N_12068,N_12602);
nand U13554 (N_13554,N_12162,N_12775);
nand U13555 (N_13555,N_12611,N_12553);
or U13556 (N_13556,N_12865,N_12952);
and U13557 (N_13557,N_12989,N_12626);
xnor U13558 (N_13558,N_12078,N_12110);
nand U13559 (N_13559,N_13142,N_12623);
and U13560 (N_13560,N_12609,N_12986);
and U13561 (N_13561,N_12916,N_12348);
nand U13562 (N_13562,N_12344,N_12509);
nor U13563 (N_13563,N_13141,N_12722);
nand U13564 (N_13564,N_12666,N_12172);
or U13565 (N_13565,N_12676,N_12143);
nand U13566 (N_13566,N_12698,N_13073);
nor U13567 (N_13567,N_12563,N_12876);
and U13568 (N_13568,N_12686,N_13097);
and U13569 (N_13569,N_12212,N_12915);
nor U13570 (N_13570,N_13076,N_12286);
nor U13571 (N_13571,N_12831,N_12590);
nand U13572 (N_13572,N_12725,N_12516);
xnor U13573 (N_13573,N_12920,N_13098);
xnor U13574 (N_13574,N_12907,N_12206);
nand U13575 (N_13575,N_12260,N_12755);
xor U13576 (N_13576,N_12758,N_12859);
or U13577 (N_13577,N_12846,N_12278);
and U13578 (N_13578,N_12979,N_12841);
xnor U13579 (N_13579,N_12552,N_13119);
xnor U13580 (N_13580,N_13059,N_12176);
or U13581 (N_13581,N_12140,N_13001);
or U13582 (N_13582,N_12268,N_12072);
and U13583 (N_13583,N_12123,N_12825);
or U13584 (N_13584,N_13191,N_12573);
nand U13585 (N_13585,N_12761,N_12304);
or U13586 (N_13586,N_12021,N_12678);
xnor U13587 (N_13587,N_12180,N_13163);
and U13588 (N_13588,N_12214,N_12780);
and U13589 (N_13589,N_12338,N_13033);
xnor U13590 (N_13590,N_12415,N_13181);
or U13591 (N_13591,N_13148,N_12772);
nor U13592 (N_13592,N_12567,N_12363);
and U13593 (N_13593,N_12018,N_12596);
or U13594 (N_13594,N_12652,N_12158);
or U13595 (N_13595,N_12470,N_12970);
nor U13596 (N_13596,N_12889,N_12540);
and U13597 (N_13597,N_12276,N_13109);
nand U13598 (N_13598,N_12945,N_12490);
or U13599 (N_13599,N_13061,N_12674);
xnor U13600 (N_13600,N_12705,N_12282);
nand U13601 (N_13601,N_12238,N_12174);
nor U13602 (N_13602,N_13005,N_13017);
nor U13603 (N_13603,N_13188,N_12231);
or U13604 (N_13604,N_13021,N_12802);
nand U13605 (N_13605,N_12324,N_12196);
xnor U13606 (N_13606,N_12638,N_12302);
nor U13607 (N_13607,N_12518,N_12860);
and U13608 (N_13608,N_12369,N_12968);
and U13609 (N_13609,N_12681,N_12070);
nand U13610 (N_13610,N_12708,N_12956);
xor U13611 (N_13611,N_12641,N_12218);
or U13612 (N_13612,N_12538,N_12942);
and U13613 (N_13613,N_12598,N_13118);
xnor U13614 (N_13614,N_12658,N_12511);
nand U13615 (N_13615,N_12497,N_12601);
nor U13616 (N_13616,N_12974,N_12294);
or U13617 (N_13617,N_12252,N_12388);
nand U13618 (N_13618,N_13199,N_12358);
or U13619 (N_13619,N_12215,N_13149);
and U13620 (N_13620,N_12423,N_12754);
or U13621 (N_13621,N_12837,N_13168);
xnor U13622 (N_13622,N_12062,N_12823);
or U13623 (N_13623,N_12265,N_13111);
xor U13624 (N_13624,N_12541,N_13078);
nor U13625 (N_13625,N_12987,N_12599);
or U13626 (N_13626,N_12854,N_12785);
xnor U13627 (N_13627,N_12323,N_12097);
nor U13628 (N_13628,N_12014,N_12230);
nand U13629 (N_13629,N_12734,N_12477);
nand U13630 (N_13630,N_12128,N_12075);
nand U13631 (N_13631,N_12131,N_13170);
nand U13632 (N_13632,N_12469,N_13043);
nor U13633 (N_13633,N_12171,N_12494);
and U13634 (N_13634,N_13198,N_13106);
xnor U13635 (N_13635,N_12740,N_12169);
nand U13636 (N_13636,N_12030,N_12484);
or U13637 (N_13637,N_12766,N_12633);
nor U13638 (N_13638,N_13006,N_12928);
nand U13639 (N_13639,N_12480,N_12095);
or U13640 (N_13640,N_13117,N_12803);
xnor U13641 (N_13641,N_13189,N_13045);
xnor U13642 (N_13642,N_12004,N_12256);
and U13643 (N_13643,N_13166,N_12774);
or U13644 (N_13644,N_12556,N_12221);
nor U13645 (N_13645,N_12713,N_12114);
or U13646 (N_13646,N_13131,N_12291);
nor U13647 (N_13647,N_12724,N_12507);
xnor U13648 (N_13648,N_12325,N_13128);
or U13649 (N_13649,N_13019,N_12613);
nand U13650 (N_13650,N_12922,N_12977);
or U13651 (N_13651,N_12409,N_12930);
nand U13652 (N_13652,N_13036,N_12738);
and U13653 (N_13653,N_12715,N_12069);
nor U13654 (N_13654,N_13002,N_12333);
xnor U13655 (N_13655,N_12496,N_12600);
or U13656 (N_13656,N_13066,N_12425);
and U13657 (N_13657,N_12377,N_12175);
nand U13658 (N_13658,N_12201,N_12869);
nor U13659 (N_13659,N_12039,N_12848);
xor U13660 (N_13660,N_13088,N_12284);
nand U13661 (N_13661,N_12760,N_12797);
nand U13662 (N_13662,N_12744,N_12589);
nand U13663 (N_13663,N_12522,N_12739);
nor U13664 (N_13664,N_12003,N_12322);
nand U13665 (N_13665,N_12386,N_12545);
nand U13666 (N_13666,N_12855,N_12181);
and U13667 (N_13667,N_12394,N_12313);
and U13668 (N_13668,N_12354,N_12966);
nand U13669 (N_13669,N_12251,N_12696);
nand U13670 (N_13670,N_13155,N_13077);
xnor U13671 (N_13671,N_12672,N_12625);
nand U13672 (N_13672,N_13194,N_13182);
nand U13673 (N_13673,N_12245,N_12213);
nor U13674 (N_13674,N_12822,N_12586);
xor U13675 (N_13675,N_12936,N_12965);
or U13676 (N_13676,N_12229,N_12126);
or U13677 (N_13677,N_12693,N_12151);
and U13678 (N_13678,N_12414,N_13065);
xnor U13679 (N_13679,N_12566,N_12684);
xnor U13680 (N_13680,N_12753,N_13160);
xnor U13681 (N_13681,N_12939,N_12500);
xor U13682 (N_13682,N_13139,N_13172);
nand U13683 (N_13683,N_12959,N_12687);
nor U13684 (N_13684,N_12933,N_12199);
nand U13685 (N_13685,N_12429,N_12521);
nor U13686 (N_13686,N_12438,N_12066);
nor U13687 (N_13687,N_12372,N_12661);
and U13688 (N_13688,N_13147,N_12076);
nand U13689 (N_13689,N_13064,N_12571);
xor U13690 (N_13690,N_12632,N_12464);
and U13691 (N_13691,N_12136,N_12893);
nand U13692 (N_13692,N_13107,N_12314);
nand U13693 (N_13693,N_12059,N_12572);
nand U13694 (N_13694,N_12353,N_12864);
or U13695 (N_13695,N_12906,N_12084);
and U13696 (N_13696,N_12366,N_12892);
nand U13697 (N_13697,N_12275,N_12685);
or U13698 (N_13698,N_12459,N_12064);
nand U13699 (N_13699,N_12937,N_12523);
xnor U13700 (N_13700,N_13138,N_12767);
nor U13701 (N_13701,N_12412,N_12913);
xor U13702 (N_13702,N_12371,N_13156);
or U13703 (N_13703,N_12071,N_12707);
xor U13704 (N_13704,N_12115,N_12771);
and U13705 (N_13705,N_12530,N_12188);
xnor U13706 (N_13706,N_12395,N_12701);
nand U13707 (N_13707,N_12258,N_12073);
nand U13708 (N_13708,N_12037,N_12648);
or U13709 (N_13709,N_13020,N_12671);
nor U13710 (N_13710,N_12270,N_13167);
nor U13711 (N_13711,N_12787,N_12117);
or U13712 (N_13712,N_12842,N_12935);
xor U13713 (N_13713,N_13007,N_12186);
nor U13714 (N_13714,N_13126,N_13092);
xnor U13715 (N_13715,N_12665,N_13029);
and U13716 (N_13716,N_12810,N_12549);
or U13717 (N_13717,N_12914,N_12243);
xor U13718 (N_13718,N_12244,N_12223);
nor U13719 (N_13719,N_12580,N_12697);
and U13720 (N_13720,N_12976,N_12926);
xnor U13721 (N_13721,N_12679,N_12351);
or U13722 (N_13722,N_12957,N_12211);
nor U13723 (N_13723,N_12178,N_12301);
or U13724 (N_13724,N_13115,N_12786);
nor U13725 (N_13725,N_12288,N_13134);
xor U13726 (N_13726,N_12680,N_12605);
nand U13727 (N_13727,N_12428,N_12617);
nand U13728 (N_13728,N_13013,N_12849);
or U13729 (N_13729,N_13049,N_12382);
xnor U13730 (N_13730,N_12969,N_12411);
nand U13731 (N_13731,N_12950,N_13187);
or U13732 (N_13732,N_13177,N_12373);
or U13733 (N_13733,N_12316,N_12646);
and U13734 (N_13734,N_12948,N_12198);
xnor U13735 (N_13735,N_12983,N_12520);
or U13736 (N_13736,N_12330,N_12890);
xnor U13737 (N_13737,N_12861,N_13081);
nand U13738 (N_13738,N_12903,N_12481);
nor U13739 (N_13739,N_12834,N_12584);
nand U13740 (N_13740,N_13034,N_12932);
nand U13741 (N_13741,N_12458,N_12525);
xor U13742 (N_13742,N_12106,N_12359);
nand U13743 (N_13743,N_12816,N_12103);
and U13744 (N_13744,N_12819,N_12604);
xnor U13745 (N_13745,N_12197,N_13176);
nand U13746 (N_13746,N_12249,N_12028);
or U13747 (N_13747,N_12074,N_12048);
or U13748 (N_13748,N_13012,N_12881);
nand U13749 (N_13749,N_12592,N_13192);
xor U13750 (N_13750,N_13089,N_13153);
nor U13751 (N_13751,N_12274,N_12506);
xor U13752 (N_13752,N_12432,N_13086);
and U13753 (N_13753,N_12120,N_12336);
or U13754 (N_13754,N_13052,N_12559);
and U13755 (N_13755,N_12909,N_12795);
xnor U13756 (N_13756,N_13000,N_12691);
nor U13757 (N_13757,N_12770,N_13071);
nand U13758 (N_13758,N_12689,N_12683);
xor U13759 (N_13759,N_12900,N_12814);
nor U13760 (N_13760,N_12526,N_12008);
nand U13761 (N_13761,N_13031,N_12762);
and U13762 (N_13762,N_13114,N_12515);
or U13763 (N_13763,N_12410,N_13180);
or U13764 (N_13764,N_12444,N_12159);
and U13765 (N_13765,N_12489,N_13069);
nor U13766 (N_13766,N_12660,N_12982);
or U13767 (N_13767,N_13015,N_12420);
xor U13768 (N_13768,N_12466,N_12550);
nand U13769 (N_13769,N_12086,N_12543);
nor U13770 (N_13770,N_12160,N_12879);
xnor U13771 (N_13771,N_12006,N_12885);
and U13772 (N_13772,N_12711,N_12163);
nand U13773 (N_13773,N_13003,N_13154);
nand U13774 (N_13774,N_12434,N_12798);
nor U13775 (N_13775,N_12467,N_12647);
nand U13776 (N_13776,N_12152,N_12504);
nand U13777 (N_13777,N_12941,N_12129);
nand U13778 (N_13778,N_12165,N_12319);
xnor U13779 (N_13779,N_12182,N_12121);
nor U13780 (N_13780,N_12544,N_12695);
nand U13781 (N_13781,N_12067,N_13074);
or U13782 (N_13782,N_12736,N_12290);
and U13783 (N_13783,N_12912,N_12501);
or U13784 (N_13784,N_12015,N_12183);
xnor U13785 (N_13785,N_12224,N_12146);
nand U13786 (N_13786,N_13039,N_12096);
nor U13787 (N_13787,N_12978,N_12153);
nand U13788 (N_13788,N_12240,N_12318);
and U13789 (N_13789,N_12949,N_12421);
and U13790 (N_13790,N_12091,N_12492);
and U13791 (N_13791,N_12634,N_12793);
nand U13792 (N_13792,N_13026,N_12863);
nand U13793 (N_13793,N_12269,N_12092);
nor U13794 (N_13794,N_12044,N_12659);
nor U13795 (N_13795,N_12727,N_12287);
or U13796 (N_13796,N_13009,N_13037);
xnor U13797 (N_13797,N_13146,N_13099);
xor U13798 (N_13798,N_12246,N_12817);
or U13799 (N_13799,N_13175,N_12512);
or U13800 (N_13800,N_12603,N_12497);
or U13801 (N_13801,N_12896,N_12952);
or U13802 (N_13802,N_12240,N_12859);
nor U13803 (N_13803,N_12999,N_12184);
and U13804 (N_13804,N_12721,N_13068);
xnor U13805 (N_13805,N_13189,N_12584);
and U13806 (N_13806,N_12901,N_13019);
xor U13807 (N_13807,N_12635,N_13184);
xor U13808 (N_13808,N_12487,N_12843);
nor U13809 (N_13809,N_12557,N_12738);
xor U13810 (N_13810,N_12210,N_13069);
xor U13811 (N_13811,N_13048,N_12480);
xor U13812 (N_13812,N_12037,N_13102);
nand U13813 (N_13813,N_12078,N_12976);
nor U13814 (N_13814,N_12872,N_12178);
or U13815 (N_13815,N_12790,N_12240);
or U13816 (N_13816,N_12366,N_12140);
nand U13817 (N_13817,N_12237,N_12857);
nand U13818 (N_13818,N_13005,N_12318);
or U13819 (N_13819,N_12444,N_12765);
or U13820 (N_13820,N_12827,N_12891);
and U13821 (N_13821,N_12732,N_13065);
nor U13822 (N_13822,N_12485,N_12158);
or U13823 (N_13823,N_12296,N_12982);
xnor U13824 (N_13824,N_12929,N_13022);
nor U13825 (N_13825,N_12638,N_12267);
nand U13826 (N_13826,N_13086,N_12800);
xor U13827 (N_13827,N_12280,N_12911);
or U13828 (N_13828,N_12485,N_12122);
nor U13829 (N_13829,N_13125,N_13185);
xor U13830 (N_13830,N_12899,N_12218);
xor U13831 (N_13831,N_12099,N_12467);
nor U13832 (N_13832,N_12092,N_12697);
and U13833 (N_13833,N_13146,N_12808);
nor U13834 (N_13834,N_12920,N_12968);
or U13835 (N_13835,N_12579,N_12562);
or U13836 (N_13836,N_12398,N_12561);
xor U13837 (N_13837,N_12160,N_12919);
and U13838 (N_13838,N_12930,N_13199);
xnor U13839 (N_13839,N_12004,N_12844);
and U13840 (N_13840,N_12539,N_12321);
and U13841 (N_13841,N_12161,N_12061);
nand U13842 (N_13842,N_12329,N_12081);
xor U13843 (N_13843,N_12048,N_12636);
xor U13844 (N_13844,N_12744,N_12797);
and U13845 (N_13845,N_12787,N_12180);
nor U13846 (N_13846,N_12570,N_13105);
nor U13847 (N_13847,N_12573,N_12394);
nor U13848 (N_13848,N_13164,N_12839);
nor U13849 (N_13849,N_12516,N_12509);
nand U13850 (N_13850,N_13002,N_12959);
or U13851 (N_13851,N_12423,N_12996);
or U13852 (N_13852,N_12100,N_12825);
nand U13853 (N_13853,N_12543,N_12516);
or U13854 (N_13854,N_12744,N_12149);
and U13855 (N_13855,N_13111,N_12128);
xor U13856 (N_13856,N_12154,N_12724);
and U13857 (N_13857,N_12117,N_13185);
nor U13858 (N_13858,N_12223,N_12369);
or U13859 (N_13859,N_13003,N_12705);
nand U13860 (N_13860,N_12397,N_12773);
and U13861 (N_13861,N_12558,N_12687);
xor U13862 (N_13862,N_12790,N_13069);
nor U13863 (N_13863,N_12831,N_12217);
xor U13864 (N_13864,N_12284,N_12214);
xor U13865 (N_13865,N_12260,N_13197);
nand U13866 (N_13866,N_12597,N_13186);
nor U13867 (N_13867,N_12297,N_13021);
nor U13868 (N_13868,N_12954,N_12116);
nor U13869 (N_13869,N_12014,N_12781);
and U13870 (N_13870,N_12880,N_12727);
nor U13871 (N_13871,N_13162,N_12393);
and U13872 (N_13872,N_12311,N_13176);
or U13873 (N_13873,N_13130,N_12833);
and U13874 (N_13874,N_12514,N_12544);
nor U13875 (N_13875,N_12924,N_12379);
nand U13876 (N_13876,N_13102,N_12858);
or U13877 (N_13877,N_12777,N_12304);
or U13878 (N_13878,N_12298,N_12810);
xor U13879 (N_13879,N_12785,N_12056);
nor U13880 (N_13880,N_12030,N_12846);
nand U13881 (N_13881,N_12427,N_13154);
nand U13882 (N_13882,N_13128,N_12846);
nor U13883 (N_13883,N_12821,N_12182);
and U13884 (N_13884,N_12329,N_12497);
or U13885 (N_13885,N_12876,N_12976);
and U13886 (N_13886,N_12265,N_12592);
and U13887 (N_13887,N_12878,N_12687);
nand U13888 (N_13888,N_12961,N_12201);
and U13889 (N_13889,N_13178,N_12597);
xnor U13890 (N_13890,N_12227,N_12188);
xor U13891 (N_13891,N_12570,N_12258);
or U13892 (N_13892,N_12407,N_12479);
or U13893 (N_13893,N_13195,N_13051);
xnor U13894 (N_13894,N_12884,N_12878);
xnor U13895 (N_13895,N_13027,N_12690);
or U13896 (N_13896,N_13148,N_12925);
or U13897 (N_13897,N_12658,N_12854);
nand U13898 (N_13898,N_12583,N_12429);
nor U13899 (N_13899,N_12043,N_12175);
nor U13900 (N_13900,N_13177,N_12727);
and U13901 (N_13901,N_13138,N_12214);
nand U13902 (N_13902,N_12692,N_12447);
nor U13903 (N_13903,N_12596,N_12296);
nor U13904 (N_13904,N_12327,N_12889);
nor U13905 (N_13905,N_12532,N_12002);
nor U13906 (N_13906,N_12914,N_12385);
xor U13907 (N_13907,N_12250,N_12121);
and U13908 (N_13908,N_12873,N_12744);
and U13909 (N_13909,N_12133,N_13031);
and U13910 (N_13910,N_12821,N_12025);
nor U13911 (N_13911,N_12248,N_12129);
nor U13912 (N_13912,N_12872,N_13068);
nand U13913 (N_13913,N_12826,N_12429);
and U13914 (N_13914,N_12518,N_12645);
and U13915 (N_13915,N_12934,N_12136);
or U13916 (N_13916,N_13111,N_12991);
xor U13917 (N_13917,N_12690,N_12862);
nor U13918 (N_13918,N_13186,N_13193);
xor U13919 (N_13919,N_12364,N_12739);
nor U13920 (N_13920,N_12259,N_12232);
or U13921 (N_13921,N_12053,N_12567);
xnor U13922 (N_13922,N_12344,N_12245);
and U13923 (N_13923,N_12681,N_12479);
and U13924 (N_13924,N_12222,N_13080);
nand U13925 (N_13925,N_13099,N_12114);
or U13926 (N_13926,N_12182,N_12581);
nor U13927 (N_13927,N_13141,N_12673);
nand U13928 (N_13928,N_13044,N_12578);
or U13929 (N_13929,N_12068,N_13066);
xor U13930 (N_13930,N_12698,N_12377);
xor U13931 (N_13931,N_12829,N_13001);
nand U13932 (N_13932,N_12636,N_12100);
and U13933 (N_13933,N_12870,N_12682);
or U13934 (N_13934,N_12058,N_12992);
or U13935 (N_13935,N_12736,N_13036);
nand U13936 (N_13936,N_12244,N_12397);
nand U13937 (N_13937,N_12790,N_12035);
nand U13938 (N_13938,N_12453,N_12822);
nor U13939 (N_13939,N_13095,N_12728);
nor U13940 (N_13940,N_12586,N_12326);
or U13941 (N_13941,N_13172,N_12394);
nor U13942 (N_13942,N_12528,N_12492);
or U13943 (N_13943,N_12019,N_12735);
nor U13944 (N_13944,N_13052,N_12779);
nand U13945 (N_13945,N_12357,N_12234);
nand U13946 (N_13946,N_12435,N_12664);
xnor U13947 (N_13947,N_12757,N_12588);
and U13948 (N_13948,N_13028,N_12888);
xor U13949 (N_13949,N_12769,N_12470);
and U13950 (N_13950,N_12791,N_12866);
and U13951 (N_13951,N_12320,N_12285);
nor U13952 (N_13952,N_12934,N_12697);
or U13953 (N_13953,N_13019,N_12847);
nor U13954 (N_13954,N_12009,N_12419);
xor U13955 (N_13955,N_12727,N_12494);
xor U13956 (N_13956,N_12730,N_12873);
nand U13957 (N_13957,N_12093,N_12345);
xor U13958 (N_13958,N_12677,N_12316);
or U13959 (N_13959,N_12964,N_12137);
xnor U13960 (N_13960,N_13034,N_12026);
and U13961 (N_13961,N_12881,N_12078);
or U13962 (N_13962,N_12555,N_12113);
xnor U13963 (N_13963,N_12577,N_12357);
and U13964 (N_13964,N_12330,N_12524);
and U13965 (N_13965,N_12123,N_12512);
nand U13966 (N_13966,N_12949,N_12263);
xor U13967 (N_13967,N_12800,N_12156);
or U13968 (N_13968,N_12293,N_12060);
nand U13969 (N_13969,N_12875,N_13082);
or U13970 (N_13970,N_12618,N_12721);
or U13971 (N_13971,N_12001,N_13108);
or U13972 (N_13972,N_12975,N_12062);
xor U13973 (N_13973,N_13110,N_12576);
or U13974 (N_13974,N_13028,N_12878);
or U13975 (N_13975,N_13063,N_13124);
nor U13976 (N_13976,N_12708,N_12777);
or U13977 (N_13977,N_12252,N_12216);
and U13978 (N_13978,N_12180,N_12009);
nor U13979 (N_13979,N_13084,N_12941);
xor U13980 (N_13980,N_12480,N_12677);
and U13981 (N_13981,N_12320,N_12785);
and U13982 (N_13982,N_12993,N_12238);
and U13983 (N_13983,N_12858,N_12468);
and U13984 (N_13984,N_13176,N_12155);
xor U13985 (N_13985,N_12184,N_12044);
nand U13986 (N_13986,N_12485,N_12410);
or U13987 (N_13987,N_12525,N_12481);
nand U13988 (N_13988,N_12244,N_12163);
nor U13989 (N_13989,N_12709,N_12901);
or U13990 (N_13990,N_13101,N_13149);
and U13991 (N_13991,N_12245,N_12888);
or U13992 (N_13992,N_12068,N_12496);
xnor U13993 (N_13993,N_13005,N_12336);
or U13994 (N_13994,N_12600,N_12536);
nand U13995 (N_13995,N_12146,N_13067);
xnor U13996 (N_13996,N_12677,N_12105);
xor U13997 (N_13997,N_12667,N_12124);
nor U13998 (N_13998,N_12674,N_12581);
or U13999 (N_13999,N_12569,N_12119);
and U14000 (N_14000,N_12577,N_12732);
or U14001 (N_14001,N_12710,N_12552);
nand U14002 (N_14002,N_12287,N_12148);
and U14003 (N_14003,N_12864,N_12306);
nand U14004 (N_14004,N_12633,N_12740);
nor U14005 (N_14005,N_12842,N_12086);
xor U14006 (N_14006,N_12904,N_13159);
nand U14007 (N_14007,N_13065,N_12633);
or U14008 (N_14008,N_13086,N_12576);
or U14009 (N_14009,N_13097,N_12850);
or U14010 (N_14010,N_12354,N_12479);
or U14011 (N_14011,N_12672,N_13109);
nor U14012 (N_14012,N_12626,N_12155);
xnor U14013 (N_14013,N_12880,N_12913);
and U14014 (N_14014,N_12754,N_12360);
xor U14015 (N_14015,N_12308,N_12416);
or U14016 (N_14016,N_13176,N_12614);
nand U14017 (N_14017,N_13103,N_12629);
or U14018 (N_14018,N_12754,N_12042);
or U14019 (N_14019,N_12314,N_13046);
nand U14020 (N_14020,N_12646,N_12131);
and U14021 (N_14021,N_13191,N_12273);
xnor U14022 (N_14022,N_12441,N_12803);
and U14023 (N_14023,N_12185,N_12269);
and U14024 (N_14024,N_12674,N_12183);
nor U14025 (N_14025,N_12158,N_12636);
or U14026 (N_14026,N_12752,N_12677);
nor U14027 (N_14027,N_12148,N_12689);
or U14028 (N_14028,N_13009,N_12748);
and U14029 (N_14029,N_12855,N_12463);
nand U14030 (N_14030,N_12389,N_12804);
and U14031 (N_14031,N_13092,N_12440);
nand U14032 (N_14032,N_12857,N_12448);
and U14033 (N_14033,N_13097,N_13018);
nor U14034 (N_14034,N_12307,N_12006);
nor U14035 (N_14035,N_12348,N_13069);
xor U14036 (N_14036,N_12293,N_12571);
nand U14037 (N_14037,N_12245,N_13060);
and U14038 (N_14038,N_12287,N_12517);
nor U14039 (N_14039,N_12064,N_13037);
xnor U14040 (N_14040,N_12950,N_12297);
and U14041 (N_14041,N_13154,N_13100);
nand U14042 (N_14042,N_12589,N_12389);
xnor U14043 (N_14043,N_12432,N_12299);
nand U14044 (N_14044,N_12539,N_12516);
xor U14045 (N_14045,N_12937,N_13172);
and U14046 (N_14046,N_12589,N_12931);
and U14047 (N_14047,N_12805,N_12986);
or U14048 (N_14048,N_12876,N_12915);
and U14049 (N_14049,N_13105,N_12528);
nor U14050 (N_14050,N_12887,N_12613);
nor U14051 (N_14051,N_13108,N_12906);
nor U14052 (N_14052,N_12692,N_12319);
nor U14053 (N_14053,N_12863,N_12952);
nand U14054 (N_14054,N_12328,N_12060);
nor U14055 (N_14055,N_12375,N_12659);
nand U14056 (N_14056,N_12750,N_12494);
and U14057 (N_14057,N_12662,N_12535);
or U14058 (N_14058,N_12547,N_12790);
or U14059 (N_14059,N_12286,N_12277);
nand U14060 (N_14060,N_12625,N_12428);
xnor U14061 (N_14061,N_13066,N_12989);
and U14062 (N_14062,N_12380,N_12284);
or U14063 (N_14063,N_12648,N_13173);
xor U14064 (N_14064,N_12921,N_12873);
or U14065 (N_14065,N_13107,N_13086);
or U14066 (N_14066,N_12337,N_12430);
nand U14067 (N_14067,N_12372,N_12510);
xnor U14068 (N_14068,N_12753,N_13143);
nand U14069 (N_14069,N_13168,N_12749);
or U14070 (N_14070,N_13152,N_13114);
xor U14071 (N_14071,N_12360,N_12111);
xnor U14072 (N_14072,N_12086,N_12644);
or U14073 (N_14073,N_12353,N_12038);
nor U14074 (N_14074,N_12425,N_12851);
nor U14075 (N_14075,N_13015,N_12861);
xor U14076 (N_14076,N_12337,N_12153);
nand U14077 (N_14077,N_12337,N_12323);
and U14078 (N_14078,N_12313,N_13027);
or U14079 (N_14079,N_12085,N_12889);
xor U14080 (N_14080,N_13068,N_12802);
and U14081 (N_14081,N_12118,N_13071);
or U14082 (N_14082,N_12185,N_12161);
nand U14083 (N_14083,N_12975,N_12633);
or U14084 (N_14084,N_12660,N_12430);
nor U14085 (N_14085,N_12080,N_12272);
and U14086 (N_14086,N_12400,N_12107);
or U14087 (N_14087,N_12674,N_12727);
or U14088 (N_14088,N_13109,N_12861);
xor U14089 (N_14089,N_12897,N_12680);
xnor U14090 (N_14090,N_12669,N_12126);
nand U14091 (N_14091,N_13122,N_12587);
nand U14092 (N_14092,N_12113,N_13025);
nand U14093 (N_14093,N_12939,N_12632);
xor U14094 (N_14094,N_12614,N_12903);
xnor U14095 (N_14095,N_13041,N_12331);
nand U14096 (N_14096,N_12289,N_12287);
nor U14097 (N_14097,N_12707,N_12300);
nand U14098 (N_14098,N_13046,N_12547);
nand U14099 (N_14099,N_12234,N_13056);
and U14100 (N_14100,N_12917,N_12307);
nand U14101 (N_14101,N_12154,N_12172);
nand U14102 (N_14102,N_12214,N_12938);
nor U14103 (N_14103,N_13076,N_12910);
nand U14104 (N_14104,N_13155,N_12901);
and U14105 (N_14105,N_12406,N_12547);
and U14106 (N_14106,N_12794,N_13084);
xnor U14107 (N_14107,N_13090,N_12713);
nand U14108 (N_14108,N_13096,N_12624);
nor U14109 (N_14109,N_12558,N_12236);
xor U14110 (N_14110,N_12410,N_12955);
nor U14111 (N_14111,N_12900,N_12343);
xnor U14112 (N_14112,N_12497,N_13111);
xnor U14113 (N_14113,N_13038,N_12153);
nand U14114 (N_14114,N_12405,N_12811);
nand U14115 (N_14115,N_12063,N_12632);
and U14116 (N_14116,N_12901,N_12745);
or U14117 (N_14117,N_12708,N_12924);
nor U14118 (N_14118,N_12091,N_12963);
xor U14119 (N_14119,N_12951,N_12557);
nand U14120 (N_14120,N_12342,N_13192);
nand U14121 (N_14121,N_12497,N_12297);
nor U14122 (N_14122,N_12833,N_12399);
xnor U14123 (N_14123,N_12354,N_12552);
or U14124 (N_14124,N_12108,N_12741);
nand U14125 (N_14125,N_12663,N_12076);
nand U14126 (N_14126,N_13007,N_12485);
or U14127 (N_14127,N_12126,N_12529);
xor U14128 (N_14128,N_12766,N_12369);
xnor U14129 (N_14129,N_12977,N_12798);
nor U14130 (N_14130,N_12162,N_12061);
nand U14131 (N_14131,N_12157,N_12804);
nand U14132 (N_14132,N_12415,N_13128);
nand U14133 (N_14133,N_12228,N_12491);
or U14134 (N_14134,N_12128,N_12026);
or U14135 (N_14135,N_12573,N_12832);
xor U14136 (N_14136,N_13001,N_12953);
xnor U14137 (N_14137,N_12319,N_12057);
or U14138 (N_14138,N_12431,N_12258);
nor U14139 (N_14139,N_12388,N_13095);
and U14140 (N_14140,N_13192,N_12858);
xnor U14141 (N_14141,N_12444,N_13121);
nor U14142 (N_14142,N_13097,N_12456);
and U14143 (N_14143,N_12082,N_12727);
nand U14144 (N_14144,N_12177,N_12897);
nor U14145 (N_14145,N_12782,N_12266);
xor U14146 (N_14146,N_12164,N_12004);
and U14147 (N_14147,N_12038,N_12446);
nor U14148 (N_14148,N_13033,N_12611);
nor U14149 (N_14149,N_12820,N_13085);
nor U14150 (N_14150,N_12640,N_12720);
or U14151 (N_14151,N_12659,N_12479);
xor U14152 (N_14152,N_12414,N_12563);
and U14153 (N_14153,N_13094,N_12109);
nand U14154 (N_14154,N_12087,N_12095);
nand U14155 (N_14155,N_12061,N_12952);
and U14156 (N_14156,N_12192,N_12121);
xor U14157 (N_14157,N_12377,N_12958);
nand U14158 (N_14158,N_12119,N_12513);
and U14159 (N_14159,N_12857,N_12568);
xnor U14160 (N_14160,N_12038,N_13010);
xnor U14161 (N_14161,N_12143,N_13094);
xor U14162 (N_14162,N_12191,N_12592);
or U14163 (N_14163,N_13017,N_12331);
or U14164 (N_14164,N_12825,N_13053);
or U14165 (N_14165,N_12991,N_12573);
and U14166 (N_14166,N_12795,N_12966);
xnor U14167 (N_14167,N_12789,N_12419);
nand U14168 (N_14168,N_12096,N_12971);
xnor U14169 (N_14169,N_12447,N_12449);
nor U14170 (N_14170,N_12222,N_13167);
or U14171 (N_14171,N_12712,N_12949);
and U14172 (N_14172,N_12580,N_12266);
or U14173 (N_14173,N_12606,N_12144);
and U14174 (N_14174,N_12883,N_13152);
xor U14175 (N_14175,N_12864,N_12392);
or U14176 (N_14176,N_12628,N_12071);
xor U14177 (N_14177,N_12455,N_12786);
and U14178 (N_14178,N_12121,N_12174);
and U14179 (N_14179,N_12985,N_13080);
nand U14180 (N_14180,N_12112,N_12839);
xor U14181 (N_14181,N_12024,N_13089);
and U14182 (N_14182,N_13149,N_12785);
nand U14183 (N_14183,N_12710,N_12848);
xor U14184 (N_14184,N_13173,N_12412);
or U14185 (N_14185,N_12287,N_13128);
xnor U14186 (N_14186,N_12765,N_12863);
nor U14187 (N_14187,N_12220,N_12743);
xor U14188 (N_14188,N_12757,N_13016);
xor U14189 (N_14189,N_12304,N_12411);
or U14190 (N_14190,N_12742,N_12911);
and U14191 (N_14191,N_13099,N_12621);
or U14192 (N_14192,N_12078,N_12483);
nand U14193 (N_14193,N_12507,N_12852);
and U14194 (N_14194,N_12976,N_12771);
nor U14195 (N_14195,N_12579,N_12542);
nand U14196 (N_14196,N_12422,N_12741);
and U14197 (N_14197,N_13168,N_12190);
xnor U14198 (N_14198,N_12673,N_12450);
nand U14199 (N_14199,N_12822,N_12889);
and U14200 (N_14200,N_12911,N_13105);
xnor U14201 (N_14201,N_12991,N_13116);
xor U14202 (N_14202,N_12788,N_12766);
nor U14203 (N_14203,N_12900,N_12898);
xnor U14204 (N_14204,N_13061,N_13081);
and U14205 (N_14205,N_12618,N_12947);
or U14206 (N_14206,N_12881,N_12641);
or U14207 (N_14207,N_12377,N_12261);
nand U14208 (N_14208,N_12451,N_13078);
nand U14209 (N_14209,N_12732,N_12874);
and U14210 (N_14210,N_12159,N_12465);
xnor U14211 (N_14211,N_12366,N_12786);
nand U14212 (N_14212,N_13010,N_12246);
nor U14213 (N_14213,N_12564,N_13145);
nor U14214 (N_14214,N_12425,N_12718);
nor U14215 (N_14215,N_12103,N_13014);
xnor U14216 (N_14216,N_12888,N_12289);
xnor U14217 (N_14217,N_12888,N_12775);
nand U14218 (N_14218,N_12288,N_12826);
nand U14219 (N_14219,N_13028,N_13114);
nand U14220 (N_14220,N_12245,N_12823);
xnor U14221 (N_14221,N_12002,N_12456);
nand U14222 (N_14222,N_13190,N_13111);
xnor U14223 (N_14223,N_13001,N_12409);
nor U14224 (N_14224,N_12461,N_12285);
and U14225 (N_14225,N_12358,N_12329);
nor U14226 (N_14226,N_12615,N_12601);
or U14227 (N_14227,N_12531,N_13024);
and U14228 (N_14228,N_12230,N_13008);
nand U14229 (N_14229,N_12604,N_12681);
and U14230 (N_14230,N_13065,N_12164);
and U14231 (N_14231,N_12626,N_12274);
nor U14232 (N_14232,N_12362,N_13118);
nor U14233 (N_14233,N_12528,N_12936);
and U14234 (N_14234,N_12334,N_12400);
nor U14235 (N_14235,N_12009,N_12919);
nand U14236 (N_14236,N_12723,N_12741);
and U14237 (N_14237,N_13147,N_12765);
or U14238 (N_14238,N_12321,N_12427);
or U14239 (N_14239,N_12380,N_12676);
nand U14240 (N_14240,N_13156,N_13162);
or U14241 (N_14241,N_12051,N_12856);
and U14242 (N_14242,N_12593,N_12363);
or U14243 (N_14243,N_12942,N_12897);
xnor U14244 (N_14244,N_12464,N_13030);
and U14245 (N_14245,N_12130,N_12735);
xor U14246 (N_14246,N_12750,N_13169);
or U14247 (N_14247,N_12817,N_12350);
xor U14248 (N_14248,N_12022,N_12487);
or U14249 (N_14249,N_12630,N_13135);
or U14250 (N_14250,N_13051,N_12951);
or U14251 (N_14251,N_12955,N_12209);
nand U14252 (N_14252,N_12851,N_12134);
nand U14253 (N_14253,N_12405,N_13157);
and U14254 (N_14254,N_12735,N_12637);
and U14255 (N_14255,N_12975,N_12193);
xor U14256 (N_14256,N_12763,N_12406);
nand U14257 (N_14257,N_13167,N_12384);
and U14258 (N_14258,N_12888,N_12619);
and U14259 (N_14259,N_12563,N_12903);
nand U14260 (N_14260,N_12756,N_12063);
nor U14261 (N_14261,N_12057,N_12571);
and U14262 (N_14262,N_12007,N_12965);
nand U14263 (N_14263,N_12079,N_12096);
nor U14264 (N_14264,N_12248,N_12661);
xor U14265 (N_14265,N_12741,N_13103);
nand U14266 (N_14266,N_12552,N_12342);
nor U14267 (N_14267,N_12652,N_12667);
nand U14268 (N_14268,N_12236,N_12179);
xor U14269 (N_14269,N_12234,N_13010);
and U14270 (N_14270,N_12822,N_12604);
nand U14271 (N_14271,N_12615,N_13054);
nand U14272 (N_14272,N_12373,N_12488);
nor U14273 (N_14273,N_12271,N_12191);
xnor U14274 (N_14274,N_12250,N_12596);
xor U14275 (N_14275,N_12460,N_12814);
and U14276 (N_14276,N_12525,N_12804);
and U14277 (N_14277,N_12014,N_12114);
and U14278 (N_14278,N_12978,N_12973);
xor U14279 (N_14279,N_12804,N_12620);
and U14280 (N_14280,N_12696,N_12598);
nor U14281 (N_14281,N_13010,N_12985);
nand U14282 (N_14282,N_12453,N_12167);
nand U14283 (N_14283,N_12434,N_12147);
xor U14284 (N_14284,N_12187,N_12288);
or U14285 (N_14285,N_12979,N_12670);
and U14286 (N_14286,N_12985,N_13190);
nand U14287 (N_14287,N_12184,N_12518);
nor U14288 (N_14288,N_12303,N_12359);
xor U14289 (N_14289,N_13173,N_12488);
and U14290 (N_14290,N_12644,N_12076);
xor U14291 (N_14291,N_12929,N_12047);
and U14292 (N_14292,N_13188,N_13095);
and U14293 (N_14293,N_12935,N_12548);
nor U14294 (N_14294,N_12367,N_12691);
xor U14295 (N_14295,N_13178,N_12119);
and U14296 (N_14296,N_12288,N_12255);
xor U14297 (N_14297,N_12505,N_12973);
xnor U14298 (N_14298,N_12064,N_12276);
and U14299 (N_14299,N_12514,N_12453);
nand U14300 (N_14300,N_12933,N_12116);
nand U14301 (N_14301,N_12555,N_12312);
and U14302 (N_14302,N_12829,N_13143);
nand U14303 (N_14303,N_13146,N_12753);
and U14304 (N_14304,N_12681,N_12520);
or U14305 (N_14305,N_12664,N_12883);
xor U14306 (N_14306,N_12993,N_12529);
and U14307 (N_14307,N_12127,N_12618);
nand U14308 (N_14308,N_12245,N_12431);
nand U14309 (N_14309,N_12260,N_12472);
nand U14310 (N_14310,N_12408,N_12522);
and U14311 (N_14311,N_12269,N_12113);
nand U14312 (N_14312,N_12965,N_12117);
nor U14313 (N_14313,N_12692,N_12079);
and U14314 (N_14314,N_13152,N_12412);
xor U14315 (N_14315,N_12987,N_12388);
xor U14316 (N_14316,N_12452,N_12066);
nand U14317 (N_14317,N_12462,N_13111);
xnor U14318 (N_14318,N_12461,N_13146);
or U14319 (N_14319,N_13041,N_12746);
nor U14320 (N_14320,N_12806,N_12745);
and U14321 (N_14321,N_12986,N_12772);
or U14322 (N_14322,N_12720,N_12971);
xor U14323 (N_14323,N_12130,N_13127);
xnor U14324 (N_14324,N_12397,N_12895);
or U14325 (N_14325,N_13028,N_12101);
nand U14326 (N_14326,N_12994,N_12442);
nor U14327 (N_14327,N_12330,N_12918);
and U14328 (N_14328,N_12376,N_12876);
or U14329 (N_14329,N_12571,N_12240);
or U14330 (N_14330,N_12004,N_12398);
and U14331 (N_14331,N_12861,N_12641);
xor U14332 (N_14332,N_12328,N_12024);
nor U14333 (N_14333,N_13197,N_13177);
or U14334 (N_14334,N_12624,N_12073);
nor U14335 (N_14335,N_12664,N_12780);
or U14336 (N_14336,N_13073,N_12882);
and U14337 (N_14337,N_12200,N_13021);
and U14338 (N_14338,N_12423,N_12070);
nand U14339 (N_14339,N_12213,N_12005);
and U14340 (N_14340,N_12459,N_13062);
xnor U14341 (N_14341,N_12071,N_12263);
xnor U14342 (N_14342,N_12359,N_12497);
xnor U14343 (N_14343,N_12230,N_12251);
nor U14344 (N_14344,N_12497,N_12554);
or U14345 (N_14345,N_12568,N_12190);
or U14346 (N_14346,N_12627,N_12949);
xor U14347 (N_14347,N_12864,N_12841);
nand U14348 (N_14348,N_12488,N_12872);
and U14349 (N_14349,N_12472,N_12774);
nand U14350 (N_14350,N_12424,N_12070);
nand U14351 (N_14351,N_12130,N_12056);
nor U14352 (N_14352,N_12904,N_13186);
or U14353 (N_14353,N_12291,N_12809);
xor U14354 (N_14354,N_12122,N_12731);
nor U14355 (N_14355,N_12686,N_12121);
nand U14356 (N_14356,N_12183,N_12220);
nor U14357 (N_14357,N_13078,N_13040);
nand U14358 (N_14358,N_12045,N_12674);
or U14359 (N_14359,N_12425,N_12389);
or U14360 (N_14360,N_12307,N_12202);
or U14361 (N_14361,N_12552,N_12156);
and U14362 (N_14362,N_12601,N_12113);
nand U14363 (N_14363,N_12973,N_12998);
xnor U14364 (N_14364,N_12608,N_12575);
and U14365 (N_14365,N_13018,N_13193);
nand U14366 (N_14366,N_12137,N_12601);
xnor U14367 (N_14367,N_13174,N_12895);
nor U14368 (N_14368,N_12253,N_12673);
or U14369 (N_14369,N_12033,N_12633);
or U14370 (N_14370,N_12709,N_13040);
nor U14371 (N_14371,N_12236,N_12056);
or U14372 (N_14372,N_13089,N_12857);
or U14373 (N_14373,N_13077,N_13194);
xnor U14374 (N_14374,N_12900,N_13194);
or U14375 (N_14375,N_12808,N_12265);
nor U14376 (N_14376,N_12346,N_12653);
or U14377 (N_14377,N_13176,N_12588);
xnor U14378 (N_14378,N_12828,N_12507);
nor U14379 (N_14379,N_12725,N_12802);
xor U14380 (N_14380,N_12522,N_13035);
and U14381 (N_14381,N_13023,N_12996);
or U14382 (N_14382,N_12202,N_12070);
nand U14383 (N_14383,N_12967,N_12979);
and U14384 (N_14384,N_12364,N_12303);
nor U14385 (N_14385,N_12531,N_13051);
nand U14386 (N_14386,N_12762,N_12790);
xnor U14387 (N_14387,N_12190,N_13029);
and U14388 (N_14388,N_12806,N_12828);
nor U14389 (N_14389,N_13148,N_12232);
nand U14390 (N_14390,N_12708,N_12660);
and U14391 (N_14391,N_12281,N_13009);
and U14392 (N_14392,N_12698,N_12792);
xor U14393 (N_14393,N_12331,N_12632);
nand U14394 (N_14394,N_12615,N_12932);
or U14395 (N_14395,N_12771,N_12721);
xnor U14396 (N_14396,N_12930,N_12054);
nand U14397 (N_14397,N_12778,N_13145);
nand U14398 (N_14398,N_13095,N_12653);
or U14399 (N_14399,N_12510,N_12527);
nand U14400 (N_14400,N_13322,N_13703);
or U14401 (N_14401,N_13873,N_13716);
or U14402 (N_14402,N_14071,N_13859);
nand U14403 (N_14403,N_13384,N_13405);
xor U14404 (N_14404,N_13363,N_13334);
nand U14405 (N_14405,N_13659,N_13840);
nor U14406 (N_14406,N_14107,N_14305);
or U14407 (N_14407,N_14054,N_14057);
xnor U14408 (N_14408,N_14256,N_13745);
or U14409 (N_14409,N_13688,N_13242);
nor U14410 (N_14410,N_13665,N_13442);
xnor U14411 (N_14411,N_14162,N_13743);
or U14412 (N_14412,N_14208,N_13722);
or U14413 (N_14413,N_14056,N_13781);
nand U14414 (N_14414,N_13890,N_13581);
nand U14415 (N_14415,N_13951,N_14258);
xor U14416 (N_14416,N_13562,N_14050);
nand U14417 (N_14417,N_13290,N_13664);
and U14418 (N_14418,N_13981,N_13495);
and U14419 (N_14419,N_14325,N_13741);
nor U14420 (N_14420,N_13862,N_13957);
and U14421 (N_14421,N_13652,N_13748);
nor U14422 (N_14422,N_13533,N_13358);
nand U14423 (N_14423,N_13385,N_13935);
or U14424 (N_14424,N_13387,N_13506);
and U14425 (N_14425,N_14275,N_13367);
xnor U14426 (N_14426,N_14194,N_13746);
and U14427 (N_14427,N_13552,N_14003);
nand U14428 (N_14428,N_13503,N_13401);
nand U14429 (N_14429,N_13956,N_13784);
and U14430 (N_14430,N_13393,N_14375);
nor U14431 (N_14431,N_14175,N_13885);
and U14432 (N_14432,N_13379,N_13430);
and U14433 (N_14433,N_14304,N_14318);
nand U14434 (N_14434,N_14079,N_14285);
nand U14435 (N_14435,N_13622,N_13501);
and U14436 (N_14436,N_14237,N_13252);
and U14437 (N_14437,N_13738,N_13250);
xor U14438 (N_14438,N_13273,N_14103);
xnor U14439 (N_14439,N_13233,N_13331);
or U14440 (N_14440,N_13473,N_14091);
or U14441 (N_14441,N_13778,N_13551);
and U14442 (N_14442,N_13677,N_14205);
and U14443 (N_14443,N_13436,N_14284);
xor U14444 (N_14444,N_13614,N_13757);
nand U14445 (N_14445,N_14131,N_13346);
or U14446 (N_14446,N_13596,N_13227);
nand U14447 (N_14447,N_13820,N_14130);
nor U14448 (N_14448,N_13921,N_13472);
nand U14449 (N_14449,N_13818,N_13924);
xnor U14450 (N_14450,N_13490,N_13431);
xor U14451 (N_14451,N_13355,N_13548);
or U14452 (N_14452,N_13940,N_13403);
nor U14453 (N_14453,N_13261,N_13296);
xor U14454 (N_14454,N_14055,N_13730);
and U14455 (N_14455,N_13587,N_14371);
or U14456 (N_14456,N_14243,N_13493);
nand U14457 (N_14457,N_14396,N_13416);
and U14458 (N_14458,N_13914,N_14180);
and U14459 (N_14459,N_13238,N_13550);
xor U14460 (N_14460,N_14366,N_14128);
or U14461 (N_14461,N_13723,N_13378);
or U14462 (N_14462,N_14352,N_14022);
nor U14463 (N_14463,N_13700,N_13661);
nand U14464 (N_14464,N_13631,N_14332);
xor U14465 (N_14465,N_14322,N_13452);
xor U14466 (N_14466,N_14141,N_13397);
and U14467 (N_14467,N_13790,N_14342);
nand U14468 (N_14468,N_13236,N_13314);
xnor U14469 (N_14469,N_14327,N_13636);
nor U14470 (N_14470,N_14093,N_13341);
nand U14471 (N_14471,N_13788,N_13642);
and U14472 (N_14472,N_14282,N_14347);
nor U14473 (N_14473,N_13698,N_13799);
xor U14474 (N_14474,N_13294,N_14334);
xnor U14475 (N_14475,N_13532,N_13374);
nor U14476 (N_14476,N_13860,N_13293);
nand U14477 (N_14477,N_14125,N_13417);
nand U14478 (N_14478,N_13595,N_13569);
nand U14479 (N_14479,N_13440,N_13360);
xor U14480 (N_14480,N_14169,N_14363);
xor U14481 (N_14481,N_13564,N_13215);
nor U14482 (N_14482,N_14254,N_14398);
and U14483 (N_14483,N_13832,N_13964);
and U14484 (N_14484,N_13710,N_13540);
and U14485 (N_14485,N_13909,N_14263);
or U14486 (N_14486,N_13444,N_13870);
nand U14487 (N_14487,N_14031,N_14348);
and U14488 (N_14488,N_13952,N_13549);
and U14489 (N_14489,N_13571,N_13381);
nand U14490 (N_14490,N_13750,N_14287);
xor U14491 (N_14491,N_14309,N_13663);
nor U14492 (N_14492,N_13866,N_13512);
and U14493 (N_14493,N_13680,N_14026);
nor U14494 (N_14494,N_13281,N_14227);
xor U14495 (N_14495,N_14321,N_14386);
nand U14496 (N_14496,N_14207,N_13829);
or U14497 (N_14497,N_14132,N_13310);
nor U14498 (N_14498,N_13773,N_13260);
or U14499 (N_14499,N_13879,N_13896);
nand U14500 (N_14500,N_13766,N_13625);
nor U14501 (N_14501,N_13299,N_14027);
nor U14502 (N_14502,N_13850,N_13447);
or U14503 (N_14503,N_14139,N_14383);
nand U14504 (N_14504,N_13612,N_13464);
xor U14505 (N_14505,N_14084,N_13992);
or U14506 (N_14506,N_14157,N_13649);
nor U14507 (N_14507,N_13209,N_13609);
nor U14508 (N_14508,N_13303,N_13971);
and U14509 (N_14509,N_13983,N_13232);
xor U14510 (N_14510,N_14115,N_14226);
and U14511 (N_14511,N_13574,N_13368);
nor U14512 (N_14512,N_13454,N_14061);
or U14513 (N_14513,N_13423,N_14264);
and U14514 (N_14514,N_13500,N_14025);
nand U14515 (N_14515,N_13205,N_13793);
and U14516 (N_14516,N_14124,N_13791);
and U14517 (N_14517,N_13223,N_14239);
nand U14518 (N_14518,N_13254,N_14001);
xor U14519 (N_14519,N_14283,N_13289);
xor U14520 (N_14520,N_13409,N_14369);
or U14521 (N_14521,N_13613,N_14095);
nand U14522 (N_14522,N_13295,N_13523);
and U14523 (N_14523,N_13491,N_13611);
nor U14524 (N_14524,N_13646,N_13243);
or U14525 (N_14525,N_14265,N_13984);
nor U14526 (N_14526,N_13208,N_13210);
nor U14527 (N_14527,N_14122,N_13561);
nor U14528 (N_14528,N_13797,N_14006);
nor U14529 (N_14529,N_13449,N_13993);
nor U14530 (N_14530,N_14087,N_14041);
and U14531 (N_14531,N_13725,N_13734);
or U14532 (N_14532,N_13383,N_14021);
xnor U14533 (N_14533,N_14364,N_14219);
xor U14534 (N_14534,N_13212,N_14242);
nor U14535 (N_14535,N_14296,N_13882);
xor U14536 (N_14536,N_13841,N_14066);
xor U14537 (N_14537,N_14229,N_14181);
xor U14538 (N_14538,N_14308,N_14004);
or U14539 (N_14539,N_13911,N_14178);
xor U14540 (N_14540,N_14261,N_13390);
xnor U14541 (N_14541,N_14397,N_14295);
or U14542 (N_14542,N_13932,N_13942);
xor U14543 (N_14543,N_13576,N_14344);
or U14544 (N_14544,N_13937,N_13831);
xor U14545 (N_14545,N_14209,N_14238);
xor U14546 (N_14546,N_13415,N_14297);
and U14547 (N_14547,N_14250,N_13749);
or U14548 (N_14548,N_14023,N_13699);
nor U14549 (N_14549,N_13286,N_14196);
xnor U14550 (N_14550,N_13967,N_13817);
nor U14551 (N_14551,N_14213,N_14349);
or U14552 (N_14552,N_14138,N_13535);
xor U14553 (N_14553,N_13708,N_13328);
nand U14554 (N_14554,N_14099,N_14255);
or U14555 (N_14555,N_13938,N_13715);
and U14556 (N_14556,N_14036,N_14279);
nor U14557 (N_14557,N_14030,N_14392);
nand U14558 (N_14558,N_13230,N_13207);
xnor U14559 (N_14559,N_13467,N_13991);
and U14560 (N_14560,N_14202,N_13568);
or U14561 (N_14561,N_13916,N_13779);
xnor U14562 (N_14562,N_14088,N_14268);
nor U14563 (N_14563,N_13451,N_13352);
xnor U14564 (N_14564,N_14230,N_14152);
or U14565 (N_14565,N_13408,N_14247);
xnor U14566 (N_14566,N_14108,N_14257);
xnor U14567 (N_14567,N_13627,N_13446);
or U14568 (N_14568,N_13908,N_14038);
or U14569 (N_14569,N_14126,N_13327);
xnor U14570 (N_14570,N_13843,N_13727);
or U14571 (N_14571,N_13350,N_14120);
nor U14572 (N_14572,N_14101,N_13563);
nand U14573 (N_14573,N_13827,N_14035);
and U14574 (N_14574,N_13789,N_13978);
xnor U14575 (N_14575,N_13284,N_13979);
nand U14576 (N_14576,N_13755,N_13487);
or U14577 (N_14577,N_14168,N_13498);
xor U14578 (N_14578,N_14359,N_13593);
or U14579 (N_14579,N_13849,N_13691);
or U14580 (N_14580,N_13411,N_13369);
and U14581 (N_14581,N_14290,N_14039);
or U14582 (N_14582,N_13783,N_13754);
or U14583 (N_14583,N_13272,N_13504);
and U14584 (N_14584,N_14377,N_13376);
or U14585 (N_14585,N_13221,N_13298);
nand U14586 (N_14586,N_13229,N_14320);
nand U14587 (N_14587,N_13982,N_13580);
xnor U14588 (N_14588,N_13427,N_13453);
and U14589 (N_14589,N_13675,N_13329);
nor U14590 (N_14590,N_14184,N_14102);
xnor U14591 (N_14591,N_14249,N_13584);
or U14592 (N_14592,N_13271,N_13657);
or U14593 (N_14593,N_14024,N_14358);
xnor U14594 (N_14594,N_14323,N_13724);
and U14595 (N_14595,N_14159,N_13960);
nand U14596 (N_14596,N_14011,N_13886);
xor U14597 (N_14597,N_13629,N_13884);
and U14598 (N_14598,N_13736,N_14013);
and U14599 (N_14599,N_13705,N_14060);
or U14600 (N_14600,N_14228,N_14374);
or U14601 (N_14601,N_13528,N_14073);
nor U14602 (N_14602,N_13547,N_13998);
and U14603 (N_14603,N_13201,N_13674);
nor U14604 (N_14604,N_13421,N_13573);
xor U14605 (N_14605,N_13362,N_14133);
nor U14606 (N_14606,N_13570,N_13428);
xnor U14607 (N_14607,N_13204,N_13412);
xor U14608 (N_14608,N_13466,N_13902);
nor U14609 (N_14609,N_13438,N_13963);
nand U14610 (N_14610,N_14203,N_13483);
nand U14611 (N_14611,N_13666,N_13263);
and U14612 (N_14612,N_13933,N_14121);
xor U14613 (N_14613,N_14075,N_13520);
nor U14614 (N_14614,N_13751,N_13333);
xnor U14615 (N_14615,N_14373,N_13364);
xor U14616 (N_14616,N_14140,N_13539);
nor U14617 (N_14617,N_13976,N_13828);
and U14618 (N_14618,N_13413,N_13988);
nor U14619 (N_14619,N_13740,N_13434);
and U14620 (N_14620,N_13653,N_14210);
or U14621 (N_14621,N_14136,N_13541);
xnor U14622 (N_14622,N_13669,N_14259);
xnor U14623 (N_14623,N_13557,N_13747);
xnor U14624 (N_14624,N_13950,N_13822);
nand U14625 (N_14625,N_13258,N_13835);
or U14626 (N_14626,N_13245,N_14063);
nand U14627 (N_14627,N_13765,N_14135);
xnor U14628 (N_14628,N_14146,N_14372);
nor U14629 (N_14629,N_13425,N_13887);
or U14630 (N_14630,N_13923,N_14389);
xor U14631 (N_14631,N_14393,N_14100);
and U14632 (N_14632,N_13519,N_13662);
nand U14633 (N_14633,N_14390,N_13899);
xor U14634 (N_14634,N_14316,N_14082);
or U14635 (N_14635,N_13762,N_14008);
nand U14636 (N_14636,N_13894,N_14232);
xor U14637 (N_14637,N_14292,N_13851);
and U14638 (N_14638,N_14160,N_13521);
nor U14639 (N_14639,N_13711,N_13544);
nor U14640 (N_14640,N_13819,N_13465);
nor U14641 (N_14641,N_13259,N_13913);
xor U14642 (N_14642,N_14089,N_13673);
and U14643 (N_14643,N_13795,N_13306);
or U14644 (N_14644,N_14299,N_13977);
xnor U14645 (N_14645,N_13257,N_14007);
nor U14646 (N_14646,N_13514,N_14064);
or U14647 (N_14647,N_14074,N_14300);
or U14648 (N_14648,N_13277,N_13463);
and U14649 (N_14649,N_13235,N_14340);
and U14650 (N_14650,N_14116,N_14307);
nand U14651 (N_14651,N_13304,N_13696);
xor U14652 (N_14652,N_14215,N_13955);
and U14653 (N_14653,N_13986,N_13315);
or U14654 (N_14654,N_13577,N_14154);
or U14655 (N_14655,N_14161,N_13839);
nand U14656 (N_14656,N_13966,N_13927);
or U14657 (N_14657,N_13482,N_14354);
nor U14658 (N_14658,N_13508,N_13947);
nand U14659 (N_14659,N_14391,N_13803);
or U14660 (N_14660,N_14179,N_14083);
xnor U14661 (N_14661,N_13837,N_13224);
nand U14662 (N_14662,N_14018,N_14142);
xor U14663 (N_14663,N_13634,N_13536);
and U14664 (N_14664,N_13400,N_13905);
or U14665 (N_14665,N_13255,N_13780);
or U14666 (N_14666,N_13985,N_14248);
nand U14667 (N_14667,N_13513,N_13624);
xor U14668 (N_14668,N_13392,N_13640);
and U14669 (N_14669,N_13953,N_14144);
nand U14670 (N_14670,N_13356,N_13647);
nor U14671 (N_14671,N_13763,N_13206);
and U14672 (N_14672,N_13237,N_13599);
or U14673 (N_14673,N_13437,N_13728);
nand U14674 (N_14674,N_13336,N_14173);
and U14675 (N_14675,N_14269,N_13433);
or U14676 (N_14676,N_13217,N_13450);
xor U14677 (N_14677,N_14153,N_14097);
nand U14678 (N_14678,N_13502,N_13214);
xor U14679 (N_14679,N_14233,N_13489);
nor U14680 (N_14680,N_13670,N_13878);
nand U14681 (N_14681,N_13658,N_14385);
nand U14682 (N_14682,N_13844,N_13726);
or U14683 (N_14683,N_13585,N_13335);
nand U14684 (N_14684,N_14311,N_13949);
and U14685 (N_14685,N_13382,N_14294);
or U14686 (N_14686,N_13994,N_13704);
and U14687 (N_14687,N_13359,N_13231);
nor U14688 (N_14688,N_13525,N_13494);
and U14689 (N_14689,N_14186,N_13815);
or U14690 (N_14690,N_13266,N_14266);
nand U14691 (N_14691,N_14353,N_14096);
and U14692 (N_14692,N_14176,N_13868);
xnor U14693 (N_14693,N_13709,N_14197);
and U14694 (N_14694,N_14267,N_13280);
or U14695 (N_14695,N_13898,N_13616);
xor U14696 (N_14696,N_13317,N_14034);
nor U14697 (N_14697,N_13347,N_14351);
and U14698 (N_14698,N_13800,N_13895);
nand U14699 (N_14699,N_13269,N_13848);
xnor U14700 (N_14700,N_13782,N_13537);
nand U14701 (N_14701,N_14337,N_13468);
xor U14702 (N_14702,N_13975,N_13253);
and U14703 (N_14703,N_13756,N_14231);
and U14704 (N_14704,N_14094,N_14235);
and U14705 (N_14705,N_13394,N_13968);
nor U14706 (N_14706,N_13961,N_14164);
or U14707 (N_14707,N_13618,N_13842);
and U14708 (N_14708,N_14360,N_14378);
xor U14709 (N_14709,N_13262,N_14183);
and U14710 (N_14710,N_13786,N_13742);
or U14711 (N_14711,N_13458,N_13319);
and U14712 (N_14712,N_13655,N_13845);
xor U14713 (N_14713,N_13684,N_13915);
nor U14714 (N_14714,N_13854,N_13804);
nor U14715 (N_14715,N_14170,N_13694);
nand U14716 (N_14716,N_13770,N_13241);
or U14717 (N_14717,N_13930,N_13302);
or U14718 (N_14718,N_13869,N_13311);
nand U14719 (N_14719,N_13488,N_13518);
xnor U14720 (N_14720,N_13889,N_13461);
nand U14721 (N_14721,N_14293,N_14067);
xnor U14722 (N_14722,N_13861,N_14106);
nand U14723 (N_14723,N_13922,N_14271);
or U14724 (N_14724,N_13496,N_14379);
nor U14725 (N_14725,N_14165,N_13247);
or U14726 (N_14726,N_13228,N_14313);
or U14727 (N_14727,N_14199,N_14076);
nor U14728 (N_14728,N_13633,N_14058);
nand U14729 (N_14729,N_14105,N_13478);
nand U14730 (N_14730,N_13660,N_13601);
and U14731 (N_14731,N_13510,N_13265);
or U14732 (N_14732,N_14047,N_13946);
nor U14733 (N_14733,N_13735,N_13492);
xnor U14734 (N_14734,N_14345,N_14338);
nand U14735 (N_14735,N_13396,N_14328);
or U14736 (N_14736,N_13338,N_13973);
or U14737 (N_14737,N_13893,N_13285);
and U14738 (N_14738,N_13202,N_13648);
xnor U14739 (N_14739,N_13366,N_13919);
nor U14740 (N_14740,N_13389,N_13481);
nand U14741 (N_14741,N_13610,N_14218);
xor U14742 (N_14742,N_13220,N_14346);
nor U14743 (N_14743,N_14356,N_14037);
nor U14744 (N_14744,N_13406,N_14220);
and U14745 (N_14745,N_13402,N_13522);
and U14746 (N_14746,N_13455,N_13853);
and U14747 (N_14747,N_13460,N_14053);
nor U14748 (N_14748,N_13941,N_13516);
nand U14749 (N_14749,N_13268,N_13559);
and U14750 (N_14750,N_14070,N_14043);
and U14751 (N_14751,N_14129,N_13486);
xnor U14752 (N_14752,N_14380,N_13872);
nor U14753 (N_14753,N_13958,N_13582);
nor U14754 (N_14754,N_13326,N_14240);
or U14755 (N_14755,N_13226,N_13744);
nand U14756 (N_14756,N_13639,N_13897);
or U14757 (N_14757,N_13880,N_13792);
nor U14758 (N_14758,N_13365,N_13904);
and U14759 (N_14759,N_14333,N_13701);
nor U14760 (N_14760,N_14381,N_13693);
and U14761 (N_14761,N_13772,N_13903);
and U14762 (N_14762,N_13240,N_13234);
nor U14763 (N_14763,N_13404,N_13211);
nor U14764 (N_14764,N_13632,N_14062);
and U14765 (N_14765,N_14357,N_13305);
nor U14766 (N_14766,N_13753,N_13989);
xnor U14767 (N_14767,N_13323,N_14010);
and U14768 (N_14768,N_14000,N_13321);
nor U14769 (N_14769,N_13638,N_13987);
or U14770 (N_14770,N_14111,N_13641);
and U14771 (N_14771,N_13300,N_13813);
and U14772 (N_14772,N_14110,N_13682);
nor U14773 (N_14773,N_14362,N_13928);
or U14774 (N_14774,N_13307,N_13370);
nand U14775 (N_14775,N_14005,N_13288);
xor U14776 (N_14776,N_14150,N_13920);
or U14777 (N_14777,N_13325,N_13477);
or U14778 (N_14778,N_13507,N_13324);
and U14779 (N_14779,N_13777,N_13714);
or U14780 (N_14780,N_14312,N_13667);
nand U14781 (N_14781,N_13429,N_13419);
nand U14782 (N_14782,N_13801,N_13936);
or U14783 (N_14783,N_14090,N_13871);
and U14784 (N_14784,N_13681,N_13420);
nor U14785 (N_14785,N_13598,N_13787);
or U14786 (N_14786,N_13316,N_13597);
nor U14787 (N_14787,N_13826,N_13200);
nor U14788 (N_14788,N_13720,N_14336);
xor U14789 (N_14789,N_13686,N_14216);
or U14790 (N_14790,N_14361,N_13697);
nand U14791 (N_14791,N_13424,N_13678);
nor U14792 (N_14792,N_13388,N_13256);
xnor U14793 (N_14793,N_13558,N_14331);
nand U14794 (N_14794,N_13555,N_14014);
and U14795 (N_14795,N_13717,N_13560);
xnor U14796 (N_14796,N_14195,N_14319);
nor U14797 (N_14797,N_13808,N_13538);
and U14798 (N_14798,N_13375,N_14212);
or U14799 (N_14799,N_13972,N_14065);
xnor U14800 (N_14800,N_13974,N_13441);
or U14801 (N_14801,N_14303,N_13471);
nor U14802 (N_14802,N_14270,N_13320);
nor U14803 (N_14803,N_14167,N_13283);
xor U14804 (N_14804,N_13497,N_13764);
nor U14805 (N_14805,N_13604,N_14281);
xnor U14806 (N_14806,N_13888,N_14211);
nand U14807 (N_14807,N_14187,N_14280);
and U14808 (N_14808,N_13630,N_14382);
or U14809 (N_14809,N_13891,N_13739);
and U14810 (N_14810,N_13264,N_13470);
xor U14811 (N_14811,N_13225,N_13836);
xor U14812 (N_14812,N_14191,N_14200);
nor U14813 (N_14813,N_13578,N_13776);
nand U14814 (N_14814,N_13918,N_13857);
and U14815 (N_14815,N_13353,N_13509);
or U14816 (N_14816,N_13203,N_14092);
or U14817 (N_14817,N_14326,N_14365);
and U14818 (N_14818,N_13798,N_14044);
nor U14819 (N_14819,N_13810,N_13399);
nor U14820 (N_14820,N_13858,N_13343);
and U14821 (N_14821,N_13372,N_14012);
xnor U14822 (N_14822,N_13589,N_13556);
nor U14823 (N_14823,N_13485,N_13856);
xnor U14824 (N_14824,N_13505,N_13594);
nand U14825 (N_14825,N_13959,N_13719);
and U14826 (N_14826,N_13695,N_13806);
or U14827 (N_14827,N_14277,N_14193);
and U14828 (N_14828,N_14223,N_13617);
nor U14829 (N_14829,N_13876,N_13469);
or U14830 (N_14830,N_13534,N_13809);
and U14831 (N_14831,N_14182,N_13654);
nand U14832 (N_14832,N_13929,N_13309);
nor U14833 (N_14833,N_13476,N_13917);
nand U14834 (N_14834,N_13925,N_13877);
or U14835 (N_14835,N_14376,N_13934);
or U14836 (N_14836,N_13308,N_13246);
nand U14837 (N_14837,N_13291,N_13279);
nor U14838 (N_14838,N_14246,N_14158);
or U14839 (N_14839,N_13566,N_14251);
nor U14840 (N_14840,N_13459,N_13270);
and U14841 (N_14841,N_14245,N_13901);
nand U14842 (N_14842,N_13759,N_13685);
nand U14843 (N_14843,N_14081,N_13637);
and U14844 (N_14844,N_13635,N_14028);
nor U14845 (N_14845,N_13676,N_14190);
nand U14846 (N_14846,N_14069,N_13999);
nand U14847 (N_14847,N_13931,N_14272);
nor U14848 (N_14848,N_13668,N_13216);
and U14849 (N_14849,N_13511,N_14214);
xnor U14850 (N_14850,N_14156,N_13865);
or U14851 (N_14851,N_14049,N_14368);
nand U14852 (N_14852,N_14278,N_14206);
nand U14853 (N_14853,N_13690,N_14324);
xor U14854 (N_14854,N_13621,N_13432);
nand U14855 (N_14855,N_13768,N_13683);
xnor U14856 (N_14856,N_14262,N_14098);
nand U14857 (N_14857,N_14341,N_14387);
nand U14858 (N_14858,N_14350,N_13970);
nand U14859 (N_14859,N_13371,N_14244);
xnor U14860 (N_14860,N_13332,N_14123);
nor U14861 (N_14861,N_13962,N_13480);
nor U14862 (N_14862,N_14330,N_13349);
nor U14863 (N_14863,N_13475,N_13954);
or U14864 (N_14864,N_14046,N_13457);
and U14865 (N_14865,N_14172,N_13628);
nor U14866 (N_14866,N_13603,N_13591);
or U14867 (N_14867,N_14163,N_13218);
or U14868 (N_14868,N_13834,N_13758);
and U14869 (N_14869,N_14253,N_13774);
xor U14870 (N_14870,N_13251,N_14306);
nor U14871 (N_14871,N_13456,N_13287);
and U14872 (N_14872,N_14201,N_14052);
and U14873 (N_14873,N_13386,N_13846);
nand U14874 (N_14874,N_13418,N_14029);
nor U14875 (N_14875,N_14204,N_13679);
xnor U14876 (N_14876,N_13656,N_14104);
nand U14877 (N_14877,N_13912,N_14384);
or U14878 (N_14878,N_13615,N_14335);
xnor U14879 (N_14879,N_14339,N_13892);
nand U14880 (N_14880,N_14015,N_13448);
or U14881 (N_14881,N_13769,N_13462);
and U14882 (N_14882,N_14317,N_14395);
or U14883 (N_14883,N_13439,N_14171);
and U14884 (N_14884,N_13301,N_13718);
nor U14885 (N_14885,N_13345,N_13811);
nor U14886 (N_14886,N_14032,N_13414);
or U14887 (N_14887,N_13608,N_13706);
nor U14888 (N_14888,N_13543,N_13565);
or U14889 (N_14889,N_14217,N_13545);
or U14890 (N_14890,N_13731,N_13297);
xnor U14891 (N_14891,N_14236,N_13244);
nor U14892 (N_14892,N_14177,N_13292);
xor U14893 (N_14893,N_14343,N_13278);
xor U14894 (N_14894,N_13713,N_14188);
and U14895 (N_14895,N_14399,N_13771);
nand U14896 (N_14896,N_14148,N_13883);
xor U14897 (N_14897,N_13602,N_13361);
xnor U14898 (N_14898,N_13814,N_13761);
xnor U14899 (N_14899,N_14147,N_13542);
nand U14900 (N_14900,N_13881,N_13380);
nand U14901 (N_14901,N_14260,N_13732);
or U14902 (N_14902,N_14117,N_13590);
or U14903 (N_14903,N_13249,N_14045);
xnor U14904 (N_14904,N_14388,N_13337);
and U14905 (N_14905,N_14080,N_14134);
nor U14906 (N_14906,N_13276,N_13479);
nor U14907 (N_14907,N_14040,N_13965);
or U14908 (N_14908,N_13515,N_13651);
nand U14909 (N_14909,N_13443,N_14314);
or U14910 (N_14910,N_13980,N_13499);
nand U14911 (N_14911,N_13526,N_13996);
nand U14912 (N_14912,N_14192,N_14143);
and U14913 (N_14913,N_13474,N_13377);
nor U14914 (N_14914,N_14166,N_13592);
xor U14915 (N_14915,N_14020,N_14051);
xnor U14916 (N_14916,N_13530,N_13864);
nand U14917 (N_14917,N_13671,N_13838);
nor U14918 (N_14918,N_13373,N_14291);
and U14919 (N_14919,N_13275,N_14042);
or U14920 (N_14920,N_14252,N_13990);
and U14921 (N_14921,N_14222,N_13619);
nand U14922 (N_14922,N_13531,N_13926);
or U14923 (N_14923,N_14033,N_13821);
nand U14924 (N_14924,N_13906,N_13948);
and U14925 (N_14925,N_13623,N_13867);
nor U14926 (N_14926,N_14198,N_14224);
xnor U14927 (N_14927,N_13944,N_13847);
nand U14928 (N_14928,N_13529,N_13852);
or U14929 (N_14929,N_14301,N_13407);
and U14930 (N_14930,N_14276,N_13620);
and U14931 (N_14931,N_13702,N_13344);
or U14932 (N_14932,N_13796,N_14085);
nor U14933 (N_14933,N_14370,N_13391);
nor U14934 (N_14934,N_13330,N_14394);
xnor U14935 (N_14935,N_13775,N_14113);
nand U14936 (N_14936,N_13833,N_14310);
and U14937 (N_14937,N_13579,N_13945);
nor U14938 (N_14938,N_14174,N_13767);
or U14939 (N_14939,N_13339,N_14329);
and U14940 (N_14940,N_13583,N_13398);
or U14941 (N_14941,N_13410,N_13554);
nand U14942 (N_14942,N_13274,N_13435);
and U14943 (N_14943,N_14112,N_13907);
xor U14944 (N_14944,N_13553,N_13312);
and U14945 (N_14945,N_13318,N_13605);
nand U14946 (N_14946,N_13282,N_13712);
nand U14947 (N_14947,N_13863,N_14048);
or U14948 (N_14948,N_13997,N_13874);
and U14949 (N_14949,N_13752,N_13348);
nor U14950 (N_14950,N_13760,N_13943);
nand U14951 (N_14951,N_13626,N_13484);
nand U14952 (N_14952,N_13572,N_13567);
and U14953 (N_14953,N_14086,N_13527);
nor U14954 (N_14954,N_13606,N_14185);
or U14955 (N_14955,N_13785,N_13969);
and U14956 (N_14956,N_13995,N_13340);
nor U14957 (N_14957,N_14302,N_13351);
or U14958 (N_14958,N_13875,N_13692);
nand U14959 (N_14959,N_14002,N_14355);
nor U14960 (N_14960,N_13600,N_14119);
and U14961 (N_14961,N_13707,N_13357);
and U14962 (N_14962,N_14149,N_13650);
nor U14963 (N_14963,N_13687,N_14155);
xnor U14964 (N_14964,N_13729,N_13689);
nand U14965 (N_14965,N_13825,N_13395);
nand U14966 (N_14966,N_14241,N_13248);
xor U14967 (N_14967,N_13816,N_14114);
nand U14968 (N_14968,N_14274,N_13645);
nand U14969 (N_14969,N_13213,N_13733);
or U14970 (N_14970,N_14286,N_13586);
xnor U14971 (N_14971,N_13855,N_13672);
nor U14972 (N_14972,N_13823,N_14077);
and U14973 (N_14973,N_13643,N_13313);
nand U14974 (N_14974,N_13422,N_13239);
xor U14975 (N_14975,N_14118,N_14109);
nand U14976 (N_14976,N_14145,N_13219);
nor U14977 (N_14977,N_14017,N_14019);
nand U14978 (N_14978,N_13222,N_14315);
nor U14979 (N_14979,N_13267,N_13575);
and U14980 (N_14980,N_13737,N_13546);
nor U14981 (N_14981,N_14273,N_14225);
xnor U14982 (N_14982,N_13342,N_14189);
or U14983 (N_14983,N_14016,N_14221);
nor U14984 (N_14984,N_14298,N_13910);
or U14985 (N_14985,N_13588,N_14137);
and U14986 (N_14986,N_13721,N_14288);
or U14987 (N_14987,N_14289,N_13354);
nand U14988 (N_14988,N_14367,N_14059);
and U14989 (N_14989,N_13426,N_13607);
nand U14990 (N_14990,N_13805,N_13812);
nor U14991 (N_14991,N_13807,N_14127);
nor U14992 (N_14992,N_13794,N_14009);
and U14993 (N_14993,N_14151,N_14078);
nand U14994 (N_14994,N_13802,N_13939);
nor U14995 (N_14995,N_13824,N_13900);
nand U14996 (N_14996,N_14234,N_14068);
nor U14997 (N_14997,N_14072,N_13830);
and U14998 (N_14998,N_13445,N_13644);
nand U14999 (N_14999,N_13524,N_13517);
nand U15000 (N_15000,N_13940,N_13778);
and U15001 (N_15001,N_13890,N_13355);
and U15002 (N_15002,N_13792,N_13383);
xnor U15003 (N_15003,N_13647,N_13532);
nand U15004 (N_15004,N_13518,N_13879);
nand U15005 (N_15005,N_13772,N_13202);
xnor U15006 (N_15006,N_13664,N_14096);
and U15007 (N_15007,N_14248,N_13390);
xnor U15008 (N_15008,N_14328,N_14234);
nand U15009 (N_15009,N_13964,N_13825);
and U15010 (N_15010,N_14318,N_13997);
and U15011 (N_15011,N_14371,N_13898);
or U15012 (N_15012,N_13410,N_13466);
or U15013 (N_15013,N_14038,N_13582);
or U15014 (N_15014,N_13496,N_13435);
xnor U15015 (N_15015,N_13444,N_13804);
nand U15016 (N_15016,N_14363,N_13710);
nand U15017 (N_15017,N_14134,N_13915);
or U15018 (N_15018,N_14334,N_13928);
or U15019 (N_15019,N_13506,N_13942);
and U15020 (N_15020,N_13635,N_13748);
nor U15021 (N_15021,N_14073,N_13483);
and U15022 (N_15022,N_13225,N_14293);
xnor U15023 (N_15023,N_13336,N_14134);
nor U15024 (N_15024,N_13829,N_14029);
nor U15025 (N_15025,N_13316,N_13393);
or U15026 (N_15026,N_13512,N_13540);
nor U15027 (N_15027,N_14064,N_13415);
nor U15028 (N_15028,N_13607,N_13381);
nor U15029 (N_15029,N_13355,N_14272);
and U15030 (N_15030,N_14202,N_13449);
or U15031 (N_15031,N_13307,N_13937);
nor U15032 (N_15032,N_14089,N_13813);
or U15033 (N_15033,N_13989,N_13752);
xor U15034 (N_15034,N_14049,N_13492);
or U15035 (N_15035,N_14310,N_13989);
or U15036 (N_15036,N_13767,N_14160);
and U15037 (N_15037,N_13430,N_14026);
or U15038 (N_15038,N_13890,N_14127);
and U15039 (N_15039,N_13237,N_13801);
xnor U15040 (N_15040,N_14330,N_13542);
or U15041 (N_15041,N_13521,N_14087);
xnor U15042 (N_15042,N_13465,N_14296);
xor U15043 (N_15043,N_13304,N_14097);
nor U15044 (N_15044,N_13317,N_13391);
nand U15045 (N_15045,N_13779,N_13919);
xor U15046 (N_15046,N_14219,N_13437);
xor U15047 (N_15047,N_13574,N_14399);
nor U15048 (N_15048,N_13795,N_13847);
nand U15049 (N_15049,N_13212,N_13451);
nor U15050 (N_15050,N_13738,N_14210);
or U15051 (N_15051,N_14282,N_13659);
or U15052 (N_15052,N_14276,N_14381);
xor U15053 (N_15053,N_13973,N_13608);
nand U15054 (N_15054,N_13420,N_14283);
or U15055 (N_15055,N_13220,N_13460);
xor U15056 (N_15056,N_14058,N_14034);
or U15057 (N_15057,N_13548,N_14188);
nor U15058 (N_15058,N_14206,N_14054);
nor U15059 (N_15059,N_14262,N_13917);
xnor U15060 (N_15060,N_13367,N_13735);
or U15061 (N_15061,N_13554,N_13764);
or U15062 (N_15062,N_13844,N_13357);
or U15063 (N_15063,N_13589,N_14383);
and U15064 (N_15064,N_13307,N_13530);
nand U15065 (N_15065,N_14035,N_13580);
and U15066 (N_15066,N_13216,N_14062);
or U15067 (N_15067,N_13485,N_14177);
xor U15068 (N_15068,N_14136,N_13946);
nor U15069 (N_15069,N_14236,N_13876);
nand U15070 (N_15070,N_13421,N_14201);
or U15071 (N_15071,N_13696,N_13237);
xnor U15072 (N_15072,N_13784,N_13423);
nand U15073 (N_15073,N_13642,N_13332);
nor U15074 (N_15074,N_13920,N_13916);
xnor U15075 (N_15075,N_13693,N_14032);
or U15076 (N_15076,N_13407,N_13257);
or U15077 (N_15077,N_13657,N_13470);
and U15078 (N_15078,N_14360,N_13698);
xnor U15079 (N_15079,N_13337,N_13412);
xor U15080 (N_15080,N_14383,N_13264);
nand U15081 (N_15081,N_13751,N_13570);
xnor U15082 (N_15082,N_13509,N_13276);
or U15083 (N_15083,N_13330,N_14053);
nand U15084 (N_15084,N_13442,N_13417);
nor U15085 (N_15085,N_13204,N_13316);
and U15086 (N_15086,N_13243,N_13340);
or U15087 (N_15087,N_13986,N_14263);
or U15088 (N_15088,N_14301,N_13262);
and U15089 (N_15089,N_13227,N_13381);
or U15090 (N_15090,N_13266,N_13839);
xor U15091 (N_15091,N_13255,N_13375);
nor U15092 (N_15092,N_13904,N_13475);
or U15093 (N_15093,N_13579,N_13623);
and U15094 (N_15094,N_14054,N_13347);
xnor U15095 (N_15095,N_13942,N_14042);
nand U15096 (N_15096,N_14071,N_14012);
nand U15097 (N_15097,N_13494,N_14343);
nor U15098 (N_15098,N_14315,N_13522);
nand U15099 (N_15099,N_13241,N_13881);
xnor U15100 (N_15100,N_13394,N_13816);
nor U15101 (N_15101,N_14106,N_13209);
and U15102 (N_15102,N_13806,N_13874);
or U15103 (N_15103,N_13534,N_13434);
or U15104 (N_15104,N_13801,N_13749);
xor U15105 (N_15105,N_13303,N_13769);
nor U15106 (N_15106,N_14225,N_13256);
nor U15107 (N_15107,N_13434,N_13484);
nand U15108 (N_15108,N_13794,N_13981);
nor U15109 (N_15109,N_13903,N_13597);
nor U15110 (N_15110,N_13761,N_13230);
and U15111 (N_15111,N_14054,N_13562);
nor U15112 (N_15112,N_14022,N_14122);
or U15113 (N_15113,N_13592,N_13752);
or U15114 (N_15114,N_14224,N_13674);
xor U15115 (N_15115,N_14223,N_13513);
nor U15116 (N_15116,N_13842,N_13669);
nand U15117 (N_15117,N_13983,N_13631);
nor U15118 (N_15118,N_13261,N_14246);
nor U15119 (N_15119,N_14128,N_14113);
nor U15120 (N_15120,N_14256,N_13813);
and U15121 (N_15121,N_14067,N_13408);
nor U15122 (N_15122,N_13742,N_13489);
nand U15123 (N_15123,N_13764,N_14215);
nand U15124 (N_15124,N_14308,N_13658);
and U15125 (N_15125,N_14339,N_13312);
nand U15126 (N_15126,N_14086,N_14021);
nand U15127 (N_15127,N_13412,N_14237);
nor U15128 (N_15128,N_13650,N_13278);
or U15129 (N_15129,N_14388,N_13384);
nand U15130 (N_15130,N_13562,N_14324);
or U15131 (N_15131,N_14222,N_13385);
xnor U15132 (N_15132,N_14243,N_13698);
and U15133 (N_15133,N_14115,N_13448);
xor U15134 (N_15134,N_13559,N_13885);
xnor U15135 (N_15135,N_14323,N_14021);
nor U15136 (N_15136,N_14347,N_14255);
nand U15137 (N_15137,N_14017,N_14356);
xnor U15138 (N_15138,N_13946,N_13874);
and U15139 (N_15139,N_14239,N_13286);
xnor U15140 (N_15140,N_13392,N_13729);
nand U15141 (N_15141,N_13439,N_13351);
nor U15142 (N_15142,N_14038,N_13922);
or U15143 (N_15143,N_13600,N_14280);
or U15144 (N_15144,N_14368,N_13473);
or U15145 (N_15145,N_13453,N_13717);
nor U15146 (N_15146,N_13412,N_14035);
nor U15147 (N_15147,N_14364,N_13388);
nand U15148 (N_15148,N_14283,N_13416);
nor U15149 (N_15149,N_14290,N_13628);
or U15150 (N_15150,N_14357,N_14053);
xor U15151 (N_15151,N_13992,N_13687);
or U15152 (N_15152,N_13468,N_13757);
nor U15153 (N_15153,N_13485,N_14186);
nand U15154 (N_15154,N_13207,N_14247);
nor U15155 (N_15155,N_13772,N_13914);
xnor U15156 (N_15156,N_13360,N_13808);
nor U15157 (N_15157,N_13304,N_13920);
and U15158 (N_15158,N_14129,N_13308);
nor U15159 (N_15159,N_13341,N_13287);
nand U15160 (N_15160,N_13531,N_13688);
xor U15161 (N_15161,N_13403,N_14150);
nor U15162 (N_15162,N_13327,N_14213);
and U15163 (N_15163,N_14380,N_13772);
nand U15164 (N_15164,N_14353,N_13399);
nand U15165 (N_15165,N_13564,N_13833);
xnor U15166 (N_15166,N_13249,N_14272);
nand U15167 (N_15167,N_13441,N_14121);
xnor U15168 (N_15168,N_13990,N_14030);
and U15169 (N_15169,N_13396,N_13827);
nor U15170 (N_15170,N_14230,N_13640);
and U15171 (N_15171,N_14001,N_14263);
and U15172 (N_15172,N_13608,N_13276);
xor U15173 (N_15173,N_13507,N_14218);
nand U15174 (N_15174,N_14078,N_13624);
xor U15175 (N_15175,N_13318,N_14199);
or U15176 (N_15176,N_14121,N_13240);
nand U15177 (N_15177,N_14160,N_13779);
nor U15178 (N_15178,N_13609,N_13248);
nand U15179 (N_15179,N_13673,N_13372);
or U15180 (N_15180,N_14304,N_13713);
xor U15181 (N_15181,N_13461,N_13320);
nor U15182 (N_15182,N_14121,N_13602);
nand U15183 (N_15183,N_13950,N_14209);
or U15184 (N_15184,N_13824,N_13881);
xnor U15185 (N_15185,N_13797,N_13915);
nor U15186 (N_15186,N_13762,N_13224);
nor U15187 (N_15187,N_13982,N_14304);
or U15188 (N_15188,N_13909,N_13673);
xor U15189 (N_15189,N_13793,N_14215);
xnor U15190 (N_15190,N_14171,N_14239);
xnor U15191 (N_15191,N_13478,N_14277);
nor U15192 (N_15192,N_14058,N_13299);
nand U15193 (N_15193,N_13713,N_13267);
and U15194 (N_15194,N_13930,N_13585);
nand U15195 (N_15195,N_13818,N_13509);
and U15196 (N_15196,N_13603,N_13865);
or U15197 (N_15197,N_14022,N_14160);
or U15198 (N_15198,N_13220,N_14345);
nor U15199 (N_15199,N_13996,N_14265);
nand U15200 (N_15200,N_14143,N_14226);
and U15201 (N_15201,N_13910,N_14029);
xor U15202 (N_15202,N_14140,N_13330);
and U15203 (N_15203,N_13558,N_13204);
nand U15204 (N_15204,N_13250,N_14024);
nand U15205 (N_15205,N_13315,N_13399);
xor U15206 (N_15206,N_14300,N_13651);
xor U15207 (N_15207,N_13403,N_14082);
and U15208 (N_15208,N_13514,N_13785);
or U15209 (N_15209,N_14231,N_13385);
nor U15210 (N_15210,N_13968,N_13633);
and U15211 (N_15211,N_14392,N_14387);
nor U15212 (N_15212,N_13434,N_13855);
or U15213 (N_15213,N_13447,N_13642);
nor U15214 (N_15214,N_13352,N_14293);
nand U15215 (N_15215,N_13604,N_13453);
or U15216 (N_15216,N_13248,N_13660);
or U15217 (N_15217,N_13959,N_14326);
nor U15218 (N_15218,N_13841,N_13701);
xnor U15219 (N_15219,N_13304,N_13237);
nor U15220 (N_15220,N_13681,N_13382);
or U15221 (N_15221,N_13249,N_13537);
nand U15222 (N_15222,N_13722,N_13765);
or U15223 (N_15223,N_14197,N_14109);
and U15224 (N_15224,N_13546,N_13911);
xnor U15225 (N_15225,N_13758,N_14133);
nor U15226 (N_15226,N_13555,N_14157);
or U15227 (N_15227,N_14277,N_13582);
nor U15228 (N_15228,N_13718,N_13713);
and U15229 (N_15229,N_13431,N_13999);
xnor U15230 (N_15230,N_13443,N_13584);
or U15231 (N_15231,N_14368,N_13272);
or U15232 (N_15232,N_13937,N_13260);
nand U15233 (N_15233,N_13287,N_13518);
nor U15234 (N_15234,N_14018,N_14159);
or U15235 (N_15235,N_13882,N_13823);
xor U15236 (N_15236,N_13484,N_13388);
or U15237 (N_15237,N_14046,N_14085);
and U15238 (N_15238,N_14271,N_13545);
nand U15239 (N_15239,N_13734,N_13532);
or U15240 (N_15240,N_14115,N_14286);
or U15241 (N_15241,N_13261,N_14334);
and U15242 (N_15242,N_13230,N_14187);
and U15243 (N_15243,N_14032,N_13658);
nand U15244 (N_15244,N_14235,N_14375);
and U15245 (N_15245,N_13597,N_14399);
xor U15246 (N_15246,N_14064,N_13588);
xor U15247 (N_15247,N_13713,N_14351);
and U15248 (N_15248,N_13888,N_13889);
nor U15249 (N_15249,N_13899,N_13579);
xor U15250 (N_15250,N_13315,N_13460);
nor U15251 (N_15251,N_13587,N_13805);
and U15252 (N_15252,N_13386,N_14050);
nor U15253 (N_15253,N_13844,N_14060);
nand U15254 (N_15254,N_14236,N_13734);
and U15255 (N_15255,N_13747,N_13719);
nand U15256 (N_15256,N_13542,N_14219);
nand U15257 (N_15257,N_13444,N_14337);
nor U15258 (N_15258,N_13826,N_14258);
nand U15259 (N_15259,N_13902,N_13993);
nor U15260 (N_15260,N_14213,N_13934);
or U15261 (N_15261,N_14256,N_14164);
nand U15262 (N_15262,N_13611,N_13418);
nor U15263 (N_15263,N_13748,N_14109);
nor U15264 (N_15264,N_13886,N_14098);
xnor U15265 (N_15265,N_14177,N_14022);
or U15266 (N_15266,N_14296,N_13220);
nand U15267 (N_15267,N_14126,N_13316);
nor U15268 (N_15268,N_13571,N_13448);
and U15269 (N_15269,N_13805,N_13570);
or U15270 (N_15270,N_13291,N_14212);
and U15271 (N_15271,N_14188,N_14085);
nand U15272 (N_15272,N_13966,N_14232);
and U15273 (N_15273,N_13678,N_13636);
nor U15274 (N_15274,N_13389,N_14115);
or U15275 (N_15275,N_13740,N_13657);
xor U15276 (N_15276,N_13461,N_13234);
nor U15277 (N_15277,N_13934,N_13884);
and U15278 (N_15278,N_14128,N_13558);
nor U15279 (N_15279,N_13678,N_13416);
or U15280 (N_15280,N_13728,N_13664);
or U15281 (N_15281,N_13685,N_13540);
nor U15282 (N_15282,N_14186,N_13722);
nor U15283 (N_15283,N_13819,N_13230);
nor U15284 (N_15284,N_13751,N_14019);
or U15285 (N_15285,N_13384,N_13745);
and U15286 (N_15286,N_14028,N_13324);
nand U15287 (N_15287,N_13834,N_14004);
xor U15288 (N_15288,N_13742,N_14131);
xor U15289 (N_15289,N_13528,N_14331);
nand U15290 (N_15290,N_13830,N_14295);
and U15291 (N_15291,N_13897,N_13637);
and U15292 (N_15292,N_13764,N_13280);
xnor U15293 (N_15293,N_13991,N_14284);
or U15294 (N_15294,N_13547,N_14368);
and U15295 (N_15295,N_13335,N_13393);
nand U15296 (N_15296,N_13375,N_13430);
and U15297 (N_15297,N_13265,N_14399);
xnor U15298 (N_15298,N_14340,N_14175);
nand U15299 (N_15299,N_13230,N_13766);
nand U15300 (N_15300,N_13354,N_14385);
xor U15301 (N_15301,N_14138,N_14329);
or U15302 (N_15302,N_13258,N_13566);
nor U15303 (N_15303,N_13519,N_14325);
and U15304 (N_15304,N_13454,N_13530);
and U15305 (N_15305,N_13571,N_13636);
xor U15306 (N_15306,N_13342,N_14262);
and U15307 (N_15307,N_14366,N_14391);
or U15308 (N_15308,N_13939,N_14033);
nor U15309 (N_15309,N_14168,N_13514);
nor U15310 (N_15310,N_13200,N_14356);
and U15311 (N_15311,N_13832,N_14077);
nand U15312 (N_15312,N_14208,N_13718);
or U15313 (N_15313,N_13238,N_13441);
xnor U15314 (N_15314,N_14234,N_13544);
or U15315 (N_15315,N_13662,N_13921);
or U15316 (N_15316,N_13207,N_13553);
and U15317 (N_15317,N_13730,N_13923);
or U15318 (N_15318,N_13375,N_13555);
and U15319 (N_15319,N_13442,N_13980);
nor U15320 (N_15320,N_14188,N_13763);
nor U15321 (N_15321,N_14242,N_13341);
xor U15322 (N_15322,N_14160,N_13629);
and U15323 (N_15323,N_13794,N_13275);
xnor U15324 (N_15324,N_13584,N_13372);
nand U15325 (N_15325,N_13352,N_13493);
or U15326 (N_15326,N_13458,N_14370);
xor U15327 (N_15327,N_13259,N_13955);
xnor U15328 (N_15328,N_13811,N_13704);
nand U15329 (N_15329,N_14061,N_14300);
and U15330 (N_15330,N_14214,N_14010);
nand U15331 (N_15331,N_13257,N_14312);
xor U15332 (N_15332,N_14158,N_14241);
xor U15333 (N_15333,N_14002,N_13332);
xnor U15334 (N_15334,N_13932,N_14172);
or U15335 (N_15335,N_13240,N_13361);
nand U15336 (N_15336,N_13908,N_13914);
and U15337 (N_15337,N_14094,N_13857);
nand U15338 (N_15338,N_14026,N_13932);
xnor U15339 (N_15339,N_13460,N_13449);
and U15340 (N_15340,N_13877,N_14041);
or U15341 (N_15341,N_14234,N_13309);
and U15342 (N_15342,N_13977,N_13205);
nor U15343 (N_15343,N_13753,N_13486);
and U15344 (N_15344,N_13807,N_13783);
or U15345 (N_15345,N_14375,N_14324);
and U15346 (N_15346,N_14053,N_13804);
xor U15347 (N_15347,N_13759,N_13933);
xnor U15348 (N_15348,N_14297,N_14112);
and U15349 (N_15349,N_13609,N_13670);
nand U15350 (N_15350,N_13873,N_13526);
nand U15351 (N_15351,N_14128,N_14297);
nor U15352 (N_15352,N_14052,N_14341);
and U15353 (N_15353,N_13258,N_13222);
nor U15354 (N_15354,N_13874,N_14265);
and U15355 (N_15355,N_13959,N_13870);
nor U15356 (N_15356,N_13730,N_13456);
nand U15357 (N_15357,N_13496,N_13967);
or U15358 (N_15358,N_13838,N_13482);
or U15359 (N_15359,N_14143,N_13930);
xor U15360 (N_15360,N_14232,N_14212);
and U15361 (N_15361,N_13841,N_13825);
nand U15362 (N_15362,N_13538,N_14009);
or U15363 (N_15363,N_14237,N_13227);
nand U15364 (N_15364,N_14154,N_13314);
and U15365 (N_15365,N_13394,N_13622);
nor U15366 (N_15366,N_13490,N_14187);
and U15367 (N_15367,N_13765,N_13526);
nand U15368 (N_15368,N_13994,N_14184);
xor U15369 (N_15369,N_14087,N_13987);
nand U15370 (N_15370,N_13752,N_13308);
xor U15371 (N_15371,N_14031,N_13266);
xnor U15372 (N_15372,N_14107,N_13478);
nor U15373 (N_15373,N_14143,N_14053);
xor U15374 (N_15374,N_13534,N_14025);
xnor U15375 (N_15375,N_14185,N_13218);
nand U15376 (N_15376,N_13262,N_14387);
xor U15377 (N_15377,N_13479,N_13501);
nand U15378 (N_15378,N_13503,N_14257);
nor U15379 (N_15379,N_14182,N_13945);
nor U15380 (N_15380,N_13249,N_13257);
xor U15381 (N_15381,N_14255,N_13728);
xor U15382 (N_15382,N_13692,N_13627);
nand U15383 (N_15383,N_13575,N_14355);
nand U15384 (N_15384,N_13904,N_13255);
nand U15385 (N_15385,N_13843,N_14147);
nand U15386 (N_15386,N_13522,N_13421);
nand U15387 (N_15387,N_13837,N_14388);
or U15388 (N_15388,N_13708,N_14170);
and U15389 (N_15389,N_14020,N_14307);
nand U15390 (N_15390,N_14016,N_13692);
and U15391 (N_15391,N_13643,N_13891);
xor U15392 (N_15392,N_14013,N_13316);
or U15393 (N_15393,N_14260,N_13765);
or U15394 (N_15394,N_13834,N_13548);
nor U15395 (N_15395,N_13684,N_13924);
nand U15396 (N_15396,N_13951,N_13366);
or U15397 (N_15397,N_14113,N_14208);
and U15398 (N_15398,N_13375,N_13808);
xor U15399 (N_15399,N_13923,N_13414);
nand U15400 (N_15400,N_13698,N_14103);
nor U15401 (N_15401,N_14069,N_13758);
and U15402 (N_15402,N_13217,N_13995);
and U15403 (N_15403,N_14020,N_14342);
or U15404 (N_15404,N_14112,N_13271);
nand U15405 (N_15405,N_13759,N_13343);
xnor U15406 (N_15406,N_13694,N_13958);
and U15407 (N_15407,N_13929,N_13207);
nand U15408 (N_15408,N_14277,N_14229);
or U15409 (N_15409,N_13823,N_13586);
nand U15410 (N_15410,N_14271,N_14073);
nor U15411 (N_15411,N_13473,N_13490);
nand U15412 (N_15412,N_13958,N_14215);
xnor U15413 (N_15413,N_13568,N_13620);
and U15414 (N_15414,N_14234,N_13304);
or U15415 (N_15415,N_13387,N_13310);
xnor U15416 (N_15416,N_13876,N_13330);
or U15417 (N_15417,N_13804,N_13492);
xor U15418 (N_15418,N_13296,N_13881);
xnor U15419 (N_15419,N_13891,N_13901);
and U15420 (N_15420,N_13711,N_13916);
or U15421 (N_15421,N_13212,N_14245);
or U15422 (N_15422,N_13717,N_13895);
nor U15423 (N_15423,N_13234,N_14019);
nand U15424 (N_15424,N_13531,N_13991);
nand U15425 (N_15425,N_13467,N_13601);
xnor U15426 (N_15426,N_13903,N_13200);
and U15427 (N_15427,N_13643,N_14337);
nand U15428 (N_15428,N_13898,N_13395);
or U15429 (N_15429,N_13876,N_13942);
or U15430 (N_15430,N_13800,N_14292);
xor U15431 (N_15431,N_13398,N_13305);
nand U15432 (N_15432,N_13833,N_13970);
nor U15433 (N_15433,N_13306,N_14378);
and U15434 (N_15434,N_13347,N_13917);
or U15435 (N_15435,N_13726,N_13472);
or U15436 (N_15436,N_13864,N_13807);
and U15437 (N_15437,N_14015,N_13376);
nand U15438 (N_15438,N_13906,N_14094);
or U15439 (N_15439,N_14172,N_13287);
nor U15440 (N_15440,N_13803,N_13262);
and U15441 (N_15441,N_13948,N_13939);
or U15442 (N_15442,N_13980,N_13983);
xnor U15443 (N_15443,N_13975,N_13748);
and U15444 (N_15444,N_13356,N_13747);
and U15445 (N_15445,N_13344,N_14125);
and U15446 (N_15446,N_13881,N_13876);
or U15447 (N_15447,N_13611,N_13844);
or U15448 (N_15448,N_13490,N_13767);
nor U15449 (N_15449,N_14114,N_13232);
nand U15450 (N_15450,N_13524,N_13218);
xor U15451 (N_15451,N_13320,N_13890);
or U15452 (N_15452,N_14238,N_14026);
and U15453 (N_15453,N_14341,N_14135);
nor U15454 (N_15454,N_13309,N_14040);
or U15455 (N_15455,N_14189,N_13939);
nand U15456 (N_15456,N_14173,N_13836);
nand U15457 (N_15457,N_13330,N_13947);
nand U15458 (N_15458,N_14260,N_13591);
or U15459 (N_15459,N_14346,N_14265);
xnor U15460 (N_15460,N_13572,N_13496);
nand U15461 (N_15461,N_13602,N_14329);
xnor U15462 (N_15462,N_13718,N_13295);
and U15463 (N_15463,N_14020,N_14366);
nor U15464 (N_15464,N_13775,N_13533);
and U15465 (N_15465,N_13956,N_13791);
xnor U15466 (N_15466,N_14224,N_13236);
nor U15467 (N_15467,N_13714,N_13601);
and U15468 (N_15468,N_13445,N_14076);
xor U15469 (N_15469,N_14387,N_14220);
nand U15470 (N_15470,N_14157,N_14313);
xor U15471 (N_15471,N_14044,N_13563);
or U15472 (N_15472,N_13408,N_13626);
xnor U15473 (N_15473,N_13357,N_13696);
nor U15474 (N_15474,N_14185,N_13389);
nor U15475 (N_15475,N_13319,N_13265);
or U15476 (N_15476,N_13232,N_13562);
and U15477 (N_15477,N_13811,N_13800);
xor U15478 (N_15478,N_13890,N_14362);
xor U15479 (N_15479,N_14196,N_14357);
nor U15480 (N_15480,N_13872,N_14345);
and U15481 (N_15481,N_13969,N_13727);
nand U15482 (N_15482,N_14067,N_13264);
and U15483 (N_15483,N_13696,N_13676);
nor U15484 (N_15484,N_13908,N_13706);
nor U15485 (N_15485,N_13941,N_13209);
nor U15486 (N_15486,N_13682,N_13946);
nand U15487 (N_15487,N_13992,N_14268);
nand U15488 (N_15488,N_13681,N_13645);
xor U15489 (N_15489,N_14028,N_13845);
and U15490 (N_15490,N_13499,N_13245);
or U15491 (N_15491,N_13773,N_13769);
and U15492 (N_15492,N_13530,N_14043);
nand U15493 (N_15493,N_13831,N_13378);
nand U15494 (N_15494,N_13839,N_13317);
nand U15495 (N_15495,N_14070,N_14125);
xnor U15496 (N_15496,N_14240,N_14075);
or U15497 (N_15497,N_13813,N_13541);
nand U15498 (N_15498,N_13986,N_13522);
nand U15499 (N_15499,N_13475,N_13971);
nor U15500 (N_15500,N_13580,N_13913);
and U15501 (N_15501,N_14011,N_13825);
nand U15502 (N_15502,N_14088,N_13807);
xor U15503 (N_15503,N_13820,N_14257);
or U15504 (N_15504,N_13412,N_13640);
xor U15505 (N_15505,N_14055,N_13521);
nor U15506 (N_15506,N_13921,N_13741);
nor U15507 (N_15507,N_14256,N_14163);
xnor U15508 (N_15508,N_13760,N_13776);
nand U15509 (N_15509,N_14129,N_13479);
nor U15510 (N_15510,N_14178,N_14239);
or U15511 (N_15511,N_13703,N_13827);
xor U15512 (N_15512,N_13950,N_14072);
or U15513 (N_15513,N_13301,N_14252);
nand U15514 (N_15514,N_13314,N_13985);
or U15515 (N_15515,N_13737,N_13853);
nand U15516 (N_15516,N_14118,N_14327);
and U15517 (N_15517,N_13576,N_13981);
or U15518 (N_15518,N_14025,N_13275);
nor U15519 (N_15519,N_14087,N_13806);
nand U15520 (N_15520,N_13863,N_14023);
xor U15521 (N_15521,N_13360,N_13401);
and U15522 (N_15522,N_14113,N_13506);
xnor U15523 (N_15523,N_13590,N_13253);
nand U15524 (N_15524,N_14283,N_13739);
xnor U15525 (N_15525,N_13634,N_13559);
nand U15526 (N_15526,N_13348,N_14062);
nand U15527 (N_15527,N_14096,N_14158);
or U15528 (N_15528,N_13858,N_14271);
nor U15529 (N_15529,N_13423,N_13292);
xor U15530 (N_15530,N_13607,N_13946);
nand U15531 (N_15531,N_13554,N_13662);
and U15532 (N_15532,N_13925,N_13793);
xor U15533 (N_15533,N_13500,N_14026);
nand U15534 (N_15534,N_13527,N_14031);
or U15535 (N_15535,N_13892,N_14049);
xnor U15536 (N_15536,N_13939,N_13346);
or U15537 (N_15537,N_14243,N_13959);
and U15538 (N_15538,N_13536,N_14363);
nand U15539 (N_15539,N_13448,N_13615);
and U15540 (N_15540,N_13929,N_14363);
nand U15541 (N_15541,N_13947,N_14032);
and U15542 (N_15542,N_13937,N_13725);
nand U15543 (N_15543,N_13252,N_14286);
xnor U15544 (N_15544,N_13343,N_13602);
xor U15545 (N_15545,N_14320,N_14107);
nand U15546 (N_15546,N_14370,N_13600);
xnor U15547 (N_15547,N_13929,N_13400);
nor U15548 (N_15548,N_13966,N_13326);
nor U15549 (N_15549,N_13859,N_13249);
nand U15550 (N_15550,N_14172,N_14281);
xnor U15551 (N_15551,N_13425,N_13583);
and U15552 (N_15552,N_14378,N_13581);
and U15553 (N_15553,N_13428,N_13293);
nor U15554 (N_15554,N_13930,N_14231);
nor U15555 (N_15555,N_14002,N_14385);
or U15556 (N_15556,N_13769,N_13523);
and U15557 (N_15557,N_13349,N_14353);
and U15558 (N_15558,N_14298,N_13393);
or U15559 (N_15559,N_14121,N_13835);
or U15560 (N_15560,N_13334,N_13530);
or U15561 (N_15561,N_13450,N_13205);
and U15562 (N_15562,N_13366,N_14172);
nand U15563 (N_15563,N_13551,N_13934);
nand U15564 (N_15564,N_14342,N_14387);
xor U15565 (N_15565,N_14138,N_14000);
nor U15566 (N_15566,N_14039,N_14346);
xnor U15567 (N_15567,N_13762,N_13776);
nand U15568 (N_15568,N_14223,N_13695);
or U15569 (N_15569,N_13374,N_14213);
or U15570 (N_15570,N_13759,N_13536);
and U15571 (N_15571,N_14353,N_13804);
xnor U15572 (N_15572,N_13266,N_13328);
xnor U15573 (N_15573,N_14390,N_13935);
and U15574 (N_15574,N_14282,N_13933);
nor U15575 (N_15575,N_14186,N_13854);
nand U15576 (N_15576,N_14211,N_13677);
and U15577 (N_15577,N_14094,N_13712);
and U15578 (N_15578,N_14016,N_14200);
or U15579 (N_15579,N_13212,N_13458);
nand U15580 (N_15580,N_13868,N_13733);
xor U15581 (N_15581,N_13397,N_13657);
nor U15582 (N_15582,N_14280,N_14160);
or U15583 (N_15583,N_13278,N_14197);
nor U15584 (N_15584,N_13387,N_13627);
nand U15585 (N_15585,N_13977,N_13872);
and U15586 (N_15586,N_14000,N_13392);
and U15587 (N_15587,N_13443,N_13652);
nor U15588 (N_15588,N_14375,N_13803);
or U15589 (N_15589,N_13512,N_14020);
and U15590 (N_15590,N_14293,N_13298);
or U15591 (N_15591,N_14239,N_13846);
xnor U15592 (N_15592,N_13896,N_14040);
or U15593 (N_15593,N_13274,N_13581);
xor U15594 (N_15594,N_13714,N_14055);
or U15595 (N_15595,N_14199,N_13419);
xor U15596 (N_15596,N_14280,N_14338);
xnor U15597 (N_15597,N_14201,N_14025);
nand U15598 (N_15598,N_13761,N_13970);
and U15599 (N_15599,N_13455,N_13841);
nand U15600 (N_15600,N_14670,N_15011);
xor U15601 (N_15601,N_15173,N_15127);
and U15602 (N_15602,N_15353,N_14913);
nor U15603 (N_15603,N_15258,N_15133);
or U15604 (N_15604,N_15002,N_14682);
or U15605 (N_15605,N_14633,N_15150);
nor U15606 (N_15606,N_15076,N_14891);
nand U15607 (N_15607,N_14622,N_14779);
nand U15608 (N_15608,N_15511,N_15325);
nor U15609 (N_15609,N_14617,N_15346);
nand U15610 (N_15610,N_15085,N_15383);
xor U15611 (N_15611,N_14515,N_15236);
or U15612 (N_15612,N_14483,N_15340);
or U15613 (N_15613,N_15341,N_14951);
nand U15614 (N_15614,N_14509,N_15196);
or U15615 (N_15615,N_15223,N_14772);
xnor U15616 (N_15616,N_14794,N_15359);
nor U15617 (N_15617,N_15301,N_14587);
xor U15618 (N_15618,N_15277,N_15303);
or U15619 (N_15619,N_15452,N_15566);
nor U15620 (N_15620,N_14853,N_14773);
or U15621 (N_15621,N_14992,N_14921);
or U15622 (N_15622,N_15414,N_15039);
xnor U15623 (N_15623,N_15220,N_14415);
and U15624 (N_15624,N_15231,N_15265);
or U15625 (N_15625,N_15191,N_14973);
and U15626 (N_15626,N_14920,N_14726);
and U15627 (N_15627,N_14742,N_14411);
nor U15628 (N_15628,N_14657,N_14807);
and U15629 (N_15629,N_14828,N_15105);
nand U15630 (N_15630,N_15262,N_14578);
nor U15631 (N_15631,N_15443,N_15015);
or U15632 (N_15632,N_14529,N_15048);
and U15633 (N_15633,N_14996,N_14881);
nor U15634 (N_15634,N_15007,N_14997);
xnor U15635 (N_15635,N_14746,N_15203);
or U15636 (N_15636,N_14601,N_14623);
nor U15637 (N_15637,N_14639,N_15115);
nand U15638 (N_15638,N_15156,N_15238);
xnor U15639 (N_15639,N_14851,N_15336);
or U15640 (N_15640,N_15142,N_14542);
nand U15641 (N_15641,N_15497,N_15531);
xor U15642 (N_15642,N_14660,N_14735);
or U15643 (N_15643,N_15058,N_14539);
xnor U15644 (N_15644,N_15400,N_14986);
nand U15645 (N_15645,N_15369,N_15013);
nand U15646 (N_15646,N_15317,N_14892);
xnor U15647 (N_15647,N_14497,N_14982);
nor U15648 (N_15648,N_15348,N_15418);
nand U15649 (N_15649,N_14655,N_14981);
and U15650 (N_15650,N_14780,N_15559);
or U15651 (N_15651,N_14778,N_14548);
nand U15652 (N_15652,N_15478,N_15561);
and U15653 (N_15653,N_14522,N_14857);
or U15654 (N_15654,N_14716,N_14987);
nor U15655 (N_15655,N_15463,N_14957);
nor U15656 (N_15656,N_14518,N_14607);
nand U15657 (N_15657,N_15001,N_14696);
nor U15658 (N_15658,N_14948,N_15054);
or U15659 (N_15659,N_14424,N_14532);
and U15660 (N_15660,N_15329,N_15404);
xnor U15661 (N_15661,N_14896,N_15392);
xor U15662 (N_15662,N_15316,N_15240);
or U15663 (N_15663,N_14612,N_15576);
nand U15664 (N_15664,N_14443,N_15368);
xor U15665 (N_15665,N_14757,N_15060);
xnor U15666 (N_15666,N_14975,N_15287);
nor U15667 (N_15667,N_14567,N_15524);
nand U15668 (N_15668,N_15206,N_15064);
xor U15669 (N_15669,N_15063,N_14688);
nor U15670 (N_15670,N_14749,N_14441);
nand U15671 (N_15671,N_14756,N_15382);
xor U15672 (N_15672,N_14668,N_15094);
nand U15673 (N_15673,N_15439,N_14444);
xor U15674 (N_15674,N_15069,N_14449);
and U15675 (N_15675,N_14827,N_14985);
nor U15676 (N_15676,N_15189,N_14915);
and U15677 (N_15677,N_15041,N_14816);
xor U15678 (N_15678,N_15185,N_14802);
nand U15679 (N_15679,N_15519,N_14481);
xnor U15680 (N_15680,N_14419,N_15098);
and U15681 (N_15681,N_14950,N_15592);
or U15682 (N_15682,N_15072,N_15153);
xnor U15683 (N_15683,N_14903,N_14909);
and U15684 (N_15684,N_15209,N_15045);
and U15685 (N_15685,N_15466,N_14648);
xor U15686 (N_15686,N_14651,N_14905);
xnor U15687 (N_15687,N_14882,N_14430);
nand U15688 (N_15688,N_15249,N_15577);
xnor U15689 (N_15689,N_14519,N_15299);
xor U15690 (N_15690,N_14761,N_14733);
or U15691 (N_15691,N_14849,N_14584);
nor U15692 (N_15692,N_14942,N_14410);
xnor U15693 (N_15693,N_14631,N_14962);
or U15694 (N_15694,N_15406,N_14573);
or U15695 (N_15695,N_15009,N_15237);
xor U15696 (N_15696,N_15527,N_14740);
nand U15697 (N_15697,N_15176,N_14721);
xor U15698 (N_15698,N_14416,N_14421);
and U15699 (N_15699,N_14686,N_14971);
nor U15700 (N_15700,N_14910,N_14654);
or U15701 (N_15701,N_14945,N_14669);
and U15702 (N_15702,N_14938,N_15071);
and U15703 (N_15703,N_14597,N_15283);
or U15704 (N_15704,N_15148,N_15145);
nor U15705 (N_15705,N_14640,N_14408);
xnor U15706 (N_15706,N_15005,N_15449);
nor U15707 (N_15707,N_15432,N_14466);
or U15708 (N_15708,N_15417,N_15456);
xor U15709 (N_15709,N_14561,N_15170);
nor U15710 (N_15710,N_15590,N_15228);
nor U15711 (N_15711,N_15377,N_15210);
or U15712 (N_15712,N_15372,N_15451);
nand U15713 (N_15713,N_15006,N_15308);
nor U15714 (N_15714,N_15583,N_15214);
nor U15715 (N_15715,N_15461,N_15518);
nor U15716 (N_15716,N_14732,N_14711);
xor U15717 (N_15717,N_14628,N_15430);
xor U15718 (N_15718,N_15345,N_15104);
and U15719 (N_15719,N_14953,N_15255);
or U15720 (N_15720,N_14439,N_14402);
xor U15721 (N_15721,N_15455,N_15057);
or U15722 (N_15722,N_15154,N_15295);
xor U15723 (N_15723,N_14646,N_14469);
nand U15724 (N_15724,N_14559,N_14712);
xor U15725 (N_15725,N_15043,N_15597);
or U15726 (N_15726,N_15163,N_15389);
nand U15727 (N_15727,N_15416,N_14693);
and U15728 (N_15728,N_15288,N_14877);
nor U15729 (N_15729,N_15136,N_15355);
nor U15730 (N_15730,N_14830,N_15207);
or U15731 (N_15731,N_14786,N_15294);
nand U15732 (N_15732,N_14453,N_14709);
nor U15733 (N_15733,N_15252,N_15164);
nor U15734 (N_15734,N_14530,N_15014);
xnor U15735 (N_15735,N_14847,N_14689);
and U15736 (N_15736,N_15268,N_15289);
nor U15737 (N_15737,N_14511,N_14999);
xor U15738 (N_15738,N_15574,N_14704);
nand U15739 (N_15739,N_15134,N_15378);
nand U15740 (N_15740,N_15211,N_14661);
nor U15741 (N_15741,N_14618,N_14609);
nor U15742 (N_15742,N_15501,N_14543);
nand U15743 (N_15743,N_15422,N_15259);
or U15744 (N_15744,N_15568,N_15110);
or U15745 (N_15745,N_15297,N_14610);
and U15746 (N_15746,N_15504,N_15050);
nand U15747 (N_15747,N_15447,N_14840);
nor U15748 (N_15748,N_14846,N_14902);
and U15749 (N_15749,N_15351,N_14884);
nand U15750 (N_15750,N_14747,N_15507);
xnor U15751 (N_15751,N_15350,N_15394);
and U15752 (N_15752,N_15281,N_15138);
xnor U15753 (N_15753,N_14484,N_14460);
or U15754 (N_15754,N_14429,N_15485);
xor U15755 (N_15755,N_14553,N_15594);
xor U15756 (N_15756,N_14538,N_15126);
nor U15757 (N_15757,N_15526,N_15251);
nor U15758 (N_15758,N_14673,N_15472);
nor U15759 (N_15759,N_14782,N_15309);
or U15760 (N_15760,N_14810,N_14671);
nor U15761 (N_15761,N_14893,N_15197);
or U15762 (N_15762,N_14722,N_14455);
xor U15763 (N_15763,N_14431,N_15547);
or U15764 (N_15764,N_14858,N_15423);
nor U15765 (N_15765,N_14477,N_15147);
and U15766 (N_15766,N_15569,N_14492);
or U15767 (N_15767,N_15062,N_15032);
nor U15768 (N_15768,N_14582,N_14546);
nand U15769 (N_15769,N_14959,N_15161);
nor U15770 (N_15770,N_15402,N_14860);
nand U15771 (N_15771,N_15356,N_14545);
nor U15772 (N_15772,N_15230,N_14754);
or U15773 (N_15773,N_15513,N_15122);
nand U15774 (N_15774,N_15084,N_14937);
xor U15775 (N_15775,N_15354,N_14621);
nand U15776 (N_15776,N_15181,N_15343);
nor U15777 (N_15777,N_15300,N_14461);
nor U15778 (N_15778,N_14974,N_14777);
xor U15779 (N_15779,N_14991,N_14656);
nor U15780 (N_15780,N_14977,N_15139);
nor U15781 (N_15781,N_15522,N_15427);
or U15782 (N_15782,N_15381,N_14895);
nand U15783 (N_15783,N_15521,N_14922);
or U15784 (N_15784,N_15362,N_14800);
and U15785 (N_15785,N_14448,N_15235);
xor U15786 (N_15786,N_15051,N_15286);
and U15787 (N_15787,N_14536,N_15208);
nand U15788 (N_15788,N_14967,N_14459);
nand U15789 (N_15789,N_15232,N_14620);
and U15790 (N_15790,N_15114,N_15487);
nand U15791 (N_15791,N_14474,N_15587);
and U15792 (N_15792,N_14580,N_14564);
nand U15793 (N_15793,N_14521,N_14739);
xnor U15794 (N_15794,N_14450,N_15412);
and U15795 (N_15795,N_15589,N_15315);
and U15796 (N_15796,N_14540,N_15118);
xnor U15797 (N_15797,N_15477,N_14947);
nor U15798 (N_15798,N_14629,N_14832);
nand U15799 (N_15799,N_15313,N_14404);
nand U15800 (N_15800,N_14728,N_14883);
nand U15801 (N_15801,N_15508,N_15549);
or U15802 (N_15802,N_15229,N_15182);
xnor U15803 (N_15803,N_14730,N_14941);
or U15804 (N_15804,N_14944,N_14720);
nor U15805 (N_15805,N_14551,N_14767);
xnor U15806 (N_15806,N_14845,N_15323);
nor U15807 (N_15807,N_15465,N_15266);
and U15808 (N_15808,N_14715,N_14650);
xor U15809 (N_15809,N_14486,N_15371);
or U15810 (N_15810,N_14939,N_15012);
nand U15811 (N_15811,N_14577,N_14598);
and U15812 (N_15812,N_15520,N_14811);
and U15813 (N_15813,N_14787,N_15111);
xor U15814 (N_15814,N_15538,N_14642);
nand U15815 (N_15815,N_15246,N_14718);
or U15816 (N_15816,N_14960,N_14914);
nand U15817 (N_15817,N_15517,N_14784);
nor U15818 (N_15818,N_15320,N_15029);
and U15819 (N_15819,N_15221,N_14501);
and U15820 (N_15820,N_14700,N_14889);
and U15821 (N_15821,N_15264,N_14979);
xnor U15822 (N_15822,N_15375,N_14769);
nor U15823 (N_15823,N_14908,N_14978);
and U15824 (N_15824,N_14652,N_14403);
nor U15825 (N_15825,N_14763,N_15448);
or U15826 (N_15826,N_15425,N_14936);
or U15827 (N_15827,N_14994,N_14468);
or U15828 (N_15828,N_15036,N_15274);
or U15829 (N_15829,N_15100,N_14758);
xnor U15830 (N_15830,N_15324,N_14581);
or U15831 (N_15831,N_15370,N_14894);
nand U15832 (N_15832,N_15505,N_14478);
nor U15833 (N_15833,N_15498,N_15494);
or U15834 (N_15834,N_15386,N_15401);
or U15835 (N_15835,N_15290,N_14886);
and U15836 (N_15836,N_14899,N_15380);
nand U15837 (N_15837,N_15088,N_14852);
or U15838 (N_15838,N_14980,N_14674);
and U15839 (N_15839,N_14644,N_15398);
and U15840 (N_15840,N_14822,N_15437);
xor U15841 (N_15841,N_15390,N_15363);
xor U15842 (N_15842,N_14645,N_15555);
nand U15843 (N_15843,N_14880,N_14666);
xnor U15844 (N_15844,N_15140,N_14890);
nor U15845 (N_15845,N_14727,N_15434);
or U15846 (N_15846,N_15040,N_14871);
nor U15847 (N_15847,N_14569,N_15467);
nor U15848 (N_15848,N_14848,N_15061);
or U15849 (N_15849,N_15541,N_15020);
or U15850 (N_15850,N_14467,N_15095);
nand U15851 (N_15851,N_14672,N_15066);
nand U15852 (N_15852,N_15585,N_15241);
nor U15853 (N_15853,N_14452,N_15244);
and U15854 (N_15854,N_14635,N_15055);
or U15855 (N_15855,N_15205,N_15364);
nand U15856 (N_15856,N_15004,N_15263);
or U15857 (N_15857,N_15128,N_14571);
nor U15858 (N_15858,N_15130,N_14574);
or U15859 (N_15859,N_14785,N_14510);
and U15860 (N_15860,N_14823,N_15296);
xnor U15861 (N_15861,N_15391,N_14753);
nand U15862 (N_15862,N_15445,N_14485);
xnor U15863 (N_15863,N_15330,N_14949);
nand U15864 (N_15864,N_15454,N_14963);
xnor U15865 (N_15865,N_14555,N_14859);
or U15866 (N_15866,N_14502,N_15405);
nand U15867 (N_15867,N_14885,N_15457);
nor U15868 (N_15868,N_14683,N_14604);
and U15869 (N_15869,N_14918,N_15464);
and U15870 (N_15870,N_15242,N_14814);
nor U15871 (N_15871,N_14888,N_14576);
and U15872 (N_15872,N_14676,N_15421);
and U15873 (N_15873,N_15204,N_15550);
nand U15874 (N_15874,N_15338,N_14589);
and U15875 (N_15875,N_14520,N_15269);
nor U15876 (N_15876,N_14926,N_15565);
or U15877 (N_15877,N_15563,N_15385);
nand U15878 (N_15878,N_14737,N_14819);
nor U15879 (N_15879,N_14413,N_14818);
and U15880 (N_15880,N_15213,N_15079);
and U15881 (N_15881,N_15166,N_15018);
and U15882 (N_15882,N_15553,N_15331);
nand U15883 (N_15883,N_14613,N_14906);
nor U15884 (N_15884,N_15124,N_14972);
nor U15885 (N_15885,N_15253,N_15149);
nor U15886 (N_15886,N_15028,N_15089);
xnor U15887 (N_15887,N_14427,N_15333);
and U15888 (N_15888,N_14471,N_14714);
nor U15889 (N_15889,N_15499,N_14901);
and U15890 (N_15890,N_14602,N_14984);
and U15891 (N_15891,N_15428,N_15158);
nand U15892 (N_15892,N_15367,N_14762);
nor U15893 (N_15893,N_15260,N_15468);
nand U15894 (N_15894,N_15169,N_14789);
xnor U15895 (N_15895,N_14697,N_14575);
nor U15896 (N_15896,N_15093,N_14964);
nand U15897 (N_15897,N_15399,N_14940);
or U15898 (N_15898,N_15082,N_14423);
nor U15899 (N_15899,N_15558,N_14765);
xor U15900 (N_15900,N_15510,N_15078);
or U15901 (N_15901,N_14562,N_15332);
or U15902 (N_15902,N_14528,N_15334);
nand U15903 (N_15903,N_15365,N_14813);
xnor U15904 (N_15904,N_14493,N_14537);
nor U15905 (N_15905,N_15073,N_15120);
nand U15906 (N_15906,N_14774,N_15270);
nor U15907 (N_15907,N_15535,N_15407);
and U15908 (N_15908,N_15017,N_14838);
and U15909 (N_15909,N_14636,N_15074);
nor U15910 (N_15910,N_14736,N_14590);
or U15911 (N_15911,N_14491,N_14911);
and U15912 (N_15912,N_14797,N_15031);
or U15913 (N_15913,N_14690,N_14508);
and U15914 (N_15914,N_14702,N_14681);
xnor U15915 (N_15915,N_15157,N_15546);
or U15916 (N_15916,N_15441,N_14592);
nand U15917 (N_15917,N_14463,N_14750);
xor U15918 (N_15918,N_14549,N_14526);
nor U15919 (N_15919,N_15033,N_14833);
or U15920 (N_15920,N_14855,N_14428);
xnor U15921 (N_15921,N_15135,N_14815);
xnor U15922 (N_15922,N_15278,N_15307);
and U15923 (N_15923,N_15579,N_15395);
nor U15924 (N_15924,N_14748,N_14619);
and U15925 (N_15925,N_14771,N_14412);
and U15926 (N_15926,N_15326,N_14879);
or U15927 (N_15927,N_14687,N_15515);
xnor U15928 (N_15928,N_15403,N_15321);
nor U15929 (N_15929,N_14904,N_15112);
or U15930 (N_15930,N_15212,N_15107);
xnor U15931 (N_15931,N_15542,N_14956);
nand U15932 (N_15932,N_14677,N_14630);
nand U15933 (N_15933,N_15475,N_15459);
xor U15934 (N_15934,N_15151,N_15159);
or U15935 (N_15935,N_14989,N_14436);
nand U15936 (N_15936,N_15424,N_14611);
and U15937 (N_15937,N_14961,N_14482);
xor U15938 (N_15938,N_15193,N_15304);
nand U15939 (N_15939,N_14834,N_15560);
xor U15940 (N_15940,N_15433,N_14557);
nor U15941 (N_15941,N_15177,N_14498);
and U15942 (N_15942,N_14456,N_14965);
nor U15943 (N_15943,N_14409,N_14864);
xor U15944 (N_15944,N_14420,N_15543);
and U15945 (N_15945,N_14837,N_14970);
and U15946 (N_15946,N_15312,N_14487);
xnor U15947 (N_15947,N_15125,N_15344);
nor U15948 (N_15948,N_15328,N_15101);
xor U15949 (N_15949,N_14887,N_15174);
and U15950 (N_15950,N_15186,N_14600);
and U15951 (N_15951,N_15167,N_15285);
nor U15952 (N_15952,N_14856,N_15552);
nand U15953 (N_15953,N_15224,N_14793);
and U15954 (N_15954,N_15119,N_14927);
and U15955 (N_15955,N_15435,N_15202);
or U15956 (N_15956,N_15257,N_15021);
nand U15957 (N_15957,N_14933,N_15171);
or U15958 (N_15958,N_14798,N_15551);
and U15959 (N_15959,N_15431,N_14931);
xor U15960 (N_15960,N_15537,N_15027);
nor U15961 (N_15961,N_14874,N_15536);
or U15962 (N_15962,N_15261,N_15109);
xor U15963 (N_15963,N_14805,N_14988);
and U15964 (N_15964,N_14465,N_14775);
or U15965 (N_15965,N_15469,N_15415);
nor U15966 (N_15966,N_15160,N_14764);
and U15967 (N_15967,N_15179,N_15096);
nand U15968 (N_15968,N_15462,N_14679);
xor U15969 (N_15969,N_14500,N_15190);
and U15970 (N_15970,N_14925,N_14505);
and U15971 (N_15971,N_15533,N_15580);
xnor U15972 (N_15972,N_15175,N_15349);
nand U15973 (N_15973,N_15491,N_14632);
xnor U15974 (N_15974,N_14801,N_15049);
xor U15975 (N_15975,N_15488,N_15271);
or U15976 (N_15976,N_15502,N_14946);
nor U15977 (N_15977,N_14932,N_15482);
and U15978 (N_15978,N_15319,N_15318);
nand U15979 (N_15979,N_14792,N_15446);
nor U15980 (N_15980,N_15077,N_14850);
or U15981 (N_15981,N_14717,N_15097);
nand U15982 (N_15982,N_15046,N_15292);
nor U15983 (N_15983,N_14706,N_14854);
xor U15984 (N_15984,N_15479,N_15024);
xor U15985 (N_15985,N_15293,N_14820);
nor U15986 (N_15986,N_15225,N_15420);
and U15987 (N_15987,N_15199,N_14768);
nor U15988 (N_15988,N_15155,N_14664);
or U15989 (N_15989,N_14418,N_15042);
nand U15990 (N_15990,N_15458,N_14930);
nor U15991 (N_15991,N_14966,N_14494);
xor U15992 (N_15992,N_15373,N_15591);
nor U15993 (N_15993,N_14568,N_15188);
or U15994 (N_15994,N_15342,N_14626);
or U15995 (N_15995,N_15586,N_14566);
or U15996 (N_15996,N_15267,N_14691);
nand U15997 (N_15997,N_15419,N_14898);
nor U15998 (N_15998,N_14867,N_14916);
and U15999 (N_15999,N_14634,N_14699);
nand U16000 (N_16000,N_15528,N_15194);
nand U16001 (N_16001,N_14755,N_14843);
or U16002 (N_16002,N_15035,N_15059);
xnor U16003 (N_16003,N_14869,N_14745);
nand U16004 (N_16004,N_15008,N_14594);
and U16005 (N_16005,N_15248,N_15471);
or U16006 (N_16006,N_15509,N_15523);
nand U16007 (N_16007,N_14897,N_15234);
or U16008 (N_16008,N_14731,N_14694);
or U16009 (N_16009,N_15056,N_15453);
nor U16010 (N_16010,N_14606,N_14625);
or U16011 (N_16011,N_15571,N_14713);
nor U16012 (N_16012,N_15557,N_15298);
nand U16013 (N_16013,N_15087,N_14701);
and U16014 (N_16014,N_15116,N_15408);
or U16015 (N_16015,N_14665,N_15180);
nand U16016 (N_16016,N_15540,N_14653);
xor U16017 (N_16017,N_15503,N_15496);
or U16018 (N_16018,N_14993,N_15493);
xnor U16019 (N_16019,N_14637,N_15121);
or U16020 (N_16020,N_14572,N_14870);
and U16021 (N_16021,N_14579,N_15279);
nand U16022 (N_16022,N_14795,N_15376);
xnor U16023 (N_16023,N_14873,N_14831);
and U16024 (N_16024,N_15593,N_15337);
or U16025 (N_16025,N_15227,N_15195);
and U16026 (N_16026,N_15137,N_14563);
nor U16027 (N_16027,N_14863,N_14451);
or U16028 (N_16028,N_15361,N_14923);
nor U16029 (N_16029,N_15183,N_15080);
nor U16030 (N_16030,N_14490,N_15545);
or U16031 (N_16031,N_15438,N_15291);
and U16032 (N_16032,N_15470,N_15102);
or U16033 (N_16033,N_15525,N_15103);
nand U16034 (N_16034,N_14599,N_14998);
xnor U16035 (N_16035,N_15016,N_14968);
nor U16036 (N_16036,N_14719,N_14710);
or U16037 (N_16037,N_14685,N_14422);
and U16038 (N_16038,N_14440,N_15339);
nand U16039 (N_16039,N_15172,N_15476);
or U16040 (N_16040,N_15366,N_15280);
nor U16041 (N_16041,N_14723,N_14835);
and U16042 (N_16042,N_14928,N_15000);
nor U16043 (N_16043,N_15396,N_14875);
and U16044 (N_16044,N_15239,N_15379);
and U16045 (N_16045,N_14458,N_14514);
and U16046 (N_16046,N_15442,N_15492);
or U16047 (N_16047,N_14614,N_15129);
nor U16048 (N_16048,N_14554,N_15514);
nor U16049 (N_16049,N_14729,N_15075);
or U16050 (N_16050,N_15529,N_14659);
and U16051 (N_16051,N_14454,N_15484);
or U16052 (N_16052,N_14791,N_14844);
or U16053 (N_16053,N_15037,N_15473);
or U16054 (N_16054,N_14534,N_15564);
nor U16055 (N_16055,N_14470,N_14550);
nor U16056 (N_16056,N_14533,N_14861);
nor U16057 (N_16057,N_15495,N_14479);
nand U16058 (N_16058,N_15314,N_14919);
nand U16059 (N_16059,N_14934,N_15243);
nor U16060 (N_16060,N_15254,N_14426);
nand U16061 (N_16061,N_15143,N_15247);
nor U16062 (N_16062,N_15335,N_15481);
nand U16063 (N_16063,N_14531,N_15250);
or U16064 (N_16064,N_14624,N_15306);
or U16065 (N_16065,N_14751,N_14990);
xor U16066 (N_16066,N_14586,N_14703);
and U16067 (N_16067,N_14806,N_14547);
nand U16068 (N_16068,N_14570,N_14595);
nand U16069 (N_16069,N_14507,N_15411);
xor U16070 (N_16070,N_15086,N_15216);
xnor U16071 (N_16071,N_15091,N_15256);
nor U16072 (N_16072,N_14995,N_15374);
xnor U16073 (N_16073,N_14523,N_15584);
and U16074 (N_16074,N_14437,N_15141);
nor U16075 (N_16075,N_14591,N_14588);
nand U16076 (N_16076,N_14684,N_14766);
nand U16077 (N_16077,N_15070,N_15165);
xor U16078 (N_16078,N_15200,N_15276);
and U16079 (N_16079,N_15410,N_15034);
or U16080 (N_16080,N_14812,N_15117);
or U16081 (N_16081,N_15460,N_14804);
nor U16082 (N_16082,N_14513,N_14662);
xor U16083 (N_16083,N_14647,N_15067);
or U16084 (N_16084,N_15201,N_14638);
nor U16085 (N_16085,N_14680,N_15409);
or U16086 (N_16086,N_15010,N_15065);
or U16087 (N_16087,N_14829,N_14565);
and U16088 (N_16088,N_14969,N_15152);
nor U16089 (N_16089,N_14759,N_14878);
or U16090 (N_16090,N_15184,N_15516);
nor U16091 (N_16091,N_14593,N_15245);
nor U16092 (N_16092,N_14865,N_14596);
xor U16093 (N_16093,N_14817,N_14503);
and U16094 (N_16094,N_14744,N_14525);
or U16095 (N_16095,N_15599,N_15450);
nor U16096 (N_16096,N_14907,N_15108);
nor U16097 (N_16097,N_15168,N_14809);
nor U16098 (N_16098,N_14556,N_15106);
or U16099 (N_16099,N_14752,N_14585);
xor U16100 (N_16100,N_14912,N_15092);
or U16101 (N_16101,N_14616,N_15215);
xnor U16102 (N_16102,N_15310,N_15578);
and U16103 (N_16103,N_14406,N_14803);
and U16104 (N_16104,N_14649,N_14445);
nand U16105 (N_16105,N_14432,N_14738);
nand U16106 (N_16106,N_14446,N_15444);
and U16107 (N_16107,N_15572,N_14929);
nor U16108 (N_16108,N_14868,N_14544);
xnor U16109 (N_16109,N_14603,N_14608);
xnor U16110 (N_16110,N_14480,N_14464);
nor U16111 (N_16111,N_14417,N_14583);
nand U16112 (N_16112,N_15123,N_14705);
xor U16113 (N_16113,N_14698,N_15132);
xnor U16114 (N_16114,N_15222,N_14917);
xor U16115 (N_16115,N_14462,N_14734);
nor U16116 (N_16116,N_15474,N_14667);
nand U16117 (N_16117,N_14788,N_14955);
nand U16118 (N_16118,N_15053,N_14842);
nand U16119 (N_16119,N_15556,N_14558);
and U16120 (N_16120,N_15500,N_15275);
nand U16121 (N_16121,N_14866,N_15598);
or U16122 (N_16122,N_14876,N_15144);
nor U16123 (N_16123,N_14527,N_15099);
nor U16124 (N_16124,N_14781,N_14790);
or U16125 (N_16125,N_14678,N_15483);
xor U16126 (N_16126,N_14475,N_14512);
and U16127 (N_16127,N_14516,N_15397);
or U16128 (N_16128,N_15030,N_15068);
or U16129 (N_16129,N_14692,N_15272);
xor U16130 (N_16130,N_14495,N_15284);
or U16131 (N_16131,N_15187,N_15548);
nor U16132 (N_16132,N_14447,N_14605);
nor U16133 (N_16133,N_14826,N_15358);
xor U16134 (N_16134,N_15302,N_14476);
xnor U16135 (N_16135,N_15413,N_15131);
xor U16136 (N_16136,N_14836,N_15026);
xnor U16137 (N_16137,N_15534,N_15083);
xnor U16138 (N_16138,N_15081,N_15282);
and U16139 (N_16139,N_15038,N_15090);
xnor U16140 (N_16140,N_14552,N_14435);
xnor U16141 (N_16141,N_14663,N_14496);
xor U16142 (N_16142,N_15022,N_14724);
nor U16143 (N_16143,N_15532,N_15352);
and U16144 (N_16144,N_15567,N_15322);
and U16145 (N_16145,N_14401,N_14442);
and U16146 (N_16146,N_14958,N_14504);
and U16147 (N_16147,N_15025,N_15192);
nand U16148 (N_16148,N_14438,N_14954);
nand U16149 (N_16149,N_14541,N_15327);
and U16150 (N_16150,N_15486,N_14707);
xnor U16151 (N_16151,N_14641,N_15047);
xnor U16152 (N_16152,N_14473,N_14821);
and U16153 (N_16153,N_15512,N_15219);
or U16154 (N_16154,N_14943,N_14434);
or U16155 (N_16155,N_15489,N_15596);
nor U16156 (N_16156,N_14675,N_15570);
nor U16157 (N_16157,N_14615,N_14796);
or U16158 (N_16158,N_15426,N_15539);
nor U16159 (N_16159,N_15146,N_14488);
nor U16160 (N_16160,N_15544,N_14658);
xor U16161 (N_16161,N_14400,N_14783);
nor U16162 (N_16162,N_15581,N_14643);
nand U16163 (N_16163,N_15429,N_14976);
nand U16164 (N_16164,N_15218,N_14407);
and U16165 (N_16165,N_14862,N_15388);
nor U16166 (N_16166,N_14741,N_15023);
nand U16167 (N_16167,N_15436,N_14872);
and U16168 (N_16168,N_14760,N_14983);
nor U16169 (N_16169,N_15178,N_14841);
xor U16170 (N_16170,N_15019,N_15233);
and U16171 (N_16171,N_15052,N_15113);
xor U16172 (N_16172,N_15198,N_14535);
nor U16173 (N_16173,N_14433,N_14414);
nor U16174 (N_16174,N_14506,N_15506);
nand U16175 (N_16175,N_15490,N_14708);
and U16176 (N_16176,N_14472,N_15217);
nand U16177 (N_16177,N_15044,N_15573);
nand U16178 (N_16178,N_15273,N_15440);
nand U16179 (N_16179,N_15595,N_15162);
or U16180 (N_16180,N_15226,N_14743);
xnor U16181 (N_16181,N_14524,N_14824);
nand U16182 (N_16182,N_14900,N_14799);
nand U16183 (N_16183,N_14517,N_15480);
and U16184 (N_16184,N_15393,N_14776);
or U16185 (N_16185,N_14839,N_14695);
nand U16186 (N_16186,N_14825,N_15357);
xnor U16187 (N_16187,N_14425,N_14952);
or U16188 (N_16188,N_14627,N_15347);
nor U16189 (N_16189,N_15588,N_15305);
and U16190 (N_16190,N_14560,N_14935);
and U16191 (N_16191,N_14924,N_14770);
or U16192 (N_16192,N_14808,N_14457);
xor U16193 (N_16193,N_15387,N_15575);
nor U16194 (N_16194,N_14725,N_15311);
and U16195 (N_16195,N_15384,N_14499);
and U16196 (N_16196,N_15554,N_14405);
nand U16197 (N_16197,N_15582,N_15562);
and U16198 (N_16198,N_15530,N_15360);
or U16199 (N_16199,N_14489,N_15003);
xor U16200 (N_16200,N_14503,N_14568);
and U16201 (N_16201,N_15456,N_15177);
and U16202 (N_16202,N_14576,N_15052);
or U16203 (N_16203,N_14888,N_14660);
nor U16204 (N_16204,N_14959,N_14641);
or U16205 (N_16205,N_14657,N_14507);
and U16206 (N_16206,N_14574,N_14427);
and U16207 (N_16207,N_14701,N_14497);
nor U16208 (N_16208,N_15554,N_14880);
and U16209 (N_16209,N_15184,N_15014);
nand U16210 (N_16210,N_14952,N_14879);
xor U16211 (N_16211,N_15464,N_15336);
xnor U16212 (N_16212,N_14819,N_15340);
nand U16213 (N_16213,N_15310,N_15526);
or U16214 (N_16214,N_14477,N_14678);
or U16215 (N_16215,N_15514,N_14639);
or U16216 (N_16216,N_14982,N_15334);
or U16217 (N_16217,N_15458,N_15264);
xor U16218 (N_16218,N_15201,N_15513);
and U16219 (N_16219,N_15181,N_14578);
or U16220 (N_16220,N_14906,N_14465);
or U16221 (N_16221,N_14888,N_15511);
nand U16222 (N_16222,N_15145,N_15390);
xor U16223 (N_16223,N_14451,N_15112);
xor U16224 (N_16224,N_15187,N_14514);
or U16225 (N_16225,N_15065,N_15550);
or U16226 (N_16226,N_14821,N_15345);
or U16227 (N_16227,N_15573,N_14724);
and U16228 (N_16228,N_14590,N_15425);
or U16229 (N_16229,N_14423,N_15139);
or U16230 (N_16230,N_15120,N_14701);
nor U16231 (N_16231,N_14463,N_14609);
nand U16232 (N_16232,N_14583,N_15146);
nand U16233 (N_16233,N_14452,N_14868);
nand U16234 (N_16234,N_14651,N_14636);
nand U16235 (N_16235,N_14573,N_14808);
nand U16236 (N_16236,N_15173,N_15575);
nor U16237 (N_16237,N_15225,N_15473);
nor U16238 (N_16238,N_15515,N_15404);
nand U16239 (N_16239,N_15202,N_14821);
nor U16240 (N_16240,N_15366,N_14722);
or U16241 (N_16241,N_15497,N_14619);
nand U16242 (N_16242,N_14642,N_14408);
and U16243 (N_16243,N_15568,N_15072);
nor U16244 (N_16244,N_14433,N_15395);
or U16245 (N_16245,N_15387,N_14411);
xnor U16246 (N_16246,N_15478,N_14666);
or U16247 (N_16247,N_14564,N_15322);
and U16248 (N_16248,N_14805,N_14716);
xor U16249 (N_16249,N_14950,N_15234);
and U16250 (N_16250,N_15558,N_15507);
or U16251 (N_16251,N_15281,N_14745);
and U16252 (N_16252,N_15527,N_14809);
xnor U16253 (N_16253,N_15452,N_15097);
and U16254 (N_16254,N_15356,N_15071);
or U16255 (N_16255,N_15013,N_14917);
nor U16256 (N_16256,N_14404,N_14868);
nand U16257 (N_16257,N_15202,N_14630);
or U16258 (N_16258,N_15490,N_15028);
and U16259 (N_16259,N_15233,N_15544);
or U16260 (N_16260,N_15079,N_15259);
and U16261 (N_16261,N_15294,N_14605);
and U16262 (N_16262,N_15088,N_15302);
nor U16263 (N_16263,N_15256,N_15383);
nor U16264 (N_16264,N_14771,N_15494);
nor U16265 (N_16265,N_15326,N_15388);
xnor U16266 (N_16266,N_15092,N_15316);
or U16267 (N_16267,N_15279,N_14664);
nand U16268 (N_16268,N_14896,N_14986);
or U16269 (N_16269,N_15103,N_15467);
nand U16270 (N_16270,N_15091,N_14652);
xor U16271 (N_16271,N_14627,N_14520);
nand U16272 (N_16272,N_15298,N_15515);
or U16273 (N_16273,N_15097,N_14806);
or U16274 (N_16274,N_15335,N_15447);
nand U16275 (N_16275,N_15529,N_14906);
xor U16276 (N_16276,N_15144,N_15007);
nand U16277 (N_16277,N_14662,N_14532);
and U16278 (N_16278,N_15011,N_14513);
and U16279 (N_16279,N_14583,N_15396);
or U16280 (N_16280,N_14585,N_14503);
and U16281 (N_16281,N_14659,N_14910);
nand U16282 (N_16282,N_15487,N_15208);
and U16283 (N_16283,N_14596,N_14679);
nand U16284 (N_16284,N_15209,N_14873);
nor U16285 (N_16285,N_15201,N_14846);
or U16286 (N_16286,N_15115,N_14430);
xnor U16287 (N_16287,N_15111,N_15396);
and U16288 (N_16288,N_14434,N_14658);
nor U16289 (N_16289,N_15594,N_15068);
nor U16290 (N_16290,N_14532,N_14489);
xor U16291 (N_16291,N_14457,N_14886);
nand U16292 (N_16292,N_14924,N_14573);
nand U16293 (N_16293,N_15352,N_14900);
xnor U16294 (N_16294,N_14681,N_15116);
nand U16295 (N_16295,N_14582,N_14413);
nor U16296 (N_16296,N_15028,N_14526);
xor U16297 (N_16297,N_15133,N_15304);
or U16298 (N_16298,N_15055,N_14960);
xor U16299 (N_16299,N_15323,N_15533);
nand U16300 (N_16300,N_14944,N_14768);
nand U16301 (N_16301,N_14731,N_15183);
nand U16302 (N_16302,N_14878,N_15021);
and U16303 (N_16303,N_15471,N_14915);
and U16304 (N_16304,N_14915,N_14964);
nand U16305 (N_16305,N_15322,N_15484);
xor U16306 (N_16306,N_15188,N_15332);
nand U16307 (N_16307,N_15333,N_14635);
and U16308 (N_16308,N_14576,N_14511);
nand U16309 (N_16309,N_15492,N_14774);
nand U16310 (N_16310,N_15430,N_14824);
nor U16311 (N_16311,N_14698,N_15245);
or U16312 (N_16312,N_15549,N_15384);
xnor U16313 (N_16313,N_15230,N_14402);
nand U16314 (N_16314,N_14483,N_15125);
nor U16315 (N_16315,N_15261,N_15047);
and U16316 (N_16316,N_15465,N_15186);
or U16317 (N_16317,N_15446,N_15151);
and U16318 (N_16318,N_14587,N_15040);
nor U16319 (N_16319,N_15070,N_14823);
or U16320 (N_16320,N_14904,N_15067);
nand U16321 (N_16321,N_14914,N_15079);
xor U16322 (N_16322,N_14548,N_15276);
nand U16323 (N_16323,N_14624,N_14837);
nor U16324 (N_16324,N_14473,N_14556);
nand U16325 (N_16325,N_14895,N_14859);
and U16326 (N_16326,N_15536,N_14678);
xor U16327 (N_16327,N_15173,N_14484);
xnor U16328 (N_16328,N_14589,N_15175);
and U16329 (N_16329,N_15011,N_14856);
and U16330 (N_16330,N_14996,N_15324);
nor U16331 (N_16331,N_14566,N_15176);
nor U16332 (N_16332,N_14825,N_14486);
nor U16333 (N_16333,N_14762,N_14564);
nor U16334 (N_16334,N_14982,N_14547);
xor U16335 (N_16335,N_15167,N_15544);
xnor U16336 (N_16336,N_15417,N_15144);
nor U16337 (N_16337,N_15559,N_15304);
nor U16338 (N_16338,N_15544,N_15469);
and U16339 (N_16339,N_15452,N_15201);
and U16340 (N_16340,N_15557,N_14676);
nand U16341 (N_16341,N_14476,N_15000);
xor U16342 (N_16342,N_15194,N_14747);
or U16343 (N_16343,N_15390,N_15242);
nor U16344 (N_16344,N_15560,N_14622);
nand U16345 (N_16345,N_14488,N_14611);
or U16346 (N_16346,N_14848,N_14882);
nand U16347 (N_16347,N_14558,N_15522);
xnor U16348 (N_16348,N_15214,N_15467);
xnor U16349 (N_16349,N_14500,N_15529);
nor U16350 (N_16350,N_14908,N_14713);
nor U16351 (N_16351,N_14621,N_14947);
and U16352 (N_16352,N_15190,N_14410);
xnor U16353 (N_16353,N_14645,N_14509);
and U16354 (N_16354,N_14931,N_14886);
or U16355 (N_16355,N_15592,N_14877);
nand U16356 (N_16356,N_15326,N_14606);
nand U16357 (N_16357,N_14967,N_14514);
nor U16358 (N_16358,N_15179,N_15579);
nor U16359 (N_16359,N_15011,N_14732);
nand U16360 (N_16360,N_15378,N_15066);
or U16361 (N_16361,N_14704,N_15398);
xnor U16362 (N_16362,N_14652,N_14506);
and U16363 (N_16363,N_14922,N_14416);
nor U16364 (N_16364,N_15065,N_14864);
nor U16365 (N_16365,N_15004,N_14449);
nor U16366 (N_16366,N_15468,N_15415);
nand U16367 (N_16367,N_15263,N_15235);
or U16368 (N_16368,N_15015,N_14831);
nand U16369 (N_16369,N_15120,N_14812);
xnor U16370 (N_16370,N_15005,N_14976);
or U16371 (N_16371,N_14932,N_14812);
xnor U16372 (N_16372,N_14918,N_15427);
or U16373 (N_16373,N_14948,N_14647);
nand U16374 (N_16374,N_14479,N_15017);
nor U16375 (N_16375,N_15353,N_14515);
nand U16376 (N_16376,N_14932,N_15144);
xnor U16377 (N_16377,N_15498,N_15041);
nor U16378 (N_16378,N_14832,N_15056);
nand U16379 (N_16379,N_14818,N_15134);
or U16380 (N_16380,N_14463,N_14782);
and U16381 (N_16381,N_15284,N_14550);
xor U16382 (N_16382,N_14658,N_15134);
and U16383 (N_16383,N_15255,N_14772);
xnor U16384 (N_16384,N_14439,N_14917);
or U16385 (N_16385,N_15043,N_15408);
and U16386 (N_16386,N_14904,N_14445);
nor U16387 (N_16387,N_15015,N_14655);
or U16388 (N_16388,N_14450,N_15310);
and U16389 (N_16389,N_14600,N_14960);
xnor U16390 (N_16390,N_15191,N_15248);
and U16391 (N_16391,N_14652,N_15582);
nand U16392 (N_16392,N_14939,N_14819);
and U16393 (N_16393,N_15427,N_14978);
and U16394 (N_16394,N_14831,N_14449);
and U16395 (N_16395,N_15243,N_14878);
nor U16396 (N_16396,N_15451,N_14745);
nor U16397 (N_16397,N_15447,N_15194);
xnor U16398 (N_16398,N_14573,N_14582);
xnor U16399 (N_16399,N_15373,N_15233);
and U16400 (N_16400,N_14566,N_14461);
and U16401 (N_16401,N_14532,N_14482);
nor U16402 (N_16402,N_15322,N_14694);
nor U16403 (N_16403,N_15335,N_14568);
and U16404 (N_16404,N_14940,N_14712);
or U16405 (N_16405,N_15360,N_14790);
nand U16406 (N_16406,N_15473,N_14468);
xnor U16407 (N_16407,N_15206,N_14588);
nor U16408 (N_16408,N_14816,N_14840);
nor U16409 (N_16409,N_15231,N_15274);
or U16410 (N_16410,N_15523,N_14797);
nand U16411 (N_16411,N_15116,N_14752);
or U16412 (N_16412,N_15215,N_14430);
or U16413 (N_16413,N_14970,N_15165);
xnor U16414 (N_16414,N_14664,N_14794);
nor U16415 (N_16415,N_14796,N_14535);
and U16416 (N_16416,N_14748,N_14848);
xor U16417 (N_16417,N_15236,N_14892);
or U16418 (N_16418,N_14814,N_15285);
or U16419 (N_16419,N_14965,N_15155);
or U16420 (N_16420,N_15204,N_14400);
nor U16421 (N_16421,N_14411,N_14815);
or U16422 (N_16422,N_14455,N_15046);
or U16423 (N_16423,N_15435,N_14527);
and U16424 (N_16424,N_15555,N_14738);
or U16425 (N_16425,N_14533,N_15446);
and U16426 (N_16426,N_15357,N_14637);
or U16427 (N_16427,N_15207,N_15444);
and U16428 (N_16428,N_15470,N_15334);
nor U16429 (N_16429,N_15352,N_14761);
and U16430 (N_16430,N_15344,N_14666);
xor U16431 (N_16431,N_14668,N_14645);
nor U16432 (N_16432,N_14478,N_15399);
and U16433 (N_16433,N_14714,N_15213);
nor U16434 (N_16434,N_15110,N_15305);
nand U16435 (N_16435,N_15380,N_14992);
and U16436 (N_16436,N_14473,N_14653);
nand U16437 (N_16437,N_14861,N_15177);
nand U16438 (N_16438,N_15227,N_15499);
and U16439 (N_16439,N_15261,N_14895);
nand U16440 (N_16440,N_14951,N_15544);
xor U16441 (N_16441,N_14703,N_14602);
xor U16442 (N_16442,N_15104,N_15165);
nand U16443 (N_16443,N_14488,N_15454);
nand U16444 (N_16444,N_15331,N_14449);
nor U16445 (N_16445,N_14481,N_14561);
xor U16446 (N_16446,N_14475,N_15568);
xor U16447 (N_16447,N_14960,N_14549);
xnor U16448 (N_16448,N_14981,N_15252);
nand U16449 (N_16449,N_14761,N_14727);
xor U16450 (N_16450,N_14950,N_15341);
nor U16451 (N_16451,N_14598,N_14654);
and U16452 (N_16452,N_15427,N_14747);
or U16453 (N_16453,N_15517,N_15071);
and U16454 (N_16454,N_14441,N_14656);
or U16455 (N_16455,N_14794,N_15151);
nand U16456 (N_16456,N_15568,N_15457);
nand U16457 (N_16457,N_14558,N_14442);
nor U16458 (N_16458,N_15423,N_14738);
or U16459 (N_16459,N_15325,N_15207);
nor U16460 (N_16460,N_14573,N_15263);
and U16461 (N_16461,N_15107,N_14540);
nand U16462 (N_16462,N_14739,N_14974);
nor U16463 (N_16463,N_14821,N_14764);
and U16464 (N_16464,N_14484,N_14485);
nor U16465 (N_16465,N_15344,N_15079);
nand U16466 (N_16466,N_15171,N_15272);
nor U16467 (N_16467,N_14597,N_14758);
nand U16468 (N_16468,N_15494,N_15342);
nand U16469 (N_16469,N_14833,N_15197);
nand U16470 (N_16470,N_15438,N_15214);
or U16471 (N_16471,N_14658,N_14740);
and U16472 (N_16472,N_15160,N_15376);
or U16473 (N_16473,N_15175,N_15417);
nand U16474 (N_16474,N_14977,N_15344);
nor U16475 (N_16475,N_14581,N_15282);
and U16476 (N_16476,N_15135,N_15039);
nand U16477 (N_16477,N_14625,N_15077);
nand U16478 (N_16478,N_14437,N_15454);
and U16479 (N_16479,N_14401,N_15278);
nand U16480 (N_16480,N_15144,N_14975);
nand U16481 (N_16481,N_14999,N_15518);
nor U16482 (N_16482,N_15338,N_14933);
and U16483 (N_16483,N_15447,N_14530);
xnor U16484 (N_16484,N_15302,N_15107);
nor U16485 (N_16485,N_15307,N_14553);
and U16486 (N_16486,N_15018,N_15435);
xnor U16487 (N_16487,N_15546,N_14416);
nor U16488 (N_16488,N_14901,N_14913);
nor U16489 (N_16489,N_14989,N_14680);
nor U16490 (N_16490,N_14978,N_14996);
or U16491 (N_16491,N_15492,N_15449);
nor U16492 (N_16492,N_14492,N_15589);
and U16493 (N_16493,N_14543,N_14964);
or U16494 (N_16494,N_14450,N_15217);
or U16495 (N_16495,N_14969,N_15561);
xor U16496 (N_16496,N_14713,N_15241);
or U16497 (N_16497,N_15539,N_14648);
and U16498 (N_16498,N_15413,N_15450);
nand U16499 (N_16499,N_14808,N_15534);
nand U16500 (N_16500,N_14557,N_14875);
xnor U16501 (N_16501,N_14425,N_14764);
nor U16502 (N_16502,N_15049,N_15533);
nor U16503 (N_16503,N_15593,N_14798);
nor U16504 (N_16504,N_14537,N_15226);
nor U16505 (N_16505,N_14863,N_15016);
xor U16506 (N_16506,N_14772,N_15232);
or U16507 (N_16507,N_14537,N_15096);
and U16508 (N_16508,N_14558,N_15008);
xor U16509 (N_16509,N_14579,N_15257);
xor U16510 (N_16510,N_15458,N_14470);
nand U16511 (N_16511,N_14514,N_14979);
or U16512 (N_16512,N_15516,N_15091);
or U16513 (N_16513,N_15293,N_14961);
or U16514 (N_16514,N_15096,N_15401);
nor U16515 (N_16515,N_15264,N_15202);
nand U16516 (N_16516,N_15474,N_15542);
xnor U16517 (N_16517,N_15177,N_14865);
xnor U16518 (N_16518,N_15147,N_14846);
xor U16519 (N_16519,N_14807,N_14417);
nor U16520 (N_16520,N_15509,N_15274);
or U16521 (N_16521,N_14417,N_14644);
and U16522 (N_16522,N_15011,N_15261);
nand U16523 (N_16523,N_15281,N_14948);
or U16524 (N_16524,N_14958,N_15163);
nor U16525 (N_16525,N_14963,N_15139);
nand U16526 (N_16526,N_15454,N_15031);
xor U16527 (N_16527,N_14474,N_15539);
or U16528 (N_16528,N_14573,N_15216);
and U16529 (N_16529,N_15212,N_14961);
or U16530 (N_16530,N_14782,N_15023);
and U16531 (N_16531,N_15381,N_15451);
xnor U16532 (N_16532,N_14659,N_15233);
and U16533 (N_16533,N_14551,N_14548);
nor U16534 (N_16534,N_14786,N_15258);
nand U16535 (N_16535,N_15454,N_15279);
xnor U16536 (N_16536,N_15528,N_15448);
nor U16537 (N_16537,N_14571,N_15297);
or U16538 (N_16538,N_14843,N_15084);
xnor U16539 (N_16539,N_14406,N_15000);
and U16540 (N_16540,N_15299,N_15510);
and U16541 (N_16541,N_15299,N_15422);
or U16542 (N_16542,N_14694,N_14499);
xor U16543 (N_16543,N_14945,N_15437);
nand U16544 (N_16544,N_14536,N_15256);
nand U16545 (N_16545,N_14762,N_14551);
or U16546 (N_16546,N_14844,N_14780);
nor U16547 (N_16547,N_15533,N_14725);
xor U16548 (N_16548,N_14589,N_14841);
and U16549 (N_16549,N_15064,N_15302);
or U16550 (N_16550,N_14947,N_14761);
nand U16551 (N_16551,N_15102,N_14801);
nor U16552 (N_16552,N_15054,N_15135);
xnor U16553 (N_16553,N_15138,N_15448);
xor U16554 (N_16554,N_15205,N_14418);
and U16555 (N_16555,N_15359,N_14694);
xnor U16556 (N_16556,N_14677,N_14896);
nand U16557 (N_16557,N_15005,N_14779);
nand U16558 (N_16558,N_14921,N_14474);
nand U16559 (N_16559,N_15051,N_15369);
nand U16560 (N_16560,N_14496,N_14747);
xor U16561 (N_16561,N_15022,N_14538);
and U16562 (N_16562,N_14561,N_15409);
or U16563 (N_16563,N_14424,N_15471);
xnor U16564 (N_16564,N_15330,N_15162);
nor U16565 (N_16565,N_15327,N_14559);
nor U16566 (N_16566,N_15599,N_15459);
nor U16567 (N_16567,N_15002,N_14826);
or U16568 (N_16568,N_15103,N_14736);
and U16569 (N_16569,N_15156,N_15038);
xor U16570 (N_16570,N_15291,N_15367);
nor U16571 (N_16571,N_15360,N_15528);
xnor U16572 (N_16572,N_15494,N_15146);
nor U16573 (N_16573,N_15435,N_14487);
nor U16574 (N_16574,N_14811,N_15241);
nor U16575 (N_16575,N_14479,N_15431);
or U16576 (N_16576,N_14747,N_14741);
and U16577 (N_16577,N_14775,N_14912);
nand U16578 (N_16578,N_14492,N_14586);
and U16579 (N_16579,N_15093,N_14965);
nor U16580 (N_16580,N_15188,N_15029);
and U16581 (N_16581,N_15083,N_15072);
nand U16582 (N_16582,N_14788,N_14904);
and U16583 (N_16583,N_14439,N_15247);
nand U16584 (N_16584,N_15031,N_15323);
and U16585 (N_16585,N_15597,N_14573);
and U16586 (N_16586,N_14461,N_15254);
nand U16587 (N_16587,N_15332,N_14466);
xnor U16588 (N_16588,N_15103,N_14922);
nand U16589 (N_16589,N_15361,N_14981);
nand U16590 (N_16590,N_15282,N_14911);
xor U16591 (N_16591,N_15458,N_15125);
and U16592 (N_16592,N_14952,N_15098);
and U16593 (N_16593,N_15345,N_15252);
or U16594 (N_16594,N_15125,N_14818);
or U16595 (N_16595,N_15086,N_14943);
and U16596 (N_16596,N_15392,N_14816);
nor U16597 (N_16597,N_14682,N_15136);
or U16598 (N_16598,N_14846,N_15584);
and U16599 (N_16599,N_14725,N_14434);
nand U16600 (N_16600,N_14536,N_14540);
or U16601 (N_16601,N_14717,N_14902);
nand U16602 (N_16602,N_15208,N_14925);
nor U16603 (N_16603,N_14964,N_15435);
and U16604 (N_16604,N_15363,N_14531);
xnor U16605 (N_16605,N_15405,N_14493);
xor U16606 (N_16606,N_15240,N_15285);
or U16607 (N_16607,N_14886,N_15243);
and U16608 (N_16608,N_15399,N_15339);
nor U16609 (N_16609,N_14423,N_14963);
or U16610 (N_16610,N_14528,N_14901);
or U16611 (N_16611,N_14886,N_14920);
nand U16612 (N_16612,N_15581,N_14630);
or U16613 (N_16613,N_15394,N_15502);
nor U16614 (N_16614,N_14603,N_14747);
nor U16615 (N_16615,N_14804,N_14565);
or U16616 (N_16616,N_15032,N_15537);
nor U16617 (N_16617,N_14692,N_15396);
and U16618 (N_16618,N_14502,N_14929);
xnor U16619 (N_16619,N_15485,N_15051);
xnor U16620 (N_16620,N_14844,N_15098);
nand U16621 (N_16621,N_14603,N_15522);
or U16622 (N_16622,N_14700,N_15366);
and U16623 (N_16623,N_14817,N_15244);
and U16624 (N_16624,N_14609,N_14623);
or U16625 (N_16625,N_14581,N_15054);
and U16626 (N_16626,N_14731,N_15538);
nand U16627 (N_16627,N_14929,N_15466);
or U16628 (N_16628,N_15409,N_14644);
and U16629 (N_16629,N_14788,N_14471);
and U16630 (N_16630,N_14736,N_15138);
xor U16631 (N_16631,N_15185,N_14536);
nand U16632 (N_16632,N_14944,N_15085);
nand U16633 (N_16633,N_15540,N_15431);
and U16634 (N_16634,N_14564,N_15158);
xnor U16635 (N_16635,N_15036,N_15235);
xnor U16636 (N_16636,N_15408,N_15060);
xnor U16637 (N_16637,N_15279,N_14887);
and U16638 (N_16638,N_15309,N_14538);
and U16639 (N_16639,N_15416,N_15429);
and U16640 (N_16640,N_15515,N_14665);
nand U16641 (N_16641,N_14655,N_14437);
xnor U16642 (N_16642,N_14855,N_14931);
and U16643 (N_16643,N_14634,N_15072);
or U16644 (N_16644,N_14725,N_15564);
and U16645 (N_16645,N_15140,N_14662);
or U16646 (N_16646,N_15347,N_15297);
nand U16647 (N_16647,N_15340,N_14876);
nand U16648 (N_16648,N_14577,N_14922);
and U16649 (N_16649,N_15395,N_14496);
nor U16650 (N_16650,N_14643,N_15367);
or U16651 (N_16651,N_14566,N_14839);
xnor U16652 (N_16652,N_15003,N_14572);
xnor U16653 (N_16653,N_14679,N_14936);
nand U16654 (N_16654,N_15365,N_14413);
or U16655 (N_16655,N_14498,N_14619);
nor U16656 (N_16656,N_15172,N_15197);
xnor U16657 (N_16657,N_14946,N_15285);
and U16658 (N_16658,N_14484,N_14836);
xor U16659 (N_16659,N_15180,N_14411);
or U16660 (N_16660,N_14668,N_15257);
and U16661 (N_16661,N_15125,N_14487);
nand U16662 (N_16662,N_14551,N_15322);
and U16663 (N_16663,N_15418,N_14623);
xnor U16664 (N_16664,N_14870,N_14899);
and U16665 (N_16665,N_14863,N_15511);
and U16666 (N_16666,N_14757,N_14550);
nand U16667 (N_16667,N_15151,N_15238);
nand U16668 (N_16668,N_15467,N_15515);
and U16669 (N_16669,N_15448,N_15435);
nand U16670 (N_16670,N_14915,N_15534);
nand U16671 (N_16671,N_15457,N_15343);
or U16672 (N_16672,N_14442,N_15483);
xnor U16673 (N_16673,N_15337,N_14445);
nand U16674 (N_16674,N_14909,N_14622);
nand U16675 (N_16675,N_15443,N_15181);
and U16676 (N_16676,N_15391,N_14930);
xnor U16677 (N_16677,N_15290,N_14402);
or U16678 (N_16678,N_14509,N_15334);
and U16679 (N_16679,N_14688,N_14537);
xor U16680 (N_16680,N_15302,N_15453);
nand U16681 (N_16681,N_14798,N_15554);
xor U16682 (N_16682,N_14754,N_15452);
nor U16683 (N_16683,N_15537,N_14483);
nand U16684 (N_16684,N_15369,N_14976);
xnor U16685 (N_16685,N_15119,N_14636);
xor U16686 (N_16686,N_15472,N_14537);
xor U16687 (N_16687,N_15099,N_14674);
xnor U16688 (N_16688,N_15574,N_15569);
xor U16689 (N_16689,N_14720,N_15418);
and U16690 (N_16690,N_15346,N_14912);
or U16691 (N_16691,N_15568,N_15244);
and U16692 (N_16692,N_14627,N_14729);
xnor U16693 (N_16693,N_14981,N_15028);
or U16694 (N_16694,N_15206,N_14576);
nand U16695 (N_16695,N_14505,N_14947);
or U16696 (N_16696,N_14577,N_15163);
or U16697 (N_16697,N_15360,N_14664);
nor U16698 (N_16698,N_14653,N_14597);
xor U16699 (N_16699,N_14510,N_15266);
xnor U16700 (N_16700,N_15583,N_14941);
nor U16701 (N_16701,N_15330,N_15410);
xnor U16702 (N_16702,N_14773,N_15356);
and U16703 (N_16703,N_14635,N_15362);
and U16704 (N_16704,N_15431,N_14796);
xnor U16705 (N_16705,N_15067,N_14533);
or U16706 (N_16706,N_15125,N_14736);
xor U16707 (N_16707,N_14965,N_14974);
xor U16708 (N_16708,N_14595,N_15019);
or U16709 (N_16709,N_14730,N_14504);
or U16710 (N_16710,N_14735,N_14547);
xnor U16711 (N_16711,N_15362,N_15246);
xor U16712 (N_16712,N_15432,N_15157);
xor U16713 (N_16713,N_14832,N_14547);
and U16714 (N_16714,N_15410,N_15215);
xnor U16715 (N_16715,N_14604,N_14812);
nor U16716 (N_16716,N_14829,N_15514);
xor U16717 (N_16717,N_15351,N_15553);
xnor U16718 (N_16718,N_14810,N_15462);
or U16719 (N_16719,N_15127,N_14528);
nor U16720 (N_16720,N_15452,N_14599);
and U16721 (N_16721,N_15050,N_15081);
xnor U16722 (N_16722,N_14769,N_15497);
and U16723 (N_16723,N_15152,N_14724);
xor U16724 (N_16724,N_15557,N_14501);
or U16725 (N_16725,N_15535,N_15034);
and U16726 (N_16726,N_14527,N_15111);
and U16727 (N_16727,N_15305,N_15395);
xnor U16728 (N_16728,N_15430,N_15298);
nor U16729 (N_16729,N_15263,N_15593);
xor U16730 (N_16730,N_14771,N_15147);
nor U16731 (N_16731,N_14439,N_15515);
nor U16732 (N_16732,N_15133,N_14406);
nor U16733 (N_16733,N_14407,N_15500);
nand U16734 (N_16734,N_15283,N_15483);
and U16735 (N_16735,N_14658,N_15173);
nor U16736 (N_16736,N_15403,N_14456);
nand U16737 (N_16737,N_15125,N_15004);
nor U16738 (N_16738,N_14905,N_14472);
and U16739 (N_16739,N_15500,N_14881);
nand U16740 (N_16740,N_14917,N_15232);
nor U16741 (N_16741,N_14988,N_14730);
xor U16742 (N_16742,N_14895,N_15148);
and U16743 (N_16743,N_15408,N_15097);
and U16744 (N_16744,N_15473,N_15057);
nand U16745 (N_16745,N_15265,N_15157);
nand U16746 (N_16746,N_14547,N_15391);
xor U16747 (N_16747,N_14927,N_14866);
xor U16748 (N_16748,N_15221,N_15081);
or U16749 (N_16749,N_15510,N_14881);
xor U16750 (N_16750,N_15376,N_14872);
xnor U16751 (N_16751,N_14997,N_15529);
nor U16752 (N_16752,N_14928,N_14641);
and U16753 (N_16753,N_14789,N_14683);
nor U16754 (N_16754,N_15175,N_14835);
xnor U16755 (N_16755,N_15321,N_14817);
xor U16756 (N_16756,N_14442,N_14699);
nand U16757 (N_16757,N_15481,N_15381);
nor U16758 (N_16758,N_15243,N_15351);
nor U16759 (N_16759,N_15462,N_14612);
xor U16760 (N_16760,N_15050,N_14502);
and U16761 (N_16761,N_14819,N_15541);
nor U16762 (N_16762,N_15246,N_15134);
nor U16763 (N_16763,N_14493,N_15296);
nor U16764 (N_16764,N_15509,N_14729);
xnor U16765 (N_16765,N_14608,N_15573);
or U16766 (N_16766,N_15526,N_14507);
xor U16767 (N_16767,N_15319,N_15178);
xor U16768 (N_16768,N_15355,N_15445);
xor U16769 (N_16769,N_14554,N_15220);
xor U16770 (N_16770,N_15455,N_14627);
or U16771 (N_16771,N_14624,N_14553);
nand U16772 (N_16772,N_15154,N_14459);
and U16773 (N_16773,N_15132,N_15562);
nor U16774 (N_16774,N_15352,N_15462);
and U16775 (N_16775,N_14589,N_14928);
or U16776 (N_16776,N_15224,N_15398);
and U16777 (N_16777,N_15169,N_14823);
nor U16778 (N_16778,N_15384,N_15238);
xor U16779 (N_16779,N_14588,N_15311);
nand U16780 (N_16780,N_14783,N_15366);
nand U16781 (N_16781,N_15282,N_14403);
nand U16782 (N_16782,N_14702,N_15171);
xnor U16783 (N_16783,N_14737,N_15534);
xor U16784 (N_16784,N_15479,N_15264);
nor U16785 (N_16785,N_14444,N_14899);
xnor U16786 (N_16786,N_15541,N_15264);
nand U16787 (N_16787,N_15171,N_15050);
and U16788 (N_16788,N_15124,N_15263);
xnor U16789 (N_16789,N_14576,N_14697);
or U16790 (N_16790,N_14477,N_14798);
nor U16791 (N_16791,N_14889,N_14600);
and U16792 (N_16792,N_15064,N_14632);
and U16793 (N_16793,N_14549,N_14636);
or U16794 (N_16794,N_14571,N_14755);
nand U16795 (N_16795,N_15583,N_15406);
xor U16796 (N_16796,N_14402,N_15530);
or U16797 (N_16797,N_15208,N_14480);
nand U16798 (N_16798,N_14556,N_14926);
nor U16799 (N_16799,N_14693,N_15399);
xnor U16800 (N_16800,N_15739,N_16151);
nand U16801 (N_16801,N_16583,N_15775);
nand U16802 (N_16802,N_16341,N_15997);
xnor U16803 (N_16803,N_16548,N_15655);
or U16804 (N_16804,N_15870,N_16142);
or U16805 (N_16805,N_16263,N_16131);
nand U16806 (N_16806,N_16010,N_15981);
or U16807 (N_16807,N_16179,N_16650);
or U16808 (N_16808,N_16289,N_15924);
nand U16809 (N_16809,N_15783,N_15601);
xor U16810 (N_16810,N_16273,N_16016);
or U16811 (N_16811,N_16314,N_16296);
or U16812 (N_16812,N_16398,N_15709);
nand U16813 (N_16813,N_15905,N_16505);
nand U16814 (N_16814,N_15842,N_15898);
and U16815 (N_16815,N_16632,N_16237);
nand U16816 (N_16816,N_16007,N_16261);
xnor U16817 (N_16817,N_16733,N_15988);
nor U16818 (N_16818,N_15718,N_16385);
xnor U16819 (N_16819,N_15611,N_16712);
nand U16820 (N_16820,N_16722,N_16424);
or U16821 (N_16821,N_16628,N_16725);
or U16822 (N_16822,N_15944,N_15770);
or U16823 (N_16823,N_16365,N_16232);
nor U16824 (N_16824,N_15614,N_16464);
nor U16825 (N_16825,N_16105,N_15874);
or U16826 (N_16826,N_16550,N_15803);
nor U16827 (N_16827,N_16213,N_15619);
nand U16828 (N_16828,N_15694,N_16114);
nor U16829 (N_16829,N_16406,N_16559);
or U16830 (N_16830,N_16674,N_16594);
and U16831 (N_16831,N_16283,N_16259);
xnor U16832 (N_16832,N_16160,N_16715);
nor U16833 (N_16833,N_16667,N_16122);
nor U16834 (N_16834,N_16293,N_15663);
or U16835 (N_16835,N_15707,N_15604);
nand U16836 (N_16836,N_15699,N_15983);
and U16837 (N_16837,N_15875,N_16230);
or U16838 (N_16838,N_16768,N_15762);
or U16839 (N_16839,N_16564,N_16692);
and U16840 (N_16840,N_15706,N_15795);
nor U16841 (N_16841,N_15643,N_16547);
and U16842 (N_16842,N_16311,N_15705);
and U16843 (N_16843,N_16689,N_15765);
nand U16844 (N_16844,N_16757,N_16143);
xor U16845 (N_16845,N_16136,N_16645);
and U16846 (N_16846,N_15646,N_15832);
or U16847 (N_16847,N_16255,N_15794);
nor U16848 (N_16848,N_16130,N_16728);
or U16849 (N_16849,N_16219,N_16767);
or U16850 (N_16850,N_16523,N_16287);
nor U16851 (N_16851,N_16388,N_15681);
xor U16852 (N_16852,N_16716,N_16599);
and U16853 (N_16853,N_15800,N_16745);
nor U16854 (N_16854,N_16379,N_16642);
nand U16855 (N_16855,N_15841,N_16119);
or U16856 (N_16856,N_16171,N_16521);
or U16857 (N_16857,N_16752,N_15847);
xnor U16858 (N_16858,N_16481,N_16309);
and U16859 (N_16859,N_16449,N_16648);
and U16860 (N_16860,N_15731,N_16605);
xor U16861 (N_16861,N_16029,N_15786);
nor U16862 (N_16862,N_16125,N_16666);
nor U16863 (N_16863,N_16206,N_16661);
or U16864 (N_16864,N_16258,N_16421);
and U16865 (N_16865,N_16133,N_15833);
xor U16866 (N_16866,N_16101,N_16377);
nor U16867 (N_16867,N_15941,N_15986);
or U16868 (N_16868,N_15761,N_15909);
and U16869 (N_16869,N_15600,N_15647);
nand U16870 (N_16870,N_16770,N_15928);
and U16871 (N_16871,N_16476,N_16773);
nand U16872 (N_16872,N_15767,N_16185);
nand U16873 (N_16873,N_15695,N_15797);
xor U16874 (N_16874,N_16199,N_16473);
or U16875 (N_16875,N_16520,N_16163);
nor U16876 (N_16876,N_16695,N_16221);
or U16877 (N_16877,N_15827,N_16228);
xnor U16878 (N_16878,N_16418,N_16531);
xnor U16879 (N_16879,N_15916,N_15808);
nand U16880 (N_16880,N_16134,N_16582);
nor U16881 (N_16881,N_15645,N_16732);
nor U16882 (N_16882,N_16623,N_16747);
xnor U16883 (N_16883,N_16404,N_16681);
xnor U16884 (N_16884,N_16382,N_15908);
or U16885 (N_16885,N_15782,N_15697);
xor U16886 (N_16886,N_16647,N_16074);
xnor U16887 (N_16887,N_16205,N_16274);
nand U16888 (N_16888,N_16708,N_15877);
and U16889 (N_16889,N_15653,N_16413);
nor U16890 (N_16890,N_16447,N_16102);
and U16891 (N_16891,N_15968,N_15788);
xnor U16892 (N_16892,N_16215,N_16718);
and U16893 (N_16893,N_16031,N_16499);
nor U16894 (N_16894,N_16729,N_16015);
or U16895 (N_16895,N_16412,N_16753);
or U16896 (N_16896,N_16442,N_16491);
xnor U16897 (N_16897,N_15667,N_16756);
nand U16898 (N_16898,N_16239,N_15603);
and U16899 (N_16899,N_15954,N_16127);
nor U16900 (N_16900,N_16370,N_15781);
and U16901 (N_16901,N_16658,N_15719);
nand U16902 (N_16902,N_15720,N_16357);
or U16903 (N_16903,N_16693,N_15756);
or U16904 (N_16904,N_16774,N_16478);
and U16905 (N_16905,N_16177,N_15766);
nand U16906 (N_16906,N_16012,N_16400);
nor U16907 (N_16907,N_16369,N_15885);
nand U16908 (N_16908,N_16158,N_16188);
nor U16909 (N_16909,N_16124,N_16036);
nor U16910 (N_16910,N_15972,N_15689);
nand U16911 (N_16911,N_16192,N_16282);
nor U16912 (N_16912,N_16086,N_15650);
nor U16913 (N_16913,N_16711,N_15796);
or U16914 (N_16914,N_16005,N_16256);
nor U16915 (N_16915,N_15973,N_15878);
and U16916 (N_16916,N_15675,N_16709);
or U16917 (N_16917,N_16619,N_16678);
or U16918 (N_16918,N_16765,N_16037);
nand U16919 (N_16919,N_16760,N_16578);
and U16920 (N_16920,N_16563,N_16116);
nand U16921 (N_16921,N_16669,N_16480);
or U16922 (N_16922,N_16522,N_16401);
xnor U16923 (N_16923,N_16097,N_16194);
nand U16924 (N_16924,N_15880,N_16062);
and U16925 (N_16925,N_16764,N_16749);
or U16926 (N_16926,N_16065,N_16509);
or U16927 (N_16927,N_15982,N_15914);
and U16928 (N_16928,N_15670,N_15886);
nor U16929 (N_16929,N_16109,N_16190);
nand U16930 (N_16930,N_16662,N_16717);
nor U16931 (N_16931,N_16025,N_16214);
nand U16932 (N_16932,N_15763,N_16141);
or U16933 (N_16933,N_16387,N_16434);
nor U16934 (N_16934,N_16300,N_16120);
nand U16935 (N_16935,N_16467,N_16275);
nand U16936 (N_16936,N_16796,N_16006);
xnor U16937 (N_16937,N_16513,N_16461);
nand U16938 (N_16938,N_16140,N_15974);
nand U16939 (N_16939,N_16448,N_15657);
and U16940 (N_16940,N_16793,N_15958);
nor U16941 (N_16941,N_16003,N_16304);
nand U16942 (N_16942,N_16542,N_15708);
nor U16943 (N_16943,N_15659,N_16574);
xnor U16944 (N_16944,N_15753,N_15679);
xnor U16945 (N_16945,N_16466,N_16298);
and U16946 (N_16946,N_16649,N_16425);
xor U16947 (N_16947,N_15764,N_16337);
and U16948 (N_16948,N_15624,N_16734);
nor U16949 (N_16949,N_16349,N_16494);
nand U16950 (N_16950,N_16433,N_15957);
xor U16951 (N_16951,N_16581,N_15779);
or U16952 (N_16952,N_16640,N_15821);
xnor U16953 (N_16953,N_15602,N_16530);
nor U16954 (N_16954,N_15934,N_16254);
nand U16955 (N_16955,N_16541,N_15899);
or U16956 (N_16956,N_15834,N_16034);
nor U16957 (N_16957,N_16705,N_15823);
nor U16958 (N_16958,N_15950,N_15726);
xor U16959 (N_16959,N_16570,N_16148);
and U16960 (N_16960,N_16685,N_16617);
or U16961 (N_16961,N_15854,N_16637);
or U16962 (N_16962,N_15838,N_16556);
and U16963 (N_16963,N_16367,N_16361);
and U16964 (N_16964,N_16222,N_16291);
nand U16965 (N_16965,N_15966,N_16393);
and U16966 (N_16966,N_15949,N_16310);
nor U16967 (N_16967,N_16061,N_16603);
nand U16968 (N_16968,N_15936,N_16202);
nand U16969 (N_16969,N_16313,N_15677);
xor U16970 (N_16970,N_16048,N_16286);
and U16971 (N_16971,N_16799,N_15751);
and U16972 (N_16972,N_15960,N_16532);
or U16973 (N_16973,N_15747,N_16653);
and U16974 (N_16974,N_16346,N_16394);
xnor U16975 (N_16975,N_16477,N_16458);
xnor U16976 (N_16976,N_16052,N_15933);
nor U16977 (N_16977,N_16064,N_16279);
and U16978 (N_16978,N_16557,N_15926);
xor U16979 (N_16979,N_16055,N_16225);
nand U16980 (N_16980,N_16396,N_16149);
and U16981 (N_16981,N_16660,N_15774);
or U16982 (N_16982,N_16409,N_15776);
nand U16983 (N_16983,N_16246,N_15861);
nand U16984 (N_16984,N_16782,N_16137);
xor U16985 (N_16985,N_15771,N_16788);
or U16986 (N_16986,N_16233,N_16781);
xnor U16987 (N_16987,N_15656,N_15809);
or U16988 (N_16988,N_16132,N_16735);
xnor U16989 (N_16989,N_16696,N_16184);
nand U16990 (N_16990,N_16615,N_16312);
xnor U16991 (N_16991,N_16634,N_16766);
nand U16992 (N_16992,N_16100,N_16288);
xnor U16993 (N_16993,N_15868,N_15851);
or U16994 (N_16994,N_15666,N_16284);
nor U16995 (N_16995,N_16572,N_15883);
xor U16996 (N_16996,N_15664,N_15849);
nand U16997 (N_16997,N_16511,N_16697);
nand U16998 (N_16998,N_15822,N_15637);
nor U16999 (N_16999,N_16479,N_16067);
xnor U17000 (N_17000,N_16644,N_16054);
xnor U17001 (N_17001,N_16414,N_16486);
xor U17002 (N_17002,N_16621,N_15992);
and U17003 (N_17003,N_15642,N_16076);
nand U17004 (N_17004,N_16032,N_16568);
nor U17005 (N_17005,N_15638,N_16000);
or U17006 (N_17006,N_16704,N_16195);
and U17007 (N_17007,N_16294,N_16707);
nand U17008 (N_17008,N_16014,N_16673);
xnor U17009 (N_17009,N_16320,N_16209);
nor U17010 (N_17010,N_16220,N_16022);
or U17011 (N_17011,N_15711,N_16210);
and U17012 (N_17012,N_16422,N_16450);
and U17013 (N_17013,N_15790,N_15943);
xor U17014 (N_17014,N_15716,N_16775);
nor U17015 (N_17015,N_16165,N_16383);
nand U17016 (N_17016,N_16651,N_15722);
nor U17017 (N_17017,N_15829,N_16200);
nand U17018 (N_17018,N_16405,N_16252);
or U17019 (N_17019,N_16562,N_15636);
or U17020 (N_17020,N_16169,N_15621);
nor U17021 (N_17021,N_16178,N_16786);
xor U17022 (N_17022,N_16295,N_16162);
nor U17023 (N_17023,N_16157,N_16703);
xnor U17024 (N_17024,N_15693,N_15629);
xnor U17025 (N_17025,N_16240,N_16071);
and U17026 (N_17026,N_16262,N_16506);
or U17027 (N_17027,N_16248,N_16595);
or U17028 (N_17028,N_15912,N_16526);
nor U17029 (N_17029,N_15999,N_16411);
or U17030 (N_17030,N_15831,N_16187);
nor U17031 (N_17031,N_16281,N_16610);
or U17032 (N_17032,N_15930,N_15613);
nor U17033 (N_17033,N_16602,N_15938);
or U17034 (N_17034,N_16677,N_16380);
nor U17035 (N_17035,N_16153,N_16445);
xor U17036 (N_17036,N_16739,N_16664);
or U17037 (N_17037,N_16710,N_16079);
nand U17038 (N_17038,N_16207,N_16198);
and U17039 (N_17039,N_15961,N_16440);
nand U17040 (N_17040,N_16107,N_16553);
xnor U17041 (N_17041,N_16652,N_16303);
xor U17042 (N_17042,N_16569,N_16290);
and U17043 (N_17043,N_15661,N_16196);
nor U17044 (N_17044,N_16686,N_15696);
nor U17045 (N_17045,N_15824,N_16112);
nor U17046 (N_17046,N_15702,N_15871);
nand U17047 (N_17047,N_16073,N_16609);
and U17048 (N_17048,N_16211,N_16001);
nand U17049 (N_17049,N_16358,N_16611);
nor U17050 (N_17050,N_16575,N_16302);
or U17051 (N_17051,N_16597,N_16191);
nor U17052 (N_17052,N_16687,N_16508);
nor U17053 (N_17053,N_16543,N_15820);
xnor U17054 (N_17054,N_15959,N_16484);
or U17055 (N_17055,N_16354,N_15625);
or U17056 (N_17056,N_15819,N_16571);
and U17057 (N_17057,N_15952,N_15806);
or U17058 (N_17058,N_16245,N_16088);
nor U17059 (N_17059,N_16671,N_16567);
nor U17060 (N_17060,N_16111,N_16672);
nor U17061 (N_17061,N_16278,N_16417);
nand U17062 (N_17062,N_15852,N_15740);
nor U17063 (N_17063,N_15994,N_16573);
or U17064 (N_17064,N_15985,N_16251);
nor U17065 (N_17065,N_16189,N_16343);
nor U17066 (N_17066,N_16454,N_15758);
or U17067 (N_17067,N_16145,N_15615);
and U17068 (N_17068,N_15630,N_16777);
nor U17069 (N_17069,N_16453,N_16545);
xor U17070 (N_17070,N_16468,N_16604);
nand U17071 (N_17071,N_16181,N_16035);
and U17072 (N_17072,N_16203,N_16011);
nand U17073 (N_17073,N_15906,N_16436);
xor U17074 (N_17074,N_16502,N_16472);
and U17075 (N_17075,N_15859,N_15889);
nand U17076 (N_17076,N_15990,N_16495);
or U17077 (N_17077,N_15759,N_16627);
and U17078 (N_17078,N_15684,N_15978);
nand U17079 (N_17079,N_15757,N_16730);
or U17080 (N_17080,N_16063,N_15680);
nand U17081 (N_17081,N_15752,N_16738);
or U17082 (N_17082,N_16056,N_15791);
xor U17083 (N_17083,N_16144,N_15872);
and U17084 (N_17084,N_16330,N_16399);
nand U17085 (N_17085,N_16460,N_16030);
nor U17086 (N_17086,N_16235,N_16498);
nor U17087 (N_17087,N_16694,N_16675);
xnor U17088 (N_17088,N_16362,N_15850);
xor U17089 (N_17089,N_15866,N_16253);
nand U17090 (N_17090,N_15727,N_15641);
nand U17091 (N_17091,N_16426,N_16561);
nand U17092 (N_17092,N_15815,N_15772);
or U17093 (N_17093,N_16376,N_15724);
and U17094 (N_17094,N_15682,N_16748);
or U17095 (N_17095,N_16699,N_15732);
nor U17096 (N_17096,N_16208,N_16438);
and U17097 (N_17097,N_16350,N_16135);
xnor U17098 (N_17098,N_16075,N_15807);
and U17099 (N_17099,N_16082,N_16635);
xor U17100 (N_17100,N_16093,N_15967);
xnor U17101 (N_17101,N_16155,N_16792);
and U17102 (N_17102,N_15890,N_15913);
nand U17103 (N_17103,N_16483,N_16322);
or U17104 (N_17104,N_16051,N_16363);
nor U17105 (N_17105,N_16428,N_15730);
xor U17106 (N_17106,N_16643,N_16586);
nand U17107 (N_17107,N_16250,N_16356);
nand U17108 (N_17108,N_15755,N_15712);
nor U17109 (N_17109,N_16243,N_16164);
nor U17110 (N_17110,N_16264,N_15998);
or U17111 (N_17111,N_15789,N_16272);
xor U17112 (N_17112,N_16338,N_16415);
xnor U17113 (N_17113,N_15749,N_16299);
nor U17114 (N_17114,N_16057,N_16497);
nand U17115 (N_17115,N_16613,N_15704);
nor U17116 (N_17116,N_16044,N_16193);
or U17117 (N_17117,N_15895,N_16359);
nand U17118 (N_17118,N_16701,N_16375);
xor U17119 (N_17119,N_15685,N_16395);
and U17120 (N_17120,N_15953,N_16683);
or U17121 (N_17121,N_15939,N_16596);
nor U17122 (N_17122,N_16049,N_16368);
and U17123 (N_17123,N_16512,N_16386);
nand U17124 (N_17124,N_16021,N_16684);
and U17125 (N_17125,N_16761,N_16126);
or U17126 (N_17126,N_16390,N_16167);
or U17127 (N_17127,N_16474,N_16465);
nor U17128 (N_17128,N_16762,N_15887);
and U17129 (N_17129,N_15669,N_16534);
nand U17130 (N_17130,N_15900,N_15743);
nor U17131 (N_17131,N_15723,N_16423);
nand U17132 (N_17132,N_16790,N_16384);
or U17133 (N_17133,N_15626,N_16047);
xor U17134 (N_17134,N_15947,N_16241);
and U17135 (N_17135,N_16089,N_15911);
or U17136 (N_17136,N_15768,N_15901);
and U17137 (N_17137,N_16459,N_16771);
or U17138 (N_17138,N_15654,N_15927);
xor U17139 (N_17139,N_16721,N_16355);
nand U17140 (N_17140,N_16754,N_15951);
nand U17141 (N_17141,N_16759,N_16551);
or U17142 (N_17142,N_15744,N_16340);
nor U17143 (N_17143,N_15632,N_16173);
xnor U17144 (N_17144,N_16755,N_15867);
nor U17145 (N_17145,N_16576,N_16389);
nor U17146 (N_17146,N_16094,N_16630);
nand U17147 (N_17147,N_15893,N_16514);
and U17148 (N_17148,N_16580,N_16794);
and U17149 (N_17149,N_16746,N_16045);
nor U17150 (N_17150,N_15814,N_16629);
nand U17151 (N_17151,N_16432,N_15920);
nor U17152 (N_17152,N_16091,N_16231);
xnor U17153 (N_17153,N_16680,N_15942);
nand U17154 (N_17154,N_16769,N_15844);
xnor U17155 (N_17155,N_16280,N_16364);
xnor U17156 (N_17156,N_16216,N_16028);
nor U17157 (N_17157,N_15692,N_15760);
nand U17158 (N_17158,N_15811,N_15640);
nand U17159 (N_17159,N_16663,N_15634);
nand U17160 (N_17160,N_16333,N_16698);
or U17161 (N_17161,N_15837,N_15660);
nor U17162 (N_17162,N_15818,N_16229);
nor U17163 (N_17163,N_16443,N_16352);
nand U17164 (N_17164,N_16566,N_16429);
or U17165 (N_17165,N_16702,N_16517);
and U17166 (N_17166,N_15826,N_16457);
xnor U17167 (N_17167,N_15616,N_16081);
nor U17168 (N_17168,N_16342,N_16763);
or U17169 (N_17169,N_16469,N_16285);
nand U17170 (N_17170,N_16587,N_15773);
nor U17171 (N_17171,N_15649,N_15792);
or U17172 (N_17172,N_15750,N_16668);
and U17173 (N_17173,N_16223,N_16268);
nand U17174 (N_17174,N_16138,N_15922);
and U17175 (N_17175,N_15633,N_16737);
xnor U17176 (N_17176,N_16482,N_15839);
nand U17177 (N_17177,N_16560,N_16544);
or U17178 (N_17178,N_16475,N_16204);
and U17179 (N_17179,N_16470,N_15793);
xnor U17180 (N_17180,N_15891,N_15698);
nor U17181 (N_17181,N_16183,N_16437);
nand U17182 (N_17182,N_16638,N_16106);
nor U17183 (N_17183,N_15665,N_15946);
or U17184 (N_17184,N_15658,N_16040);
xnor U17185 (N_17185,N_16787,N_16128);
or U17186 (N_17186,N_16226,N_16758);
and U17187 (N_17187,N_16507,N_16374);
nand U17188 (N_17188,N_15907,N_15945);
nand U17189 (N_17189,N_16224,N_15923);
xor U17190 (N_17190,N_15962,N_16121);
xor U17191 (N_17191,N_16345,N_16740);
nand U17192 (N_17192,N_16026,N_16182);
and U17193 (N_17193,N_16515,N_15987);
or U17194 (N_17194,N_16257,N_16113);
and U17195 (N_17195,N_16176,N_16403);
and U17196 (N_17196,N_15862,N_16778);
and U17197 (N_17197,N_15855,N_15713);
xnor U17198 (N_17198,N_16315,N_16622);
and U17199 (N_17199,N_16351,N_15873);
and U17200 (N_17200,N_16555,N_15607);
xnor U17201 (N_17201,N_16462,N_15892);
and U17202 (N_17202,N_16227,N_16714);
nor U17203 (N_17203,N_16123,N_15863);
or U17204 (N_17204,N_15688,N_15628);
and U17205 (N_17205,N_15802,N_16641);
nor U17206 (N_17206,N_16439,N_16490);
xor U17207 (N_17207,N_16744,N_15620);
nand U17208 (N_17208,N_16277,N_16174);
and U17209 (N_17209,N_16419,N_16552);
nand U17210 (N_17210,N_15948,N_16318);
nand U17211 (N_17211,N_15989,N_15672);
xor U17212 (N_17212,N_15686,N_16307);
xor U17213 (N_17213,N_15976,N_15980);
xnor U17214 (N_17214,N_16736,N_15879);
and U17215 (N_17215,N_16452,N_16301);
nand U17216 (N_17216,N_16485,N_16727);
nand U17217 (N_17217,N_16046,N_15921);
nand U17218 (N_17218,N_15700,N_16008);
nand U17219 (N_17219,N_15996,N_15780);
or U17220 (N_17220,N_15639,N_16618);
or U17221 (N_17221,N_15652,N_16270);
xnor U17222 (N_17222,N_16489,N_15882);
or U17223 (N_17223,N_15622,N_16540);
xnor U17224 (N_17224,N_16620,N_16070);
nor U17225 (N_17225,N_15671,N_16724);
and U17226 (N_17226,N_16095,N_15965);
nand U17227 (N_17227,N_15857,N_16271);
nor U17228 (N_17228,N_16039,N_15674);
and U17229 (N_17229,N_16050,N_16041);
xor U17230 (N_17230,N_16017,N_16083);
xor U17231 (N_17231,N_16679,N_15612);
or U17232 (N_17232,N_16772,N_16516);
or U17233 (N_17233,N_16719,N_16463);
nand U17234 (N_17234,N_16317,N_16150);
and U17235 (N_17235,N_15623,N_16146);
nor U17236 (N_17236,N_16348,N_16068);
nor U17237 (N_17237,N_15840,N_16161);
and U17238 (N_17238,N_16528,N_16159);
nor U17239 (N_17239,N_15631,N_16579);
and U17240 (N_17240,N_15701,N_15728);
nor U17241 (N_17241,N_16323,N_16612);
nand U17242 (N_17242,N_16538,N_16713);
and U17243 (N_17243,N_16780,N_15737);
or U17244 (N_17244,N_16218,N_16510);
or U17245 (N_17245,N_15617,N_15846);
or U17246 (N_17246,N_16529,N_16392);
xnor U17247 (N_17247,N_16108,N_16098);
and U17248 (N_17248,N_16750,N_16002);
and U17249 (N_17249,N_16503,N_16043);
or U17250 (N_17250,N_15673,N_16328);
nand U17251 (N_17251,N_15865,N_16493);
nand U17252 (N_17252,N_16776,N_16535);
xor U17253 (N_17253,N_16496,N_16360);
nand U17254 (N_17254,N_16332,N_16269);
and U17255 (N_17255,N_16410,N_16166);
nand U17256 (N_17256,N_15777,N_15746);
nor U17257 (N_17257,N_16616,N_15937);
nor U17258 (N_17258,N_15676,N_16156);
and U17259 (N_17259,N_16455,N_16584);
and U17260 (N_17260,N_16327,N_15799);
and U17261 (N_17261,N_16416,N_15856);
and U17262 (N_17262,N_16785,N_16518);
nor U17263 (N_17263,N_16319,N_15940);
nand U17264 (N_17264,N_16297,N_15644);
nand U17265 (N_17265,N_15969,N_15609);
or U17266 (N_17266,N_16607,N_16598);
xnor U17267 (N_17267,N_15816,N_16670);
nand U17268 (N_17268,N_15817,N_16519);
nand U17269 (N_17269,N_16731,N_16266);
or U17270 (N_17270,N_16691,N_16069);
and U17271 (N_17271,N_15741,N_15919);
xnor U17272 (N_17272,N_16391,N_15825);
or U17273 (N_17273,N_16018,N_15931);
or U17274 (N_17274,N_15714,N_15888);
and U17275 (N_17275,N_16741,N_16625);
or U17276 (N_17276,N_15910,N_16308);
xnor U17277 (N_17277,N_16080,N_15860);
xnor U17278 (N_17278,N_16633,N_16329);
nor U17279 (N_17279,N_16353,N_16038);
and U17280 (N_17280,N_16451,N_16639);
xnor U17281 (N_17281,N_16608,N_15869);
xor U17282 (N_17282,N_16152,N_16795);
or U17283 (N_17283,N_15836,N_16092);
or U17284 (N_17284,N_16659,N_16554);
and U17285 (N_17285,N_16058,N_15984);
nor U17286 (N_17286,N_15835,N_16078);
nand U17287 (N_17287,N_16614,N_15683);
nor U17288 (N_17288,N_15687,N_16537);
nor U17289 (N_17289,N_15991,N_15894);
nand U17290 (N_17290,N_15668,N_16217);
xor U17291 (N_17291,N_16084,N_15956);
and U17292 (N_17292,N_16726,N_15858);
nor U17293 (N_17293,N_16316,N_16129);
and U17294 (N_17294,N_16441,N_15902);
xor U17295 (N_17295,N_15610,N_15917);
or U17296 (N_17296,N_16456,N_16558);
or U17297 (N_17297,N_15735,N_15662);
and U17298 (N_17298,N_15691,N_16238);
xnor U17299 (N_17299,N_16372,N_15918);
xnor U17300 (N_17300,N_16751,N_16276);
or U17301 (N_17301,N_16381,N_16743);
nand U17302 (N_17302,N_16626,N_15715);
and U17303 (N_17303,N_16631,N_16706);
nand U17304 (N_17304,N_15678,N_16201);
and U17305 (N_17305,N_16791,N_16600);
xor U17306 (N_17306,N_16407,N_16117);
nand U17307 (N_17307,N_16234,N_16427);
and U17308 (N_17308,N_16103,N_16096);
nor U17309 (N_17309,N_16072,N_15805);
nor U17310 (N_17310,N_16019,N_15925);
nor U17311 (N_17311,N_15975,N_15804);
and U17312 (N_17312,N_16784,N_15995);
nor U17313 (N_17313,N_15864,N_16665);
nor U17314 (N_17314,N_16085,N_15848);
xor U17315 (N_17315,N_16260,N_15963);
xnor U17316 (N_17316,N_16335,N_16066);
nand U17317 (N_17317,N_15742,N_16249);
or U17318 (N_17318,N_16004,N_15729);
nand U17319 (N_17319,N_16588,N_15785);
nor U17320 (N_17320,N_16624,N_15784);
and U17321 (N_17321,N_16657,N_16536);
and U17322 (N_17322,N_16186,N_15745);
or U17323 (N_17323,N_16060,N_16306);
and U17324 (N_17324,N_16592,N_15738);
nor U17325 (N_17325,N_16446,N_15903);
and U17326 (N_17326,N_16789,N_16042);
and U17327 (N_17327,N_15787,N_16525);
xnor U17328 (N_17328,N_16504,N_16435);
nor U17329 (N_17329,N_15884,N_15798);
xnor U17330 (N_17330,N_15845,N_15648);
and U17331 (N_17331,N_16053,N_16646);
xnor U17332 (N_17332,N_16471,N_16334);
or U17333 (N_17333,N_15977,N_16797);
nor U17334 (N_17334,N_16378,N_16154);
or U17335 (N_17335,N_16676,N_15690);
xnor U17336 (N_17336,N_15876,N_15843);
nor U17337 (N_17337,N_16589,N_15721);
and U17338 (N_17338,N_16344,N_16347);
xnor U17339 (N_17339,N_15810,N_16524);
nand U17340 (N_17340,N_15881,N_16527);
xor U17341 (N_17341,N_16321,N_16655);
or U17342 (N_17342,N_16533,N_16723);
nand U17343 (N_17343,N_16212,N_16324);
nor U17344 (N_17344,N_16371,N_16024);
nand U17345 (N_17345,N_16577,N_16549);
nand U17346 (N_17346,N_16366,N_16009);
xor U17347 (N_17347,N_16326,N_15717);
xor U17348 (N_17348,N_16488,N_16180);
or U17349 (N_17349,N_15964,N_16170);
or U17350 (N_17350,N_15734,N_16090);
nand U17351 (N_17351,N_16267,N_16242);
or U17352 (N_17352,N_16139,N_16033);
xnor U17353 (N_17353,N_16601,N_15897);
or U17354 (N_17354,N_16027,N_15830);
or U17355 (N_17355,N_16500,N_16197);
nand U17356 (N_17356,N_16373,N_16336);
nand U17357 (N_17357,N_16420,N_15932);
or U17358 (N_17358,N_16431,N_16236);
nand U17359 (N_17359,N_16244,N_15904);
or U17360 (N_17360,N_15853,N_16172);
or U17361 (N_17361,N_16402,N_15618);
nand U17362 (N_17362,N_15736,N_15935);
xnor U17363 (N_17363,N_16087,N_15748);
and U17364 (N_17364,N_16305,N_15955);
nor U17365 (N_17365,N_15651,N_16585);
nor U17366 (N_17366,N_16168,N_16487);
nand U17367 (N_17367,N_15929,N_15725);
nand U17368 (N_17368,N_16339,N_15608);
or U17369 (N_17369,N_15754,N_15828);
nand U17370 (N_17370,N_15801,N_16700);
nand U17371 (N_17371,N_16636,N_16606);
nand U17372 (N_17372,N_15769,N_15703);
or U17373 (N_17373,N_15915,N_15993);
nor U17374 (N_17374,N_15778,N_16325);
xor U17375 (N_17375,N_16408,N_16265);
nand U17376 (N_17376,N_16742,N_15733);
nand U17377 (N_17377,N_16720,N_15979);
nor U17378 (N_17378,N_16656,N_16331);
nand U17379 (N_17379,N_16013,N_15971);
nand U17380 (N_17380,N_15627,N_16247);
nand U17381 (N_17381,N_16059,N_16175);
nor U17382 (N_17382,N_16104,N_15635);
nand U17383 (N_17383,N_16397,N_16688);
or U17384 (N_17384,N_15813,N_16492);
nand U17385 (N_17385,N_15606,N_16539);
or U17386 (N_17386,N_16292,N_16590);
and U17387 (N_17387,N_16147,N_16779);
nor U17388 (N_17388,N_16020,N_16077);
nor U17389 (N_17389,N_15812,N_16798);
nor U17390 (N_17390,N_16593,N_16430);
and U17391 (N_17391,N_15896,N_16099);
nand U17392 (N_17392,N_16654,N_16110);
nor U17393 (N_17393,N_16023,N_16591);
nand U17394 (N_17394,N_16682,N_16783);
or U17395 (N_17395,N_16444,N_15710);
and U17396 (N_17396,N_16690,N_15970);
xnor U17397 (N_17397,N_16118,N_16115);
nor U17398 (N_17398,N_16565,N_15605);
nor U17399 (N_17399,N_16546,N_16501);
xnor U17400 (N_17400,N_15856,N_16113);
or U17401 (N_17401,N_15884,N_15611);
or U17402 (N_17402,N_16131,N_16469);
or U17403 (N_17403,N_16710,N_15786);
and U17404 (N_17404,N_15616,N_15754);
or U17405 (N_17405,N_16427,N_16403);
or U17406 (N_17406,N_16142,N_15611);
or U17407 (N_17407,N_16281,N_16306);
and U17408 (N_17408,N_15955,N_16726);
or U17409 (N_17409,N_15875,N_16036);
and U17410 (N_17410,N_16097,N_16014);
nand U17411 (N_17411,N_16217,N_16319);
and U17412 (N_17412,N_15984,N_16485);
nor U17413 (N_17413,N_16422,N_15635);
or U17414 (N_17414,N_16675,N_15656);
and U17415 (N_17415,N_16213,N_16175);
xnor U17416 (N_17416,N_16414,N_16495);
nand U17417 (N_17417,N_16788,N_15864);
xor U17418 (N_17418,N_16753,N_16193);
nand U17419 (N_17419,N_16649,N_16139);
nand U17420 (N_17420,N_16479,N_16374);
xor U17421 (N_17421,N_16064,N_16744);
or U17422 (N_17422,N_16660,N_16288);
and U17423 (N_17423,N_16518,N_15936);
nor U17424 (N_17424,N_16722,N_16032);
or U17425 (N_17425,N_16610,N_16464);
xor U17426 (N_17426,N_16019,N_16031);
xor U17427 (N_17427,N_16688,N_16459);
xnor U17428 (N_17428,N_15829,N_16602);
nor U17429 (N_17429,N_16065,N_16433);
and U17430 (N_17430,N_16558,N_16622);
and U17431 (N_17431,N_15874,N_16035);
and U17432 (N_17432,N_16208,N_16534);
nand U17433 (N_17433,N_15883,N_16458);
or U17434 (N_17434,N_15797,N_16586);
nand U17435 (N_17435,N_15636,N_16294);
xor U17436 (N_17436,N_16744,N_15751);
xor U17437 (N_17437,N_16117,N_16082);
and U17438 (N_17438,N_15926,N_15808);
or U17439 (N_17439,N_15649,N_16050);
xor U17440 (N_17440,N_16314,N_16640);
xor U17441 (N_17441,N_15792,N_16409);
nand U17442 (N_17442,N_15816,N_15934);
or U17443 (N_17443,N_15893,N_16586);
and U17444 (N_17444,N_16432,N_16576);
nor U17445 (N_17445,N_16495,N_16629);
xnor U17446 (N_17446,N_16748,N_15857);
nor U17447 (N_17447,N_15727,N_16129);
or U17448 (N_17448,N_15605,N_16207);
or U17449 (N_17449,N_15874,N_15764);
nor U17450 (N_17450,N_16245,N_16791);
nand U17451 (N_17451,N_16233,N_16429);
or U17452 (N_17452,N_16218,N_15779);
and U17453 (N_17453,N_16246,N_15753);
or U17454 (N_17454,N_16307,N_16152);
xnor U17455 (N_17455,N_15748,N_16085);
nor U17456 (N_17456,N_15623,N_15846);
nor U17457 (N_17457,N_16757,N_15619);
nand U17458 (N_17458,N_15617,N_16179);
xnor U17459 (N_17459,N_16190,N_16471);
nand U17460 (N_17460,N_15882,N_16518);
nor U17461 (N_17461,N_16508,N_15800);
xnor U17462 (N_17462,N_15686,N_16613);
or U17463 (N_17463,N_16509,N_15632);
nor U17464 (N_17464,N_15654,N_16266);
or U17465 (N_17465,N_16112,N_16338);
xor U17466 (N_17466,N_16228,N_15897);
xor U17467 (N_17467,N_15906,N_16165);
or U17468 (N_17468,N_15971,N_15679);
xor U17469 (N_17469,N_16018,N_16385);
and U17470 (N_17470,N_16028,N_15838);
and U17471 (N_17471,N_16722,N_16085);
and U17472 (N_17472,N_16587,N_16047);
nor U17473 (N_17473,N_15869,N_15606);
nor U17474 (N_17474,N_16451,N_16131);
or U17475 (N_17475,N_15779,N_15799);
and U17476 (N_17476,N_16290,N_16568);
nor U17477 (N_17477,N_15792,N_16308);
or U17478 (N_17478,N_16136,N_16519);
and U17479 (N_17479,N_15811,N_16775);
nand U17480 (N_17480,N_16476,N_15846);
and U17481 (N_17481,N_15763,N_16570);
and U17482 (N_17482,N_15749,N_16729);
xnor U17483 (N_17483,N_16555,N_16111);
xnor U17484 (N_17484,N_16082,N_16738);
nand U17485 (N_17485,N_15650,N_15898);
nand U17486 (N_17486,N_16095,N_16617);
and U17487 (N_17487,N_16293,N_15727);
nor U17488 (N_17488,N_16517,N_16366);
and U17489 (N_17489,N_16056,N_15688);
or U17490 (N_17490,N_15760,N_16751);
and U17491 (N_17491,N_15902,N_15896);
and U17492 (N_17492,N_16571,N_15852);
nand U17493 (N_17493,N_16747,N_16041);
xor U17494 (N_17494,N_16067,N_15723);
nor U17495 (N_17495,N_15864,N_16088);
nand U17496 (N_17496,N_16391,N_16659);
or U17497 (N_17497,N_16602,N_15698);
nand U17498 (N_17498,N_16067,N_16275);
nand U17499 (N_17499,N_16255,N_16730);
nand U17500 (N_17500,N_15750,N_15992);
or U17501 (N_17501,N_16623,N_16536);
or U17502 (N_17502,N_16479,N_15999);
and U17503 (N_17503,N_16508,N_15680);
nand U17504 (N_17504,N_15777,N_16024);
nor U17505 (N_17505,N_16047,N_16139);
nand U17506 (N_17506,N_15904,N_16678);
nand U17507 (N_17507,N_15987,N_16264);
nor U17508 (N_17508,N_16256,N_16598);
nor U17509 (N_17509,N_16405,N_16290);
nor U17510 (N_17510,N_16190,N_16157);
or U17511 (N_17511,N_16590,N_16743);
nand U17512 (N_17512,N_16159,N_15957);
xnor U17513 (N_17513,N_15967,N_16058);
or U17514 (N_17514,N_15825,N_15634);
or U17515 (N_17515,N_15620,N_16724);
xor U17516 (N_17516,N_16013,N_15722);
nor U17517 (N_17517,N_16507,N_16528);
and U17518 (N_17518,N_15752,N_16071);
nor U17519 (N_17519,N_16233,N_15845);
nor U17520 (N_17520,N_16765,N_16591);
nand U17521 (N_17521,N_16359,N_16243);
xor U17522 (N_17522,N_16362,N_15695);
and U17523 (N_17523,N_15981,N_16406);
and U17524 (N_17524,N_16534,N_16509);
xor U17525 (N_17525,N_16694,N_16186);
and U17526 (N_17526,N_15715,N_16202);
and U17527 (N_17527,N_16175,N_15689);
nand U17528 (N_17528,N_16198,N_15655);
nand U17529 (N_17529,N_16009,N_16010);
nor U17530 (N_17530,N_16048,N_16629);
nor U17531 (N_17531,N_16488,N_16360);
and U17532 (N_17532,N_15801,N_16284);
and U17533 (N_17533,N_15612,N_15935);
nand U17534 (N_17534,N_16192,N_15696);
or U17535 (N_17535,N_15730,N_15947);
nor U17536 (N_17536,N_16690,N_16196);
or U17537 (N_17537,N_15900,N_16166);
and U17538 (N_17538,N_16489,N_16128);
xnor U17539 (N_17539,N_16788,N_15813);
nor U17540 (N_17540,N_15867,N_16265);
xor U17541 (N_17541,N_16756,N_16027);
nor U17542 (N_17542,N_16178,N_16025);
or U17543 (N_17543,N_15761,N_16764);
or U17544 (N_17544,N_15864,N_15777);
and U17545 (N_17545,N_16466,N_15755);
nor U17546 (N_17546,N_16596,N_16798);
nor U17547 (N_17547,N_15966,N_16542);
nor U17548 (N_17548,N_16293,N_16753);
nor U17549 (N_17549,N_16219,N_16232);
nor U17550 (N_17550,N_16438,N_16601);
and U17551 (N_17551,N_15779,N_16745);
nand U17552 (N_17552,N_16503,N_15638);
nand U17553 (N_17553,N_15874,N_15712);
xnor U17554 (N_17554,N_16588,N_16027);
and U17555 (N_17555,N_16718,N_15653);
or U17556 (N_17556,N_16573,N_16105);
xor U17557 (N_17557,N_15856,N_16172);
nor U17558 (N_17558,N_15761,N_16552);
or U17559 (N_17559,N_16749,N_16607);
xor U17560 (N_17560,N_15672,N_15715);
and U17561 (N_17561,N_16000,N_15869);
nor U17562 (N_17562,N_16485,N_16657);
xnor U17563 (N_17563,N_16658,N_15837);
xor U17564 (N_17564,N_16614,N_16432);
and U17565 (N_17565,N_15895,N_16331);
xor U17566 (N_17566,N_16236,N_16659);
or U17567 (N_17567,N_15932,N_16486);
nor U17568 (N_17568,N_15947,N_16145);
xor U17569 (N_17569,N_16698,N_16238);
or U17570 (N_17570,N_16123,N_16365);
or U17571 (N_17571,N_15956,N_16678);
and U17572 (N_17572,N_15764,N_15835);
or U17573 (N_17573,N_16726,N_16259);
or U17574 (N_17574,N_16217,N_16168);
or U17575 (N_17575,N_16152,N_16246);
xor U17576 (N_17576,N_16111,N_15861);
nor U17577 (N_17577,N_16489,N_16288);
nor U17578 (N_17578,N_16340,N_15985);
and U17579 (N_17579,N_16638,N_16791);
or U17580 (N_17580,N_16535,N_15982);
nor U17581 (N_17581,N_15717,N_15631);
nor U17582 (N_17582,N_16143,N_16527);
nand U17583 (N_17583,N_15649,N_15651);
xor U17584 (N_17584,N_15753,N_15621);
or U17585 (N_17585,N_15681,N_15891);
nand U17586 (N_17586,N_15774,N_15940);
xor U17587 (N_17587,N_15717,N_16799);
xnor U17588 (N_17588,N_15985,N_16609);
and U17589 (N_17589,N_16155,N_16101);
or U17590 (N_17590,N_15737,N_15759);
nand U17591 (N_17591,N_16026,N_15704);
and U17592 (N_17592,N_16517,N_16101);
and U17593 (N_17593,N_16439,N_16416);
and U17594 (N_17594,N_15872,N_15960);
nor U17595 (N_17595,N_16532,N_16444);
nor U17596 (N_17596,N_16683,N_16544);
or U17597 (N_17597,N_16771,N_15990);
xnor U17598 (N_17598,N_16466,N_16729);
nor U17599 (N_17599,N_16407,N_16508);
and U17600 (N_17600,N_16684,N_16617);
xor U17601 (N_17601,N_16489,N_15698);
nor U17602 (N_17602,N_16120,N_15755);
xnor U17603 (N_17603,N_15998,N_16528);
xor U17604 (N_17604,N_15879,N_16081);
and U17605 (N_17605,N_16727,N_16421);
nand U17606 (N_17606,N_15819,N_15794);
or U17607 (N_17607,N_16667,N_16272);
or U17608 (N_17608,N_16079,N_16179);
xor U17609 (N_17609,N_16271,N_15763);
nor U17610 (N_17610,N_16794,N_15991);
xnor U17611 (N_17611,N_16491,N_16690);
nand U17612 (N_17612,N_16660,N_15640);
xnor U17613 (N_17613,N_15825,N_16601);
nor U17614 (N_17614,N_16155,N_15948);
nor U17615 (N_17615,N_16026,N_16292);
xnor U17616 (N_17616,N_15781,N_16054);
and U17617 (N_17617,N_16350,N_16611);
and U17618 (N_17618,N_16492,N_16411);
nand U17619 (N_17619,N_16099,N_16584);
and U17620 (N_17620,N_15873,N_16449);
or U17621 (N_17621,N_16089,N_16366);
xnor U17622 (N_17622,N_16712,N_15723);
nor U17623 (N_17623,N_16178,N_15960);
and U17624 (N_17624,N_16373,N_15916);
nor U17625 (N_17625,N_16190,N_16563);
xnor U17626 (N_17626,N_16463,N_16150);
and U17627 (N_17627,N_16329,N_15983);
nand U17628 (N_17628,N_16207,N_16258);
nand U17629 (N_17629,N_15781,N_16652);
nor U17630 (N_17630,N_16480,N_15854);
nand U17631 (N_17631,N_16097,N_16261);
nor U17632 (N_17632,N_16539,N_16674);
nor U17633 (N_17633,N_16025,N_16335);
xor U17634 (N_17634,N_16312,N_16550);
or U17635 (N_17635,N_16275,N_15673);
xnor U17636 (N_17636,N_16430,N_16620);
or U17637 (N_17637,N_16597,N_16178);
or U17638 (N_17638,N_15742,N_15712);
and U17639 (N_17639,N_16547,N_16331);
nand U17640 (N_17640,N_16486,N_15905);
nand U17641 (N_17641,N_15710,N_15912);
and U17642 (N_17642,N_16207,N_15881);
or U17643 (N_17643,N_16728,N_15764);
xnor U17644 (N_17644,N_16742,N_15643);
nor U17645 (N_17645,N_16216,N_15718);
or U17646 (N_17646,N_16648,N_16037);
xnor U17647 (N_17647,N_15906,N_15861);
xnor U17648 (N_17648,N_15768,N_16376);
and U17649 (N_17649,N_16696,N_16382);
nand U17650 (N_17650,N_15703,N_15965);
nand U17651 (N_17651,N_16711,N_15959);
nand U17652 (N_17652,N_16502,N_16320);
or U17653 (N_17653,N_16270,N_16501);
and U17654 (N_17654,N_16605,N_16164);
or U17655 (N_17655,N_15645,N_16418);
xnor U17656 (N_17656,N_15717,N_16622);
xor U17657 (N_17657,N_16271,N_16798);
and U17658 (N_17658,N_15847,N_16323);
xnor U17659 (N_17659,N_16049,N_16745);
and U17660 (N_17660,N_16147,N_16262);
and U17661 (N_17661,N_15895,N_15736);
nand U17662 (N_17662,N_16091,N_15934);
xor U17663 (N_17663,N_16559,N_15614);
xnor U17664 (N_17664,N_16711,N_16182);
nor U17665 (N_17665,N_15612,N_15817);
or U17666 (N_17666,N_16658,N_16692);
xor U17667 (N_17667,N_15648,N_16365);
nor U17668 (N_17668,N_15761,N_15906);
nand U17669 (N_17669,N_16199,N_16697);
nor U17670 (N_17670,N_16070,N_16000);
or U17671 (N_17671,N_16212,N_16092);
xor U17672 (N_17672,N_16593,N_16193);
xnor U17673 (N_17673,N_16316,N_16470);
and U17674 (N_17674,N_16250,N_16568);
nor U17675 (N_17675,N_15747,N_16546);
or U17676 (N_17676,N_15678,N_16461);
and U17677 (N_17677,N_15708,N_16345);
nor U17678 (N_17678,N_15918,N_15635);
xor U17679 (N_17679,N_16270,N_15696);
xnor U17680 (N_17680,N_15907,N_16278);
nor U17681 (N_17681,N_15928,N_16041);
xor U17682 (N_17682,N_16731,N_15733);
and U17683 (N_17683,N_16784,N_15639);
nor U17684 (N_17684,N_16092,N_15859);
or U17685 (N_17685,N_15731,N_15793);
or U17686 (N_17686,N_16508,N_15995);
or U17687 (N_17687,N_15629,N_15692);
or U17688 (N_17688,N_15919,N_16670);
or U17689 (N_17689,N_15777,N_16118);
and U17690 (N_17690,N_16438,N_16036);
xor U17691 (N_17691,N_16131,N_16122);
and U17692 (N_17692,N_16559,N_15714);
nor U17693 (N_17693,N_16353,N_16452);
xnor U17694 (N_17694,N_15994,N_16518);
or U17695 (N_17695,N_15601,N_16588);
or U17696 (N_17696,N_16294,N_16072);
xor U17697 (N_17697,N_16624,N_15983);
nand U17698 (N_17698,N_16793,N_16385);
and U17699 (N_17699,N_16271,N_16014);
or U17700 (N_17700,N_16229,N_16025);
nand U17701 (N_17701,N_15713,N_16782);
nor U17702 (N_17702,N_16250,N_16138);
or U17703 (N_17703,N_16516,N_15953);
and U17704 (N_17704,N_16586,N_16027);
nor U17705 (N_17705,N_15721,N_16132);
or U17706 (N_17706,N_15835,N_16460);
or U17707 (N_17707,N_16662,N_16189);
and U17708 (N_17708,N_16778,N_16525);
and U17709 (N_17709,N_16256,N_16150);
or U17710 (N_17710,N_16328,N_16507);
and U17711 (N_17711,N_16145,N_16345);
or U17712 (N_17712,N_16699,N_16012);
or U17713 (N_17713,N_15986,N_15876);
and U17714 (N_17714,N_15921,N_16617);
nor U17715 (N_17715,N_16229,N_16734);
nand U17716 (N_17716,N_15675,N_16126);
nor U17717 (N_17717,N_15713,N_16382);
or U17718 (N_17718,N_16239,N_16388);
nor U17719 (N_17719,N_16153,N_16617);
or U17720 (N_17720,N_15852,N_15707);
nand U17721 (N_17721,N_15776,N_16363);
nor U17722 (N_17722,N_16353,N_15964);
and U17723 (N_17723,N_16152,N_15727);
and U17724 (N_17724,N_16426,N_15713);
xnor U17725 (N_17725,N_16759,N_15973);
and U17726 (N_17726,N_16716,N_16176);
xnor U17727 (N_17727,N_15991,N_16643);
xnor U17728 (N_17728,N_16036,N_15963);
or U17729 (N_17729,N_16444,N_16104);
nand U17730 (N_17730,N_15629,N_15925);
and U17731 (N_17731,N_15983,N_16785);
nor U17732 (N_17732,N_15771,N_16670);
nor U17733 (N_17733,N_15830,N_15796);
xnor U17734 (N_17734,N_15969,N_16011);
nand U17735 (N_17735,N_16089,N_15731);
xor U17736 (N_17736,N_16649,N_15694);
nand U17737 (N_17737,N_16276,N_16471);
and U17738 (N_17738,N_15826,N_16227);
nor U17739 (N_17739,N_15938,N_16510);
xnor U17740 (N_17740,N_16298,N_16538);
xor U17741 (N_17741,N_16556,N_16184);
nor U17742 (N_17742,N_16707,N_16346);
nand U17743 (N_17743,N_15712,N_16717);
or U17744 (N_17744,N_16053,N_15637);
xor U17745 (N_17745,N_16001,N_15721);
and U17746 (N_17746,N_16779,N_16295);
xor U17747 (N_17747,N_15628,N_15684);
nor U17748 (N_17748,N_16143,N_15636);
xnor U17749 (N_17749,N_16113,N_15789);
nor U17750 (N_17750,N_15893,N_16154);
and U17751 (N_17751,N_16155,N_16617);
xor U17752 (N_17752,N_16592,N_16458);
xnor U17753 (N_17753,N_16188,N_16415);
or U17754 (N_17754,N_15650,N_16601);
nor U17755 (N_17755,N_16695,N_16505);
and U17756 (N_17756,N_16776,N_16042);
xnor U17757 (N_17757,N_15758,N_16128);
and U17758 (N_17758,N_15762,N_16730);
nor U17759 (N_17759,N_16788,N_16499);
nand U17760 (N_17760,N_16338,N_16735);
or U17761 (N_17761,N_16290,N_16093);
and U17762 (N_17762,N_15765,N_15990);
or U17763 (N_17763,N_16060,N_16243);
nor U17764 (N_17764,N_16561,N_16651);
xnor U17765 (N_17765,N_15617,N_16641);
and U17766 (N_17766,N_16317,N_15693);
xor U17767 (N_17767,N_15707,N_16351);
xnor U17768 (N_17768,N_16693,N_16231);
xnor U17769 (N_17769,N_16122,N_16045);
and U17770 (N_17770,N_16087,N_15750);
xnor U17771 (N_17771,N_15731,N_15939);
or U17772 (N_17772,N_15946,N_16297);
xnor U17773 (N_17773,N_15749,N_16371);
xor U17774 (N_17774,N_16478,N_15770);
or U17775 (N_17775,N_16090,N_16432);
xnor U17776 (N_17776,N_16384,N_16648);
or U17777 (N_17777,N_16553,N_16320);
or U17778 (N_17778,N_16072,N_16233);
nor U17779 (N_17779,N_16044,N_16594);
nor U17780 (N_17780,N_16703,N_15936);
nor U17781 (N_17781,N_16331,N_16137);
nor U17782 (N_17782,N_15856,N_15906);
nor U17783 (N_17783,N_15891,N_16183);
or U17784 (N_17784,N_16534,N_16269);
nor U17785 (N_17785,N_15735,N_15657);
nor U17786 (N_17786,N_16319,N_16474);
or U17787 (N_17787,N_16560,N_15983);
nand U17788 (N_17788,N_16119,N_16574);
xor U17789 (N_17789,N_16578,N_16214);
and U17790 (N_17790,N_15863,N_15619);
or U17791 (N_17791,N_16371,N_16725);
xor U17792 (N_17792,N_15674,N_16200);
nand U17793 (N_17793,N_15610,N_16763);
or U17794 (N_17794,N_16143,N_15947);
and U17795 (N_17795,N_16182,N_16561);
and U17796 (N_17796,N_16234,N_16125);
nand U17797 (N_17797,N_16441,N_16086);
nor U17798 (N_17798,N_16473,N_16510);
nor U17799 (N_17799,N_15957,N_16580);
nand U17800 (N_17800,N_16612,N_16044);
nand U17801 (N_17801,N_15925,N_16038);
nand U17802 (N_17802,N_15996,N_16118);
xnor U17803 (N_17803,N_16285,N_16380);
xnor U17804 (N_17804,N_16021,N_15964);
nand U17805 (N_17805,N_16185,N_16732);
xnor U17806 (N_17806,N_16171,N_16499);
and U17807 (N_17807,N_16232,N_15823);
xnor U17808 (N_17808,N_16046,N_15667);
nor U17809 (N_17809,N_16551,N_16628);
and U17810 (N_17810,N_15931,N_15780);
nor U17811 (N_17811,N_15901,N_16603);
or U17812 (N_17812,N_16124,N_16691);
and U17813 (N_17813,N_16485,N_15626);
nand U17814 (N_17814,N_15875,N_16218);
xor U17815 (N_17815,N_16493,N_15966);
nor U17816 (N_17816,N_16321,N_16547);
and U17817 (N_17817,N_16756,N_16057);
or U17818 (N_17818,N_16416,N_15763);
xnor U17819 (N_17819,N_16108,N_16270);
nor U17820 (N_17820,N_16456,N_16688);
nor U17821 (N_17821,N_16536,N_16176);
xnor U17822 (N_17822,N_16660,N_16285);
nand U17823 (N_17823,N_15967,N_16617);
and U17824 (N_17824,N_16456,N_15872);
nor U17825 (N_17825,N_16307,N_15720);
nand U17826 (N_17826,N_15649,N_15848);
xor U17827 (N_17827,N_16257,N_16484);
and U17828 (N_17828,N_16132,N_15810);
and U17829 (N_17829,N_15815,N_15604);
and U17830 (N_17830,N_16126,N_16757);
or U17831 (N_17831,N_16146,N_16747);
or U17832 (N_17832,N_16305,N_16128);
xnor U17833 (N_17833,N_15899,N_15720);
and U17834 (N_17834,N_16350,N_16224);
nor U17835 (N_17835,N_15970,N_15701);
xnor U17836 (N_17836,N_16400,N_15683);
xnor U17837 (N_17837,N_15977,N_16119);
nor U17838 (N_17838,N_16575,N_16409);
nor U17839 (N_17839,N_15709,N_16003);
nor U17840 (N_17840,N_16078,N_16547);
or U17841 (N_17841,N_16489,N_16215);
nor U17842 (N_17842,N_16684,N_16022);
or U17843 (N_17843,N_15930,N_16545);
or U17844 (N_17844,N_16160,N_16169);
nor U17845 (N_17845,N_16409,N_16196);
nand U17846 (N_17846,N_16479,N_16153);
and U17847 (N_17847,N_16585,N_16327);
and U17848 (N_17848,N_15839,N_16332);
nand U17849 (N_17849,N_15790,N_15608);
xor U17850 (N_17850,N_16367,N_15914);
nand U17851 (N_17851,N_15729,N_16402);
nand U17852 (N_17852,N_16214,N_16088);
and U17853 (N_17853,N_15708,N_16674);
nor U17854 (N_17854,N_16218,N_15961);
xnor U17855 (N_17855,N_16464,N_15898);
or U17856 (N_17856,N_16733,N_16029);
or U17857 (N_17857,N_16298,N_16724);
nand U17858 (N_17858,N_16563,N_16176);
nor U17859 (N_17859,N_16239,N_15693);
xor U17860 (N_17860,N_15685,N_16714);
or U17861 (N_17861,N_16231,N_15997);
xnor U17862 (N_17862,N_16242,N_16597);
or U17863 (N_17863,N_16555,N_16553);
nand U17864 (N_17864,N_16664,N_16021);
nor U17865 (N_17865,N_16232,N_16030);
or U17866 (N_17866,N_16187,N_16494);
nor U17867 (N_17867,N_16214,N_16055);
nand U17868 (N_17868,N_16521,N_15662);
xor U17869 (N_17869,N_15817,N_16755);
or U17870 (N_17870,N_15860,N_16223);
nor U17871 (N_17871,N_15802,N_16512);
or U17872 (N_17872,N_15730,N_16566);
xor U17873 (N_17873,N_16000,N_15754);
and U17874 (N_17874,N_16749,N_15656);
nand U17875 (N_17875,N_16277,N_16620);
xnor U17876 (N_17876,N_16646,N_16153);
xnor U17877 (N_17877,N_16200,N_15789);
or U17878 (N_17878,N_16429,N_16130);
nor U17879 (N_17879,N_15884,N_15856);
nor U17880 (N_17880,N_16165,N_16478);
nor U17881 (N_17881,N_16146,N_16750);
or U17882 (N_17882,N_15719,N_15692);
or U17883 (N_17883,N_15896,N_15615);
nor U17884 (N_17884,N_16515,N_16458);
xor U17885 (N_17885,N_16719,N_15735);
and U17886 (N_17886,N_15600,N_15898);
and U17887 (N_17887,N_15687,N_16056);
or U17888 (N_17888,N_16278,N_16545);
xnor U17889 (N_17889,N_16502,N_15668);
nor U17890 (N_17890,N_16600,N_16072);
nor U17891 (N_17891,N_15770,N_16174);
xnor U17892 (N_17892,N_16426,N_16291);
xor U17893 (N_17893,N_16379,N_16322);
nor U17894 (N_17894,N_16612,N_15845);
or U17895 (N_17895,N_16750,N_16116);
or U17896 (N_17896,N_15934,N_15875);
nor U17897 (N_17897,N_15823,N_16143);
or U17898 (N_17898,N_15783,N_16246);
or U17899 (N_17899,N_15984,N_16450);
and U17900 (N_17900,N_16368,N_15619);
nor U17901 (N_17901,N_15724,N_15747);
and U17902 (N_17902,N_16498,N_16461);
nor U17903 (N_17903,N_16769,N_15656);
or U17904 (N_17904,N_16249,N_16129);
nor U17905 (N_17905,N_15928,N_16365);
or U17906 (N_17906,N_15611,N_15923);
and U17907 (N_17907,N_16457,N_16397);
xor U17908 (N_17908,N_16319,N_16723);
and U17909 (N_17909,N_15909,N_15799);
and U17910 (N_17910,N_16575,N_16379);
nor U17911 (N_17911,N_16360,N_15973);
nand U17912 (N_17912,N_16719,N_15847);
nand U17913 (N_17913,N_15900,N_16210);
nor U17914 (N_17914,N_16188,N_16588);
and U17915 (N_17915,N_16114,N_15918);
and U17916 (N_17916,N_16007,N_15745);
nor U17917 (N_17917,N_16673,N_16210);
and U17918 (N_17918,N_16587,N_16040);
nand U17919 (N_17919,N_15756,N_15810);
xnor U17920 (N_17920,N_16087,N_16248);
or U17921 (N_17921,N_15879,N_16023);
and U17922 (N_17922,N_15775,N_15914);
xor U17923 (N_17923,N_16403,N_16166);
and U17924 (N_17924,N_15615,N_16227);
nor U17925 (N_17925,N_16197,N_16396);
nor U17926 (N_17926,N_16719,N_16095);
xnor U17927 (N_17927,N_16377,N_16512);
and U17928 (N_17928,N_16344,N_16044);
xor U17929 (N_17929,N_16138,N_16624);
or U17930 (N_17930,N_16060,N_15972);
nand U17931 (N_17931,N_16315,N_15945);
nor U17932 (N_17932,N_16091,N_16159);
nand U17933 (N_17933,N_15734,N_16064);
nor U17934 (N_17934,N_15752,N_16131);
nor U17935 (N_17935,N_16421,N_16063);
xnor U17936 (N_17936,N_15873,N_16691);
nor U17937 (N_17937,N_15643,N_16185);
xnor U17938 (N_17938,N_16726,N_15963);
xor U17939 (N_17939,N_16051,N_16245);
nand U17940 (N_17940,N_16775,N_16110);
nor U17941 (N_17941,N_16517,N_16389);
xor U17942 (N_17942,N_15651,N_15618);
nand U17943 (N_17943,N_15945,N_16537);
and U17944 (N_17944,N_16357,N_15916);
nand U17945 (N_17945,N_15688,N_15983);
nand U17946 (N_17946,N_15834,N_16155);
xor U17947 (N_17947,N_15649,N_15974);
nor U17948 (N_17948,N_16620,N_15843);
xor U17949 (N_17949,N_15755,N_16600);
or U17950 (N_17950,N_16697,N_16421);
nand U17951 (N_17951,N_16781,N_15681);
and U17952 (N_17952,N_15993,N_15739);
nand U17953 (N_17953,N_16132,N_15975);
or U17954 (N_17954,N_16568,N_16037);
and U17955 (N_17955,N_16625,N_16038);
or U17956 (N_17956,N_15691,N_15809);
nor U17957 (N_17957,N_16428,N_16785);
and U17958 (N_17958,N_15884,N_16390);
nor U17959 (N_17959,N_16671,N_16297);
xor U17960 (N_17960,N_15729,N_16648);
and U17961 (N_17961,N_15993,N_16283);
and U17962 (N_17962,N_15636,N_15856);
nor U17963 (N_17963,N_16538,N_15682);
and U17964 (N_17964,N_16696,N_16202);
and U17965 (N_17965,N_16006,N_15782);
nand U17966 (N_17966,N_15904,N_15605);
nor U17967 (N_17967,N_16245,N_16307);
and U17968 (N_17968,N_16005,N_16136);
xor U17969 (N_17969,N_15888,N_16274);
xnor U17970 (N_17970,N_16140,N_15718);
xor U17971 (N_17971,N_15880,N_16447);
nand U17972 (N_17972,N_15954,N_16694);
nor U17973 (N_17973,N_16108,N_16419);
xnor U17974 (N_17974,N_16662,N_15870);
or U17975 (N_17975,N_16741,N_16627);
or U17976 (N_17976,N_16579,N_15684);
or U17977 (N_17977,N_16493,N_16300);
and U17978 (N_17978,N_16085,N_16698);
and U17979 (N_17979,N_16301,N_16367);
nand U17980 (N_17980,N_16537,N_16051);
nor U17981 (N_17981,N_16383,N_15882);
xnor U17982 (N_17982,N_16235,N_16479);
or U17983 (N_17983,N_15638,N_16635);
or U17984 (N_17984,N_16043,N_15640);
nor U17985 (N_17985,N_16601,N_16327);
nand U17986 (N_17986,N_16185,N_15722);
xor U17987 (N_17987,N_16311,N_15735);
and U17988 (N_17988,N_15734,N_16557);
and U17989 (N_17989,N_16660,N_15993);
and U17990 (N_17990,N_16325,N_16220);
or U17991 (N_17991,N_16196,N_16338);
nand U17992 (N_17992,N_16049,N_15999);
and U17993 (N_17993,N_15909,N_16191);
xnor U17994 (N_17994,N_16476,N_16162);
nand U17995 (N_17995,N_15942,N_15882);
and U17996 (N_17996,N_16360,N_16416);
xnor U17997 (N_17997,N_16053,N_16064);
xnor U17998 (N_17998,N_16021,N_16402);
xnor U17999 (N_17999,N_15693,N_15888);
or U18000 (N_18000,N_17432,N_17947);
nor U18001 (N_18001,N_17266,N_16973);
nand U18002 (N_18002,N_17951,N_17176);
and U18003 (N_18003,N_17654,N_17684);
or U18004 (N_18004,N_17337,N_17930);
xnor U18005 (N_18005,N_17300,N_17236);
and U18006 (N_18006,N_17203,N_17994);
nor U18007 (N_18007,N_16980,N_17000);
or U18008 (N_18008,N_16808,N_17573);
nor U18009 (N_18009,N_17928,N_17604);
xnor U18010 (N_18010,N_17957,N_16959);
nor U18011 (N_18011,N_17486,N_17144);
and U18012 (N_18012,N_17755,N_16816);
xnor U18013 (N_18013,N_17088,N_17105);
and U18014 (N_18014,N_17991,N_17931);
nand U18015 (N_18015,N_17914,N_17122);
nor U18016 (N_18016,N_17079,N_17652);
xnor U18017 (N_18017,N_17075,N_17511);
and U18018 (N_18018,N_17466,N_17966);
nor U18019 (N_18019,N_17155,N_17864);
xor U18020 (N_18020,N_17272,N_17160);
nor U18021 (N_18021,N_17166,N_16809);
nand U18022 (N_18022,N_17926,N_17482);
xor U18023 (N_18023,N_17238,N_17935);
or U18024 (N_18024,N_16845,N_17901);
or U18025 (N_18025,N_16911,N_17233);
nand U18026 (N_18026,N_17006,N_16918);
xnor U18027 (N_18027,N_17336,N_17567);
nand U18028 (N_18028,N_17642,N_17761);
nand U18029 (N_18029,N_17998,N_17577);
nand U18030 (N_18030,N_17237,N_17867);
or U18031 (N_18031,N_17841,N_17764);
nor U18032 (N_18032,N_17177,N_17164);
nand U18033 (N_18033,N_17549,N_17054);
xnor U18034 (N_18034,N_16938,N_17838);
nand U18035 (N_18035,N_17501,N_17769);
xor U18036 (N_18036,N_17607,N_17110);
nand U18037 (N_18037,N_17396,N_17284);
nand U18038 (N_18038,N_17219,N_17081);
and U18039 (N_18039,N_17025,N_16928);
nand U18040 (N_18040,N_16860,N_17814);
nand U18041 (N_18041,N_17545,N_17460);
nand U18042 (N_18042,N_17475,N_17473);
nand U18043 (N_18043,N_17368,N_17133);
or U18044 (N_18044,N_17766,N_17859);
nand U18045 (N_18045,N_17318,N_17039);
or U18046 (N_18046,N_17314,N_17708);
or U18047 (N_18047,N_17463,N_17013);
and U18048 (N_18048,N_17468,N_16818);
nor U18049 (N_18049,N_17269,N_17832);
nand U18050 (N_18050,N_17023,N_17274);
xor U18051 (N_18051,N_17627,N_17303);
xor U18052 (N_18052,N_16810,N_17772);
nor U18053 (N_18053,N_17228,N_16800);
nand U18054 (N_18054,N_17608,N_17297);
nor U18055 (N_18055,N_17896,N_16830);
nor U18056 (N_18056,N_17637,N_17397);
xor U18057 (N_18057,N_16812,N_17257);
nor U18058 (N_18058,N_17096,N_17724);
and U18059 (N_18059,N_17165,N_17571);
and U18060 (N_18060,N_17622,N_17973);
nand U18061 (N_18061,N_17844,N_17967);
xnor U18062 (N_18062,N_17391,N_17097);
xor U18063 (N_18063,N_17854,N_17375);
and U18064 (N_18064,N_17884,N_17737);
and U18065 (N_18065,N_17002,N_17268);
xnor U18066 (N_18066,N_17270,N_17941);
or U18067 (N_18067,N_17979,N_17090);
or U18068 (N_18068,N_17344,N_17467);
xor U18069 (N_18069,N_17371,N_16965);
and U18070 (N_18070,N_17835,N_17358);
xnor U18071 (N_18071,N_17619,N_17181);
and U18072 (N_18072,N_17395,N_17848);
nand U18073 (N_18073,N_17028,N_17906);
nand U18074 (N_18074,N_17639,N_17856);
nand U18075 (N_18075,N_17083,N_17647);
or U18076 (N_18076,N_17971,N_17044);
xor U18077 (N_18077,N_17161,N_17156);
nor U18078 (N_18078,N_17747,N_17311);
and U18079 (N_18079,N_17863,N_17184);
or U18080 (N_18080,N_17064,N_17768);
nand U18081 (N_18081,N_17005,N_17965);
xor U18082 (N_18082,N_17646,N_17182);
or U18083 (N_18083,N_17940,N_17774);
nor U18084 (N_18084,N_17046,N_17406);
and U18085 (N_18085,N_16881,N_16984);
and U18086 (N_18086,N_17449,N_17056);
xor U18087 (N_18087,N_17052,N_17362);
or U18088 (N_18088,N_17826,N_17218);
or U18089 (N_18089,N_16912,N_17992);
nand U18090 (N_18090,N_17405,N_16992);
xnor U18091 (N_18091,N_16892,N_17869);
or U18092 (N_18092,N_17602,N_17943);
or U18093 (N_18093,N_17656,N_17249);
or U18094 (N_18094,N_17040,N_17464);
nand U18095 (N_18095,N_17618,N_17436);
and U18096 (N_18096,N_17180,N_17886);
nand U18097 (N_18097,N_17323,N_17235);
xor U18098 (N_18098,N_17102,N_17938);
and U18099 (N_18099,N_17111,N_17820);
nand U18100 (N_18100,N_17733,N_17600);
nor U18101 (N_18101,N_17365,N_17601);
and U18102 (N_18102,N_17158,N_16893);
nor U18103 (N_18103,N_17198,N_17698);
xor U18104 (N_18104,N_17433,N_17725);
or U18105 (N_18105,N_17765,N_17553);
and U18106 (N_18106,N_16967,N_16932);
or U18107 (N_18107,N_17092,N_17551);
xnor U18108 (N_18108,N_17528,N_17359);
and U18109 (N_18109,N_17702,N_17649);
and U18110 (N_18110,N_17374,N_17418);
xor U18111 (N_18111,N_17977,N_17167);
nand U18112 (N_18112,N_17487,N_17072);
xor U18113 (N_18113,N_16941,N_17932);
nand U18114 (N_18114,N_16856,N_17690);
nor U18115 (N_18115,N_16957,N_17787);
nand U18116 (N_18116,N_17445,N_17470);
nor U18117 (N_18117,N_17253,N_17714);
and U18118 (N_18118,N_17369,N_17512);
or U18119 (N_18119,N_17021,N_17254);
nand U18120 (N_18120,N_16852,N_17523);
nand U18121 (N_18121,N_17675,N_17663);
or U18122 (N_18122,N_17408,N_17767);
xnor U18123 (N_18123,N_16970,N_17824);
xnor U18124 (N_18124,N_17471,N_16850);
and U18125 (N_18125,N_16962,N_17557);
nor U18126 (N_18126,N_17214,N_16991);
xnor U18127 (N_18127,N_17340,N_16875);
or U18128 (N_18128,N_17258,N_17658);
or U18129 (N_18129,N_17380,N_17407);
nand U18130 (N_18130,N_17558,N_17587);
or U18131 (N_18131,N_17756,N_17026);
nor U18132 (N_18132,N_17829,N_17148);
and U18133 (N_18133,N_17672,N_17332);
nand U18134 (N_18134,N_17715,N_17648);
nand U18135 (N_18135,N_17506,N_17354);
xnor U18136 (N_18136,N_17862,N_17498);
nand U18137 (N_18137,N_17377,N_17655);
xor U18138 (N_18138,N_17413,N_17596);
nand U18139 (N_18139,N_17908,N_17923);
nor U18140 (N_18140,N_17221,N_16833);
and U18141 (N_18141,N_17172,N_17041);
nor U18142 (N_18142,N_16815,N_16937);
nor U18143 (N_18143,N_16993,N_17055);
or U18144 (N_18144,N_17985,N_16897);
nor U18145 (N_18145,N_16895,N_17252);
xor U18146 (N_18146,N_17222,N_17282);
xnor U18147 (N_18147,N_16996,N_17705);
and U18148 (N_18148,N_17179,N_16806);
nand U18149 (N_18149,N_16872,N_17997);
nor U18150 (N_18150,N_17280,N_17423);
xnor U18151 (N_18151,N_17146,N_17461);
or U18152 (N_18152,N_17849,N_17409);
xor U18153 (N_18153,N_17921,N_17500);
or U18154 (N_18154,N_17846,N_17411);
or U18155 (N_18155,N_17738,N_17566);
nor U18156 (N_18156,N_17630,N_17902);
or U18157 (N_18157,N_17858,N_16926);
nor U18158 (N_18158,N_16976,N_17312);
nor U18159 (N_18159,N_17799,N_17749);
nand U18160 (N_18160,N_17352,N_17924);
or U18161 (N_18161,N_16844,N_17806);
xor U18162 (N_18162,N_17792,N_17537);
nand U18163 (N_18163,N_17212,N_17350);
nor U18164 (N_18164,N_17533,N_17718);
nand U18165 (N_18165,N_17812,N_17907);
nand U18166 (N_18166,N_16819,N_17098);
nand U18167 (N_18167,N_17990,N_17011);
xnor U18168 (N_18168,N_17050,N_17825);
and U18169 (N_18169,N_17495,N_17509);
nor U18170 (N_18170,N_17584,N_17968);
or U18171 (N_18171,N_17682,N_17494);
xnor U18172 (N_18172,N_17978,N_17163);
or U18173 (N_18173,N_16989,N_16886);
nor U18174 (N_18174,N_17834,N_17527);
and U18175 (N_18175,N_17197,N_16823);
nand U18176 (N_18176,N_17568,N_17925);
xnor U18177 (N_18177,N_17817,N_17113);
nor U18178 (N_18178,N_17448,N_16825);
nand U18179 (N_18179,N_17692,N_17481);
and U18180 (N_18180,N_17583,N_17480);
and U18181 (N_18181,N_17561,N_17964);
nor U18182 (N_18182,N_17898,N_17091);
xor U18183 (N_18183,N_17136,N_17731);
nand U18184 (N_18184,N_16822,N_16807);
xnor U18185 (N_18185,N_17911,N_17681);
nor U18186 (N_18186,N_17211,N_17114);
xor U18187 (N_18187,N_17525,N_17572);
and U18188 (N_18188,N_17119,N_17239);
nor U18189 (N_18189,N_17469,N_17813);
xnor U18190 (N_18190,N_17539,N_17289);
and U18191 (N_18191,N_17707,N_17808);
nand U18192 (N_18192,N_17351,N_17744);
or U18193 (N_18193,N_17443,N_17868);
nor U18194 (N_18194,N_17309,N_17620);
and U18195 (N_18195,N_17983,N_17379);
xnor U18196 (N_18196,N_16944,N_17229);
nand U18197 (N_18197,N_16862,N_17195);
and U18198 (N_18198,N_17123,N_17430);
and U18199 (N_18199,N_17012,N_17259);
nand U18200 (N_18200,N_16972,N_17325);
nand U18201 (N_18201,N_17169,N_17945);
nand U18202 (N_18202,N_17936,N_16958);
and U18203 (N_18203,N_16885,N_17067);
or U18204 (N_18204,N_17191,N_16848);
xor U18205 (N_18205,N_17010,N_17700);
or U18206 (N_18206,N_17816,N_17209);
or U18207 (N_18207,N_16922,N_17771);
nor U18208 (N_18208,N_17783,N_17544);
or U18209 (N_18209,N_17192,N_16975);
and U18210 (N_18210,N_17697,N_17240);
nand U18211 (N_18211,N_17126,N_17538);
xnor U18212 (N_18212,N_17415,N_17989);
nor U18213 (N_18213,N_17950,N_17283);
nor U18214 (N_18214,N_16920,N_17555);
nor U18215 (N_18215,N_17428,N_17033);
nand U18216 (N_18216,N_17030,N_17419);
nand U18217 (N_18217,N_17821,N_16909);
or U18218 (N_18218,N_17120,N_17676);
and U18219 (N_18219,N_17094,N_17503);
nand U18220 (N_18220,N_17758,N_17706);
nor U18221 (N_18221,N_17810,N_17807);
nand U18222 (N_18222,N_17962,N_16884);
nor U18223 (N_18223,N_17459,N_17691);
or U18224 (N_18224,N_17735,N_17322);
and U18225 (N_18225,N_17306,N_17770);
nand U18226 (N_18226,N_17290,N_17404);
nor U18227 (N_18227,N_17069,N_17581);
or U18228 (N_18228,N_16969,N_17385);
xor U18229 (N_18229,N_17640,N_17717);
or U18230 (N_18230,N_17417,N_17795);
nand U18231 (N_18231,N_17324,N_17004);
nand U18232 (N_18232,N_17232,N_17298);
or U18233 (N_18233,N_17696,N_16947);
or U18234 (N_18234,N_17546,N_17815);
xor U18235 (N_18235,N_17650,N_17559);
or U18236 (N_18236,N_17248,N_17890);
nor U18237 (N_18237,N_17877,N_17759);
or U18238 (N_18238,N_17876,N_17887);
nor U18239 (N_18239,N_16841,N_17830);
or U18240 (N_18240,N_16814,N_17634);
nor U18241 (N_18241,N_16880,N_17153);
or U18242 (N_18242,N_17134,N_17420);
xnor U18243 (N_18243,N_17505,N_17127);
xnor U18244 (N_18244,N_17739,N_17593);
nor U18245 (N_18245,N_17920,N_17393);
nor U18246 (N_18246,N_17210,N_16840);
xnor U18247 (N_18247,N_17918,N_17281);
xor U18248 (N_18248,N_17980,N_17595);
and U18249 (N_18249,N_17029,N_17905);
nor U18250 (N_18250,N_16832,N_17818);
xnor U18251 (N_18251,N_17387,N_17226);
and U18252 (N_18252,N_17410,N_16857);
nand U18253 (N_18253,N_16900,N_17900);
or U18254 (N_18254,N_16820,N_16999);
nand U18255 (N_18255,N_17591,N_17394);
and U18256 (N_18256,N_17014,N_17302);
nor U18257 (N_18257,N_17588,N_17452);
or U18258 (N_18258,N_17401,N_17893);
or U18259 (N_18259,N_16869,N_17889);
xor U18260 (N_18260,N_17047,N_17776);
or U18261 (N_18261,N_17491,N_17129);
and U18262 (N_18262,N_17709,N_17521);
nor U18263 (N_18263,N_16935,N_17355);
and U18264 (N_18264,N_17386,N_17330);
or U18265 (N_18265,N_17204,N_17636);
nand U18266 (N_18266,N_17366,N_17037);
nor U18267 (N_18267,N_17534,N_17597);
nand U18268 (N_18268,N_17353,N_17952);
nor U18269 (N_18269,N_17716,N_16858);
xor U18270 (N_18270,N_16916,N_17215);
nor U18271 (N_18271,N_17960,N_16802);
xnor U18272 (N_18272,N_17308,N_17851);
nand U18273 (N_18273,N_17343,N_17483);
or U18274 (N_18274,N_16877,N_17199);
nor U18275 (N_18275,N_17699,N_17036);
xor U18276 (N_18276,N_17916,N_16834);
xor U18277 (N_18277,N_16963,N_16936);
nor U18278 (N_18278,N_17242,N_17563);
xnor U18279 (N_18279,N_17296,N_17873);
and U18280 (N_18280,N_17256,N_17154);
or U18281 (N_18281,N_17103,N_17076);
or U18282 (N_18282,N_17187,N_17686);
and U18283 (N_18283,N_17424,N_17565);
or U18284 (N_18284,N_16889,N_17852);
or U18285 (N_18285,N_16966,N_17578);
xor U18286 (N_18286,N_17885,N_17245);
xor U18287 (N_18287,N_17271,N_16942);
nor U18288 (N_18288,N_17456,N_17661);
and U18289 (N_18289,N_16851,N_17513);
nand U18290 (N_18290,N_16867,N_17502);
xnor U18291 (N_18291,N_16952,N_17730);
xnor U18292 (N_18292,N_17562,N_17305);
nand U18293 (N_18293,N_17688,N_17683);
nor U18294 (N_18294,N_17579,N_17086);
nand U18295 (N_18295,N_17058,N_17760);
nor U18296 (N_18296,N_16994,N_17974);
and U18297 (N_18297,N_17342,N_17929);
nor U18298 (N_18298,N_17605,N_17291);
and U18299 (N_18299,N_17429,N_16955);
and U18300 (N_18300,N_17106,N_17141);
xor U18301 (N_18301,N_17987,N_17611);
or U18302 (N_18302,N_17477,N_17757);
or U18303 (N_18303,N_17454,N_17152);
or U18304 (N_18304,N_17594,N_17643);
nor U18305 (N_18305,N_17972,N_16882);
or U18306 (N_18306,N_16977,N_17363);
nand U18307 (N_18307,N_17694,N_17678);
xnor U18308 (N_18308,N_17223,N_17024);
nor U18309 (N_18309,N_17524,N_16817);
or U18310 (N_18310,N_16824,N_17328);
nand U18311 (N_18311,N_17061,N_17231);
xor U18312 (N_18312,N_16934,N_17117);
and U18313 (N_18313,N_17384,N_17984);
or U18314 (N_18314,N_17250,N_17208);
nand U18315 (N_18315,N_16871,N_17178);
nand U18316 (N_18316,N_16953,N_17162);
or U18317 (N_18317,N_16929,N_17334);
xnor U18318 (N_18318,N_17736,N_17059);
nand U18319 (N_18319,N_16925,N_17638);
nand U18320 (N_18320,N_17919,N_17084);
nand U18321 (N_18321,N_17586,N_17981);
nand U18322 (N_18322,N_17361,N_17399);
xor U18323 (N_18323,N_17788,N_17139);
and U18324 (N_18324,N_17132,N_16821);
or U18325 (N_18325,N_17552,N_17367);
or U18326 (N_18326,N_17213,N_17975);
nand U18327 (N_18327,N_17339,N_17453);
nand U18328 (N_18328,N_17777,N_17712);
xor U18329 (N_18329,N_17999,N_16843);
and U18330 (N_18330,N_17882,N_17115);
xnor U18331 (N_18331,N_17629,N_17427);
nor U18332 (N_18332,N_17216,N_17750);
nand U18333 (N_18333,N_17138,N_17934);
xor U18334 (N_18334,N_17704,N_16837);
or U18335 (N_18335,N_17437,N_17001);
nand U18336 (N_18336,N_17944,N_17288);
nor U18337 (N_18337,N_17616,N_17837);
xnor U18338 (N_18338,N_17194,N_17112);
nor U18339 (N_18339,N_16861,N_17492);
or U18340 (N_18340,N_17631,N_17617);
nand U18341 (N_18341,N_17099,N_17078);
or U18342 (N_18342,N_17752,N_17171);
xnor U18343 (N_18343,N_16986,N_17299);
and U18344 (N_18344,N_17917,N_17360);
nand U18345 (N_18345,N_16982,N_17939);
or U18346 (N_18346,N_17493,N_17442);
nor U18347 (N_18347,N_17937,N_16805);
nor U18348 (N_18348,N_17196,N_17895);
or U18349 (N_18349,N_17279,N_17400);
nand U18350 (N_18350,N_16887,N_17734);
nor U18351 (N_18351,N_17320,N_17791);
xnor U18352 (N_18352,N_17632,N_17273);
and U18353 (N_18353,N_17474,N_16946);
and U18354 (N_18354,N_17261,N_17653);
or U18355 (N_18355,N_17819,N_17635);
nand U18356 (N_18356,N_16829,N_17881);
or U18357 (N_18357,N_17892,N_17349);
or U18358 (N_18358,N_17986,N_17357);
and U18359 (N_18359,N_17836,N_17912);
nand U18360 (N_18360,N_17220,N_17319);
nor U18361 (N_18361,N_17671,N_17721);
xnor U18362 (N_18362,N_16971,N_17743);
or U18363 (N_18363,N_17243,N_17802);
nand U18364 (N_18364,N_17251,N_17020);
nor U18365 (N_18365,N_17711,N_17333);
nor U18366 (N_18366,N_17034,N_17548);
xnor U18367 (N_18367,N_17953,N_17225);
and U18368 (N_18368,N_17062,N_17621);
and U18369 (N_18369,N_17080,N_17897);
nand U18370 (N_18370,N_16968,N_17140);
and U18371 (N_18371,N_17489,N_17241);
and U18372 (N_18372,N_17070,N_16974);
and U18373 (N_18373,N_17190,N_17403);
or U18374 (N_18374,N_17753,N_17170);
or U18375 (N_18375,N_17189,N_17556);
and U18376 (N_18376,N_17713,N_16988);
and U18377 (N_18377,N_17060,N_17693);
or U18378 (N_18378,N_17441,N_17292);
xor U18379 (N_18379,N_17200,N_16855);
or U18380 (N_18380,N_17032,N_16896);
and U18381 (N_18381,N_17507,N_17077);
nor U18382 (N_18382,N_17183,N_17286);
and U18383 (N_18383,N_16853,N_16847);
xnor U18384 (N_18384,N_16883,N_17402);
nor U18385 (N_18385,N_16866,N_17599);
xor U18386 (N_18386,N_17125,N_17440);
xnor U18387 (N_18387,N_16899,N_17536);
nor U18388 (N_18388,N_17958,N_17276);
nor U18389 (N_18389,N_17662,N_17612);
nor U18390 (N_18390,N_16888,N_16835);
nand U18391 (N_18391,N_16870,N_17370);
and U18392 (N_18392,N_17496,N_17007);
and U18393 (N_18393,N_16813,N_17444);
nand U18394 (N_18394,N_17027,N_17626);
nor U18395 (N_18395,N_17346,N_17378);
and U18396 (N_18396,N_17870,N_16903);
nand U18397 (N_18397,N_17842,N_16979);
nor U18398 (N_18398,N_17022,N_16990);
nor U18399 (N_18399,N_17147,N_16940);
xor U18400 (N_18400,N_17703,N_17174);
or U18401 (N_18401,N_17186,N_17425);
and U18402 (N_18402,N_17674,N_17840);
and U18403 (N_18403,N_16854,N_17118);
or U18404 (N_18404,N_16836,N_17845);
or U18405 (N_18405,N_17657,N_17398);
and U18406 (N_18406,N_17828,N_16985);
nor U18407 (N_18407,N_17315,N_17942);
nand U18408 (N_18408,N_16997,N_17295);
nand U18409 (N_18409,N_17478,N_17455);
and U18410 (N_18410,N_17850,N_17063);
or U18411 (N_18411,N_17504,N_17540);
and U18412 (N_18412,N_16919,N_16804);
xnor U18413 (N_18413,N_17293,N_17175);
and U18414 (N_18414,N_17613,N_17742);
and U18415 (N_18415,N_17388,N_17159);
nor U18416 (N_18416,N_17285,N_17988);
xnor U18417 (N_18417,N_16839,N_17948);
nor U18418 (N_18418,N_17719,N_17899);
nand U18419 (N_18419,N_17121,N_17701);
nand U18420 (N_18420,N_16924,N_17476);
and U18421 (N_18421,N_17963,N_17909);
nor U18422 (N_18422,N_16868,N_17526);
nor U18423 (N_18423,N_16927,N_17053);
nand U18424 (N_18424,N_17341,N_17434);
xor U18425 (N_18425,N_17479,N_17458);
xor U18426 (N_18426,N_16842,N_17193);
or U18427 (N_18427,N_17781,N_17670);
nand U18428 (N_18428,N_17530,N_17575);
or U18429 (N_18429,N_17101,N_17224);
nand U18430 (N_18430,N_16983,N_17313);
nor U18431 (N_18431,N_16954,N_17762);
nor U18432 (N_18432,N_17687,N_17801);
nor U18433 (N_18433,N_17933,N_17438);
xnor U18434 (N_18434,N_17462,N_17982);
nor U18435 (N_18435,N_17922,N_17093);
and U18436 (N_18436,N_17710,N_17839);
nor U18437 (N_18437,N_17137,N_17517);
and U18438 (N_18438,N_17015,N_17008);
nand U18439 (N_18439,N_17490,N_16811);
and U18440 (N_18440,N_17592,N_16874);
xor U18441 (N_18441,N_17570,N_17522);
nor U18442 (N_18442,N_17157,N_17915);
nor U18443 (N_18443,N_17880,N_17109);
and U18444 (N_18444,N_17100,N_17531);
xor U18445 (N_18445,N_17085,N_17317);
xnor U18446 (N_18446,N_17874,N_17450);
nor U18447 (N_18447,N_17580,N_17412);
nand U18448 (N_18448,N_17472,N_17894);
and U18449 (N_18449,N_16960,N_17797);
nor U18450 (N_18450,N_17207,N_17878);
nand U18451 (N_18451,N_17035,N_17651);
or U18452 (N_18452,N_17741,N_17264);
xor U18453 (N_18453,N_17327,N_17446);
nor U18454 (N_18454,N_17543,N_17628);
and U18455 (N_18455,N_17860,N_16923);
xor U18456 (N_18456,N_17746,N_17488);
or U18457 (N_18457,N_17665,N_16961);
and U18458 (N_18458,N_16831,N_17541);
or U18459 (N_18459,N_17373,N_17255);
nor U18460 (N_18460,N_17664,N_16863);
xor U18461 (N_18461,N_16879,N_17135);
or U18462 (N_18462,N_17206,N_17372);
nand U18463 (N_18463,N_17451,N_17485);
or U18464 (N_18464,N_17392,N_16950);
xnor U18465 (N_18465,N_17667,N_17589);
nor U18466 (N_18466,N_17532,N_17585);
xnor U18467 (N_18467,N_16803,N_17310);
and U18468 (N_18468,N_17104,N_17390);
and U18469 (N_18469,N_17049,N_17497);
or U18470 (N_18470,N_16956,N_17574);
nand U18471 (N_18471,N_17499,N_17018);
nand U18472 (N_18472,N_17645,N_17603);
nor U18473 (N_18473,N_16894,N_17726);
xor U18474 (N_18474,N_17376,N_17805);
nand U18475 (N_18475,N_17927,N_17843);
nor U18476 (N_18476,N_17904,N_17009);
xor U18477 (N_18477,N_17508,N_17073);
nand U18478 (N_18478,N_16890,N_17623);
or U18479 (N_18479,N_17042,N_17205);
xnor U18480 (N_18480,N_17969,N_16998);
or U18481 (N_18481,N_17857,N_17872);
nor U18482 (N_18482,N_17677,N_17875);
or U18483 (N_18483,N_16995,N_17883);
nand U18484 (N_18484,N_17130,N_17065);
or U18485 (N_18485,N_17732,N_17262);
nor U18486 (N_18486,N_16801,N_17910);
xnor U18487 (N_18487,N_17800,N_17202);
xnor U18488 (N_18488,N_16902,N_17959);
and U18489 (N_18489,N_16915,N_16891);
and U18490 (N_18490,N_17775,N_17529);
or U18491 (N_18491,N_17230,N_17865);
nor U18492 (N_18492,N_16913,N_17431);
nand U18493 (N_18493,N_16914,N_16901);
xnor U18494 (N_18494,N_17149,N_17263);
or U18495 (N_18495,N_16930,N_17793);
xor U18496 (N_18496,N_17913,N_17294);
or U18497 (N_18497,N_17381,N_16864);
or U18498 (N_18498,N_16981,N_17057);
nor U18499 (N_18499,N_17803,N_17168);
and U18500 (N_18500,N_17773,N_17779);
xnor U18501 (N_18501,N_17831,N_17519);
nand U18502 (N_18502,N_16921,N_17903);
and U18503 (N_18503,N_17641,N_17510);
xor U18504 (N_18504,N_16978,N_17329);
xor U18505 (N_18505,N_17659,N_17082);
xor U18506 (N_18506,N_17569,N_17383);
nand U18507 (N_18507,N_16907,N_17201);
xnor U18508 (N_18508,N_17422,N_16948);
xnor U18509 (N_18509,N_17321,N_17689);
or U18510 (N_18510,N_17188,N_17789);
and U18511 (N_18511,N_17751,N_17518);
or U18512 (N_18512,N_17625,N_17108);
and U18513 (N_18513,N_17277,N_17031);
and U18514 (N_18514,N_17465,N_17554);
nand U18515 (N_18515,N_17326,N_17345);
nand U18516 (N_18516,N_17823,N_17389);
xnor U18517 (N_18517,N_17609,N_17457);
nor U18518 (N_18518,N_17784,N_16917);
xor U18519 (N_18519,N_17949,N_17666);
and U18520 (N_18520,N_17891,N_17866);
or U18521 (N_18521,N_17287,N_17019);
and U18522 (N_18522,N_17847,N_17068);
nand U18523 (N_18523,N_17804,N_17071);
nor U18524 (N_18524,N_17542,N_17364);
and U18525 (N_18525,N_17016,N_17822);
xnor U18526 (N_18526,N_17782,N_16939);
and U18527 (N_18527,N_17048,N_17143);
and U18528 (N_18528,N_17045,N_17560);
nand U18529 (N_18529,N_17685,N_17038);
and U18530 (N_18530,N_17644,N_17331);
nor U18531 (N_18531,N_17275,N_16951);
xnor U18532 (N_18532,N_17888,N_17116);
nor U18533 (N_18533,N_17680,N_17260);
or U18534 (N_18534,N_17576,N_17633);
nand U18535 (N_18535,N_17778,N_17435);
and U18536 (N_18536,N_16876,N_17142);
or U18537 (N_18537,N_16898,N_17796);
and U18538 (N_18538,N_17348,N_17614);
nor U18539 (N_18539,N_16878,N_17234);
nand U18540 (N_18540,N_17763,N_17955);
or U18541 (N_18541,N_17151,N_17003);
xor U18542 (N_18542,N_17679,N_17439);
and U18543 (N_18543,N_17745,N_17043);
and U18544 (N_18544,N_17729,N_17615);
nor U18545 (N_18545,N_16987,N_17307);
nor U18546 (N_18546,N_17173,N_16827);
nor U18547 (N_18547,N_17811,N_17660);
and U18548 (N_18548,N_17246,N_17267);
xor U18549 (N_18549,N_17720,N_17853);
xnor U18550 (N_18550,N_17780,N_17107);
nor U18551 (N_18551,N_17416,N_16910);
or U18552 (N_18552,N_17809,N_16859);
xnor U18553 (N_18553,N_16945,N_17871);
and U18554 (N_18554,N_17669,N_17879);
and U18555 (N_18555,N_17335,N_17740);
nand U18556 (N_18556,N_16931,N_17074);
and U18557 (N_18557,N_17786,N_17976);
nor U18558 (N_18558,N_17550,N_17582);
or U18559 (N_18559,N_17993,N_17535);
xnor U18560 (N_18560,N_16838,N_17278);
or U18561 (N_18561,N_16904,N_16943);
and U18562 (N_18562,N_17382,N_16949);
xor U18563 (N_18563,N_17785,N_17754);
or U18564 (N_18564,N_17265,N_16964);
or U18565 (N_18565,N_17790,N_17244);
xnor U18566 (N_18566,N_17185,N_17748);
nand U18567 (N_18567,N_17217,N_17598);
and U18568 (N_18568,N_16846,N_17316);
nor U18569 (N_18569,N_17150,N_17827);
xnor U18570 (N_18570,N_16826,N_17301);
and U18571 (N_18571,N_17668,N_17484);
and U18572 (N_18572,N_17961,N_17946);
nor U18573 (N_18573,N_17727,N_17606);
xor U18574 (N_18574,N_17414,N_16828);
nor U18575 (N_18575,N_17066,N_17095);
nor U18576 (N_18576,N_17590,N_17723);
and U18577 (N_18577,N_17304,N_17855);
nor U18578 (N_18578,N_17426,N_16865);
nand U18579 (N_18579,N_17051,N_17695);
or U18580 (N_18580,N_17996,N_17516);
nand U18581 (N_18581,N_16906,N_17356);
nand U18582 (N_18582,N_17515,N_17610);
nor U18583 (N_18583,N_17564,N_17547);
and U18584 (N_18584,N_17954,N_17995);
or U18585 (N_18585,N_17728,N_17338);
nor U18586 (N_18586,N_17447,N_16908);
nand U18587 (N_18587,N_17956,N_17520);
xor U18588 (N_18588,N_17347,N_17145);
xor U18589 (N_18589,N_16849,N_17970);
nor U18590 (N_18590,N_17861,N_17128);
xor U18591 (N_18591,N_17798,N_17131);
nand U18592 (N_18592,N_16905,N_17227);
xor U18593 (N_18593,N_17514,N_17089);
nand U18594 (N_18594,N_17421,N_17624);
nand U18595 (N_18595,N_16933,N_17794);
xor U18596 (N_18596,N_17722,N_17124);
nand U18597 (N_18597,N_17017,N_16873);
nor U18598 (N_18598,N_17087,N_17833);
or U18599 (N_18599,N_17673,N_17247);
and U18600 (N_18600,N_17267,N_16840);
nor U18601 (N_18601,N_17059,N_17596);
or U18602 (N_18602,N_16835,N_16857);
xnor U18603 (N_18603,N_17949,N_17990);
xnor U18604 (N_18604,N_16892,N_17313);
nor U18605 (N_18605,N_17913,N_17855);
xnor U18606 (N_18606,N_17123,N_16810);
nor U18607 (N_18607,N_17593,N_17527);
xnor U18608 (N_18608,N_17778,N_17533);
and U18609 (N_18609,N_17492,N_17381);
nor U18610 (N_18610,N_17190,N_16833);
nor U18611 (N_18611,N_17883,N_17940);
nor U18612 (N_18612,N_17742,N_17788);
or U18613 (N_18613,N_17912,N_17881);
xor U18614 (N_18614,N_16849,N_17329);
and U18615 (N_18615,N_17728,N_17729);
xnor U18616 (N_18616,N_17626,N_17093);
nand U18617 (N_18617,N_17910,N_17232);
xor U18618 (N_18618,N_17053,N_17420);
and U18619 (N_18619,N_16898,N_17434);
xor U18620 (N_18620,N_17735,N_17562);
and U18621 (N_18621,N_17480,N_17260);
nand U18622 (N_18622,N_17385,N_17783);
xnor U18623 (N_18623,N_17221,N_17503);
xor U18624 (N_18624,N_17655,N_17107);
and U18625 (N_18625,N_17782,N_17349);
xor U18626 (N_18626,N_17948,N_17094);
and U18627 (N_18627,N_17293,N_16874);
xnor U18628 (N_18628,N_17728,N_16996);
and U18629 (N_18629,N_17991,N_17060);
or U18630 (N_18630,N_17613,N_17721);
xor U18631 (N_18631,N_17489,N_17318);
or U18632 (N_18632,N_16801,N_17481);
xnor U18633 (N_18633,N_17415,N_17912);
nor U18634 (N_18634,N_17566,N_17444);
xnor U18635 (N_18635,N_16836,N_17471);
xor U18636 (N_18636,N_17821,N_17746);
xor U18637 (N_18637,N_16834,N_17925);
nand U18638 (N_18638,N_17947,N_17825);
nor U18639 (N_18639,N_17635,N_16847);
xnor U18640 (N_18640,N_17766,N_17862);
or U18641 (N_18641,N_17098,N_17210);
nor U18642 (N_18642,N_17845,N_16840);
and U18643 (N_18643,N_17158,N_17817);
xnor U18644 (N_18644,N_17559,N_17393);
or U18645 (N_18645,N_17038,N_17307);
nor U18646 (N_18646,N_17965,N_17774);
nand U18647 (N_18647,N_16912,N_17681);
xnor U18648 (N_18648,N_16899,N_17903);
nor U18649 (N_18649,N_17733,N_17110);
nor U18650 (N_18650,N_17034,N_17892);
nor U18651 (N_18651,N_17014,N_17356);
and U18652 (N_18652,N_17238,N_17164);
xor U18653 (N_18653,N_17277,N_17559);
or U18654 (N_18654,N_17421,N_17278);
and U18655 (N_18655,N_16976,N_17947);
xor U18656 (N_18656,N_17803,N_17498);
nor U18657 (N_18657,N_17790,N_17724);
or U18658 (N_18658,N_17617,N_17246);
or U18659 (N_18659,N_17297,N_17011);
xnor U18660 (N_18660,N_17175,N_16965);
nor U18661 (N_18661,N_17614,N_17451);
and U18662 (N_18662,N_16985,N_17570);
nor U18663 (N_18663,N_17539,N_17706);
or U18664 (N_18664,N_17297,N_17361);
and U18665 (N_18665,N_17505,N_17525);
or U18666 (N_18666,N_17363,N_17147);
or U18667 (N_18667,N_17266,N_17343);
xor U18668 (N_18668,N_16961,N_16877);
xor U18669 (N_18669,N_17301,N_17532);
nor U18670 (N_18670,N_17616,N_16991);
nand U18671 (N_18671,N_17238,N_17274);
or U18672 (N_18672,N_17239,N_17118);
nor U18673 (N_18673,N_17849,N_17989);
or U18674 (N_18674,N_17949,N_17470);
or U18675 (N_18675,N_17767,N_17464);
nand U18676 (N_18676,N_17358,N_17656);
and U18677 (N_18677,N_17273,N_16884);
nand U18678 (N_18678,N_17521,N_17227);
or U18679 (N_18679,N_16886,N_17541);
nand U18680 (N_18680,N_16877,N_17448);
xnor U18681 (N_18681,N_16869,N_17420);
xor U18682 (N_18682,N_17387,N_17091);
xor U18683 (N_18683,N_17603,N_17776);
nand U18684 (N_18684,N_17126,N_17278);
and U18685 (N_18685,N_17520,N_17239);
and U18686 (N_18686,N_17302,N_16958);
or U18687 (N_18687,N_17575,N_17894);
or U18688 (N_18688,N_17628,N_17777);
xor U18689 (N_18689,N_17499,N_16844);
or U18690 (N_18690,N_16955,N_17077);
and U18691 (N_18691,N_16946,N_17791);
nor U18692 (N_18692,N_17207,N_17039);
nor U18693 (N_18693,N_17555,N_17715);
or U18694 (N_18694,N_17203,N_17146);
and U18695 (N_18695,N_17819,N_16987);
nand U18696 (N_18696,N_17091,N_17008);
and U18697 (N_18697,N_17611,N_16844);
and U18698 (N_18698,N_16953,N_16825);
nand U18699 (N_18699,N_17023,N_16945);
nor U18700 (N_18700,N_16810,N_17910);
and U18701 (N_18701,N_17230,N_17114);
or U18702 (N_18702,N_17212,N_16932);
xnor U18703 (N_18703,N_17360,N_17972);
and U18704 (N_18704,N_17975,N_17615);
nor U18705 (N_18705,N_17863,N_17501);
nor U18706 (N_18706,N_17492,N_17052);
and U18707 (N_18707,N_17288,N_17703);
nand U18708 (N_18708,N_17988,N_17917);
or U18709 (N_18709,N_17994,N_17138);
nand U18710 (N_18710,N_17456,N_17309);
nand U18711 (N_18711,N_17878,N_17180);
nor U18712 (N_18712,N_17347,N_17602);
and U18713 (N_18713,N_17668,N_17256);
xnor U18714 (N_18714,N_16838,N_17562);
xnor U18715 (N_18715,N_17172,N_17390);
nand U18716 (N_18716,N_17103,N_17584);
nor U18717 (N_18717,N_17492,N_17426);
or U18718 (N_18718,N_17411,N_17744);
nand U18719 (N_18719,N_17423,N_17595);
and U18720 (N_18720,N_17254,N_16864);
nor U18721 (N_18721,N_16819,N_17550);
nand U18722 (N_18722,N_17690,N_17698);
nand U18723 (N_18723,N_17131,N_17485);
or U18724 (N_18724,N_17236,N_16816);
or U18725 (N_18725,N_16871,N_17131);
xnor U18726 (N_18726,N_17730,N_17991);
or U18727 (N_18727,N_17407,N_17245);
and U18728 (N_18728,N_16867,N_17383);
xnor U18729 (N_18729,N_17425,N_17454);
nor U18730 (N_18730,N_17474,N_17889);
nand U18731 (N_18731,N_17816,N_17043);
nand U18732 (N_18732,N_17621,N_17032);
and U18733 (N_18733,N_17753,N_17672);
nand U18734 (N_18734,N_17757,N_17817);
or U18735 (N_18735,N_17600,N_16883);
and U18736 (N_18736,N_17348,N_17473);
xor U18737 (N_18737,N_17050,N_17923);
and U18738 (N_18738,N_16894,N_17069);
xor U18739 (N_18739,N_16900,N_17337);
or U18740 (N_18740,N_17995,N_17772);
nand U18741 (N_18741,N_17846,N_17810);
nor U18742 (N_18742,N_16950,N_17922);
nand U18743 (N_18743,N_17596,N_17239);
nand U18744 (N_18744,N_17613,N_17824);
or U18745 (N_18745,N_17804,N_17802);
xor U18746 (N_18746,N_17852,N_17135);
and U18747 (N_18747,N_17211,N_17450);
nor U18748 (N_18748,N_16922,N_17435);
nand U18749 (N_18749,N_16830,N_17098);
and U18750 (N_18750,N_17223,N_17674);
nand U18751 (N_18751,N_16962,N_16964);
xor U18752 (N_18752,N_17494,N_17939);
and U18753 (N_18753,N_17761,N_17237);
nand U18754 (N_18754,N_17867,N_16973);
nor U18755 (N_18755,N_17893,N_17943);
and U18756 (N_18756,N_17052,N_17389);
and U18757 (N_18757,N_16908,N_17445);
nand U18758 (N_18758,N_17191,N_17877);
or U18759 (N_18759,N_17517,N_17436);
or U18760 (N_18760,N_17782,N_17130);
xor U18761 (N_18761,N_16932,N_16842);
xor U18762 (N_18762,N_17510,N_17122);
and U18763 (N_18763,N_17872,N_17610);
nand U18764 (N_18764,N_17563,N_17743);
nand U18765 (N_18765,N_17143,N_17584);
or U18766 (N_18766,N_17178,N_17543);
nand U18767 (N_18767,N_17494,N_17109);
or U18768 (N_18768,N_17513,N_17393);
xor U18769 (N_18769,N_16956,N_17761);
xor U18770 (N_18770,N_17244,N_17634);
or U18771 (N_18771,N_17184,N_17477);
xnor U18772 (N_18772,N_17028,N_17969);
xor U18773 (N_18773,N_17257,N_16809);
nor U18774 (N_18774,N_17801,N_17710);
and U18775 (N_18775,N_17205,N_17274);
nand U18776 (N_18776,N_17122,N_17393);
or U18777 (N_18777,N_17487,N_17491);
and U18778 (N_18778,N_16927,N_17661);
xor U18779 (N_18779,N_17849,N_16814);
or U18780 (N_18780,N_17119,N_16987);
nand U18781 (N_18781,N_16940,N_17903);
nor U18782 (N_18782,N_16990,N_16985);
or U18783 (N_18783,N_17012,N_17016);
or U18784 (N_18784,N_17576,N_16957);
nand U18785 (N_18785,N_17396,N_17793);
nand U18786 (N_18786,N_17757,N_17060);
and U18787 (N_18787,N_16980,N_17954);
nor U18788 (N_18788,N_17910,N_17857);
xor U18789 (N_18789,N_17298,N_17701);
nand U18790 (N_18790,N_17328,N_17456);
xor U18791 (N_18791,N_17505,N_16800);
or U18792 (N_18792,N_16931,N_17689);
nand U18793 (N_18793,N_17756,N_17361);
nor U18794 (N_18794,N_17489,N_17809);
nand U18795 (N_18795,N_17365,N_17420);
or U18796 (N_18796,N_17283,N_16969);
nor U18797 (N_18797,N_16954,N_17849);
and U18798 (N_18798,N_17448,N_16918);
nand U18799 (N_18799,N_17301,N_17928);
or U18800 (N_18800,N_17547,N_17360);
nand U18801 (N_18801,N_17191,N_17663);
or U18802 (N_18802,N_17893,N_17119);
or U18803 (N_18803,N_17638,N_17165);
nand U18804 (N_18804,N_17379,N_17204);
xnor U18805 (N_18805,N_17854,N_17609);
nand U18806 (N_18806,N_17638,N_17478);
and U18807 (N_18807,N_17220,N_17269);
or U18808 (N_18808,N_17681,N_17005);
nand U18809 (N_18809,N_16839,N_17528);
xor U18810 (N_18810,N_17232,N_17419);
nand U18811 (N_18811,N_17497,N_17750);
and U18812 (N_18812,N_17920,N_16831);
nor U18813 (N_18813,N_17668,N_16960);
or U18814 (N_18814,N_17945,N_17261);
or U18815 (N_18815,N_17850,N_17277);
nand U18816 (N_18816,N_17806,N_17702);
xor U18817 (N_18817,N_17443,N_17230);
nand U18818 (N_18818,N_17753,N_16899);
nand U18819 (N_18819,N_17892,N_17428);
xnor U18820 (N_18820,N_17688,N_16902);
nor U18821 (N_18821,N_16999,N_17811);
xor U18822 (N_18822,N_17121,N_17265);
or U18823 (N_18823,N_17766,N_16804);
and U18824 (N_18824,N_16917,N_17113);
nand U18825 (N_18825,N_16825,N_17750);
xor U18826 (N_18826,N_17225,N_17785);
nand U18827 (N_18827,N_17165,N_17854);
or U18828 (N_18828,N_17388,N_17758);
and U18829 (N_18829,N_17709,N_17909);
and U18830 (N_18830,N_17797,N_17021);
xnor U18831 (N_18831,N_17766,N_17017);
or U18832 (N_18832,N_17355,N_17700);
xor U18833 (N_18833,N_17738,N_17289);
and U18834 (N_18834,N_16819,N_17658);
nand U18835 (N_18835,N_16813,N_17394);
or U18836 (N_18836,N_17451,N_17128);
or U18837 (N_18837,N_17043,N_17977);
nor U18838 (N_18838,N_17698,N_17377);
and U18839 (N_18839,N_17652,N_17319);
and U18840 (N_18840,N_17510,N_16902);
nor U18841 (N_18841,N_17150,N_17492);
xnor U18842 (N_18842,N_16939,N_17568);
xor U18843 (N_18843,N_17632,N_17000);
and U18844 (N_18844,N_17219,N_16950);
xor U18845 (N_18845,N_17580,N_16970);
nor U18846 (N_18846,N_17485,N_16952);
nor U18847 (N_18847,N_17634,N_17444);
and U18848 (N_18848,N_16924,N_17368);
and U18849 (N_18849,N_17011,N_17281);
or U18850 (N_18850,N_17189,N_17922);
nand U18851 (N_18851,N_17365,N_17563);
nor U18852 (N_18852,N_17364,N_17624);
nand U18853 (N_18853,N_16860,N_17604);
nand U18854 (N_18854,N_17048,N_17337);
or U18855 (N_18855,N_17877,N_17677);
xnor U18856 (N_18856,N_17077,N_17547);
xnor U18857 (N_18857,N_17548,N_17443);
xnor U18858 (N_18858,N_17372,N_17725);
or U18859 (N_18859,N_16878,N_17551);
nor U18860 (N_18860,N_17827,N_16858);
xor U18861 (N_18861,N_17270,N_17776);
and U18862 (N_18862,N_17622,N_17876);
and U18863 (N_18863,N_17769,N_17304);
or U18864 (N_18864,N_16840,N_17390);
nand U18865 (N_18865,N_17144,N_16910);
xnor U18866 (N_18866,N_17180,N_17700);
or U18867 (N_18867,N_17022,N_17111);
or U18868 (N_18868,N_17922,N_17330);
and U18869 (N_18869,N_16894,N_16995);
nand U18870 (N_18870,N_17160,N_17610);
or U18871 (N_18871,N_17950,N_16969);
nand U18872 (N_18872,N_17488,N_17535);
nor U18873 (N_18873,N_17174,N_17522);
nor U18874 (N_18874,N_17449,N_17031);
xor U18875 (N_18875,N_17801,N_17053);
nand U18876 (N_18876,N_17204,N_17493);
nor U18877 (N_18877,N_17357,N_17530);
and U18878 (N_18878,N_17371,N_17609);
or U18879 (N_18879,N_16801,N_17691);
or U18880 (N_18880,N_17268,N_17970);
nand U18881 (N_18881,N_17294,N_17694);
or U18882 (N_18882,N_16908,N_17687);
nand U18883 (N_18883,N_17342,N_17716);
nor U18884 (N_18884,N_17947,N_16939);
and U18885 (N_18885,N_17465,N_17432);
xor U18886 (N_18886,N_17714,N_17414);
nor U18887 (N_18887,N_17172,N_17263);
xor U18888 (N_18888,N_17617,N_17484);
nand U18889 (N_18889,N_17919,N_17252);
nand U18890 (N_18890,N_17593,N_17803);
and U18891 (N_18891,N_17208,N_16861);
and U18892 (N_18892,N_17746,N_17870);
nand U18893 (N_18893,N_17494,N_17592);
xnor U18894 (N_18894,N_17091,N_17735);
nor U18895 (N_18895,N_16948,N_16839);
nor U18896 (N_18896,N_17043,N_17577);
and U18897 (N_18897,N_16910,N_17990);
or U18898 (N_18898,N_16819,N_17943);
and U18899 (N_18899,N_17574,N_16802);
xor U18900 (N_18900,N_17853,N_17951);
or U18901 (N_18901,N_17754,N_17602);
nand U18902 (N_18902,N_17357,N_17788);
or U18903 (N_18903,N_16852,N_17893);
xnor U18904 (N_18904,N_17494,N_17764);
or U18905 (N_18905,N_17613,N_17944);
or U18906 (N_18906,N_17228,N_16900);
and U18907 (N_18907,N_17505,N_17938);
and U18908 (N_18908,N_17729,N_17810);
and U18909 (N_18909,N_17060,N_17318);
and U18910 (N_18910,N_16853,N_17624);
and U18911 (N_18911,N_17663,N_17134);
nand U18912 (N_18912,N_17182,N_17682);
nand U18913 (N_18913,N_17456,N_17041);
nand U18914 (N_18914,N_17640,N_17015);
and U18915 (N_18915,N_17097,N_16836);
nor U18916 (N_18916,N_17645,N_17985);
and U18917 (N_18917,N_17612,N_17704);
and U18918 (N_18918,N_17338,N_17518);
and U18919 (N_18919,N_17377,N_16916);
or U18920 (N_18920,N_17586,N_17767);
and U18921 (N_18921,N_17774,N_17906);
or U18922 (N_18922,N_17638,N_17486);
and U18923 (N_18923,N_17383,N_17398);
and U18924 (N_18924,N_17354,N_17862);
xor U18925 (N_18925,N_17629,N_17590);
or U18926 (N_18926,N_17139,N_17582);
and U18927 (N_18927,N_17310,N_17461);
nand U18928 (N_18928,N_17638,N_17503);
nand U18929 (N_18929,N_17705,N_17631);
xor U18930 (N_18930,N_17064,N_17956);
xor U18931 (N_18931,N_17873,N_17298);
xnor U18932 (N_18932,N_17143,N_17639);
xnor U18933 (N_18933,N_17341,N_17128);
or U18934 (N_18934,N_17038,N_17258);
or U18935 (N_18935,N_17421,N_16896);
or U18936 (N_18936,N_17684,N_17146);
nand U18937 (N_18937,N_17857,N_16809);
or U18938 (N_18938,N_17095,N_17415);
and U18939 (N_18939,N_17591,N_17682);
xnor U18940 (N_18940,N_17832,N_17567);
xor U18941 (N_18941,N_17917,N_17304);
and U18942 (N_18942,N_17913,N_17609);
nor U18943 (N_18943,N_17562,N_17194);
nor U18944 (N_18944,N_16821,N_17007);
and U18945 (N_18945,N_17034,N_17588);
nand U18946 (N_18946,N_17380,N_17275);
nand U18947 (N_18947,N_17858,N_17552);
or U18948 (N_18948,N_17354,N_17965);
xor U18949 (N_18949,N_17971,N_17462);
nor U18950 (N_18950,N_16947,N_17904);
and U18951 (N_18951,N_17123,N_17649);
or U18952 (N_18952,N_17013,N_17666);
nor U18953 (N_18953,N_17301,N_17506);
or U18954 (N_18954,N_16863,N_17738);
nor U18955 (N_18955,N_17840,N_16907);
and U18956 (N_18956,N_17287,N_17110);
or U18957 (N_18957,N_16935,N_17598);
nor U18958 (N_18958,N_17194,N_17170);
nand U18959 (N_18959,N_17023,N_17521);
or U18960 (N_18960,N_17775,N_17949);
nor U18961 (N_18961,N_17653,N_17048);
nand U18962 (N_18962,N_17871,N_16878);
nand U18963 (N_18963,N_17394,N_17928);
nand U18964 (N_18964,N_17371,N_16989);
xor U18965 (N_18965,N_17874,N_17905);
xor U18966 (N_18966,N_16814,N_17965);
xor U18967 (N_18967,N_17719,N_17465);
or U18968 (N_18968,N_17816,N_16898);
xnor U18969 (N_18969,N_17208,N_17688);
or U18970 (N_18970,N_17068,N_17690);
nor U18971 (N_18971,N_17681,N_17751);
or U18972 (N_18972,N_17768,N_17042);
nand U18973 (N_18973,N_17267,N_17953);
or U18974 (N_18974,N_17551,N_16928);
nor U18975 (N_18975,N_17910,N_17532);
or U18976 (N_18976,N_17797,N_17772);
nand U18977 (N_18977,N_17095,N_16940);
nor U18978 (N_18978,N_17774,N_17519);
nand U18979 (N_18979,N_17313,N_17381);
xor U18980 (N_18980,N_17198,N_16827);
nand U18981 (N_18981,N_17144,N_16879);
xnor U18982 (N_18982,N_17645,N_17498);
xor U18983 (N_18983,N_17294,N_17654);
xnor U18984 (N_18984,N_16995,N_17395);
xor U18985 (N_18985,N_17827,N_17878);
nor U18986 (N_18986,N_17650,N_16963);
xnor U18987 (N_18987,N_16946,N_17359);
or U18988 (N_18988,N_17488,N_17887);
nand U18989 (N_18989,N_16824,N_17171);
nand U18990 (N_18990,N_17748,N_17350);
nor U18991 (N_18991,N_17911,N_16966);
or U18992 (N_18992,N_17655,N_17261);
and U18993 (N_18993,N_17985,N_17001);
and U18994 (N_18994,N_17207,N_16887);
and U18995 (N_18995,N_16834,N_17637);
nor U18996 (N_18996,N_16814,N_17174);
and U18997 (N_18997,N_17740,N_17654);
nor U18998 (N_18998,N_17354,N_17319);
xnor U18999 (N_18999,N_17188,N_16990);
nor U19000 (N_19000,N_17288,N_17078);
and U19001 (N_19001,N_17266,N_17129);
or U19002 (N_19002,N_17273,N_16987);
and U19003 (N_19003,N_17849,N_17178);
or U19004 (N_19004,N_17009,N_17556);
xnor U19005 (N_19005,N_17044,N_17474);
nand U19006 (N_19006,N_17297,N_17807);
nand U19007 (N_19007,N_17664,N_17312);
or U19008 (N_19008,N_17506,N_17746);
or U19009 (N_19009,N_16820,N_17659);
nor U19010 (N_19010,N_17307,N_16997);
nor U19011 (N_19011,N_17678,N_17616);
nand U19012 (N_19012,N_17935,N_17269);
or U19013 (N_19013,N_16842,N_16973);
nand U19014 (N_19014,N_17237,N_16852);
nand U19015 (N_19015,N_17639,N_17021);
or U19016 (N_19016,N_17513,N_17262);
xnor U19017 (N_19017,N_17735,N_16898);
or U19018 (N_19018,N_17088,N_17894);
nand U19019 (N_19019,N_17730,N_17476);
nor U19020 (N_19020,N_17568,N_17187);
and U19021 (N_19021,N_17367,N_17805);
nand U19022 (N_19022,N_16902,N_16942);
and U19023 (N_19023,N_17469,N_17785);
and U19024 (N_19024,N_17576,N_17765);
nand U19025 (N_19025,N_17122,N_17309);
or U19026 (N_19026,N_17213,N_17244);
xor U19027 (N_19027,N_17201,N_17827);
nand U19028 (N_19028,N_17240,N_17246);
and U19029 (N_19029,N_17801,N_17220);
nor U19030 (N_19030,N_17583,N_17318);
nand U19031 (N_19031,N_17845,N_17302);
nand U19032 (N_19032,N_17137,N_17353);
xor U19033 (N_19033,N_16908,N_17874);
xnor U19034 (N_19034,N_17094,N_17789);
nor U19035 (N_19035,N_17156,N_16952);
xnor U19036 (N_19036,N_17645,N_17032);
nand U19037 (N_19037,N_17121,N_16848);
nand U19038 (N_19038,N_17125,N_17285);
nor U19039 (N_19039,N_17589,N_17591);
nand U19040 (N_19040,N_17336,N_17559);
nand U19041 (N_19041,N_17258,N_17796);
nor U19042 (N_19042,N_17530,N_17824);
or U19043 (N_19043,N_16988,N_16866);
nor U19044 (N_19044,N_16901,N_17186);
nand U19045 (N_19045,N_17606,N_16877);
nand U19046 (N_19046,N_17411,N_17225);
nor U19047 (N_19047,N_17469,N_16950);
xnor U19048 (N_19048,N_17810,N_17508);
xnor U19049 (N_19049,N_17318,N_17194);
and U19050 (N_19050,N_17763,N_17282);
and U19051 (N_19051,N_17985,N_16977);
nand U19052 (N_19052,N_17040,N_16810);
nor U19053 (N_19053,N_17813,N_17007);
and U19054 (N_19054,N_16903,N_17385);
nor U19055 (N_19055,N_16850,N_17347);
xnor U19056 (N_19056,N_17978,N_17499);
nor U19057 (N_19057,N_17490,N_17925);
and U19058 (N_19058,N_16913,N_17365);
nand U19059 (N_19059,N_16804,N_17727);
and U19060 (N_19060,N_17625,N_17603);
xnor U19061 (N_19061,N_16913,N_17191);
or U19062 (N_19062,N_17988,N_17502);
nor U19063 (N_19063,N_17324,N_17692);
nand U19064 (N_19064,N_17367,N_17358);
and U19065 (N_19065,N_17195,N_17179);
nand U19066 (N_19066,N_16956,N_17906);
or U19067 (N_19067,N_17536,N_17973);
and U19068 (N_19068,N_17792,N_17383);
nand U19069 (N_19069,N_17090,N_17949);
and U19070 (N_19070,N_17823,N_16976);
or U19071 (N_19071,N_16877,N_17609);
and U19072 (N_19072,N_17322,N_17326);
nand U19073 (N_19073,N_17018,N_17851);
nand U19074 (N_19074,N_17105,N_17857);
xnor U19075 (N_19075,N_17764,N_17661);
nand U19076 (N_19076,N_17580,N_17552);
or U19077 (N_19077,N_17659,N_17475);
or U19078 (N_19078,N_17655,N_17638);
nor U19079 (N_19079,N_17227,N_17074);
xnor U19080 (N_19080,N_17206,N_17396);
and U19081 (N_19081,N_16937,N_17423);
or U19082 (N_19082,N_17493,N_17904);
xor U19083 (N_19083,N_17754,N_17798);
or U19084 (N_19084,N_17573,N_16835);
and U19085 (N_19085,N_17918,N_17710);
nand U19086 (N_19086,N_17610,N_17852);
or U19087 (N_19087,N_17090,N_16868);
or U19088 (N_19088,N_17640,N_16866);
nor U19089 (N_19089,N_17406,N_16881);
nand U19090 (N_19090,N_17560,N_17699);
and U19091 (N_19091,N_17535,N_17122);
and U19092 (N_19092,N_17257,N_16990);
nand U19093 (N_19093,N_17895,N_17194);
xnor U19094 (N_19094,N_17626,N_17953);
nand U19095 (N_19095,N_17695,N_17595);
xnor U19096 (N_19096,N_16992,N_17896);
xnor U19097 (N_19097,N_17359,N_17670);
xnor U19098 (N_19098,N_17674,N_17078);
nand U19099 (N_19099,N_17451,N_17531);
or U19100 (N_19100,N_17190,N_17298);
xnor U19101 (N_19101,N_17493,N_17276);
nand U19102 (N_19102,N_16818,N_17937);
nor U19103 (N_19103,N_17341,N_17427);
nand U19104 (N_19104,N_17270,N_16877);
nand U19105 (N_19105,N_17073,N_17777);
xnor U19106 (N_19106,N_17702,N_17152);
and U19107 (N_19107,N_17072,N_17493);
and U19108 (N_19108,N_17209,N_17733);
xnor U19109 (N_19109,N_17330,N_17387);
or U19110 (N_19110,N_17709,N_17800);
xnor U19111 (N_19111,N_17869,N_16872);
xor U19112 (N_19112,N_17289,N_17550);
nand U19113 (N_19113,N_17849,N_17976);
nand U19114 (N_19114,N_17182,N_17063);
xnor U19115 (N_19115,N_16976,N_17876);
nand U19116 (N_19116,N_17709,N_17827);
nand U19117 (N_19117,N_17639,N_16933);
and U19118 (N_19118,N_17046,N_16881);
or U19119 (N_19119,N_17754,N_17407);
nor U19120 (N_19120,N_17834,N_16930);
nor U19121 (N_19121,N_17465,N_16997);
xor U19122 (N_19122,N_17421,N_17658);
nor U19123 (N_19123,N_17042,N_17696);
xnor U19124 (N_19124,N_17175,N_17335);
nor U19125 (N_19125,N_17051,N_16889);
nand U19126 (N_19126,N_16921,N_17921);
nor U19127 (N_19127,N_17429,N_17545);
nand U19128 (N_19128,N_16943,N_17709);
nand U19129 (N_19129,N_16873,N_17073);
and U19130 (N_19130,N_17735,N_17720);
nor U19131 (N_19131,N_17057,N_17505);
or U19132 (N_19132,N_17545,N_17164);
nand U19133 (N_19133,N_16808,N_17857);
or U19134 (N_19134,N_17037,N_17620);
and U19135 (N_19135,N_17397,N_17085);
or U19136 (N_19136,N_17315,N_17110);
or U19137 (N_19137,N_17267,N_17495);
nand U19138 (N_19138,N_17675,N_17890);
nand U19139 (N_19139,N_17192,N_16896);
and U19140 (N_19140,N_17687,N_17471);
or U19141 (N_19141,N_17022,N_17702);
nor U19142 (N_19142,N_17942,N_17856);
nor U19143 (N_19143,N_17955,N_16913);
xnor U19144 (N_19144,N_17768,N_17285);
xnor U19145 (N_19145,N_17589,N_17620);
nand U19146 (N_19146,N_17647,N_17425);
nand U19147 (N_19147,N_16845,N_17359);
or U19148 (N_19148,N_17358,N_17185);
nor U19149 (N_19149,N_17420,N_17114);
nand U19150 (N_19150,N_17402,N_17643);
nor U19151 (N_19151,N_17072,N_16906);
nor U19152 (N_19152,N_17456,N_17263);
and U19153 (N_19153,N_17196,N_17632);
nand U19154 (N_19154,N_16954,N_17138);
or U19155 (N_19155,N_17530,N_17839);
nor U19156 (N_19156,N_17352,N_16928);
xnor U19157 (N_19157,N_17230,N_17709);
and U19158 (N_19158,N_17015,N_17515);
and U19159 (N_19159,N_17143,N_17734);
nand U19160 (N_19160,N_17190,N_17386);
nor U19161 (N_19161,N_17287,N_17261);
and U19162 (N_19162,N_17093,N_17327);
nand U19163 (N_19163,N_17322,N_17421);
and U19164 (N_19164,N_17358,N_17061);
or U19165 (N_19165,N_17912,N_17699);
or U19166 (N_19166,N_17532,N_17443);
xnor U19167 (N_19167,N_17477,N_17408);
nand U19168 (N_19168,N_17158,N_17243);
xor U19169 (N_19169,N_17519,N_17577);
and U19170 (N_19170,N_17027,N_17278);
xnor U19171 (N_19171,N_17729,N_17255);
xor U19172 (N_19172,N_17219,N_17598);
or U19173 (N_19173,N_16883,N_16870);
xor U19174 (N_19174,N_17136,N_16935);
nand U19175 (N_19175,N_17692,N_17352);
nand U19176 (N_19176,N_17824,N_17924);
nor U19177 (N_19177,N_17586,N_17229);
and U19178 (N_19178,N_17590,N_16998);
xnor U19179 (N_19179,N_17649,N_16933);
xor U19180 (N_19180,N_16973,N_17477);
nand U19181 (N_19181,N_17346,N_17771);
or U19182 (N_19182,N_17768,N_17399);
or U19183 (N_19183,N_17730,N_17287);
xor U19184 (N_19184,N_17288,N_17088);
or U19185 (N_19185,N_16839,N_17523);
nor U19186 (N_19186,N_17322,N_16943);
nand U19187 (N_19187,N_16923,N_17478);
and U19188 (N_19188,N_16892,N_17010);
nand U19189 (N_19189,N_17872,N_17846);
or U19190 (N_19190,N_16968,N_17561);
nand U19191 (N_19191,N_17774,N_17839);
and U19192 (N_19192,N_17459,N_17945);
nand U19193 (N_19193,N_17815,N_16809);
nand U19194 (N_19194,N_16984,N_16800);
nand U19195 (N_19195,N_17183,N_17712);
nand U19196 (N_19196,N_17809,N_16857);
or U19197 (N_19197,N_17154,N_17215);
or U19198 (N_19198,N_17279,N_17147);
and U19199 (N_19199,N_17378,N_17938);
nand U19200 (N_19200,N_19103,N_18813);
and U19201 (N_19201,N_18775,N_18200);
nor U19202 (N_19202,N_19097,N_18456);
and U19203 (N_19203,N_18249,N_18018);
nor U19204 (N_19204,N_18535,N_18133);
nand U19205 (N_19205,N_19095,N_18966);
or U19206 (N_19206,N_19140,N_19108);
nand U19207 (N_19207,N_18494,N_19154);
nand U19208 (N_19208,N_18783,N_18577);
xnor U19209 (N_19209,N_18284,N_18657);
nor U19210 (N_19210,N_19015,N_18526);
nand U19211 (N_19211,N_18585,N_18914);
xor U19212 (N_19212,N_18641,N_18916);
xor U19213 (N_19213,N_18727,N_18237);
nand U19214 (N_19214,N_18286,N_18685);
nand U19215 (N_19215,N_18501,N_19037);
nor U19216 (N_19216,N_18189,N_19033);
nor U19217 (N_19217,N_18077,N_18398);
and U19218 (N_19218,N_18959,N_18785);
or U19219 (N_19219,N_18755,N_18465);
nor U19220 (N_19220,N_18961,N_18873);
and U19221 (N_19221,N_19068,N_19001);
xor U19222 (N_19222,N_18661,N_18696);
nand U19223 (N_19223,N_19113,N_18055);
nor U19224 (N_19224,N_18253,N_18498);
nor U19225 (N_19225,N_19170,N_19142);
and U19226 (N_19226,N_18850,N_18404);
nor U19227 (N_19227,N_18593,N_18699);
nor U19228 (N_19228,N_18715,N_18514);
and U19229 (N_19229,N_18969,N_18680);
or U19230 (N_19230,N_18995,N_18683);
nor U19231 (N_19231,N_18230,N_18483);
xor U19232 (N_19232,N_19180,N_18104);
nor U19233 (N_19233,N_18938,N_18983);
or U19234 (N_19234,N_18626,N_18168);
or U19235 (N_19235,N_18220,N_18152);
nand U19236 (N_19236,N_18310,N_18158);
nor U19237 (N_19237,N_19036,N_19003);
xor U19238 (N_19238,N_18043,N_19058);
nor U19239 (N_19239,N_19199,N_18028);
nand U19240 (N_19240,N_19185,N_18438);
or U19241 (N_19241,N_19073,N_18853);
and U19242 (N_19242,N_18108,N_18663);
and U19243 (N_19243,N_18815,N_18917);
nand U19244 (N_19244,N_18072,N_18651);
nand U19245 (N_19245,N_19169,N_18433);
and U19246 (N_19246,N_18709,N_19105);
xor U19247 (N_19247,N_18892,N_18376);
nor U19248 (N_19248,N_18437,N_18215);
or U19249 (N_19249,N_18326,N_18106);
or U19250 (N_19250,N_18855,N_18321);
or U19251 (N_19251,N_18274,N_18466);
nand U19252 (N_19252,N_18265,N_18188);
nand U19253 (N_19253,N_18298,N_18455);
nand U19254 (N_19254,N_18163,N_18328);
xnor U19255 (N_19255,N_19125,N_18381);
xnor U19256 (N_19256,N_19178,N_19196);
and U19257 (N_19257,N_18777,N_18493);
nor U19258 (N_19258,N_18839,N_18830);
or U19259 (N_19259,N_18567,N_18036);
or U19260 (N_19260,N_18782,N_18954);
xor U19261 (N_19261,N_18009,N_18492);
nand U19262 (N_19262,N_18716,N_18377);
nor U19263 (N_19263,N_18902,N_18833);
nor U19264 (N_19264,N_19076,N_18659);
nand U19265 (N_19265,N_18093,N_18632);
nand U19266 (N_19266,N_18861,N_19006);
xor U19267 (N_19267,N_18978,N_19116);
nor U19268 (N_19268,N_18046,N_18471);
xor U19269 (N_19269,N_18788,N_18637);
xor U19270 (N_19270,N_19102,N_18633);
and U19271 (N_19271,N_18880,N_18197);
and U19272 (N_19272,N_18283,N_18473);
and U19273 (N_19273,N_19109,N_18330);
nand U19274 (N_19274,N_19048,N_18089);
xnor U19275 (N_19275,N_19043,N_18031);
and U19276 (N_19276,N_18900,N_19039);
nor U19277 (N_19277,N_18219,N_18135);
and U19278 (N_19278,N_19188,N_18458);
xnor U19279 (N_19279,N_18142,N_18828);
xor U19280 (N_19280,N_19115,N_18110);
nand U19281 (N_19281,N_18000,N_18267);
nand U19282 (N_19282,N_18134,N_18315);
nand U19283 (N_19283,N_18743,N_18226);
and U19284 (N_19284,N_18837,N_18533);
nor U19285 (N_19285,N_19072,N_18384);
nand U19286 (N_19286,N_18371,N_18705);
xor U19287 (N_19287,N_18216,N_18447);
nor U19288 (N_19288,N_18428,N_19078);
nand U19289 (N_19289,N_18446,N_18047);
nand U19290 (N_19290,N_18268,N_19163);
nand U19291 (N_19291,N_19069,N_18545);
nand U19292 (N_19292,N_19092,N_18453);
or U19293 (N_19293,N_18309,N_18085);
and U19294 (N_19294,N_18987,N_18757);
xnor U19295 (N_19295,N_18479,N_18392);
nor U19296 (N_19296,N_18347,N_18940);
and U19297 (N_19297,N_18957,N_18974);
and U19298 (N_19298,N_18736,N_18173);
or U19299 (N_19299,N_18746,N_18124);
or U19300 (N_19300,N_19182,N_18534);
and U19301 (N_19301,N_18930,N_18594);
or U19302 (N_19302,N_18962,N_18964);
or U19303 (N_19303,N_19002,N_18794);
nor U19304 (N_19304,N_18870,N_18649);
and U19305 (N_19305,N_18116,N_18920);
or U19306 (N_19306,N_18279,N_18883);
and U19307 (N_19307,N_19064,N_19009);
nor U19308 (N_19308,N_18178,N_18643);
or U19309 (N_19309,N_18067,N_18587);
or U19310 (N_19310,N_18337,N_19186);
nor U19311 (N_19311,N_18305,N_18574);
xnor U19312 (N_19312,N_18723,N_18350);
and U19313 (N_19313,N_18580,N_18712);
xor U19314 (N_19314,N_19047,N_18516);
nand U19315 (N_19315,N_18692,N_19138);
or U19316 (N_19316,N_19010,N_18035);
or U19317 (N_19317,N_18238,N_18767);
nand U19318 (N_19318,N_18729,N_18291);
xor U19319 (N_19319,N_18496,N_18431);
nor U19320 (N_19320,N_18477,N_18248);
xor U19321 (N_19321,N_18784,N_18896);
nor U19322 (N_19322,N_19106,N_18497);
nor U19323 (N_19323,N_18003,N_18597);
xnor U19324 (N_19324,N_18034,N_18327);
nand U19325 (N_19325,N_18734,N_18925);
or U19326 (N_19326,N_18354,N_18906);
nand U19327 (N_19327,N_18811,N_18943);
nor U19328 (N_19328,N_19152,N_18014);
nand U19329 (N_19329,N_18169,N_18988);
or U19330 (N_19330,N_18460,N_18285);
nor U19331 (N_19331,N_18251,N_18541);
or U19332 (N_19332,N_18203,N_19011);
xnor U19333 (N_19333,N_19066,N_19021);
xnor U19334 (N_19334,N_18138,N_18985);
nand U19335 (N_19335,N_18835,N_18807);
nand U19336 (N_19336,N_18667,N_19016);
xnor U19337 (N_19337,N_19181,N_18751);
nand U19338 (N_19338,N_18927,N_18418);
nand U19339 (N_19339,N_18139,N_18707);
and U19340 (N_19340,N_18847,N_18159);
or U19341 (N_19341,N_18419,N_18684);
and U19342 (N_19342,N_18143,N_18092);
or U19343 (N_19343,N_18128,N_18314);
or U19344 (N_19344,N_18980,N_19091);
nand U19345 (N_19345,N_18011,N_18592);
nor U19346 (N_19346,N_18366,N_19085);
and U19347 (N_19347,N_18505,N_18166);
nor U19348 (N_19348,N_18120,N_18700);
and U19349 (N_19349,N_18703,N_18955);
nand U19350 (N_19350,N_18866,N_18397);
xor U19351 (N_19351,N_18281,N_18878);
and U19352 (N_19352,N_18395,N_18806);
or U19353 (N_19353,N_18081,N_18903);
nor U19354 (N_19354,N_18464,N_18559);
and U19355 (N_19355,N_18161,N_18293);
or U19356 (N_19356,N_18472,N_18386);
xnor U19357 (N_19357,N_18517,N_18513);
xor U19358 (N_19358,N_18414,N_18631);
nand U19359 (N_19359,N_18656,N_18059);
or U19360 (N_19360,N_18886,N_19081);
and U19361 (N_19361,N_18240,N_18894);
xnor U19362 (N_19362,N_19045,N_18766);
or U19363 (N_19363,N_18524,N_19017);
and U19364 (N_19364,N_18311,N_18345);
nand U19365 (N_19365,N_19060,N_18838);
nor U19366 (N_19366,N_18801,N_18698);
xnor U19367 (N_19367,N_19027,N_18280);
and U19368 (N_19368,N_18679,N_18664);
nand U19369 (N_19369,N_18489,N_19136);
or U19370 (N_19370,N_18970,N_18167);
xnor U19371 (N_19371,N_18502,N_19122);
and U19372 (N_19372,N_18048,N_19179);
xnor U19373 (N_19373,N_18484,N_18565);
xnor U19374 (N_19374,N_18261,N_18302);
nand U19375 (N_19375,N_19114,N_18387);
xor U19376 (N_19376,N_19139,N_19054);
nor U19377 (N_19377,N_18671,N_18053);
and U19378 (N_19378,N_18074,N_18140);
and U19379 (N_19379,N_18208,N_18403);
or U19380 (N_19380,N_18851,N_18881);
nor U19381 (N_19381,N_18192,N_18439);
or U19382 (N_19382,N_18058,N_18681);
or U19383 (N_19383,N_18407,N_18951);
and U19384 (N_19384,N_18444,N_18171);
and U19385 (N_19385,N_18911,N_18107);
nor U19386 (N_19386,N_18589,N_18061);
nor U19387 (N_19387,N_18122,N_18101);
or U19388 (N_19388,N_18020,N_18441);
xor U19389 (N_19389,N_18029,N_18442);
and U19390 (N_19390,N_18854,N_18213);
and U19391 (N_19391,N_19146,N_18144);
xor U19392 (N_19392,N_19133,N_18629);
and U19393 (N_19393,N_19143,N_18972);
xor U19394 (N_19394,N_18979,N_18673);
nor U19395 (N_19395,N_18005,N_18724);
xnor U19396 (N_19396,N_18946,N_18542);
xnor U19397 (N_19397,N_18748,N_18634);
or U19398 (N_19398,N_18269,N_19023);
nor U19399 (N_19399,N_19013,N_18778);
nor U19400 (N_19400,N_18688,N_18976);
and U19401 (N_19401,N_19148,N_18195);
xnor U19402 (N_19402,N_18531,N_18223);
or U19403 (N_19403,N_18202,N_18997);
or U19404 (N_19404,N_18888,N_19187);
nor U19405 (N_19405,N_18764,N_18373);
or U19406 (N_19406,N_18155,N_19191);
and U19407 (N_19407,N_18153,N_18227);
nor U19408 (N_19408,N_18602,N_18319);
and U19409 (N_19409,N_18015,N_19065);
xnor U19410 (N_19410,N_18994,N_19135);
or U19411 (N_19411,N_18875,N_18992);
and U19412 (N_19412,N_19131,N_18620);
nand U19413 (N_19413,N_19034,N_18605);
or U19414 (N_19414,N_18065,N_18332);
nand U19415 (N_19415,N_19195,N_18409);
or U19416 (N_19416,N_18677,N_18079);
xnor U19417 (N_19417,N_18174,N_18868);
and U19418 (N_19418,N_18608,N_18741);
and U19419 (N_19419,N_18889,N_18747);
nor U19420 (N_19420,N_18480,N_18538);
nor U19421 (N_19421,N_18300,N_18389);
nor U19422 (N_19422,N_18521,N_18410);
and U19423 (N_19423,N_18432,N_19025);
and U19424 (N_19424,N_18753,N_18205);
or U19425 (N_19425,N_18926,N_18372);
or U19426 (N_19426,N_18086,N_18390);
and U19427 (N_19427,N_18207,N_19177);
nand U19428 (N_19428,N_18612,N_18999);
xnor U19429 (N_19429,N_18749,N_18733);
xnor U19430 (N_19430,N_18770,N_18162);
and U19431 (N_19431,N_18952,N_18278);
nor U19432 (N_19432,N_18325,N_18958);
nand U19433 (N_19433,N_18164,N_18495);
nor U19434 (N_19434,N_18735,N_18127);
and U19435 (N_19435,N_18790,N_18342);
and U19436 (N_19436,N_19050,N_18033);
xnor U19437 (N_19437,N_18359,N_18413);
nand U19438 (N_19438,N_18831,N_18858);
and U19439 (N_19439,N_18012,N_18027);
xnor U19440 (N_19440,N_19088,N_18179);
or U19441 (N_19441,N_18818,N_18040);
and U19442 (N_19442,N_18827,N_19168);
and U19443 (N_19443,N_18848,N_18119);
or U19444 (N_19444,N_18105,N_18897);
nor U19445 (N_19445,N_18975,N_19067);
or U19446 (N_19446,N_18187,N_19159);
or U19447 (N_19447,N_18662,N_18949);
or U19448 (N_19448,N_18774,N_18804);
xnor U19449 (N_19449,N_19038,N_18022);
and U19450 (N_19450,N_18343,N_18862);
nand U19451 (N_19451,N_19145,N_18242);
and U19452 (N_19452,N_19173,N_18504);
nand U19453 (N_19453,N_18379,N_19110);
nand U19454 (N_19454,N_18355,N_18125);
nor U19455 (N_19455,N_18401,N_18102);
or U19456 (N_19456,N_19007,N_18146);
nand U19457 (N_19457,N_18536,N_18623);
or U19458 (N_19458,N_18588,N_18360);
or U19459 (N_19459,N_18918,N_19161);
nand U19460 (N_19460,N_18841,N_18156);
or U19461 (N_19461,N_18845,N_18088);
or U19462 (N_19462,N_19087,N_18181);
nand U19463 (N_19463,N_18944,N_18071);
nor U19464 (N_19464,N_18935,N_18579);
nor U19465 (N_19465,N_18010,N_18895);
nor U19466 (N_19466,N_18287,N_18292);
xor U19467 (N_19467,N_18184,N_18448);
and U19468 (N_19468,N_18416,N_18443);
xnor U19469 (N_19469,N_18672,N_18898);
xor U19470 (N_19470,N_19190,N_18218);
or U19471 (N_19471,N_18313,N_19134);
and U19472 (N_19472,N_18056,N_18942);
and U19473 (N_19473,N_18511,N_18430);
xor U19474 (N_19474,N_19099,N_18998);
and U19475 (N_19475,N_18260,N_18212);
nor U19476 (N_19476,N_18126,N_18196);
and U19477 (N_19477,N_18400,N_18756);
nand U19478 (N_19478,N_18586,N_18396);
nor U19479 (N_19479,N_18924,N_18136);
xnor U19480 (N_19480,N_19014,N_18570);
nor U19481 (N_19481,N_19111,N_18475);
and U19482 (N_19482,N_18739,N_18947);
and U19483 (N_19483,N_19121,N_18154);
nand U19484 (N_19484,N_18083,N_18819);
nand U19485 (N_19485,N_18646,N_18021);
xor U19486 (N_19486,N_18129,N_19155);
xnor U19487 (N_19487,N_18348,N_18109);
and U19488 (N_19488,N_18091,N_19120);
and U19489 (N_19489,N_19100,N_18199);
xnor U19490 (N_19490,N_18795,N_18694);
xnor U19491 (N_19491,N_18039,N_18619);
or U19492 (N_19492,N_18320,N_18561);
xnor U19493 (N_19493,N_19057,N_18370);
or U19494 (N_19494,N_18262,N_18598);
nand U19495 (N_19495,N_18527,N_18984);
or U19496 (N_19496,N_18130,N_18094);
nand U19497 (N_19497,N_18434,N_19184);
xnor U19498 (N_19498,N_18993,N_18540);
or U19499 (N_19499,N_18457,N_18647);
xor U19500 (N_19500,N_18427,N_18754);
and U19501 (N_19501,N_19026,N_18301);
xor U19502 (N_19502,N_18004,N_18485);
or U19503 (N_19503,N_19162,N_18426);
or U19504 (N_19504,N_18702,N_18652);
nor U19505 (N_19505,N_18113,N_18805);
or U19506 (N_19506,N_18193,N_18779);
nand U19507 (N_19507,N_19123,N_18714);
and U19508 (N_19508,N_18335,N_18600);
nor U19509 (N_19509,N_18329,N_18668);
nand U19510 (N_19510,N_18429,N_18243);
nand U19511 (N_19511,N_18740,N_18568);
nand U19512 (N_19512,N_18628,N_18941);
nor U19513 (N_19513,N_18191,N_18204);
nor U19514 (N_19514,N_19193,N_18141);
and U19515 (N_19515,N_18933,N_18554);
nor U19516 (N_19516,N_18551,N_19128);
nand U19517 (N_19517,N_18422,N_18923);
nand U19518 (N_19518,N_18613,N_18254);
nand U19519 (N_19519,N_18147,N_18463);
nand U19520 (N_19520,N_18415,N_19056);
and U19521 (N_19521,N_18391,N_18050);
or U19522 (N_19522,N_18282,N_18915);
and U19523 (N_19523,N_18290,N_18640);
xor U19524 (N_19524,N_18417,N_18808);
nand U19525 (N_19525,N_18771,N_18864);
or U19526 (N_19526,N_19000,N_18564);
or U19527 (N_19527,N_18201,N_18383);
xor U19528 (N_19528,N_19004,N_18601);
or U19529 (N_19529,N_18257,N_18222);
xnor U19530 (N_19530,N_19096,N_19053);
nor U19531 (N_19531,N_18611,N_19077);
or U19532 (N_19532,N_18582,N_18233);
or U19533 (N_19533,N_18745,N_18338);
nor U19534 (N_19534,N_18803,N_19080);
and U19535 (N_19535,N_18500,N_18791);
and U19536 (N_19536,N_19028,N_18622);
nor U19537 (N_19537,N_18322,N_19063);
nand U19538 (N_19538,N_18185,N_18708);
or U19539 (N_19539,N_18731,N_18137);
or U19540 (N_19540,N_18175,N_19165);
xor U19541 (N_19541,N_18701,N_19062);
nor U19542 (N_19542,N_18859,N_19046);
nor U19543 (N_19543,N_18510,N_19059);
or U19544 (N_19544,N_18369,N_19167);
and U19545 (N_19545,N_18210,N_18636);
nor U19546 (N_19546,N_18451,N_18931);
xnor U19547 (N_19547,N_19192,N_18760);
xnor U19548 (N_19548,N_18863,N_18073);
and U19549 (N_19549,N_18800,N_19127);
nand U19550 (N_19550,N_18963,N_18644);
xnor U19551 (N_19551,N_18989,N_18068);
and U19552 (N_19552,N_18971,N_19150);
and U19553 (N_19553,N_18856,N_18362);
or U19554 (N_19554,N_18277,N_18045);
or U19555 (N_19555,N_18857,N_18973);
nand U19556 (N_19556,N_18236,N_18097);
xor U19557 (N_19557,N_18490,N_18645);
xor U19558 (N_19558,N_18177,N_18420);
and U19559 (N_19559,N_18810,N_18796);
xor U19560 (N_19560,N_18333,N_18530);
and U19561 (N_19561,N_18049,N_18732);
nand U19562 (N_19562,N_18548,N_18761);
or U19563 (N_19563,N_18340,N_18312);
nand U19564 (N_19564,N_18006,N_18607);
nand U19565 (N_19565,N_18722,N_18697);
nor U19566 (N_19566,N_19070,N_18515);
nand U19567 (N_19567,N_18406,N_18344);
or U19568 (N_19568,N_18872,N_18604);
nor U19569 (N_19569,N_18635,N_18306);
nor U19570 (N_19570,N_18007,N_18596);
nand U19571 (N_19571,N_19030,N_18445);
xor U19572 (N_19572,N_19147,N_18151);
xor U19573 (N_19573,N_18773,N_18725);
nand U19574 (N_19574,N_18666,N_19024);
xor U19575 (N_19575,N_19124,N_18507);
and U19576 (N_19576,N_18052,N_18730);
or U19577 (N_19577,N_18491,N_18317);
or U19578 (N_19578,N_19055,N_18423);
and U19579 (N_19579,N_18408,N_18132);
and U19580 (N_19580,N_18272,N_18625);
and U19581 (N_19581,N_18512,N_18578);
or U19582 (N_19582,N_18547,N_18799);
nand U19583 (N_19583,N_18241,N_19164);
or U19584 (N_19584,N_18270,N_18331);
or U19585 (N_19585,N_18225,N_18421);
nor U19586 (N_19586,N_19119,N_19035);
and U19587 (N_19587,N_18871,N_18318);
nor U19588 (N_19588,N_18539,N_18209);
or U19589 (N_19589,N_18103,N_19082);
nand U19590 (N_19590,N_18726,N_18563);
or U19591 (N_19591,N_18581,N_18402);
nor U19592 (N_19592,N_18678,N_18956);
and U19593 (N_19593,N_18520,N_18273);
xnor U19594 (N_19594,N_18616,N_18412);
nor U19595 (N_19595,N_18653,N_18440);
or U19596 (N_19596,N_18621,N_18967);
xor U19597 (N_19597,N_18648,N_18711);
or U19598 (N_19598,N_19012,N_18758);
and U19599 (N_19599,N_18537,N_19101);
and U19600 (N_19600,N_19022,N_18885);
or U19601 (N_19601,N_18070,N_19008);
or U19602 (N_19602,N_18436,N_18939);
and U19603 (N_19603,N_18584,N_18041);
and U19604 (N_19604,N_18614,N_18772);
xnor U19605 (N_19605,N_18303,N_18829);
nor U19606 (N_19606,N_18549,N_18675);
nand U19607 (N_19607,N_18781,N_18114);
xor U19608 (N_19608,N_18255,N_19094);
xor U19609 (N_19609,N_18710,N_19198);
or U19610 (N_19610,N_18590,N_18509);
and U19611 (N_19611,N_18288,N_18555);
and U19612 (N_19612,N_18001,N_18229);
nand U19613 (N_19613,N_18025,N_18096);
nor U19614 (N_19614,N_18349,N_18660);
and U19615 (N_19615,N_18468,N_18235);
nor U19616 (N_19616,N_19156,N_18160);
nand U19617 (N_19617,N_18953,N_18525);
xor U19618 (N_19618,N_19194,N_18738);
or U19619 (N_19619,N_18246,N_18172);
nor U19620 (N_19620,N_18353,N_18670);
nand U19621 (N_19621,N_19158,N_18150);
nor U19622 (N_19622,N_18720,N_18186);
or U19623 (N_19623,N_18913,N_18435);
and U19624 (N_19624,N_18907,N_18843);
nor U19625 (N_19625,N_18385,N_18481);
xor U19626 (N_19626,N_18111,N_18893);
or U19627 (N_19627,N_18658,N_18295);
xnor U19628 (N_19628,N_18965,N_18308);
and U19629 (N_19629,N_19032,N_18488);
and U19630 (N_19630,N_18522,N_18909);
nand U19631 (N_19631,N_18296,N_18532);
xnor U19632 (N_19632,N_18304,N_18276);
nand U19633 (N_19633,N_18252,N_18224);
xor U19634 (N_19634,N_18919,N_19098);
or U19635 (N_19635,N_18098,N_18546);
nand U19636 (N_19636,N_18454,N_18769);
nor U19637 (N_19637,N_18686,N_18380);
nor U19638 (N_19638,N_18183,N_18075);
nor U19639 (N_19639,N_18776,N_18339);
or U19640 (N_19640,N_18131,N_19197);
nand U19641 (N_19641,N_18609,N_18057);
nand U19642 (N_19642,N_18467,N_18575);
xnor U19643 (N_19643,N_18798,N_19144);
nand U19644 (N_19644,N_19189,N_18706);
nor U19645 (N_19645,N_19129,N_18316);
or U19646 (N_19646,N_19172,N_18836);
and U19647 (N_19647,N_18650,N_18695);
xnor U19648 (N_19648,N_18825,N_18411);
nor U19649 (N_19649,N_18874,N_18569);
xor U19650 (N_19650,N_18066,N_18228);
nand U19651 (N_19651,N_18948,N_18840);
nor U19652 (N_19652,N_18750,N_18610);
nor U19653 (N_19653,N_19183,N_18865);
nor U19654 (N_19654,N_18912,N_18910);
and U19655 (N_19655,N_18936,N_18363);
xnor U19656 (N_19656,N_18624,N_18786);
or U19657 (N_19657,N_18324,N_18069);
nor U19658 (N_19658,N_18690,N_18508);
or U19659 (N_19659,N_18562,N_18064);
and U19660 (N_19660,N_18713,N_18486);
nand U19661 (N_19661,N_19020,N_18573);
nor U19662 (N_19662,N_18117,N_19018);
nor U19663 (N_19663,N_19090,N_18932);
nor U19664 (N_19664,N_18506,N_18470);
nor U19665 (N_19665,N_18817,N_18263);
nand U19666 (N_19666,N_19176,N_18346);
and U19667 (N_19667,N_18780,N_18860);
or U19668 (N_19668,N_19171,N_18459);
nor U19669 (N_19669,N_18869,N_18388);
nand U19670 (N_19670,N_18182,N_18982);
nor U19671 (N_19671,N_18876,N_18639);
nand U19672 (N_19672,N_19019,N_18921);
xnor U19673 (N_19673,N_18595,N_18618);
or U19674 (N_19674,N_18642,N_18566);
or U19675 (N_19675,N_18019,N_18945);
xor U19676 (N_19676,N_18929,N_18449);
nand U19677 (N_19677,N_19149,N_18051);
or U19678 (N_19678,N_18908,N_18665);
nor U19679 (N_19679,N_18937,N_19093);
or U19680 (N_19680,N_18793,N_18572);
xor U19681 (N_19681,N_18452,N_18529);
nand U19682 (N_19682,N_18844,N_18968);
nor U19683 (N_19683,N_18336,N_18742);
nand U19684 (N_19684,N_19049,N_18478);
and U19685 (N_19685,N_18002,N_18239);
xor U19686 (N_19686,N_18294,N_18206);
nor U19687 (N_19687,N_18687,N_18519);
nand U19688 (N_19688,N_19126,N_18180);
and U19689 (N_19689,N_18100,N_18356);
or U19690 (N_19690,N_18042,N_18842);
and U19691 (N_19691,N_18121,N_18374);
nand U19692 (N_19692,N_18244,N_18543);
nand U19693 (N_19693,N_18060,N_18528);
nand U19694 (N_19694,N_18518,N_18832);
and U19695 (N_19695,N_18905,N_19117);
nor U19696 (N_19696,N_18038,N_18030);
and U19697 (N_19697,N_18368,N_18165);
or U19698 (N_19698,N_18655,N_18032);
or U19699 (N_19699,N_19112,N_18615);
nand U19700 (N_19700,N_18899,N_18405);
nand U19701 (N_19701,N_18476,N_19005);
xor U19702 (N_19702,N_18689,N_18960);
xor U19703 (N_19703,N_18789,N_18013);
nor U19704 (N_19704,N_18375,N_18591);
or U19705 (N_19705,N_18024,N_18087);
and U19706 (N_19706,N_18234,N_18928);
xor U19707 (N_19707,N_18271,N_18763);
and U19708 (N_19708,N_18812,N_18834);
or U19709 (N_19709,N_18078,N_18638);
and U19710 (N_19710,N_18214,N_18719);
and U19711 (N_19711,N_18095,N_18148);
and U19712 (N_19712,N_18289,N_18482);
nor U19713 (N_19713,N_19074,N_18461);
and U19714 (N_19714,N_19042,N_18630);
nor U19715 (N_19715,N_18090,N_18762);
nand U19716 (N_19716,N_19118,N_18654);
or U19717 (N_19717,N_19079,N_18231);
nand U19718 (N_19718,N_18361,N_18523);
or U19719 (N_19719,N_18487,N_18752);
xor U19720 (N_19720,N_18365,N_18849);
and U19721 (N_19721,N_18728,N_18768);
nand U19722 (N_19722,N_18721,N_18552);
and U19723 (N_19723,N_18682,N_18852);
xnor U19724 (N_19724,N_18082,N_19044);
nor U19725 (N_19725,N_19083,N_19052);
nor U19726 (N_19726,N_19137,N_18157);
xor U19727 (N_19727,N_18393,N_18922);
nor U19728 (N_19728,N_18358,N_18550);
nand U19729 (N_19729,N_18986,N_18822);
nand U19730 (N_19730,N_18826,N_18991);
nand U19731 (N_19731,N_18266,N_18737);
nor U19732 (N_19732,N_18990,N_18341);
and U19733 (N_19733,N_18217,N_18145);
nor U19734 (N_19734,N_18996,N_18044);
or U19735 (N_19735,N_18367,N_18334);
or U19736 (N_19736,N_18256,N_19075);
and U19737 (N_19737,N_18693,N_18016);
and U19738 (N_19738,N_18809,N_18323);
xnor U19739 (N_19739,N_18364,N_18797);
nand U19740 (N_19740,N_19104,N_18378);
nand U19741 (N_19741,N_18887,N_18583);
or U19742 (N_19742,N_18558,N_18669);
nor U19743 (N_19743,N_19084,N_18264);
nor U19744 (N_19744,N_18823,N_18394);
nor U19745 (N_19745,N_18882,N_18977);
and U19746 (N_19746,N_18557,N_18792);
and U19747 (N_19747,N_18824,N_18821);
and U19748 (N_19748,N_18099,N_19151);
nor U19749 (N_19749,N_18802,N_19166);
nor U19750 (N_19750,N_18718,N_18425);
nor U19751 (N_19751,N_19160,N_19132);
nor U19752 (N_19752,N_18877,N_19031);
nand U19753 (N_19753,N_18704,N_18867);
or U19754 (N_19754,N_18576,N_18080);
and U19755 (N_19755,N_18176,N_19130);
or U19756 (N_19756,N_18307,N_18063);
and U19757 (N_19757,N_18627,N_18950);
and U19758 (N_19758,N_18717,N_18054);
nor U19759 (N_19759,N_18846,N_18245);
nor U19760 (N_19760,N_18211,N_18115);
or U19761 (N_19761,N_18553,N_18462);
and U19762 (N_19762,N_18499,N_18275);
xnor U19763 (N_19763,N_18297,N_18062);
nand U19764 (N_19764,N_18076,N_18424);
and U19765 (N_19765,N_19141,N_18879);
and U19766 (N_19766,N_18820,N_18232);
or U19767 (N_19767,N_18891,N_18676);
nor U19768 (N_19768,N_19174,N_19041);
xor U19769 (N_19769,N_18674,N_18221);
nand U19770 (N_19770,N_19157,N_18503);
nor U19771 (N_19771,N_19040,N_18259);
xor U19772 (N_19772,N_18560,N_19153);
or U19773 (N_19773,N_18901,N_18450);
and U19774 (N_19774,N_19051,N_19089);
and U19775 (N_19775,N_18544,N_18981);
xnor U19776 (N_19776,N_18765,N_18190);
or U19777 (N_19777,N_18556,N_18934);
nand U19778 (N_19778,N_18814,N_18258);
or U19779 (N_19779,N_18787,N_19086);
or U19780 (N_19780,N_18691,N_18357);
nor U19781 (N_19781,N_18149,N_18194);
or U19782 (N_19782,N_18037,N_18816);
xor U19783 (N_19783,N_18118,N_18351);
xor U19784 (N_19784,N_18023,N_18112);
nand U19785 (N_19785,N_19061,N_19071);
xor U19786 (N_19786,N_19107,N_18744);
xor U19787 (N_19787,N_18382,N_18299);
nand U19788 (N_19788,N_18198,N_18606);
nand U19789 (N_19789,N_19029,N_18469);
xor U19790 (N_19790,N_18399,N_18026);
and U19791 (N_19791,N_18250,N_18474);
nand U19792 (N_19792,N_18603,N_18571);
xor U19793 (N_19793,N_18759,N_18084);
and U19794 (N_19794,N_18599,N_18123);
xor U19795 (N_19795,N_18890,N_18904);
or U19796 (N_19796,N_18352,N_18247);
xor U19797 (N_19797,N_18884,N_18008);
nand U19798 (N_19798,N_18017,N_18170);
nor U19799 (N_19799,N_18617,N_19175);
and U19800 (N_19800,N_18673,N_18517);
xnor U19801 (N_19801,N_18902,N_18585);
or U19802 (N_19802,N_18015,N_18809);
or U19803 (N_19803,N_18062,N_18324);
nor U19804 (N_19804,N_18318,N_18825);
and U19805 (N_19805,N_18660,N_18580);
xnor U19806 (N_19806,N_18539,N_18096);
xor U19807 (N_19807,N_18087,N_19081);
and U19808 (N_19808,N_18988,N_18825);
or U19809 (N_19809,N_18513,N_18395);
xor U19810 (N_19810,N_18115,N_18341);
nand U19811 (N_19811,N_18171,N_18564);
xnor U19812 (N_19812,N_18303,N_18340);
nand U19813 (N_19813,N_18517,N_18236);
xor U19814 (N_19814,N_18089,N_19165);
nor U19815 (N_19815,N_18455,N_18211);
nor U19816 (N_19816,N_19054,N_18397);
xor U19817 (N_19817,N_19092,N_18730);
and U19818 (N_19818,N_18452,N_18545);
nand U19819 (N_19819,N_18977,N_18756);
and U19820 (N_19820,N_19146,N_18451);
or U19821 (N_19821,N_18907,N_18867);
xor U19822 (N_19822,N_19082,N_18004);
or U19823 (N_19823,N_19026,N_18350);
nor U19824 (N_19824,N_18976,N_18738);
xnor U19825 (N_19825,N_18283,N_18747);
and U19826 (N_19826,N_18647,N_18552);
nand U19827 (N_19827,N_18488,N_18079);
xor U19828 (N_19828,N_18148,N_18777);
nand U19829 (N_19829,N_18873,N_18230);
xnor U19830 (N_19830,N_18686,N_18694);
nor U19831 (N_19831,N_18446,N_18708);
or U19832 (N_19832,N_18065,N_18126);
nor U19833 (N_19833,N_18159,N_18357);
nand U19834 (N_19834,N_18308,N_19016);
and U19835 (N_19835,N_18862,N_19056);
and U19836 (N_19836,N_18164,N_18971);
and U19837 (N_19837,N_18269,N_19183);
and U19838 (N_19838,N_18853,N_18298);
or U19839 (N_19839,N_19043,N_19031);
nor U19840 (N_19840,N_18337,N_18954);
and U19841 (N_19841,N_18205,N_18664);
nand U19842 (N_19842,N_19023,N_18341);
and U19843 (N_19843,N_18224,N_18209);
or U19844 (N_19844,N_18949,N_18600);
or U19845 (N_19845,N_18815,N_19096);
or U19846 (N_19846,N_19163,N_18713);
nand U19847 (N_19847,N_18607,N_18295);
and U19848 (N_19848,N_18094,N_18167);
nand U19849 (N_19849,N_18007,N_19103);
and U19850 (N_19850,N_18949,N_18697);
xnor U19851 (N_19851,N_18014,N_18416);
xnor U19852 (N_19852,N_18179,N_18562);
or U19853 (N_19853,N_19003,N_18055);
or U19854 (N_19854,N_18061,N_18936);
or U19855 (N_19855,N_18875,N_19072);
or U19856 (N_19856,N_18470,N_18439);
xor U19857 (N_19857,N_19190,N_18820);
and U19858 (N_19858,N_18864,N_19006);
nor U19859 (N_19859,N_18501,N_19084);
xnor U19860 (N_19860,N_18955,N_18849);
and U19861 (N_19861,N_18656,N_18982);
xor U19862 (N_19862,N_18748,N_19152);
xor U19863 (N_19863,N_18598,N_18657);
or U19864 (N_19864,N_19174,N_18143);
nand U19865 (N_19865,N_18578,N_18300);
and U19866 (N_19866,N_18905,N_18760);
xnor U19867 (N_19867,N_18188,N_19076);
nor U19868 (N_19868,N_18331,N_19060);
xnor U19869 (N_19869,N_19013,N_18114);
xnor U19870 (N_19870,N_18666,N_18408);
nor U19871 (N_19871,N_18236,N_18079);
nor U19872 (N_19872,N_18907,N_18896);
or U19873 (N_19873,N_18413,N_18021);
nand U19874 (N_19874,N_19074,N_18327);
xor U19875 (N_19875,N_18412,N_18081);
or U19876 (N_19876,N_19076,N_18332);
xnor U19877 (N_19877,N_18694,N_18611);
nand U19878 (N_19878,N_18745,N_18070);
and U19879 (N_19879,N_18645,N_18763);
xnor U19880 (N_19880,N_18425,N_18264);
nand U19881 (N_19881,N_18120,N_18145);
and U19882 (N_19882,N_18622,N_18280);
nand U19883 (N_19883,N_18238,N_18394);
nor U19884 (N_19884,N_19093,N_18569);
or U19885 (N_19885,N_18940,N_18301);
xnor U19886 (N_19886,N_18678,N_19178);
and U19887 (N_19887,N_18231,N_18402);
nand U19888 (N_19888,N_18316,N_18081);
and U19889 (N_19889,N_18518,N_18341);
nor U19890 (N_19890,N_18017,N_18763);
nor U19891 (N_19891,N_18356,N_18965);
nand U19892 (N_19892,N_18177,N_18961);
or U19893 (N_19893,N_18157,N_18648);
nand U19894 (N_19894,N_18756,N_18669);
xnor U19895 (N_19895,N_18435,N_18968);
or U19896 (N_19896,N_18894,N_18435);
xnor U19897 (N_19897,N_19194,N_18579);
or U19898 (N_19898,N_18147,N_18013);
and U19899 (N_19899,N_18978,N_19126);
or U19900 (N_19900,N_18102,N_18498);
nor U19901 (N_19901,N_18212,N_18662);
nor U19902 (N_19902,N_18377,N_18712);
nor U19903 (N_19903,N_18049,N_18647);
nor U19904 (N_19904,N_18758,N_18089);
nand U19905 (N_19905,N_18410,N_18859);
nor U19906 (N_19906,N_18024,N_18347);
or U19907 (N_19907,N_18631,N_18820);
nor U19908 (N_19908,N_18296,N_18408);
xor U19909 (N_19909,N_18286,N_18262);
or U19910 (N_19910,N_18151,N_19187);
or U19911 (N_19911,N_18250,N_19063);
and U19912 (N_19912,N_18404,N_18871);
nor U19913 (N_19913,N_18504,N_18958);
or U19914 (N_19914,N_19062,N_18127);
xnor U19915 (N_19915,N_18497,N_18038);
or U19916 (N_19916,N_18481,N_18471);
or U19917 (N_19917,N_18218,N_18691);
or U19918 (N_19918,N_18397,N_18538);
nor U19919 (N_19919,N_19176,N_18821);
xor U19920 (N_19920,N_18815,N_18695);
nor U19921 (N_19921,N_18971,N_19124);
nand U19922 (N_19922,N_18828,N_18353);
and U19923 (N_19923,N_18511,N_18984);
nand U19924 (N_19924,N_19191,N_18276);
or U19925 (N_19925,N_18755,N_18731);
nand U19926 (N_19926,N_18225,N_18527);
xor U19927 (N_19927,N_18181,N_18433);
nor U19928 (N_19928,N_19154,N_18169);
xnor U19929 (N_19929,N_19101,N_18504);
or U19930 (N_19930,N_18673,N_18509);
nor U19931 (N_19931,N_18017,N_18357);
nand U19932 (N_19932,N_18407,N_19079);
nand U19933 (N_19933,N_18476,N_18546);
nand U19934 (N_19934,N_18759,N_18563);
nand U19935 (N_19935,N_18853,N_18005);
or U19936 (N_19936,N_18227,N_18068);
nand U19937 (N_19937,N_18198,N_18364);
nand U19938 (N_19938,N_18504,N_18967);
xnor U19939 (N_19939,N_19115,N_18843);
or U19940 (N_19940,N_19170,N_18789);
xnor U19941 (N_19941,N_18353,N_18329);
nor U19942 (N_19942,N_18560,N_18820);
xnor U19943 (N_19943,N_18348,N_18144);
and U19944 (N_19944,N_19116,N_18489);
xor U19945 (N_19945,N_19088,N_19075);
nand U19946 (N_19946,N_19023,N_18897);
xnor U19947 (N_19947,N_19155,N_19113);
nand U19948 (N_19948,N_18805,N_18659);
and U19949 (N_19949,N_19188,N_18083);
xor U19950 (N_19950,N_19118,N_19102);
nor U19951 (N_19951,N_18215,N_18207);
nand U19952 (N_19952,N_18417,N_19114);
or U19953 (N_19953,N_19197,N_19175);
nor U19954 (N_19954,N_18984,N_18364);
nand U19955 (N_19955,N_18331,N_18236);
or U19956 (N_19956,N_18011,N_19088);
or U19957 (N_19957,N_18153,N_18872);
nor U19958 (N_19958,N_18791,N_18244);
or U19959 (N_19959,N_19037,N_18491);
and U19960 (N_19960,N_18561,N_18108);
nor U19961 (N_19961,N_18816,N_18307);
or U19962 (N_19962,N_18024,N_18597);
nor U19963 (N_19963,N_18938,N_18007);
nand U19964 (N_19964,N_18264,N_18099);
nand U19965 (N_19965,N_18620,N_18418);
xnor U19966 (N_19966,N_18091,N_18074);
or U19967 (N_19967,N_18037,N_18722);
xnor U19968 (N_19968,N_18770,N_18695);
and U19969 (N_19969,N_18110,N_18408);
xor U19970 (N_19970,N_18736,N_18375);
xor U19971 (N_19971,N_18925,N_19012);
or U19972 (N_19972,N_18218,N_19109);
nor U19973 (N_19973,N_18617,N_18221);
xor U19974 (N_19974,N_18616,N_18921);
and U19975 (N_19975,N_18836,N_18556);
xnor U19976 (N_19976,N_18486,N_18740);
nand U19977 (N_19977,N_18338,N_18709);
or U19978 (N_19978,N_18534,N_18510);
nor U19979 (N_19979,N_18781,N_18043);
and U19980 (N_19980,N_18608,N_19090);
or U19981 (N_19981,N_18111,N_18823);
xnor U19982 (N_19982,N_19080,N_18698);
or U19983 (N_19983,N_19125,N_18480);
and U19984 (N_19984,N_18638,N_18487);
or U19985 (N_19985,N_18295,N_18464);
and U19986 (N_19986,N_18438,N_18101);
nor U19987 (N_19987,N_18532,N_19062);
nor U19988 (N_19988,N_18351,N_18404);
nand U19989 (N_19989,N_18882,N_18903);
and U19990 (N_19990,N_19161,N_19057);
xor U19991 (N_19991,N_18097,N_18276);
nor U19992 (N_19992,N_19157,N_19195);
and U19993 (N_19993,N_18340,N_18118);
nor U19994 (N_19994,N_19165,N_19128);
nand U19995 (N_19995,N_18655,N_18736);
xor U19996 (N_19996,N_18921,N_18314);
and U19997 (N_19997,N_18053,N_18892);
nor U19998 (N_19998,N_18148,N_18604);
and U19999 (N_19999,N_18734,N_18163);
xor U20000 (N_20000,N_18287,N_18401);
nor U20001 (N_20001,N_19128,N_18483);
nand U20002 (N_20002,N_18803,N_19150);
and U20003 (N_20003,N_18729,N_19051);
and U20004 (N_20004,N_18001,N_18522);
xnor U20005 (N_20005,N_18697,N_18340);
xnor U20006 (N_20006,N_18951,N_18712);
nand U20007 (N_20007,N_18579,N_18581);
and U20008 (N_20008,N_18632,N_18625);
or U20009 (N_20009,N_18811,N_18587);
and U20010 (N_20010,N_18500,N_18161);
and U20011 (N_20011,N_18831,N_18662);
nor U20012 (N_20012,N_18530,N_18214);
and U20013 (N_20013,N_18358,N_18341);
nor U20014 (N_20014,N_18653,N_19113);
xor U20015 (N_20015,N_18428,N_18623);
or U20016 (N_20016,N_18185,N_18749);
nor U20017 (N_20017,N_18541,N_18764);
and U20018 (N_20018,N_18326,N_18339);
and U20019 (N_20019,N_18885,N_19164);
nor U20020 (N_20020,N_18283,N_18587);
or U20021 (N_20021,N_18438,N_18838);
nor U20022 (N_20022,N_18721,N_19118);
nand U20023 (N_20023,N_18744,N_19134);
nor U20024 (N_20024,N_18533,N_18444);
or U20025 (N_20025,N_18829,N_18559);
xor U20026 (N_20026,N_18511,N_18423);
nor U20027 (N_20027,N_18663,N_18147);
and U20028 (N_20028,N_18099,N_18035);
nand U20029 (N_20029,N_18796,N_18365);
nand U20030 (N_20030,N_18281,N_18662);
nand U20031 (N_20031,N_18619,N_18320);
or U20032 (N_20032,N_18491,N_18809);
and U20033 (N_20033,N_18407,N_18157);
and U20034 (N_20034,N_18777,N_18097);
nor U20035 (N_20035,N_18548,N_18279);
and U20036 (N_20036,N_18802,N_18458);
nor U20037 (N_20037,N_18119,N_18157);
xnor U20038 (N_20038,N_18766,N_18394);
nor U20039 (N_20039,N_18922,N_18284);
xor U20040 (N_20040,N_18698,N_18630);
nand U20041 (N_20041,N_18039,N_18461);
nor U20042 (N_20042,N_18381,N_18876);
nor U20043 (N_20043,N_18236,N_18661);
and U20044 (N_20044,N_18193,N_19110);
or U20045 (N_20045,N_18148,N_18368);
nand U20046 (N_20046,N_18162,N_18868);
and U20047 (N_20047,N_18365,N_18130);
nand U20048 (N_20048,N_18286,N_18939);
xor U20049 (N_20049,N_18622,N_18472);
or U20050 (N_20050,N_18406,N_18166);
xor U20051 (N_20051,N_18078,N_18225);
xor U20052 (N_20052,N_18411,N_18052);
or U20053 (N_20053,N_18332,N_18787);
and U20054 (N_20054,N_18802,N_18187);
nand U20055 (N_20055,N_18622,N_19070);
nor U20056 (N_20056,N_18138,N_18715);
nand U20057 (N_20057,N_18322,N_18787);
nor U20058 (N_20058,N_18815,N_18310);
and U20059 (N_20059,N_18828,N_19010);
or U20060 (N_20060,N_19025,N_18282);
nand U20061 (N_20061,N_18701,N_18936);
xnor U20062 (N_20062,N_18190,N_18163);
and U20063 (N_20063,N_18312,N_18500);
or U20064 (N_20064,N_18491,N_18434);
and U20065 (N_20065,N_18768,N_18515);
or U20066 (N_20066,N_18870,N_18537);
xnor U20067 (N_20067,N_18220,N_18415);
or U20068 (N_20068,N_18802,N_18388);
xor U20069 (N_20069,N_18941,N_18936);
or U20070 (N_20070,N_19118,N_18807);
or U20071 (N_20071,N_18303,N_19042);
or U20072 (N_20072,N_19036,N_19073);
and U20073 (N_20073,N_19144,N_19047);
or U20074 (N_20074,N_18574,N_18430);
xnor U20075 (N_20075,N_18055,N_18625);
and U20076 (N_20076,N_19100,N_18794);
nor U20077 (N_20077,N_18082,N_18323);
nand U20078 (N_20078,N_18267,N_18002);
and U20079 (N_20079,N_18541,N_18530);
nand U20080 (N_20080,N_18054,N_19186);
nor U20081 (N_20081,N_18443,N_18782);
xor U20082 (N_20082,N_18484,N_18745);
or U20083 (N_20083,N_18919,N_18481);
xor U20084 (N_20084,N_18675,N_18755);
nor U20085 (N_20085,N_18814,N_18731);
and U20086 (N_20086,N_18049,N_18423);
nand U20087 (N_20087,N_19004,N_18610);
nor U20088 (N_20088,N_18656,N_18965);
xor U20089 (N_20089,N_18226,N_18353);
xnor U20090 (N_20090,N_18556,N_18579);
or U20091 (N_20091,N_18809,N_18778);
nor U20092 (N_20092,N_18414,N_18682);
nor U20093 (N_20093,N_19114,N_18839);
or U20094 (N_20094,N_18890,N_19112);
and U20095 (N_20095,N_18506,N_18026);
nor U20096 (N_20096,N_19194,N_18648);
xnor U20097 (N_20097,N_18406,N_18695);
xor U20098 (N_20098,N_18319,N_19042);
nand U20099 (N_20099,N_18109,N_18192);
or U20100 (N_20100,N_18700,N_18969);
and U20101 (N_20101,N_18758,N_18136);
nand U20102 (N_20102,N_18658,N_18729);
nand U20103 (N_20103,N_18267,N_18780);
nand U20104 (N_20104,N_18707,N_18915);
nand U20105 (N_20105,N_18881,N_18068);
nand U20106 (N_20106,N_18353,N_18367);
nor U20107 (N_20107,N_18155,N_18567);
or U20108 (N_20108,N_18196,N_18920);
and U20109 (N_20109,N_18911,N_18492);
nand U20110 (N_20110,N_18629,N_18131);
nor U20111 (N_20111,N_18363,N_18065);
or U20112 (N_20112,N_18685,N_19078);
or U20113 (N_20113,N_18591,N_18561);
nor U20114 (N_20114,N_18805,N_18369);
xnor U20115 (N_20115,N_18017,N_18397);
and U20116 (N_20116,N_18529,N_18439);
nor U20117 (N_20117,N_18587,N_18984);
nor U20118 (N_20118,N_18274,N_18093);
nand U20119 (N_20119,N_18791,N_18845);
or U20120 (N_20120,N_18788,N_18210);
nand U20121 (N_20121,N_18080,N_18771);
nand U20122 (N_20122,N_18580,N_18716);
xnor U20123 (N_20123,N_18730,N_18244);
nand U20124 (N_20124,N_18548,N_18448);
xnor U20125 (N_20125,N_18076,N_18259);
and U20126 (N_20126,N_18637,N_19041);
or U20127 (N_20127,N_18214,N_18731);
nand U20128 (N_20128,N_18696,N_18643);
nor U20129 (N_20129,N_18407,N_18473);
xnor U20130 (N_20130,N_18954,N_19050);
xor U20131 (N_20131,N_18855,N_18728);
and U20132 (N_20132,N_18211,N_18777);
nand U20133 (N_20133,N_18259,N_18304);
nor U20134 (N_20134,N_18322,N_18244);
or U20135 (N_20135,N_18998,N_18195);
nand U20136 (N_20136,N_18022,N_18852);
or U20137 (N_20137,N_18444,N_18008);
xor U20138 (N_20138,N_18958,N_18524);
and U20139 (N_20139,N_18903,N_18957);
nor U20140 (N_20140,N_18031,N_18873);
xor U20141 (N_20141,N_18157,N_18670);
and U20142 (N_20142,N_18958,N_18185);
nor U20143 (N_20143,N_18513,N_18255);
nand U20144 (N_20144,N_18404,N_18406);
or U20145 (N_20145,N_18165,N_19056);
or U20146 (N_20146,N_18545,N_18830);
nor U20147 (N_20147,N_19199,N_19030);
and U20148 (N_20148,N_18883,N_18531);
or U20149 (N_20149,N_18636,N_18913);
nand U20150 (N_20150,N_18619,N_18844);
and U20151 (N_20151,N_18750,N_18110);
nor U20152 (N_20152,N_19157,N_18167);
xnor U20153 (N_20153,N_18019,N_18477);
and U20154 (N_20154,N_18908,N_18363);
nor U20155 (N_20155,N_19068,N_19091);
xnor U20156 (N_20156,N_18391,N_18801);
nor U20157 (N_20157,N_18267,N_18071);
xnor U20158 (N_20158,N_18395,N_18549);
nand U20159 (N_20159,N_18761,N_18574);
xnor U20160 (N_20160,N_18801,N_18159);
nand U20161 (N_20161,N_18135,N_18337);
nand U20162 (N_20162,N_18232,N_18480);
and U20163 (N_20163,N_19108,N_18795);
nand U20164 (N_20164,N_18293,N_19060);
nor U20165 (N_20165,N_18916,N_18430);
xnor U20166 (N_20166,N_18447,N_18883);
nor U20167 (N_20167,N_18309,N_18998);
xnor U20168 (N_20168,N_18733,N_18582);
and U20169 (N_20169,N_18254,N_18499);
or U20170 (N_20170,N_18522,N_18831);
nand U20171 (N_20171,N_18018,N_18836);
nand U20172 (N_20172,N_18572,N_19042);
and U20173 (N_20173,N_18763,N_18536);
xnor U20174 (N_20174,N_19004,N_18868);
and U20175 (N_20175,N_18580,N_19110);
nor U20176 (N_20176,N_18759,N_18637);
and U20177 (N_20177,N_18504,N_18202);
and U20178 (N_20178,N_18847,N_18587);
or U20179 (N_20179,N_19078,N_18636);
xor U20180 (N_20180,N_18518,N_19073);
xnor U20181 (N_20181,N_18700,N_18539);
nand U20182 (N_20182,N_18931,N_18830);
or U20183 (N_20183,N_19069,N_18386);
and U20184 (N_20184,N_18049,N_18565);
nand U20185 (N_20185,N_18222,N_18910);
or U20186 (N_20186,N_18342,N_19196);
nand U20187 (N_20187,N_19177,N_18192);
nand U20188 (N_20188,N_18008,N_18957);
or U20189 (N_20189,N_18574,N_18942);
or U20190 (N_20190,N_18975,N_18276);
xnor U20191 (N_20191,N_18244,N_18819);
or U20192 (N_20192,N_19178,N_18685);
and U20193 (N_20193,N_18410,N_18533);
xnor U20194 (N_20194,N_18943,N_18601);
and U20195 (N_20195,N_18698,N_19190);
xnor U20196 (N_20196,N_18080,N_18418);
and U20197 (N_20197,N_18741,N_18133);
and U20198 (N_20198,N_19152,N_18974);
or U20199 (N_20199,N_18589,N_18184);
xor U20200 (N_20200,N_18517,N_18939);
nor U20201 (N_20201,N_18453,N_18721);
and U20202 (N_20202,N_18004,N_18827);
and U20203 (N_20203,N_18719,N_18869);
xor U20204 (N_20204,N_18192,N_18847);
nand U20205 (N_20205,N_18159,N_18664);
and U20206 (N_20206,N_19125,N_18478);
xnor U20207 (N_20207,N_18062,N_18162);
or U20208 (N_20208,N_19080,N_19038);
and U20209 (N_20209,N_18511,N_19173);
or U20210 (N_20210,N_18332,N_19141);
nor U20211 (N_20211,N_18566,N_18320);
nor U20212 (N_20212,N_18918,N_19027);
nand U20213 (N_20213,N_18377,N_18710);
xor U20214 (N_20214,N_19108,N_18774);
and U20215 (N_20215,N_18787,N_18590);
nand U20216 (N_20216,N_18739,N_18617);
nand U20217 (N_20217,N_18295,N_18353);
or U20218 (N_20218,N_18148,N_18008);
nand U20219 (N_20219,N_18683,N_18143);
nand U20220 (N_20220,N_18722,N_18486);
or U20221 (N_20221,N_18899,N_18266);
and U20222 (N_20222,N_19175,N_18740);
or U20223 (N_20223,N_18795,N_18359);
and U20224 (N_20224,N_18938,N_18148);
xor U20225 (N_20225,N_18251,N_18835);
xnor U20226 (N_20226,N_18450,N_18052);
nor U20227 (N_20227,N_18028,N_18461);
xor U20228 (N_20228,N_18133,N_18653);
or U20229 (N_20229,N_18473,N_18900);
and U20230 (N_20230,N_18939,N_18015);
and U20231 (N_20231,N_19033,N_19077);
nand U20232 (N_20232,N_18063,N_19115);
nor U20233 (N_20233,N_18948,N_18692);
xor U20234 (N_20234,N_18524,N_18082);
nand U20235 (N_20235,N_18805,N_18004);
nand U20236 (N_20236,N_18173,N_18186);
nand U20237 (N_20237,N_18760,N_19013);
nor U20238 (N_20238,N_18269,N_18198);
xnor U20239 (N_20239,N_18750,N_18176);
xnor U20240 (N_20240,N_18532,N_18949);
nand U20241 (N_20241,N_18075,N_18174);
xor U20242 (N_20242,N_18719,N_18806);
nand U20243 (N_20243,N_18052,N_18736);
xor U20244 (N_20244,N_18892,N_18886);
nand U20245 (N_20245,N_18296,N_18129);
and U20246 (N_20246,N_18663,N_18352);
or U20247 (N_20247,N_18579,N_18164);
or U20248 (N_20248,N_18696,N_18054);
or U20249 (N_20249,N_18243,N_18577);
nor U20250 (N_20250,N_18704,N_18506);
or U20251 (N_20251,N_18081,N_18057);
nor U20252 (N_20252,N_19049,N_18181);
and U20253 (N_20253,N_19161,N_18443);
or U20254 (N_20254,N_18131,N_18190);
or U20255 (N_20255,N_18440,N_18975);
and U20256 (N_20256,N_18854,N_18427);
xor U20257 (N_20257,N_18938,N_19164);
or U20258 (N_20258,N_19141,N_18753);
and U20259 (N_20259,N_18542,N_18824);
xor U20260 (N_20260,N_18083,N_19135);
nor U20261 (N_20261,N_19072,N_18873);
or U20262 (N_20262,N_18197,N_18009);
xnor U20263 (N_20263,N_18545,N_18221);
or U20264 (N_20264,N_18382,N_18380);
or U20265 (N_20265,N_18899,N_18641);
or U20266 (N_20266,N_18567,N_18712);
nand U20267 (N_20267,N_18693,N_18304);
nand U20268 (N_20268,N_18973,N_18826);
xnor U20269 (N_20269,N_18956,N_18633);
and U20270 (N_20270,N_18698,N_18201);
nand U20271 (N_20271,N_18803,N_18936);
and U20272 (N_20272,N_19050,N_18493);
and U20273 (N_20273,N_18426,N_18803);
or U20274 (N_20274,N_18745,N_18776);
nor U20275 (N_20275,N_18450,N_18261);
and U20276 (N_20276,N_18755,N_19102);
nand U20277 (N_20277,N_19127,N_18610);
nor U20278 (N_20278,N_19120,N_18813);
nand U20279 (N_20279,N_18972,N_18212);
nor U20280 (N_20280,N_19067,N_18976);
nand U20281 (N_20281,N_18378,N_18006);
nor U20282 (N_20282,N_18672,N_18060);
and U20283 (N_20283,N_19165,N_18544);
and U20284 (N_20284,N_19097,N_18601);
nand U20285 (N_20285,N_18761,N_18173);
nor U20286 (N_20286,N_18594,N_18961);
or U20287 (N_20287,N_18814,N_19088);
and U20288 (N_20288,N_18201,N_18529);
and U20289 (N_20289,N_18775,N_18479);
nor U20290 (N_20290,N_18544,N_18382);
xnor U20291 (N_20291,N_18375,N_18249);
nor U20292 (N_20292,N_19057,N_18711);
and U20293 (N_20293,N_18784,N_18280);
nand U20294 (N_20294,N_18615,N_18568);
nor U20295 (N_20295,N_18401,N_18188);
and U20296 (N_20296,N_19015,N_18415);
xor U20297 (N_20297,N_18401,N_18166);
nor U20298 (N_20298,N_18169,N_18575);
nand U20299 (N_20299,N_18366,N_18798);
or U20300 (N_20300,N_18507,N_18540);
and U20301 (N_20301,N_19143,N_18113);
nor U20302 (N_20302,N_18933,N_18569);
nand U20303 (N_20303,N_18407,N_18322);
xnor U20304 (N_20304,N_18383,N_19119);
nand U20305 (N_20305,N_18873,N_18007);
xor U20306 (N_20306,N_18391,N_18182);
xor U20307 (N_20307,N_18730,N_18603);
nor U20308 (N_20308,N_18085,N_18058);
nor U20309 (N_20309,N_18381,N_18331);
or U20310 (N_20310,N_18819,N_18508);
nor U20311 (N_20311,N_18860,N_18355);
xnor U20312 (N_20312,N_19059,N_18779);
xnor U20313 (N_20313,N_18535,N_18554);
and U20314 (N_20314,N_18777,N_18020);
nand U20315 (N_20315,N_18400,N_18548);
or U20316 (N_20316,N_18711,N_18689);
nand U20317 (N_20317,N_19054,N_18349);
xor U20318 (N_20318,N_19054,N_18031);
xor U20319 (N_20319,N_18673,N_18552);
nor U20320 (N_20320,N_18911,N_19055);
nor U20321 (N_20321,N_18444,N_18758);
and U20322 (N_20322,N_19139,N_19013);
nor U20323 (N_20323,N_18969,N_18617);
nand U20324 (N_20324,N_19142,N_18713);
xor U20325 (N_20325,N_18401,N_18542);
nor U20326 (N_20326,N_19006,N_18910);
nand U20327 (N_20327,N_18575,N_18646);
and U20328 (N_20328,N_19163,N_19025);
and U20329 (N_20329,N_18101,N_18964);
and U20330 (N_20330,N_18400,N_18857);
nor U20331 (N_20331,N_19129,N_18925);
and U20332 (N_20332,N_18303,N_18980);
or U20333 (N_20333,N_19078,N_18011);
xor U20334 (N_20334,N_18855,N_19107);
nor U20335 (N_20335,N_18992,N_18208);
or U20336 (N_20336,N_18557,N_18996);
xor U20337 (N_20337,N_18080,N_18931);
or U20338 (N_20338,N_18896,N_18671);
and U20339 (N_20339,N_18486,N_18207);
nor U20340 (N_20340,N_19157,N_18445);
nor U20341 (N_20341,N_18437,N_18316);
nor U20342 (N_20342,N_18497,N_18007);
nand U20343 (N_20343,N_18212,N_18137);
nand U20344 (N_20344,N_19135,N_18449);
or U20345 (N_20345,N_18877,N_19113);
or U20346 (N_20346,N_18511,N_19178);
xor U20347 (N_20347,N_18325,N_18414);
and U20348 (N_20348,N_18293,N_18598);
xnor U20349 (N_20349,N_18369,N_18172);
nand U20350 (N_20350,N_18909,N_18929);
or U20351 (N_20351,N_19197,N_18189);
and U20352 (N_20352,N_18249,N_18049);
nand U20353 (N_20353,N_18455,N_19124);
nand U20354 (N_20354,N_18739,N_18664);
nand U20355 (N_20355,N_18398,N_19168);
nand U20356 (N_20356,N_18664,N_18336);
nand U20357 (N_20357,N_18911,N_18016);
or U20358 (N_20358,N_19091,N_18745);
nor U20359 (N_20359,N_19054,N_19143);
nand U20360 (N_20360,N_19005,N_18875);
or U20361 (N_20361,N_18732,N_18253);
nand U20362 (N_20362,N_18133,N_18204);
nor U20363 (N_20363,N_18072,N_19126);
nand U20364 (N_20364,N_18563,N_18781);
xor U20365 (N_20365,N_18952,N_18461);
xor U20366 (N_20366,N_19114,N_18831);
and U20367 (N_20367,N_18541,N_18740);
and U20368 (N_20368,N_18316,N_19065);
nand U20369 (N_20369,N_18484,N_19100);
nand U20370 (N_20370,N_18354,N_18607);
and U20371 (N_20371,N_18818,N_18386);
xor U20372 (N_20372,N_19164,N_19124);
xnor U20373 (N_20373,N_19097,N_18472);
and U20374 (N_20374,N_18432,N_18428);
nor U20375 (N_20375,N_18698,N_18549);
nor U20376 (N_20376,N_18041,N_18220);
nand U20377 (N_20377,N_19196,N_18202);
xor U20378 (N_20378,N_18366,N_18521);
nor U20379 (N_20379,N_18294,N_19029);
nand U20380 (N_20380,N_18091,N_18282);
xnor U20381 (N_20381,N_18169,N_18231);
nor U20382 (N_20382,N_18847,N_18324);
xnor U20383 (N_20383,N_18639,N_18109);
nand U20384 (N_20384,N_18101,N_18903);
xor U20385 (N_20385,N_18419,N_19174);
nand U20386 (N_20386,N_18367,N_18143);
nand U20387 (N_20387,N_18279,N_18248);
or U20388 (N_20388,N_18810,N_18046);
or U20389 (N_20389,N_18931,N_18660);
nand U20390 (N_20390,N_18388,N_18841);
xor U20391 (N_20391,N_18067,N_18156);
nand U20392 (N_20392,N_18445,N_18567);
nand U20393 (N_20393,N_18088,N_18674);
nand U20394 (N_20394,N_18879,N_18540);
and U20395 (N_20395,N_18804,N_18136);
xor U20396 (N_20396,N_18423,N_18808);
and U20397 (N_20397,N_18338,N_18115);
nor U20398 (N_20398,N_19199,N_19171);
xor U20399 (N_20399,N_18935,N_18987);
nand U20400 (N_20400,N_19897,N_20203);
or U20401 (N_20401,N_19265,N_20335);
and U20402 (N_20402,N_20373,N_19636);
xor U20403 (N_20403,N_19713,N_20370);
or U20404 (N_20404,N_20323,N_19230);
xnor U20405 (N_20405,N_19612,N_19760);
nand U20406 (N_20406,N_20114,N_19876);
xnor U20407 (N_20407,N_19562,N_20033);
nand U20408 (N_20408,N_20354,N_19238);
nor U20409 (N_20409,N_19768,N_19848);
nor U20410 (N_20410,N_19305,N_19381);
nand U20411 (N_20411,N_19700,N_19289);
xnor U20412 (N_20412,N_19383,N_19797);
nand U20413 (N_20413,N_19386,N_19791);
or U20414 (N_20414,N_20379,N_20130);
nor U20415 (N_20415,N_20342,N_19615);
nand U20416 (N_20416,N_19972,N_19762);
and U20417 (N_20417,N_19516,N_19501);
or U20418 (N_20418,N_19417,N_20350);
xnor U20419 (N_20419,N_19464,N_19853);
or U20420 (N_20420,N_20080,N_19888);
nand U20421 (N_20421,N_19886,N_20262);
and U20422 (N_20422,N_19767,N_20004);
xnor U20423 (N_20423,N_19217,N_19505);
nor U20424 (N_20424,N_20123,N_19325);
nand U20425 (N_20425,N_19926,N_19517);
xor U20426 (N_20426,N_19406,N_20113);
nor U20427 (N_20427,N_19653,N_20239);
xor U20428 (N_20428,N_19327,N_20027);
nand U20429 (N_20429,N_19293,N_19777);
and U20430 (N_20430,N_19795,N_19958);
nand U20431 (N_20431,N_19640,N_20233);
nand U20432 (N_20432,N_19874,N_19409);
or U20433 (N_20433,N_20244,N_19870);
nor U20434 (N_20434,N_19969,N_19712);
nor U20435 (N_20435,N_19538,N_19428);
or U20436 (N_20436,N_20234,N_19576);
or U20437 (N_20437,N_20115,N_20394);
or U20438 (N_20438,N_19260,N_19203);
and U20439 (N_20439,N_19366,N_19866);
nor U20440 (N_20440,N_20199,N_19492);
nand U20441 (N_20441,N_19588,N_19745);
nor U20442 (N_20442,N_19607,N_19865);
and U20443 (N_20443,N_19323,N_19833);
nor U20444 (N_20444,N_19765,N_19707);
and U20445 (N_20445,N_20003,N_19533);
nand U20446 (N_20446,N_20051,N_20336);
and U20447 (N_20447,N_20015,N_20277);
nand U20448 (N_20448,N_19288,N_19262);
nor U20449 (N_20449,N_19592,N_20014);
xnor U20450 (N_20450,N_19316,N_20363);
or U20451 (N_20451,N_20361,N_19726);
xor U20452 (N_20452,N_19559,N_19749);
and U20453 (N_20453,N_20393,N_19264);
xnor U20454 (N_20454,N_19678,N_20388);
or U20455 (N_20455,N_19626,N_19877);
nand U20456 (N_20456,N_19318,N_19365);
xor U20457 (N_20457,N_20073,N_19580);
xnor U20458 (N_20458,N_19332,N_19402);
nand U20459 (N_20459,N_19385,N_19404);
nand U20460 (N_20460,N_19393,N_19359);
or U20461 (N_20461,N_20134,N_20349);
or U20462 (N_20462,N_19670,N_20387);
or U20463 (N_20463,N_20315,N_20137);
nor U20464 (N_20464,N_20043,N_19963);
or U20465 (N_20465,N_20328,N_19210);
xor U20466 (N_20466,N_19589,N_20374);
and U20467 (N_20467,N_19493,N_20170);
nand U20468 (N_20468,N_19574,N_19910);
or U20469 (N_20469,N_19380,N_20305);
and U20470 (N_20470,N_19556,N_19583);
or U20471 (N_20471,N_19675,N_20299);
or U20472 (N_20472,N_19875,N_19689);
or U20473 (N_20473,N_19304,N_19807);
nand U20474 (N_20474,N_19457,N_19526);
and U20475 (N_20475,N_19803,N_19237);
xor U20476 (N_20476,N_19548,N_19256);
nor U20477 (N_20477,N_19328,N_19962);
xnor U20478 (N_20478,N_19826,N_19337);
nand U20479 (N_20479,N_19776,N_19672);
nand U20480 (N_20480,N_19280,N_20297);
nand U20481 (N_20481,N_20242,N_19602);
nand U20482 (N_20482,N_20337,N_19658);
xor U20483 (N_20483,N_19463,N_19285);
nor U20484 (N_20484,N_19269,N_20247);
xor U20485 (N_20485,N_19449,N_19849);
or U20486 (N_20486,N_19993,N_19697);
or U20487 (N_20487,N_19277,N_20389);
or U20488 (N_20488,N_19647,N_19551);
xor U20489 (N_20489,N_19416,N_20365);
and U20490 (N_20490,N_19223,N_20183);
nand U20491 (N_20491,N_19593,N_19465);
nor U20492 (N_20492,N_19818,N_19834);
and U20493 (N_20493,N_19934,N_19349);
and U20494 (N_20494,N_19775,N_19307);
nor U20495 (N_20495,N_19825,N_19632);
or U20496 (N_20496,N_20212,N_19793);
nand U20497 (N_20497,N_19320,N_19233);
xnor U20498 (N_20498,N_20097,N_20283);
and U20499 (N_20499,N_20284,N_20383);
nor U20500 (N_20500,N_19927,N_20108);
nand U20501 (N_20501,N_19893,N_19213);
and U20502 (N_20502,N_19604,N_20111);
xor U20503 (N_20503,N_19701,N_19204);
and U20504 (N_20504,N_19451,N_19840);
nand U20505 (N_20505,N_19659,N_19908);
nand U20506 (N_20506,N_20346,N_19510);
nor U20507 (N_20507,N_20044,N_19944);
nor U20508 (N_20508,N_19430,N_20359);
or U20509 (N_20509,N_19437,N_19747);
and U20510 (N_20510,N_19873,N_19567);
nor U20511 (N_20511,N_20240,N_19633);
or U20512 (N_20512,N_19374,N_19480);
and U20513 (N_20513,N_20188,N_20232);
nand U20514 (N_20514,N_19912,N_19804);
and U20515 (N_20515,N_19751,N_20301);
or U20516 (N_20516,N_19508,N_19554);
nand U20517 (N_20517,N_19940,N_20302);
or U20518 (N_20518,N_19988,N_20165);
nand U20519 (N_20519,N_19757,N_19945);
xor U20520 (N_20520,N_20160,N_20088);
and U20521 (N_20521,N_19829,N_19992);
xnor U20522 (N_20522,N_20078,N_19263);
nor U20523 (N_20523,N_19234,N_20371);
xor U20524 (N_20524,N_20006,N_19918);
nand U20525 (N_20525,N_20202,N_20071);
xnor U20526 (N_20526,N_19235,N_20169);
and U20527 (N_20527,N_19929,N_20321);
and U20528 (N_20528,N_19355,N_19858);
nor U20529 (N_20529,N_19856,N_19577);
and U20530 (N_20530,N_19925,N_20171);
nor U20531 (N_20531,N_19652,N_19980);
nor U20532 (N_20532,N_20200,N_20372);
xnor U20533 (N_20533,N_19321,N_19471);
and U20534 (N_20534,N_20107,N_19419);
or U20535 (N_20535,N_20102,N_19843);
or U20536 (N_20536,N_19522,N_19738);
or U20537 (N_20537,N_19821,N_20220);
or U20538 (N_20538,N_19692,N_19601);
xnor U20539 (N_20539,N_20013,N_19789);
nor U20540 (N_20540,N_19693,N_20204);
nand U20541 (N_20541,N_20266,N_19206);
nand U20542 (N_20542,N_19823,N_19442);
or U20543 (N_20543,N_19744,N_20235);
nand U20544 (N_20544,N_20101,N_19345);
nand U20545 (N_20545,N_19618,N_20042);
xor U20546 (N_20546,N_20077,N_20012);
xnor U20547 (N_20547,N_20360,N_20248);
xor U20548 (N_20548,N_19362,N_19390);
xor U20549 (N_20549,N_20369,N_20243);
and U20550 (N_20550,N_19252,N_19654);
or U20551 (N_20551,N_19590,N_20106);
or U20552 (N_20552,N_19450,N_20192);
and U20553 (N_20553,N_19754,N_20019);
nor U20554 (N_20554,N_19524,N_19688);
nor U20555 (N_20555,N_19731,N_19903);
xor U20556 (N_20556,N_19594,N_19569);
or U20557 (N_20557,N_19790,N_19857);
or U20558 (N_20558,N_19528,N_19224);
or U20559 (N_20559,N_19244,N_20245);
and U20560 (N_20560,N_19837,N_20206);
nand U20561 (N_20561,N_19617,N_19846);
nor U20562 (N_20562,N_19911,N_20303);
xnor U20563 (N_20563,N_19625,N_19724);
and U20564 (N_20564,N_19591,N_20050);
nor U20565 (N_20565,N_20332,N_19811);
nand U20566 (N_20566,N_19281,N_19624);
or U20567 (N_20567,N_20310,N_19202);
or U20568 (N_20568,N_20161,N_20195);
or U20569 (N_20569,N_19801,N_19350);
and U20570 (N_20570,N_20076,N_19919);
or U20571 (N_20571,N_19597,N_20309);
and U20572 (N_20572,N_20023,N_19728);
nor U20573 (N_20573,N_20162,N_20344);
nor U20574 (N_20574,N_19951,N_19581);
and U20575 (N_20575,N_19663,N_19308);
xor U20576 (N_20576,N_19921,N_19805);
nand U20577 (N_20577,N_19816,N_19555);
and U20578 (N_20578,N_20037,N_19536);
or U20579 (N_20579,N_20246,N_20380);
nor U20580 (N_20580,N_20020,N_19466);
nand U20581 (N_20581,N_20083,N_19907);
nand U20582 (N_20582,N_20109,N_19324);
nor U20583 (N_20583,N_19884,N_19302);
or U20584 (N_20584,N_20213,N_19674);
nand U20585 (N_20585,N_19820,N_19950);
nor U20586 (N_20586,N_19844,N_19788);
and U20587 (N_20587,N_20357,N_19309);
nand U20588 (N_20588,N_20312,N_20053);
xnor U20589 (N_20589,N_19706,N_20105);
or U20590 (N_20590,N_19571,N_20172);
nor U20591 (N_20591,N_19671,N_19900);
xnor U20592 (N_20592,N_19369,N_20047);
and U20593 (N_20593,N_19985,N_20175);
or U20594 (N_20594,N_20093,N_20264);
nor U20595 (N_20595,N_19455,N_20021);
nand U20596 (N_20596,N_19232,N_20186);
and U20597 (N_20597,N_19438,N_19412);
nor U20598 (N_20598,N_20227,N_19483);
nand U20599 (N_20599,N_20024,N_20280);
xnor U20600 (N_20600,N_19936,N_20112);
or U20601 (N_20601,N_19655,N_19974);
or U20602 (N_20602,N_19892,N_20367);
nand U20603 (N_20603,N_19429,N_19787);
or U20604 (N_20604,N_19394,N_19322);
nand U20605 (N_20605,N_20348,N_20296);
xnor U20606 (N_20606,N_19913,N_20355);
and U20607 (N_20607,N_19400,N_19753);
xor U20608 (N_20608,N_19312,N_20000);
nand U20609 (N_20609,N_19682,N_20125);
nor U20610 (N_20610,N_20045,N_20174);
or U20611 (N_20611,N_19373,N_19372);
nand U20612 (N_20612,N_19499,N_19651);
nor U20613 (N_20613,N_20258,N_20218);
nand U20614 (N_20614,N_19553,N_20215);
xor U20615 (N_20615,N_20168,N_19251);
nor U20616 (N_20616,N_19491,N_19519);
and U20617 (N_20617,N_19573,N_20399);
or U20618 (N_20618,N_19964,N_19299);
nor U20619 (N_20619,N_19422,N_20103);
nand U20620 (N_20620,N_19578,N_19294);
xnor U20621 (N_20621,N_20256,N_19965);
nand U20622 (N_20622,N_19758,N_19781);
xnor U20623 (N_20623,N_19405,N_20250);
or U20624 (N_20624,N_19894,N_19595);
nand U20625 (N_20625,N_19836,N_19421);
or U20626 (N_20626,N_19520,N_19859);
and U20627 (N_20627,N_19411,N_20099);
xnor U20628 (N_20628,N_20353,N_20163);
nand U20629 (N_20629,N_20398,N_19266);
xnor U20630 (N_20630,N_20153,N_19333);
nor U20631 (N_20631,N_19699,N_20236);
or U20632 (N_20632,N_19246,N_20298);
xor U20633 (N_20633,N_19761,N_19496);
and U20634 (N_20634,N_19879,N_19639);
nor U20635 (N_20635,N_19782,N_20056);
or U20636 (N_20636,N_20282,N_19249);
or U20637 (N_20637,N_20146,N_20176);
nor U20638 (N_20638,N_19346,N_19764);
nor U20639 (N_20639,N_19730,N_19397);
xnor U20640 (N_20640,N_20230,N_19971);
xor U20641 (N_20641,N_19257,N_20141);
and U20642 (N_20642,N_19741,N_20136);
nand U20643 (N_20643,N_19975,N_19637);
xor U20644 (N_20644,N_20126,N_19432);
or U20645 (N_20645,N_19564,N_20090);
nor U20646 (N_20646,N_19622,N_19623);
nor U20647 (N_20647,N_19255,N_20209);
or U20648 (N_20648,N_19772,N_19947);
and U20649 (N_20649,N_19240,N_19502);
nor U20650 (N_20650,N_19661,N_19225);
or U20651 (N_20651,N_20274,N_20098);
nor U20652 (N_20652,N_20259,N_19287);
nor U20653 (N_20653,N_19960,N_19243);
and U20654 (N_20654,N_19851,N_19838);
xnor U20655 (N_20655,N_19719,N_20253);
xnor U20656 (N_20656,N_19798,N_20314);
and U20657 (N_20657,N_19420,N_19935);
nor U20658 (N_20658,N_20167,N_19469);
or U20659 (N_20659,N_20094,N_19282);
nor U20660 (N_20660,N_19315,N_19665);
nand U20661 (N_20661,N_20049,N_20265);
nor U20662 (N_20662,N_19854,N_20217);
nand U20663 (N_20663,N_20022,N_20198);
xnor U20664 (N_20664,N_19645,N_20179);
nor U20665 (N_20665,N_19286,N_19331);
xnor U20666 (N_20666,N_19391,N_19382);
or U20667 (N_20667,N_20397,N_19931);
and U20668 (N_20668,N_20341,N_19619);
nor U20669 (N_20669,N_19314,N_20347);
nor U20670 (N_20670,N_20178,N_19495);
or U20671 (N_20671,N_20325,N_19218);
and U20672 (N_20672,N_20276,N_19515);
nor U20673 (N_20673,N_19710,N_19222);
nor U20674 (N_20674,N_20320,N_19679);
nor U20675 (N_20675,N_20138,N_20194);
xor U20676 (N_20676,N_19871,N_19709);
xnor U20677 (N_20677,N_19447,N_19418);
xnor U20678 (N_20678,N_19933,N_19867);
nand U20679 (N_20679,N_19431,N_19458);
and U20680 (N_20680,N_19895,N_19997);
nand U20681 (N_20681,N_20364,N_19860);
nand U20682 (N_20682,N_19354,N_19605);
nand U20683 (N_20683,N_19375,N_19814);
and U20684 (N_20684,N_19497,N_19644);
nand U20685 (N_20685,N_20228,N_20281);
or U20686 (N_20686,N_19778,N_19667);
or U20687 (N_20687,N_20173,N_19334);
and U20688 (N_20688,N_19298,N_19486);
and U20689 (N_20689,N_19676,N_20016);
or U20690 (N_20690,N_19714,N_19850);
nand U20691 (N_20691,N_19736,N_19403);
or U20692 (N_20692,N_20100,N_19891);
xnor U20693 (N_20693,N_19371,N_20152);
nand U20694 (N_20694,N_19530,N_19459);
nand U20695 (N_20695,N_20092,N_20311);
nor U20696 (N_20696,N_19698,N_19991);
or U20697 (N_20697,N_19660,N_19467);
nor U20698 (N_20698,N_20142,N_20133);
or U20699 (N_20699,N_19513,N_20313);
and U20700 (N_20700,N_19769,N_20229);
and U20701 (N_20701,N_20289,N_19609);
or U20702 (N_20702,N_20261,N_20070);
nor U20703 (N_20703,N_19544,N_19389);
xnor U20704 (N_20704,N_19869,N_19852);
and U20705 (N_20705,N_20300,N_20316);
nand U20706 (N_20706,N_19957,N_19441);
nand U20707 (N_20707,N_19473,N_19606);
and U20708 (N_20708,N_19300,N_20224);
xor U20709 (N_20709,N_19247,N_20005);
nor U20710 (N_20710,N_19995,N_19446);
xor U20711 (N_20711,N_20317,N_19407);
or U20712 (N_20712,N_19915,N_19468);
xnor U20713 (N_20713,N_19529,N_19342);
nor U20714 (N_20714,N_19922,N_20011);
or U20715 (N_20715,N_19424,N_19311);
xor U20716 (N_20716,N_19329,N_20269);
xor U20717 (N_20717,N_19872,N_19426);
or U20718 (N_20718,N_19771,N_19461);
nor U20719 (N_20719,N_19792,N_19684);
and U20720 (N_20720,N_20061,N_19408);
and U20721 (N_20721,N_20164,N_20046);
or U20722 (N_20722,N_20018,N_20395);
and U20723 (N_20723,N_19648,N_20009);
xor U20724 (N_20724,N_19662,N_19396);
and U20725 (N_20725,N_19864,N_19268);
or U20726 (N_20726,N_19630,N_20382);
and U20727 (N_20727,N_19242,N_19585);
nand U20728 (N_20728,N_19568,N_20340);
xnor U20729 (N_20729,N_19948,N_19509);
or U20730 (N_20730,N_19348,N_20075);
or U20731 (N_20731,N_19208,N_20377);
nor U20732 (N_20732,N_19220,N_19587);
and U20733 (N_20733,N_19550,N_19696);
nor U20734 (N_20734,N_20193,N_19503);
nand U20735 (N_20735,N_19253,N_19832);
or U20736 (N_20736,N_19462,N_20308);
or U20737 (N_20737,N_19506,N_20197);
nor U20738 (N_20738,N_19427,N_19472);
xor U20739 (N_20739,N_19664,N_19310);
xor U20740 (N_20740,N_19376,N_20041);
xor U20741 (N_20741,N_19808,N_19668);
xnor U20742 (N_20742,N_19279,N_19540);
xor U20743 (N_20743,N_19566,N_20329);
nand U20744 (N_20744,N_19284,N_20362);
and U20745 (N_20745,N_20008,N_19953);
xor U20746 (N_20746,N_19259,N_19477);
nand U20747 (N_20747,N_19815,N_19341);
and U20748 (N_20748,N_19827,N_20072);
or U20749 (N_20749,N_20145,N_19534);
nor U20750 (N_20750,N_19868,N_19835);
nor U20751 (N_20751,N_20275,N_19977);
nand U20752 (N_20752,N_19638,N_19543);
and U20753 (N_20753,N_19786,N_19436);
xor U20754 (N_20754,N_19614,N_19558);
nand U20755 (N_20755,N_20208,N_19889);
xor U20756 (N_20756,N_20286,N_19546);
or U20757 (N_20757,N_20029,N_20118);
or U20758 (N_20758,N_19987,N_19968);
and U20759 (N_20759,N_20214,N_20159);
nand U20760 (N_20760,N_20324,N_20120);
or U20761 (N_20761,N_20196,N_19862);
and U20762 (N_20762,N_20376,N_19941);
or U20763 (N_20763,N_20226,N_19642);
and U20764 (N_20764,N_19780,N_19494);
and U20765 (N_20765,N_19914,N_19549);
and U20766 (N_20766,N_19330,N_20122);
and U20767 (N_20767,N_19563,N_19979);
nand U20768 (N_20768,N_20063,N_19500);
nand U20769 (N_20769,N_19338,N_19433);
nand U20770 (N_20770,N_19319,N_19966);
and U20771 (N_20771,N_20288,N_19207);
or U20772 (N_20772,N_19596,N_19474);
nand U20773 (N_20773,N_19512,N_20358);
xnor U20774 (N_20774,N_19335,N_19401);
and U20775 (N_20775,N_20292,N_19657);
nand U20776 (N_20776,N_19610,N_19641);
nand U20777 (N_20777,N_19507,N_20263);
xor U20778 (N_20778,N_19742,N_20327);
or U20779 (N_20779,N_19887,N_19275);
nand U20780 (N_20780,N_19479,N_19802);
xor U20781 (N_20781,N_20338,N_19978);
nor U20782 (N_20782,N_19750,N_19398);
and U20783 (N_20783,N_19221,N_19236);
nand U20784 (N_20784,N_19690,N_19627);
xor U20785 (N_20785,N_20254,N_19514);
nand U20786 (N_20786,N_19650,N_20082);
nand U20787 (N_20787,N_19521,N_20057);
xnor U20788 (N_20788,N_19229,N_19785);
and U20789 (N_20789,N_20375,N_19537);
and U20790 (N_20790,N_19228,N_20052);
xor U20791 (N_20791,N_19248,N_20287);
nor U20792 (N_20792,N_19219,N_20095);
xor U20793 (N_20793,N_19928,N_19478);
and U20794 (N_20794,N_19796,N_19600);
xnor U20795 (N_20795,N_20293,N_20396);
nand U20796 (N_20796,N_20030,N_19608);
xor U20797 (N_20797,N_20270,N_19685);
or U20798 (N_20798,N_19364,N_19841);
or U20799 (N_20799,N_19909,N_19952);
nor U20800 (N_20800,N_20066,N_19292);
nand U20801 (N_20801,N_20185,N_20386);
and U20802 (N_20802,N_19949,N_19484);
nand U20803 (N_20803,N_19806,N_19504);
or U20804 (N_20804,N_19643,N_19254);
or U20805 (N_20805,N_20251,N_19634);
xor U20806 (N_20806,N_20059,N_19711);
nand U20807 (N_20807,N_19705,N_19340);
nor U20808 (N_20808,N_19923,N_19475);
nand U20809 (N_20809,N_19445,N_19582);
xnor U20810 (N_20810,N_19983,N_20110);
nand U20811 (N_20811,N_19687,N_19347);
and U20812 (N_20812,N_19939,N_19721);
xor U20813 (N_20813,N_19488,N_19613);
nor U20814 (N_20814,N_20064,N_20366);
nand U20815 (N_20815,N_20104,N_19902);
and U20816 (N_20816,N_19215,N_20117);
nor U20817 (N_20817,N_20166,N_20290);
nand U20818 (N_20818,N_20237,N_19456);
and U20819 (N_20819,N_19822,N_19905);
and U20820 (N_20820,N_19920,N_19273);
and U20821 (N_20821,N_20306,N_19924);
nand U20822 (N_20822,N_20087,N_19881);
xnor U20823 (N_20823,N_19239,N_19628);
and U20824 (N_20824,N_20119,N_20028);
nand U20825 (N_20825,N_20238,N_20149);
xnor U20826 (N_20826,N_19527,N_20055);
nand U20827 (N_20827,N_19946,N_19882);
xnor U20828 (N_20828,N_19973,N_19970);
nor U20829 (N_20829,N_20268,N_19646);
or U20830 (N_20830,N_19677,N_19276);
xnor U20831 (N_20831,N_19784,N_19227);
nor U20832 (N_20832,N_19363,N_20158);
nand U20833 (N_20833,N_20255,N_19998);
or U20834 (N_20834,N_20326,N_19565);
nor U20835 (N_20835,N_19766,N_19379);
nor U20836 (N_20836,N_20144,N_19722);
nand U20837 (N_20837,N_20121,N_19317);
nand U20838 (N_20838,N_19387,N_20307);
xor U20839 (N_20839,N_19370,N_19367);
nor U20840 (N_20840,N_19388,N_19733);
nand U20841 (N_20841,N_20150,N_19414);
nand U20842 (N_20842,N_20091,N_19831);
or U20843 (N_20843,N_19226,N_20054);
xnor U20844 (N_20844,N_20128,N_19976);
nand U20845 (N_20845,N_19425,N_20007);
nor U20846 (N_20846,N_19301,N_20089);
nand U20847 (N_20847,N_19523,N_19603);
nand U20848 (N_20848,N_20257,N_19720);
xor U20849 (N_20849,N_19616,N_20086);
xnor U20850 (N_20850,N_20390,N_19673);
nor U20851 (N_20851,N_19539,N_19454);
xor U20852 (N_20852,N_20143,N_20260);
and U20853 (N_20853,N_19800,N_19635);
nand U20854 (N_20854,N_20180,N_19755);
or U20855 (N_20855,N_19353,N_19413);
nor U20856 (N_20856,N_19377,N_20002);
and U20857 (N_20857,N_19930,N_19989);
nor U20858 (N_20858,N_20392,N_20356);
or U20859 (N_20859,N_19448,N_19216);
xor U20860 (N_20860,N_19250,N_19271);
or U20861 (N_20861,N_19984,N_20210);
xor U20862 (N_20862,N_19901,N_19541);
xor U20863 (N_20863,N_19579,N_19368);
xnor U20864 (N_20864,N_19681,N_20249);
nor U20865 (N_20865,N_19904,N_20148);
and U20866 (N_20866,N_20241,N_20060);
nor U20867 (N_20867,N_19440,N_19231);
nor U20868 (N_20868,N_20222,N_19740);
and U20869 (N_20869,N_19295,N_19545);
xor U20870 (N_20870,N_20334,N_20271);
and U20871 (N_20871,N_20036,N_20096);
xnor U20872 (N_20872,N_19961,N_20156);
nand U20873 (N_20873,N_19525,N_20010);
or U20874 (N_20874,N_19666,N_19278);
nand U20875 (N_20875,N_19272,N_19205);
or U20876 (N_20876,N_19611,N_19476);
nor U20877 (N_20877,N_19990,N_20040);
nor U20878 (N_20878,N_20368,N_20333);
nor U20879 (N_20879,N_19982,N_20322);
nand U20880 (N_20880,N_19727,N_19942);
and U20881 (N_20881,N_20139,N_19290);
and U20882 (N_20882,N_19861,N_19956);
and U20883 (N_20883,N_20351,N_19932);
nand U20884 (N_20884,N_19774,N_19737);
nor U20885 (N_20885,N_19906,N_20181);
nor U20886 (N_20886,N_19986,N_20079);
xnor U20887 (N_20887,N_19686,N_20343);
or U20888 (N_20888,N_20062,N_19855);
and U20889 (N_20889,N_19880,N_19715);
xnor U20890 (N_20890,N_19303,N_19959);
nand U20891 (N_20891,N_19415,N_19680);
and U20892 (N_20892,N_19584,N_19702);
and U20893 (N_20893,N_19211,N_19570);
or U20894 (N_20894,N_20385,N_19485);
xor U20895 (N_20895,N_19890,N_20039);
and U20896 (N_20896,N_20304,N_20184);
nor U20897 (N_20897,N_20318,N_20155);
and U20898 (N_20898,N_20378,N_19621);
nand U20899 (N_20899,N_19824,N_19481);
nor U20900 (N_20900,N_20127,N_19352);
or U20901 (N_20901,N_20031,N_19356);
or U20902 (N_20902,N_19898,N_19732);
or U20903 (N_20903,N_20273,N_19885);
or U20904 (N_20904,N_20331,N_20081);
nor U20905 (N_20905,N_19981,N_19734);
nor U20906 (N_20906,N_19384,N_20345);
and U20907 (N_20907,N_20285,N_20391);
nor U20908 (N_20908,N_19490,N_19511);
nand U20909 (N_20909,N_20157,N_19336);
and U20910 (N_20910,N_19470,N_19810);
nand U20911 (N_20911,N_19756,N_19830);
and U20912 (N_20912,N_20201,N_20182);
xnor U20913 (N_20913,N_20116,N_19967);
and U20914 (N_20914,N_20223,N_20017);
nor U20915 (N_20915,N_20048,N_19779);
or U20916 (N_20916,N_19717,N_19725);
xnor U20917 (N_20917,N_19708,N_19245);
or U20918 (N_20918,N_19656,N_20025);
and U20919 (N_20919,N_19683,N_19410);
and U20920 (N_20920,N_19954,N_20026);
nor U20921 (N_20921,N_19955,N_19817);
nand U20922 (N_20922,N_19839,N_20069);
or U20923 (N_20923,N_19718,N_19439);
nand U20924 (N_20924,N_19241,N_19599);
or U20925 (N_20925,N_20189,N_20084);
or U20926 (N_20926,N_19794,N_19274);
or U20927 (N_20927,N_19297,N_19392);
and U20928 (N_20928,N_19812,N_19452);
xor U20929 (N_20929,N_19560,N_19916);
nand U20930 (N_20930,N_20177,N_19994);
and U20931 (N_20931,N_19899,N_19552);
nor U20932 (N_20932,N_20035,N_20219);
or U20933 (N_20933,N_20278,N_19723);
xnor U20934 (N_20934,N_20221,N_20065);
or U20935 (N_20935,N_19489,N_19214);
nor U20936 (N_20936,N_20132,N_19399);
and U20937 (N_20937,N_20001,N_19518);
xnor U20938 (N_20938,N_19999,N_19575);
or U20939 (N_20939,N_20154,N_20140);
and U20940 (N_20940,N_19783,N_19532);
and U20941 (N_20941,N_19201,N_19453);
nand U20942 (N_20942,N_19443,N_20034);
nor U20943 (N_20943,N_19631,N_19743);
and U20944 (N_20944,N_20381,N_20330);
xnor U20945 (N_20945,N_20147,N_20085);
xor U20946 (N_20946,N_19360,N_19395);
nand U20947 (N_20947,N_19498,N_19669);
or U20948 (N_20948,N_19842,N_19813);
xnor U20949 (N_20949,N_19444,N_19809);
nor U20950 (N_20950,N_20294,N_20231);
or U20951 (N_20951,N_19694,N_20058);
nand U20952 (N_20952,N_19620,N_19547);
nor U20953 (N_20953,N_20216,N_19598);
nor U20954 (N_20954,N_20279,N_20151);
or U20955 (N_20955,N_19763,N_19883);
xor U20956 (N_20956,N_19212,N_20295);
nand U20957 (N_20957,N_19258,N_20207);
or U20958 (N_20958,N_19487,N_19748);
nand U20959 (N_20959,N_20267,N_19344);
nand U20960 (N_20960,N_19535,N_20190);
xnor U20961 (N_20961,N_19695,N_19326);
or U20962 (N_20962,N_19313,N_20191);
nand U20963 (N_20963,N_19209,N_20067);
nand U20964 (N_20964,N_19586,N_20225);
xor U20965 (N_20965,N_20211,N_20187);
or U20966 (N_20966,N_19557,N_19729);
xor U20967 (N_20967,N_19270,N_19343);
nor U20968 (N_20968,N_20131,N_19896);
and U20969 (N_20969,N_19200,N_19291);
nor U20970 (N_20970,N_19351,N_19339);
and U20971 (N_20971,N_19283,N_19572);
and U20972 (N_20972,N_20384,N_19704);
xor U20973 (N_20973,N_19703,N_19799);
or U20974 (N_20974,N_19746,N_19938);
nand U20975 (N_20975,N_20129,N_19460);
nand U20976 (N_20976,N_20124,N_19629);
xnor U20977 (N_20977,N_19819,N_19716);
and U20978 (N_20978,N_19752,N_20352);
and U20979 (N_20979,N_19996,N_19773);
and U20980 (N_20980,N_19845,N_19561);
nor U20981 (N_20981,N_19878,N_19847);
xnor U20982 (N_20982,N_19691,N_20032);
nand U20983 (N_20983,N_19863,N_19943);
or U20984 (N_20984,N_20272,N_19361);
nor U20985 (N_20985,N_19482,N_19296);
nand U20986 (N_20986,N_20252,N_19357);
xnor U20987 (N_20987,N_19531,N_19759);
or U20988 (N_20988,N_19735,N_20074);
nor U20989 (N_20989,N_19423,N_19306);
or U20990 (N_20990,N_19267,N_19828);
nand U20991 (N_20991,N_19770,N_19917);
xnor U20992 (N_20992,N_20205,N_20339);
or U20993 (N_20993,N_19434,N_19358);
or U20994 (N_20994,N_20319,N_20068);
or U20995 (N_20995,N_19435,N_20135);
or U20996 (N_20996,N_19378,N_19649);
nor U20997 (N_20997,N_19261,N_19739);
or U20998 (N_20998,N_19937,N_19542);
and U20999 (N_20999,N_20038,N_20291);
and U21000 (N_21000,N_19838,N_20015);
nor U21001 (N_21001,N_19558,N_19370);
or U21002 (N_21002,N_20038,N_19477);
nor U21003 (N_21003,N_19271,N_19918);
xor U21004 (N_21004,N_20004,N_20217);
xnor U21005 (N_21005,N_20270,N_19554);
and U21006 (N_21006,N_20386,N_19722);
nand U21007 (N_21007,N_19872,N_19638);
xor U21008 (N_21008,N_19612,N_19971);
or U21009 (N_21009,N_19217,N_19468);
xor U21010 (N_21010,N_19454,N_19600);
and U21011 (N_21011,N_19945,N_19631);
or U21012 (N_21012,N_19517,N_19411);
nor U21013 (N_21013,N_19928,N_20306);
xor U21014 (N_21014,N_19816,N_19354);
or U21015 (N_21015,N_20024,N_19543);
nand U21016 (N_21016,N_19203,N_19930);
nor U21017 (N_21017,N_19578,N_19540);
nand U21018 (N_21018,N_20312,N_20158);
nor U21019 (N_21019,N_19565,N_20131);
xnor U21020 (N_21020,N_19881,N_19403);
xor U21021 (N_21021,N_19862,N_19716);
and U21022 (N_21022,N_19966,N_20129);
and U21023 (N_21023,N_19405,N_20398);
or U21024 (N_21024,N_19759,N_19981);
nor U21025 (N_21025,N_20247,N_19454);
and U21026 (N_21026,N_19910,N_19440);
nand U21027 (N_21027,N_19465,N_19800);
or U21028 (N_21028,N_19970,N_19698);
nand U21029 (N_21029,N_19902,N_19608);
or U21030 (N_21030,N_19841,N_19257);
or U21031 (N_21031,N_19331,N_19950);
xor U21032 (N_21032,N_19732,N_20386);
or U21033 (N_21033,N_20371,N_19469);
or U21034 (N_21034,N_19731,N_19773);
and U21035 (N_21035,N_20000,N_19788);
xor U21036 (N_21036,N_19229,N_19880);
nand U21037 (N_21037,N_20099,N_19897);
nand U21038 (N_21038,N_19243,N_19554);
xor U21039 (N_21039,N_19226,N_20032);
and U21040 (N_21040,N_19898,N_20027);
xor U21041 (N_21041,N_19463,N_19577);
or U21042 (N_21042,N_19622,N_19816);
nor U21043 (N_21043,N_19520,N_19554);
xnor U21044 (N_21044,N_19679,N_20331);
xor U21045 (N_21045,N_20118,N_19742);
nor U21046 (N_21046,N_19535,N_19512);
and U21047 (N_21047,N_20165,N_19913);
nor U21048 (N_21048,N_19543,N_20028);
nand U21049 (N_21049,N_19791,N_19303);
and U21050 (N_21050,N_19297,N_20061);
nor U21051 (N_21051,N_19441,N_20210);
nand U21052 (N_21052,N_20284,N_19649);
and U21053 (N_21053,N_20355,N_19881);
or U21054 (N_21054,N_19329,N_19619);
xnor U21055 (N_21055,N_20289,N_19438);
or U21056 (N_21056,N_19997,N_19618);
nor U21057 (N_21057,N_19962,N_19790);
nor U21058 (N_21058,N_19747,N_19518);
nor U21059 (N_21059,N_19375,N_19329);
or U21060 (N_21060,N_19217,N_19396);
xnor U21061 (N_21061,N_19485,N_19810);
nor U21062 (N_21062,N_20029,N_20051);
and U21063 (N_21063,N_19823,N_19308);
nor U21064 (N_21064,N_19200,N_19202);
nand U21065 (N_21065,N_19460,N_20118);
or U21066 (N_21066,N_19495,N_19454);
nand U21067 (N_21067,N_19905,N_19424);
xnor U21068 (N_21068,N_20250,N_19893);
nor U21069 (N_21069,N_19802,N_19938);
and U21070 (N_21070,N_19755,N_19842);
nor U21071 (N_21071,N_19868,N_20164);
xor U21072 (N_21072,N_20146,N_19222);
nor U21073 (N_21073,N_19258,N_19447);
nand U21074 (N_21074,N_20014,N_19865);
nor U21075 (N_21075,N_19443,N_20155);
nand U21076 (N_21076,N_19648,N_19779);
nor U21077 (N_21077,N_19647,N_19402);
xnor U21078 (N_21078,N_20122,N_19967);
and U21079 (N_21079,N_19693,N_19524);
nor U21080 (N_21080,N_19730,N_20215);
or U21081 (N_21081,N_19503,N_19636);
nand U21082 (N_21082,N_20283,N_19622);
and U21083 (N_21083,N_20323,N_20297);
or U21084 (N_21084,N_20047,N_19315);
xor U21085 (N_21085,N_19413,N_20394);
or U21086 (N_21086,N_19257,N_19431);
or U21087 (N_21087,N_19544,N_19788);
nand U21088 (N_21088,N_20089,N_19892);
nand U21089 (N_21089,N_19312,N_19458);
and U21090 (N_21090,N_19276,N_20092);
xnor U21091 (N_21091,N_20034,N_20217);
nand U21092 (N_21092,N_19570,N_19339);
nand U21093 (N_21093,N_19772,N_19881);
nor U21094 (N_21094,N_19493,N_19583);
nor U21095 (N_21095,N_19228,N_19473);
and U21096 (N_21096,N_20166,N_19657);
xor U21097 (N_21097,N_19963,N_19414);
xor U21098 (N_21098,N_20158,N_19216);
and U21099 (N_21099,N_20018,N_20269);
and U21100 (N_21100,N_20195,N_19712);
nor U21101 (N_21101,N_20220,N_20236);
nor U21102 (N_21102,N_19306,N_19740);
nand U21103 (N_21103,N_20108,N_19449);
or U21104 (N_21104,N_20196,N_20004);
and U21105 (N_21105,N_19676,N_20050);
xnor U21106 (N_21106,N_19636,N_20222);
or U21107 (N_21107,N_19717,N_19489);
or U21108 (N_21108,N_19577,N_20112);
and U21109 (N_21109,N_19967,N_20094);
nand U21110 (N_21110,N_19821,N_19601);
or U21111 (N_21111,N_19327,N_20170);
and U21112 (N_21112,N_19843,N_20179);
or U21113 (N_21113,N_19976,N_19431);
and U21114 (N_21114,N_20363,N_19839);
and U21115 (N_21115,N_19954,N_19235);
nand U21116 (N_21116,N_20079,N_19343);
nand U21117 (N_21117,N_20339,N_19483);
and U21118 (N_21118,N_19777,N_19470);
or U21119 (N_21119,N_19938,N_19202);
nand U21120 (N_21120,N_19733,N_19521);
xnor U21121 (N_21121,N_19702,N_19435);
or U21122 (N_21122,N_19491,N_19839);
xor U21123 (N_21123,N_19896,N_19673);
nand U21124 (N_21124,N_19923,N_20345);
and U21125 (N_21125,N_19361,N_19629);
or U21126 (N_21126,N_20066,N_19601);
xnor U21127 (N_21127,N_19901,N_20295);
nand U21128 (N_21128,N_19390,N_19612);
xor U21129 (N_21129,N_19361,N_19265);
nor U21130 (N_21130,N_20332,N_20256);
nor U21131 (N_21131,N_19649,N_19856);
and U21132 (N_21132,N_20005,N_19924);
nand U21133 (N_21133,N_19411,N_20078);
and U21134 (N_21134,N_19783,N_20016);
and U21135 (N_21135,N_19821,N_19246);
xor U21136 (N_21136,N_19627,N_20124);
or U21137 (N_21137,N_19294,N_19910);
nor U21138 (N_21138,N_20201,N_19902);
or U21139 (N_21139,N_20065,N_20070);
nor U21140 (N_21140,N_19323,N_20060);
nor U21141 (N_21141,N_19934,N_19809);
and U21142 (N_21142,N_19229,N_19754);
nor U21143 (N_21143,N_20323,N_20148);
nand U21144 (N_21144,N_19502,N_19832);
nor U21145 (N_21145,N_19497,N_19733);
nand U21146 (N_21146,N_20208,N_19303);
or U21147 (N_21147,N_19917,N_19772);
or U21148 (N_21148,N_20008,N_19816);
and U21149 (N_21149,N_19802,N_19231);
and U21150 (N_21150,N_19794,N_19752);
nand U21151 (N_21151,N_20193,N_20179);
nor U21152 (N_21152,N_20072,N_19572);
nand U21153 (N_21153,N_20021,N_20397);
nor U21154 (N_21154,N_20348,N_20195);
xnor U21155 (N_21155,N_20324,N_19358);
nor U21156 (N_21156,N_19861,N_20053);
nor U21157 (N_21157,N_19818,N_19932);
or U21158 (N_21158,N_20364,N_19259);
nor U21159 (N_21159,N_19591,N_19785);
and U21160 (N_21160,N_19963,N_20329);
xnor U21161 (N_21161,N_20101,N_19856);
nand U21162 (N_21162,N_19420,N_19246);
xor U21163 (N_21163,N_19822,N_19503);
and U21164 (N_21164,N_19702,N_19707);
nor U21165 (N_21165,N_19832,N_20154);
xnor U21166 (N_21166,N_20197,N_19508);
and U21167 (N_21167,N_20179,N_19754);
or U21168 (N_21168,N_20222,N_19625);
nand U21169 (N_21169,N_20279,N_19785);
xor U21170 (N_21170,N_19602,N_19649);
nor U21171 (N_21171,N_20018,N_19933);
and U21172 (N_21172,N_19429,N_20108);
nor U21173 (N_21173,N_19473,N_20374);
or U21174 (N_21174,N_19410,N_19454);
nand U21175 (N_21175,N_19220,N_19725);
nor U21176 (N_21176,N_19548,N_20101);
or U21177 (N_21177,N_19307,N_19896);
and U21178 (N_21178,N_19461,N_19907);
nand U21179 (N_21179,N_20186,N_19505);
nand U21180 (N_21180,N_19763,N_20348);
nor U21181 (N_21181,N_20162,N_20294);
or U21182 (N_21182,N_19508,N_19790);
nand U21183 (N_21183,N_19722,N_20276);
and U21184 (N_21184,N_19216,N_20092);
or U21185 (N_21185,N_20277,N_20000);
xnor U21186 (N_21186,N_19492,N_19898);
nor U21187 (N_21187,N_19497,N_19665);
nor U21188 (N_21188,N_19830,N_19869);
nand U21189 (N_21189,N_20100,N_20068);
xnor U21190 (N_21190,N_19835,N_19755);
nand U21191 (N_21191,N_20192,N_19752);
nand U21192 (N_21192,N_20131,N_19686);
or U21193 (N_21193,N_19942,N_19714);
nand U21194 (N_21194,N_19889,N_19925);
xnor U21195 (N_21195,N_19312,N_19920);
xor U21196 (N_21196,N_19828,N_19680);
nor U21197 (N_21197,N_19295,N_19902);
and U21198 (N_21198,N_20066,N_19442);
nor U21199 (N_21199,N_19533,N_19717);
xor U21200 (N_21200,N_20285,N_20058);
xnor U21201 (N_21201,N_19279,N_19308);
and U21202 (N_21202,N_19238,N_20301);
nor U21203 (N_21203,N_19342,N_20362);
xnor U21204 (N_21204,N_19263,N_20316);
xnor U21205 (N_21205,N_19967,N_19648);
nor U21206 (N_21206,N_19338,N_19238);
nand U21207 (N_21207,N_19684,N_20361);
nand U21208 (N_21208,N_20271,N_20266);
or U21209 (N_21209,N_20349,N_19201);
xor U21210 (N_21210,N_20229,N_20304);
xnor U21211 (N_21211,N_20057,N_19896);
nand U21212 (N_21212,N_19942,N_19687);
nand U21213 (N_21213,N_19912,N_19633);
and U21214 (N_21214,N_19334,N_19652);
nor U21215 (N_21215,N_19543,N_20025);
nand U21216 (N_21216,N_20259,N_20073);
nand U21217 (N_21217,N_19832,N_20198);
nand U21218 (N_21218,N_19753,N_19552);
nor U21219 (N_21219,N_19974,N_19262);
and U21220 (N_21220,N_19434,N_19582);
and U21221 (N_21221,N_19933,N_19473);
or U21222 (N_21222,N_19800,N_19444);
or U21223 (N_21223,N_19522,N_20101);
nand U21224 (N_21224,N_19681,N_19337);
nor U21225 (N_21225,N_20103,N_20062);
or U21226 (N_21226,N_19217,N_20194);
nand U21227 (N_21227,N_20218,N_20162);
and U21228 (N_21228,N_19218,N_20141);
and U21229 (N_21229,N_19517,N_19850);
nor U21230 (N_21230,N_19798,N_19415);
and U21231 (N_21231,N_19456,N_19782);
or U21232 (N_21232,N_19358,N_20238);
xor U21233 (N_21233,N_20023,N_19874);
nand U21234 (N_21234,N_19553,N_20020);
xnor U21235 (N_21235,N_19688,N_20146);
nand U21236 (N_21236,N_19728,N_19393);
xnor U21237 (N_21237,N_19484,N_19324);
nor U21238 (N_21238,N_20080,N_20310);
xnor U21239 (N_21239,N_19756,N_20141);
or U21240 (N_21240,N_20132,N_20399);
nand U21241 (N_21241,N_19628,N_20280);
nand U21242 (N_21242,N_19282,N_20340);
or U21243 (N_21243,N_19715,N_19490);
nand U21244 (N_21244,N_19507,N_19919);
nor U21245 (N_21245,N_20281,N_19427);
nand U21246 (N_21246,N_20226,N_19903);
xor U21247 (N_21247,N_19917,N_19208);
xor U21248 (N_21248,N_20310,N_19337);
and U21249 (N_21249,N_19777,N_20245);
nand U21250 (N_21250,N_20133,N_19488);
xor U21251 (N_21251,N_20302,N_19439);
nand U21252 (N_21252,N_20208,N_19291);
and U21253 (N_21253,N_19592,N_20093);
and U21254 (N_21254,N_19307,N_20148);
nand U21255 (N_21255,N_19641,N_19790);
or U21256 (N_21256,N_20163,N_19290);
nand U21257 (N_21257,N_19206,N_19357);
or U21258 (N_21258,N_20361,N_20114);
and U21259 (N_21259,N_19488,N_19951);
nor U21260 (N_21260,N_19987,N_19380);
and U21261 (N_21261,N_19869,N_20193);
nor U21262 (N_21262,N_19218,N_19978);
nand U21263 (N_21263,N_19946,N_20112);
nand U21264 (N_21264,N_20093,N_19336);
or U21265 (N_21265,N_19656,N_20366);
nand U21266 (N_21266,N_19217,N_19211);
xnor U21267 (N_21267,N_19561,N_20074);
or U21268 (N_21268,N_20144,N_20054);
nand U21269 (N_21269,N_19891,N_19317);
xor U21270 (N_21270,N_20030,N_19300);
or U21271 (N_21271,N_19518,N_19700);
or U21272 (N_21272,N_19371,N_19949);
xor U21273 (N_21273,N_19237,N_19547);
nand U21274 (N_21274,N_20157,N_20100);
or U21275 (N_21275,N_20285,N_20078);
nor U21276 (N_21276,N_19545,N_19480);
nor U21277 (N_21277,N_20218,N_19459);
nand U21278 (N_21278,N_19477,N_19391);
or U21279 (N_21279,N_20171,N_20205);
or U21280 (N_21280,N_20340,N_20109);
nand U21281 (N_21281,N_20128,N_19597);
xnor U21282 (N_21282,N_19947,N_20070);
nor U21283 (N_21283,N_19578,N_20327);
xor U21284 (N_21284,N_20371,N_19566);
or U21285 (N_21285,N_20069,N_19544);
nor U21286 (N_21286,N_20144,N_19945);
or U21287 (N_21287,N_19382,N_20262);
and U21288 (N_21288,N_19361,N_19496);
nand U21289 (N_21289,N_19808,N_19457);
nor U21290 (N_21290,N_20294,N_20006);
and U21291 (N_21291,N_19853,N_20064);
or U21292 (N_21292,N_20101,N_19917);
xnor U21293 (N_21293,N_19935,N_20094);
nor U21294 (N_21294,N_19867,N_19240);
or U21295 (N_21295,N_19518,N_19436);
nand U21296 (N_21296,N_19234,N_19607);
or U21297 (N_21297,N_19329,N_19507);
nor U21298 (N_21298,N_20236,N_19821);
and U21299 (N_21299,N_19242,N_20325);
nor U21300 (N_21300,N_19784,N_19309);
nor U21301 (N_21301,N_19525,N_19288);
xor U21302 (N_21302,N_19676,N_19441);
xor U21303 (N_21303,N_19268,N_19315);
nor U21304 (N_21304,N_19639,N_19755);
and U21305 (N_21305,N_20247,N_19920);
and U21306 (N_21306,N_19458,N_19435);
xnor U21307 (N_21307,N_19444,N_19387);
xnor U21308 (N_21308,N_19607,N_20115);
and U21309 (N_21309,N_19252,N_20207);
and U21310 (N_21310,N_19450,N_19469);
and U21311 (N_21311,N_19914,N_19240);
nor U21312 (N_21312,N_19760,N_19455);
or U21313 (N_21313,N_19835,N_19973);
and U21314 (N_21314,N_19319,N_19304);
xnor U21315 (N_21315,N_19342,N_19858);
nor U21316 (N_21316,N_20260,N_19552);
xnor U21317 (N_21317,N_19451,N_19719);
and U21318 (N_21318,N_19840,N_19974);
xnor U21319 (N_21319,N_20292,N_20052);
nand U21320 (N_21320,N_19561,N_20203);
or U21321 (N_21321,N_20297,N_19781);
or U21322 (N_21322,N_19558,N_19450);
xnor U21323 (N_21323,N_19279,N_20007);
xnor U21324 (N_21324,N_19239,N_19974);
or U21325 (N_21325,N_19446,N_20099);
xor U21326 (N_21326,N_19659,N_19808);
nor U21327 (N_21327,N_19409,N_19977);
and U21328 (N_21328,N_19652,N_20324);
xnor U21329 (N_21329,N_19536,N_19460);
and U21330 (N_21330,N_19942,N_20247);
nor U21331 (N_21331,N_19723,N_19295);
nand U21332 (N_21332,N_19650,N_19527);
nor U21333 (N_21333,N_19332,N_19484);
and U21334 (N_21334,N_19775,N_19666);
nor U21335 (N_21335,N_20087,N_19982);
nand U21336 (N_21336,N_19766,N_20292);
and U21337 (N_21337,N_19396,N_19723);
nor U21338 (N_21338,N_20011,N_19219);
nand U21339 (N_21339,N_19374,N_20273);
xnor U21340 (N_21340,N_20025,N_19560);
or U21341 (N_21341,N_19625,N_20057);
and U21342 (N_21342,N_19883,N_20199);
nand U21343 (N_21343,N_19552,N_19641);
nand U21344 (N_21344,N_19843,N_19236);
and U21345 (N_21345,N_20397,N_20094);
or U21346 (N_21346,N_19800,N_19878);
or U21347 (N_21347,N_19602,N_19435);
nand U21348 (N_21348,N_20299,N_19472);
and U21349 (N_21349,N_19541,N_19516);
and U21350 (N_21350,N_19391,N_19640);
nand U21351 (N_21351,N_20010,N_19242);
and U21352 (N_21352,N_19270,N_19699);
and U21353 (N_21353,N_19632,N_20349);
or U21354 (N_21354,N_19626,N_20142);
xnor U21355 (N_21355,N_19870,N_20328);
and U21356 (N_21356,N_20175,N_20018);
xnor U21357 (N_21357,N_19919,N_19385);
nand U21358 (N_21358,N_19301,N_19562);
xor U21359 (N_21359,N_19589,N_20343);
nand U21360 (N_21360,N_19251,N_20322);
or U21361 (N_21361,N_19326,N_19777);
and U21362 (N_21362,N_20002,N_19654);
nor U21363 (N_21363,N_19665,N_20297);
xnor U21364 (N_21364,N_20141,N_19328);
and U21365 (N_21365,N_20128,N_19497);
xnor U21366 (N_21366,N_19806,N_19793);
nor U21367 (N_21367,N_19914,N_19310);
or U21368 (N_21368,N_19701,N_19602);
and U21369 (N_21369,N_19765,N_20041);
xnor U21370 (N_21370,N_20227,N_19676);
nand U21371 (N_21371,N_19462,N_19402);
or U21372 (N_21372,N_20222,N_20009);
or U21373 (N_21373,N_19744,N_19644);
and U21374 (N_21374,N_19508,N_20381);
xnor U21375 (N_21375,N_19325,N_19733);
nor U21376 (N_21376,N_19436,N_19308);
and U21377 (N_21377,N_19276,N_19632);
and U21378 (N_21378,N_19638,N_20245);
nand U21379 (N_21379,N_19315,N_19537);
nand U21380 (N_21380,N_20182,N_20280);
xnor U21381 (N_21381,N_20058,N_19479);
xor U21382 (N_21382,N_20266,N_19380);
xnor U21383 (N_21383,N_19550,N_19945);
and U21384 (N_21384,N_19649,N_20063);
and U21385 (N_21385,N_19521,N_20317);
xnor U21386 (N_21386,N_20067,N_19242);
nand U21387 (N_21387,N_19418,N_20315);
and U21388 (N_21388,N_19581,N_19823);
and U21389 (N_21389,N_19389,N_19597);
xnor U21390 (N_21390,N_20266,N_19597);
and U21391 (N_21391,N_20152,N_20294);
and U21392 (N_21392,N_20093,N_19265);
or U21393 (N_21393,N_19505,N_19226);
or U21394 (N_21394,N_19844,N_20148);
or U21395 (N_21395,N_20012,N_19550);
nor U21396 (N_21396,N_19404,N_19487);
and U21397 (N_21397,N_20379,N_19639);
nor U21398 (N_21398,N_19408,N_19399);
and U21399 (N_21399,N_20248,N_20392);
nor U21400 (N_21400,N_19373,N_19815);
xor U21401 (N_21401,N_20348,N_19880);
xor U21402 (N_21402,N_19746,N_19907);
and U21403 (N_21403,N_19207,N_19405);
and U21404 (N_21404,N_20264,N_19782);
xor U21405 (N_21405,N_19596,N_20024);
nor U21406 (N_21406,N_19446,N_20344);
nor U21407 (N_21407,N_19713,N_19912);
or U21408 (N_21408,N_19311,N_19234);
nor U21409 (N_21409,N_19958,N_19205);
and U21410 (N_21410,N_20394,N_19997);
or U21411 (N_21411,N_19884,N_19734);
nor U21412 (N_21412,N_19731,N_20342);
nor U21413 (N_21413,N_19973,N_19988);
nor U21414 (N_21414,N_20344,N_19718);
xor U21415 (N_21415,N_19440,N_19508);
nand U21416 (N_21416,N_19560,N_19469);
and U21417 (N_21417,N_19996,N_20313);
xnor U21418 (N_21418,N_19643,N_19990);
nor U21419 (N_21419,N_20310,N_20095);
nor U21420 (N_21420,N_19915,N_20074);
and U21421 (N_21421,N_19858,N_19922);
or U21422 (N_21422,N_19805,N_19427);
or U21423 (N_21423,N_20315,N_20046);
nor U21424 (N_21424,N_19230,N_19917);
xnor U21425 (N_21425,N_19861,N_20186);
nor U21426 (N_21426,N_20066,N_19263);
nor U21427 (N_21427,N_19227,N_19342);
xor U21428 (N_21428,N_20014,N_19981);
xnor U21429 (N_21429,N_19243,N_20196);
or U21430 (N_21430,N_19627,N_20255);
or U21431 (N_21431,N_19328,N_20253);
nor U21432 (N_21432,N_19787,N_19684);
or U21433 (N_21433,N_19535,N_20026);
nand U21434 (N_21434,N_19229,N_19490);
xnor U21435 (N_21435,N_19490,N_19705);
nor U21436 (N_21436,N_19221,N_19474);
nand U21437 (N_21437,N_19342,N_20044);
and U21438 (N_21438,N_19421,N_20341);
nand U21439 (N_21439,N_20138,N_19700);
nand U21440 (N_21440,N_19646,N_19748);
nor U21441 (N_21441,N_19631,N_19267);
nor U21442 (N_21442,N_19512,N_20310);
and U21443 (N_21443,N_19551,N_19399);
or U21444 (N_21444,N_20248,N_19308);
and U21445 (N_21445,N_20008,N_19226);
and U21446 (N_21446,N_20094,N_19215);
nand U21447 (N_21447,N_19595,N_19643);
xor U21448 (N_21448,N_19296,N_19964);
nor U21449 (N_21449,N_19971,N_19461);
nor U21450 (N_21450,N_19376,N_19367);
or U21451 (N_21451,N_20016,N_20199);
nand U21452 (N_21452,N_19627,N_20045);
and U21453 (N_21453,N_19807,N_19859);
nor U21454 (N_21454,N_20258,N_19493);
or U21455 (N_21455,N_19438,N_19674);
and U21456 (N_21456,N_20132,N_19202);
or U21457 (N_21457,N_19200,N_19835);
or U21458 (N_21458,N_20121,N_19301);
nand U21459 (N_21459,N_19758,N_19221);
xnor U21460 (N_21460,N_19237,N_19979);
xor U21461 (N_21461,N_19381,N_20391);
or U21462 (N_21462,N_19604,N_19257);
nand U21463 (N_21463,N_19566,N_19614);
and U21464 (N_21464,N_19691,N_19646);
and U21465 (N_21465,N_19761,N_20009);
or U21466 (N_21466,N_20260,N_19309);
and U21467 (N_21467,N_19893,N_19818);
nand U21468 (N_21468,N_20169,N_20124);
nand U21469 (N_21469,N_19343,N_19589);
nand U21470 (N_21470,N_19593,N_19286);
xor U21471 (N_21471,N_19510,N_20013);
nand U21472 (N_21472,N_20092,N_20214);
or U21473 (N_21473,N_19567,N_19250);
and U21474 (N_21474,N_19333,N_19673);
and U21475 (N_21475,N_19927,N_19626);
nor U21476 (N_21476,N_19825,N_19439);
and U21477 (N_21477,N_20096,N_20147);
and U21478 (N_21478,N_20333,N_19770);
xnor U21479 (N_21479,N_20069,N_20379);
xnor U21480 (N_21480,N_19793,N_19386);
and U21481 (N_21481,N_19684,N_19927);
nand U21482 (N_21482,N_19823,N_19923);
or U21483 (N_21483,N_19431,N_20358);
or U21484 (N_21484,N_19839,N_19702);
xor U21485 (N_21485,N_19621,N_20225);
xnor U21486 (N_21486,N_19345,N_19552);
nor U21487 (N_21487,N_20030,N_19221);
nor U21488 (N_21488,N_20013,N_19591);
xnor U21489 (N_21489,N_19215,N_19655);
xor U21490 (N_21490,N_19824,N_20073);
xnor U21491 (N_21491,N_20151,N_19536);
or U21492 (N_21492,N_20007,N_19980);
nand U21493 (N_21493,N_20112,N_19903);
nand U21494 (N_21494,N_19943,N_20369);
xor U21495 (N_21495,N_19464,N_19294);
xnor U21496 (N_21496,N_19865,N_19851);
or U21497 (N_21497,N_19931,N_19778);
xor U21498 (N_21498,N_20151,N_19494);
xor U21499 (N_21499,N_20270,N_19541);
nand U21500 (N_21500,N_20229,N_19659);
nor U21501 (N_21501,N_20192,N_19717);
and U21502 (N_21502,N_20373,N_19956);
xnor U21503 (N_21503,N_20150,N_20034);
nand U21504 (N_21504,N_20187,N_19879);
or U21505 (N_21505,N_19895,N_19752);
nor U21506 (N_21506,N_19921,N_20268);
and U21507 (N_21507,N_19318,N_19456);
nand U21508 (N_21508,N_19396,N_19961);
nand U21509 (N_21509,N_19725,N_19259);
or U21510 (N_21510,N_19246,N_19355);
or U21511 (N_21511,N_19457,N_20331);
and U21512 (N_21512,N_19423,N_19489);
and U21513 (N_21513,N_20216,N_19400);
or U21514 (N_21514,N_20290,N_19309);
xor U21515 (N_21515,N_19724,N_19474);
nand U21516 (N_21516,N_20227,N_19261);
nand U21517 (N_21517,N_19217,N_19291);
xnor U21518 (N_21518,N_19671,N_19221);
and U21519 (N_21519,N_19412,N_19748);
nand U21520 (N_21520,N_20013,N_19451);
or U21521 (N_21521,N_19248,N_19289);
nor U21522 (N_21522,N_19490,N_19916);
nor U21523 (N_21523,N_20241,N_19322);
nand U21524 (N_21524,N_20049,N_19816);
or U21525 (N_21525,N_19603,N_20253);
xnor U21526 (N_21526,N_20109,N_19725);
nor U21527 (N_21527,N_20045,N_19354);
and U21528 (N_21528,N_19708,N_20182);
and U21529 (N_21529,N_20349,N_19968);
nand U21530 (N_21530,N_20270,N_19236);
nand U21531 (N_21531,N_20132,N_19641);
and U21532 (N_21532,N_20308,N_19988);
and U21533 (N_21533,N_19403,N_19583);
and U21534 (N_21534,N_20205,N_19499);
nand U21535 (N_21535,N_20206,N_19773);
and U21536 (N_21536,N_20299,N_19946);
and U21537 (N_21537,N_19996,N_19540);
nand U21538 (N_21538,N_19445,N_19555);
nand U21539 (N_21539,N_19788,N_20119);
nand U21540 (N_21540,N_19370,N_19820);
or U21541 (N_21541,N_20369,N_20263);
or U21542 (N_21542,N_19774,N_19710);
nand U21543 (N_21543,N_19723,N_20154);
and U21544 (N_21544,N_19686,N_19516);
nor U21545 (N_21545,N_19641,N_19780);
nor U21546 (N_21546,N_19211,N_20307);
xor U21547 (N_21547,N_19499,N_20299);
nor U21548 (N_21548,N_19653,N_19561);
and U21549 (N_21549,N_20237,N_20024);
and U21550 (N_21550,N_19711,N_19657);
and U21551 (N_21551,N_19449,N_20372);
or U21552 (N_21552,N_20342,N_20171);
xnor U21553 (N_21553,N_20385,N_19908);
nor U21554 (N_21554,N_19787,N_19439);
xnor U21555 (N_21555,N_19339,N_19631);
xor U21556 (N_21556,N_19448,N_20034);
or U21557 (N_21557,N_19330,N_20329);
nand U21558 (N_21558,N_20137,N_19887);
nand U21559 (N_21559,N_20256,N_19822);
or U21560 (N_21560,N_19291,N_19230);
nand U21561 (N_21561,N_19488,N_19361);
nor U21562 (N_21562,N_19659,N_20368);
and U21563 (N_21563,N_19887,N_20264);
or U21564 (N_21564,N_19514,N_20328);
nor U21565 (N_21565,N_19745,N_20373);
xor U21566 (N_21566,N_19844,N_20086);
nor U21567 (N_21567,N_20392,N_19931);
nor U21568 (N_21568,N_20191,N_19619);
and U21569 (N_21569,N_19881,N_19718);
xor U21570 (N_21570,N_19560,N_19262);
and U21571 (N_21571,N_19494,N_19598);
or U21572 (N_21572,N_19556,N_19926);
nand U21573 (N_21573,N_20288,N_20312);
nand U21574 (N_21574,N_19987,N_19718);
nor U21575 (N_21575,N_20041,N_19538);
xnor U21576 (N_21576,N_19594,N_20290);
nand U21577 (N_21577,N_20089,N_19986);
xor U21578 (N_21578,N_19445,N_19399);
and U21579 (N_21579,N_19648,N_19820);
nand U21580 (N_21580,N_19907,N_19781);
xnor U21581 (N_21581,N_20122,N_20343);
or U21582 (N_21582,N_19502,N_19889);
nor U21583 (N_21583,N_19394,N_20089);
xnor U21584 (N_21584,N_19950,N_19577);
nand U21585 (N_21585,N_19688,N_19433);
xnor U21586 (N_21586,N_19740,N_20317);
nand U21587 (N_21587,N_20247,N_19552);
nand U21588 (N_21588,N_19600,N_20013);
nand U21589 (N_21589,N_20182,N_20188);
xor U21590 (N_21590,N_19967,N_19578);
and U21591 (N_21591,N_19502,N_19492);
nand U21592 (N_21592,N_19755,N_20022);
xnor U21593 (N_21593,N_19397,N_19887);
nand U21594 (N_21594,N_19349,N_19799);
or U21595 (N_21595,N_19586,N_19489);
xor U21596 (N_21596,N_19790,N_19377);
xnor U21597 (N_21597,N_19661,N_20277);
and U21598 (N_21598,N_19722,N_19963);
or U21599 (N_21599,N_19269,N_19828);
xor U21600 (N_21600,N_21541,N_21228);
xor U21601 (N_21601,N_20415,N_21148);
nor U21602 (N_21602,N_21050,N_20629);
xor U21603 (N_21603,N_21127,N_21464);
xnor U21604 (N_21604,N_20738,N_20481);
and U21605 (N_21605,N_20659,N_21491);
xnor U21606 (N_21606,N_21255,N_21135);
xnor U21607 (N_21607,N_21471,N_20803);
nor U21608 (N_21608,N_21022,N_20864);
nor U21609 (N_21609,N_21566,N_20714);
and U21610 (N_21610,N_21118,N_21174);
and U21611 (N_21611,N_20882,N_20939);
xor U21612 (N_21612,N_20911,N_20751);
xor U21613 (N_21613,N_20463,N_20887);
xnor U21614 (N_21614,N_21121,N_20908);
or U21615 (N_21615,N_20573,N_21401);
xor U21616 (N_21616,N_21262,N_20971);
or U21617 (N_21617,N_20792,N_21529);
nor U21618 (N_21618,N_21131,N_20921);
and U21619 (N_21619,N_21216,N_21545);
or U21620 (N_21620,N_21247,N_21291);
xnor U21621 (N_21621,N_20757,N_20853);
and U21622 (N_21622,N_20407,N_20692);
and U21623 (N_21623,N_20974,N_21501);
and U21624 (N_21624,N_20427,N_20733);
nand U21625 (N_21625,N_21152,N_20471);
nor U21626 (N_21626,N_21368,N_21272);
or U21627 (N_21627,N_21147,N_20483);
nand U21628 (N_21628,N_20851,N_20867);
xnor U21629 (N_21629,N_21017,N_21108);
xor U21630 (N_21630,N_21018,N_21385);
or U21631 (N_21631,N_21354,N_20615);
or U21632 (N_21632,N_21151,N_20500);
xor U21633 (N_21633,N_20596,N_20540);
xor U21634 (N_21634,N_21286,N_21473);
or U21635 (N_21635,N_21078,N_20591);
nor U21636 (N_21636,N_21067,N_21163);
nand U21637 (N_21637,N_20608,N_20409);
nand U21638 (N_21638,N_21103,N_21096);
nor U21639 (N_21639,N_21425,N_21371);
xor U21640 (N_21640,N_20616,N_20889);
xor U21641 (N_21641,N_21577,N_20750);
and U21642 (N_21642,N_21249,N_21170);
and U21643 (N_21643,N_20675,N_21155);
or U21644 (N_21644,N_21567,N_20775);
xor U21645 (N_21645,N_21191,N_21474);
nor U21646 (N_21646,N_20571,N_21421);
xnor U21647 (N_21647,N_20744,N_21455);
or U21648 (N_21648,N_21012,N_20532);
nand U21649 (N_21649,N_21408,N_21362);
xor U21650 (N_21650,N_21063,N_20606);
nand U21651 (N_21651,N_21231,N_20612);
xnor U21652 (N_21652,N_20888,N_21429);
nor U21653 (N_21653,N_21102,N_20569);
nor U21654 (N_21654,N_20490,N_21356);
nand U21655 (N_21655,N_21350,N_20900);
xor U21656 (N_21656,N_20735,N_20802);
xor U21657 (N_21657,N_21260,N_20949);
nand U21658 (N_21658,N_21119,N_20998);
and U21659 (N_21659,N_20894,N_20437);
and U21660 (N_21660,N_20979,N_21418);
and U21661 (N_21661,N_21046,N_20715);
or U21662 (N_21662,N_20996,N_20443);
nand U21663 (N_21663,N_20458,N_20712);
and U21664 (N_21664,N_21482,N_21070);
and U21665 (N_21665,N_21332,N_21523);
nand U21666 (N_21666,N_20776,N_21279);
xor U21667 (N_21667,N_21428,N_21261);
nor U21668 (N_21668,N_21171,N_20574);
or U21669 (N_21669,N_21192,N_21179);
nand U21670 (N_21670,N_21109,N_21056);
nor U21671 (N_21671,N_20972,N_21485);
nor U21672 (N_21672,N_21316,N_20405);
or U21673 (N_21673,N_21410,N_21466);
or U21674 (N_21674,N_20603,N_21568);
nand U21675 (N_21675,N_20997,N_20788);
nand U21676 (N_21676,N_20565,N_21374);
xor U21677 (N_21677,N_21513,N_20594);
nand U21678 (N_21678,N_21288,N_21169);
nand U21679 (N_21679,N_20640,N_21526);
or U21680 (N_21680,N_20966,N_21312);
nor U21681 (N_21681,N_21595,N_21562);
xor U21682 (N_21682,N_21042,N_20946);
nand U21683 (N_21683,N_21413,N_20741);
nor U21684 (N_21684,N_20843,N_21598);
or U21685 (N_21685,N_21328,N_20786);
and U21686 (N_21686,N_21003,N_21185);
and U21687 (N_21687,N_21301,N_21424);
nor U21688 (N_21688,N_21481,N_20507);
xor U21689 (N_21689,N_20558,N_20819);
and U21690 (N_21690,N_20417,N_21435);
xnor U21691 (N_21691,N_21405,N_20766);
nor U21692 (N_21692,N_21539,N_21265);
and U21693 (N_21693,N_21536,N_21537);
nor U21694 (N_21694,N_20890,N_20456);
and U21695 (N_21695,N_21433,N_21584);
nand U21696 (N_21696,N_20736,N_20893);
xor U21697 (N_21697,N_20680,N_21549);
and U21698 (N_21698,N_20431,N_20572);
xnor U21699 (N_21699,N_21086,N_20812);
or U21700 (N_21700,N_21520,N_20805);
nand U21701 (N_21701,N_21285,N_20948);
or U21702 (N_21702,N_20761,N_21190);
nor U21703 (N_21703,N_20722,N_21394);
and U21704 (N_21704,N_21519,N_21334);
or U21705 (N_21705,N_20925,N_20632);
xor U21706 (N_21706,N_20600,N_21033);
or U21707 (N_21707,N_20713,N_21074);
nor U21708 (N_21708,N_20570,N_21547);
and U21709 (N_21709,N_21194,N_20683);
and U21710 (N_21710,N_21061,N_20917);
nor U21711 (N_21711,N_20672,N_20447);
nand U21712 (N_21712,N_20716,N_20418);
xor U21713 (N_21713,N_21300,N_21069);
nor U21714 (N_21714,N_21092,N_20771);
nor U21715 (N_21715,N_21530,N_21227);
nand U21716 (N_21716,N_20462,N_20541);
or U21717 (N_21717,N_20476,N_21158);
xnor U21718 (N_21718,N_20673,N_20414);
xnor U21719 (N_21719,N_21237,N_20486);
and U21720 (N_21720,N_20701,N_21202);
or U21721 (N_21721,N_20633,N_20472);
and U21722 (N_21722,N_20995,N_21367);
nand U21723 (N_21723,N_21244,N_21306);
nor U21724 (N_21724,N_21098,N_20793);
or U21725 (N_21725,N_20860,N_20953);
nand U21726 (N_21726,N_21437,N_20937);
or U21727 (N_21727,N_20724,N_21522);
xnor U21728 (N_21728,N_21207,N_21273);
and U21729 (N_21729,N_20556,N_21357);
nand U21730 (N_21730,N_21318,N_20576);
and U21731 (N_21731,N_20808,N_20625);
or U21732 (N_21732,N_21383,N_20469);
or U21733 (N_21733,N_20601,N_21477);
and U21734 (N_21734,N_20526,N_21309);
or U21735 (N_21735,N_21442,N_21351);
or U21736 (N_21736,N_21591,N_21507);
xnor U21737 (N_21737,N_20833,N_21219);
nand U21738 (N_21738,N_21540,N_20696);
nand U21739 (N_21739,N_20797,N_20992);
and U21740 (N_21740,N_20484,N_20988);
and U21741 (N_21741,N_20678,N_21426);
and U21742 (N_21742,N_20538,N_20627);
or U21743 (N_21743,N_21387,N_21274);
and U21744 (N_21744,N_21439,N_21082);
or U21745 (N_21745,N_20912,N_20823);
xor U21746 (N_21746,N_21494,N_20896);
or U21747 (N_21747,N_21006,N_21326);
xnor U21748 (N_21748,N_21596,N_20674);
xnor U21749 (N_21749,N_20957,N_21499);
and U21750 (N_21750,N_21027,N_21456);
xor U21751 (N_21751,N_21248,N_21110);
nand U21752 (N_21752,N_20461,N_20589);
and U21753 (N_21753,N_20487,N_21432);
nor U21754 (N_21754,N_20906,N_21088);
nor U21755 (N_21755,N_21535,N_20991);
xnor U21756 (N_21756,N_20969,N_20813);
and U21757 (N_21757,N_21122,N_20955);
or U21758 (N_21758,N_20559,N_21370);
nor U21759 (N_21759,N_21233,N_20704);
or U21760 (N_21760,N_20563,N_20514);
and U21761 (N_21761,N_21214,N_20784);
and U21762 (N_21762,N_21176,N_21514);
or U21763 (N_21763,N_20438,N_21250);
nor U21764 (N_21764,N_20518,N_21222);
xnor U21765 (N_21765,N_21283,N_21182);
and U21766 (N_21766,N_20944,N_20497);
nor U21767 (N_21767,N_21509,N_21024);
and U21768 (N_21768,N_21565,N_20516);
xor U21769 (N_21769,N_21040,N_20650);
nand U21770 (N_21770,N_21445,N_21489);
nand U21771 (N_21771,N_20587,N_20897);
or U21772 (N_21772,N_21329,N_20468);
and U21773 (N_21773,N_21105,N_20910);
or U21774 (N_21774,N_21215,N_20816);
or U21775 (N_21775,N_21259,N_20429);
and U21776 (N_21776,N_20865,N_21314);
nand U21777 (N_21777,N_20847,N_21303);
xor U21778 (N_21778,N_21007,N_20830);
or U21779 (N_21779,N_20474,N_20475);
and U21780 (N_21780,N_20492,N_20842);
nand U21781 (N_21781,N_21353,N_20795);
nor U21782 (N_21782,N_21008,N_21266);
xor U21783 (N_21783,N_21452,N_20607);
xnor U21784 (N_21784,N_20413,N_21583);
or U21785 (N_21785,N_20857,N_20765);
nor U21786 (N_21786,N_21313,N_20705);
nand U21787 (N_21787,N_20502,N_21071);
nand U21788 (N_21788,N_20513,N_21278);
or U21789 (N_21789,N_21576,N_20654);
or U21790 (N_21790,N_21402,N_21484);
xnor U21791 (N_21791,N_21430,N_20772);
nor U21792 (N_21792,N_21159,N_21220);
and U21793 (N_21793,N_21138,N_21079);
nor U21794 (N_21794,N_21123,N_21563);
or U21795 (N_21795,N_20480,N_21443);
nand U21796 (N_21796,N_21375,N_20613);
or U21797 (N_21797,N_20598,N_21459);
and U21798 (N_21798,N_20838,N_20455);
nor U21799 (N_21799,N_21327,N_21243);
or U21800 (N_21800,N_20404,N_21156);
nand U21801 (N_21801,N_20769,N_21420);
xnor U21802 (N_21802,N_21204,N_21073);
and U21803 (N_21803,N_20872,N_21582);
nand U21804 (N_21804,N_20647,N_20835);
xor U21805 (N_21805,N_21229,N_20602);
and U21806 (N_21806,N_20543,N_21406);
or U21807 (N_21807,N_20728,N_21412);
or U21808 (N_21808,N_21095,N_20534);
and U21809 (N_21809,N_20503,N_20667);
nand U21810 (N_21810,N_20987,N_20562);
nor U21811 (N_21811,N_20903,N_21077);
nor U21812 (N_21812,N_20530,N_21113);
xnor U21813 (N_21813,N_20928,N_21487);
or U21814 (N_21814,N_20653,N_21270);
or U21815 (N_21815,N_20690,N_20536);
nor U21816 (N_21816,N_20439,N_20902);
and U21817 (N_21817,N_21427,N_21001);
xnor U21818 (N_21818,N_21005,N_20403);
nor U21819 (N_21819,N_20796,N_21524);
xnor U21820 (N_21820,N_20981,N_20986);
xnor U21821 (N_21821,N_21245,N_20552);
and U21822 (N_21822,N_20620,N_21373);
xor U21823 (N_21823,N_21500,N_20916);
and U21824 (N_21824,N_20926,N_21546);
or U21825 (N_21825,N_20510,N_21035);
nand U21826 (N_21826,N_21325,N_21302);
xor U21827 (N_21827,N_21168,N_21030);
xnor U21828 (N_21828,N_21052,N_21101);
xnor U21829 (N_21829,N_21396,N_20764);
or U21830 (N_21830,N_21308,N_20436);
or U21831 (N_21831,N_20555,N_20913);
nand U21832 (N_21832,N_20901,N_21454);
nor U21833 (N_21833,N_20762,N_21355);
or U21834 (N_21834,N_20718,N_21269);
nor U21835 (N_21835,N_20952,N_21049);
nor U21836 (N_21836,N_21256,N_21587);
xnor U21837 (N_21837,N_20548,N_21180);
nor U21838 (N_21838,N_21000,N_20852);
nor U21839 (N_21839,N_20945,N_21034);
nor U21840 (N_21840,N_20628,N_21187);
xor U21841 (N_21841,N_21496,N_20870);
and U21842 (N_21842,N_21107,N_20664);
nor U21843 (N_21843,N_21146,N_21076);
or U21844 (N_21844,N_20482,N_20978);
nand U21845 (N_21845,N_20609,N_20670);
xor U21846 (N_21846,N_21493,N_20660);
nand U21847 (N_21847,N_21065,N_21381);
xor U21848 (N_21848,N_20557,N_20528);
nor U21849 (N_21849,N_21142,N_21495);
xor U21850 (N_21850,N_20631,N_20809);
nor U21851 (N_21851,N_20723,N_20621);
nor U21852 (N_21852,N_21114,N_20535);
nor U21853 (N_21853,N_21388,N_21206);
xor U21854 (N_21854,N_21297,N_20959);
nor U21855 (N_21855,N_20515,N_20963);
nor U21856 (N_21856,N_21166,N_21343);
and U21857 (N_21857,N_20801,N_21289);
nand U21858 (N_21858,N_20420,N_20970);
nand U21859 (N_21859,N_21497,N_21465);
nor U21860 (N_21860,N_21483,N_20410);
nor U21861 (N_21861,N_21311,N_20467);
or U21862 (N_21862,N_21181,N_20743);
nand U21863 (N_21863,N_20505,N_21199);
or U21864 (N_21864,N_21136,N_21277);
and U21865 (N_21865,N_20459,N_20798);
xor U21866 (N_21866,N_21440,N_21010);
nand U21867 (N_21867,N_21450,N_21157);
nor U21868 (N_21868,N_20539,N_21039);
and U21869 (N_21869,N_20691,N_21223);
or U21870 (N_21870,N_21060,N_20524);
or U21871 (N_21871,N_21287,N_21338);
and U21872 (N_21872,N_20779,N_21559);
xor U21873 (N_21873,N_21246,N_20432);
nand U21874 (N_21874,N_21209,N_21324);
xnor U21875 (N_21875,N_21436,N_21478);
or U21876 (N_21876,N_20422,N_20841);
nand U21877 (N_21877,N_20639,N_21134);
nand U21878 (N_21878,N_20523,N_21153);
xor U21879 (N_21879,N_21208,N_20730);
xor U21880 (N_21880,N_21239,N_21543);
and U21881 (N_21881,N_21363,N_20840);
or U21882 (N_21882,N_20700,N_21139);
xnor U21883 (N_21883,N_21475,N_21575);
and U21884 (N_21884,N_21143,N_21461);
nor U21885 (N_21885,N_21032,N_20419);
xor U21886 (N_21886,N_21218,N_20470);
nor U21887 (N_21887,N_20734,N_20520);
or U21888 (N_21888,N_20837,N_21469);
nand U21889 (N_21889,N_20745,N_20582);
nand U21890 (N_21890,N_21479,N_21556);
or U21891 (N_21891,N_21048,N_21282);
nand U21892 (N_21892,N_20618,N_21083);
xnor U21893 (N_21893,N_21062,N_20876);
nand U21894 (N_21894,N_20960,N_21149);
nand U21895 (N_21895,N_21066,N_20810);
nor U21896 (N_21896,N_20477,N_21037);
and U21897 (N_21897,N_20811,N_20623);
or U21898 (N_21898,N_21054,N_21460);
xor U21899 (N_21899,N_21293,N_21574);
xor U21900 (N_21900,N_20521,N_20923);
xor U21901 (N_21901,N_20711,N_20662);
or U21902 (N_21902,N_20531,N_20693);
or U21903 (N_21903,N_20435,N_21593);
and U21904 (N_21904,N_20434,N_21415);
xor U21905 (N_21905,N_20780,N_20815);
nor U21906 (N_21906,N_21296,N_20428);
or U21907 (N_21907,N_21570,N_20465);
nand U21908 (N_21908,N_21364,N_20554);
xnor U21909 (N_21909,N_21226,N_21389);
nor U21910 (N_21910,N_20655,N_20832);
xor U21911 (N_21911,N_20827,N_20657);
nand U21912 (N_21912,N_21064,N_20892);
and U21913 (N_21913,N_20644,N_21145);
or U21914 (N_21914,N_20433,N_20989);
nand U21915 (N_21915,N_20578,N_20982);
xnor U21916 (N_21916,N_21085,N_21112);
or U21917 (N_21917,N_21586,N_21038);
xor U21918 (N_21918,N_20599,N_20707);
or U21919 (N_21919,N_20643,N_20994);
or U21920 (N_21920,N_20583,N_21133);
nand U21921 (N_21921,N_20777,N_21120);
nand U21922 (N_21922,N_21104,N_20512);
xnor U21923 (N_21923,N_20854,N_20703);
or U21924 (N_21924,N_21476,N_21451);
or U21925 (N_21925,N_21011,N_20421);
nand U21926 (N_21926,N_20710,N_21594);
xnor U21927 (N_21927,N_20983,N_20499);
xnor U21928 (N_21928,N_21203,N_20590);
and U21929 (N_21929,N_20423,N_21407);
and U21930 (N_21930,N_20856,N_20965);
or U21931 (N_21931,N_20624,N_21013);
xor U21932 (N_21932,N_20742,N_20767);
and U21933 (N_21933,N_20758,N_20855);
nor U21934 (N_21934,N_21453,N_21380);
xnor U21935 (N_21935,N_21253,N_21094);
nand U21936 (N_21936,N_20498,N_20506);
or U21937 (N_21937,N_20977,N_20942);
or U21938 (N_21938,N_20586,N_20579);
nor U21939 (N_21939,N_20719,N_21264);
nor U21940 (N_21940,N_20412,N_20877);
xnor U21941 (N_21941,N_21590,N_20935);
xor U21942 (N_21942,N_20938,N_20936);
nor U21943 (N_21943,N_20649,N_21177);
xnor U21944 (N_21944,N_20951,N_20411);
xor U21945 (N_21945,N_21533,N_21555);
nand U21946 (N_21946,N_21463,N_20858);
xor U21947 (N_21947,N_21100,N_20814);
nor U21948 (N_21948,N_21553,N_20821);
nor U21949 (N_21949,N_21068,N_20501);
xor U21950 (N_21950,N_20879,N_20773);
or U21951 (N_21951,N_21564,N_20749);
and U21952 (N_21952,N_20478,N_21390);
or U21953 (N_21953,N_21572,N_21090);
nand U21954 (N_21954,N_20416,N_20768);
xor U21955 (N_21955,N_21538,N_21081);
nor U21956 (N_21956,N_21506,N_21267);
nor U21957 (N_21957,N_21195,N_20706);
or U21958 (N_21958,N_21305,N_20493);
nor U21959 (N_21959,N_21345,N_20676);
nor U21960 (N_21960,N_21560,N_21057);
xor U21961 (N_21961,N_21240,N_20976);
or U21962 (N_21962,N_20575,N_21234);
xnor U21963 (N_21963,N_21550,N_21201);
or U21964 (N_21964,N_20962,N_21551);
xor U21965 (N_21965,N_20922,N_21213);
and U21966 (N_21966,N_20929,N_20993);
nand U21967 (N_21967,N_20581,N_21331);
nor U21968 (N_21968,N_20895,N_20604);
nor U21969 (N_21969,N_20442,N_21045);
nor U21970 (N_21970,N_20708,N_20635);
xor U21971 (N_21971,N_21080,N_21016);
nand U21972 (N_21972,N_20485,N_21597);
xnor U21973 (N_21973,N_21409,N_21391);
or U21974 (N_21974,N_21275,N_20561);
nand U21975 (N_21975,N_21580,N_21115);
and U21976 (N_21976,N_20580,N_21292);
xor U21977 (N_21977,N_20785,N_20566);
xnor U21978 (N_21978,N_20592,N_21571);
and U21979 (N_21979,N_21480,N_21504);
nor U21980 (N_21980,N_21124,N_20460);
or U21981 (N_21981,N_21447,N_20509);
nand U21982 (N_21982,N_20905,N_20783);
nand U21983 (N_21983,N_20778,N_21026);
or U21984 (N_21984,N_20519,N_20697);
or U21985 (N_21985,N_20464,N_21554);
and U21986 (N_21986,N_21025,N_21031);
xnor U21987 (N_21987,N_20669,N_21020);
nand U21988 (N_21988,N_21585,N_20831);
nor U21989 (N_21989,N_20954,N_21150);
nand U21990 (N_21990,N_21352,N_21341);
and U21991 (N_21991,N_21360,N_20850);
or U21992 (N_21992,N_20875,N_21377);
or U21993 (N_21993,N_20898,N_21211);
xor U21994 (N_21994,N_20822,N_21236);
or U21995 (N_21995,N_20577,N_20522);
nor U21996 (N_21996,N_21014,N_20975);
and U21997 (N_21997,N_21492,N_21276);
nor U21998 (N_21998,N_20756,N_20451);
nand U21999 (N_21999,N_20448,N_21058);
nor U22000 (N_22000,N_20927,N_20863);
nor U22001 (N_22001,N_20425,N_21457);
nand U22002 (N_22002,N_20839,N_20652);
xor U22003 (N_22003,N_21470,N_20958);
nor U22004 (N_22004,N_20961,N_20637);
nor U22005 (N_22005,N_20868,N_20862);
or U22006 (N_22006,N_21335,N_20907);
nor U22007 (N_22007,N_20781,N_21393);
nand U22008 (N_22008,N_21431,N_20614);
nand U22009 (N_22009,N_20800,N_20806);
nand U22010 (N_22010,N_21392,N_20956);
nor U22011 (N_22011,N_21561,N_20844);
nand U22012 (N_22012,N_21417,N_20924);
or U22013 (N_22013,N_21111,N_21254);
nand U22014 (N_22014,N_21212,N_20651);
xnor U22015 (N_22015,N_21379,N_21449);
or U22016 (N_22016,N_21528,N_20681);
xnor U22017 (N_22017,N_21295,N_21029);
or U22018 (N_22018,N_20934,N_21330);
or U22019 (N_22019,N_21251,N_21548);
xor U22020 (N_22020,N_21041,N_21544);
and U22021 (N_22021,N_21186,N_21144);
nor U22022 (N_22022,N_20774,N_21021);
nand U22023 (N_22023,N_21106,N_20665);
and U22024 (N_22024,N_21175,N_20918);
nor U22025 (N_22025,N_20638,N_21198);
or U22026 (N_22026,N_20440,N_21339);
xnor U22027 (N_22027,N_21395,N_20904);
nand U22028 (N_22028,N_21444,N_20845);
nor U22029 (N_22029,N_21337,N_20595);
nand U22030 (N_22030,N_20914,N_21200);
nor U22031 (N_22031,N_20940,N_20537);
and U22032 (N_22032,N_21441,N_20964);
and U22033 (N_22033,N_20999,N_21304);
nor U22034 (N_22034,N_20824,N_20909);
nor U22035 (N_22035,N_21116,N_20656);
and U22036 (N_22036,N_20568,N_20545);
nand U22037 (N_22037,N_21376,N_21230);
or U22038 (N_22038,N_21252,N_20729);
nand U22039 (N_22039,N_20542,N_20426);
or U22040 (N_22040,N_20679,N_21358);
xnor U22041 (N_22041,N_21404,N_21579);
or U22042 (N_22042,N_21498,N_20817);
or U22043 (N_22043,N_20689,N_20885);
or U22044 (N_22044,N_20770,N_20611);
or U22045 (N_22045,N_20661,N_21340);
and U22046 (N_22046,N_20699,N_21322);
or U22047 (N_22047,N_21400,N_21378);
nor U22048 (N_22048,N_21023,N_20605);
and U22049 (N_22049,N_20884,N_20666);
nor U22050 (N_22050,N_21511,N_20544);
xor U22051 (N_22051,N_20932,N_20759);
nor U22052 (N_22052,N_20849,N_21342);
nand U22053 (N_22053,N_20760,N_21310);
or U22054 (N_22054,N_21055,N_20726);
or U22055 (N_22055,N_20504,N_21210);
and U22056 (N_22056,N_20799,N_21346);
nor U22057 (N_22057,N_20846,N_20702);
and U22058 (N_22058,N_21581,N_20984);
nor U22059 (N_22059,N_20630,N_20446);
xor U22060 (N_22060,N_21224,N_20682);
or U22061 (N_22061,N_21419,N_20551);
xor U22062 (N_22062,N_21004,N_21508);
or U22063 (N_22063,N_20727,N_21160);
xnor U22064 (N_22064,N_21002,N_20720);
nor U22065 (N_22065,N_21281,N_20968);
or U22066 (N_22066,N_21165,N_20457);
or U22067 (N_22067,N_20866,N_20491);
nor U22068 (N_22068,N_20930,N_20560);
nor U22069 (N_22069,N_20400,N_21438);
or U22070 (N_22070,N_21599,N_20794);
xnor U22071 (N_22071,N_20489,N_20517);
xnor U22072 (N_22072,N_20891,N_20488);
xor U22073 (N_22073,N_21414,N_20547);
and U22074 (N_22074,N_20973,N_21347);
nor U22075 (N_22075,N_20619,N_20453);
xnor U22076 (N_22076,N_21129,N_21140);
nand U22077 (N_22077,N_21384,N_20642);
and U22078 (N_22078,N_20698,N_21503);
xor U22079 (N_22079,N_21518,N_21084);
nor U22080 (N_22080,N_20444,N_20441);
xor U22081 (N_22081,N_20454,N_21172);
xor U22082 (N_22082,N_20646,N_20828);
nor U22083 (N_22083,N_21510,N_20430);
nand U22084 (N_22084,N_21532,N_21386);
xor U22085 (N_22085,N_20584,N_21557);
xor U22086 (N_22086,N_20947,N_21569);
xnor U22087 (N_22087,N_21323,N_21242);
nand U22088 (N_22088,N_21019,N_21028);
nand U22089 (N_22089,N_21137,N_21588);
nand U22090 (N_22090,N_21263,N_20445);
or U22091 (N_22091,N_21486,N_21154);
nand U22092 (N_22092,N_20466,N_21099);
or U22093 (N_22093,N_20747,N_20748);
or U22094 (N_22094,N_21189,N_21258);
xor U22095 (N_22095,N_21036,N_21531);
nor U22096 (N_22096,N_20479,N_21126);
and U22097 (N_22097,N_20826,N_21372);
nand U22098 (N_22098,N_20943,N_21197);
and U22099 (N_22099,N_21589,N_20790);
and U22100 (N_22100,N_20641,N_21205);
and U22101 (N_22101,N_21167,N_20585);
or U22102 (N_22102,N_21552,N_21221);
and U22103 (N_22103,N_20634,N_21462);
or U22104 (N_22104,N_20950,N_21044);
nand U22105 (N_22105,N_21515,N_21578);
or U22106 (N_22106,N_21294,N_21009);
nand U22107 (N_22107,N_20529,N_20804);
nand U22108 (N_22108,N_20754,N_20588);
nor U22109 (N_22109,N_20967,N_20617);
or U22110 (N_22110,N_20553,N_21361);
and U22111 (N_22111,N_21525,N_20874);
xor U22112 (N_22112,N_20402,N_20406);
and U22113 (N_22113,N_21043,N_20597);
or U22114 (N_22114,N_21117,N_21434);
nand U22115 (N_22115,N_20622,N_20687);
xor U22116 (N_22116,N_20686,N_21321);
and U22117 (N_22117,N_21299,N_20825);
and U22118 (N_22118,N_21132,N_20818);
and U22119 (N_22119,N_20546,N_20671);
xnor U22120 (N_22120,N_20648,N_21319);
or U22121 (N_22121,N_21333,N_20593);
xnor U22122 (N_22122,N_20450,N_20527);
xor U22123 (N_22123,N_21097,N_21225);
nand U22124 (N_22124,N_20834,N_20449);
nor U22125 (N_22125,N_21184,N_20740);
and U22126 (N_22126,N_20915,N_20871);
and U22127 (N_22127,N_21257,N_20549);
or U22128 (N_22128,N_21592,N_21349);
xor U22129 (N_22129,N_20886,N_20732);
nand U22130 (N_22130,N_20873,N_20985);
nor U22131 (N_22131,N_21162,N_21173);
nand U22132 (N_22132,N_20791,N_21512);
or U22133 (N_22133,N_20525,N_21521);
nor U22134 (N_22134,N_21183,N_21178);
xor U22135 (N_22135,N_20881,N_21093);
or U22136 (N_22136,N_21089,N_21467);
xnor U22137 (N_22137,N_20807,N_20645);
or U22138 (N_22138,N_21542,N_21336);
nand U22139 (N_22139,N_21403,N_20668);
xor U22140 (N_22140,N_21235,N_21307);
or U22141 (N_22141,N_21141,N_21188);
nand U22142 (N_22142,N_20752,N_20880);
xnor U22143 (N_22143,N_21558,N_20731);
nand U22144 (N_22144,N_20452,N_20980);
and U22145 (N_22145,N_20746,N_20658);
or U22146 (N_22146,N_21161,N_21369);
nor U22147 (N_22147,N_20920,N_21472);
xnor U22148 (N_22148,N_20859,N_21446);
xor U22149 (N_22149,N_20494,N_21051);
and U22150 (N_22150,N_20755,N_21366);
and U22151 (N_22151,N_20473,N_21468);
and U22152 (N_22152,N_20721,N_21458);
nor U22153 (N_22153,N_20878,N_20789);
or U22154 (N_22154,N_20883,N_21241);
or U22155 (N_22155,N_21516,N_20610);
or U22156 (N_22156,N_20694,N_21268);
nand U22157 (N_22157,N_20869,N_21284);
or U22158 (N_22158,N_20564,N_20931);
nor U22159 (N_22159,N_21075,N_20919);
nand U22160 (N_22160,N_20753,N_21348);
and U22161 (N_22161,N_20709,N_20663);
or U22162 (N_22162,N_20787,N_21365);
xor U22163 (N_22163,N_21193,N_20829);
nand U22164 (N_22164,N_21271,N_21059);
and U22165 (N_22165,N_20990,N_21164);
nor U22166 (N_22166,N_21317,N_20626);
nor U22167 (N_22167,N_20941,N_21280);
nand U22168 (N_22168,N_21047,N_20820);
xnor U22169 (N_22169,N_20401,N_21359);
or U22170 (N_22170,N_20763,N_21573);
nand U22171 (N_22171,N_21411,N_21128);
xnor U22172 (N_22172,N_21398,N_20737);
and U22173 (N_22173,N_20408,N_21232);
nand U22174 (N_22174,N_21091,N_21217);
or U22175 (N_22175,N_20836,N_21298);
xor U22176 (N_22176,N_21488,N_20567);
and U22177 (N_22177,N_21382,N_21125);
nand U22178 (N_22178,N_20685,N_21320);
nand U22179 (N_22179,N_20684,N_21505);
nor U22180 (N_22180,N_21238,N_21196);
and U22181 (N_22181,N_21399,N_21315);
xor U22182 (N_22182,N_20424,N_21397);
xor U22183 (N_22183,N_20933,N_20636);
nand U22184 (N_22184,N_20677,N_21072);
or U22185 (N_22185,N_20695,N_20861);
nand U22186 (N_22186,N_21422,N_20782);
nand U22187 (N_22187,N_21015,N_21448);
nand U22188 (N_22188,N_20533,N_21344);
and U22189 (N_22189,N_21416,N_20508);
nand U22190 (N_22190,N_21290,N_20725);
or U22191 (N_22191,N_21130,N_21517);
nor U22192 (N_22192,N_21053,N_20717);
nand U22193 (N_22193,N_21502,N_21087);
xnor U22194 (N_22194,N_21527,N_21423);
and U22195 (N_22195,N_21534,N_20739);
or U22196 (N_22196,N_20688,N_20899);
xnor U22197 (N_22197,N_21490,N_20495);
nor U22198 (N_22198,N_20496,N_20848);
xor U22199 (N_22199,N_20511,N_20550);
nand U22200 (N_22200,N_21170,N_21243);
or U22201 (N_22201,N_21222,N_21320);
xnor U22202 (N_22202,N_20405,N_20525);
nor U22203 (N_22203,N_21575,N_20949);
or U22204 (N_22204,N_20916,N_20586);
or U22205 (N_22205,N_21321,N_21232);
nand U22206 (N_22206,N_20489,N_20732);
nand U22207 (N_22207,N_20689,N_21170);
nand U22208 (N_22208,N_21369,N_20713);
or U22209 (N_22209,N_21211,N_20486);
or U22210 (N_22210,N_21555,N_20920);
and U22211 (N_22211,N_20626,N_21507);
and U22212 (N_22212,N_20648,N_20543);
xor U22213 (N_22213,N_21158,N_20538);
and U22214 (N_22214,N_20947,N_21098);
and U22215 (N_22215,N_20998,N_20957);
nor U22216 (N_22216,N_21287,N_21544);
nor U22217 (N_22217,N_20562,N_21009);
and U22218 (N_22218,N_20476,N_20450);
nor U22219 (N_22219,N_21268,N_21066);
xnor U22220 (N_22220,N_20485,N_21573);
xor U22221 (N_22221,N_21373,N_20639);
and U22222 (N_22222,N_20822,N_21524);
nor U22223 (N_22223,N_21325,N_20890);
xnor U22224 (N_22224,N_20700,N_21264);
or U22225 (N_22225,N_21332,N_21098);
nor U22226 (N_22226,N_21311,N_20891);
or U22227 (N_22227,N_21283,N_20476);
and U22228 (N_22228,N_20896,N_21556);
xor U22229 (N_22229,N_21399,N_21473);
xnor U22230 (N_22230,N_20477,N_20910);
xor U22231 (N_22231,N_20847,N_20645);
xor U22232 (N_22232,N_21334,N_21549);
nand U22233 (N_22233,N_20564,N_21403);
nor U22234 (N_22234,N_21041,N_20584);
nor U22235 (N_22235,N_21417,N_20782);
xnor U22236 (N_22236,N_20887,N_20687);
xor U22237 (N_22237,N_20539,N_20749);
or U22238 (N_22238,N_20788,N_20862);
nand U22239 (N_22239,N_21198,N_20515);
and U22240 (N_22240,N_20918,N_21106);
or U22241 (N_22241,N_21153,N_20620);
nand U22242 (N_22242,N_21114,N_20774);
and U22243 (N_22243,N_21575,N_20458);
nand U22244 (N_22244,N_20790,N_20479);
xor U22245 (N_22245,N_20905,N_21398);
nor U22246 (N_22246,N_21258,N_20744);
or U22247 (N_22247,N_21260,N_20898);
nand U22248 (N_22248,N_20969,N_20800);
and U22249 (N_22249,N_20615,N_20603);
nand U22250 (N_22250,N_20504,N_21056);
and U22251 (N_22251,N_21354,N_20401);
xor U22252 (N_22252,N_20961,N_20979);
xnor U22253 (N_22253,N_21370,N_21128);
nor U22254 (N_22254,N_20881,N_21012);
nand U22255 (N_22255,N_20663,N_21151);
xnor U22256 (N_22256,N_21141,N_20686);
and U22257 (N_22257,N_20638,N_20976);
nand U22258 (N_22258,N_21440,N_20413);
and U22259 (N_22259,N_20553,N_20997);
nor U22260 (N_22260,N_21511,N_20849);
xnor U22261 (N_22261,N_20573,N_21231);
nand U22262 (N_22262,N_20630,N_21348);
and U22263 (N_22263,N_21446,N_20550);
or U22264 (N_22264,N_20437,N_20725);
nor U22265 (N_22265,N_21445,N_21042);
nand U22266 (N_22266,N_21479,N_21037);
and U22267 (N_22267,N_21538,N_21055);
nand U22268 (N_22268,N_20805,N_21403);
and U22269 (N_22269,N_20404,N_21163);
or U22270 (N_22270,N_21209,N_21472);
nor U22271 (N_22271,N_21135,N_20689);
and U22272 (N_22272,N_20621,N_21130);
nor U22273 (N_22273,N_20758,N_20461);
and U22274 (N_22274,N_20987,N_21543);
nor U22275 (N_22275,N_20423,N_21223);
nand U22276 (N_22276,N_21385,N_20543);
or U22277 (N_22277,N_21207,N_21325);
or U22278 (N_22278,N_20667,N_21477);
xor U22279 (N_22279,N_21431,N_21010);
and U22280 (N_22280,N_20685,N_20997);
nor U22281 (N_22281,N_21007,N_20680);
xnor U22282 (N_22282,N_20884,N_21287);
and U22283 (N_22283,N_21470,N_21364);
nor U22284 (N_22284,N_21476,N_21154);
nor U22285 (N_22285,N_21488,N_20813);
or U22286 (N_22286,N_21127,N_21412);
and U22287 (N_22287,N_20749,N_20738);
nand U22288 (N_22288,N_21540,N_21283);
nor U22289 (N_22289,N_21062,N_21130);
or U22290 (N_22290,N_20825,N_21223);
nand U22291 (N_22291,N_21194,N_20694);
nor U22292 (N_22292,N_20473,N_20727);
nand U22293 (N_22293,N_21273,N_21196);
xor U22294 (N_22294,N_20767,N_21465);
nand U22295 (N_22295,N_20463,N_21551);
nor U22296 (N_22296,N_21257,N_21581);
xnor U22297 (N_22297,N_21219,N_21056);
nand U22298 (N_22298,N_20941,N_20578);
nor U22299 (N_22299,N_20993,N_20509);
nand U22300 (N_22300,N_21289,N_20985);
nand U22301 (N_22301,N_20448,N_20925);
nor U22302 (N_22302,N_21037,N_20662);
or U22303 (N_22303,N_20785,N_21491);
or U22304 (N_22304,N_20980,N_21586);
and U22305 (N_22305,N_20542,N_21536);
nand U22306 (N_22306,N_20744,N_21080);
nand U22307 (N_22307,N_20727,N_20952);
and U22308 (N_22308,N_20631,N_21506);
xnor U22309 (N_22309,N_20722,N_21492);
nor U22310 (N_22310,N_21064,N_21253);
and U22311 (N_22311,N_20787,N_20495);
xnor U22312 (N_22312,N_21247,N_20477);
and U22313 (N_22313,N_20561,N_20933);
xor U22314 (N_22314,N_20947,N_20584);
and U22315 (N_22315,N_20924,N_21342);
nor U22316 (N_22316,N_21050,N_20434);
nor U22317 (N_22317,N_21014,N_21224);
nand U22318 (N_22318,N_21002,N_20963);
nor U22319 (N_22319,N_21138,N_20490);
or U22320 (N_22320,N_20883,N_20725);
and U22321 (N_22321,N_20656,N_20829);
nand U22322 (N_22322,N_20517,N_21098);
or U22323 (N_22323,N_20953,N_21019);
xor U22324 (N_22324,N_21150,N_21349);
or U22325 (N_22325,N_21430,N_20423);
nand U22326 (N_22326,N_21504,N_20918);
or U22327 (N_22327,N_21289,N_20803);
or U22328 (N_22328,N_20959,N_21198);
nand U22329 (N_22329,N_20790,N_20591);
and U22330 (N_22330,N_20904,N_20676);
and U22331 (N_22331,N_20943,N_21493);
xor U22332 (N_22332,N_20898,N_20779);
nor U22333 (N_22333,N_21513,N_20679);
and U22334 (N_22334,N_21304,N_21017);
and U22335 (N_22335,N_20820,N_20655);
xor U22336 (N_22336,N_20772,N_20982);
nand U22337 (N_22337,N_21018,N_21408);
xor U22338 (N_22338,N_20540,N_20997);
nand U22339 (N_22339,N_21112,N_20988);
and U22340 (N_22340,N_21091,N_20933);
or U22341 (N_22341,N_20818,N_21386);
or U22342 (N_22342,N_21239,N_20849);
xor U22343 (N_22343,N_20942,N_21367);
or U22344 (N_22344,N_21495,N_20535);
nand U22345 (N_22345,N_21444,N_20529);
and U22346 (N_22346,N_21178,N_20549);
nor U22347 (N_22347,N_20981,N_20817);
or U22348 (N_22348,N_20518,N_20490);
xor U22349 (N_22349,N_20450,N_21334);
nand U22350 (N_22350,N_21404,N_21066);
and U22351 (N_22351,N_21468,N_21545);
xnor U22352 (N_22352,N_20483,N_20574);
and U22353 (N_22353,N_20602,N_20505);
nand U22354 (N_22354,N_20837,N_21122);
nand U22355 (N_22355,N_20903,N_20712);
xnor U22356 (N_22356,N_20847,N_20953);
nand U22357 (N_22357,N_20951,N_20541);
nor U22358 (N_22358,N_20425,N_21551);
or U22359 (N_22359,N_20477,N_20458);
and U22360 (N_22360,N_21379,N_20611);
nand U22361 (N_22361,N_20818,N_20957);
or U22362 (N_22362,N_21333,N_20569);
nor U22363 (N_22363,N_21349,N_20986);
xnor U22364 (N_22364,N_20833,N_21265);
nor U22365 (N_22365,N_20486,N_21203);
xnor U22366 (N_22366,N_20564,N_21008);
nand U22367 (N_22367,N_21513,N_20560);
xor U22368 (N_22368,N_21482,N_20823);
nand U22369 (N_22369,N_20487,N_21384);
xor U22370 (N_22370,N_20686,N_20862);
nor U22371 (N_22371,N_20694,N_21362);
nand U22372 (N_22372,N_21077,N_20569);
or U22373 (N_22373,N_21449,N_21357);
and U22374 (N_22374,N_20611,N_21385);
nor U22375 (N_22375,N_21389,N_21283);
nor U22376 (N_22376,N_21599,N_20906);
and U22377 (N_22377,N_21344,N_20891);
xor U22378 (N_22378,N_20721,N_21481);
nand U22379 (N_22379,N_21518,N_20592);
xnor U22380 (N_22380,N_21445,N_20616);
xnor U22381 (N_22381,N_21345,N_20850);
and U22382 (N_22382,N_21420,N_21466);
or U22383 (N_22383,N_21586,N_21518);
xnor U22384 (N_22384,N_21304,N_21424);
nor U22385 (N_22385,N_20465,N_21494);
or U22386 (N_22386,N_21065,N_20794);
and U22387 (N_22387,N_20515,N_21320);
nor U22388 (N_22388,N_21254,N_20540);
nand U22389 (N_22389,N_21498,N_20961);
nand U22390 (N_22390,N_21334,N_21064);
and U22391 (N_22391,N_21540,N_20795);
or U22392 (N_22392,N_20540,N_21431);
nor U22393 (N_22393,N_20953,N_21400);
xor U22394 (N_22394,N_21259,N_20736);
or U22395 (N_22395,N_20409,N_21556);
nand U22396 (N_22396,N_20597,N_20909);
xor U22397 (N_22397,N_21173,N_20461);
and U22398 (N_22398,N_20946,N_20811);
or U22399 (N_22399,N_20871,N_20448);
nor U22400 (N_22400,N_20840,N_21374);
or U22401 (N_22401,N_20975,N_20544);
and U22402 (N_22402,N_20497,N_20771);
xnor U22403 (N_22403,N_21392,N_21247);
and U22404 (N_22404,N_20980,N_20400);
xnor U22405 (N_22405,N_20573,N_20863);
xnor U22406 (N_22406,N_21146,N_21599);
nand U22407 (N_22407,N_20885,N_20986);
nand U22408 (N_22408,N_21585,N_21113);
nand U22409 (N_22409,N_21459,N_20566);
xor U22410 (N_22410,N_20989,N_21045);
and U22411 (N_22411,N_21007,N_21338);
xor U22412 (N_22412,N_21083,N_21107);
nor U22413 (N_22413,N_21014,N_20548);
nand U22414 (N_22414,N_21570,N_21262);
nor U22415 (N_22415,N_21167,N_21220);
and U22416 (N_22416,N_21451,N_20989);
and U22417 (N_22417,N_20732,N_21194);
nand U22418 (N_22418,N_20659,N_20576);
and U22419 (N_22419,N_20890,N_20571);
or U22420 (N_22420,N_21050,N_21352);
xor U22421 (N_22421,N_21493,N_21511);
or U22422 (N_22422,N_20567,N_20518);
and U22423 (N_22423,N_20783,N_21290);
xor U22424 (N_22424,N_21317,N_21467);
or U22425 (N_22425,N_20734,N_21053);
or U22426 (N_22426,N_21294,N_20922);
nor U22427 (N_22427,N_21284,N_21292);
nand U22428 (N_22428,N_21359,N_20973);
xnor U22429 (N_22429,N_20993,N_20571);
nand U22430 (N_22430,N_21288,N_21399);
xnor U22431 (N_22431,N_21269,N_21042);
nor U22432 (N_22432,N_20864,N_20525);
or U22433 (N_22433,N_21253,N_21320);
nor U22434 (N_22434,N_20690,N_21160);
nand U22435 (N_22435,N_21312,N_20801);
nand U22436 (N_22436,N_20411,N_21542);
nor U22437 (N_22437,N_21403,N_21267);
and U22438 (N_22438,N_21007,N_20879);
and U22439 (N_22439,N_21177,N_20931);
nor U22440 (N_22440,N_21441,N_20481);
nor U22441 (N_22441,N_20735,N_20689);
nand U22442 (N_22442,N_20822,N_20524);
and U22443 (N_22443,N_20488,N_21305);
xor U22444 (N_22444,N_21177,N_20501);
nor U22445 (N_22445,N_20884,N_20594);
xor U22446 (N_22446,N_20665,N_20768);
and U22447 (N_22447,N_20537,N_21217);
or U22448 (N_22448,N_20985,N_20652);
or U22449 (N_22449,N_21059,N_20430);
or U22450 (N_22450,N_21179,N_21375);
xor U22451 (N_22451,N_20774,N_20466);
nor U22452 (N_22452,N_20870,N_21234);
nor U22453 (N_22453,N_20962,N_21433);
xnor U22454 (N_22454,N_20627,N_21399);
or U22455 (N_22455,N_21118,N_21014);
and U22456 (N_22456,N_21487,N_20762);
and U22457 (N_22457,N_21155,N_21216);
or U22458 (N_22458,N_20801,N_20683);
or U22459 (N_22459,N_20766,N_20983);
and U22460 (N_22460,N_21445,N_20505);
xor U22461 (N_22461,N_20948,N_20994);
or U22462 (N_22462,N_21027,N_20772);
nand U22463 (N_22463,N_21289,N_21355);
nand U22464 (N_22464,N_21537,N_20966);
nor U22465 (N_22465,N_21252,N_21352);
or U22466 (N_22466,N_21074,N_21425);
or U22467 (N_22467,N_20680,N_21038);
and U22468 (N_22468,N_20860,N_20698);
and U22469 (N_22469,N_21133,N_21231);
nand U22470 (N_22470,N_20700,N_21326);
nand U22471 (N_22471,N_20771,N_20756);
nand U22472 (N_22472,N_20501,N_20967);
or U22473 (N_22473,N_20436,N_20885);
and U22474 (N_22474,N_20481,N_20539);
nand U22475 (N_22475,N_20740,N_20670);
xor U22476 (N_22476,N_20882,N_20895);
xnor U22477 (N_22477,N_20760,N_21450);
nor U22478 (N_22478,N_21449,N_20521);
nand U22479 (N_22479,N_20553,N_21511);
nand U22480 (N_22480,N_20967,N_20887);
and U22481 (N_22481,N_21242,N_20576);
nor U22482 (N_22482,N_21089,N_21415);
xnor U22483 (N_22483,N_20805,N_20903);
nand U22484 (N_22484,N_21271,N_21168);
nand U22485 (N_22485,N_20684,N_20822);
nor U22486 (N_22486,N_20754,N_20599);
nand U22487 (N_22487,N_20784,N_20480);
and U22488 (N_22488,N_20470,N_20433);
and U22489 (N_22489,N_21205,N_21322);
xnor U22490 (N_22490,N_21087,N_20874);
nor U22491 (N_22491,N_20506,N_21381);
xor U22492 (N_22492,N_21182,N_21396);
nand U22493 (N_22493,N_21423,N_20470);
or U22494 (N_22494,N_20841,N_21010);
xor U22495 (N_22495,N_20728,N_21269);
or U22496 (N_22496,N_20880,N_21278);
nor U22497 (N_22497,N_20407,N_21278);
and U22498 (N_22498,N_21340,N_21058);
nand U22499 (N_22499,N_20751,N_21311);
xnor U22500 (N_22500,N_20538,N_20737);
xnor U22501 (N_22501,N_21556,N_21083);
or U22502 (N_22502,N_21286,N_21568);
nor U22503 (N_22503,N_21163,N_20436);
xor U22504 (N_22504,N_21065,N_20432);
nor U22505 (N_22505,N_20874,N_20855);
and U22506 (N_22506,N_20797,N_20820);
xnor U22507 (N_22507,N_21481,N_20514);
xnor U22508 (N_22508,N_21103,N_20807);
nand U22509 (N_22509,N_21594,N_20651);
and U22510 (N_22510,N_21112,N_20767);
nor U22511 (N_22511,N_20440,N_21003);
and U22512 (N_22512,N_20586,N_21127);
and U22513 (N_22513,N_21125,N_20701);
nand U22514 (N_22514,N_21597,N_20702);
or U22515 (N_22515,N_21522,N_20545);
and U22516 (N_22516,N_20446,N_21598);
and U22517 (N_22517,N_21528,N_21030);
xor U22518 (N_22518,N_21580,N_20419);
nand U22519 (N_22519,N_21030,N_21266);
xnor U22520 (N_22520,N_20430,N_21262);
and U22521 (N_22521,N_20605,N_21308);
nand U22522 (N_22522,N_20486,N_20909);
xor U22523 (N_22523,N_20488,N_21115);
nand U22524 (N_22524,N_21418,N_20798);
xor U22525 (N_22525,N_20956,N_20950);
nand U22526 (N_22526,N_20946,N_21047);
nor U22527 (N_22527,N_20634,N_20712);
nor U22528 (N_22528,N_21574,N_21188);
nor U22529 (N_22529,N_21079,N_20486);
xor U22530 (N_22530,N_21417,N_21438);
nor U22531 (N_22531,N_21371,N_20404);
and U22532 (N_22532,N_20529,N_20488);
xnor U22533 (N_22533,N_20908,N_20438);
or U22534 (N_22534,N_20472,N_21429);
xor U22535 (N_22535,N_21301,N_20913);
and U22536 (N_22536,N_20641,N_20670);
nor U22537 (N_22537,N_20555,N_20682);
xnor U22538 (N_22538,N_21044,N_21400);
xnor U22539 (N_22539,N_20883,N_21262);
nor U22540 (N_22540,N_21083,N_21088);
nor U22541 (N_22541,N_21010,N_20660);
or U22542 (N_22542,N_21559,N_20585);
or U22543 (N_22543,N_20806,N_21114);
or U22544 (N_22544,N_20883,N_21400);
nor U22545 (N_22545,N_21053,N_21397);
and U22546 (N_22546,N_21490,N_20408);
or U22547 (N_22547,N_21514,N_20899);
and U22548 (N_22548,N_20961,N_20468);
xnor U22549 (N_22549,N_20864,N_20579);
nor U22550 (N_22550,N_20940,N_21033);
and U22551 (N_22551,N_20816,N_20517);
or U22552 (N_22552,N_21314,N_21421);
and U22553 (N_22553,N_21341,N_20415);
or U22554 (N_22554,N_20697,N_20430);
nand U22555 (N_22555,N_20861,N_21182);
or U22556 (N_22556,N_21569,N_21528);
xor U22557 (N_22557,N_20516,N_20410);
and U22558 (N_22558,N_21236,N_20736);
and U22559 (N_22559,N_21125,N_21582);
nor U22560 (N_22560,N_21075,N_21003);
xnor U22561 (N_22561,N_20857,N_20981);
or U22562 (N_22562,N_21507,N_21339);
xor U22563 (N_22563,N_20737,N_20460);
nand U22564 (N_22564,N_21541,N_20542);
nand U22565 (N_22565,N_21285,N_20729);
xor U22566 (N_22566,N_20771,N_20846);
xnor U22567 (N_22567,N_20903,N_20708);
nand U22568 (N_22568,N_21147,N_20680);
nor U22569 (N_22569,N_21051,N_20763);
or U22570 (N_22570,N_20588,N_20503);
or U22571 (N_22571,N_20784,N_20921);
nand U22572 (N_22572,N_21097,N_20512);
or U22573 (N_22573,N_20455,N_20664);
and U22574 (N_22574,N_21139,N_20729);
xor U22575 (N_22575,N_21163,N_21304);
or U22576 (N_22576,N_21416,N_20525);
xor U22577 (N_22577,N_21374,N_20918);
nor U22578 (N_22578,N_20472,N_20632);
or U22579 (N_22579,N_21165,N_21218);
or U22580 (N_22580,N_20997,N_21478);
nand U22581 (N_22581,N_21084,N_20858);
nand U22582 (N_22582,N_21492,N_20583);
nand U22583 (N_22583,N_21358,N_21372);
or U22584 (N_22584,N_21552,N_20529);
or U22585 (N_22585,N_20923,N_20907);
and U22586 (N_22586,N_21313,N_21097);
xor U22587 (N_22587,N_21456,N_20932);
nor U22588 (N_22588,N_21461,N_21499);
xor U22589 (N_22589,N_21565,N_20954);
xnor U22590 (N_22590,N_21209,N_20892);
and U22591 (N_22591,N_21127,N_20687);
nor U22592 (N_22592,N_21377,N_20868);
xnor U22593 (N_22593,N_20563,N_21424);
nor U22594 (N_22594,N_21457,N_20484);
or U22595 (N_22595,N_20779,N_20514);
and U22596 (N_22596,N_20500,N_20807);
or U22597 (N_22597,N_20666,N_21372);
nor U22598 (N_22598,N_21127,N_21577);
and U22599 (N_22599,N_20801,N_20823);
and U22600 (N_22600,N_20965,N_20826);
and U22601 (N_22601,N_21184,N_21358);
or U22602 (N_22602,N_21243,N_21180);
xor U22603 (N_22603,N_21375,N_21193);
or U22604 (N_22604,N_20554,N_21341);
or U22605 (N_22605,N_21305,N_21177);
or U22606 (N_22606,N_21597,N_20761);
xnor U22607 (N_22607,N_21286,N_20668);
nand U22608 (N_22608,N_21509,N_21529);
and U22609 (N_22609,N_21305,N_20543);
nor U22610 (N_22610,N_21544,N_20978);
xnor U22611 (N_22611,N_21261,N_20817);
nor U22612 (N_22612,N_21085,N_21361);
and U22613 (N_22613,N_20857,N_20575);
xor U22614 (N_22614,N_20529,N_20725);
and U22615 (N_22615,N_21518,N_21119);
or U22616 (N_22616,N_20438,N_21091);
and U22617 (N_22617,N_20934,N_20806);
nand U22618 (N_22618,N_21568,N_21562);
nor U22619 (N_22619,N_21210,N_20491);
nand U22620 (N_22620,N_21232,N_20493);
xnor U22621 (N_22621,N_20471,N_20819);
nand U22622 (N_22622,N_20536,N_20954);
nand U22623 (N_22623,N_20932,N_20788);
xor U22624 (N_22624,N_21273,N_21051);
nand U22625 (N_22625,N_21585,N_21328);
xnor U22626 (N_22626,N_21356,N_20927);
and U22627 (N_22627,N_20444,N_20711);
and U22628 (N_22628,N_21315,N_21246);
nand U22629 (N_22629,N_21460,N_20873);
and U22630 (N_22630,N_20971,N_20789);
and U22631 (N_22631,N_21254,N_20940);
nor U22632 (N_22632,N_20983,N_21537);
or U22633 (N_22633,N_21138,N_20466);
nor U22634 (N_22634,N_20479,N_21547);
nor U22635 (N_22635,N_21434,N_20547);
nand U22636 (N_22636,N_20646,N_20533);
nor U22637 (N_22637,N_21524,N_21219);
and U22638 (N_22638,N_21269,N_21363);
and U22639 (N_22639,N_21465,N_21238);
or U22640 (N_22640,N_20699,N_21161);
nand U22641 (N_22641,N_21159,N_21230);
and U22642 (N_22642,N_21494,N_21304);
xor U22643 (N_22643,N_20601,N_20589);
or U22644 (N_22644,N_21548,N_20648);
and U22645 (N_22645,N_21178,N_21208);
xor U22646 (N_22646,N_20581,N_20910);
nand U22647 (N_22647,N_21547,N_20674);
or U22648 (N_22648,N_21164,N_21214);
nand U22649 (N_22649,N_21349,N_20603);
nor U22650 (N_22650,N_21166,N_21371);
or U22651 (N_22651,N_20459,N_21334);
and U22652 (N_22652,N_20544,N_21151);
xor U22653 (N_22653,N_20602,N_21169);
and U22654 (N_22654,N_21483,N_21312);
or U22655 (N_22655,N_21555,N_20726);
nand U22656 (N_22656,N_21468,N_20576);
xor U22657 (N_22657,N_21504,N_21577);
xor U22658 (N_22658,N_21207,N_21304);
and U22659 (N_22659,N_21471,N_20850);
nand U22660 (N_22660,N_21422,N_20931);
nand U22661 (N_22661,N_21432,N_20761);
nand U22662 (N_22662,N_20880,N_20956);
nand U22663 (N_22663,N_21112,N_20801);
or U22664 (N_22664,N_21349,N_20717);
and U22665 (N_22665,N_20859,N_20784);
and U22666 (N_22666,N_21144,N_21530);
and U22667 (N_22667,N_20764,N_20867);
or U22668 (N_22668,N_20799,N_21274);
nand U22669 (N_22669,N_21042,N_21355);
nand U22670 (N_22670,N_20991,N_20413);
xnor U22671 (N_22671,N_20891,N_20508);
nand U22672 (N_22672,N_21297,N_20411);
and U22673 (N_22673,N_21228,N_21566);
and U22674 (N_22674,N_21338,N_21495);
nor U22675 (N_22675,N_20969,N_20540);
nor U22676 (N_22676,N_20814,N_20479);
nor U22677 (N_22677,N_21423,N_21169);
or U22678 (N_22678,N_20605,N_20684);
nor U22679 (N_22679,N_21245,N_21215);
xnor U22680 (N_22680,N_20921,N_21094);
nor U22681 (N_22681,N_21139,N_21264);
or U22682 (N_22682,N_21577,N_21227);
nor U22683 (N_22683,N_21446,N_21089);
or U22684 (N_22684,N_20419,N_21071);
nand U22685 (N_22685,N_21393,N_21361);
and U22686 (N_22686,N_20536,N_20433);
xnor U22687 (N_22687,N_20523,N_20533);
or U22688 (N_22688,N_21323,N_20435);
xnor U22689 (N_22689,N_21367,N_21035);
or U22690 (N_22690,N_20523,N_21232);
nor U22691 (N_22691,N_21574,N_21237);
nand U22692 (N_22692,N_21129,N_20969);
xor U22693 (N_22693,N_21250,N_21325);
nand U22694 (N_22694,N_21407,N_20641);
xor U22695 (N_22695,N_21356,N_20920);
nand U22696 (N_22696,N_20826,N_21453);
nor U22697 (N_22697,N_21272,N_20436);
nor U22698 (N_22698,N_21190,N_21415);
nand U22699 (N_22699,N_21042,N_20903);
nand U22700 (N_22700,N_21556,N_20841);
nor U22701 (N_22701,N_20790,N_20548);
xnor U22702 (N_22702,N_21270,N_21010);
nor U22703 (N_22703,N_20718,N_21131);
and U22704 (N_22704,N_20726,N_21453);
or U22705 (N_22705,N_21569,N_21545);
nor U22706 (N_22706,N_20674,N_21311);
and U22707 (N_22707,N_21452,N_20861);
nand U22708 (N_22708,N_20544,N_20420);
nor U22709 (N_22709,N_21149,N_21581);
xnor U22710 (N_22710,N_20475,N_21060);
xnor U22711 (N_22711,N_21570,N_21010);
or U22712 (N_22712,N_20621,N_21471);
nor U22713 (N_22713,N_20583,N_21518);
or U22714 (N_22714,N_21455,N_21463);
nand U22715 (N_22715,N_20912,N_21289);
xor U22716 (N_22716,N_21313,N_20769);
and U22717 (N_22717,N_20796,N_20932);
and U22718 (N_22718,N_21433,N_20506);
nor U22719 (N_22719,N_21445,N_20838);
nand U22720 (N_22720,N_21255,N_21034);
and U22721 (N_22721,N_20662,N_20445);
and U22722 (N_22722,N_21484,N_21340);
nand U22723 (N_22723,N_20428,N_20540);
or U22724 (N_22724,N_20822,N_21005);
nand U22725 (N_22725,N_21263,N_21531);
xnor U22726 (N_22726,N_20724,N_21327);
nand U22727 (N_22727,N_21573,N_21141);
nor U22728 (N_22728,N_20636,N_21396);
or U22729 (N_22729,N_21298,N_21369);
and U22730 (N_22730,N_20747,N_20993);
xnor U22731 (N_22731,N_20893,N_20976);
nor U22732 (N_22732,N_20653,N_20827);
nor U22733 (N_22733,N_20765,N_20792);
or U22734 (N_22734,N_20581,N_20525);
nand U22735 (N_22735,N_20580,N_20706);
xor U22736 (N_22736,N_20976,N_20405);
or U22737 (N_22737,N_21392,N_21114);
nand U22738 (N_22738,N_20999,N_21490);
or U22739 (N_22739,N_21526,N_21238);
nand U22740 (N_22740,N_20684,N_21243);
and U22741 (N_22741,N_21307,N_21191);
and U22742 (N_22742,N_20928,N_21347);
or U22743 (N_22743,N_20986,N_20487);
nand U22744 (N_22744,N_21459,N_21589);
xnor U22745 (N_22745,N_20981,N_21065);
nand U22746 (N_22746,N_20764,N_21306);
nor U22747 (N_22747,N_20757,N_21070);
nand U22748 (N_22748,N_20930,N_21063);
nor U22749 (N_22749,N_21419,N_20870);
nor U22750 (N_22750,N_20963,N_20740);
xor U22751 (N_22751,N_20742,N_20591);
or U22752 (N_22752,N_20724,N_20674);
or U22753 (N_22753,N_21494,N_21534);
xor U22754 (N_22754,N_20549,N_21012);
xor U22755 (N_22755,N_21062,N_21077);
nor U22756 (N_22756,N_21482,N_21295);
xor U22757 (N_22757,N_21503,N_20636);
or U22758 (N_22758,N_21018,N_21258);
nor U22759 (N_22759,N_21481,N_21586);
and U22760 (N_22760,N_20974,N_21091);
and U22761 (N_22761,N_20987,N_21459);
and U22762 (N_22762,N_21053,N_20970);
nor U22763 (N_22763,N_20987,N_20731);
nor U22764 (N_22764,N_21258,N_21576);
and U22765 (N_22765,N_21270,N_20599);
or U22766 (N_22766,N_21013,N_20456);
and U22767 (N_22767,N_21284,N_20865);
xor U22768 (N_22768,N_21256,N_20563);
or U22769 (N_22769,N_20954,N_21057);
xor U22770 (N_22770,N_20474,N_20936);
nor U22771 (N_22771,N_20530,N_21589);
xnor U22772 (N_22772,N_21337,N_20588);
and U22773 (N_22773,N_20497,N_20438);
and U22774 (N_22774,N_21466,N_20641);
nor U22775 (N_22775,N_21325,N_20665);
or U22776 (N_22776,N_21147,N_21314);
nor U22777 (N_22777,N_20435,N_21228);
xor U22778 (N_22778,N_20820,N_20534);
nor U22779 (N_22779,N_20845,N_20806);
xnor U22780 (N_22780,N_20920,N_20965);
or U22781 (N_22781,N_20645,N_20710);
xnor U22782 (N_22782,N_21066,N_20965);
nand U22783 (N_22783,N_21333,N_20660);
xnor U22784 (N_22784,N_20537,N_20809);
xor U22785 (N_22785,N_21471,N_21175);
or U22786 (N_22786,N_20753,N_20877);
xnor U22787 (N_22787,N_20703,N_20758);
or U22788 (N_22788,N_20571,N_21213);
nand U22789 (N_22789,N_21569,N_20872);
and U22790 (N_22790,N_20466,N_21353);
nand U22791 (N_22791,N_21177,N_21514);
nand U22792 (N_22792,N_20760,N_21555);
xnor U22793 (N_22793,N_21042,N_20621);
or U22794 (N_22794,N_21528,N_20778);
nor U22795 (N_22795,N_20769,N_20540);
and U22796 (N_22796,N_21218,N_20713);
nand U22797 (N_22797,N_20980,N_21391);
nand U22798 (N_22798,N_21254,N_20651);
or U22799 (N_22799,N_21554,N_21363);
xor U22800 (N_22800,N_22145,N_22006);
and U22801 (N_22801,N_21642,N_22666);
xnor U22802 (N_22802,N_21719,N_22517);
xor U22803 (N_22803,N_22080,N_22622);
xor U22804 (N_22804,N_22166,N_22263);
nand U22805 (N_22805,N_22093,N_22001);
nand U22806 (N_22806,N_21757,N_22062);
nor U22807 (N_22807,N_21639,N_22060);
xor U22808 (N_22808,N_22641,N_22402);
or U22809 (N_22809,N_21792,N_21980);
nor U22810 (N_22810,N_22662,N_22432);
nor U22811 (N_22811,N_21838,N_22475);
and U22812 (N_22812,N_22204,N_22528);
or U22813 (N_22813,N_22621,N_22000);
or U22814 (N_22814,N_22683,N_21773);
and U22815 (N_22815,N_22125,N_21798);
nand U22816 (N_22816,N_22045,N_22678);
nor U22817 (N_22817,N_21795,N_22746);
nor U22818 (N_22818,N_21731,N_21820);
nand U22819 (N_22819,N_22680,N_21600);
nand U22820 (N_22820,N_21660,N_22293);
and U22821 (N_22821,N_22154,N_22282);
nor U22822 (N_22822,N_22525,N_22403);
and U22823 (N_22823,N_22146,N_22753);
or U22824 (N_22824,N_21834,N_22454);
and U22825 (N_22825,N_22655,N_21830);
nand U22826 (N_22826,N_22118,N_22371);
or U22827 (N_22827,N_22373,N_22259);
and U22828 (N_22828,N_21961,N_22257);
nor U22829 (N_22829,N_22554,N_22742);
and U22830 (N_22830,N_22094,N_21990);
xnor U22831 (N_22831,N_21770,N_22553);
or U22832 (N_22832,N_21790,N_21666);
nor U22833 (N_22833,N_21939,N_22791);
xor U22834 (N_22834,N_21669,N_21744);
xor U22835 (N_22835,N_22123,N_22012);
nor U22836 (N_22836,N_22441,N_22430);
nand U22837 (N_22837,N_21747,N_22550);
or U22838 (N_22838,N_21813,N_22053);
nor U22839 (N_22839,N_22215,N_22479);
nand U22840 (N_22840,N_22505,N_22458);
nand U22841 (N_22841,N_21614,N_22738);
or U22842 (N_22842,N_22075,N_21951);
and U22843 (N_22843,N_22609,N_22568);
nand U22844 (N_22844,N_21636,N_22198);
nor U22845 (N_22845,N_21877,N_22730);
xnor U22846 (N_22846,N_22321,N_21685);
nor U22847 (N_22847,N_21687,N_22179);
nor U22848 (N_22848,N_21756,N_22377);
xnor U22849 (N_22849,N_21616,N_21917);
nor U22850 (N_22850,N_21948,N_21721);
and U22851 (N_22851,N_21858,N_22063);
or U22852 (N_22852,N_22197,N_22460);
or U22853 (N_22853,N_22795,N_22133);
nand U22854 (N_22854,N_22563,N_21787);
or U22855 (N_22855,N_21649,N_22055);
and U22856 (N_22856,N_22391,N_22231);
xnor U22857 (N_22857,N_21698,N_22237);
nor U22858 (N_22858,N_22392,N_22346);
nor U22859 (N_22859,N_22155,N_22462);
or U22860 (N_22860,N_22589,N_21882);
xnor U22861 (N_22861,N_22591,N_22054);
xnor U22862 (N_22862,N_21899,N_21689);
or U22863 (N_22863,N_22124,N_22461);
xor U22864 (N_22864,N_22630,N_22511);
or U22865 (N_22865,N_22538,N_22775);
nor U22866 (N_22866,N_21761,N_22233);
or U22867 (N_22867,N_22411,N_22760);
nand U22868 (N_22868,N_22032,N_21849);
and U22869 (N_22869,N_21654,N_22141);
nand U22870 (N_22870,N_22797,N_21743);
nand U22871 (N_22871,N_21662,N_21690);
xnor U22872 (N_22872,N_21791,N_22018);
xor U22873 (N_22873,N_22472,N_22407);
or U22874 (N_22874,N_22670,N_22028);
nor U22875 (N_22875,N_22681,N_22169);
xnor U22876 (N_22876,N_21863,N_22184);
or U22877 (N_22877,N_22485,N_22449);
xor U22878 (N_22878,N_22529,N_22111);
or U22879 (N_22879,N_22225,N_22544);
nand U22880 (N_22880,N_21665,N_22576);
and U22881 (N_22881,N_22369,N_22116);
and U22882 (N_22882,N_22380,N_22719);
and U22883 (N_22883,N_22716,N_21755);
and U22884 (N_22884,N_21811,N_22552);
nand U22885 (N_22885,N_21776,N_21602);
or U22886 (N_22886,N_21752,N_22177);
xor U22887 (N_22887,N_22510,N_22439);
nor U22888 (N_22888,N_22273,N_22261);
nand U22889 (N_22889,N_22319,N_21793);
xnor U22890 (N_22890,N_21728,N_21851);
or U22891 (N_22891,N_21855,N_21641);
or U22892 (N_22892,N_22498,N_22624);
xor U22893 (N_22893,N_22309,N_22556);
or U22894 (N_22894,N_22634,N_22672);
nor U22895 (N_22895,N_22307,N_22252);
xnor U22896 (N_22896,N_22159,N_22256);
or U22897 (N_22897,N_22682,N_22691);
and U22898 (N_22898,N_22151,N_22561);
nor U22899 (N_22899,N_22639,N_22577);
nor U22900 (N_22900,N_21624,N_21722);
nor U22901 (N_22901,N_21700,N_22378);
nor U22902 (N_22902,N_22705,N_22564);
nor U22903 (N_22903,N_22372,N_22539);
nand U22904 (N_22904,N_22438,N_22569);
nor U22905 (N_22905,N_22776,N_22696);
nand U22906 (N_22906,N_22777,N_21983);
xor U22907 (N_22907,N_21869,N_22183);
and U22908 (N_22908,N_22469,N_22192);
xnor U22909 (N_22909,N_22444,N_22101);
xor U22910 (N_22910,N_21883,N_21868);
nand U22911 (N_22911,N_22203,N_22542);
nor U22912 (N_22912,N_22779,N_21936);
xnor U22913 (N_22913,N_22036,N_22326);
or U22914 (N_22914,N_21764,N_22484);
nand U22915 (N_22915,N_21908,N_22153);
nor U22916 (N_22916,N_22697,N_21736);
nand U22917 (N_22917,N_21769,N_21780);
or U22918 (N_22918,N_22205,N_22115);
nand U22919 (N_22919,N_22656,N_22686);
nor U22920 (N_22920,N_22074,N_22463);
nand U22921 (N_22921,N_22446,N_21796);
xor U22922 (N_22922,N_22174,N_22781);
or U22923 (N_22923,N_22489,N_22370);
and U22924 (N_22924,N_22052,N_21784);
nand U22925 (N_22925,N_21766,N_22745);
or U22926 (N_22926,N_21625,N_21872);
nand U22927 (N_22927,N_21867,N_21896);
or U22928 (N_22928,N_22114,N_22186);
nand U22929 (N_22929,N_22787,N_22758);
and U22930 (N_22930,N_22132,N_21930);
nand U22931 (N_22931,N_21652,N_22314);
nor U22932 (N_22932,N_22566,N_22305);
xnor U22933 (N_22933,N_22456,N_22037);
nand U22934 (N_22934,N_22384,N_22281);
nor U22935 (N_22935,N_21841,N_22532);
or U22936 (N_22936,N_21901,N_21732);
xnor U22937 (N_22937,N_22021,N_22669);
and U22938 (N_22938,N_22612,N_22303);
nand U22939 (N_22939,N_21950,N_22158);
nand U22940 (N_22940,N_21812,N_22148);
xor U22941 (N_22941,N_22199,N_21783);
nand U22942 (N_22942,N_22535,N_22249);
and U22943 (N_22943,N_22718,N_22286);
and U22944 (N_22944,N_21692,N_22499);
nor U22945 (N_22945,N_21965,N_22332);
xor U22946 (N_22946,N_21847,N_22657);
or U22947 (N_22947,N_22279,N_22193);
or U22948 (N_22948,N_21828,N_22424);
or U22949 (N_22949,N_22418,N_22503);
nor U22950 (N_22950,N_22262,N_22011);
and U22951 (N_22951,N_22022,N_22120);
nor U22952 (N_22952,N_22619,N_22049);
and U22953 (N_22953,N_21920,N_22520);
nand U22954 (N_22954,N_22057,N_22731);
xnor U22955 (N_22955,N_22239,N_22690);
and U22956 (N_22956,N_22355,N_22200);
or U22957 (N_22957,N_21688,N_21745);
nor U22958 (N_22958,N_21762,N_22756);
or U22959 (N_22959,N_21767,N_22422);
nor U22960 (N_22960,N_22635,N_21891);
and U22961 (N_22961,N_21984,N_22616);
or U22962 (N_22962,N_22401,N_21964);
xnor U22963 (N_22963,N_22429,N_21737);
nand U22964 (N_22964,N_21630,N_22008);
xnor U22965 (N_22965,N_22390,N_22724);
nor U22966 (N_22966,N_22064,N_21749);
and U22967 (N_22967,N_22389,N_22220);
and U22968 (N_22968,N_21963,N_21754);
xor U22969 (N_22969,N_21680,N_22222);
and U22970 (N_22970,N_21782,N_22216);
nand U22971 (N_22971,N_22692,N_21724);
or U22972 (N_22972,N_22598,N_22398);
nand U22973 (N_22973,N_22768,N_22604);
nor U22974 (N_22974,N_22406,N_22350);
nor U22975 (N_22975,N_22091,N_22530);
nor U22976 (N_22976,N_22014,N_21972);
nand U22977 (N_22977,N_22409,N_22653);
nor U22978 (N_22978,N_22702,N_22477);
xnor U22979 (N_22979,N_21935,N_22786);
nor U22980 (N_22980,N_22487,N_22104);
xor U22981 (N_22981,N_21681,N_21938);
nand U22982 (N_22982,N_22291,N_22476);
nand U22983 (N_22983,N_22089,N_21873);
xor U22984 (N_22984,N_22707,N_21673);
nand U22985 (N_22985,N_21661,N_21871);
nand U22986 (N_22986,N_21985,N_21703);
xor U22987 (N_22987,N_22481,N_22752);
nand U22988 (N_22988,N_21907,N_22061);
nor U22989 (N_22989,N_22365,N_22796);
xor U22990 (N_22990,N_22574,N_21640);
xnor U22991 (N_22991,N_22443,N_22207);
or U22992 (N_22992,N_21620,N_22755);
and U22993 (N_22993,N_22726,N_22764);
nor U22994 (N_22994,N_21827,N_21678);
nand U22995 (N_22995,N_22783,N_21663);
nor U22996 (N_22996,N_22560,N_22241);
or U22997 (N_22997,N_22152,N_22329);
or U22998 (N_22998,N_22607,N_22181);
and U22999 (N_22999,N_22306,N_22296);
xor U23000 (N_23000,N_21991,N_21959);
nor U23001 (N_23001,N_21889,N_21768);
nor U23002 (N_23002,N_21894,N_22229);
and U23003 (N_23003,N_22570,N_22171);
xor U23004 (N_23004,N_21676,N_22349);
xor U23005 (N_23005,N_22005,N_22173);
xor U23006 (N_23006,N_22297,N_22397);
nor U23007 (N_23007,N_22142,N_22227);
and U23008 (N_23008,N_21606,N_22450);
xor U23009 (N_23009,N_21805,N_21941);
and U23010 (N_23010,N_22362,N_21904);
nand U23011 (N_23011,N_22357,N_21881);
or U23012 (N_23012,N_21840,N_22625);
nor U23013 (N_23013,N_21940,N_22260);
nand U23014 (N_23014,N_22295,N_22134);
xor U23015 (N_23015,N_22799,N_22209);
and U23016 (N_23016,N_22067,N_22234);
nand U23017 (N_23017,N_22368,N_22717);
and U23018 (N_23018,N_21800,N_22773);
nand U23019 (N_23019,N_22191,N_22493);
and U23020 (N_23020,N_22747,N_22351);
xnor U23021 (N_23021,N_22269,N_22533);
and U23022 (N_23022,N_22601,N_21954);
and U23023 (N_23023,N_22386,N_22046);
nor U23024 (N_23024,N_22405,N_22311);
nor U23025 (N_23025,N_22253,N_21746);
and U23026 (N_23026,N_22595,N_22770);
or U23027 (N_23027,N_22754,N_21926);
nand U23028 (N_23028,N_22650,N_22188);
and U23029 (N_23029,N_21903,N_22693);
and U23030 (N_23030,N_21897,N_21878);
and U23031 (N_23031,N_22587,N_21706);
and U23032 (N_23032,N_21704,N_22023);
nor U23033 (N_23033,N_22393,N_22341);
nor U23034 (N_23034,N_21699,N_22593);
and U23035 (N_23035,N_22292,N_21657);
nor U23036 (N_23036,N_22482,N_22108);
nor U23037 (N_23037,N_22739,N_22122);
and U23038 (N_23038,N_22050,N_21843);
or U23039 (N_23039,N_22255,N_22661);
and U23040 (N_23040,N_22626,N_22526);
xor U23041 (N_23041,N_22013,N_21802);
nor U23042 (N_23042,N_21694,N_21819);
nor U23043 (N_23043,N_22778,N_21741);
or U23044 (N_23044,N_21646,N_22496);
xor U23045 (N_23045,N_21603,N_22425);
and U23046 (N_23046,N_22644,N_22737);
nand U23047 (N_23047,N_21919,N_22506);
xor U23048 (N_23048,N_21982,N_22264);
xor U23049 (N_23049,N_21957,N_22009);
or U23050 (N_23050,N_22160,N_22504);
or U23051 (N_23051,N_22521,N_22043);
xor U23052 (N_23052,N_21804,N_21932);
nor U23053 (N_23053,N_22047,N_22268);
nand U23054 (N_23054,N_21845,N_22408);
nand U23055 (N_23055,N_22361,N_22290);
nand U23056 (N_23056,N_22694,N_22343);
nor U23057 (N_23057,N_21672,N_22792);
nor U23058 (N_23058,N_22614,N_21609);
nor U23059 (N_23059,N_22066,N_22344);
or U23060 (N_23060,N_22095,N_22038);
xnor U23061 (N_23061,N_21921,N_21727);
and U23062 (N_23062,N_22338,N_22789);
nor U23063 (N_23063,N_21627,N_22208);
or U23064 (N_23064,N_22794,N_22647);
nor U23065 (N_23065,N_22143,N_22761);
nor U23066 (N_23066,N_21997,N_21969);
and U23067 (N_23067,N_21635,N_21677);
nand U23068 (N_23068,N_22112,N_22762);
or U23069 (N_23069,N_21816,N_22410);
and U23070 (N_23070,N_21610,N_22494);
and U23071 (N_23071,N_22163,N_22790);
xnor U23072 (N_23072,N_22740,N_21684);
or U23073 (N_23073,N_22082,N_22618);
xnor U23074 (N_23074,N_22793,N_21993);
and U23075 (N_23075,N_22435,N_22218);
xor U23076 (N_23076,N_21848,N_21717);
nand U23077 (N_23077,N_21996,N_21623);
xor U23078 (N_23078,N_22715,N_22258);
nand U23079 (N_23079,N_22396,N_21695);
or U23080 (N_23080,N_21622,N_22774);
and U23081 (N_23081,N_22523,N_21708);
and U23082 (N_23082,N_22381,N_21975);
nor U23083 (N_23083,N_21825,N_22628);
or U23084 (N_23084,N_21826,N_22072);
nand U23085 (N_23085,N_21857,N_22376);
xor U23086 (N_23086,N_22562,N_22310);
xor U23087 (N_23087,N_22327,N_22097);
nand U23088 (N_23088,N_22785,N_22301);
xnor U23089 (N_23089,N_22394,N_22058);
or U23090 (N_23090,N_22375,N_22352);
xor U23091 (N_23091,N_22024,N_22027);
xor U23092 (N_23092,N_22335,N_22345);
xor U23093 (N_23093,N_21705,N_22323);
and U23094 (N_23094,N_22098,N_22507);
and U23095 (N_23095,N_22480,N_21810);
xor U23096 (N_23096,N_22664,N_21852);
xnor U23097 (N_23097,N_22748,N_22202);
xnor U23098 (N_23098,N_22266,N_21906);
and U23099 (N_23099,N_21905,N_22219);
xnor U23100 (N_23100,N_21937,N_22404);
or U23101 (N_23101,N_22743,N_22276);
xor U23102 (N_23102,N_21807,N_22320);
nor U23103 (N_23103,N_22236,N_22168);
or U23104 (N_23104,N_22280,N_21621);
nor U23105 (N_23105,N_21831,N_22497);
xor U23106 (N_23106,N_22190,N_22649);
or U23107 (N_23107,N_21750,N_21892);
nand U23108 (N_23108,N_22182,N_22637);
nor U23109 (N_23109,N_22540,N_22710);
or U23110 (N_23110,N_21888,N_21927);
nor U23111 (N_23111,N_22581,N_22623);
nand U23112 (N_23112,N_22685,N_22069);
xnor U23113 (N_23113,N_22423,N_21853);
nor U23114 (N_23114,N_22632,N_22445);
nor U23115 (N_23115,N_21879,N_21947);
or U23116 (N_23116,N_22788,N_22689);
xnor U23117 (N_23117,N_22287,N_21909);
and U23118 (N_23118,N_21815,N_22735);
nor U23119 (N_23119,N_22642,N_22638);
and U23120 (N_23120,N_22465,N_22033);
or U23121 (N_23121,N_21914,N_21976);
and U23122 (N_23122,N_22714,N_22107);
and U23123 (N_23123,N_22703,N_22782);
nor U23124 (N_23124,N_22363,N_21945);
and U23125 (N_23125,N_21647,N_21675);
or U23126 (N_23126,N_22590,N_22744);
or U23127 (N_23127,N_22100,N_22336);
and U23128 (N_23128,N_22414,N_21775);
xnor U23129 (N_23129,N_22277,N_22360);
nand U23130 (N_23130,N_22078,N_22272);
nand U23131 (N_23131,N_22725,N_22347);
nand U23132 (N_23132,N_22223,N_22478);
xnor U23133 (N_23133,N_22048,N_22084);
or U23134 (N_23134,N_22238,N_22374);
nand U23135 (N_23135,N_22288,N_21748);
and U23136 (N_23136,N_22473,N_21794);
xnor U23137 (N_23137,N_22537,N_22640);
or U23138 (N_23138,N_22767,N_22051);
and U23139 (N_23139,N_21726,N_22633);
and U23140 (N_23140,N_22077,N_22135);
and U23141 (N_23141,N_21833,N_21738);
or U23142 (N_23142,N_21786,N_22600);
or U23143 (N_23143,N_22490,N_22212);
nor U23144 (N_23144,N_21886,N_21763);
or U23145 (N_23145,N_22565,N_21682);
nand U23146 (N_23146,N_21758,N_22240);
xnor U23147 (N_23147,N_22663,N_22721);
or U23148 (N_23148,N_21922,N_22426);
nand U23149 (N_23149,N_21884,N_21801);
and U23150 (N_23150,N_22417,N_21697);
xor U23151 (N_23151,N_22147,N_22090);
nor U23152 (N_23152,N_22610,N_22500);
or U23153 (N_23153,N_22019,N_21977);
and U23154 (N_23154,N_22501,N_22210);
nand U23155 (N_23155,N_22102,N_22035);
or U23156 (N_23156,N_22096,N_21615);
nor U23157 (N_23157,N_22534,N_21765);
xor U23158 (N_23158,N_21668,N_22733);
nor U23159 (N_23159,N_22217,N_21618);
or U23160 (N_23160,N_22364,N_21788);
xnor U23161 (N_23161,N_21928,N_22545);
xor U23162 (N_23162,N_22455,N_21846);
nor U23163 (N_23163,N_22315,N_22187);
or U23164 (N_23164,N_22156,N_22085);
nand U23165 (N_23165,N_21995,N_22588);
nor U23166 (N_23166,N_22483,N_22519);
and U23167 (N_23167,N_22088,N_22486);
xnor U23168 (N_23168,N_22602,N_21751);
or U23169 (N_23169,N_22359,N_22068);
nor U23170 (N_23170,N_22004,N_22723);
xor U23171 (N_23171,N_22643,N_21629);
nor U23172 (N_23172,N_22571,N_22214);
xor U23173 (N_23173,N_22342,N_22749);
and U23174 (N_23174,N_21774,N_22667);
nand U23175 (N_23175,N_22245,N_22573);
nand U23176 (N_23176,N_21865,N_22695);
nor U23177 (N_23177,N_22235,N_22129);
and U23178 (N_23178,N_22491,N_22140);
nand U23179 (N_23179,N_22558,N_22447);
or U23180 (N_23180,N_22474,N_22031);
and U23181 (N_23181,N_21978,N_22603);
nand U23182 (N_23182,N_21814,N_21955);
nand U23183 (N_23183,N_22629,N_22071);
xor U23184 (N_23184,N_21943,N_22457);
xor U23185 (N_23185,N_22388,N_21832);
nand U23186 (N_23186,N_21718,N_22294);
xor U23187 (N_23187,N_22110,N_21876);
or U23188 (N_23188,N_21842,N_21651);
xor U23189 (N_23189,N_22299,N_21902);
nor U23190 (N_23190,N_21915,N_21979);
nor U23191 (N_23191,N_21956,N_22221);
and U23192 (N_23192,N_21981,N_22196);
nor U23193 (N_23193,N_21725,N_22065);
xnor U23194 (N_23194,N_22244,N_22555);
or U23195 (N_23195,N_22167,N_22466);
nor U23196 (N_23196,N_22699,N_22366);
nor U23197 (N_23197,N_22766,N_22322);
nor U23198 (N_23198,N_22284,N_22759);
xnor U23199 (N_23199,N_21971,N_22251);
nor U23200 (N_23200,N_22324,N_21670);
and U23201 (N_23201,N_22654,N_22549);
nand U23202 (N_23202,N_21890,N_22003);
nor U23203 (N_23203,N_21910,N_21716);
or U23204 (N_23204,N_21987,N_21715);
nor U23205 (N_23205,N_21809,N_22226);
xnor U23206 (N_23206,N_21683,N_22105);
nor U23207 (N_23207,N_21656,N_21870);
nand U23208 (N_23208,N_22211,N_21854);
xnor U23209 (N_23209,N_21759,N_22613);
or U23210 (N_23210,N_21604,N_22677);
nand U23211 (N_23211,N_22527,N_21818);
nand U23212 (N_23212,N_22687,N_22605);
nor U23213 (N_23213,N_22492,N_21925);
nand U23214 (N_23214,N_22771,N_22660);
nand U23215 (N_23215,N_22467,N_22232);
nor U23216 (N_23216,N_22722,N_22387);
and U23217 (N_23217,N_22340,N_22353);
xor U23218 (N_23218,N_22385,N_22034);
or U23219 (N_23219,N_21839,N_21994);
and U23220 (N_23220,N_21992,N_22383);
xnor U23221 (N_23221,N_22599,N_22313);
and U23222 (N_23222,N_22448,N_22586);
nand U23223 (N_23223,N_22070,N_22304);
or U23224 (N_23224,N_21929,N_21626);
or U23225 (N_23225,N_22337,N_21822);
nand U23226 (N_23226,N_22164,N_22606);
nor U23227 (N_23227,N_22416,N_22452);
xor U23228 (N_23228,N_22578,N_22488);
xnor U23229 (N_23229,N_21799,N_22395);
xor U23230 (N_23230,N_21710,N_22029);
xor U23231 (N_23231,N_22042,N_22318);
nor U23232 (N_23232,N_21734,N_22645);
xor U23233 (N_23233,N_21924,N_22413);
and U23234 (N_23234,N_22150,N_22617);
xor U23235 (N_23235,N_22016,N_21967);
xor U23236 (N_23236,N_22228,N_21898);
and U23237 (N_23237,N_21880,N_21671);
xor U23238 (N_23238,N_22325,N_21911);
xnor U23239 (N_23239,N_22684,N_22017);
xor U23240 (N_23240,N_22180,N_22400);
and U23241 (N_23241,N_22531,N_21946);
nand U23242 (N_23242,N_22583,N_22316);
nor U23243 (N_23243,N_22139,N_22596);
nor U23244 (N_23244,N_22274,N_22128);
xor U23245 (N_23245,N_22170,N_21709);
or U23246 (N_23246,N_22436,N_21931);
xnor U23247 (N_23247,N_22185,N_22428);
nor U23248 (N_23248,N_21753,N_22769);
and U23249 (N_23249,N_22119,N_21658);
nor U23250 (N_23250,N_21777,N_21691);
nand U23251 (N_23251,N_22471,N_21797);
nor U23252 (N_23252,N_22516,N_22379);
and U23253 (N_23253,N_21866,N_22083);
nand U23254 (N_23254,N_21960,N_22470);
nor U23255 (N_23255,N_22092,N_22712);
or U23256 (N_23256,N_21942,N_21631);
and U23257 (N_23257,N_22044,N_21862);
or U23258 (N_23258,N_22248,N_22736);
or U23259 (N_23259,N_22144,N_22594);
nand U23260 (N_23260,N_22007,N_21893);
xor U23261 (N_23261,N_22464,N_21844);
nor U23262 (N_23262,N_22131,N_21612);
nor U23263 (N_23263,N_22551,N_22206);
or U23264 (N_23264,N_22130,N_22412);
nor U23265 (N_23265,N_22230,N_22572);
and U23266 (N_23266,N_22059,N_22433);
nand U23267 (N_23267,N_21986,N_22298);
xor U23268 (N_23268,N_22704,N_21895);
and U23269 (N_23269,N_21772,N_22729);
xnor U23270 (N_23270,N_22700,N_22627);
nand U23271 (N_23271,N_21633,N_22162);
nor U23272 (N_23272,N_22431,N_21701);
and U23273 (N_23273,N_21958,N_22176);
nand U23274 (N_23274,N_21861,N_21949);
or U23275 (N_23275,N_22440,N_22679);
xor U23276 (N_23276,N_21785,N_22224);
and U23277 (N_23277,N_22136,N_22512);
and U23278 (N_23278,N_22015,N_22330);
xnor U23279 (N_23279,N_22127,N_22751);
or U23280 (N_23280,N_22161,N_21803);
or U23281 (N_23281,N_21634,N_21730);
xor U23282 (N_23282,N_21740,N_22246);
nor U23283 (N_23283,N_22040,N_22673);
nor U23284 (N_23284,N_22113,N_22317);
nand U23285 (N_23285,N_21659,N_21711);
xor U23286 (N_23286,N_22757,N_22250);
and U23287 (N_23287,N_22103,N_22584);
xnor U23288 (N_23288,N_22646,N_22727);
xnor U23289 (N_23289,N_21944,N_21988);
nand U23290 (N_23290,N_21645,N_21613);
or U23291 (N_23291,N_22039,N_22459);
nor U23292 (N_23292,N_21973,N_22495);
or U23293 (N_23293,N_22367,N_22138);
nor U23294 (N_23294,N_22126,N_22300);
and U23295 (N_23295,N_21912,N_21760);
or U23296 (N_23296,N_22709,N_22720);
nor U23297 (N_23297,N_21653,N_22348);
xnor U23298 (N_23298,N_22149,N_22765);
or U23299 (N_23299,N_22592,N_22419);
or U23300 (N_23300,N_21605,N_21608);
and U23301 (N_23301,N_21970,N_22213);
nor U23302 (N_23302,N_21900,N_22763);
and U23303 (N_23303,N_22026,N_21714);
or U23304 (N_23304,N_22275,N_22010);
and U23305 (N_23305,N_22620,N_21729);
and U23306 (N_23306,N_22175,N_22442);
or U23307 (N_23307,N_22076,N_21655);
nor U23308 (N_23308,N_22399,N_21934);
or U23309 (N_23309,N_21679,N_22041);
nor U23310 (N_23310,N_22597,N_22741);
or U23311 (N_23311,N_21859,N_22784);
nand U23312 (N_23312,N_21824,N_21723);
nand U23313 (N_23313,N_22580,N_22536);
or U23314 (N_23314,N_22308,N_22165);
or U23315 (N_23315,N_22178,N_21601);
and U23316 (N_23316,N_21707,N_22451);
or U23317 (N_23317,N_21742,N_22087);
and U23318 (N_23318,N_22508,N_22585);
nand U23319 (N_23319,N_22109,N_21778);
nand U23320 (N_23320,N_22713,N_21650);
and U23321 (N_23321,N_22254,N_22137);
nand U23322 (N_23322,N_21617,N_21962);
and U23323 (N_23323,N_22468,N_22522);
nor U23324 (N_23324,N_22651,N_21674);
or U23325 (N_23325,N_21686,N_22427);
nand U23326 (N_23326,N_22195,N_22665);
nor U23327 (N_23327,N_21713,N_22708);
and U23328 (N_23328,N_22652,N_22636);
xor U23329 (N_23329,N_21702,N_21712);
nand U23330 (N_23330,N_21664,N_21918);
xnor U23331 (N_23331,N_21781,N_22271);
nand U23332 (N_23332,N_22732,N_22658);
nor U23333 (N_23333,N_22201,N_22081);
nor U23334 (N_23334,N_21916,N_21733);
xor U23335 (N_23335,N_22121,N_21644);
or U23336 (N_23336,N_22547,N_22056);
nand U23337 (N_23337,N_22420,N_22541);
nand U23338 (N_23338,N_21696,N_22073);
and U23339 (N_23339,N_22631,N_22002);
or U23340 (N_23340,N_21607,N_21998);
xnor U23341 (N_23341,N_22515,N_21637);
nand U23342 (N_23342,N_21952,N_21875);
nand U23343 (N_23343,N_21933,N_21887);
nand U23344 (N_23344,N_21974,N_22189);
and U23345 (N_23345,N_22676,N_22772);
and U23346 (N_23346,N_22706,N_22567);
nand U23347 (N_23347,N_22312,N_21837);
and U23348 (N_23348,N_22334,N_21968);
nand U23349 (N_23349,N_22265,N_21806);
nor U23350 (N_23350,N_22750,N_22099);
nor U23351 (N_23351,N_22415,N_21864);
nor U23352 (N_23352,N_22328,N_22020);
xnor U23353 (N_23353,N_22608,N_22780);
or U23354 (N_23354,N_22698,N_21823);
or U23355 (N_23355,N_22659,N_22243);
nand U23356 (N_23356,N_22283,N_21874);
nand U23357 (N_23357,N_22106,N_21860);
nor U23358 (N_23358,N_21735,N_22582);
and U23359 (N_23359,N_21779,N_22157);
nor U23360 (N_23360,N_21789,N_22382);
or U23361 (N_23361,N_22711,N_22194);
xnor U23362 (N_23362,N_22453,N_22728);
xor U23363 (N_23363,N_21739,N_21966);
xnor U23364 (N_23364,N_22278,N_22267);
xnor U23365 (N_23365,N_22242,N_21808);
nand U23366 (N_23366,N_22798,N_21667);
xor U23367 (N_23367,N_22421,N_22524);
and U23368 (N_23368,N_22543,N_22333);
and U23369 (N_23369,N_22285,N_22289);
nand U23370 (N_23370,N_21771,N_22509);
nor U23371 (N_23371,N_21619,N_21693);
nand U23372 (N_23372,N_22356,N_21913);
nand U23373 (N_23373,N_22734,N_22270);
and U23374 (N_23374,N_22339,N_22548);
nor U23375 (N_23375,N_21923,N_21836);
and U23376 (N_23376,N_22025,N_21885);
nor U23377 (N_23377,N_22668,N_21829);
xor U23378 (N_23378,N_21835,N_22518);
nand U23379 (N_23379,N_21632,N_22117);
nand U23380 (N_23380,N_22675,N_22086);
or U23381 (N_23381,N_21850,N_22611);
and U23382 (N_23382,N_22358,N_22079);
or U23383 (N_23383,N_22648,N_22502);
xor U23384 (N_23384,N_21856,N_22674);
or U23385 (N_23385,N_21999,N_22437);
nor U23386 (N_23386,N_22546,N_22514);
nor U23387 (N_23387,N_22559,N_22331);
or U23388 (N_23388,N_21821,N_22172);
nor U23389 (N_23389,N_22615,N_21643);
xnor U23390 (N_23390,N_22302,N_21989);
xor U23391 (N_23391,N_21648,N_22557);
and U23392 (N_23392,N_22701,N_22513);
xnor U23393 (N_23393,N_22688,N_22030);
or U23394 (N_23394,N_22579,N_22434);
xnor U23395 (N_23395,N_21817,N_21628);
or U23396 (N_23396,N_22575,N_22247);
and U23397 (N_23397,N_21720,N_21953);
nor U23398 (N_23398,N_21638,N_22354);
xnor U23399 (N_23399,N_21611,N_22671);
and U23400 (N_23400,N_21947,N_22540);
nand U23401 (N_23401,N_22162,N_21677);
xnor U23402 (N_23402,N_22395,N_22658);
or U23403 (N_23403,N_22088,N_22361);
nor U23404 (N_23404,N_21884,N_22537);
xor U23405 (N_23405,N_22740,N_21749);
nand U23406 (N_23406,N_22767,N_22480);
or U23407 (N_23407,N_22558,N_22508);
nand U23408 (N_23408,N_22371,N_21930);
and U23409 (N_23409,N_22429,N_22319);
nand U23410 (N_23410,N_22362,N_22211);
or U23411 (N_23411,N_22058,N_22665);
nor U23412 (N_23412,N_22768,N_22004);
and U23413 (N_23413,N_21722,N_21956);
or U23414 (N_23414,N_22288,N_22324);
nor U23415 (N_23415,N_22353,N_22738);
and U23416 (N_23416,N_21924,N_22428);
nor U23417 (N_23417,N_22194,N_21656);
nor U23418 (N_23418,N_22107,N_22147);
and U23419 (N_23419,N_22277,N_22451);
xnor U23420 (N_23420,N_21829,N_22478);
nor U23421 (N_23421,N_22691,N_22020);
and U23422 (N_23422,N_22275,N_22713);
xnor U23423 (N_23423,N_22152,N_22239);
nor U23424 (N_23424,N_22484,N_22506);
xor U23425 (N_23425,N_22185,N_21659);
or U23426 (N_23426,N_22156,N_22763);
and U23427 (N_23427,N_22498,N_22296);
and U23428 (N_23428,N_21779,N_22401);
nand U23429 (N_23429,N_22135,N_21981);
nand U23430 (N_23430,N_22054,N_22098);
nor U23431 (N_23431,N_21817,N_21948);
or U23432 (N_23432,N_22413,N_21654);
xor U23433 (N_23433,N_22192,N_21914);
and U23434 (N_23434,N_22063,N_22547);
nor U23435 (N_23435,N_22285,N_22344);
xnor U23436 (N_23436,N_22583,N_22542);
or U23437 (N_23437,N_22153,N_21767);
nand U23438 (N_23438,N_22150,N_22672);
nand U23439 (N_23439,N_21684,N_21853);
nand U23440 (N_23440,N_22685,N_22404);
nand U23441 (N_23441,N_21873,N_22112);
or U23442 (N_23442,N_22794,N_22176);
and U23443 (N_23443,N_21846,N_22562);
or U23444 (N_23444,N_22588,N_22668);
or U23445 (N_23445,N_21881,N_22484);
nand U23446 (N_23446,N_22642,N_21731);
xor U23447 (N_23447,N_21808,N_22163);
and U23448 (N_23448,N_22760,N_22164);
xor U23449 (N_23449,N_21779,N_21977);
and U23450 (N_23450,N_22399,N_22086);
xor U23451 (N_23451,N_21642,N_21772);
xnor U23452 (N_23452,N_22278,N_22072);
nand U23453 (N_23453,N_22617,N_21740);
and U23454 (N_23454,N_21694,N_22295);
nor U23455 (N_23455,N_21993,N_22243);
and U23456 (N_23456,N_22578,N_22590);
and U23457 (N_23457,N_22125,N_22382);
xnor U23458 (N_23458,N_22213,N_21679);
and U23459 (N_23459,N_22691,N_21666);
nand U23460 (N_23460,N_21972,N_21628);
xor U23461 (N_23461,N_22742,N_22630);
and U23462 (N_23462,N_22217,N_22771);
nor U23463 (N_23463,N_21794,N_22095);
and U23464 (N_23464,N_22063,N_22462);
nor U23465 (N_23465,N_21725,N_21753);
and U23466 (N_23466,N_22791,N_22432);
nor U23467 (N_23467,N_21940,N_22230);
and U23468 (N_23468,N_22642,N_21609);
or U23469 (N_23469,N_22457,N_22132);
and U23470 (N_23470,N_22124,N_21967);
xnor U23471 (N_23471,N_22427,N_22524);
nand U23472 (N_23472,N_22409,N_21888);
or U23473 (N_23473,N_22115,N_22191);
and U23474 (N_23474,N_21954,N_22745);
nor U23475 (N_23475,N_22332,N_21977);
xnor U23476 (N_23476,N_21782,N_22234);
and U23477 (N_23477,N_21931,N_21918);
and U23478 (N_23478,N_21954,N_21931);
or U23479 (N_23479,N_22005,N_22464);
xnor U23480 (N_23480,N_22097,N_22436);
and U23481 (N_23481,N_22329,N_22355);
xnor U23482 (N_23482,N_22244,N_22481);
nand U23483 (N_23483,N_22279,N_22252);
or U23484 (N_23484,N_21821,N_21932);
and U23485 (N_23485,N_21624,N_22560);
nor U23486 (N_23486,N_22411,N_22144);
nor U23487 (N_23487,N_21969,N_21986);
and U23488 (N_23488,N_21716,N_21885);
or U23489 (N_23489,N_21787,N_22265);
and U23490 (N_23490,N_22180,N_21610);
or U23491 (N_23491,N_21704,N_22654);
xor U23492 (N_23492,N_22299,N_21736);
nor U23493 (N_23493,N_22522,N_22739);
or U23494 (N_23494,N_22367,N_22186);
or U23495 (N_23495,N_21736,N_21915);
nand U23496 (N_23496,N_22663,N_22246);
or U23497 (N_23497,N_22183,N_22256);
and U23498 (N_23498,N_22360,N_22392);
or U23499 (N_23499,N_22087,N_22614);
nand U23500 (N_23500,N_22469,N_22366);
xor U23501 (N_23501,N_22765,N_21701);
xor U23502 (N_23502,N_22667,N_22599);
or U23503 (N_23503,N_22377,N_21652);
nand U23504 (N_23504,N_22681,N_21629);
and U23505 (N_23505,N_22131,N_22644);
and U23506 (N_23506,N_22051,N_22681);
and U23507 (N_23507,N_21664,N_21758);
nor U23508 (N_23508,N_22570,N_22640);
xnor U23509 (N_23509,N_22071,N_22259);
xor U23510 (N_23510,N_22547,N_22424);
or U23511 (N_23511,N_21708,N_22757);
xnor U23512 (N_23512,N_22558,N_22330);
or U23513 (N_23513,N_22466,N_22427);
nor U23514 (N_23514,N_22103,N_21759);
and U23515 (N_23515,N_22567,N_21983);
and U23516 (N_23516,N_22791,N_22221);
and U23517 (N_23517,N_22324,N_21858);
xnor U23518 (N_23518,N_21946,N_21765);
or U23519 (N_23519,N_22572,N_22430);
nand U23520 (N_23520,N_22308,N_22157);
xor U23521 (N_23521,N_22595,N_22168);
and U23522 (N_23522,N_22105,N_21831);
xnor U23523 (N_23523,N_22218,N_22206);
or U23524 (N_23524,N_22231,N_22224);
nor U23525 (N_23525,N_22760,N_21659);
or U23526 (N_23526,N_21780,N_22436);
or U23527 (N_23527,N_21622,N_22439);
nand U23528 (N_23528,N_22467,N_22569);
xnor U23529 (N_23529,N_21983,N_22522);
and U23530 (N_23530,N_22080,N_22770);
or U23531 (N_23531,N_22406,N_22600);
and U23532 (N_23532,N_21661,N_22090);
or U23533 (N_23533,N_22178,N_22055);
nand U23534 (N_23534,N_22479,N_21902);
nor U23535 (N_23535,N_22265,N_22649);
nor U23536 (N_23536,N_22518,N_21605);
xnor U23537 (N_23537,N_22625,N_21728);
nor U23538 (N_23538,N_21671,N_22652);
xor U23539 (N_23539,N_22098,N_21832);
nand U23540 (N_23540,N_22043,N_22228);
and U23541 (N_23541,N_22438,N_21603);
nand U23542 (N_23542,N_22777,N_22113);
nor U23543 (N_23543,N_22158,N_22056);
nand U23544 (N_23544,N_22146,N_22586);
nor U23545 (N_23545,N_22202,N_22515);
and U23546 (N_23546,N_22183,N_21910);
nand U23547 (N_23547,N_21712,N_22788);
or U23548 (N_23548,N_22155,N_22521);
xnor U23549 (N_23549,N_21966,N_21831);
nand U23550 (N_23550,N_21868,N_21827);
or U23551 (N_23551,N_21770,N_22660);
nand U23552 (N_23552,N_22087,N_22385);
or U23553 (N_23553,N_21782,N_22135);
nor U23554 (N_23554,N_22591,N_22250);
xor U23555 (N_23555,N_22438,N_22114);
nor U23556 (N_23556,N_22161,N_22297);
nor U23557 (N_23557,N_22523,N_22732);
and U23558 (N_23558,N_22016,N_21883);
xor U23559 (N_23559,N_22488,N_21881);
and U23560 (N_23560,N_22482,N_22634);
xor U23561 (N_23561,N_22296,N_21872);
xor U23562 (N_23562,N_22454,N_22630);
and U23563 (N_23563,N_22117,N_22684);
nor U23564 (N_23564,N_21691,N_22659);
or U23565 (N_23565,N_22315,N_22389);
and U23566 (N_23566,N_21685,N_22091);
and U23567 (N_23567,N_22196,N_22667);
and U23568 (N_23568,N_22518,N_21981);
and U23569 (N_23569,N_22591,N_22045);
and U23570 (N_23570,N_22004,N_22735);
or U23571 (N_23571,N_22617,N_22710);
nor U23572 (N_23572,N_21754,N_21837);
xor U23573 (N_23573,N_22082,N_21885);
xnor U23574 (N_23574,N_22426,N_21986);
xor U23575 (N_23575,N_22605,N_22381);
nor U23576 (N_23576,N_21688,N_22400);
or U23577 (N_23577,N_22730,N_21648);
and U23578 (N_23578,N_22129,N_21695);
xor U23579 (N_23579,N_21854,N_22250);
and U23580 (N_23580,N_22655,N_21630);
xnor U23581 (N_23581,N_21946,N_21841);
or U23582 (N_23582,N_22479,N_22138);
nor U23583 (N_23583,N_22687,N_22639);
xor U23584 (N_23584,N_22481,N_22568);
xnor U23585 (N_23585,N_21802,N_21704);
or U23586 (N_23586,N_21853,N_22277);
nand U23587 (N_23587,N_22694,N_21899);
or U23588 (N_23588,N_21987,N_22064);
nand U23589 (N_23589,N_22139,N_21641);
nand U23590 (N_23590,N_22629,N_22586);
and U23591 (N_23591,N_21787,N_22003);
or U23592 (N_23592,N_21697,N_22386);
nor U23593 (N_23593,N_21847,N_22345);
xnor U23594 (N_23594,N_22363,N_22358);
and U23595 (N_23595,N_22464,N_22313);
nand U23596 (N_23596,N_22583,N_22732);
and U23597 (N_23597,N_22500,N_22069);
or U23598 (N_23598,N_22429,N_22058);
nand U23599 (N_23599,N_22510,N_21826);
and U23600 (N_23600,N_22102,N_21798);
or U23601 (N_23601,N_21831,N_21807);
and U23602 (N_23602,N_22148,N_22344);
and U23603 (N_23603,N_22193,N_22231);
nor U23604 (N_23604,N_21607,N_22764);
xor U23605 (N_23605,N_22474,N_22691);
nand U23606 (N_23606,N_22441,N_21884);
xnor U23607 (N_23607,N_21612,N_22565);
and U23608 (N_23608,N_21884,N_22214);
or U23609 (N_23609,N_22183,N_21987);
nor U23610 (N_23610,N_21647,N_21762);
and U23611 (N_23611,N_22457,N_21745);
xor U23612 (N_23612,N_22739,N_21894);
xor U23613 (N_23613,N_22603,N_21823);
xor U23614 (N_23614,N_22612,N_22311);
xnor U23615 (N_23615,N_22738,N_21900);
nand U23616 (N_23616,N_22550,N_22597);
xnor U23617 (N_23617,N_21983,N_21774);
nand U23618 (N_23618,N_22390,N_22007);
nand U23619 (N_23619,N_22454,N_21766);
and U23620 (N_23620,N_22454,N_22223);
xor U23621 (N_23621,N_22453,N_22403);
xor U23622 (N_23622,N_22776,N_22016);
or U23623 (N_23623,N_22488,N_22145);
or U23624 (N_23624,N_22644,N_21654);
or U23625 (N_23625,N_22353,N_22342);
and U23626 (N_23626,N_21728,N_22010);
and U23627 (N_23627,N_21861,N_22608);
nand U23628 (N_23628,N_22762,N_21997);
or U23629 (N_23629,N_21628,N_22054);
nand U23630 (N_23630,N_21828,N_22417);
xor U23631 (N_23631,N_22660,N_22048);
nor U23632 (N_23632,N_22300,N_22718);
or U23633 (N_23633,N_22152,N_22467);
and U23634 (N_23634,N_22327,N_22135);
and U23635 (N_23635,N_22096,N_22494);
xnor U23636 (N_23636,N_22774,N_22402);
xnor U23637 (N_23637,N_22606,N_22200);
or U23638 (N_23638,N_21980,N_21905);
nand U23639 (N_23639,N_22762,N_21976);
and U23640 (N_23640,N_21857,N_22427);
xnor U23641 (N_23641,N_21926,N_22041);
nor U23642 (N_23642,N_22183,N_22776);
and U23643 (N_23643,N_21912,N_22230);
nand U23644 (N_23644,N_22477,N_22630);
nand U23645 (N_23645,N_22485,N_21689);
nand U23646 (N_23646,N_22201,N_21692);
xor U23647 (N_23647,N_22573,N_21951);
and U23648 (N_23648,N_21763,N_21686);
xnor U23649 (N_23649,N_22592,N_21752);
and U23650 (N_23650,N_22413,N_22652);
or U23651 (N_23651,N_21600,N_22394);
nand U23652 (N_23652,N_22781,N_22056);
and U23653 (N_23653,N_22440,N_22680);
and U23654 (N_23654,N_22438,N_22101);
nor U23655 (N_23655,N_21990,N_21634);
and U23656 (N_23656,N_22694,N_21755);
nor U23657 (N_23657,N_22308,N_22303);
xor U23658 (N_23658,N_22630,N_21889);
or U23659 (N_23659,N_22043,N_22663);
or U23660 (N_23660,N_22614,N_21674);
and U23661 (N_23661,N_21868,N_22332);
xor U23662 (N_23662,N_22025,N_22394);
nor U23663 (N_23663,N_22737,N_22252);
xnor U23664 (N_23664,N_21897,N_22263);
nand U23665 (N_23665,N_22530,N_21973);
nand U23666 (N_23666,N_22571,N_21885);
and U23667 (N_23667,N_21763,N_21608);
and U23668 (N_23668,N_21788,N_22032);
xnor U23669 (N_23669,N_22790,N_21801);
nor U23670 (N_23670,N_22438,N_21851);
and U23671 (N_23671,N_21704,N_22697);
or U23672 (N_23672,N_21727,N_22403);
nand U23673 (N_23673,N_22796,N_22450);
xor U23674 (N_23674,N_21926,N_22495);
xor U23675 (N_23675,N_22006,N_22324);
nor U23676 (N_23676,N_22593,N_22403);
or U23677 (N_23677,N_22349,N_22231);
xor U23678 (N_23678,N_22364,N_22244);
nor U23679 (N_23679,N_21754,N_22099);
or U23680 (N_23680,N_22216,N_21962);
nand U23681 (N_23681,N_21615,N_22333);
nand U23682 (N_23682,N_22517,N_21787);
nor U23683 (N_23683,N_22399,N_21787);
and U23684 (N_23684,N_21779,N_21915);
or U23685 (N_23685,N_22525,N_22699);
or U23686 (N_23686,N_22452,N_21842);
and U23687 (N_23687,N_21685,N_21666);
nand U23688 (N_23688,N_22138,N_22450);
or U23689 (N_23689,N_21881,N_22093);
nand U23690 (N_23690,N_22022,N_22592);
nor U23691 (N_23691,N_22626,N_22031);
or U23692 (N_23692,N_22439,N_22111);
and U23693 (N_23693,N_22203,N_21848);
xnor U23694 (N_23694,N_21603,N_21963);
nand U23695 (N_23695,N_22030,N_22672);
xnor U23696 (N_23696,N_21682,N_22392);
or U23697 (N_23697,N_22630,N_22764);
or U23698 (N_23698,N_22219,N_21685);
nor U23699 (N_23699,N_22265,N_22362);
or U23700 (N_23700,N_21984,N_22218);
nand U23701 (N_23701,N_22376,N_22097);
xnor U23702 (N_23702,N_22260,N_22540);
and U23703 (N_23703,N_22469,N_21992);
or U23704 (N_23704,N_22334,N_22488);
or U23705 (N_23705,N_22226,N_22079);
nand U23706 (N_23706,N_22117,N_22261);
and U23707 (N_23707,N_22474,N_21693);
or U23708 (N_23708,N_22705,N_22326);
nor U23709 (N_23709,N_21672,N_22410);
nor U23710 (N_23710,N_21820,N_22177);
xnor U23711 (N_23711,N_21688,N_21706);
or U23712 (N_23712,N_21654,N_22591);
and U23713 (N_23713,N_22228,N_21755);
xnor U23714 (N_23714,N_22024,N_22789);
or U23715 (N_23715,N_21625,N_22622);
xor U23716 (N_23716,N_21640,N_22057);
nor U23717 (N_23717,N_22401,N_22535);
and U23718 (N_23718,N_22162,N_22730);
and U23719 (N_23719,N_22595,N_22235);
or U23720 (N_23720,N_21995,N_21745);
and U23721 (N_23721,N_22269,N_22209);
xnor U23722 (N_23722,N_22514,N_22390);
and U23723 (N_23723,N_21726,N_21987);
nor U23724 (N_23724,N_22674,N_22485);
nand U23725 (N_23725,N_22332,N_22482);
nand U23726 (N_23726,N_22771,N_22282);
xor U23727 (N_23727,N_21941,N_21866);
nor U23728 (N_23728,N_22141,N_22243);
nand U23729 (N_23729,N_21766,N_22179);
nor U23730 (N_23730,N_22610,N_21757);
nor U23731 (N_23731,N_21744,N_22276);
or U23732 (N_23732,N_22522,N_22093);
nand U23733 (N_23733,N_22008,N_22111);
nand U23734 (N_23734,N_21763,N_21951);
nor U23735 (N_23735,N_21790,N_21837);
or U23736 (N_23736,N_22394,N_21692);
xor U23737 (N_23737,N_22253,N_21859);
and U23738 (N_23738,N_21952,N_21688);
xnor U23739 (N_23739,N_22171,N_22629);
nor U23740 (N_23740,N_22285,N_21814);
xor U23741 (N_23741,N_22449,N_22513);
xor U23742 (N_23742,N_21828,N_22145);
nand U23743 (N_23743,N_21809,N_22107);
nand U23744 (N_23744,N_22741,N_22795);
xnor U23745 (N_23745,N_22017,N_21898);
or U23746 (N_23746,N_22358,N_22160);
xnor U23747 (N_23747,N_21657,N_21787);
or U23748 (N_23748,N_21687,N_21650);
xor U23749 (N_23749,N_22585,N_22203);
and U23750 (N_23750,N_22664,N_21753);
xor U23751 (N_23751,N_21607,N_21842);
and U23752 (N_23752,N_22163,N_21955);
nor U23753 (N_23753,N_22085,N_21636);
xnor U23754 (N_23754,N_21878,N_21911);
nor U23755 (N_23755,N_22237,N_22232);
or U23756 (N_23756,N_22293,N_21965);
nor U23757 (N_23757,N_22317,N_22412);
nand U23758 (N_23758,N_21895,N_22654);
nor U23759 (N_23759,N_22134,N_22586);
xor U23760 (N_23760,N_21726,N_22597);
nor U23761 (N_23761,N_21843,N_21762);
or U23762 (N_23762,N_22496,N_22215);
xor U23763 (N_23763,N_22146,N_21944);
nor U23764 (N_23764,N_22020,N_22660);
and U23765 (N_23765,N_22256,N_21754);
or U23766 (N_23766,N_22221,N_22570);
or U23767 (N_23767,N_22169,N_22321);
nor U23768 (N_23768,N_22181,N_21835);
or U23769 (N_23769,N_21964,N_22299);
or U23770 (N_23770,N_21729,N_22297);
nand U23771 (N_23771,N_21614,N_21675);
or U23772 (N_23772,N_22401,N_22247);
or U23773 (N_23773,N_22211,N_22414);
nand U23774 (N_23774,N_22542,N_21999);
nor U23775 (N_23775,N_21842,N_22676);
and U23776 (N_23776,N_21985,N_21790);
nand U23777 (N_23777,N_22158,N_22223);
nand U23778 (N_23778,N_21844,N_22519);
nand U23779 (N_23779,N_21795,N_21630);
nand U23780 (N_23780,N_22354,N_21611);
nor U23781 (N_23781,N_21725,N_22285);
nand U23782 (N_23782,N_22648,N_21758);
xor U23783 (N_23783,N_22276,N_21638);
nor U23784 (N_23784,N_22299,N_21883);
nand U23785 (N_23785,N_22796,N_22272);
nand U23786 (N_23786,N_22649,N_22199);
and U23787 (N_23787,N_22268,N_22396);
and U23788 (N_23788,N_21981,N_21813);
nand U23789 (N_23789,N_22586,N_21704);
or U23790 (N_23790,N_22096,N_22280);
nand U23791 (N_23791,N_22209,N_22232);
and U23792 (N_23792,N_21972,N_21786);
nand U23793 (N_23793,N_22356,N_22150);
and U23794 (N_23794,N_21899,N_22419);
nand U23795 (N_23795,N_22662,N_22761);
xnor U23796 (N_23796,N_21854,N_22700);
or U23797 (N_23797,N_22151,N_22534);
and U23798 (N_23798,N_22748,N_22517);
xnor U23799 (N_23799,N_22508,N_21993);
or U23800 (N_23800,N_22757,N_22235);
or U23801 (N_23801,N_21973,N_22632);
xor U23802 (N_23802,N_22406,N_22207);
nand U23803 (N_23803,N_22555,N_21761);
or U23804 (N_23804,N_22047,N_22794);
nand U23805 (N_23805,N_22393,N_21850);
nand U23806 (N_23806,N_22105,N_21648);
xnor U23807 (N_23807,N_22384,N_21709);
nand U23808 (N_23808,N_22335,N_22782);
xor U23809 (N_23809,N_21962,N_22703);
or U23810 (N_23810,N_22402,N_22677);
xor U23811 (N_23811,N_22221,N_21663);
nand U23812 (N_23812,N_22145,N_22097);
and U23813 (N_23813,N_22535,N_22091);
nand U23814 (N_23814,N_21723,N_22203);
nor U23815 (N_23815,N_21972,N_22450);
xor U23816 (N_23816,N_22002,N_22335);
nor U23817 (N_23817,N_21908,N_21748);
and U23818 (N_23818,N_22372,N_22436);
xor U23819 (N_23819,N_22409,N_22581);
nor U23820 (N_23820,N_22760,N_22465);
nor U23821 (N_23821,N_22569,N_21830);
nor U23822 (N_23822,N_21775,N_22537);
nand U23823 (N_23823,N_22547,N_22115);
and U23824 (N_23824,N_21843,N_22130);
or U23825 (N_23825,N_21646,N_22521);
nand U23826 (N_23826,N_22335,N_21627);
and U23827 (N_23827,N_22231,N_22265);
or U23828 (N_23828,N_22403,N_22538);
and U23829 (N_23829,N_22375,N_22035);
and U23830 (N_23830,N_21622,N_22489);
and U23831 (N_23831,N_22676,N_21609);
nand U23832 (N_23832,N_22309,N_22747);
and U23833 (N_23833,N_22368,N_21941);
and U23834 (N_23834,N_22720,N_21615);
or U23835 (N_23835,N_21693,N_22101);
xor U23836 (N_23836,N_22565,N_22024);
xnor U23837 (N_23837,N_21609,N_22492);
nor U23838 (N_23838,N_22725,N_22148);
and U23839 (N_23839,N_21837,N_22789);
xor U23840 (N_23840,N_21765,N_22352);
nand U23841 (N_23841,N_21766,N_21674);
nand U23842 (N_23842,N_22579,N_21731);
nand U23843 (N_23843,N_22613,N_22391);
or U23844 (N_23844,N_22136,N_22717);
and U23845 (N_23845,N_22684,N_22793);
or U23846 (N_23846,N_21770,N_21685);
and U23847 (N_23847,N_21985,N_22240);
and U23848 (N_23848,N_22749,N_22521);
and U23849 (N_23849,N_22171,N_21954);
and U23850 (N_23850,N_22728,N_22527);
or U23851 (N_23851,N_22113,N_22082);
or U23852 (N_23852,N_22517,N_22753);
and U23853 (N_23853,N_22059,N_22606);
nand U23854 (N_23854,N_22207,N_22545);
or U23855 (N_23855,N_21996,N_22519);
or U23856 (N_23856,N_21640,N_22486);
xor U23857 (N_23857,N_21671,N_22516);
and U23858 (N_23858,N_22012,N_22627);
nand U23859 (N_23859,N_22533,N_21646);
xor U23860 (N_23860,N_21684,N_22175);
and U23861 (N_23861,N_22103,N_21764);
nor U23862 (N_23862,N_22050,N_22618);
nor U23863 (N_23863,N_22410,N_22477);
nand U23864 (N_23864,N_22099,N_21908);
or U23865 (N_23865,N_22548,N_21821);
or U23866 (N_23866,N_22662,N_22410);
xor U23867 (N_23867,N_21711,N_21963);
nand U23868 (N_23868,N_22092,N_22225);
nor U23869 (N_23869,N_22770,N_22550);
nand U23870 (N_23870,N_22171,N_21813);
and U23871 (N_23871,N_22663,N_22794);
nand U23872 (N_23872,N_22495,N_21664);
and U23873 (N_23873,N_21792,N_22724);
and U23874 (N_23874,N_22475,N_22007);
or U23875 (N_23875,N_22132,N_21819);
or U23876 (N_23876,N_22361,N_21728);
nor U23877 (N_23877,N_22624,N_22090);
xor U23878 (N_23878,N_22443,N_22278);
nand U23879 (N_23879,N_22671,N_22422);
and U23880 (N_23880,N_22174,N_21858);
or U23881 (N_23881,N_22573,N_21924);
nor U23882 (N_23882,N_22511,N_22595);
nand U23883 (N_23883,N_22428,N_22594);
nand U23884 (N_23884,N_22257,N_22516);
or U23885 (N_23885,N_21803,N_22433);
nand U23886 (N_23886,N_21917,N_22420);
nand U23887 (N_23887,N_22692,N_21694);
xor U23888 (N_23888,N_21752,N_21663);
or U23889 (N_23889,N_21866,N_22300);
nand U23890 (N_23890,N_22424,N_22322);
or U23891 (N_23891,N_22610,N_22490);
and U23892 (N_23892,N_21927,N_22484);
and U23893 (N_23893,N_21689,N_22735);
nand U23894 (N_23894,N_22036,N_21606);
xnor U23895 (N_23895,N_22694,N_21948);
nand U23896 (N_23896,N_22235,N_22492);
xnor U23897 (N_23897,N_22629,N_22442);
nand U23898 (N_23898,N_22714,N_22603);
or U23899 (N_23899,N_22619,N_22179);
nand U23900 (N_23900,N_22709,N_21833);
nor U23901 (N_23901,N_21753,N_22165);
nand U23902 (N_23902,N_22685,N_22088);
and U23903 (N_23903,N_21879,N_21699);
or U23904 (N_23904,N_22267,N_22214);
xor U23905 (N_23905,N_21876,N_22216);
nor U23906 (N_23906,N_22406,N_22515);
xor U23907 (N_23907,N_22003,N_22109);
xnor U23908 (N_23908,N_22765,N_22018);
nand U23909 (N_23909,N_22138,N_22017);
nor U23910 (N_23910,N_21869,N_22187);
nand U23911 (N_23911,N_22199,N_21758);
and U23912 (N_23912,N_22657,N_21829);
xor U23913 (N_23913,N_21740,N_22754);
and U23914 (N_23914,N_22199,N_22027);
xor U23915 (N_23915,N_21981,N_22600);
nand U23916 (N_23916,N_22375,N_22192);
nor U23917 (N_23917,N_22498,N_21968);
nand U23918 (N_23918,N_22182,N_22359);
and U23919 (N_23919,N_22320,N_22255);
nor U23920 (N_23920,N_22035,N_22396);
and U23921 (N_23921,N_22026,N_21679);
nand U23922 (N_23922,N_22007,N_21966);
and U23923 (N_23923,N_21738,N_21867);
or U23924 (N_23924,N_21824,N_22693);
and U23925 (N_23925,N_22330,N_22291);
nor U23926 (N_23926,N_22640,N_22220);
xnor U23927 (N_23927,N_22466,N_22414);
nand U23928 (N_23928,N_22408,N_22730);
and U23929 (N_23929,N_22763,N_22662);
or U23930 (N_23930,N_22150,N_21787);
and U23931 (N_23931,N_22443,N_21827);
nand U23932 (N_23932,N_22792,N_22689);
and U23933 (N_23933,N_22786,N_21668);
nor U23934 (N_23934,N_21769,N_22295);
and U23935 (N_23935,N_22589,N_21992);
or U23936 (N_23936,N_21796,N_22552);
nand U23937 (N_23937,N_21848,N_22787);
xor U23938 (N_23938,N_22101,N_22172);
or U23939 (N_23939,N_22545,N_22747);
or U23940 (N_23940,N_22421,N_22742);
or U23941 (N_23941,N_21803,N_22051);
nor U23942 (N_23942,N_21796,N_22556);
and U23943 (N_23943,N_22580,N_21661);
nor U23944 (N_23944,N_21623,N_21914);
xnor U23945 (N_23945,N_21822,N_21782);
nor U23946 (N_23946,N_22543,N_22736);
or U23947 (N_23947,N_22622,N_22028);
and U23948 (N_23948,N_21908,N_22581);
nand U23949 (N_23949,N_22459,N_21846);
or U23950 (N_23950,N_22354,N_22592);
xnor U23951 (N_23951,N_21885,N_22233);
nor U23952 (N_23952,N_21957,N_22488);
nand U23953 (N_23953,N_22587,N_21915);
nor U23954 (N_23954,N_22250,N_21746);
xor U23955 (N_23955,N_21954,N_22300);
nor U23956 (N_23956,N_22233,N_22526);
and U23957 (N_23957,N_22323,N_22285);
nor U23958 (N_23958,N_22011,N_22419);
xor U23959 (N_23959,N_21616,N_22027);
and U23960 (N_23960,N_22629,N_22409);
xor U23961 (N_23961,N_22754,N_22257);
nor U23962 (N_23962,N_22019,N_21603);
nand U23963 (N_23963,N_21844,N_22770);
and U23964 (N_23964,N_22108,N_22781);
nand U23965 (N_23965,N_21661,N_22723);
and U23966 (N_23966,N_22175,N_21672);
or U23967 (N_23967,N_22173,N_22451);
nand U23968 (N_23968,N_22576,N_21658);
or U23969 (N_23969,N_22134,N_22362);
nor U23970 (N_23970,N_22157,N_22321);
nand U23971 (N_23971,N_22106,N_22232);
xor U23972 (N_23972,N_22494,N_22413);
nand U23973 (N_23973,N_22650,N_22294);
nand U23974 (N_23974,N_22512,N_22469);
nand U23975 (N_23975,N_22446,N_22583);
xnor U23976 (N_23976,N_22429,N_22517);
nand U23977 (N_23977,N_22432,N_22777);
or U23978 (N_23978,N_22059,N_21821);
xor U23979 (N_23979,N_22187,N_22137);
and U23980 (N_23980,N_21932,N_22038);
nor U23981 (N_23981,N_21841,N_22097);
xnor U23982 (N_23982,N_22428,N_22174);
or U23983 (N_23983,N_22468,N_22039);
nand U23984 (N_23984,N_22006,N_21607);
and U23985 (N_23985,N_22217,N_22547);
nand U23986 (N_23986,N_22153,N_21779);
nor U23987 (N_23987,N_22602,N_22209);
or U23988 (N_23988,N_22043,N_22218);
nor U23989 (N_23989,N_22562,N_22294);
and U23990 (N_23990,N_21683,N_21809);
xor U23991 (N_23991,N_22748,N_22070);
nand U23992 (N_23992,N_22163,N_22642);
xor U23993 (N_23993,N_22027,N_22694);
or U23994 (N_23994,N_21975,N_22023);
and U23995 (N_23995,N_21874,N_21930);
nand U23996 (N_23996,N_22125,N_22474);
nand U23997 (N_23997,N_22521,N_21849);
nand U23998 (N_23998,N_21969,N_21771);
or U23999 (N_23999,N_22108,N_21897);
or U24000 (N_24000,N_23208,N_23201);
xor U24001 (N_24001,N_23041,N_23516);
and U24002 (N_24002,N_23794,N_23589);
nand U24003 (N_24003,N_23407,N_23043);
and U24004 (N_24004,N_23062,N_23129);
or U24005 (N_24005,N_23312,N_23469);
and U24006 (N_24006,N_22871,N_23136);
xor U24007 (N_24007,N_23333,N_23602);
or U24008 (N_24008,N_23953,N_22837);
nor U24009 (N_24009,N_23834,N_23566);
or U24010 (N_24010,N_23527,N_23993);
nand U24011 (N_24011,N_23188,N_23619);
nor U24012 (N_24012,N_23678,N_23500);
nand U24013 (N_24013,N_23263,N_23587);
and U24014 (N_24014,N_23276,N_23184);
or U24015 (N_24015,N_23542,N_22948);
or U24016 (N_24016,N_23326,N_23650);
xor U24017 (N_24017,N_23811,N_23091);
nor U24018 (N_24018,N_23557,N_22829);
nor U24019 (N_24019,N_22889,N_23064);
or U24020 (N_24020,N_23777,N_23849);
and U24021 (N_24021,N_23252,N_23710);
and U24022 (N_24022,N_23440,N_22885);
and U24023 (N_24023,N_23689,N_23969);
nand U24024 (N_24024,N_23306,N_23726);
nor U24025 (N_24025,N_23102,N_22944);
nand U24026 (N_24026,N_22857,N_23829);
nor U24027 (N_24027,N_23693,N_22867);
nor U24028 (N_24028,N_23765,N_23686);
or U24029 (N_24029,N_23768,N_22888);
xnor U24030 (N_24030,N_23151,N_23809);
or U24031 (N_24031,N_23004,N_23304);
xnor U24032 (N_24032,N_23732,N_23265);
nand U24033 (N_24033,N_23892,N_22905);
nand U24034 (N_24034,N_23808,N_23747);
xor U24035 (N_24035,N_23198,N_23165);
or U24036 (N_24036,N_22864,N_23416);
and U24037 (N_24037,N_23528,N_23127);
or U24038 (N_24038,N_23438,N_23949);
xnor U24039 (N_24039,N_23753,N_23121);
nand U24040 (N_24040,N_23696,N_23011);
or U24041 (N_24041,N_23523,N_22813);
nand U24042 (N_24042,N_23393,N_23670);
and U24043 (N_24043,N_23618,N_22958);
or U24044 (N_24044,N_23508,N_23124);
xor U24045 (N_24045,N_23952,N_23613);
nand U24046 (N_24046,N_23632,N_23712);
and U24047 (N_24047,N_23247,N_23044);
or U24048 (N_24048,N_23234,N_23430);
and U24049 (N_24049,N_23140,N_22818);
or U24050 (N_24050,N_23189,N_23859);
nor U24051 (N_24051,N_23793,N_23708);
xor U24052 (N_24052,N_23106,N_22927);
nor U24053 (N_24053,N_23873,N_23323);
xor U24054 (N_24054,N_23420,N_23085);
xor U24055 (N_24055,N_23958,N_23588);
and U24056 (N_24056,N_23431,N_23212);
and U24057 (N_24057,N_23956,N_23100);
and U24058 (N_24058,N_23244,N_23453);
and U24059 (N_24059,N_22843,N_23770);
xnor U24060 (N_24060,N_23219,N_23042);
or U24061 (N_24061,N_23422,N_23680);
xor U24062 (N_24062,N_23965,N_22940);
and U24063 (N_24063,N_23296,N_23737);
or U24064 (N_24064,N_22982,N_23446);
xnor U24065 (N_24065,N_23423,N_23402);
and U24066 (N_24066,N_23351,N_22997);
or U24067 (N_24067,N_22898,N_23027);
nor U24068 (N_24068,N_23851,N_23384);
or U24069 (N_24069,N_22956,N_23985);
and U24070 (N_24070,N_23633,N_23917);
or U24071 (N_24071,N_23879,N_23719);
nand U24072 (N_24072,N_23551,N_23149);
xor U24073 (N_24073,N_23659,N_22988);
and U24074 (N_24074,N_23382,N_23331);
and U24075 (N_24075,N_23218,N_23979);
and U24076 (N_24076,N_23321,N_23534);
or U24077 (N_24077,N_23720,N_23311);
or U24078 (N_24078,N_22833,N_22930);
or U24079 (N_24079,N_23817,N_22943);
or U24080 (N_24080,N_23825,N_23377);
xor U24081 (N_24081,N_23517,N_22968);
nand U24082 (N_24082,N_23303,N_22907);
and U24083 (N_24083,N_23773,N_23550);
xnor U24084 (N_24084,N_23223,N_23146);
nor U24085 (N_24085,N_23577,N_23891);
and U24086 (N_24086,N_22990,N_23068);
nand U24087 (N_24087,N_23755,N_23795);
or U24088 (N_24088,N_23474,N_22860);
nor U24089 (N_24089,N_23485,N_22935);
nor U24090 (N_24090,N_22804,N_23666);
nor U24091 (N_24091,N_23052,N_23139);
and U24092 (N_24092,N_23622,N_23275);
or U24093 (N_24093,N_23886,N_23270);
xnor U24094 (N_24094,N_23461,N_23803);
or U24095 (N_24095,N_23078,N_23575);
nor U24096 (N_24096,N_23338,N_23473);
nand U24097 (N_24097,N_23487,N_23850);
xor U24098 (N_24098,N_23537,N_23204);
nand U24099 (N_24099,N_23114,N_23977);
nor U24100 (N_24100,N_23974,N_23012);
or U24101 (N_24101,N_23049,N_23955);
xnor U24102 (N_24102,N_23681,N_23230);
and U24103 (N_24103,N_22895,N_23273);
and U24104 (N_24104,N_23490,N_22932);
or U24105 (N_24105,N_23518,N_23111);
xor U24106 (N_24106,N_23653,N_23397);
or U24107 (N_24107,N_23168,N_23801);
and U24108 (N_24108,N_22917,N_23771);
and U24109 (N_24109,N_23606,N_23635);
nor U24110 (N_24110,N_23443,N_23983);
or U24111 (N_24111,N_23480,N_22892);
and U24112 (N_24112,N_23307,N_23617);
nor U24113 (N_24113,N_22815,N_23915);
nor U24114 (N_24114,N_23791,N_22900);
nand U24115 (N_24115,N_23596,N_22811);
nor U24116 (N_24116,N_22937,N_23746);
nand U24117 (N_24117,N_23002,N_23269);
or U24118 (N_24118,N_23000,N_23649);
or U24119 (N_24119,N_23141,N_23187);
nor U24120 (N_24120,N_23353,N_23769);
nor U24121 (N_24121,N_23468,N_23137);
xnor U24122 (N_24122,N_23799,N_23001);
and U24123 (N_24123,N_23903,N_23036);
xnor U24124 (N_24124,N_23229,N_23564);
xor U24125 (N_24125,N_23539,N_23594);
xor U24126 (N_24126,N_23990,N_22903);
or U24127 (N_24127,N_23170,N_23220);
and U24128 (N_24128,N_23336,N_23023);
nand U24129 (N_24129,N_23939,N_23287);
xnor U24130 (N_24130,N_23017,N_23261);
xnor U24131 (N_24131,N_23571,N_22945);
or U24132 (N_24132,N_23660,N_22883);
nand U24133 (N_24133,N_23267,N_22819);
and U24134 (N_24134,N_23583,N_23194);
and U24135 (N_24135,N_23254,N_23626);
or U24136 (N_24136,N_22872,N_23764);
nand U24137 (N_24137,N_23463,N_22994);
nand U24138 (N_24138,N_22830,N_23822);
nor U24139 (N_24139,N_23010,N_23724);
nand U24140 (N_24140,N_23604,N_23869);
xnor U24141 (N_24141,N_22931,N_23329);
nor U24142 (N_24142,N_23699,N_23569);
or U24143 (N_24143,N_23365,N_23585);
and U24144 (N_24144,N_23655,N_23414);
nand U24145 (N_24145,N_23887,N_23228);
nand U24146 (N_24146,N_23152,N_23345);
or U24147 (N_24147,N_23846,N_23148);
or U24148 (N_24148,N_23386,N_23629);
nand U24149 (N_24149,N_23196,N_23783);
nand U24150 (N_24150,N_23242,N_22803);
nand U24151 (N_24151,N_23005,N_22971);
nand U24152 (N_24152,N_23996,N_23909);
nand U24153 (N_24153,N_23798,N_23502);
and U24154 (N_24154,N_23081,N_22925);
nor U24155 (N_24155,N_23894,N_23631);
nor U24156 (N_24156,N_23421,N_23530);
and U24157 (N_24157,N_23716,N_23174);
and U24158 (N_24158,N_23082,N_23535);
or U24159 (N_24159,N_22896,N_23922);
and U24160 (N_24160,N_23452,N_23221);
xor U24161 (N_24161,N_22894,N_23366);
and U24162 (N_24162,N_23982,N_23153);
and U24163 (N_24163,N_23839,N_23630);
and U24164 (N_24164,N_23524,N_23738);
nand U24165 (N_24165,N_23734,N_23231);
nand U24166 (N_24166,N_23507,N_23086);
nand U24167 (N_24167,N_23740,N_23498);
and U24168 (N_24168,N_23973,N_23159);
or U24169 (N_24169,N_23505,N_23390);
or U24170 (N_24170,N_23035,N_23818);
nor U24171 (N_24171,N_23093,N_23685);
nand U24172 (N_24172,N_23047,N_23059);
nor U24173 (N_24173,N_23492,N_23928);
or U24174 (N_24174,N_23672,N_22936);
nand U24175 (N_24175,N_23009,N_23522);
or U24176 (N_24176,N_23709,N_23135);
nand U24177 (N_24177,N_23360,N_23006);
and U24178 (N_24178,N_23417,N_22828);
or U24179 (N_24179,N_23991,N_23462);
nor U24180 (N_24180,N_22866,N_23936);
and U24181 (N_24181,N_23282,N_23897);
or U24182 (N_24182,N_23259,N_22916);
and U24183 (N_24183,N_23579,N_23130);
nand U24184 (N_24184,N_22950,N_23520);
nand U24185 (N_24185,N_23727,N_23866);
xor U24186 (N_24186,N_22942,N_23389);
or U24187 (N_24187,N_23144,N_23968);
xor U24188 (N_24188,N_23646,N_22823);
and U24189 (N_24189,N_23156,N_23202);
nor U24190 (N_24190,N_22875,N_23702);
xor U24191 (N_24191,N_23959,N_23056);
or U24192 (N_24192,N_23620,N_23090);
nor U24193 (N_24193,N_23495,N_23429);
nor U24194 (N_24194,N_23458,N_23815);
or U24195 (N_24195,N_23257,N_22868);
or U24196 (N_24196,N_23444,N_23749);
nor U24197 (N_24197,N_23852,N_23833);
nand U24198 (N_24198,N_23033,N_23804);
nand U24199 (N_24199,N_23970,N_23120);
nor U24200 (N_24200,N_23847,N_23119);
or U24201 (N_24201,N_23711,N_23154);
xnor U24202 (N_24202,N_23280,N_23122);
xor U24203 (N_24203,N_22959,N_23929);
nor U24204 (N_24204,N_23067,N_23391);
xor U24205 (N_24205,N_23316,N_23298);
nand U24206 (N_24206,N_23895,N_23224);
or U24207 (N_24207,N_23434,N_23032);
or U24208 (N_24208,N_23193,N_23941);
and U24209 (N_24209,N_23476,N_23126);
xnor U24210 (N_24210,N_23568,N_23459);
nor U24211 (N_24211,N_23790,N_22963);
nor U24212 (N_24212,N_22999,N_23662);
xor U24213 (N_24213,N_23872,N_23245);
and U24214 (N_24214,N_23694,N_22834);
and U24215 (N_24215,N_23371,N_23383);
and U24216 (N_24216,N_23018,N_23488);
nand U24217 (N_24217,N_23576,N_23132);
nor U24218 (N_24218,N_22810,N_23713);
or U24219 (N_24219,N_23021,N_23639);
nor U24220 (N_24220,N_23561,N_22922);
nor U24221 (N_24221,N_22861,N_23055);
nand U24222 (N_24222,N_23258,N_23923);
or U24223 (N_24223,N_23937,N_23848);
xor U24224 (N_24224,N_23820,N_23641);
or U24225 (N_24225,N_23880,N_22879);
xor U24226 (N_24226,N_23946,N_23368);
or U24227 (N_24227,N_23378,N_23862);
or U24228 (N_24228,N_23310,N_22941);
nor U24229 (N_24229,N_22981,N_23858);
xnor U24230 (N_24230,N_23782,N_23200);
nor U24231 (N_24231,N_23447,N_23874);
and U24232 (N_24232,N_23098,N_23293);
xnor U24233 (N_24233,N_22876,N_22980);
and U24234 (N_24234,N_23735,N_23241);
nand U24235 (N_24235,N_22924,N_23664);
and U24236 (N_24236,N_23095,N_23819);
or U24237 (N_24237,N_22846,N_23262);
and U24238 (N_24238,N_22840,N_23644);
xnor U24239 (N_24239,N_23865,N_23134);
nor U24240 (N_24240,N_23363,N_23173);
or U24241 (N_24241,N_23687,N_23741);
nand U24242 (N_24242,N_23405,N_23558);
nand U24243 (N_24243,N_22954,N_23981);
xnor U24244 (N_24244,N_23654,N_23288);
and U24245 (N_24245,N_23905,N_23210);
and U24246 (N_24246,N_23342,N_23785);
nand U24247 (N_24247,N_23911,N_23404);
or U24248 (N_24248,N_23706,N_23250);
and U24249 (N_24249,N_23277,N_22807);
or U24250 (N_24250,N_23669,N_23966);
nor U24251 (N_24251,N_23999,N_22904);
nor U24252 (N_24252,N_23544,N_23657);
nand U24253 (N_24253,N_23623,N_23445);
or U24254 (N_24254,N_23893,N_23112);
xnor U24255 (N_24255,N_23070,N_23835);
nand U24256 (N_24256,N_23456,N_22928);
and U24257 (N_24257,N_23074,N_23533);
nor U24258 (N_24258,N_23489,N_23698);
nor U24259 (N_24259,N_22938,N_23092);
xor U24260 (N_24260,N_23089,N_23933);
nand U24261 (N_24261,N_23932,N_23155);
or U24262 (N_24262,N_22870,N_22949);
xor U24263 (N_24263,N_23169,N_23029);
and U24264 (N_24264,N_23163,N_23354);
or U24265 (N_24265,N_23038,N_23529);
nand U24266 (N_24266,N_23103,N_23305);
or U24267 (N_24267,N_23573,N_22910);
and U24268 (N_24268,N_23142,N_23235);
xnor U24269 (N_24269,N_23079,N_23906);
xnor U24270 (N_24270,N_23295,N_23123);
nand U24271 (N_24271,N_23256,N_23889);
xnor U24272 (N_24272,N_22974,N_23367);
and U24273 (N_24273,N_23061,N_22801);
nand U24274 (N_24274,N_23682,N_23403);
nand U24275 (N_24275,N_23695,N_23478);
and U24276 (N_24276,N_23538,N_23586);
nand U24277 (N_24277,N_23552,N_22998);
nor U24278 (N_24278,N_23546,N_23215);
and U24279 (N_24279,N_22878,N_23379);
xnor U24280 (N_24280,N_23322,N_23388);
and U24281 (N_24281,N_23692,N_22850);
nor U24282 (N_24282,N_22884,N_23612);
nor U24283 (N_24283,N_22893,N_23209);
and U24284 (N_24284,N_23251,N_23031);
nor U24285 (N_24285,N_23045,N_23940);
xor U24286 (N_24286,N_23472,N_23823);
nand U24287 (N_24287,N_23494,N_23395);
or U24288 (N_24288,N_23249,N_23745);
and U24289 (N_24289,N_23016,N_23113);
nor U24290 (N_24290,N_23598,N_23330);
nand U24291 (N_24291,N_23868,N_22906);
nor U24292 (N_24292,N_23904,N_22964);
nand U24293 (N_24293,N_23385,N_23222);
or U24294 (N_24294,N_23088,N_23285);
nand U24295 (N_24295,N_23656,N_22955);
or U24296 (N_24296,N_23962,N_23691);
xor U24297 (N_24297,N_23470,N_22824);
and U24298 (N_24298,N_23638,N_22845);
and U24299 (N_24299,N_23743,N_23763);
nand U24300 (N_24300,N_23506,N_23784);
and U24301 (N_24301,N_23286,N_22817);
nor U24302 (N_24302,N_23118,N_23493);
xnor U24303 (N_24303,N_23651,N_23992);
nand U24304 (N_24304,N_23677,N_23611);
or U24305 (N_24305,N_23607,N_23357);
and U24306 (N_24306,N_23239,N_23896);
or U24307 (N_24307,N_23615,N_23813);
nor U24308 (N_24308,N_23827,N_23150);
and U24309 (N_24309,N_23674,N_23128);
and U24310 (N_24310,N_23975,N_22809);
nor U24311 (N_24311,N_23545,N_23671);
nor U24312 (N_24312,N_23172,N_22886);
xor U24313 (N_24313,N_23854,N_23690);
or U24314 (N_24314,N_23274,N_23521);
and U24315 (N_24315,N_22920,N_22918);
nand U24316 (N_24316,N_23549,N_23308);
nor U24317 (N_24317,N_23913,N_23084);
and U24318 (N_24318,N_23957,N_23037);
xor U24319 (N_24319,N_23246,N_23328);
and U24320 (N_24320,N_22902,N_23760);
and U24321 (N_24321,N_23503,N_23272);
nand U24322 (N_24322,N_22851,N_23951);
nor U24323 (N_24323,N_22908,N_23185);
or U24324 (N_24324,N_23908,N_23451);
nand U24325 (N_24325,N_22993,N_23800);
nor U24326 (N_24326,N_23810,N_23750);
nor U24327 (N_24327,N_23838,N_23663);
xor U24328 (N_24328,N_23536,N_23730);
xnor U24329 (N_24329,N_23332,N_23901);
nor U24330 (N_24330,N_22890,N_23721);
nor U24331 (N_24331,N_22996,N_23464);
nand U24332 (N_24332,N_23197,N_23271);
nor U24333 (N_24333,N_23051,N_22976);
or U24334 (N_24334,N_23976,N_23824);
nor U24335 (N_24335,N_23460,N_23679);
or U24336 (N_24336,N_23343,N_23013);
nand U24337 (N_24337,N_23624,N_23175);
and U24338 (N_24338,N_23014,N_23515);
nor U24339 (N_24339,N_23176,N_23164);
or U24340 (N_24340,N_23284,N_23065);
nand U24341 (N_24341,N_23299,N_22827);
or U24342 (N_24342,N_23807,N_23039);
nor U24343 (N_24343,N_22989,N_22808);
xnor U24344 (N_24344,N_23780,N_23614);
or U24345 (N_24345,N_23877,N_23410);
and U24346 (N_24346,N_23581,N_22858);
xnor U24347 (N_24347,N_23723,N_23814);
and U24348 (N_24348,N_23504,N_23399);
nor U24349 (N_24349,N_23412,N_23279);
nor U24350 (N_24350,N_23349,N_22985);
nand U24351 (N_24351,N_23024,N_23436);
or U24352 (N_24352,N_23752,N_23560);
nand U24353 (N_24353,N_22946,N_23980);
or U24354 (N_24354,N_23610,N_23356);
and U24355 (N_24355,N_23348,N_22979);
nor U24356 (N_24356,N_23454,N_23717);
or U24357 (N_24357,N_23358,N_23914);
xnor U24358 (N_24358,N_23158,N_23844);
and U24359 (N_24359,N_22826,N_22991);
xnor U24360 (N_24360,N_23455,N_23778);
and U24361 (N_24361,N_22842,N_23370);
and U24362 (N_24362,N_23359,N_23240);
and U24363 (N_24363,N_23510,N_23313);
and U24364 (N_24364,N_23961,N_23860);
nor U24365 (N_24365,N_22831,N_23543);
xor U24366 (N_24366,N_23876,N_23177);
nand U24367 (N_24367,N_23411,N_23971);
or U24368 (N_24368,N_23145,N_23419);
xnor U24369 (N_24369,N_22970,N_23943);
nand U24370 (N_24370,N_23015,N_23479);
or U24371 (N_24371,N_23392,N_23593);
or U24372 (N_24372,N_22969,N_23645);
xor U24373 (N_24373,N_23739,N_23167);
nand U24374 (N_24374,N_23776,N_22881);
nand U24375 (N_24375,N_23772,N_23268);
xor U24376 (N_24376,N_23574,N_23183);
or U24377 (N_24377,N_23930,N_23863);
and U24378 (N_24378,N_22882,N_23281);
xor U24379 (N_24379,N_23563,N_23314);
nor U24380 (N_24380,N_23190,N_23634);
nor U24381 (N_24381,N_23040,N_23319);
and U24382 (N_24382,N_23987,N_23206);
xnor U24383 (N_24383,N_23548,N_23439);
or U24384 (N_24384,N_23105,N_23570);
or U24385 (N_24385,N_22921,N_23432);
and U24386 (N_24386,N_23248,N_23216);
and U24387 (N_24387,N_23580,N_22849);
or U24388 (N_24388,N_23797,N_23448);
nand U24389 (N_24389,N_23108,N_23374);
nor U24390 (N_24390,N_23661,N_23703);
xor U24391 (N_24391,N_23087,N_23290);
and U24392 (N_24392,N_23054,N_23449);
xnor U24393 (N_24393,N_22841,N_23668);
xnor U24394 (N_24394,N_22961,N_23578);
nand U24395 (N_24395,N_23066,N_23162);
xor U24396 (N_24396,N_22806,N_23707);
or U24397 (N_24397,N_23950,N_22978);
nand U24398 (N_24398,N_22832,N_23401);
nand U24399 (N_24399,N_23109,N_22844);
or U24400 (N_24400,N_23882,N_23442);
nand U24401 (N_24401,N_23166,N_23705);
or U24402 (N_24402,N_23335,N_22805);
nand U24403 (N_24403,N_23555,N_23283);
xnor U24404 (N_24404,N_23910,N_23097);
and U24405 (N_24405,N_23369,N_23337);
nor U24406 (N_24406,N_23101,N_23861);
xnor U24407 (N_24407,N_22859,N_23704);
and U24408 (N_24408,N_23441,N_23227);
nand U24409 (N_24409,N_23898,N_22952);
nand U24410 (N_24410,N_23019,N_23171);
and U24411 (N_24411,N_23963,N_23609);
nand U24412 (N_24412,N_23071,N_23253);
xor U24413 (N_24413,N_22947,N_23553);
or U24414 (N_24414,N_23766,N_23857);
nor U24415 (N_24415,N_23942,N_23541);
nand U24416 (N_24416,N_23255,N_23324);
nor U24417 (N_24417,N_23796,N_22835);
and U24418 (N_24418,N_23821,N_22847);
or U24419 (N_24419,N_22960,N_23603);
nand U24420 (N_24420,N_23192,N_22995);
and U24421 (N_24421,N_23920,N_23072);
xor U24422 (N_24422,N_23232,N_23069);
xor U24423 (N_24423,N_23075,N_23935);
nor U24424 (N_24424,N_23058,N_23540);
nand U24425 (N_24425,N_23346,N_23289);
and U24426 (N_24426,N_23931,N_23762);
and U24427 (N_24427,N_23060,N_23497);
nand U24428 (N_24428,N_23499,N_22951);
nand U24429 (N_24429,N_23380,N_22915);
or U24430 (N_24430,N_22853,N_23722);
nor U24431 (N_24431,N_23592,N_23073);
nor U24432 (N_24432,N_23836,N_23225);
and U24433 (N_24433,N_23531,N_23104);
and U24434 (N_24434,N_23890,N_23948);
or U24435 (N_24435,N_23309,N_23582);
nand U24436 (N_24436,N_23214,N_23595);
nor U24437 (N_24437,N_23756,N_23138);
and U24438 (N_24438,N_22874,N_23885);
nor U24439 (N_24439,N_23475,N_23978);
nor U24440 (N_24440,N_23554,N_23924);
nand U24441 (N_24441,N_23427,N_23781);
and U24442 (N_24442,N_23748,N_22848);
nor U24443 (N_24443,N_23921,N_22877);
nand U24444 (N_24444,N_23562,N_23509);
nor U24445 (N_24445,N_23376,N_22800);
nor U24446 (N_24446,N_23731,N_23292);
or U24447 (N_24447,N_23925,N_22869);
and U24448 (N_24448,N_23237,N_23046);
and U24449 (N_24449,N_23375,N_23556);
nor U24450 (N_24450,N_23372,N_23779);
nand U24451 (N_24451,N_23116,N_23387);
nor U24452 (N_24452,N_23967,N_23355);
or U24453 (N_24453,N_23008,N_23026);
xnor U24454 (N_24454,N_22891,N_23621);
nor U24455 (N_24455,N_23806,N_23334);
xor U24456 (N_24456,N_23787,N_23157);
xnor U24457 (N_24457,N_23466,N_23684);
xnor U24458 (N_24458,N_23718,N_23117);
and U24459 (N_24459,N_23652,N_23243);
nor U24460 (N_24460,N_23643,N_23057);
and U24461 (N_24461,N_23767,N_22977);
nor U24462 (N_24462,N_22957,N_23742);
and U24463 (N_24463,N_22816,N_23022);
xor U24464 (N_24464,N_23003,N_23491);
or U24465 (N_24465,N_23400,N_23180);
or U24466 (N_24466,N_23302,N_23907);
or U24467 (N_24467,N_23178,N_23147);
nor U24468 (N_24468,N_22873,N_23426);
nand U24469 (N_24469,N_22962,N_23076);
nor U24470 (N_24470,N_23916,N_23217);
and U24471 (N_24471,N_23688,N_23758);
nand U24472 (N_24472,N_22923,N_23339);
nor U24473 (N_24473,N_23927,N_22862);
nor U24474 (N_24474,N_23317,N_23077);
or U24475 (N_24475,N_22855,N_22965);
xnor U24476 (N_24476,N_23658,N_23418);
nand U24477 (N_24477,N_23465,N_23842);
nor U24478 (N_24478,N_23774,N_23841);
nor U24479 (N_24479,N_23291,N_22967);
or U24480 (N_24480,N_23636,N_23761);
nor U24481 (N_24481,N_23213,N_22854);
and U24482 (N_24482,N_23511,N_22899);
nand U24483 (N_24483,N_23757,N_23428);
nand U24484 (N_24484,N_22856,N_23627);
xor U24485 (N_24485,N_23828,N_23467);
and U24486 (N_24486,N_23572,N_22909);
and U24487 (N_24487,N_23816,N_22838);
and U24488 (N_24488,N_23883,N_23048);
xnor U24489 (N_24489,N_23315,N_23301);
nor U24490 (N_24490,N_22865,N_23884);
nand U24491 (N_24491,N_23394,N_23115);
and U24492 (N_24492,N_23986,N_22863);
and U24493 (N_24493,N_23030,N_22926);
or U24494 (N_24494,N_23725,N_23673);
nor U24495 (N_24495,N_23450,N_23437);
and U24496 (N_24496,N_22992,N_23300);
xnor U24497 (N_24497,N_23398,N_23133);
nor U24498 (N_24498,N_23028,N_22836);
and U24499 (N_24499,N_23361,N_23988);
nand U24500 (N_24500,N_23094,N_23775);
nor U24501 (N_24501,N_23728,N_23871);
nor U24502 (N_24502,N_23792,N_23477);
and U24503 (N_24503,N_23864,N_23888);
nand U24504 (N_24504,N_23266,N_23182);
or U24505 (N_24505,N_23675,N_22929);
and U24506 (N_24506,N_23855,N_23640);
or U24507 (N_24507,N_23853,N_23984);
nor U24508 (N_24508,N_23179,N_22914);
or U24509 (N_24509,N_23902,N_23063);
nand U24510 (N_24510,N_23812,N_23195);
nand U24511 (N_24511,N_22822,N_23754);
nor U24512 (N_24512,N_22975,N_22802);
nand U24513 (N_24513,N_22912,N_22814);
xor U24514 (N_24514,N_23362,N_23826);
nand U24515 (N_24515,N_23605,N_23482);
nor U24516 (N_24516,N_23733,N_23294);
xnor U24517 (N_24517,N_22986,N_23020);
and U24518 (N_24518,N_23637,N_23994);
or U24519 (N_24519,N_23701,N_23205);
or U24520 (N_24520,N_22966,N_23080);
nor U24521 (N_24521,N_22984,N_23759);
xnor U24522 (N_24522,N_23007,N_23233);
and U24523 (N_24523,N_23945,N_23424);
and U24524 (N_24524,N_22933,N_22972);
nand U24525 (N_24525,N_23736,N_23260);
nand U24526 (N_24526,N_23514,N_23457);
and U24527 (N_24527,N_23341,N_22911);
xnor U24528 (N_24528,N_23944,N_23496);
xnor U24529 (N_24529,N_23408,N_23525);
or U24530 (N_24530,N_23802,N_23972);
and U24531 (N_24531,N_23900,N_23203);
xnor U24532 (N_24532,N_23484,N_23347);
nor U24533 (N_24533,N_23471,N_23926);
or U24534 (N_24534,N_23559,N_23513);
nor U24535 (N_24535,N_23099,N_23938);
xor U24536 (N_24536,N_23107,N_23715);
and U24537 (N_24537,N_22973,N_23584);
or U24538 (N_24538,N_23875,N_23034);
nor U24539 (N_24539,N_23325,N_23856);
nor U24540 (N_24540,N_23714,N_23110);
nand U24541 (N_24541,N_22919,N_23665);
nand U24542 (N_24542,N_23616,N_23934);
xnor U24543 (N_24543,N_23486,N_22897);
or U24544 (N_24544,N_23700,N_23409);
nor U24545 (N_24545,N_22983,N_22812);
nor U24546 (N_24546,N_23867,N_23532);
and U24547 (N_24547,N_23238,N_23697);
xnor U24548 (N_24548,N_23512,N_23870);
or U24549 (N_24549,N_23519,N_23278);
or U24550 (N_24550,N_23160,N_23199);
and U24551 (N_24551,N_23053,N_22852);
nand U24552 (N_24552,N_23608,N_23186);
xnor U24553 (N_24553,N_23989,N_23845);
and U24554 (N_24554,N_23918,N_23373);
xor U24555 (N_24555,N_23483,N_23161);
nand U24556 (N_24556,N_23318,N_23083);
and U24557 (N_24557,N_23676,N_23667);
or U24558 (N_24558,N_23912,N_23590);
and U24559 (N_24559,N_22913,N_23350);
nor U24560 (N_24560,N_23181,N_23096);
and U24561 (N_24561,N_23788,N_23947);
and U24562 (N_24562,N_23600,N_23191);
or U24563 (N_24563,N_23995,N_23327);
nor U24564 (N_24564,N_23881,N_22839);
and U24565 (N_24565,N_23805,N_23501);
or U24566 (N_24566,N_23396,N_23131);
xor U24567 (N_24567,N_23344,N_23919);
nand U24568 (N_24568,N_23413,N_23381);
xnor U24569 (N_24569,N_23647,N_23211);
nand U24570 (N_24570,N_23751,N_23406);
nand U24571 (N_24571,N_23830,N_23831);
xor U24572 (N_24572,N_23547,N_23415);
xor U24573 (N_24573,N_23628,N_23352);
nor U24574 (N_24574,N_23143,N_23591);
or U24575 (N_24575,N_23964,N_23648);
and U24576 (N_24576,N_23236,N_22825);
nor U24577 (N_24577,N_23683,N_23625);
nand U24578 (N_24578,N_22887,N_23297);
nor U24579 (N_24579,N_23481,N_23597);
xnor U24580 (N_24580,N_23565,N_22953);
nor U24581 (N_24581,N_23878,N_23960);
nand U24582 (N_24582,N_23425,N_23050);
nor U24583 (N_24583,N_23840,N_23025);
or U24584 (N_24584,N_23998,N_23364);
nand U24585 (N_24585,N_23433,N_23786);
xor U24586 (N_24586,N_23997,N_23320);
nand U24587 (N_24587,N_23226,N_23526);
or U24588 (N_24588,N_23832,N_23954);
and U24589 (N_24589,N_23843,N_22820);
nor U24590 (N_24590,N_23744,N_23125);
and U24591 (N_24591,N_23837,N_22934);
xnor U24592 (N_24592,N_23642,N_23899);
xnor U24593 (N_24593,N_23789,N_23207);
and U24594 (N_24594,N_23729,N_23264);
and U24595 (N_24595,N_22880,N_23567);
xnor U24596 (N_24596,N_22939,N_23435);
or U24597 (N_24597,N_22821,N_23601);
nand U24598 (N_24598,N_22901,N_23599);
nor U24599 (N_24599,N_22987,N_23340);
and U24600 (N_24600,N_23956,N_22829);
and U24601 (N_24601,N_22938,N_22832);
or U24602 (N_24602,N_22933,N_23441);
or U24603 (N_24603,N_22954,N_22963);
and U24604 (N_24604,N_23369,N_23841);
or U24605 (N_24605,N_23541,N_23416);
and U24606 (N_24606,N_22905,N_22977);
nor U24607 (N_24607,N_23323,N_23173);
or U24608 (N_24608,N_23463,N_23352);
nor U24609 (N_24609,N_22997,N_23093);
nand U24610 (N_24610,N_23548,N_22904);
nor U24611 (N_24611,N_22866,N_22919);
xnor U24612 (N_24612,N_23450,N_23473);
and U24613 (N_24613,N_23312,N_23515);
xor U24614 (N_24614,N_22820,N_23728);
and U24615 (N_24615,N_23138,N_23591);
xor U24616 (N_24616,N_23272,N_23668);
and U24617 (N_24617,N_23859,N_23987);
xor U24618 (N_24618,N_23238,N_23408);
xor U24619 (N_24619,N_23514,N_23116);
and U24620 (N_24620,N_22908,N_23754);
and U24621 (N_24621,N_22895,N_23419);
and U24622 (N_24622,N_23783,N_23142);
or U24623 (N_24623,N_23021,N_23558);
and U24624 (N_24624,N_23162,N_23301);
and U24625 (N_24625,N_23435,N_23781);
nor U24626 (N_24626,N_23574,N_23518);
nand U24627 (N_24627,N_23354,N_23107);
nand U24628 (N_24628,N_23216,N_23116);
or U24629 (N_24629,N_22820,N_23136);
or U24630 (N_24630,N_23630,N_23339);
xor U24631 (N_24631,N_23025,N_22819);
or U24632 (N_24632,N_23281,N_23555);
or U24633 (N_24633,N_23746,N_23472);
xnor U24634 (N_24634,N_23407,N_23108);
nor U24635 (N_24635,N_23863,N_23389);
nor U24636 (N_24636,N_23139,N_23650);
and U24637 (N_24637,N_23967,N_22855);
or U24638 (N_24638,N_23802,N_23292);
nor U24639 (N_24639,N_23546,N_23417);
and U24640 (N_24640,N_22945,N_23308);
and U24641 (N_24641,N_23045,N_23173);
nand U24642 (N_24642,N_23607,N_23842);
xnor U24643 (N_24643,N_23136,N_23540);
xor U24644 (N_24644,N_23256,N_23563);
and U24645 (N_24645,N_22871,N_23177);
or U24646 (N_24646,N_22932,N_23251);
nand U24647 (N_24647,N_23229,N_23253);
and U24648 (N_24648,N_23888,N_23366);
and U24649 (N_24649,N_23636,N_23385);
nor U24650 (N_24650,N_23609,N_23600);
nor U24651 (N_24651,N_23519,N_23025);
and U24652 (N_24652,N_23709,N_23717);
xor U24653 (N_24653,N_23453,N_23590);
or U24654 (N_24654,N_22884,N_23650);
nand U24655 (N_24655,N_23418,N_22944);
and U24656 (N_24656,N_23390,N_23339);
and U24657 (N_24657,N_23988,N_23754);
nor U24658 (N_24658,N_23361,N_23076);
or U24659 (N_24659,N_22845,N_22895);
or U24660 (N_24660,N_23908,N_23619);
xor U24661 (N_24661,N_23791,N_23569);
or U24662 (N_24662,N_22942,N_22822);
and U24663 (N_24663,N_23133,N_23936);
nor U24664 (N_24664,N_23142,N_23810);
nand U24665 (N_24665,N_23522,N_23092);
xor U24666 (N_24666,N_23406,N_22916);
or U24667 (N_24667,N_23098,N_23552);
nor U24668 (N_24668,N_23955,N_22826);
and U24669 (N_24669,N_23966,N_22952);
xnor U24670 (N_24670,N_23409,N_23174);
xor U24671 (N_24671,N_23143,N_23663);
xnor U24672 (N_24672,N_23872,N_22915);
nor U24673 (N_24673,N_23457,N_23319);
or U24674 (N_24674,N_23256,N_23040);
and U24675 (N_24675,N_23264,N_23847);
and U24676 (N_24676,N_23752,N_23706);
or U24677 (N_24677,N_23762,N_22940);
xor U24678 (N_24678,N_23636,N_23697);
xor U24679 (N_24679,N_23547,N_23260);
and U24680 (N_24680,N_22846,N_22849);
xnor U24681 (N_24681,N_23494,N_23229);
nand U24682 (N_24682,N_23124,N_23716);
nand U24683 (N_24683,N_23964,N_22845);
nor U24684 (N_24684,N_23101,N_22909);
or U24685 (N_24685,N_23194,N_23056);
nor U24686 (N_24686,N_23001,N_23175);
nand U24687 (N_24687,N_23757,N_23892);
or U24688 (N_24688,N_23252,N_23676);
xor U24689 (N_24689,N_23421,N_22926);
or U24690 (N_24690,N_23156,N_23343);
and U24691 (N_24691,N_22821,N_23509);
or U24692 (N_24692,N_23821,N_23632);
xor U24693 (N_24693,N_23940,N_23521);
and U24694 (N_24694,N_23248,N_22935);
or U24695 (N_24695,N_23189,N_23397);
xor U24696 (N_24696,N_23536,N_23418);
and U24697 (N_24697,N_23823,N_23036);
xnor U24698 (N_24698,N_23620,N_23281);
nand U24699 (N_24699,N_23949,N_23417);
and U24700 (N_24700,N_23726,N_23312);
or U24701 (N_24701,N_23287,N_23930);
and U24702 (N_24702,N_23123,N_23166);
nand U24703 (N_24703,N_23154,N_23271);
nor U24704 (N_24704,N_23181,N_22904);
nand U24705 (N_24705,N_22947,N_23234);
and U24706 (N_24706,N_23509,N_23221);
or U24707 (N_24707,N_23798,N_23729);
and U24708 (N_24708,N_23587,N_23903);
nand U24709 (N_24709,N_23707,N_23359);
nor U24710 (N_24710,N_23202,N_22803);
nand U24711 (N_24711,N_22947,N_23230);
nor U24712 (N_24712,N_23144,N_22834);
xor U24713 (N_24713,N_22857,N_23054);
or U24714 (N_24714,N_23320,N_23261);
nor U24715 (N_24715,N_22808,N_23329);
or U24716 (N_24716,N_22820,N_23334);
and U24717 (N_24717,N_23521,N_23863);
nand U24718 (N_24718,N_23238,N_23625);
xnor U24719 (N_24719,N_23746,N_23848);
nand U24720 (N_24720,N_22931,N_22971);
nor U24721 (N_24721,N_23038,N_23520);
xor U24722 (N_24722,N_23414,N_23026);
and U24723 (N_24723,N_22927,N_23194);
nor U24724 (N_24724,N_23932,N_23328);
xor U24725 (N_24725,N_23353,N_23882);
and U24726 (N_24726,N_23756,N_23095);
xnor U24727 (N_24727,N_23531,N_23905);
or U24728 (N_24728,N_23567,N_23632);
xor U24729 (N_24729,N_23395,N_23908);
xnor U24730 (N_24730,N_23418,N_23886);
nor U24731 (N_24731,N_23921,N_23908);
nand U24732 (N_24732,N_23889,N_23373);
and U24733 (N_24733,N_23805,N_22991);
nand U24734 (N_24734,N_23994,N_22925);
or U24735 (N_24735,N_23886,N_23080);
and U24736 (N_24736,N_23737,N_22923);
nor U24737 (N_24737,N_23227,N_22920);
nand U24738 (N_24738,N_23526,N_23471);
xor U24739 (N_24739,N_22850,N_23125);
nand U24740 (N_24740,N_23031,N_23801);
xnor U24741 (N_24741,N_23369,N_23679);
nand U24742 (N_24742,N_22868,N_23149);
nand U24743 (N_24743,N_22880,N_23102);
nand U24744 (N_24744,N_23179,N_23249);
nor U24745 (N_24745,N_23007,N_23114);
nor U24746 (N_24746,N_22827,N_23971);
nor U24747 (N_24747,N_23490,N_23442);
xnor U24748 (N_24748,N_23067,N_22945);
nand U24749 (N_24749,N_23944,N_23866);
nand U24750 (N_24750,N_23972,N_23866);
nor U24751 (N_24751,N_23917,N_23943);
or U24752 (N_24752,N_23647,N_22915);
xor U24753 (N_24753,N_22895,N_23295);
nand U24754 (N_24754,N_23404,N_23926);
xor U24755 (N_24755,N_23878,N_23449);
nand U24756 (N_24756,N_23882,N_23481);
nand U24757 (N_24757,N_23356,N_23062);
nor U24758 (N_24758,N_22952,N_23761);
or U24759 (N_24759,N_23307,N_23943);
or U24760 (N_24760,N_23806,N_23824);
nor U24761 (N_24761,N_22841,N_23809);
xnor U24762 (N_24762,N_23847,N_23370);
and U24763 (N_24763,N_22826,N_22951);
and U24764 (N_24764,N_23349,N_23326);
nor U24765 (N_24765,N_23823,N_23301);
nor U24766 (N_24766,N_23259,N_22882);
or U24767 (N_24767,N_23235,N_23628);
nand U24768 (N_24768,N_23365,N_23256);
and U24769 (N_24769,N_23623,N_23069);
nand U24770 (N_24770,N_23942,N_23173);
nor U24771 (N_24771,N_22955,N_23688);
xor U24772 (N_24772,N_22806,N_23561);
xor U24773 (N_24773,N_23422,N_23314);
nand U24774 (N_24774,N_23848,N_23918);
or U24775 (N_24775,N_23258,N_23879);
nor U24776 (N_24776,N_23868,N_23746);
nor U24777 (N_24777,N_23491,N_22943);
xor U24778 (N_24778,N_23530,N_23938);
or U24779 (N_24779,N_23098,N_23776);
nor U24780 (N_24780,N_23608,N_23311);
nand U24781 (N_24781,N_23059,N_23541);
or U24782 (N_24782,N_23326,N_23352);
nor U24783 (N_24783,N_23667,N_23768);
or U24784 (N_24784,N_23371,N_23038);
and U24785 (N_24785,N_23041,N_23101);
nor U24786 (N_24786,N_23314,N_22887);
nand U24787 (N_24787,N_22898,N_23840);
nand U24788 (N_24788,N_23177,N_23762);
nand U24789 (N_24789,N_22826,N_23249);
and U24790 (N_24790,N_23909,N_23442);
or U24791 (N_24791,N_23853,N_23432);
or U24792 (N_24792,N_23916,N_23976);
or U24793 (N_24793,N_23389,N_23255);
xnor U24794 (N_24794,N_23281,N_23908);
xor U24795 (N_24795,N_22824,N_23425);
nand U24796 (N_24796,N_23136,N_23489);
nand U24797 (N_24797,N_23456,N_22848);
nand U24798 (N_24798,N_23319,N_23326);
nand U24799 (N_24799,N_23934,N_23374);
xor U24800 (N_24800,N_23683,N_23094);
nand U24801 (N_24801,N_23216,N_23387);
or U24802 (N_24802,N_23923,N_23295);
nand U24803 (N_24803,N_23192,N_23763);
nor U24804 (N_24804,N_23973,N_22836);
xnor U24805 (N_24805,N_23078,N_23104);
nor U24806 (N_24806,N_23721,N_23885);
and U24807 (N_24807,N_23829,N_23996);
or U24808 (N_24808,N_23242,N_22962);
nand U24809 (N_24809,N_22959,N_23204);
xor U24810 (N_24810,N_23903,N_22940);
xor U24811 (N_24811,N_23192,N_23163);
and U24812 (N_24812,N_23320,N_23024);
or U24813 (N_24813,N_23135,N_23707);
or U24814 (N_24814,N_23596,N_23901);
nor U24815 (N_24815,N_23174,N_22817);
nor U24816 (N_24816,N_23460,N_23515);
nand U24817 (N_24817,N_23336,N_23112);
or U24818 (N_24818,N_23102,N_23342);
nor U24819 (N_24819,N_22916,N_23044);
or U24820 (N_24820,N_23327,N_23218);
xor U24821 (N_24821,N_23182,N_23074);
nor U24822 (N_24822,N_23140,N_23052);
nand U24823 (N_24823,N_22921,N_22859);
xnor U24824 (N_24824,N_23950,N_23753);
nor U24825 (N_24825,N_23271,N_23975);
xnor U24826 (N_24826,N_22910,N_23009);
or U24827 (N_24827,N_23036,N_23467);
nand U24828 (N_24828,N_23620,N_22929);
xor U24829 (N_24829,N_23588,N_23604);
and U24830 (N_24830,N_23436,N_23715);
xor U24831 (N_24831,N_23180,N_23411);
or U24832 (N_24832,N_23691,N_23161);
xor U24833 (N_24833,N_23889,N_23755);
nand U24834 (N_24834,N_22954,N_23652);
nand U24835 (N_24835,N_22919,N_23371);
nand U24836 (N_24836,N_23673,N_23767);
nand U24837 (N_24837,N_23095,N_22902);
nor U24838 (N_24838,N_23360,N_23974);
or U24839 (N_24839,N_23118,N_22981);
nor U24840 (N_24840,N_23885,N_22860);
or U24841 (N_24841,N_23860,N_23084);
nor U24842 (N_24842,N_23008,N_23711);
xnor U24843 (N_24843,N_22983,N_23057);
or U24844 (N_24844,N_23600,N_23618);
or U24845 (N_24845,N_22886,N_22957);
xor U24846 (N_24846,N_22916,N_22900);
nor U24847 (N_24847,N_22978,N_23041);
and U24848 (N_24848,N_23938,N_23903);
or U24849 (N_24849,N_22819,N_23225);
and U24850 (N_24850,N_23394,N_22871);
or U24851 (N_24851,N_23547,N_22855);
xor U24852 (N_24852,N_23782,N_23692);
nor U24853 (N_24853,N_23658,N_22966);
xnor U24854 (N_24854,N_23830,N_23722);
xnor U24855 (N_24855,N_23773,N_23969);
or U24856 (N_24856,N_23699,N_23941);
or U24857 (N_24857,N_23640,N_23496);
nand U24858 (N_24858,N_23217,N_23958);
nand U24859 (N_24859,N_23030,N_23455);
and U24860 (N_24860,N_23192,N_23969);
xor U24861 (N_24861,N_23162,N_23358);
nand U24862 (N_24862,N_23082,N_23311);
nor U24863 (N_24863,N_22814,N_23992);
xnor U24864 (N_24864,N_23855,N_23429);
xnor U24865 (N_24865,N_23838,N_23165);
nand U24866 (N_24866,N_23713,N_23594);
nand U24867 (N_24867,N_23394,N_23418);
xnor U24868 (N_24868,N_22935,N_23693);
and U24869 (N_24869,N_23173,N_23890);
nor U24870 (N_24870,N_23890,N_23351);
or U24871 (N_24871,N_23558,N_23406);
nor U24872 (N_24872,N_23193,N_23295);
xor U24873 (N_24873,N_23397,N_22872);
and U24874 (N_24874,N_23933,N_23613);
and U24875 (N_24875,N_23472,N_23685);
nor U24876 (N_24876,N_23102,N_22808);
or U24877 (N_24877,N_23755,N_23986);
or U24878 (N_24878,N_23432,N_23490);
xor U24879 (N_24879,N_23952,N_23457);
xor U24880 (N_24880,N_23966,N_23558);
nor U24881 (N_24881,N_23653,N_23153);
nand U24882 (N_24882,N_23562,N_23738);
nand U24883 (N_24883,N_23498,N_23009);
nand U24884 (N_24884,N_23375,N_23250);
or U24885 (N_24885,N_23354,N_23266);
nand U24886 (N_24886,N_23088,N_23634);
or U24887 (N_24887,N_23110,N_22844);
or U24888 (N_24888,N_23168,N_22839);
and U24889 (N_24889,N_23008,N_23298);
nand U24890 (N_24890,N_23073,N_23467);
xnor U24891 (N_24891,N_23046,N_23703);
xnor U24892 (N_24892,N_23431,N_23846);
nand U24893 (N_24893,N_23559,N_22803);
xor U24894 (N_24894,N_23874,N_22879);
or U24895 (N_24895,N_22902,N_22891);
nor U24896 (N_24896,N_23441,N_23699);
nor U24897 (N_24897,N_23319,N_23378);
and U24898 (N_24898,N_22924,N_23538);
or U24899 (N_24899,N_23305,N_23638);
or U24900 (N_24900,N_23973,N_23865);
and U24901 (N_24901,N_23048,N_23726);
nand U24902 (N_24902,N_23576,N_22914);
nor U24903 (N_24903,N_22965,N_23240);
nor U24904 (N_24904,N_23640,N_23805);
nand U24905 (N_24905,N_23904,N_23211);
xor U24906 (N_24906,N_23365,N_22869);
or U24907 (N_24907,N_23913,N_23390);
and U24908 (N_24908,N_23514,N_22925);
and U24909 (N_24909,N_22847,N_22868);
xnor U24910 (N_24910,N_23469,N_23855);
nor U24911 (N_24911,N_23263,N_23087);
nor U24912 (N_24912,N_23961,N_23743);
xnor U24913 (N_24913,N_23017,N_23211);
nand U24914 (N_24914,N_22851,N_23339);
nor U24915 (N_24915,N_23855,N_23737);
or U24916 (N_24916,N_23490,N_23904);
nand U24917 (N_24917,N_23058,N_22939);
and U24918 (N_24918,N_23733,N_22960);
xnor U24919 (N_24919,N_23179,N_23387);
nor U24920 (N_24920,N_23478,N_23967);
or U24921 (N_24921,N_23332,N_23635);
or U24922 (N_24922,N_23227,N_23798);
xnor U24923 (N_24923,N_22804,N_23761);
nand U24924 (N_24924,N_23750,N_23368);
xor U24925 (N_24925,N_23283,N_23605);
nor U24926 (N_24926,N_23967,N_23435);
and U24927 (N_24927,N_23667,N_23123);
nor U24928 (N_24928,N_23054,N_22959);
nand U24929 (N_24929,N_23819,N_23655);
or U24930 (N_24930,N_23486,N_23748);
or U24931 (N_24931,N_23998,N_23682);
or U24932 (N_24932,N_22896,N_23288);
or U24933 (N_24933,N_23671,N_23586);
xnor U24934 (N_24934,N_23572,N_23118);
or U24935 (N_24935,N_23913,N_23414);
or U24936 (N_24936,N_23642,N_23674);
or U24937 (N_24937,N_23860,N_23511);
xnor U24938 (N_24938,N_23578,N_23407);
or U24939 (N_24939,N_22997,N_23778);
or U24940 (N_24940,N_23175,N_23194);
and U24941 (N_24941,N_23596,N_23985);
nor U24942 (N_24942,N_22854,N_23025);
and U24943 (N_24943,N_23711,N_23347);
and U24944 (N_24944,N_23405,N_23846);
or U24945 (N_24945,N_23018,N_23440);
and U24946 (N_24946,N_23825,N_23304);
and U24947 (N_24947,N_23350,N_23368);
nand U24948 (N_24948,N_23161,N_23862);
nor U24949 (N_24949,N_23826,N_23687);
or U24950 (N_24950,N_23055,N_23791);
nand U24951 (N_24951,N_23693,N_23148);
xnor U24952 (N_24952,N_23696,N_23949);
and U24953 (N_24953,N_23646,N_23199);
and U24954 (N_24954,N_23438,N_22822);
nand U24955 (N_24955,N_23133,N_23441);
or U24956 (N_24956,N_23802,N_22960);
nand U24957 (N_24957,N_23570,N_23594);
or U24958 (N_24958,N_23626,N_23538);
xnor U24959 (N_24959,N_23445,N_23650);
and U24960 (N_24960,N_23080,N_22926);
nand U24961 (N_24961,N_23784,N_23202);
or U24962 (N_24962,N_23855,N_22884);
and U24963 (N_24963,N_22823,N_22856);
or U24964 (N_24964,N_23557,N_23568);
nor U24965 (N_24965,N_23936,N_23980);
and U24966 (N_24966,N_23300,N_23006);
xnor U24967 (N_24967,N_23047,N_23001);
or U24968 (N_24968,N_23199,N_23424);
nand U24969 (N_24969,N_23810,N_23840);
xor U24970 (N_24970,N_23136,N_23518);
nor U24971 (N_24971,N_23845,N_22957);
nand U24972 (N_24972,N_23696,N_23836);
nand U24973 (N_24973,N_22897,N_22903);
nand U24974 (N_24974,N_23406,N_23888);
or U24975 (N_24975,N_23208,N_23630);
nand U24976 (N_24976,N_23838,N_23835);
or U24977 (N_24977,N_22926,N_23649);
xnor U24978 (N_24978,N_23655,N_23067);
or U24979 (N_24979,N_23107,N_23969);
nor U24980 (N_24980,N_23003,N_23904);
nor U24981 (N_24981,N_22863,N_23718);
and U24982 (N_24982,N_23809,N_23615);
nor U24983 (N_24983,N_23849,N_22818);
nand U24984 (N_24984,N_22851,N_23270);
or U24985 (N_24985,N_23661,N_23494);
or U24986 (N_24986,N_23970,N_22886);
xnor U24987 (N_24987,N_22970,N_22960);
nor U24988 (N_24988,N_23445,N_23612);
and U24989 (N_24989,N_23165,N_23896);
and U24990 (N_24990,N_23947,N_23114);
nor U24991 (N_24991,N_23695,N_23915);
nand U24992 (N_24992,N_23782,N_23196);
nand U24993 (N_24993,N_23787,N_23017);
nand U24994 (N_24994,N_23096,N_23412);
or U24995 (N_24995,N_23937,N_23454);
xnor U24996 (N_24996,N_23659,N_23821);
nand U24997 (N_24997,N_23042,N_23918);
and U24998 (N_24998,N_23860,N_23766);
xor U24999 (N_24999,N_23979,N_23381);
xor U25000 (N_25000,N_23581,N_23784);
xor U25001 (N_25001,N_23505,N_23933);
nand U25002 (N_25002,N_23369,N_23903);
and U25003 (N_25003,N_23571,N_23608);
nor U25004 (N_25004,N_23685,N_23918);
nor U25005 (N_25005,N_23187,N_23276);
or U25006 (N_25006,N_23482,N_23442);
xnor U25007 (N_25007,N_23485,N_23222);
nor U25008 (N_25008,N_23359,N_23859);
and U25009 (N_25009,N_23217,N_23570);
and U25010 (N_25010,N_22835,N_23472);
nand U25011 (N_25011,N_23456,N_22806);
or U25012 (N_25012,N_23582,N_23166);
nand U25013 (N_25013,N_22814,N_22954);
nor U25014 (N_25014,N_23591,N_22870);
nor U25015 (N_25015,N_22894,N_22860);
nor U25016 (N_25016,N_23909,N_23270);
nand U25017 (N_25017,N_23530,N_23745);
nand U25018 (N_25018,N_22932,N_23651);
nand U25019 (N_25019,N_23637,N_23323);
nor U25020 (N_25020,N_23932,N_23557);
xnor U25021 (N_25021,N_23901,N_23156);
and U25022 (N_25022,N_22936,N_23846);
nor U25023 (N_25023,N_23771,N_23433);
and U25024 (N_25024,N_23455,N_23825);
nand U25025 (N_25025,N_22903,N_23780);
nor U25026 (N_25026,N_23798,N_23925);
nor U25027 (N_25027,N_23315,N_23295);
and U25028 (N_25028,N_23437,N_23660);
nand U25029 (N_25029,N_23738,N_23186);
nor U25030 (N_25030,N_23980,N_23801);
nand U25031 (N_25031,N_23055,N_23374);
or U25032 (N_25032,N_23810,N_22952);
and U25033 (N_25033,N_23139,N_23870);
nor U25034 (N_25034,N_23621,N_23863);
nand U25035 (N_25035,N_23304,N_23842);
nor U25036 (N_25036,N_22810,N_23620);
or U25037 (N_25037,N_23916,N_23424);
or U25038 (N_25038,N_23351,N_22973);
or U25039 (N_25039,N_23870,N_23208);
and U25040 (N_25040,N_23992,N_23893);
or U25041 (N_25041,N_23105,N_23772);
nor U25042 (N_25042,N_23507,N_23375);
or U25043 (N_25043,N_23910,N_23110);
nor U25044 (N_25044,N_22809,N_23789);
or U25045 (N_25045,N_23067,N_23018);
and U25046 (N_25046,N_22960,N_23431);
and U25047 (N_25047,N_23529,N_23882);
xnor U25048 (N_25048,N_23416,N_23251);
or U25049 (N_25049,N_23831,N_23625);
xnor U25050 (N_25050,N_23111,N_23879);
nor U25051 (N_25051,N_22893,N_23422);
nor U25052 (N_25052,N_23502,N_23136);
xor U25053 (N_25053,N_23024,N_23397);
nor U25054 (N_25054,N_23758,N_23712);
nand U25055 (N_25055,N_23858,N_22892);
xor U25056 (N_25056,N_23730,N_23138);
xnor U25057 (N_25057,N_23921,N_22834);
xor U25058 (N_25058,N_23676,N_23405);
nor U25059 (N_25059,N_23981,N_23101);
nand U25060 (N_25060,N_23878,N_23796);
xnor U25061 (N_25061,N_22930,N_23472);
or U25062 (N_25062,N_23120,N_23389);
and U25063 (N_25063,N_23284,N_23990);
nand U25064 (N_25064,N_23831,N_23396);
or U25065 (N_25065,N_23401,N_23998);
nand U25066 (N_25066,N_23771,N_23373);
or U25067 (N_25067,N_23822,N_23367);
and U25068 (N_25068,N_23958,N_23111);
nor U25069 (N_25069,N_23544,N_22823);
xnor U25070 (N_25070,N_23277,N_23114);
nor U25071 (N_25071,N_23356,N_23393);
or U25072 (N_25072,N_23596,N_23567);
and U25073 (N_25073,N_22884,N_22890);
and U25074 (N_25074,N_23677,N_23213);
or U25075 (N_25075,N_23207,N_23227);
nor U25076 (N_25076,N_23356,N_23487);
nor U25077 (N_25077,N_23826,N_23388);
nor U25078 (N_25078,N_23482,N_22900);
or U25079 (N_25079,N_23582,N_22815);
and U25080 (N_25080,N_23045,N_23769);
nor U25081 (N_25081,N_23244,N_23527);
xnor U25082 (N_25082,N_23988,N_22992);
nand U25083 (N_25083,N_23423,N_23035);
xnor U25084 (N_25084,N_23831,N_22857);
nand U25085 (N_25085,N_23859,N_22932);
xor U25086 (N_25086,N_23668,N_22860);
nor U25087 (N_25087,N_23777,N_23584);
xor U25088 (N_25088,N_22892,N_23906);
nor U25089 (N_25089,N_22962,N_23020);
or U25090 (N_25090,N_23010,N_23874);
xnor U25091 (N_25091,N_23735,N_23194);
nand U25092 (N_25092,N_23079,N_22915);
nand U25093 (N_25093,N_22825,N_23771);
nor U25094 (N_25094,N_23774,N_23744);
or U25095 (N_25095,N_23937,N_22932);
nor U25096 (N_25096,N_23397,N_23286);
nand U25097 (N_25097,N_23520,N_23208);
nor U25098 (N_25098,N_23158,N_23411);
or U25099 (N_25099,N_23509,N_22900);
nand U25100 (N_25100,N_23691,N_22981);
or U25101 (N_25101,N_23113,N_23370);
nor U25102 (N_25102,N_23382,N_23573);
nand U25103 (N_25103,N_23794,N_23495);
or U25104 (N_25104,N_23458,N_23376);
nor U25105 (N_25105,N_23803,N_23044);
and U25106 (N_25106,N_23094,N_23252);
xnor U25107 (N_25107,N_23438,N_23290);
nand U25108 (N_25108,N_23299,N_23875);
and U25109 (N_25109,N_22861,N_23157);
and U25110 (N_25110,N_22963,N_23658);
nand U25111 (N_25111,N_23685,N_23821);
nor U25112 (N_25112,N_23154,N_23952);
and U25113 (N_25113,N_23547,N_23957);
nand U25114 (N_25114,N_22936,N_23251);
xor U25115 (N_25115,N_23544,N_22874);
xnor U25116 (N_25116,N_23872,N_23151);
nand U25117 (N_25117,N_23971,N_23410);
nor U25118 (N_25118,N_23136,N_23320);
or U25119 (N_25119,N_23634,N_23755);
xnor U25120 (N_25120,N_23763,N_23374);
and U25121 (N_25121,N_23736,N_23238);
nand U25122 (N_25122,N_23172,N_23501);
nand U25123 (N_25123,N_22890,N_23199);
xor U25124 (N_25124,N_23550,N_23013);
nand U25125 (N_25125,N_23809,N_23656);
nand U25126 (N_25126,N_23625,N_23257);
nor U25127 (N_25127,N_23868,N_23375);
nand U25128 (N_25128,N_23926,N_22873);
xnor U25129 (N_25129,N_23029,N_23034);
and U25130 (N_25130,N_23492,N_23428);
or U25131 (N_25131,N_23533,N_23576);
nand U25132 (N_25132,N_23601,N_23334);
xnor U25133 (N_25133,N_23988,N_23497);
nor U25134 (N_25134,N_23543,N_23174);
or U25135 (N_25135,N_23673,N_23442);
nor U25136 (N_25136,N_23522,N_23225);
xor U25137 (N_25137,N_23033,N_23467);
nor U25138 (N_25138,N_23605,N_23065);
and U25139 (N_25139,N_23152,N_23147);
or U25140 (N_25140,N_23680,N_23615);
and U25141 (N_25141,N_22976,N_23781);
or U25142 (N_25142,N_23849,N_22998);
nor U25143 (N_25143,N_23057,N_23249);
xor U25144 (N_25144,N_23893,N_22830);
or U25145 (N_25145,N_22872,N_23038);
or U25146 (N_25146,N_23135,N_23632);
or U25147 (N_25147,N_23000,N_23694);
nor U25148 (N_25148,N_23927,N_22800);
or U25149 (N_25149,N_23057,N_23237);
and U25150 (N_25150,N_23975,N_23436);
or U25151 (N_25151,N_23116,N_23675);
xor U25152 (N_25152,N_23881,N_23581);
and U25153 (N_25153,N_23964,N_23225);
and U25154 (N_25154,N_22998,N_22852);
and U25155 (N_25155,N_23214,N_23847);
xnor U25156 (N_25156,N_23000,N_23203);
nand U25157 (N_25157,N_23022,N_23472);
nand U25158 (N_25158,N_22891,N_23919);
and U25159 (N_25159,N_22824,N_23583);
nor U25160 (N_25160,N_23545,N_22913);
or U25161 (N_25161,N_23501,N_23387);
xnor U25162 (N_25162,N_23568,N_23655);
nor U25163 (N_25163,N_23295,N_23916);
xnor U25164 (N_25164,N_22987,N_23568);
nand U25165 (N_25165,N_23246,N_23078);
nand U25166 (N_25166,N_23501,N_23124);
nor U25167 (N_25167,N_22873,N_23192);
xnor U25168 (N_25168,N_23586,N_23851);
nor U25169 (N_25169,N_23397,N_23192);
nor U25170 (N_25170,N_22834,N_23781);
or U25171 (N_25171,N_23934,N_23434);
or U25172 (N_25172,N_22962,N_23178);
nor U25173 (N_25173,N_23444,N_22876);
xor U25174 (N_25174,N_23412,N_23246);
nand U25175 (N_25175,N_23213,N_22806);
and U25176 (N_25176,N_23474,N_23410);
nor U25177 (N_25177,N_23461,N_22919);
xnor U25178 (N_25178,N_23476,N_23152);
nand U25179 (N_25179,N_22825,N_23244);
and U25180 (N_25180,N_23041,N_23461);
and U25181 (N_25181,N_23152,N_22871);
or U25182 (N_25182,N_23214,N_22913);
nand U25183 (N_25183,N_22822,N_23933);
xnor U25184 (N_25184,N_23934,N_23585);
xnor U25185 (N_25185,N_23382,N_23440);
nand U25186 (N_25186,N_23826,N_23341);
nand U25187 (N_25187,N_23008,N_22967);
and U25188 (N_25188,N_22967,N_23906);
and U25189 (N_25189,N_23830,N_23283);
or U25190 (N_25190,N_23428,N_23358);
nand U25191 (N_25191,N_23212,N_23886);
nor U25192 (N_25192,N_23715,N_23748);
nor U25193 (N_25193,N_23167,N_23259);
or U25194 (N_25194,N_23819,N_23699);
and U25195 (N_25195,N_23442,N_23895);
and U25196 (N_25196,N_23506,N_23822);
nand U25197 (N_25197,N_23889,N_23590);
xnor U25198 (N_25198,N_23483,N_23627);
nor U25199 (N_25199,N_23191,N_23531);
nand U25200 (N_25200,N_24600,N_24170);
nand U25201 (N_25201,N_24276,N_24283);
or U25202 (N_25202,N_24397,N_24369);
nand U25203 (N_25203,N_24336,N_24771);
nand U25204 (N_25204,N_24874,N_25048);
and U25205 (N_25205,N_25199,N_24153);
nand U25206 (N_25206,N_24197,N_24304);
nand U25207 (N_25207,N_24021,N_25065);
or U25208 (N_25208,N_24866,N_24297);
nor U25209 (N_25209,N_24694,N_24615);
nand U25210 (N_25210,N_24623,N_25044);
xor U25211 (N_25211,N_24830,N_24638);
or U25212 (N_25212,N_24541,N_24504);
and U25213 (N_25213,N_25186,N_24692);
nor U25214 (N_25214,N_24554,N_24570);
or U25215 (N_25215,N_24741,N_24838);
nor U25216 (N_25216,N_24005,N_24666);
and U25217 (N_25217,N_24140,N_25035);
nor U25218 (N_25218,N_24661,N_25087);
nor U25219 (N_25219,N_24743,N_24392);
nand U25220 (N_25220,N_24934,N_24267);
nor U25221 (N_25221,N_24904,N_24577);
and U25222 (N_25222,N_24821,N_24245);
and U25223 (N_25223,N_24427,N_24470);
nor U25224 (N_25224,N_24557,N_24752);
nand U25225 (N_25225,N_24842,N_24362);
nor U25226 (N_25226,N_24313,N_24522);
nor U25227 (N_25227,N_25144,N_25115);
or U25228 (N_25228,N_24176,N_24691);
or U25229 (N_25229,N_24498,N_25066);
and U25230 (N_25230,N_25107,N_24344);
xnor U25231 (N_25231,N_25088,N_24293);
nor U25232 (N_25232,N_24973,N_24211);
xor U25233 (N_25233,N_24308,N_24490);
or U25234 (N_25234,N_25069,N_24257);
and U25235 (N_25235,N_25197,N_24697);
xor U25236 (N_25236,N_24647,N_24596);
nor U25237 (N_25237,N_25021,N_24894);
xor U25238 (N_25238,N_24151,N_24612);
or U25239 (N_25239,N_24889,N_24418);
or U25240 (N_25240,N_24289,N_24062);
nor U25241 (N_25241,N_24837,N_24566);
nor U25242 (N_25242,N_25194,N_25170);
or U25243 (N_25243,N_24291,N_24368);
or U25244 (N_25244,N_24201,N_24032);
and U25245 (N_25245,N_25143,N_25051);
nor U25246 (N_25246,N_24952,N_24869);
and U25247 (N_25247,N_25156,N_24801);
nor U25248 (N_25248,N_25191,N_24488);
and U25249 (N_25249,N_24388,N_24559);
nand U25250 (N_25250,N_25128,N_24177);
nand U25251 (N_25251,N_24063,N_24004);
nor U25252 (N_25252,N_24654,N_24426);
nand U25253 (N_25253,N_24909,N_24811);
nor U25254 (N_25254,N_24215,N_24746);
and U25255 (N_25255,N_24797,N_24054);
and U25256 (N_25256,N_25080,N_24945);
and U25257 (N_25257,N_24482,N_24076);
xnor U25258 (N_25258,N_24936,N_25060);
nor U25259 (N_25259,N_24493,N_24980);
and U25260 (N_25260,N_24673,N_24444);
nor U25261 (N_25261,N_24066,N_24331);
xnor U25262 (N_25262,N_24718,N_24687);
nor U25263 (N_25263,N_24593,N_24068);
or U25264 (N_25264,N_24385,N_24650);
xor U25265 (N_25265,N_24027,N_24480);
and U25266 (N_25266,N_25047,N_25120);
nor U25267 (N_25267,N_24376,N_24337);
xnor U25268 (N_25268,N_24784,N_24648);
or U25269 (N_25269,N_25054,N_24191);
xnor U25270 (N_25270,N_24759,N_24355);
xnor U25271 (N_25271,N_24792,N_24766);
and U25272 (N_25272,N_24014,N_24202);
or U25273 (N_25273,N_24637,N_24079);
nand U25274 (N_25274,N_24679,N_24805);
and U25275 (N_25275,N_24281,N_24102);
xnor U25276 (N_25276,N_24359,N_24535);
nor U25277 (N_25277,N_24192,N_24505);
and U25278 (N_25278,N_25058,N_24720);
nand U25279 (N_25279,N_24431,N_24982);
nor U25280 (N_25280,N_24851,N_24603);
or U25281 (N_25281,N_24058,N_24745);
nor U25282 (N_25282,N_24828,N_25000);
xnor U25283 (N_25283,N_24083,N_24879);
nor U25284 (N_25284,N_24437,N_24015);
or U25285 (N_25285,N_24365,N_24978);
xnor U25286 (N_25286,N_24877,N_24783);
nand U25287 (N_25287,N_24409,N_24234);
nor U25288 (N_25288,N_24601,N_24387);
nand U25289 (N_25289,N_25002,N_24921);
xnor U25290 (N_25290,N_24017,N_24611);
xor U25291 (N_25291,N_24918,N_24757);
xnor U25292 (N_25292,N_24206,N_24056);
xor U25293 (N_25293,N_24499,N_24575);
nor U25294 (N_25294,N_25032,N_24574);
or U25295 (N_25295,N_25159,N_24350);
and U25296 (N_25296,N_24737,N_25020);
or U25297 (N_25297,N_24824,N_24629);
nand U25298 (N_25298,N_25071,N_24342);
xor U25299 (N_25299,N_25050,N_24906);
nand U25300 (N_25300,N_25057,N_24925);
nor U25301 (N_25301,N_24028,N_24724);
and U25302 (N_25302,N_24972,N_24424);
nor U25303 (N_25303,N_24163,N_24962);
and U25304 (N_25304,N_24545,N_24061);
and U25305 (N_25305,N_24303,N_24793);
or U25306 (N_25306,N_24011,N_24338);
nand U25307 (N_25307,N_24576,N_25140);
nand U25308 (N_25308,N_24562,N_25151);
or U25309 (N_25309,N_24731,N_24872);
nand U25310 (N_25310,N_24560,N_25135);
xnor U25311 (N_25311,N_24209,N_24179);
xnor U25312 (N_25312,N_24619,N_24332);
or U25313 (N_25313,N_25097,N_25001);
nor U25314 (N_25314,N_24117,N_24977);
and U25315 (N_25315,N_25009,N_25185);
xor U25316 (N_25316,N_24002,N_24836);
xor U25317 (N_25317,N_24243,N_24573);
xor U25318 (N_25318,N_24530,N_24935);
nand U25319 (N_25319,N_24966,N_24967);
nand U25320 (N_25320,N_24280,N_24550);
or U25321 (N_25321,N_24226,N_24684);
nor U25322 (N_25322,N_24279,N_24441);
nand U25323 (N_25323,N_24510,N_24398);
and U25324 (N_25324,N_24404,N_25043);
nand U25325 (N_25325,N_25068,N_24779);
or U25326 (N_25326,N_25030,N_24951);
and U25327 (N_25327,N_24379,N_25034);
xnor U25328 (N_25328,N_24826,N_25125);
nand U25329 (N_25329,N_24009,N_24610);
xor U25330 (N_25330,N_25136,N_25090);
nor U25331 (N_25331,N_24440,N_24264);
xnor U25332 (N_25332,N_24908,N_24517);
xor U25333 (N_25333,N_24306,N_24655);
nand U25334 (N_25334,N_24091,N_24118);
nor U25335 (N_25335,N_24685,N_24583);
nor U25336 (N_25336,N_25134,N_24780);
nand U25337 (N_25337,N_24592,N_24100);
and U25338 (N_25338,N_24662,N_24782);
or U25339 (N_25339,N_24563,N_24549);
and U25340 (N_25340,N_24558,N_25130);
nor U25341 (N_25341,N_24300,N_24660);
or U25342 (N_25342,N_24185,N_24806);
and U25343 (N_25343,N_24723,N_24137);
xor U25344 (N_25344,N_24178,N_25164);
nand U25345 (N_25345,N_24030,N_24224);
xor U25346 (N_25346,N_24210,N_25129);
or U25347 (N_25347,N_24298,N_24423);
and U25348 (N_25348,N_24328,N_24835);
nand U25349 (N_25349,N_24204,N_25019);
nor U25350 (N_25350,N_25056,N_24503);
or U25351 (N_25351,N_24325,N_24753);
nor U25352 (N_25352,N_24653,N_24479);
or U25353 (N_25353,N_24950,N_25049);
nand U25354 (N_25354,N_24247,N_24820);
xnor U25355 (N_25355,N_24106,N_24683);
nor U25356 (N_25356,N_24873,N_24349);
nand U25357 (N_25357,N_24116,N_24773);
nand U25358 (N_25358,N_24269,N_24096);
and U25359 (N_25359,N_24719,N_24326);
and U25360 (N_25360,N_24235,N_24284);
xor U25361 (N_25361,N_24103,N_24233);
or U25362 (N_25362,N_24844,N_24940);
nor U25363 (N_25363,N_24274,N_24513);
or U25364 (N_25364,N_24133,N_25036);
nand U25365 (N_25365,N_24120,N_24891);
nand U25366 (N_25366,N_24165,N_24132);
or U25367 (N_25367,N_24788,N_24931);
nand U25368 (N_25368,N_25055,N_24639);
and U25369 (N_25369,N_25138,N_24157);
xor U25370 (N_25370,N_24682,N_24255);
or U25371 (N_25371,N_24082,N_24594);
and U25372 (N_25372,N_24394,N_24277);
nor U25373 (N_25373,N_24714,N_24036);
and U25374 (N_25374,N_24406,N_24670);
and U25375 (N_25375,N_24749,N_24067);
xor U25376 (N_25376,N_24074,N_25193);
nor U25377 (N_25377,N_25196,N_24136);
nor U25378 (N_25378,N_24126,N_24466);
xor U25379 (N_25379,N_25133,N_24794);
or U25380 (N_25380,N_24171,N_24196);
xor U25381 (N_25381,N_24436,N_25079);
or U25382 (N_25382,N_24785,N_24711);
nand U25383 (N_25383,N_24238,N_24640);
nor U25384 (N_25384,N_24567,N_24726);
nor U25385 (N_25385,N_25084,N_24857);
or U25386 (N_25386,N_25073,N_25100);
or U25387 (N_25387,N_24981,N_24420);
nor U25388 (N_25388,N_24569,N_24667);
nand U25389 (N_25389,N_25010,N_25027);
and U25390 (N_25390,N_24018,N_24327);
or U25391 (N_25391,N_24769,N_24875);
nor U25392 (N_25392,N_24789,N_24833);
nand U25393 (N_25393,N_24003,N_24703);
and U25394 (N_25394,N_24887,N_24860);
nand U25395 (N_25395,N_24502,N_24346);
and U25396 (N_25396,N_24781,N_24104);
or U25397 (N_25397,N_24910,N_25007);
xnor U25398 (N_25398,N_24294,N_25198);
nand U25399 (N_25399,N_24135,N_25141);
or U25400 (N_25400,N_24777,N_24963);
xor U25401 (N_25401,N_24770,N_24045);
nor U25402 (N_25402,N_24495,N_24501);
and U25403 (N_25403,N_24485,N_24472);
nor U25404 (N_25404,N_24162,N_24627);
nor U25405 (N_25405,N_24526,N_24086);
or U25406 (N_25406,N_25145,N_25040);
or U25407 (N_25407,N_24845,N_25174);
nor U25408 (N_25408,N_24383,N_24022);
or U25409 (N_25409,N_24544,N_24145);
or U25410 (N_25410,N_24421,N_24871);
xnor U25411 (N_25411,N_24047,N_24902);
xnor U25412 (N_25412,N_24214,N_24849);
xnor U25413 (N_25413,N_24194,N_24360);
nand U25414 (N_25414,N_24917,N_24285);
and U25415 (N_25415,N_24863,N_24416);
or U25416 (N_25416,N_25158,N_24055);
xnor U25417 (N_25417,N_24377,N_24795);
xnor U25418 (N_25418,N_24217,N_24552);
nor U25419 (N_25419,N_24919,N_24626);
nand U25420 (N_25420,N_24861,N_24671);
or U25421 (N_25421,N_24099,N_24748);
and U25422 (N_25422,N_24129,N_24578);
and U25423 (N_25423,N_24776,N_24310);
nand U25424 (N_25424,N_25154,N_24515);
nor U25425 (N_25425,N_24609,N_24335);
nor U25426 (N_25426,N_24579,N_25082);
and U25427 (N_25427,N_25184,N_24881);
or U25428 (N_25428,N_24270,N_24649);
nor U25429 (N_25429,N_24001,N_25016);
or U25430 (N_25430,N_24373,N_24744);
xor U25431 (N_25431,N_25085,N_24189);
nor U25432 (N_25432,N_25108,N_24324);
or U25433 (N_25433,N_24075,N_25180);
xor U25434 (N_25434,N_24758,N_24669);
and U25435 (N_25435,N_24168,N_24097);
nand U25436 (N_25436,N_24763,N_25192);
xor U25437 (N_25437,N_24531,N_24699);
nor U25438 (N_25438,N_25045,N_24876);
and U25439 (N_25439,N_25162,N_24494);
nor U25440 (N_25440,N_24605,N_24419);
and U25441 (N_25441,N_24943,N_24266);
nand U25442 (N_25442,N_24546,N_24898);
nor U25443 (N_25443,N_24812,N_24613);
nor U25444 (N_25444,N_24395,N_24125);
xor U25445 (N_25445,N_24946,N_24668);
nor U25446 (N_25446,N_24432,N_24542);
or U25447 (N_25447,N_24822,N_25139);
nand U25448 (N_25448,N_24109,N_24856);
and U25449 (N_25449,N_24476,N_24329);
and U25450 (N_25450,N_25083,N_24451);
nor U25451 (N_25451,N_24455,N_24461);
and U25452 (N_25452,N_24534,N_24853);
nor U25453 (N_25453,N_24469,N_24708);
or U25454 (N_25454,N_24568,N_24511);
or U25455 (N_25455,N_24536,N_24174);
xor U25456 (N_25456,N_24598,N_24516);
and U25457 (N_25457,N_24259,N_24307);
and U25458 (N_25458,N_24070,N_24019);
or U25459 (N_25459,N_24721,N_24452);
nand U25460 (N_25460,N_24314,N_24686);
nor U25461 (N_25461,N_24957,N_24315);
xor U25462 (N_25462,N_24216,N_24913);
nor U25463 (N_25463,N_24706,N_24924);
nand U25464 (N_25464,N_24616,N_24870);
and U25465 (N_25465,N_24039,N_25005);
or U25466 (N_25466,N_24084,N_24435);
nor U25467 (N_25467,N_24242,N_24363);
or U25468 (N_25468,N_24345,N_24240);
xor U25469 (N_25469,N_24087,N_24540);
and U25470 (N_25470,N_25175,N_24664);
or U25471 (N_25471,N_24868,N_24353);
or U25472 (N_25472,N_24282,N_24762);
and U25473 (N_25473,N_24339,N_25099);
nor U25474 (N_25474,N_24987,N_24159);
or U25475 (N_25475,N_24712,N_24333);
and U25476 (N_25476,N_24035,N_24029);
xor U25477 (N_25477,N_24646,N_24088);
xor U25478 (N_25478,N_24374,N_24895);
xor U25479 (N_25479,N_24768,N_24900);
nand U25480 (N_25480,N_24393,N_24186);
nor U25481 (N_25481,N_24905,N_24636);
or U25482 (N_25482,N_25092,N_24674);
nand U25483 (N_25483,N_25124,N_24481);
or U25484 (N_25484,N_24190,N_24134);
nor U25485 (N_25485,N_24254,N_24149);
and U25486 (N_25486,N_24523,N_24886);
xor U25487 (N_25487,N_25106,N_24010);
or U25488 (N_25488,N_24413,N_24341);
nand U25489 (N_25489,N_25132,N_24941);
nor U25490 (N_25490,N_24740,N_24312);
or U25491 (N_25491,N_24474,N_25038);
xor U25492 (N_25492,N_25119,N_24043);
nor U25493 (N_25493,N_24319,N_24976);
nand U25494 (N_25494,N_24700,N_24180);
or U25495 (N_25495,N_24220,N_25042);
or U25496 (N_25496,N_24767,N_24525);
nor U25497 (N_25497,N_24754,N_24878);
nor U25498 (N_25498,N_24890,N_25155);
nand U25499 (N_25499,N_24829,N_24831);
and U25500 (N_25500,N_25122,N_24581);
or U25501 (N_25501,N_24446,N_24954);
nand U25502 (N_25502,N_24286,N_24487);
nand U25503 (N_25503,N_24738,N_24808);
xor U25504 (N_25504,N_24704,N_24624);
and U25505 (N_25505,N_25183,N_25094);
nand U25506 (N_25506,N_24497,N_24848);
nor U25507 (N_25507,N_24729,N_24473);
or U25508 (N_25508,N_24996,N_24000);
nor U25509 (N_25509,N_24926,N_25188);
or U25510 (N_25510,N_24391,N_24361);
xor U25511 (N_25511,N_24929,N_24632);
or U25512 (N_25512,N_24443,N_24024);
xnor U25513 (N_25513,N_24475,N_24939);
nor U25514 (N_25514,N_24477,N_24960);
and U25515 (N_25515,N_24364,N_24652);
and U25516 (N_25516,N_24089,N_24663);
nand U25517 (N_25517,N_24439,N_24903);
nand U25518 (N_25518,N_24340,N_24617);
and U25519 (N_25519,N_24454,N_24053);
and U25520 (N_25520,N_24986,N_24457);
nand U25521 (N_25521,N_25025,N_24261);
nand U25522 (N_25522,N_24899,N_24884);
xor U25523 (N_25523,N_24271,N_24071);
nor U25524 (N_25524,N_24356,N_24816);
and U25525 (N_25525,N_24352,N_25160);
and U25526 (N_25526,N_24641,N_24146);
nand U25527 (N_25527,N_25150,N_24205);
xnor U25528 (N_25528,N_24532,N_25110);
nand U25529 (N_25529,N_24519,N_24048);
or U25530 (N_25530,N_24302,N_24916);
nor U25531 (N_25531,N_24250,N_24130);
xor U25532 (N_25532,N_24888,N_24371);
and U25533 (N_25533,N_24739,N_24907);
nor U25534 (N_25534,N_24858,N_25116);
or U25535 (N_25535,N_24221,N_24173);
or U25536 (N_25536,N_24644,N_24260);
xnor U25537 (N_25537,N_24651,N_24597);
nor U25538 (N_25538,N_24778,N_24923);
nand U25539 (N_25539,N_24543,N_24599);
nand U25540 (N_25540,N_24533,N_24405);
nor U25541 (N_25541,N_24803,N_24678);
and U25542 (N_25542,N_24411,N_24722);
xor U25543 (N_25543,N_24154,N_25026);
nor U25544 (N_25544,N_24462,N_25163);
xor U25545 (N_25545,N_25111,N_24584);
nor U25546 (N_25546,N_24456,N_24990);
or U25547 (N_25547,N_24232,N_24412);
or U25548 (N_25548,N_24832,N_24183);
xnor U25549 (N_25549,N_24296,N_24725);
nor U25550 (N_25550,N_24228,N_24122);
xnor U25551 (N_25551,N_24657,N_24867);
or U25552 (N_25552,N_24509,N_24244);
nand U25553 (N_25553,N_24357,N_24484);
or U25554 (N_25554,N_24807,N_25113);
xor U25555 (N_25555,N_25061,N_24538);
or U25556 (N_25556,N_24930,N_25123);
or U25557 (N_25557,N_25109,N_24492);
and U25558 (N_25558,N_24548,N_25102);
or U25559 (N_25559,N_24222,N_25014);
and U25560 (N_25560,N_24425,N_25146);
nor U25561 (N_25561,N_24897,N_24292);
or U25562 (N_25562,N_24968,N_24995);
nand U25563 (N_25563,N_24236,N_24827);
and U25564 (N_25564,N_24370,N_24311);
and U25565 (N_25565,N_24317,N_24105);
or U25566 (N_25566,N_25172,N_24169);
nand U25567 (N_25567,N_24944,N_24007);
or U25568 (N_25568,N_25029,N_25095);
nor U25569 (N_25569,N_24702,N_24823);
and U25570 (N_25570,N_24367,N_24156);
nand U25571 (N_25571,N_24561,N_25070);
xnor U25572 (N_25572,N_24988,N_24251);
and U25573 (N_25573,N_24813,N_24320);
and U25574 (N_25574,N_24072,N_24152);
or U25575 (N_25575,N_24429,N_24942);
xnor U25576 (N_25576,N_24248,N_24471);
nor U25577 (N_25577,N_24031,N_25168);
xor U25578 (N_25578,N_24016,N_24127);
nor U25579 (N_25579,N_24442,N_25182);
xnor U25580 (N_25580,N_24933,N_24880);
and U25581 (N_25581,N_24677,N_25173);
or U25582 (N_25582,N_24050,N_24959);
xnor U25583 (N_25583,N_24334,N_25105);
nand U25584 (N_25584,N_25031,N_24108);
nand U25585 (N_25585,N_25017,N_25190);
nor U25586 (N_25586,N_24564,N_24733);
or U25587 (N_25587,N_24809,N_24166);
or U25588 (N_25588,N_25033,N_25195);
nor U25589 (N_25589,N_24920,N_24551);
nand U25590 (N_25590,N_24110,N_24124);
and U25591 (N_25591,N_24184,N_24642);
nor U25592 (N_25592,N_24539,N_24458);
nor U25593 (N_25593,N_24938,N_25103);
or U25594 (N_25594,N_24607,N_24882);
and U25595 (N_25595,N_25153,N_24449);
and U25596 (N_25596,N_24148,N_25077);
nor U25597 (N_25597,N_25081,N_24730);
nand U25598 (N_25598,N_25089,N_24843);
nand U25599 (N_25599,N_24696,N_24046);
nor U25600 (N_25600,N_24198,N_24098);
nor U25601 (N_25601,N_24992,N_24112);
or U25602 (N_25602,N_24630,N_24464);
or U25603 (N_25603,N_25022,N_24382);
nor U25604 (N_25604,N_24524,N_25112);
and U25605 (N_25605,N_24804,N_24203);
nand U25606 (N_25606,N_25152,N_24528);
nor U25607 (N_25607,N_24199,N_24188);
or U25608 (N_25608,N_24911,N_24852);
nand U25609 (N_25609,N_24761,N_24059);
or U25610 (N_25610,N_24410,N_24288);
xor U25611 (N_25611,N_24512,N_24727);
xnor U25612 (N_25612,N_24862,N_24085);
xnor U25613 (N_25613,N_25075,N_24764);
nor U25614 (N_25614,N_24508,N_24675);
or U25615 (N_25615,N_24756,N_24167);
nand U25616 (N_25616,N_24659,N_24975);
nor U25617 (N_25617,N_24791,N_24113);
and U25618 (N_25618,N_24064,N_24521);
and U25619 (N_25619,N_24855,N_24081);
nor U25620 (N_25620,N_24347,N_24321);
nor U25621 (N_25621,N_24268,N_24212);
and U25622 (N_25622,N_24396,N_25046);
nor U25623 (N_25623,N_24138,N_24077);
xnor U25624 (N_25624,N_24953,N_24690);
and U25625 (N_25625,N_24263,N_24323);
and U25626 (N_25626,N_24590,N_24013);
nor U25627 (N_25627,N_24621,N_25171);
nor U25628 (N_25628,N_24207,N_24802);
or U25629 (N_25629,N_24408,N_24052);
or U25630 (N_25630,N_24854,N_24040);
nand U25631 (N_25631,N_25096,N_24556);
nand U25632 (N_25632,N_24101,N_24229);
nor U25633 (N_25633,N_25086,N_24841);
or U25634 (N_25634,N_24527,N_24817);
nand U25635 (N_25635,N_25117,N_24810);
nor U25636 (N_25636,N_24565,N_25006);
and U25637 (N_25637,N_24914,N_24625);
and U25638 (N_25638,N_24864,N_24932);
xor U25639 (N_25639,N_24815,N_24380);
nand U25640 (N_25640,N_24262,N_24709);
nor U25641 (N_25641,N_25165,N_24728);
and U25642 (N_25642,N_25093,N_25074);
and U25643 (N_25643,N_24734,N_24705);
xnor U25644 (N_25644,N_24023,N_25091);
and U25645 (N_25645,N_24008,N_24998);
and U25646 (N_25646,N_24645,N_25179);
and U25647 (N_25647,N_25161,N_24537);
xor U25648 (N_25648,N_24384,N_24131);
and U25649 (N_25649,N_24713,N_24468);
xor U25650 (N_25650,N_24239,N_24847);
and U25651 (N_25651,N_24114,N_25149);
nand U25652 (N_25652,N_25098,N_24463);
or U25653 (N_25653,N_24478,N_24786);
nor U25654 (N_25654,N_24164,N_24272);
nand U25655 (N_25655,N_24614,N_24073);
or U25656 (N_25656,N_24119,N_25187);
xnor U25657 (N_25657,N_24586,N_24514);
and U25658 (N_25658,N_24372,N_24253);
xnor U25659 (N_25659,N_24287,N_24839);
nor U25660 (N_25660,N_24717,N_24275);
and U25661 (N_25661,N_24618,N_24927);
or U25662 (N_25662,N_24467,N_24695);
or U25663 (N_25663,N_24735,N_24892);
nand U25664 (N_25664,N_24760,N_24643);
and U25665 (N_25665,N_24606,N_25013);
xnor U25666 (N_25666,N_24750,N_24366);
and U25667 (N_25667,N_24922,N_25039);
nor U25668 (N_25668,N_25004,N_24460);
nand U25669 (N_25669,N_24399,N_24547);
nor U25670 (N_25670,N_24883,N_24249);
nand U25671 (N_25671,N_24459,N_24265);
nor U25672 (N_25672,N_24378,N_24489);
or U25673 (N_25673,N_24520,N_25011);
or U25674 (N_25674,N_24620,N_24330);
and U25675 (N_25675,N_24796,N_25118);
nor U25676 (N_25676,N_24375,N_24223);
nor U25677 (N_25677,N_24107,N_24080);
nand U25678 (N_25678,N_24231,N_24258);
nand U25679 (N_25679,N_24819,N_24969);
and U25680 (N_25680,N_24182,N_25166);
nand U25681 (N_25681,N_24486,N_24983);
and U25682 (N_25682,N_25053,N_24672);
nor U25683 (N_25683,N_24580,N_25037);
nand U25684 (N_25684,N_24219,N_24985);
nand U25685 (N_25685,N_24295,N_24438);
xor U25686 (N_25686,N_24025,N_24688);
nand U25687 (N_25687,N_24111,N_24041);
nand U25688 (N_25688,N_24230,N_24358);
nand U25689 (N_25689,N_24160,N_25127);
nand U25690 (N_25690,N_24093,N_24123);
nor U25691 (N_25691,N_25157,N_25177);
nand U25692 (N_25692,N_24587,N_24430);
and U25693 (N_25693,N_25104,N_24747);
or U25694 (N_25694,N_24090,N_24422);
or U25695 (N_25695,N_24033,N_24896);
and U25696 (N_25696,N_24814,N_24755);
or U25697 (N_25697,N_24401,N_24390);
xnor U25698 (N_25698,N_24447,N_25101);
or U25699 (N_25699,N_24885,N_24225);
xnor U25700 (N_25700,N_24144,N_24800);
xor U25701 (N_25701,N_24915,N_24970);
xnor U25702 (N_25702,N_24991,N_24246);
or U25703 (N_25703,N_24553,N_24187);
nor U25704 (N_25704,N_24850,N_24020);
nand U25705 (N_25705,N_24034,N_24094);
nand U25706 (N_25706,N_24964,N_24937);
nor U25707 (N_25707,N_24381,N_24961);
xnor U25708 (N_25708,N_24354,N_24057);
nor U25709 (N_25709,N_24588,N_24128);
nand U25710 (N_25710,N_24060,N_24434);
xor U25711 (N_25711,N_24445,N_24252);
nand U25712 (N_25712,N_24971,N_24608);
xor U25713 (N_25713,N_24751,N_24433);
nand U25714 (N_25714,N_25147,N_24115);
nand U25715 (N_25715,N_24965,N_24500);
nor U25716 (N_25716,N_24218,N_24604);
xnor U25717 (N_25717,N_24496,N_24631);
xnor U25718 (N_25718,N_25064,N_24507);
nor U25719 (N_25719,N_24774,N_24979);
xnor U25720 (N_25720,N_24958,N_24227);
or U25721 (N_25721,N_24309,N_25137);
and U25722 (N_25722,N_24710,N_24465);
nor U25723 (N_25723,N_24491,N_24997);
nor U25724 (N_25724,N_24448,N_24141);
nor U25725 (N_25725,N_24316,N_25176);
nand U25726 (N_25726,N_25167,N_24037);
and U25727 (N_25727,N_24078,N_25142);
nand U25728 (N_25728,N_24181,N_24042);
and U25729 (N_25729,N_25052,N_24665);
xor U25730 (N_25730,N_24984,N_24044);
xor U25731 (N_25731,N_24676,N_24483);
and U25732 (N_25732,N_25072,N_24241);
nor U25733 (N_25733,N_25015,N_24846);
xor U25734 (N_25734,N_24840,N_24453);
xor U25735 (N_25735,N_24142,N_24121);
and U25736 (N_25736,N_24278,N_24947);
and U25737 (N_25737,N_24989,N_24999);
xnor U25738 (N_25738,N_24693,N_24305);
or U25739 (N_25739,N_24161,N_24742);
nand U25740 (N_25740,N_24402,N_24591);
nand U25741 (N_25741,N_24012,N_25028);
or U25742 (N_25742,N_24428,N_24139);
xor U25743 (N_25743,N_25181,N_24318);
and U25744 (N_25744,N_24656,N_24901);
and U25745 (N_25745,N_25062,N_24301);
nand U25746 (N_25746,N_24818,N_25063);
xor U25747 (N_25747,N_24143,N_25059);
nor U25748 (N_25748,N_24993,N_24707);
xnor U25749 (N_25749,N_24912,N_25189);
xor U25750 (N_25750,N_24506,N_24213);
and U25751 (N_25751,N_24582,N_24955);
and U25752 (N_25752,N_24956,N_24765);
nor U25753 (N_25753,N_24628,N_24150);
nor U25754 (N_25754,N_24635,N_24208);
xnor U25755 (N_25755,N_25024,N_24732);
nand U25756 (N_25756,N_24589,N_24417);
nor U25757 (N_25757,N_24736,N_24974);
nand U25758 (N_25758,N_25148,N_25114);
nand U25759 (N_25759,N_24237,N_24658);
and U25760 (N_25760,N_24572,N_24200);
and U25761 (N_25761,N_24689,N_24299);
nand U25762 (N_25762,N_24389,N_24787);
xnor U25763 (N_25763,N_24256,N_24715);
xnor U25764 (N_25764,N_24147,N_24834);
nor U25765 (N_25765,N_24415,N_24414);
nor U25766 (N_25766,N_24290,N_24633);
nor U25767 (N_25767,N_24772,N_24518);
nor U25768 (N_25768,N_24348,N_24049);
and U25769 (N_25769,N_24158,N_24006);
and U25770 (N_25770,N_24195,N_24193);
or U25771 (N_25771,N_24865,N_24273);
nor U25772 (N_25772,N_24038,N_24716);
xnor U25773 (N_25773,N_25169,N_24859);
xnor U25774 (N_25774,N_25067,N_24634);
or U25775 (N_25775,N_24450,N_25008);
nor U25776 (N_25776,N_24681,N_24602);
nand U25777 (N_25777,N_24928,N_25018);
or U25778 (N_25778,N_24698,N_24994);
or U25779 (N_25779,N_24949,N_24529);
xnor U25780 (N_25780,N_24799,N_24555);
or U25781 (N_25781,N_24069,N_24585);
and U25782 (N_25782,N_24825,N_25023);
nand U25783 (N_25783,N_25078,N_24351);
nand U25784 (N_25784,N_24701,N_24400);
or U25785 (N_25785,N_25041,N_24155);
nor U25786 (N_25786,N_25121,N_24175);
or U25787 (N_25787,N_25003,N_24403);
nand U25788 (N_25788,N_24948,N_24775);
xnor U25789 (N_25789,N_25076,N_24571);
or U25790 (N_25790,N_24065,N_24095);
or U25791 (N_25791,N_24386,N_24092);
nand U25792 (N_25792,N_24798,N_25178);
nand U25793 (N_25793,N_24322,N_24790);
nor U25794 (N_25794,N_25012,N_24026);
nand U25795 (N_25795,N_25131,N_24172);
and U25796 (N_25796,N_24407,N_24893);
xor U25797 (N_25797,N_24051,N_25126);
xor U25798 (N_25798,N_24622,N_24343);
nor U25799 (N_25799,N_24680,N_24595);
and U25800 (N_25800,N_24151,N_25049);
or U25801 (N_25801,N_25114,N_24818);
nand U25802 (N_25802,N_24556,N_24046);
nor U25803 (N_25803,N_24645,N_24155);
xnor U25804 (N_25804,N_24021,N_24704);
or U25805 (N_25805,N_24277,N_24981);
and U25806 (N_25806,N_24131,N_24698);
nor U25807 (N_25807,N_24316,N_24542);
and U25808 (N_25808,N_24926,N_24368);
nand U25809 (N_25809,N_24499,N_24923);
or U25810 (N_25810,N_24038,N_24445);
nand U25811 (N_25811,N_24500,N_24045);
or U25812 (N_25812,N_24392,N_24797);
or U25813 (N_25813,N_24036,N_24909);
nand U25814 (N_25814,N_24586,N_24163);
and U25815 (N_25815,N_25009,N_25155);
or U25816 (N_25816,N_24733,N_25157);
or U25817 (N_25817,N_24656,N_24662);
nand U25818 (N_25818,N_24366,N_24789);
nor U25819 (N_25819,N_24156,N_24735);
nor U25820 (N_25820,N_24617,N_25118);
nor U25821 (N_25821,N_24159,N_24163);
or U25822 (N_25822,N_24236,N_24259);
or U25823 (N_25823,N_25184,N_24180);
nor U25824 (N_25824,N_24565,N_24237);
nor U25825 (N_25825,N_24350,N_24713);
and U25826 (N_25826,N_24295,N_24561);
nand U25827 (N_25827,N_24594,N_24794);
and U25828 (N_25828,N_24207,N_24249);
and U25829 (N_25829,N_24928,N_24729);
nor U25830 (N_25830,N_25187,N_24415);
nor U25831 (N_25831,N_24616,N_24627);
or U25832 (N_25832,N_24687,N_25090);
nor U25833 (N_25833,N_25130,N_24867);
xnor U25834 (N_25834,N_24515,N_24072);
nand U25835 (N_25835,N_24817,N_24448);
or U25836 (N_25836,N_25119,N_24375);
xnor U25837 (N_25837,N_24923,N_24735);
or U25838 (N_25838,N_25138,N_24762);
xor U25839 (N_25839,N_24657,N_24592);
and U25840 (N_25840,N_24742,N_24859);
nor U25841 (N_25841,N_24544,N_24708);
or U25842 (N_25842,N_24274,N_25157);
nor U25843 (N_25843,N_24839,N_24771);
xnor U25844 (N_25844,N_25053,N_24643);
or U25845 (N_25845,N_24641,N_25006);
nand U25846 (N_25846,N_24268,N_25021);
nor U25847 (N_25847,N_24467,N_24722);
nand U25848 (N_25848,N_25158,N_24919);
or U25849 (N_25849,N_24925,N_24102);
or U25850 (N_25850,N_24169,N_24595);
or U25851 (N_25851,N_24796,N_24048);
nor U25852 (N_25852,N_24313,N_25068);
nor U25853 (N_25853,N_24747,N_24560);
xor U25854 (N_25854,N_24191,N_24299);
xnor U25855 (N_25855,N_24319,N_24382);
and U25856 (N_25856,N_24655,N_24960);
nand U25857 (N_25857,N_24482,N_24824);
and U25858 (N_25858,N_25023,N_25056);
or U25859 (N_25859,N_24143,N_25032);
or U25860 (N_25860,N_24585,N_24134);
nor U25861 (N_25861,N_25088,N_24354);
nand U25862 (N_25862,N_25043,N_25001);
nor U25863 (N_25863,N_24252,N_24073);
and U25864 (N_25864,N_24508,N_24521);
nand U25865 (N_25865,N_24893,N_24268);
nor U25866 (N_25866,N_24873,N_24238);
nand U25867 (N_25867,N_24721,N_24139);
xnor U25868 (N_25868,N_24975,N_24904);
nor U25869 (N_25869,N_24166,N_25115);
nor U25870 (N_25870,N_24286,N_24149);
and U25871 (N_25871,N_24950,N_24658);
nor U25872 (N_25872,N_24548,N_25175);
xnor U25873 (N_25873,N_24137,N_24503);
or U25874 (N_25874,N_24317,N_24412);
or U25875 (N_25875,N_24588,N_24413);
nand U25876 (N_25876,N_24741,N_24920);
xor U25877 (N_25877,N_25190,N_24062);
nor U25878 (N_25878,N_24648,N_25006);
or U25879 (N_25879,N_24058,N_24523);
and U25880 (N_25880,N_24132,N_24931);
nor U25881 (N_25881,N_25175,N_24371);
or U25882 (N_25882,N_24366,N_24719);
and U25883 (N_25883,N_24523,N_24760);
and U25884 (N_25884,N_25023,N_24981);
and U25885 (N_25885,N_24293,N_24799);
xor U25886 (N_25886,N_24379,N_24147);
nor U25887 (N_25887,N_24122,N_24317);
and U25888 (N_25888,N_24184,N_24603);
nand U25889 (N_25889,N_24261,N_24682);
or U25890 (N_25890,N_24458,N_24674);
nand U25891 (N_25891,N_24437,N_24609);
or U25892 (N_25892,N_24989,N_24553);
xor U25893 (N_25893,N_24088,N_24308);
xnor U25894 (N_25894,N_24662,N_24007);
nand U25895 (N_25895,N_25060,N_24116);
and U25896 (N_25896,N_24011,N_25075);
and U25897 (N_25897,N_24291,N_25153);
nor U25898 (N_25898,N_24423,N_24217);
and U25899 (N_25899,N_24605,N_24764);
nand U25900 (N_25900,N_24596,N_25127);
nor U25901 (N_25901,N_24704,N_25010);
nor U25902 (N_25902,N_24236,N_24494);
nand U25903 (N_25903,N_24849,N_24411);
or U25904 (N_25904,N_24305,N_25198);
and U25905 (N_25905,N_25127,N_24601);
xnor U25906 (N_25906,N_24020,N_24744);
xnor U25907 (N_25907,N_25089,N_24842);
xnor U25908 (N_25908,N_24561,N_24065);
nor U25909 (N_25909,N_24845,N_24358);
nand U25910 (N_25910,N_24023,N_24153);
and U25911 (N_25911,N_25197,N_24769);
nor U25912 (N_25912,N_24612,N_24672);
or U25913 (N_25913,N_25121,N_24467);
nand U25914 (N_25914,N_24222,N_24540);
xor U25915 (N_25915,N_25085,N_24445);
nor U25916 (N_25916,N_25031,N_24055);
nor U25917 (N_25917,N_24404,N_24980);
nor U25918 (N_25918,N_24948,N_24625);
or U25919 (N_25919,N_24099,N_24491);
nor U25920 (N_25920,N_25023,N_24317);
xor U25921 (N_25921,N_24411,N_24562);
or U25922 (N_25922,N_24378,N_24444);
xnor U25923 (N_25923,N_24011,N_24597);
nor U25924 (N_25924,N_24244,N_24888);
nor U25925 (N_25925,N_24644,N_24978);
and U25926 (N_25926,N_24977,N_24690);
xor U25927 (N_25927,N_24326,N_24218);
xor U25928 (N_25928,N_25175,N_24632);
nand U25929 (N_25929,N_24281,N_25171);
nor U25930 (N_25930,N_24705,N_24064);
or U25931 (N_25931,N_24722,N_24928);
and U25932 (N_25932,N_24446,N_24782);
xnor U25933 (N_25933,N_24317,N_24021);
nor U25934 (N_25934,N_24466,N_25057);
or U25935 (N_25935,N_24571,N_24002);
nand U25936 (N_25936,N_24301,N_24368);
xnor U25937 (N_25937,N_24366,N_24990);
and U25938 (N_25938,N_24906,N_24984);
and U25939 (N_25939,N_24772,N_24779);
or U25940 (N_25940,N_24131,N_25022);
xnor U25941 (N_25941,N_24347,N_24799);
and U25942 (N_25942,N_24677,N_24491);
xnor U25943 (N_25943,N_24480,N_24787);
or U25944 (N_25944,N_24897,N_24702);
nor U25945 (N_25945,N_24107,N_25149);
and U25946 (N_25946,N_24362,N_25151);
xor U25947 (N_25947,N_24377,N_24812);
nand U25948 (N_25948,N_24395,N_24049);
nor U25949 (N_25949,N_24884,N_25166);
or U25950 (N_25950,N_24855,N_24550);
or U25951 (N_25951,N_24464,N_24943);
xor U25952 (N_25952,N_24074,N_24130);
nand U25953 (N_25953,N_24822,N_24520);
or U25954 (N_25954,N_25193,N_24445);
nor U25955 (N_25955,N_24679,N_24278);
and U25956 (N_25956,N_24866,N_24916);
nor U25957 (N_25957,N_24204,N_24557);
nor U25958 (N_25958,N_24513,N_24264);
and U25959 (N_25959,N_25187,N_24730);
or U25960 (N_25960,N_24409,N_24607);
and U25961 (N_25961,N_25113,N_24294);
and U25962 (N_25962,N_24210,N_24750);
xnor U25963 (N_25963,N_25085,N_24117);
nand U25964 (N_25964,N_24201,N_25127);
nor U25965 (N_25965,N_25124,N_24443);
xnor U25966 (N_25966,N_24106,N_25135);
or U25967 (N_25967,N_24953,N_24564);
or U25968 (N_25968,N_25023,N_24010);
and U25969 (N_25969,N_24915,N_24306);
xor U25970 (N_25970,N_24479,N_25140);
nor U25971 (N_25971,N_25040,N_24031);
and U25972 (N_25972,N_24214,N_24732);
and U25973 (N_25973,N_24948,N_24515);
and U25974 (N_25974,N_24817,N_25135);
xor U25975 (N_25975,N_24010,N_24522);
xor U25976 (N_25976,N_24917,N_24683);
or U25977 (N_25977,N_24785,N_24708);
nand U25978 (N_25978,N_25034,N_24849);
xnor U25979 (N_25979,N_24315,N_25015);
or U25980 (N_25980,N_24932,N_25137);
nand U25981 (N_25981,N_24267,N_24517);
nand U25982 (N_25982,N_24996,N_24999);
nand U25983 (N_25983,N_24243,N_24773);
nor U25984 (N_25984,N_24844,N_25120);
xnor U25985 (N_25985,N_24566,N_24066);
or U25986 (N_25986,N_24555,N_24518);
xor U25987 (N_25987,N_24155,N_25049);
nand U25988 (N_25988,N_24244,N_24555);
or U25989 (N_25989,N_24086,N_24607);
and U25990 (N_25990,N_24017,N_24987);
nor U25991 (N_25991,N_24099,N_24706);
nor U25992 (N_25992,N_24802,N_24233);
and U25993 (N_25993,N_24157,N_25081);
xnor U25994 (N_25994,N_24134,N_24985);
nand U25995 (N_25995,N_24419,N_24188);
xor U25996 (N_25996,N_24046,N_24540);
xnor U25997 (N_25997,N_24422,N_25145);
nand U25998 (N_25998,N_25179,N_24118);
nand U25999 (N_25999,N_25164,N_24940);
or U26000 (N_26000,N_24974,N_25046);
or U26001 (N_26001,N_25193,N_24996);
nand U26002 (N_26002,N_24118,N_24305);
or U26003 (N_26003,N_24903,N_24485);
and U26004 (N_26004,N_24443,N_24997);
xnor U26005 (N_26005,N_24258,N_24701);
xor U26006 (N_26006,N_24190,N_24318);
nand U26007 (N_26007,N_24976,N_24448);
xor U26008 (N_26008,N_24485,N_24980);
or U26009 (N_26009,N_24009,N_24617);
or U26010 (N_26010,N_24121,N_24877);
xnor U26011 (N_26011,N_24836,N_24598);
or U26012 (N_26012,N_24653,N_24194);
xnor U26013 (N_26013,N_24220,N_25067);
and U26014 (N_26014,N_24110,N_24704);
nand U26015 (N_26015,N_24932,N_24225);
xor U26016 (N_26016,N_24718,N_24732);
nand U26017 (N_26017,N_24054,N_24674);
xnor U26018 (N_26018,N_25065,N_24916);
nor U26019 (N_26019,N_24312,N_24353);
nand U26020 (N_26020,N_24437,N_24349);
nor U26021 (N_26021,N_24655,N_24193);
or U26022 (N_26022,N_25124,N_24116);
xnor U26023 (N_26023,N_24278,N_24399);
xnor U26024 (N_26024,N_24028,N_24572);
nand U26025 (N_26025,N_24401,N_24191);
nor U26026 (N_26026,N_24716,N_25190);
or U26027 (N_26027,N_24120,N_24151);
xnor U26028 (N_26028,N_24621,N_24545);
xnor U26029 (N_26029,N_24495,N_25182);
or U26030 (N_26030,N_24297,N_24619);
nand U26031 (N_26031,N_25035,N_24455);
and U26032 (N_26032,N_24182,N_24457);
nor U26033 (N_26033,N_24503,N_24075);
nand U26034 (N_26034,N_24267,N_24264);
and U26035 (N_26035,N_24048,N_24676);
and U26036 (N_26036,N_25137,N_24315);
or U26037 (N_26037,N_24717,N_24255);
nor U26038 (N_26038,N_24457,N_24866);
and U26039 (N_26039,N_24993,N_24014);
or U26040 (N_26040,N_24326,N_24867);
or U26041 (N_26041,N_24200,N_24987);
nand U26042 (N_26042,N_24416,N_24133);
nand U26043 (N_26043,N_24956,N_24044);
or U26044 (N_26044,N_24897,N_24846);
or U26045 (N_26045,N_25014,N_24893);
or U26046 (N_26046,N_24448,N_24728);
and U26047 (N_26047,N_24974,N_24762);
nor U26048 (N_26048,N_24813,N_25108);
and U26049 (N_26049,N_24531,N_25088);
nand U26050 (N_26050,N_24465,N_24493);
and U26051 (N_26051,N_24205,N_24594);
and U26052 (N_26052,N_24951,N_24033);
and U26053 (N_26053,N_24137,N_24582);
nor U26054 (N_26054,N_25188,N_24070);
nand U26055 (N_26055,N_24490,N_24781);
or U26056 (N_26056,N_24080,N_25126);
xnor U26057 (N_26057,N_24948,N_24120);
or U26058 (N_26058,N_24661,N_24957);
or U26059 (N_26059,N_24005,N_24986);
and U26060 (N_26060,N_24402,N_24101);
nor U26061 (N_26061,N_24264,N_24851);
or U26062 (N_26062,N_24328,N_24308);
xor U26063 (N_26063,N_24279,N_24541);
nor U26064 (N_26064,N_24687,N_24375);
nor U26065 (N_26065,N_24935,N_24625);
xnor U26066 (N_26066,N_24375,N_24335);
nor U26067 (N_26067,N_24363,N_24676);
or U26068 (N_26068,N_24286,N_24772);
xnor U26069 (N_26069,N_25061,N_24297);
nor U26070 (N_26070,N_24006,N_24782);
nor U26071 (N_26071,N_24453,N_24927);
and U26072 (N_26072,N_24555,N_25175);
xor U26073 (N_26073,N_24388,N_24820);
xnor U26074 (N_26074,N_25042,N_24060);
nor U26075 (N_26075,N_24059,N_25109);
and U26076 (N_26076,N_24252,N_24793);
nor U26077 (N_26077,N_24690,N_24413);
xnor U26078 (N_26078,N_24734,N_24627);
xnor U26079 (N_26079,N_24370,N_24949);
nor U26080 (N_26080,N_24524,N_24471);
and U26081 (N_26081,N_24440,N_24203);
or U26082 (N_26082,N_24282,N_25132);
nand U26083 (N_26083,N_24697,N_24928);
xnor U26084 (N_26084,N_24868,N_24517);
nand U26085 (N_26085,N_24167,N_24383);
nor U26086 (N_26086,N_24573,N_24885);
nor U26087 (N_26087,N_24628,N_24622);
and U26088 (N_26088,N_24774,N_24274);
nand U26089 (N_26089,N_24696,N_24543);
nand U26090 (N_26090,N_25165,N_24454);
xor U26091 (N_26091,N_24016,N_25079);
and U26092 (N_26092,N_24889,N_24963);
and U26093 (N_26093,N_25032,N_24283);
xnor U26094 (N_26094,N_24194,N_25030);
nand U26095 (N_26095,N_24261,N_25013);
or U26096 (N_26096,N_24874,N_24480);
nand U26097 (N_26097,N_24847,N_24936);
and U26098 (N_26098,N_24731,N_24821);
and U26099 (N_26099,N_24703,N_24397);
nor U26100 (N_26100,N_24792,N_25173);
xnor U26101 (N_26101,N_24260,N_24695);
xnor U26102 (N_26102,N_24326,N_24997);
nor U26103 (N_26103,N_24816,N_24298);
nand U26104 (N_26104,N_24102,N_24198);
nand U26105 (N_26105,N_25073,N_24685);
xnor U26106 (N_26106,N_24749,N_24949);
nor U26107 (N_26107,N_24115,N_24933);
xnor U26108 (N_26108,N_24924,N_24441);
or U26109 (N_26109,N_24759,N_24392);
nand U26110 (N_26110,N_24691,N_24183);
nand U26111 (N_26111,N_24929,N_25029);
nor U26112 (N_26112,N_24666,N_24759);
or U26113 (N_26113,N_24366,N_24821);
or U26114 (N_26114,N_24228,N_24445);
nor U26115 (N_26115,N_25000,N_24591);
nand U26116 (N_26116,N_24041,N_25171);
nand U26117 (N_26117,N_24209,N_24109);
and U26118 (N_26118,N_24606,N_24093);
xor U26119 (N_26119,N_24931,N_24463);
nand U26120 (N_26120,N_24360,N_24482);
xnor U26121 (N_26121,N_25194,N_24920);
nor U26122 (N_26122,N_24779,N_25108);
nor U26123 (N_26123,N_24353,N_24761);
and U26124 (N_26124,N_24478,N_24711);
xnor U26125 (N_26125,N_24368,N_25047);
nor U26126 (N_26126,N_24038,N_24750);
nor U26127 (N_26127,N_24338,N_24265);
xor U26128 (N_26128,N_24141,N_24626);
or U26129 (N_26129,N_24145,N_24631);
nand U26130 (N_26130,N_24731,N_24213);
or U26131 (N_26131,N_24836,N_24708);
xnor U26132 (N_26132,N_24604,N_24325);
xor U26133 (N_26133,N_24932,N_24152);
nand U26134 (N_26134,N_24130,N_24360);
or U26135 (N_26135,N_25113,N_24210);
nand U26136 (N_26136,N_24192,N_25019);
nand U26137 (N_26137,N_24425,N_24358);
or U26138 (N_26138,N_24571,N_24589);
nand U26139 (N_26139,N_24414,N_25105);
nor U26140 (N_26140,N_24202,N_24820);
or U26141 (N_26141,N_24757,N_24747);
xor U26142 (N_26142,N_24148,N_24502);
or U26143 (N_26143,N_24288,N_24155);
nand U26144 (N_26144,N_24618,N_24821);
nand U26145 (N_26145,N_24662,N_24754);
or U26146 (N_26146,N_24017,N_24540);
nor U26147 (N_26147,N_24978,N_24326);
nand U26148 (N_26148,N_24191,N_24792);
or U26149 (N_26149,N_24344,N_24561);
xnor U26150 (N_26150,N_24277,N_24084);
or U26151 (N_26151,N_25014,N_24083);
or U26152 (N_26152,N_24381,N_24288);
nor U26153 (N_26153,N_24176,N_24061);
nand U26154 (N_26154,N_24817,N_24811);
nor U26155 (N_26155,N_24965,N_24940);
or U26156 (N_26156,N_24515,N_24392);
nor U26157 (N_26157,N_24702,N_24917);
and U26158 (N_26158,N_24789,N_24521);
and U26159 (N_26159,N_24175,N_24975);
nor U26160 (N_26160,N_24113,N_25050);
and U26161 (N_26161,N_24888,N_24621);
xnor U26162 (N_26162,N_24825,N_24082);
and U26163 (N_26163,N_25050,N_24919);
or U26164 (N_26164,N_25058,N_25198);
or U26165 (N_26165,N_24508,N_24631);
nand U26166 (N_26166,N_24652,N_24306);
nor U26167 (N_26167,N_25094,N_25149);
xor U26168 (N_26168,N_24248,N_24201);
and U26169 (N_26169,N_24709,N_24367);
or U26170 (N_26170,N_24067,N_24995);
nor U26171 (N_26171,N_24531,N_24789);
nor U26172 (N_26172,N_25169,N_24521);
or U26173 (N_26173,N_24349,N_25068);
or U26174 (N_26174,N_24994,N_24992);
xnor U26175 (N_26175,N_25178,N_24186);
nand U26176 (N_26176,N_24013,N_24043);
nand U26177 (N_26177,N_25072,N_24123);
xnor U26178 (N_26178,N_24267,N_24810);
xor U26179 (N_26179,N_24423,N_24500);
nand U26180 (N_26180,N_24655,N_24480);
xor U26181 (N_26181,N_24476,N_24868);
nand U26182 (N_26182,N_24194,N_25169);
xor U26183 (N_26183,N_24404,N_25077);
and U26184 (N_26184,N_24289,N_24925);
nand U26185 (N_26185,N_24521,N_24932);
and U26186 (N_26186,N_24897,N_24142);
or U26187 (N_26187,N_25175,N_24239);
xor U26188 (N_26188,N_24795,N_25087);
nor U26189 (N_26189,N_24390,N_24694);
nand U26190 (N_26190,N_24701,N_24952);
xnor U26191 (N_26191,N_24987,N_24985);
nor U26192 (N_26192,N_24413,N_24858);
nor U26193 (N_26193,N_24689,N_24391);
nand U26194 (N_26194,N_24741,N_24058);
or U26195 (N_26195,N_24585,N_24264);
or U26196 (N_26196,N_24574,N_25067);
or U26197 (N_26197,N_24755,N_24098);
nor U26198 (N_26198,N_24056,N_25060);
xnor U26199 (N_26199,N_24070,N_24552);
xor U26200 (N_26200,N_24171,N_24830);
nand U26201 (N_26201,N_24067,N_25042);
xnor U26202 (N_26202,N_24954,N_25098);
xnor U26203 (N_26203,N_24944,N_24510);
nor U26204 (N_26204,N_24417,N_25191);
or U26205 (N_26205,N_24555,N_24615);
nor U26206 (N_26206,N_24698,N_24087);
nor U26207 (N_26207,N_25074,N_24155);
nand U26208 (N_26208,N_24985,N_24386);
xor U26209 (N_26209,N_25052,N_24563);
nor U26210 (N_26210,N_24430,N_24652);
nand U26211 (N_26211,N_24942,N_24570);
nor U26212 (N_26212,N_24416,N_24380);
and U26213 (N_26213,N_24291,N_24679);
or U26214 (N_26214,N_24132,N_24577);
or U26215 (N_26215,N_24656,N_25169);
and U26216 (N_26216,N_24230,N_24103);
and U26217 (N_26217,N_24718,N_24636);
xor U26218 (N_26218,N_24387,N_25077);
nand U26219 (N_26219,N_24323,N_24890);
nor U26220 (N_26220,N_24286,N_24599);
or U26221 (N_26221,N_24149,N_24715);
xor U26222 (N_26222,N_24143,N_24987);
or U26223 (N_26223,N_24690,N_24786);
or U26224 (N_26224,N_24682,N_24073);
nand U26225 (N_26225,N_24902,N_25101);
and U26226 (N_26226,N_24822,N_24014);
nand U26227 (N_26227,N_25130,N_25147);
or U26228 (N_26228,N_24691,N_25126);
xnor U26229 (N_26229,N_24994,N_24894);
nor U26230 (N_26230,N_24935,N_24843);
and U26231 (N_26231,N_24563,N_24579);
xor U26232 (N_26232,N_25127,N_24743);
and U26233 (N_26233,N_24186,N_24254);
xor U26234 (N_26234,N_24952,N_24617);
xnor U26235 (N_26235,N_24708,N_24446);
and U26236 (N_26236,N_24485,N_24535);
nand U26237 (N_26237,N_24843,N_24735);
nor U26238 (N_26238,N_24860,N_24645);
or U26239 (N_26239,N_24571,N_24957);
nand U26240 (N_26240,N_24232,N_24359);
and U26241 (N_26241,N_24675,N_25129);
xor U26242 (N_26242,N_24479,N_24139);
or U26243 (N_26243,N_24187,N_24574);
nand U26244 (N_26244,N_25154,N_24294);
or U26245 (N_26245,N_24564,N_24159);
or U26246 (N_26246,N_24158,N_24658);
or U26247 (N_26247,N_24306,N_24773);
or U26248 (N_26248,N_24544,N_25069);
xnor U26249 (N_26249,N_24207,N_24321);
nor U26250 (N_26250,N_24153,N_24464);
and U26251 (N_26251,N_25073,N_25174);
nor U26252 (N_26252,N_24757,N_24733);
nor U26253 (N_26253,N_24636,N_24993);
and U26254 (N_26254,N_24143,N_24895);
nor U26255 (N_26255,N_24651,N_24789);
xor U26256 (N_26256,N_24572,N_25141);
nor U26257 (N_26257,N_24622,N_24144);
xor U26258 (N_26258,N_24378,N_24637);
xor U26259 (N_26259,N_24286,N_24111);
and U26260 (N_26260,N_24236,N_24921);
nor U26261 (N_26261,N_24083,N_24484);
or U26262 (N_26262,N_24497,N_24819);
nand U26263 (N_26263,N_24710,N_24164);
nor U26264 (N_26264,N_24346,N_24906);
nand U26265 (N_26265,N_24723,N_24983);
nand U26266 (N_26266,N_24637,N_25134);
nand U26267 (N_26267,N_24365,N_25067);
or U26268 (N_26268,N_24030,N_24413);
nand U26269 (N_26269,N_24480,N_24070);
and U26270 (N_26270,N_24445,N_24913);
or U26271 (N_26271,N_24290,N_24043);
nand U26272 (N_26272,N_24904,N_24530);
xor U26273 (N_26273,N_24891,N_24995);
xnor U26274 (N_26274,N_24624,N_24817);
nand U26275 (N_26275,N_24917,N_24092);
nand U26276 (N_26276,N_24341,N_24213);
xnor U26277 (N_26277,N_24002,N_24623);
nor U26278 (N_26278,N_24763,N_24287);
and U26279 (N_26279,N_24711,N_24293);
or U26280 (N_26280,N_24437,N_25027);
and U26281 (N_26281,N_25099,N_24567);
nand U26282 (N_26282,N_24992,N_24152);
xnor U26283 (N_26283,N_24864,N_25178);
or U26284 (N_26284,N_24192,N_25078);
nor U26285 (N_26285,N_24953,N_25111);
nand U26286 (N_26286,N_24960,N_24336);
xor U26287 (N_26287,N_24457,N_24322);
and U26288 (N_26288,N_24511,N_24274);
and U26289 (N_26289,N_24241,N_25087);
or U26290 (N_26290,N_24183,N_24212);
and U26291 (N_26291,N_24120,N_24144);
and U26292 (N_26292,N_25102,N_24091);
and U26293 (N_26293,N_24824,N_25110);
or U26294 (N_26294,N_24706,N_24428);
xor U26295 (N_26295,N_24824,N_24464);
xor U26296 (N_26296,N_24408,N_24848);
xnor U26297 (N_26297,N_24668,N_24347);
nor U26298 (N_26298,N_25038,N_25069);
and U26299 (N_26299,N_24521,N_24304);
nand U26300 (N_26300,N_24063,N_24447);
nor U26301 (N_26301,N_24369,N_24162);
or U26302 (N_26302,N_25063,N_24597);
nor U26303 (N_26303,N_25127,N_24790);
or U26304 (N_26304,N_24223,N_24481);
and U26305 (N_26305,N_24678,N_24554);
and U26306 (N_26306,N_24415,N_25001);
and U26307 (N_26307,N_24831,N_24211);
nand U26308 (N_26308,N_24513,N_25166);
xnor U26309 (N_26309,N_24673,N_24753);
xor U26310 (N_26310,N_24679,N_24758);
or U26311 (N_26311,N_24199,N_24580);
nand U26312 (N_26312,N_24416,N_25159);
nand U26313 (N_26313,N_24396,N_24997);
or U26314 (N_26314,N_24620,N_25012);
and U26315 (N_26315,N_24238,N_24757);
or U26316 (N_26316,N_24811,N_24511);
or U26317 (N_26317,N_25139,N_24556);
or U26318 (N_26318,N_24552,N_24259);
or U26319 (N_26319,N_24953,N_25009);
nand U26320 (N_26320,N_24123,N_24079);
nor U26321 (N_26321,N_24672,N_24538);
and U26322 (N_26322,N_25184,N_24412);
or U26323 (N_26323,N_24194,N_25173);
nor U26324 (N_26324,N_25064,N_24214);
and U26325 (N_26325,N_24719,N_24636);
and U26326 (N_26326,N_25050,N_24116);
nand U26327 (N_26327,N_24565,N_25175);
xor U26328 (N_26328,N_24367,N_24855);
xor U26329 (N_26329,N_25051,N_24518);
xor U26330 (N_26330,N_25066,N_24313);
or U26331 (N_26331,N_24493,N_24451);
or U26332 (N_26332,N_24209,N_24776);
xor U26333 (N_26333,N_24240,N_24843);
and U26334 (N_26334,N_24786,N_24925);
and U26335 (N_26335,N_24014,N_24618);
or U26336 (N_26336,N_24897,N_24783);
xor U26337 (N_26337,N_24565,N_25053);
or U26338 (N_26338,N_24128,N_24123);
nand U26339 (N_26339,N_24509,N_24881);
xnor U26340 (N_26340,N_24625,N_25009);
or U26341 (N_26341,N_24646,N_24401);
nor U26342 (N_26342,N_24491,N_24493);
xor U26343 (N_26343,N_25024,N_24476);
xor U26344 (N_26344,N_25145,N_24745);
and U26345 (N_26345,N_24342,N_24678);
nand U26346 (N_26346,N_24295,N_24754);
and U26347 (N_26347,N_24611,N_24013);
and U26348 (N_26348,N_24182,N_24754);
nor U26349 (N_26349,N_24328,N_24116);
nor U26350 (N_26350,N_24260,N_24425);
nor U26351 (N_26351,N_24560,N_25184);
nand U26352 (N_26352,N_24931,N_24015);
nand U26353 (N_26353,N_24629,N_24793);
or U26354 (N_26354,N_24110,N_24113);
nor U26355 (N_26355,N_24928,N_25135);
nor U26356 (N_26356,N_25076,N_24682);
and U26357 (N_26357,N_24266,N_25021);
and U26358 (N_26358,N_24559,N_24892);
or U26359 (N_26359,N_24882,N_24342);
xnor U26360 (N_26360,N_24108,N_25089);
xor U26361 (N_26361,N_24234,N_24406);
and U26362 (N_26362,N_24407,N_24592);
xor U26363 (N_26363,N_24834,N_24532);
nor U26364 (N_26364,N_24678,N_24067);
and U26365 (N_26365,N_24109,N_25006);
nand U26366 (N_26366,N_24459,N_24922);
or U26367 (N_26367,N_24730,N_24351);
and U26368 (N_26368,N_25023,N_25063);
nor U26369 (N_26369,N_24167,N_24864);
nor U26370 (N_26370,N_24793,N_24082);
and U26371 (N_26371,N_24764,N_24056);
or U26372 (N_26372,N_24048,N_24569);
xnor U26373 (N_26373,N_24858,N_24855);
xnor U26374 (N_26374,N_24372,N_24217);
xor U26375 (N_26375,N_24040,N_25169);
nor U26376 (N_26376,N_24170,N_24068);
or U26377 (N_26377,N_24915,N_25124);
and U26378 (N_26378,N_24583,N_24503);
nand U26379 (N_26379,N_24425,N_25096);
nand U26380 (N_26380,N_24988,N_25080);
or U26381 (N_26381,N_24117,N_24729);
nand U26382 (N_26382,N_24594,N_24494);
and U26383 (N_26383,N_24525,N_25082);
nand U26384 (N_26384,N_24955,N_24787);
xor U26385 (N_26385,N_24459,N_24612);
nand U26386 (N_26386,N_24182,N_24440);
nor U26387 (N_26387,N_24798,N_25172);
and U26388 (N_26388,N_25194,N_25106);
nand U26389 (N_26389,N_24144,N_25040);
and U26390 (N_26390,N_24067,N_24892);
and U26391 (N_26391,N_24094,N_24092);
and U26392 (N_26392,N_25116,N_24939);
nor U26393 (N_26393,N_24524,N_24065);
nor U26394 (N_26394,N_24423,N_24509);
nor U26395 (N_26395,N_24773,N_25147);
and U26396 (N_26396,N_24382,N_24889);
or U26397 (N_26397,N_24831,N_24565);
nand U26398 (N_26398,N_24561,N_24130);
nor U26399 (N_26399,N_24658,N_24623);
nor U26400 (N_26400,N_26066,N_26377);
nor U26401 (N_26401,N_25807,N_25719);
xnor U26402 (N_26402,N_25291,N_26269);
and U26403 (N_26403,N_25588,N_25279);
nand U26404 (N_26404,N_26178,N_25322);
xnor U26405 (N_26405,N_26232,N_25312);
and U26406 (N_26406,N_25419,N_25288);
or U26407 (N_26407,N_25367,N_25543);
nor U26408 (N_26408,N_25989,N_25800);
nand U26409 (N_26409,N_25804,N_26194);
or U26410 (N_26410,N_25587,N_25517);
nor U26411 (N_26411,N_25942,N_25349);
or U26412 (N_26412,N_25230,N_25325);
and U26413 (N_26413,N_25846,N_25458);
nand U26414 (N_26414,N_25764,N_26349);
nand U26415 (N_26415,N_25902,N_25286);
xor U26416 (N_26416,N_26311,N_26216);
nor U26417 (N_26417,N_25865,N_25538);
nor U26418 (N_26418,N_25690,N_25614);
nor U26419 (N_26419,N_25631,N_25997);
nand U26420 (N_26420,N_25969,N_26204);
or U26421 (N_26421,N_25555,N_26354);
or U26422 (N_26422,N_25248,N_25472);
and U26423 (N_26423,N_25670,N_25818);
nor U26424 (N_26424,N_26372,N_25966);
and U26425 (N_26425,N_25316,N_25999);
or U26426 (N_26426,N_26367,N_26389);
and U26427 (N_26427,N_25205,N_26391);
nor U26428 (N_26428,N_25988,N_25730);
xnor U26429 (N_26429,N_25598,N_26081);
xnor U26430 (N_26430,N_25605,N_25787);
xnor U26431 (N_26431,N_25431,N_26057);
xnor U26432 (N_26432,N_26308,N_26225);
nand U26433 (N_26433,N_25695,N_26370);
nand U26434 (N_26434,N_25613,N_25998);
and U26435 (N_26435,N_25811,N_25772);
xnor U26436 (N_26436,N_25739,N_25806);
nand U26437 (N_26437,N_25977,N_26340);
and U26438 (N_26438,N_25218,N_25845);
xnor U26439 (N_26439,N_25823,N_25584);
nor U26440 (N_26440,N_26338,N_25246);
nor U26441 (N_26441,N_25812,N_25825);
or U26442 (N_26442,N_25888,N_26380);
or U26443 (N_26443,N_26016,N_25450);
nor U26444 (N_26444,N_25463,N_25677);
xnor U26445 (N_26445,N_25401,N_25925);
xnor U26446 (N_26446,N_26227,N_26385);
nor U26447 (N_26447,N_25426,N_26241);
and U26448 (N_26448,N_25526,N_25896);
nor U26449 (N_26449,N_26257,N_25630);
nor U26450 (N_26450,N_26063,N_25547);
xnor U26451 (N_26451,N_25870,N_25652);
and U26452 (N_26452,N_25382,N_25849);
or U26453 (N_26453,N_25669,N_26327);
or U26454 (N_26454,N_25619,N_25601);
xor U26455 (N_26455,N_25241,N_25898);
xor U26456 (N_26456,N_26160,N_25485);
or U26457 (N_26457,N_25792,N_25892);
xor U26458 (N_26458,N_25894,N_25329);
or U26459 (N_26459,N_25817,N_25257);
nor U26460 (N_26460,N_25374,N_25226);
and U26461 (N_26461,N_25834,N_25227);
nand U26462 (N_26462,N_25891,N_26076);
or U26463 (N_26463,N_26215,N_26127);
nor U26464 (N_26464,N_26201,N_26210);
xor U26465 (N_26465,N_26369,N_25466);
or U26466 (N_26466,N_25498,N_26271);
nand U26467 (N_26467,N_25737,N_26398);
or U26468 (N_26468,N_25213,N_25990);
xor U26469 (N_26469,N_25317,N_25810);
nand U26470 (N_26470,N_26067,N_25581);
nor U26471 (N_26471,N_25635,N_26299);
or U26472 (N_26472,N_26009,N_25250);
or U26473 (N_26473,N_25831,N_26285);
xor U26474 (N_26474,N_25369,N_25343);
or U26475 (N_26475,N_25913,N_25955);
xnor U26476 (N_26476,N_26310,N_26283);
nor U26477 (N_26477,N_25909,N_25615);
and U26478 (N_26478,N_26314,N_25713);
or U26479 (N_26479,N_25394,N_26119);
nand U26480 (N_26480,N_26136,N_26366);
and U26481 (N_26481,N_25822,N_25916);
xnor U26482 (N_26482,N_26267,N_25646);
nor U26483 (N_26483,N_26021,N_25596);
and U26484 (N_26484,N_25599,N_25327);
nor U26485 (N_26485,N_25741,N_26237);
nand U26486 (N_26486,N_25774,N_26234);
nand U26487 (N_26487,N_25956,N_25788);
or U26488 (N_26488,N_25287,N_25697);
nor U26489 (N_26489,N_25272,N_25769);
and U26490 (N_26490,N_25465,N_25520);
and U26491 (N_26491,N_25621,N_25360);
nand U26492 (N_26492,N_25524,N_26280);
and U26493 (N_26493,N_25964,N_26233);
xor U26494 (N_26494,N_25427,N_25848);
nand U26495 (N_26495,N_26382,N_25840);
nor U26496 (N_26496,N_25500,N_25239);
nor U26497 (N_26497,N_26182,N_25400);
or U26498 (N_26498,N_25981,N_26022);
nor U26499 (N_26499,N_26296,N_25662);
nor U26500 (N_26500,N_25324,N_26006);
nor U26501 (N_26501,N_25667,N_25345);
xor U26502 (N_26502,N_26064,N_26036);
or U26503 (N_26503,N_25391,N_25968);
and U26504 (N_26504,N_26074,N_25654);
or U26505 (N_26505,N_26352,N_25928);
or U26506 (N_26506,N_26272,N_25771);
nand U26507 (N_26507,N_25686,N_26120);
xor U26508 (N_26508,N_25820,N_26360);
nand U26509 (N_26509,N_25930,N_26281);
or U26510 (N_26510,N_25918,N_25970);
nor U26511 (N_26511,N_25885,N_25442);
and U26512 (N_26512,N_25805,N_26348);
nor U26513 (N_26513,N_25573,N_25236);
nand U26514 (N_26514,N_25882,N_25570);
and U26515 (N_26515,N_26094,N_25304);
xnor U26516 (N_26516,N_25333,N_26023);
nor U26517 (N_26517,N_25815,N_26019);
xnor U26518 (N_26518,N_26174,N_26350);
nand U26519 (N_26519,N_25347,N_26202);
xor U26520 (N_26520,N_25362,N_25574);
and U26521 (N_26521,N_25430,N_25684);
xor U26522 (N_26522,N_25577,N_26316);
nor U26523 (N_26523,N_25734,N_25864);
nor U26524 (N_26524,N_26060,N_25782);
or U26525 (N_26525,N_26167,N_26291);
nand U26526 (N_26526,N_26042,N_26219);
xnor U26527 (N_26527,N_26214,N_25600);
or U26528 (N_26528,N_25611,N_25486);
and U26529 (N_26529,N_25532,N_26293);
xnor U26530 (N_26530,N_25490,N_25277);
or U26531 (N_26531,N_25428,N_26115);
or U26532 (N_26532,N_26325,N_25844);
xnor U26533 (N_26533,N_26087,N_25244);
xnor U26534 (N_26534,N_26286,N_25664);
nand U26535 (N_26535,N_25379,N_25773);
and U26536 (N_26536,N_25617,N_25854);
xnor U26537 (N_26537,N_25853,N_25872);
and U26538 (N_26538,N_26289,N_25414);
nand U26539 (N_26539,N_26231,N_26034);
or U26540 (N_26540,N_25960,N_25623);
and U26541 (N_26541,N_25412,N_26331);
or U26542 (N_26542,N_25560,N_25328);
nor U26543 (N_26543,N_25273,N_26361);
or U26544 (N_26544,N_26169,N_26079);
or U26545 (N_26545,N_25991,N_25957);
nand U26546 (N_26546,N_26328,N_25627);
or U26547 (N_26547,N_26149,N_25881);
and U26548 (N_26548,N_25386,N_25476);
and U26549 (N_26549,N_25985,N_25473);
xnor U26550 (N_26550,N_26362,N_25732);
xnor U26551 (N_26551,N_26154,N_26018);
nand U26552 (N_26552,N_25309,N_25559);
xor U26553 (N_26553,N_25456,N_25280);
nand U26554 (N_26554,N_25220,N_26224);
xor U26555 (N_26555,N_26085,N_26309);
nor U26556 (N_26556,N_26374,N_25571);
nor U26557 (N_26557,N_26226,N_26083);
or U26558 (N_26558,N_25266,N_25487);
nand U26559 (N_26559,N_25833,N_25721);
nor U26560 (N_26560,N_26254,N_25206);
xor U26561 (N_26561,N_26105,N_25278);
xor U26562 (N_26562,N_26108,N_25945);
nand U26563 (N_26563,N_25434,N_26275);
or U26564 (N_26564,N_26193,N_25384);
xor U26565 (N_26565,N_25668,N_26270);
xnor U26566 (N_26566,N_26199,N_25780);
and U26567 (N_26567,N_25620,N_25504);
xnor U26568 (N_26568,N_26103,N_25828);
xor U26569 (N_26569,N_25261,N_26242);
or U26570 (N_26570,N_25331,N_26159);
nor U26571 (N_26571,N_25380,N_25424);
or U26572 (N_26572,N_25422,N_25665);
nor U26573 (N_26573,N_25460,N_25535);
or U26574 (N_26574,N_25726,N_25565);
xor U26575 (N_26575,N_26134,N_25582);
xor U26576 (N_26576,N_25508,N_25529);
nand U26577 (N_26577,N_26040,N_25742);
and U26578 (N_26578,N_25269,N_25728);
or U26579 (N_26579,N_26097,N_25372);
nor U26580 (N_26580,N_26260,N_25495);
and U26581 (N_26581,N_26046,N_25980);
nand U26582 (N_26582,N_25501,N_25377);
nor U26583 (N_26583,N_25222,N_26185);
or U26584 (N_26584,N_25941,N_26013);
and U26585 (N_26585,N_25260,N_25553);
nor U26586 (N_26586,N_25685,N_25900);
nand U26587 (N_26587,N_25461,N_25709);
and U26588 (N_26588,N_25202,N_25784);
nand U26589 (N_26589,N_25363,N_25311);
or U26590 (N_26590,N_25489,N_25416);
or U26591 (N_26591,N_26157,N_26138);
or U26592 (N_26592,N_25642,N_25542);
nor U26593 (N_26593,N_25539,N_25357);
xor U26594 (N_26594,N_25418,N_25994);
nor U26595 (N_26595,N_25440,N_26171);
nand U26596 (N_26596,N_25284,N_25392);
and U26597 (N_26597,N_25403,N_25704);
nand U26598 (N_26598,N_25975,N_26161);
nor U26599 (N_26599,N_25908,N_25245);
and U26600 (N_26600,N_25264,N_26276);
and U26601 (N_26601,N_26106,N_25733);
xor U26602 (N_26602,N_25449,N_25231);
nand U26603 (N_26603,N_25758,N_25455);
and U26604 (N_26604,N_26323,N_26033);
nor U26605 (N_26605,N_25626,N_26287);
xor U26606 (N_26606,N_26277,N_25874);
xor U26607 (N_26607,N_25549,N_26062);
and U26608 (N_26608,N_26306,N_25335);
xnor U26609 (N_26609,N_25711,N_26353);
xor U26610 (N_26610,N_25203,N_26025);
nand U26611 (N_26611,N_25415,N_26107);
nor U26612 (N_26612,N_26304,N_25338);
nor U26613 (N_26613,N_26326,N_25358);
or U26614 (N_26614,N_25658,N_25683);
nand U26615 (N_26615,N_25289,N_26315);
or U26616 (N_26616,N_25656,N_26031);
nor U26617 (N_26617,N_25779,N_25629);
xnor U26618 (N_26618,N_26121,N_25432);
nand U26619 (N_26619,N_25373,N_25612);
and U26620 (N_26620,N_25447,N_25454);
xor U26621 (N_26621,N_26387,N_25212);
and U26622 (N_26622,N_25527,N_26086);
or U26623 (N_26623,N_26004,N_25491);
and U26624 (N_26624,N_26320,N_25562);
nor U26625 (N_26625,N_25344,N_25361);
nor U26626 (N_26626,N_26187,N_25748);
nand U26627 (N_26627,N_26200,N_25306);
nand U26628 (N_26628,N_25963,N_26313);
nand U26629 (N_26629,N_26239,N_25936);
nor U26630 (N_26630,N_25798,N_26262);
and U26631 (N_26631,N_26152,N_25469);
and U26632 (N_26632,N_26162,N_26395);
nor U26633 (N_26633,N_25420,N_25735);
and U26634 (N_26634,N_26029,N_25947);
or U26635 (N_26635,N_26295,N_25271);
xor U26636 (N_26636,N_25481,N_26365);
xnor U26637 (N_26637,N_25672,N_26051);
nand U26638 (N_26638,N_25330,N_26118);
or U26639 (N_26639,N_26045,N_25754);
nand U26640 (N_26640,N_26123,N_25567);
nand U26641 (N_26641,N_25568,N_25483);
and U26642 (N_26642,N_25267,N_25767);
nand U26643 (N_26643,N_25521,N_25350);
xnor U26644 (N_26644,N_26091,N_25889);
or U26645 (N_26645,N_25351,N_25640);
nand U26646 (N_26646,N_25530,N_26339);
or U26647 (N_26647,N_25710,N_25240);
or U26648 (N_26648,N_25839,N_25750);
nand U26649 (N_26649,N_26388,N_26026);
or U26650 (N_26650,N_25776,N_25905);
nand U26651 (N_26651,N_26396,N_25786);
or U26652 (N_26652,N_25857,N_26212);
nor U26653 (N_26653,N_26071,N_25283);
xor U26654 (N_26654,N_25301,N_26122);
nand U26655 (N_26655,N_26346,N_25698);
nand U26656 (N_26656,N_25842,N_26132);
or U26657 (N_26657,N_25318,N_25768);
nor U26658 (N_26658,N_25356,N_25211);
nor U26659 (N_26659,N_26273,N_25216);
xor U26660 (N_26660,N_25474,N_26264);
xnor U26661 (N_26661,N_25247,N_25649);
or U26662 (N_26662,N_26052,N_26243);
nand U26663 (N_26663,N_26302,N_26392);
nand U26664 (N_26664,N_25932,N_26318);
nor U26665 (N_26665,N_25224,N_26125);
xor U26666 (N_26666,N_25421,N_25228);
and U26667 (N_26667,N_25877,N_25855);
xor U26668 (N_26668,N_26049,N_26165);
xor U26669 (N_26669,N_26355,N_25838);
nor U26670 (N_26670,N_25973,N_26082);
or U26671 (N_26671,N_25528,N_26142);
nand U26672 (N_26672,N_25545,N_25893);
or U26673 (N_26673,N_26113,N_25883);
xnor U26674 (N_26674,N_25408,N_26324);
and U26675 (N_26675,N_26180,N_25441);
and U26676 (N_26676,N_25225,N_25340);
nor U26677 (N_26677,N_26363,N_25799);
or U26678 (N_26678,N_25402,N_26061);
xor U26679 (N_26679,N_25836,N_25869);
or U26680 (N_26680,N_26027,N_26196);
or U26681 (N_26681,N_26047,N_25609);
nor U26682 (N_26682,N_26069,N_25861);
nor U26683 (N_26683,N_26096,N_25731);
and U26684 (N_26684,N_26351,N_25992);
nand U26685 (N_26685,N_25355,N_25544);
nand U26686 (N_26686,N_25346,N_25715);
xor U26687 (N_26687,N_25365,N_26141);
and U26688 (N_26688,N_25931,N_25850);
nand U26689 (N_26689,N_25866,N_25912);
and U26690 (N_26690,N_25569,N_25636);
or U26691 (N_26691,N_26189,N_25860);
and U26692 (N_26692,N_25515,N_25593);
or U26693 (N_26693,N_26209,N_25702);
or U26694 (N_26694,N_26028,N_25717);
xnor U26695 (N_26695,N_26101,N_25759);
and U26696 (N_26696,N_26333,N_25522);
nand U26697 (N_26697,N_26104,N_25478);
nor U26698 (N_26698,N_25298,N_25911);
or U26699 (N_26699,N_26386,N_25607);
and U26700 (N_26700,N_25681,N_25645);
and U26701 (N_26701,N_26203,N_25464);
xor U26702 (N_26702,N_25778,N_26336);
xnor U26703 (N_26703,N_25313,N_25540);
or U26704 (N_26704,N_25755,N_25701);
xnor U26705 (N_26705,N_25659,N_26089);
xnor U26706 (N_26706,N_25972,N_25761);
and U26707 (N_26707,N_25687,N_25935);
nor U26708 (N_26708,N_25680,N_25796);
or U26709 (N_26709,N_25274,N_25661);
xnor U26710 (N_26710,N_25534,N_25655);
or U26711 (N_26711,N_25319,N_26130);
nand U26712 (N_26712,N_26394,N_25740);
nor U26713 (N_26713,N_25906,N_25305);
nand U26714 (N_26714,N_25310,N_25604);
nor U26715 (N_26715,N_26190,N_25830);
nor U26716 (N_26716,N_25747,N_25622);
nand U26717 (N_26717,N_25376,N_26117);
nor U26718 (N_26718,N_25953,N_25899);
and U26719 (N_26719,N_25923,N_26256);
and U26720 (N_26720,N_25252,N_25411);
nand U26721 (N_26721,N_25359,N_26146);
nor U26722 (N_26722,N_25725,N_25497);
nand U26723 (N_26723,N_25480,N_26073);
or U26724 (N_26724,N_25585,N_25897);
and U26725 (N_26725,N_25858,N_25675);
nor U26726 (N_26726,N_26017,N_26265);
and U26727 (N_26727,N_25462,N_25457);
nand U26728 (N_26728,N_25390,N_26223);
nand U26729 (N_26729,N_25890,N_25643);
nor U26730 (N_26730,N_26173,N_25868);
or U26731 (N_26731,N_26059,N_25751);
xor U26732 (N_26732,N_25647,N_25689);
nor U26733 (N_26733,N_25965,N_26359);
and U26734 (N_26734,N_25275,N_25723);
nor U26735 (N_26735,N_25215,N_25297);
nor U26736 (N_26736,N_25378,N_25207);
or U26737 (N_26737,N_26221,N_25259);
and U26738 (N_26738,N_25907,N_26246);
nor U26739 (N_26739,N_26095,N_25949);
xnor U26740 (N_26740,N_26288,N_26156);
and U26741 (N_26741,N_26211,N_25803);
nand U26742 (N_26742,N_25494,N_26010);
nor U26743 (N_26743,N_25837,N_26005);
xor U26744 (N_26744,N_25597,N_25639);
nand U26745 (N_26745,N_25509,N_25625);
and U26746 (N_26746,N_25948,N_26344);
or U26747 (N_26747,N_25694,N_26112);
nand U26748 (N_26748,N_25586,N_25375);
and U26749 (N_26749,N_25499,N_25398);
or U26750 (N_26750,N_25475,N_26100);
nor U26751 (N_26751,N_25789,N_25393);
xnor U26752 (N_26752,N_26139,N_25299);
and U26753 (N_26753,N_25663,N_25887);
or U26754 (N_26754,N_25255,N_26150);
nand U26755 (N_26755,N_26218,N_26321);
nand U26756 (N_26756,N_25221,N_26206);
and U26757 (N_26757,N_25282,N_25952);
nor U26758 (N_26758,N_25632,N_25433);
xnor U26759 (N_26759,N_26056,N_25303);
xnor U26760 (N_26760,N_26102,N_25589);
or U26761 (N_26761,N_25700,N_25342);
xor U26762 (N_26762,N_25841,N_26249);
nor U26763 (N_26763,N_25525,N_25962);
and U26764 (N_26764,N_25429,N_26259);
xnor U26765 (N_26765,N_25405,N_25813);
nand U26766 (N_26766,N_25753,N_25691);
nor U26767 (N_26767,N_26038,N_25396);
and U26768 (N_26768,N_26261,N_25856);
or U26769 (N_26769,N_25939,N_25832);
nand U26770 (N_26770,N_26368,N_26084);
nand U26771 (N_26771,N_25785,N_25388);
and U26772 (N_26772,N_26222,N_25482);
or U26773 (N_26773,N_26000,N_26217);
nor U26774 (N_26774,N_26020,N_26250);
nand U26775 (N_26775,N_26114,N_26168);
xor U26776 (N_26776,N_25638,N_26172);
or U26777 (N_26777,N_26303,N_26044);
and U26778 (N_26778,N_25917,N_26191);
nor U26779 (N_26779,N_25666,N_25413);
xnor U26780 (N_26780,N_25924,N_26305);
and U26781 (N_26781,N_25707,N_25219);
or U26782 (N_26782,N_25852,N_25556);
or U26783 (N_26783,N_25682,N_26133);
nor U26784 (N_26784,N_25699,N_25334);
xnor U26785 (N_26785,N_25467,N_25518);
nand U26786 (N_26786,N_25519,N_25943);
and U26787 (N_26787,N_26247,N_25443);
or U26788 (N_26788,N_26379,N_25703);
and U26789 (N_26789,N_25763,N_25976);
nor U26790 (N_26790,N_25903,N_25802);
xor U26791 (N_26791,N_25348,N_26307);
nor U26792 (N_26792,N_25337,N_26177);
nand U26793 (N_26793,N_25503,N_25404);
nand U26794 (N_26794,N_25204,N_25738);
nand U26795 (N_26795,N_26183,N_25961);
nand U26796 (N_26796,N_25249,N_25451);
nor U26797 (N_26797,N_25744,N_26399);
nor U26798 (N_26798,N_26111,N_25300);
and U26799 (N_26799,N_25752,N_25712);
or U26800 (N_26800,N_25914,N_25827);
xor U26801 (N_26801,N_26298,N_25851);
xnor U26802 (N_26802,N_25438,N_26131);
or U26803 (N_26803,N_26050,N_25383);
or U26804 (N_26804,N_26375,N_26110);
xor U26805 (N_26805,N_25826,N_25502);
nor U26806 (N_26806,N_26228,N_26390);
nor U26807 (N_26807,N_26163,N_26319);
and U26808 (N_26808,N_25716,N_26093);
nor U26809 (N_26809,N_25505,N_26024);
and U26810 (N_26810,N_26158,N_26003);
and U26811 (N_26811,N_25238,N_26041);
and U26812 (N_26812,N_25321,N_26263);
xor U26813 (N_26813,N_25552,N_26383);
nand U26814 (N_26814,N_25217,N_25944);
and U26815 (N_26815,N_25863,N_25705);
xor U26816 (N_26816,N_25579,N_25644);
nor U26817 (N_26817,N_25634,N_26070);
or U26818 (N_26818,N_26205,N_26137);
and U26819 (N_26819,N_25293,N_25770);
nor U26820 (N_26820,N_26384,N_25276);
xnor U26821 (N_26821,N_25816,N_25242);
and U26822 (N_26822,N_25341,N_25676);
and U26823 (N_26823,N_26048,N_26078);
xor U26824 (N_26824,N_25651,N_25507);
nor U26825 (N_26825,N_26335,N_26294);
and U26826 (N_26826,N_25233,N_25484);
nor U26827 (N_26827,N_26072,N_25884);
nand U26828 (N_26828,N_25336,N_25381);
nand U26829 (N_26829,N_25302,N_25446);
and U26830 (N_26830,N_26364,N_26282);
nor U26831 (N_26831,N_26236,N_25958);
nor U26832 (N_26832,N_26011,N_26068);
xor U26833 (N_26833,N_25513,N_25326);
xnor U26834 (N_26834,N_26393,N_25417);
nand U26835 (N_26835,N_25468,N_25445);
xnor U26836 (N_26836,N_25364,N_25425);
nand U26837 (N_26837,N_25922,N_26002);
nor U26838 (N_26838,N_25592,N_25867);
nand U26839 (N_26839,N_25624,N_25488);
or U26840 (N_26840,N_25722,N_25214);
nand U26841 (N_26841,N_26278,N_25510);
xor U26842 (N_26842,N_26342,N_25974);
or U26843 (N_26843,N_25843,N_25616);
nand U26844 (N_26844,N_26358,N_25253);
nor U26845 (N_26845,N_26055,N_25550);
or U26846 (N_26846,N_25746,N_26098);
nor U26847 (N_26847,N_25594,N_26186);
or U26848 (N_26848,N_25354,N_26181);
or U26849 (N_26849,N_25436,N_26170);
and U26850 (N_26850,N_25564,N_25371);
and U26851 (N_26851,N_25696,N_25523);
and U26852 (N_26852,N_26166,N_26268);
nand U26853 (N_26853,N_25650,N_25875);
xnor U26854 (N_26854,N_25575,N_26015);
nor U26855 (N_26855,N_26357,N_25910);
nor U26856 (N_26856,N_26126,N_25793);
nor U26857 (N_26857,N_25946,N_25477);
and U26858 (N_26858,N_25847,N_25984);
or U26859 (N_26859,N_25660,N_25618);
nand U26860 (N_26860,N_25558,N_25862);
and U26861 (N_26861,N_25368,N_26244);
nor U26862 (N_26862,N_26207,N_26037);
xnor U26863 (N_26863,N_26088,N_25366);
nor U26864 (N_26864,N_25762,N_25516);
and U26865 (N_26865,N_25996,N_25983);
xor U26866 (N_26866,N_25671,N_25339);
nand U26867 (N_26867,N_25982,N_25979);
xor U26868 (N_26868,N_26030,N_26322);
xnor U26869 (N_26869,N_25938,N_25536);
and U26870 (N_26870,N_25232,N_26253);
or U26871 (N_26871,N_26274,N_26240);
nand U26872 (N_26872,N_25954,N_25653);
and U26873 (N_26873,N_26039,N_26129);
nor U26874 (N_26874,N_25256,N_25637);
nand U26875 (N_26875,N_25235,N_25409);
xnor U26876 (N_26876,N_26337,N_26008);
nor U26877 (N_26877,N_25251,N_26378);
nor U26878 (N_26878,N_26065,N_26229);
xor U26879 (N_26879,N_26035,N_26279);
and U26880 (N_26880,N_26109,N_25679);
or U26881 (N_26881,N_25859,N_25808);
or U26882 (N_26882,N_25223,N_26356);
nor U26883 (N_26883,N_25878,N_25603);
and U26884 (N_26884,N_26341,N_25323);
xor U26885 (N_26885,N_25967,N_25879);
nor U26886 (N_26886,N_25243,N_26147);
xor U26887 (N_26887,N_26238,N_25729);
and U26888 (N_26888,N_26058,N_25229);
nand U26889 (N_26889,N_25745,N_25285);
nand U26890 (N_26890,N_25533,N_25435);
xnor U26891 (N_26891,N_25775,N_25353);
nor U26892 (N_26892,N_25270,N_26376);
and U26893 (N_26893,N_25692,N_26235);
xor U26894 (N_26894,N_25537,N_25410);
and U26895 (N_26895,N_26297,N_25886);
nor U26896 (N_26896,N_26373,N_25263);
nor U26897 (N_26897,N_25929,N_26381);
or U26898 (N_26898,N_25781,N_25254);
xor U26899 (N_26899,N_25541,N_25736);
nand U26900 (N_26900,N_25934,N_26343);
nor U26901 (N_26901,N_25352,N_25399);
xor U26902 (N_26902,N_25718,N_25407);
and U26903 (N_26903,N_25765,N_25437);
or U26904 (N_26904,N_25880,N_26345);
and U26905 (N_26905,N_25610,N_25756);
nor U26906 (N_26906,N_25557,N_25757);
nor U26907 (N_26907,N_25959,N_25628);
nor U26908 (N_26908,N_26258,N_25395);
nor U26909 (N_26909,N_25724,N_25265);
or U26910 (N_26910,N_26128,N_26140);
nor U26911 (N_26911,N_25572,N_25951);
and U26912 (N_26912,N_26220,N_25208);
and U26913 (N_26913,N_25459,N_25821);
and U26914 (N_26914,N_25210,N_25546);
or U26915 (N_26915,N_25307,N_25281);
nand U26916 (N_26916,N_25308,N_25641);
xnor U26917 (N_26917,N_25648,N_25777);
xor U26918 (N_26918,N_26371,N_25602);
or U26919 (N_26919,N_25563,N_25766);
and U26920 (N_26920,N_26090,N_25290);
nand U26921 (N_26921,N_26317,N_25835);
nor U26922 (N_26922,N_25406,N_25200);
xor U26923 (N_26923,N_26290,N_25678);
nand U26924 (N_26924,N_25444,N_25673);
or U26925 (N_26925,N_26284,N_26077);
or U26926 (N_26926,N_25814,N_26300);
or U26927 (N_26927,N_26043,N_26188);
or U26928 (N_26928,N_25471,N_26334);
and U26929 (N_26929,N_25470,N_26164);
xor U26930 (N_26930,N_25797,N_25506);
nand U26931 (N_26931,N_25531,N_25608);
or U26932 (N_26932,N_25453,N_26145);
xnor U26933 (N_26933,N_25633,N_25294);
nand U26934 (N_26934,N_26184,N_25370);
nor U26935 (N_26935,N_25387,N_26255);
or U26936 (N_26936,N_26192,N_25693);
xnor U26937 (N_26937,N_26213,N_25926);
and U26938 (N_26938,N_25514,N_25915);
nor U26939 (N_26939,N_25971,N_25933);
and U26940 (N_26940,N_26251,N_25688);
and U26941 (N_26941,N_25548,N_25389);
or U26942 (N_26942,N_26153,N_25749);
and U26943 (N_26943,N_25871,N_26329);
or U26944 (N_26944,N_25987,N_25580);
nand U26945 (N_26945,N_25578,N_25978);
nand U26946 (N_26946,N_25727,N_25492);
nor U26947 (N_26947,N_25511,N_26155);
xor U26948 (N_26948,N_26099,N_25595);
and U26949 (N_26949,N_26144,N_25706);
or U26950 (N_26950,N_25904,N_26248);
and U26951 (N_26951,N_25819,N_25296);
xnor U26952 (N_26952,N_26347,N_25720);
nand U26953 (N_26953,N_25790,N_25940);
nor U26954 (N_26954,N_25561,N_25332);
nor U26955 (N_26955,N_25809,N_26179);
or U26956 (N_26956,N_25801,N_26332);
nand U26957 (N_26957,N_25921,N_25708);
or U26958 (N_26958,N_25320,N_25986);
nor U26959 (N_26959,N_25760,N_25824);
or U26960 (N_26960,N_25479,N_25554);
and U26961 (N_26961,N_25295,N_26208);
xor U26962 (N_26962,N_25315,N_26116);
nand U26963 (N_26963,N_26012,N_26197);
nand U26964 (N_26964,N_26245,N_25937);
and U26965 (N_26965,N_25262,N_25901);
and U26966 (N_26966,N_25674,N_25397);
nor U26967 (N_26967,N_26124,N_26292);
nor U26968 (N_26968,N_26195,N_25795);
nor U26969 (N_26969,N_25237,N_25590);
nand U26970 (N_26970,N_26252,N_25496);
or U26971 (N_26971,N_25743,N_25576);
and U26972 (N_26972,N_26148,N_25927);
nor U26973 (N_26973,N_25292,N_25452);
nor U26974 (N_26974,N_26230,N_25258);
xnor U26975 (N_26975,N_25423,N_25268);
xnor U26976 (N_26976,N_26092,N_26032);
or U26977 (N_26977,N_26014,N_26330);
and U26978 (N_26978,N_25895,N_25209);
and U26979 (N_26979,N_26176,N_25591);
and U26980 (N_26980,N_25995,N_25566);
nor U26981 (N_26981,N_25919,N_25448);
or U26982 (N_26982,N_25439,N_25385);
xnor U26983 (N_26983,N_26266,N_26151);
and U26984 (N_26984,N_26001,N_25791);
xor U26985 (N_26985,N_25657,N_25950);
nand U26986 (N_26986,N_25993,N_26397);
nand U26987 (N_26987,N_26312,N_25201);
xnor U26988 (N_26988,N_25512,N_25873);
nand U26989 (N_26989,N_26054,N_25234);
or U26990 (N_26990,N_25583,N_26175);
or U26991 (N_26991,N_26053,N_25829);
or U26992 (N_26992,N_25314,N_26075);
xor U26993 (N_26993,N_25606,N_26198);
xnor U26994 (N_26994,N_25794,N_25783);
nand U26995 (N_26995,N_26135,N_25551);
and U26996 (N_26996,N_25714,N_26301);
or U26997 (N_26997,N_25920,N_26143);
and U26998 (N_26998,N_25493,N_26080);
nand U26999 (N_26999,N_26007,N_25876);
nand U27000 (N_27000,N_25803,N_25782);
and U27001 (N_27001,N_25524,N_25818);
and U27002 (N_27002,N_25955,N_25677);
nor U27003 (N_27003,N_25322,N_25979);
and U27004 (N_27004,N_25527,N_26137);
and U27005 (N_27005,N_25969,N_25812);
or U27006 (N_27006,N_25655,N_25429);
nand U27007 (N_27007,N_25652,N_25711);
xor U27008 (N_27008,N_26085,N_25329);
and U27009 (N_27009,N_25329,N_26180);
xor U27010 (N_27010,N_26378,N_25213);
or U27011 (N_27011,N_25977,N_25335);
and U27012 (N_27012,N_26377,N_25336);
xor U27013 (N_27013,N_26229,N_25303);
and U27014 (N_27014,N_25423,N_25730);
nor U27015 (N_27015,N_25646,N_25604);
nor U27016 (N_27016,N_25632,N_25680);
nor U27017 (N_27017,N_26162,N_26314);
nand U27018 (N_27018,N_25735,N_26362);
or U27019 (N_27019,N_25613,N_25411);
nand U27020 (N_27020,N_25724,N_25755);
or U27021 (N_27021,N_25239,N_26191);
nor U27022 (N_27022,N_25853,N_25897);
or U27023 (N_27023,N_25523,N_25519);
nor U27024 (N_27024,N_26398,N_26378);
xor U27025 (N_27025,N_25948,N_26187);
and U27026 (N_27026,N_25726,N_25353);
xnor U27027 (N_27027,N_25405,N_26176);
xnor U27028 (N_27028,N_26284,N_25312);
nor U27029 (N_27029,N_25211,N_26036);
nor U27030 (N_27030,N_25903,N_26254);
nor U27031 (N_27031,N_25684,N_26343);
and U27032 (N_27032,N_25743,N_26229);
nand U27033 (N_27033,N_25818,N_25927);
nand U27034 (N_27034,N_25959,N_26309);
or U27035 (N_27035,N_26368,N_25537);
nor U27036 (N_27036,N_26335,N_25410);
nand U27037 (N_27037,N_25646,N_25251);
xor U27038 (N_27038,N_26288,N_26114);
and U27039 (N_27039,N_25592,N_25902);
and U27040 (N_27040,N_25604,N_25596);
xnor U27041 (N_27041,N_25563,N_26012);
and U27042 (N_27042,N_25942,N_25311);
and U27043 (N_27043,N_25828,N_25824);
and U27044 (N_27044,N_26265,N_25500);
xnor U27045 (N_27045,N_26043,N_25885);
nand U27046 (N_27046,N_25990,N_25392);
nand U27047 (N_27047,N_25887,N_25722);
xor U27048 (N_27048,N_25620,N_25661);
nand U27049 (N_27049,N_26273,N_25294);
nand U27050 (N_27050,N_26084,N_26306);
xnor U27051 (N_27051,N_25651,N_25405);
and U27052 (N_27052,N_25531,N_25586);
or U27053 (N_27053,N_26064,N_25802);
nor U27054 (N_27054,N_25782,N_26058);
nand U27055 (N_27055,N_25284,N_25247);
xnor U27056 (N_27056,N_25944,N_25893);
nand U27057 (N_27057,N_25307,N_25430);
nor U27058 (N_27058,N_26039,N_26335);
nand U27059 (N_27059,N_25718,N_25274);
xor U27060 (N_27060,N_25869,N_26212);
xnor U27061 (N_27061,N_25753,N_25303);
xnor U27062 (N_27062,N_25970,N_25366);
or U27063 (N_27063,N_25246,N_25582);
nor U27064 (N_27064,N_26206,N_26268);
nand U27065 (N_27065,N_25503,N_26215);
nand U27066 (N_27066,N_25833,N_25937);
nor U27067 (N_27067,N_25484,N_25538);
and U27068 (N_27068,N_25622,N_26350);
xor U27069 (N_27069,N_25507,N_26311);
nor U27070 (N_27070,N_26245,N_26164);
xor U27071 (N_27071,N_25897,N_26269);
or U27072 (N_27072,N_26174,N_26054);
or U27073 (N_27073,N_25970,N_26359);
nand U27074 (N_27074,N_25254,N_25478);
xnor U27075 (N_27075,N_25213,N_26368);
or U27076 (N_27076,N_26271,N_25988);
nor U27077 (N_27077,N_25595,N_25755);
or U27078 (N_27078,N_25987,N_25657);
and U27079 (N_27079,N_25504,N_26291);
nand U27080 (N_27080,N_25429,N_25865);
nand U27081 (N_27081,N_26306,N_25583);
or U27082 (N_27082,N_26367,N_25903);
xor U27083 (N_27083,N_25351,N_26265);
nor U27084 (N_27084,N_25832,N_25355);
nor U27085 (N_27085,N_26267,N_25662);
nand U27086 (N_27086,N_25408,N_26278);
nor U27087 (N_27087,N_25348,N_25856);
nor U27088 (N_27088,N_26003,N_25850);
nand U27089 (N_27089,N_26295,N_25546);
and U27090 (N_27090,N_25741,N_25215);
xor U27091 (N_27091,N_25661,N_26035);
xor U27092 (N_27092,N_25566,N_25821);
nand U27093 (N_27093,N_25629,N_26113);
and U27094 (N_27094,N_25807,N_26390);
and U27095 (N_27095,N_25388,N_25844);
or U27096 (N_27096,N_26118,N_26297);
nand U27097 (N_27097,N_25716,N_25768);
and U27098 (N_27098,N_26077,N_25709);
and U27099 (N_27099,N_25623,N_26341);
or U27100 (N_27100,N_25849,N_25602);
or U27101 (N_27101,N_26141,N_25930);
or U27102 (N_27102,N_25430,N_26302);
and U27103 (N_27103,N_26025,N_26039);
and U27104 (N_27104,N_25362,N_26031);
or U27105 (N_27105,N_26141,N_25960);
xor U27106 (N_27106,N_26200,N_25541);
xnor U27107 (N_27107,N_25717,N_25842);
xor U27108 (N_27108,N_25565,N_25242);
nand U27109 (N_27109,N_25592,N_25429);
nor U27110 (N_27110,N_25381,N_26320);
and U27111 (N_27111,N_25590,N_26111);
and U27112 (N_27112,N_26044,N_25794);
nand U27113 (N_27113,N_25502,N_25704);
xnor U27114 (N_27114,N_25847,N_25222);
and U27115 (N_27115,N_26111,N_25491);
xnor U27116 (N_27116,N_25653,N_25568);
and U27117 (N_27117,N_26306,N_26350);
or U27118 (N_27118,N_26225,N_25555);
xor U27119 (N_27119,N_25693,N_25896);
nand U27120 (N_27120,N_26351,N_25514);
nand U27121 (N_27121,N_25202,N_25754);
or U27122 (N_27122,N_25643,N_25918);
nor U27123 (N_27123,N_25525,N_25849);
nor U27124 (N_27124,N_25537,N_25607);
and U27125 (N_27125,N_25742,N_25549);
nor U27126 (N_27126,N_25921,N_25529);
nand U27127 (N_27127,N_25745,N_26379);
or U27128 (N_27128,N_25462,N_25941);
and U27129 (N_27129,N_26277,N_26173);
xnor U27130 (N_27130,N_25921,N_26353);
or U27131 (N_27131,N_26180,N_25782);
nand U27132 (N_27132,N_26071,N_25970);
xor U27133 (N_27133,N_25228,N_25382);
or U27134 (N_27134,N_26171,N_25281);
nand U27135 (N_27135,N_25892,N_26350);
nor U27136 (N_27136,N_25689,N_25404);
and U27137 (N_27137,N_26286,N_25490);
xnor U27138 (N_27138,N_25202,N_26049);
nand U27139 (N_27139,N_26340,N_25670);
or U27140 (N_27140,N_25874,N_26146);
xnor U27141 (N_27141,N_25766,N_25647);
or U27142 (N_27142,N_26288,N_25753);
or U27143 (N_27143,N_25206,N_26390);
xor U27144 (N_27144,N_25202,N_26191);
nor U27145 (N_27145,N_25489,N_26391);
nand U27146 (N_27146,N_26346,N_25638);
xnor U27147 (N_27147,N_26028,N_25550);
nand U27148 (N_27148,N_25606,N_25797);
or U27149 (N_27149,N_25685,N_25319);
nand U27150 (N_27150,N_25712,N_26059);
nor U27151 (N_27151,N_26355,N_26017);
or U27152 (N_27152,N_25738,N_25531);
nand U27153 (N_27153,N_25918,N_25340);
xor U27154 (N_27154,N_25424,N_25773);
nand U27155 (N_27155,N_26303,N_25652);
or U27156 (N_27156,N_25556,N_25753);
nor U27157 (N_27157,N_25939,N_25730);
nor U27158 (N_27158,N_25885,N_25815);
and U27159 (N_27159,N_25714,N_25494);
and U27160 (N_27160,N_25700,N_25575);
or U27161 (N_27161,N_26155,N_26069);
nor U27162 (N_27162,N_26312,N_26315);
nor U27163 (N_27163,N_26257,N_25807);
or U27164 (N_27164,N_25435,N_25538);
and U27165 (N_27165,N_25991,N_25453);
and U27166 (N_27166,N_25206,N_26118);
or U27167 (N_27167,N_25293,N_26180);
xnor U27168 (N_27168,N_26264,N_25671);
nor U27169 (N_27169,N_25667,N_25679);
and U27170 (N_27170,N_25654,N_25563);
xor U27171 (N_27171,N_25265,N_25467);
and U27172 (N_27172,N_25412,N_25701);
and U27173 (N_27173,N_26183,N_25379);
nand U27174 (N_27174,N_26133,N_26228);
nand U27175 (N_27175,N_25849,N_26042);
or U27176 (N_27176,N_25810,N_25755);
nand U27177 (N_27177,N_26105,N_25953);
and U27178 (N_27178,N_25585,N_25428);
nand U27179 (N_27179,N_25675,N_25566);
nor U27180 (N_27180,N_25836,N_25343);
xnor U27181 (N_27181,N_26245,N_25434);
nor U27182 (N_27182,N_26123,N_25281);
nor U27183 (N_27183,N_25713,N_26210);
nor U27184 (N_27184,N_26310,N_25675);
or U27185 (N_27185,N_25213,N_25736);
xnor U27186 (N_27186,N_26308,N_25228);
or U27187 (N_27187,N_25455,N_25354);
nor U27188 (N_27188,N_25748,N_25462);
nand U27189 (N_27189,N_26032,N_25297);
xor U27190 (N_27190,N_26255,N_25926);
and U27191 (N_27191,N_25845,N_26025);
or U27192 (N_27192,N_25689,N_26192);
and U27193 (N_27193,N_25599,N_25409);
or U27194 (N_27194,N_25598,N_25828);
xnor U27195 (N_27195,N_25988,N_26063);
nand U27196 (N_27196,N_26024,N_25488);
or U27197 (N_27197,N_25504,N_25426);
and U27198 (N_27198,N_26168,N_26083);
nand U27199 (N_27199,N_25774,N_25222);
and U27200 (N_27200,N_26076,N_25344);
nand U27201 (N_27201,N_25961,N_25396);
nand U27202 (N_27202,N_25785,N_26067);
nor U27203 (N_27203,N_25341,N_25305);
and U27204 (N_27204,N_26198,N_25480);
nor U27205 (N_27205,N_26127,N_26116);
nor U27206 (N_27206,N_25422,N_25754);
and U27207 (N_27207,N_25705,N_25992);
nor U27208 (N_27208,N_25938,N_26299);
xnor U27209 (N_27209,N_25637,N_26038);
xnor U27210 (N_27210,N_26372,N_25871);
nor U27211 (N_27211,N_25777,N_25431);
nor U27212 (N_27212,N_25646,N_26285);
nor U27213 (N_27213,N_25526,N_25407);
xnor U27214 (N_27214,N_26022,N_25932);
or U27215 (N_27215,N_25202,N_26263);
nand U27216 (N_27216,N_26052,N_25394);
nor U27217 (N_27217,N_25317,N_25307);
nand U27218 (N_27218,N_25534,N_25452);
and U27219 (N_27219,N_25933,N_25585);
or U27220 (N_27220,N_26164,N_26137);
nand U27221 (N_27221,N_25605,N_26013);
xor U27222 (N_27222,N_26030,N_26179);
nor U27223 (N_27223,N_26385,N_25802);
nand U27224 (N_27224,N_25308,N_25396);
nor U27225 (N_27225,N_26369,N_25726);
and U27226 (N_27226,N_25297,N_26384);
nand U27227 (N_27227,N_25372,N_25950);
nand U27228 (N_27228,N_26304,N_25507);
nand U27229 (N_27229,N_25608,N_26294);
xor U27230 (N_27230,N_25243,N_25787);
nand U27231 (N_27231,N_25459,N_25915);
and U27232 (N_27232,N_26022,N_26311);
nand U27233 (N_27233,N_25213,N_25303);
nor U27234 (N_27234,N_25730,N_25270);
nand U27235 (N_27235,N_26322,N_26162);
nand U27236 (N_27236,N_26361,N_26120);
or U27237 (N_27237,N_25549,N_26005);
nand U27238 (N_27238,N_25444,N_25842);
and U27239 (N_27239,N_25640,N_25293);
xor U27240 (N_27240,N_25869,N_26154);
nor U27241 (N_27241,N_26133,N_26350);
nor U27242 (N_27242,N_25948,N_25795);
and U27243 (N_27243,N_25561,N_26249);
nor U27244 (N_27244,N_26295,N_25814);
and U27245 (N_27245,N_25843,N_25550);
or U27246 (N_27246,N_26349,N_26002);
or U27247 (N_27247,N_25634,N_25441);
or U27248 (N_27248,N_26034,N_25596);
or U27249 (N_27249,N_25207,N_25895);
xor U27250 (N_27250,N_26058,N_25725);
nor U27251 (N_27251,N_25897,N_25746);
or U27252 (N_27252,N_25962,N_25294);
and U27253 (N_27253,N_25239,N_25350);
or U27254 (N_27254,N_25200,N_26211);
or U27255 (N_27255,N_25513,N_25845);
and U27256 (N_27256,N_26289,N_26310);
nor U27257 (N_27257,N_25878,N_26368);
nor U27258 (N_27258,N_25803,N_25348);
and U27259 (N_27259,N_25612,N_26346);
and U27260 (N_27260,N_25971,N_25258);
nand U27261 (N_27261,N_26205,N_25803);
and U27262 (N_27262,N_26292,N_25731);
or U27263 (N_27263,N_25378,N_26338);
or U27264 (N_27264,N_25472,N_26120);
and U27265 (N_27265,N_25214,N_26154);
nor U27266 (N_27266,N_26148,N_25585);
nand U27267 (N_27267,N_25506,N_26081);
or U27268 (N_27268,N_25292,N_25346);
and U27269 (N_27269,N_25746,N_25531);
nand U27270 (N_27270,N_25732,N_25270);
and U27271 (N_27271,N_25666,N_25284);
xnor U27272 (N_27272,N_25868,N_26209);
xor U27273 (N_27273,N_26278,N_25523);
xor U27274 (N_27274,N_25241,N_26069);
xnor U27275 (N_27275,N_25879,N_25530);
xnor U27276 (N_27276,N_25331,N_25392);
or U27277 (N_27277,N_25291,N_25262);
or U27278 (N_27278,N_26242,N_26209);
nor U27279 (N_27279,N_26171,N_26209);
xnor U27280 (N_27280,N_25632,N_26181);
nor U27281 (N_27281,N_26217,N_26185);
nand U27282 (N_27282,N_25583,N_25500);
or U27283 (N_27283,N_26159,N_25339);
nor U27284 (N_27284,N_25447,N_26226);
nand U27285 (N_27285,N_25295,N_25526);
xnor U27286 (N_27286,N_26066,N_25674);
nand U27287 (N_27287,N_26297,N_26253);
and U27288 (N_27288,N_26384,N_26269);
xnor U27289 (N_27289,N_25832,N_25632);
nand U27290 (N_27290,N_25427,N_26085);
nor U27291 (N_27291,N_26378,N_26001);
nand U27292 (N_27292,N_25982,N_25508);
nand U27293 (N_27293,N_26224,N_25326);
nand U27294 (N_27294,N_25340,N_25590);
nor U27295 (N_27295,N_26348,N_26390);
xor U27296 (N_27296,N_25467,N_25961);
nor U27297 (N_27297,N_26251,N_26194);
nor U27298 (N_27298,N_25482,N_25845);
nor U27299 (N_27299,N_25569,N_25922);
nor U27300 (N_27300,N_25672,N_25761);
xor U27301 (N_27301,N_26359,N_26074);
nand U27302 (N_27302,N_25962,N_25795);
nor U27303 (N_27303,N_26097,N_25864);
or U27304 (N_27304,N_25300,N_25239);
nor U27305 (N_27305,N_25452,N_25952);
xnor U27306 (N_27306,N_25371,N_26311);
and U27307 (N_27307,N_26297,N_25857);
xor U27308 (N_27308,N_25499,N_26317);
and U27309 (N_27309,N_25615,N_25975);
and U27310 (N_27310,N_25201,N_25766);
and U27311 (N_27311,N_25765,N_26100);
nor U27312 (N_27312,N_26363,N_25964);
nor U27313 (N_27313,N_26260,N_25742);
nor U27314 (N_27314,N_25692,N_25251);
and U27315 (N_27315,N_26367,N_25901);
nor U27316 (N_27316,N_25615,N_26189);
or U27317 (N_27317,N_26330,N_25280);
or U27318 (N_27318,N_25603,N_26379);
xnor U27319 (N_27319,N_26109,N_26301);
or U27320 (N_27320,N_25762,N_25538);
and U27321 (N_27321,N_26183,N_25990);
or U27322 (N_27322,N_25992,N_26141);
nor U27323 (N_27323,N_25272,N_25717);
nand U27324 (N_27324,N_25268,N_26272);
nor U27325 (N_27325,N_25978,N_25596);
xnor U27326 (N_27326,N_26153,N_26385);
or U27327 (N_27327,N_25627,N_25606);
nor U27328 (N_27328,N_25368,N_25755);
and U27329 (N_27329,N_26352,N_26060);
xnor U27330 (N_27330,N_26107,N_25824);
xor U27331 (N_27331,N_25785,N_25263);
xor U27332 (N_27332,N_26129,N_26124);
nand U27333 (N_27333,N_26307,N_26320);
or U27334 (N_27334,N_26093,N_25343);
and U27335 (N_27335,N_26344,N_26383);
or U27336 (N_27336,N_25386,N_26285);
nand U27337 (N_27337,N_25214,N_25824);
nor U27338 (N_27338,N_26092,N_25899);
nand U27339 (N_27339,N_25519,N_25273);
and U27340 (N_27340,N_25344,N_25348);
and U27341 (N_27341,N_25281,N_25652);
xor U27342 (N_27342,N_25293,N_25290);
or U27343 (N_27343,N_26134,N_26028);
nand U27344 (N_27344,N_26288,N_25347);
nor U27345 (N_27345,N_25551,N_26005);
or U27346 (N_27346,N_25699,N_26094);
or U27347 (N_27347,N_25232,N_26218);
and U27348 (N_27348,N_25635,N_25374);
xor U27349 (N_27349,N_26318,N_26192);
and U27350 (N_27350,N_25352,N_25479);
xnor U27351 (N_27351,N_25391,N_25404);
nor U27352 (N_27352,N_25816,N_26333);
xor U27353 (N_27353,N_25730,N_25844);
nand U27354 (N_27354,N_25396,N_26254);
nor U27355 (N_27355,N_25981,N_25507);
nand U27356 (N_27356,N_26345,N_25597);
nor U27357 (N_27357,N_25765,N_25383);
nor U27358 (N_27358,N_25307,N_25490);
or U27359 (N_27359,N_25664,N_25708);
nand U27360 (N_27360,N_25942,N_25884);
and U27361 (N_27361,N_25942,N_26268);
xor U27362 (N_27362,N_26023,N_26314);
nor U27363 (N_27363,N_26111,N_25921);
and U27364 (N_27364,N_25755,N_25444);
xnor U27365 (N_27365,N_25264,N_25782);
nor U27366 (N_27366,N_25384,N_26163);
nor U27367 (N_27367,N_25465,N_25956);
or U27368 (N_27368,N_25265,N_26246);
or U27369 (N_27369,N_26315,N_25771);
or U27370 (N_27370,N_25210,N_25392);
nand U27371 (N_27371,N_26159,N_26284);
or U27372 (N_27372,N_25948,N_25436);
or U27373 (N_27373,N_26037,N_25710);
or U27374 (N_27374,N_26318,N_25649);
nand U27375 (N_27375,N_25478,N_26070);
and U27376 (N_27376,N_25380,N_26081);
nand U27377 (N_27377,N_25224,N_25809);
and U27378 (N_27378,N_25787,N_26022);
xnor U27379 (N_27379,N_25494,N_25349);
nor U27380 (N_27380,N_25567,N_25860);
nor U27381 (N_27381,N_25295,N_25824);
and U27382 (N_27382,N_25926,N_25459);
xnor U27383 (N_27383,N_25525,N_25393);
and U27384 (N_27384,N_25887,N_25714);
nor U27385 (N_27385,N_25960,N_26365);
or U27386 (N_27386,N_25651,N_26297);
and U27387 (N_27387,N_25533,N_26066);
and U27388 (N_27388,N_26237,N_26205);
and U27389 (N_27389,N_25844,N_25885);
xnor U27390 (N_27390,N_26386,N_26332);
and U27391 (N_27391,N_25621,N_26376);
nor U27392 (N_27392,N_26384,N_25779);
nand U27393 (N_27393,N_25735,N_26374);
or U27394 (N_27394,N_25415,N_25725);
nor U27395 (N_27395,N_26356,N_25793);
or U27396 (N_27396,N_26048,N_25595);
nor U27397 (N_27397,N_26284,N_25387);
and U27398 (N_27398,N_26190,N_25720);
nand U27399 (N_27399,N_25442,N_25210);
xnor U27400 (N_27400,N_26282,N_26291);
nand U27401 (N_27401,N_25659,N_25982);
nor U27402 (N_27402,N_25951,N_26131);
nand U27403 (N_27403,N_26134,N_25929);
xor U27404 (N_27404,N_26015,N_25396);
or U27405 (N_27405,N_25388,N_25454);
xor U27406 (N_27406,N_26256,N_25549);
or U27407 (N_27407,N_25712,N_25873);
xor U27408 (N_27408,N_26232,N_26008);
nand U27409 (N_27409,N_25575,N_25369);
nor U27410 (N_27410,N_26308,N_25350);
nor U27411 (N_27411,N_25480,N_25799);
and U27412 (N_27412,N_26287,N_25211);
xor U27413 (N_27413,N_26289,N_25672);
and U27414 (N_27414,N_26000,N_25787);
or U27415 (N_27415,N_25311,N_25607);
or U27416 (N_27416,N_25998,N_26130);
nor U27417 (N_27417,N_25887,N_25222);
xnor U27418 (N_27418,N_25536,N_25220);
xnor U27419 (N_27419,N_26207,N_26392);
or U27420 (N_27420,N_25952,N_25270);
xnor U27421 (N_27421,N_25221,N_25579);
xor U27422 (N_27422,N_25271,N_26000);
xor U27423 (N_27423,N_26290,N_25713);
or U27424 (N_27424,N_26258,N_25988);
and U27425 (N_27425,N_25216,N_25793);
nor U27426 (N_27426,N_25331,N_26275);
and U27427 (N_27427,N_25914,N_25486);
or U27428 (N_27428,N_25925,N_25330);
xnor U27429 (N_27429,N_26323,N_25492);
and U27430 (N_27430,N_26236,N_25438);
xnor U27431 (N_27431,N_26150,N_25360);
nand U27432 (N_27432,N_25288,N_25215);
nor U27433 (N_27433,N_25251,N_25321);
and U27434 (N_27434,N_25659,N_26080);
nand U27435 (N_27435,N_25219,N_26179);
or U27436 (N_27436,N_26038,N_25474);
and U27437 (N_27437,N_25779,N_25433);
or U27438 (N_27438,N_26178,N_25289);
nand U27439 (N_27439,N_26299,N_25827);
xnor U27440 (N_27440,N_26173,N_26349);
xnor U27441 (N_27441,N_25499,N_25843);
nand U27442 (N_27442,N_26228,N_26206);
nor U27443 (N_27443,N_26285,N_25886);
nor U27444 (N_27444,N_25642,N_26343);
or U27445 (N_27445,N_25957,N_26137);
xor U27446 (N_27446,N_25712,N_25410);
and U27447 (N_27447,N_25717,N_25260);
xnor U27448 (N_27448,N_25324,N_26363);
nand U27449 (N_27449,N_25616,N_25387);
nand U27450 (N_27450,N_25737,N_25612);
or U27451 (N_27451,N_26034,N_25662);
and U27452 (N_27452,N_26006,N_25440);
xnor U27453 (N_27453,N_25899,N_25600);
nor U27454 (N_27454,N_25959,N_26195);
and U27455 (N_27455,N_25982,N_25516);
nor U27456 (N_27456,N_25540,N_25367);
nor U27457 (N_27457,N_26367,N_25593);
xnor U27458 (N_27458,N_25642,N_25514);
nand U27459 (N_27459,N_25392,N_25887);
or U27460 (N_27460,N_25784,N_26335);
or U27461 (N_27461,N_25485,N_25981);
xnor U27462 (N_27462,N_25686,N_25549);
nand U27463 (N_27463,N_26344,N_25892);
nand U27464 (N_27464,N_25299,N_25470);
or U27465 (N_27465,N_25278,N_25270);
xnor U27466 (N_27466,N_25449,N_25844);
or U27467 (N_27467,N_25834,N_25703);
and U27468 (N_27468,N_25390,N_25603);
and U27469 (N_27469,N_26254,N_25274);
and U27470 (N_27470,N_25482,N_26210);
or U27471 (N_27471,N_25972,N_25868);
or U27472 (N_27472,N_26375,N_25762);
nand U27473 (N_27473,N_25548,N_25888);
nand U27474 (N_27474,N_25833,N_25255);
or U27475 (N_27475,N_25819,N_25788);
or U27476 (N_27476,N_25740,N_25973);
nand U27477 (N_27477,N_26064,N_25457);
nand U27478 (N_27478,N_25990,N_26126);
nand U27479 (N_27479,N_26342,N_25909);
xnor U27480 (N_27480,N_26122,N_25538);
and U27481 (N_27481,N_26190,N_26306);
or U27482 (N_27482,N_26216,N_25290);
nand U27483 (N_27483,N_25506,N_26088);
nand U27484 (N_27484,N_25845,N_25447);
or U27485 (N_27485,N_25562,N_25915);
nor U27486 (N_27486,N_25438,N_26295);
and U27487 (N_27487,N_26303,N_25727);
xor U27488 (N_27488,N_25335,N_25737);
nand U27489 (N_27489,N_26278,N_26288);
xnor U27490 (N_27490,N_25467,N_26083);
nand U27491 (N_27491,N_25718,N_25637);
nand U27492 (N_27492,N_26333,N_25787);
or U27493 (N_27493,N_26314,N_25508);
xor U27494 (N_27494,N_25384,N_26184);
nand U27495 (N_27495,N_25697,N_26395);
nand U27496 (N_27496,N_25865,N_26031);
or U27497 (N_27497,N_26049,N_26035);
nor U27498 (N_27498,N_25990,N_25488);
nand U27499 (N_27499,N_26038,N_25857);
nand U27500 (N_27500,N_25531,N_25843);
or U27501 (N_27501,N_26312,N_26135);
nand U27502 (N_27502,N_25891,N_26095);
xor U27503 (N_27503,N_25585,N_25985);
and U27504 (N_27504,N_25856,N_25726);
or U27505 (N_27505,N_25364,N_25384);
nand U27506 (N_27506,N_26198,N_25549);
or U27507 (N_27507,N_25237,N_26178);
xor U27508 (N_27508,N_26368,N_25624);
nand U27509 (N_27509,N_25694,N_25330);
or U27510 (N_27510,N_26266,N_25290);
xnor U27511 (N_27511,N_25508,N_25574);
and U27512 (N_27512,N_25842,N_25228);
and U27513 (N_27513,N_25604,N_25528);
xor U27514 (N_27514,N_26054,N_26073);
nor U27515 (N_27515,N_25968,N_26159);
nor U27516 (N_27516,N_25301,N_26333);
nor U27517 (N_27517,N_26010,N_26270);
nand U27518 (N_27518,N_26225,N_25678);
xnor U27519 (N_27519,N_25395,N_25411);
xnor U27520 (N_27520,N_25318,N_25557);
nor U27521 (N_27521,N_25553,N_25695);
nand U27522 (N_27522,N_25263,N_25467);
xor U27523 (N_27523,N_25785,N_26174);
and U27524 (N_27524,N_25586,N_26075);
or U27525 (N_27525,N_26279,N_25240);
and U27526 (N_27526,N_26325,N_26301);
or U27527 (N_27527,N_26035,N_25734);
xnor U27528 (N_27528,N_25933,N_25893);
nand U27529 (N_27529,N_25602,N_25554);
nand U27530 (N_27530,N_26129,N_25601);
or U27531 (N_27531,N_26210,N_26369);
xnor U27532 (N_27532,N_25327,N_25707);
and U27533 (N_27533,N_26373,N_25824);
xnor U27534 (N_27534,N_25467,N_26387);
nor U27535 (N_27535,N_25644,N_26225);
nand U27536 (N_27536,N_25885,N_26233);
or U27537 (N_27537,N_26342,N_25856);
and U27538 (N_27538,N_25420,N_25267);
nor U27539 (N_27539,N_25468,N_25991);
xnor U27540 (N_27540,N_25224,N_25620);
xor U27541 (N_27541,N_25592,N_25664);
and U27542 (N_27542,N_25961,N_26153);
nand U27543 (N_27543,N_25540,N_25229);
or U27544 (N_27544,N_25516,N_25423);
and U27545 (N_27545,N_26086,N_26281);
xor U27546 (N_27546,N_25208,N_25318);
or U27547 (N_27547,N_25500,N_25494);
nand U27548 (N_27548,N_25519,N_26184);
nor U27549 (N_27549,N_25888,N_25808);
xor U27550 (N_27550,N_25522,N_25407);
xor U27551 (N_27551,N_26003,N_25974);
nor U27552 (N_27552,N_25993,N_25919);
or U27553 (N_27553,N_25914,N_25423);
nand U27554 (N_27554,N_26115,N_25786);
and U27555 (N_27555,N_26225,N_26044);
xor U27556 (N_27556,N_25300,N_25812);
xor U27557 (N_27557,N_25779,N_26330);
or U27558 (N_27558,N_25279,N_25243);
or U27559 (N_27559,N_25639,N_25625);
and U27560 (N_27560,N_25629,N_25656);
xnor U27561 (N_27561,N_25343,N_26085);
and U27562 (N_27562,N_25652,N_25372);
or U27563 (N_27563,N_25451,N_26063);
nand U27564 (N_27564,N_25289,N_25290);
nand U27565 (N_27565,N_25272,N_25932);
nand U27566 (N_27566,N_25451,N_25623);
xor U27567 (N_27567,N_26387,N_26290);
xor U27568 (N_27568,N_25812,N_26152);
and U27569 (N_27569,N_25459,N_25902);
xor U27570 (N_27570,N_26103,N_25604);
or U27571 (N_27571,N_25215,N_25871);
and U27572 (N_27572,N_25901,N_25845);
or U27573 (N_27573,N_25830,N_26213);
xnor U27574 (N_27574,N_25732,N_26153);
xnor U27575 (N_27575,N_26093,N_26167);
or U27576 (N_27576,N_25244,N_26050);
xor U27577 (N_27577,N_25847,N_25211);
nand U27578 (N_27578,N_25525,N_25385);
and U27579 (N_27579,N_25388,N_25367);
xor U27580 (N_27580,N_25993,N_25764);
xor U27581 (N_27581,N_25767,N_25788);
nor U27582 (N_27582,N_25922,N_26274);
or U27583 (N_27583,N_26338,N_25422);
nor U27584 (N_27584,N_25323,N_25511);
xor U27585 (N_27585,N_26151,N_25433);
and U27586 (N_27586,N_25776,N_25566);
or U27587 (N_27587,N_25673,N_26160);
or U27588 (N_27588,N_25446,N_25423);
nand U27589 (N_27589,N_26399,N_25557);
nand U27590 (N_27590,N_26059,N_25490);
nand U27591 (N_27591,N_25376,N_26243);
nor U27592 (N_27592,N_25916,N_25586);
xor U27593 (N_27593,N_25496,N_25301);
xnor U27594 (N_27594,N_26002,N_25237);
or U27595 (N_27595,N_25401,N_26183);
and U27596 (N_27596,N_25811,N_25676);
or U27597 (N_27597,N_25625,N_25901);
nand U27598 (N_27598,N_26201,N_25863);
and U27599 (N_27599,N_25460,N_26292);
nor U27600 (N_27600,N_27375,N_26772);
nand U27601 (N_27601,N_27146,N_27154);
and U27602 (N_27602,N_27156,N_26683);
nor U27603 (N_27603,N_27041,N_27524);
nand U27604 (N_27604,N_27172,N_26703);
nor U27605 (N_27605,N_27000,N_26681);
or U27606 (N_27606,N_26668,N_27461);
or U27607 (N_27607,N_26822,N_27169);
xor U27608 (N_27608,N_26891,N_27356);
nand U27609 (N_27609,N_27022,N_26675);
nor U27610 (N_27610,N_27152,N_26485);
nor U27611 (N_27611,N_27181,N_26856);
xnor U27612 (N_27612,N_26526,N_26748);
or U27613 (N_27613,N_26679,N_26446);
or U27614 (N_27614,N_27373,N_27199);
nand U27615 (N_27615,N_26985,N_26933);
or U27616 (N_27616,N_26569,N_27405);
nor U27617 (N_27617,N_26945,N_27572);
xor U27618 (N_27618,N_26466,N_27585);
and U27619 (N_27619,N_26862,N_27299);
xnor U27620 (N_27620,N_27473,N_26570);
or U27621 (N_27621,N_26966,N_26801);
nand U27622 (N_27622,N_26875,N_26723);
nor U27623 (N_27623,N_26749,N_27072);
xor U27624 (N_27624,N_26475,N_27224);
and U27625 (N_27625,N_26881,N_26908);
nand U27626 (N_27626,N_26480,N_27414);
xnor U27627 (N_27627,N_26976,N_26951);
nor U27628 (N_27628,N_27031,N_27326);
or U27629 (N_27629,N_27013,N_26869);
nand U27630 (N_27630,N_27471,N_26661);
xnor U27631 (N_27631,N_26560,N_26437);
nor U27632 (N_27632,N_26702,N_26435);
or U27633 (N_27633,N_26664,N_27558);
xnor U27634 (N_27634,N_27376,N_27204);
nand U27635 (N_27635,N_27451,N_27313);
or U27636 (N_27636,N_26708,N_27305);
nor U27637 (N_27637,N_26781,N_27162);
and U27638 (N_27638,N_26717,N_26500);
nor U27639 (N_27639,N_26863,N_27590);
or U27640 (N_27640,N_27278,N_27424);
nand U27641 (N_27641,N_27077,N_26799);
xor U27642 (N_27642,N_27186,N_26828);
nand U27643 (N_27643,N_26740,N_26665);
or U27644 (N_27644,N_27068,N_27467);
or U27645 (N_27645,N_26496,N_26741);
xor U27646 (N_27646,N_27233,N_27063);
xor U27647 (N_27647,N_26796,N_26906);
and U27648 (N_27648,N_27534,N_27272);
xor U27649 (N_27649,N_26402,N_26980);
and U27650 (N_27650,N_27381,N_26459);
nor U27651 (N_27651,N_26688,N_26759);
nand U27652 (N_27652,N_27258,N_26979);
nor U27653 (N_27653,N_27098,N_27443);
xor U27654 (N_27654,N_26921,N_27331);
or U27655 (N_27655,N_27480,N_26880);
and U27656 (N_27656,N_26499,N_26685);
or U27657 (N_27657,N_26425,N_27141);
xor U27658 (N_27658,N_26785,N_27274);
nor U27659 (N_27659,N_26438,N_26696);
nor U27660 (N_27660,N_27266,N_27478);
and U27661 (N_27661,N_26483,N_27001);
or U27662 (N_27662,N_26449,N_26479);
xor U27663 (N_27663,N_27412,N_27328);
xor U27664 (N_27664,N_27486,N_26607);
nand U27665 (N_27665,N_27066,N_27521);
xor U27666 (N_27666,N_27588,N_27545);
and U27667 (N_27667,N_26554,N_26501);
nand U27668 (N_27668,N_26883,N_27007);
nand U27669 (N_27669,N_26729,N_26902);
nor U27670 (N_27670,N_27229,N_27538);
and U27671 (N_27671,N_27416,N_27002);
nor U27672 (N_27672,N_27102,N_26533);
nand U27673 (N_27673,N_27354,N_26733);
and U27674 (N_27674,N_26415,N_26847);
nor U27675 (N_27675,N_27500,N_27113);
or U27676 (N_27676,N_27234,N_26783);
nor U27677 (N_27677,N_27308,N_26580);
or U27678 (N_27678,N_27401,N_27025);
xor U27679 (N_27679,N_27061,N_27554);
and U27680 (N_27680,N_26901,N_26495);
and U27681 (N_27681,N_26414,N_26837);
nand U27682 (N_27682,N_26518,N_27158);
nor U27683 (N_27683,N_26430,N_27338);
nor U27684 (N_27684,N_26897,N_26470);
or U27685 (N_27685,N_26697,N_27073);
nor U27686 (N_27686,N_26874,N_26990);
nor U27687 (N_27687,N_26886,N_26768);
xor U27688 (N_27688,N_27231,N_27460);
xnor U27689 (N_27689,N_27133,N_26407);
nand U27690 (N_27690,N_26877,N_27127);
xor U27691 (N_27691,N_27097,N_26761);
and U27692 (N_27692,N_27295,N_26916);
nand U27693 (N_27693,N_26509,N_27253);
or U27694 (N_27694,N_26581,N_26728);
or U27695 (N_27695,N_27265,N_26556);
nand U27696 (N_27696,N_27254,N_26885);
and U27697 (N_27697,N_26907,N_26807);
or U27698 (N_27698,N_27410,N_26421);
xnor U27699 (N_27699,N_27245,N_27288);
xnor U27700 (N_27700,N_27351,N_27557);
nand U27701 (N_27701,N_27419,N_27241);
nor U27702 (N_27702,N_26974,N_27028);
nor U27703 (N_27703,N_26704,N_26598);
or U27704 (N_27704,N_26644,N_27393);
or U27705 (N_27705,N_27014,N_27309);
nand U27706 (N_27706,N_26462,N_26623);
and U27707 (N_27707,N_26525,N_27446);
nand U27708 (N_27708,N_27251,N_27088);
or U27709 (N_27709,N_26550,N_27128);
and U27710 (N_27710,N_27193,N_26636);
xor U27711 (N_27711,N_27380,N_27277);
xnor U27712 (N_27712,N_27280,N_27391);
nor U27713 (N_27713,N_27173,N_26818);
xnor U27714 (N_27714,N_26516,N_27399);
and U27715 (N_27715,N_27357,N_26695);
nand U27716 (N_27716,N_27397,N_26724);
nand U27717 (N_27717,N_27287,N_26784);
nand U27718 (N_27718,N_26409,N_27155);
and U27719 (N_27719,N_27114,N_26476);
nor U27720 (N_27720,N_27327,N_26978);
and U27721 (N_27721,N_27171,N_27188);
or U27722 (N_27722,N_27503,N_26586);
and U27723 (N_27723,N_27055,N_26443);
or U27724 (N_27724,N_27544,N_27440);
and U27725 (N_27725,N_27372,N_26953);
nor U27726 (N_27726,N_26868,N_27131);
nand U27727 (N_27727,N_27122,N_26492);
nand U27728 (N_27728,N_27067,N_26743);
xnor U27729 (N_27729,N_26531,N_26417);
nor U27730 (N_27730,N_27513,N_26848);
nand U27731 (N_27731,N_26436,N_27275);
nor U27732 (N_27732,N_27353,N_26538);
nand U27733 (N_27733,N_26789,N_26987);
or U27734 (N_27734,N_27337,N_27165);
nor U27735 (N_27735,N_26558,N_27575);
nor U27736 (N_27736,N_27542,N_27011);
xor U27737 (N_27737,N_27520,N_26963);
nand U27738 (N_27738,N_27487,N_27095);
or U27739 (N_27739,N_27382,N_26737);
and U27740 (N_27740,N_26660,N_26502);
nor U27741 (N_27741,N_26893,N_26400);
nor U27742 (N_27742,N_27048,N_26972);
or U27743 (N_27743,N_27358,N_26653);
nand U27744 (N_27744,N_27569,N_26730);
nor U27745 (N_27745,N_27045,N_26962);
nor U27746 (N_27746,N_27053,N_27285);
nand U27747 (N_27747,N_27056,N_27361);
nor U27748 (N_27748,N_26454,N_26684);
and U27749 (N_27749,N_27227,N_27168);
xor U27750 (N_27750,N_26746,N_27383);
and U27751 (N_27751,N_26544,N_27510);
nor U27752 (N_27752,N_26530,N_26814);
nand U27753 (N_27753,N_27016,N_26849);
nand U27754 (N_27754,N_26488,N_27195);
and U27755 (N_27755,N_26678,N_26843);
nand U27756 (N_27756,N_27250,N_27344);
or U27757 (N_27757,N_26770,N_26461);
nand U27758 (N_27758,N_27599,N_27054);
xor U27759 (N_27759,N_27093,N_27321);
nand U27760 (N_27760,N_27591,N_27075);
xor U27761 (N_27761,N_27504,N_26521);
and U27762 (N_27762,N_27592,N_26934);
nor U27763 (N_27763,N_26810,N_27336);
or U27764 (N_27764,N_27252,N_27150);
or U27765 (N_27765,N_27444,N_27530);
nand U27766 (N_27766,N_26497,N_27580);
or U27767 (N_27767,N_27064,N_26540);
xnor U27768 (N_27768,N_27247,N_26899);
and U27769 (N_27769,N_26692,N_26715);
and U27770 (N_27770,N_27525,N_26403);
nor U27771 (N_27771,N_27598,N_26769);
or U27772 (N_27772,N_27333,N_26835);
xnor U27773 (N_27773,N_27347,N_26790);
and U27774 (N_27774,N_27106,N_26523);
nor U27775 (N_27775,N_26505,N_26656);
and U27776 (N_27776,N_26764,N_26611);
xor U27777 (N_27777,N_26830,N_27573);
nand U27778 (N_27778,N_27187,N_27197);
or U27779 (N_27779,N_27293,N_26813);
xor U27780 (N_27780,N_27581,N_27453);
xnor U27781 (N_27781,N_26924,N_27047);
nand U27782 (N_27782,N_26944,N_27540);
xor U27783 (N_27783,N_27220,N_26453);
and U27784 (N_27784,N_27078,N_26508);
nand U27785 (N_27785,N_26662,N_27240);
or U27786 (N_27786,N_26424,N_27322);
nor U27787 (N_27787,N_26426,N_27135);
nand U27788 (N_27788,N_27519,N_27470);
and U27789 (N_27789,N_27059,N_26510);
and U27790 (N_27790,N_27472,N_27089);
and U27791 (N_27791,N_26853,N_27069);
or U27792 (N_27792,N_27300,N_26745);
or U27793 (N_27793,N_27085,N_27107);
and U27794 (N_27794,N_26973,N_27341);
nor U27795 (N_27795,N_26725,N_27298);
xor U27796 (N_27796,N_27566,N_26522);
xnor U27797 (N_27797,N_27317,N_27130);
nor U27798 (N_27798,N_27226,N_26777);
and U27799 (N_27799,N_26797,N_27213);
or U27800 (N_27800,N_27597,N_27284);
nor U27801 (N_27801,N_26969,N_27535);
nor U27802 (N_27802,N_27511,N_27352);
nor U27803 (N_27803,N_27369,N_26706);
and U27804 (N_27804,N_27483,N_26616);
or U27805 (N_27805,N_27475,N_27311);
xnor U27806 (N_27806,N_26992,N_27484);
nand U27807 (N_27807,N_26536,N_26800);
and U27808 (N_27808,N_27105,N_27457);
xor U27809 (N_27809,N_26646,N_26631);
and U27810 (N_27810,N_26619,N_26782);
nand U27811 (N_27811,N_26961,N_27035);
nand U27812 (N_27812,N_27196,N_27547);
nand U27813 (N_27813,N_26610,N_27541);
or U27814 (N_27814,N_26858,N_26941);
or U27815 (N_27815,N_26836,N_26870);
nand U27816 (N_27816,N_26567,N_26788);
xnor U27817 (N_27817,N_26983,N_27297);
nand U27818 (N_27818,N_27218,N_27394);
nand U27819 (N_27819,N_27008,N_26892);
xnor U27820 (N_27820,N_27190,N_26829);
and U27821 (N_27821,N_26658,N_27390);
xnor U27822 (N_27822,N_27413,N_27215);
nand U27823 (N_27823,N_27009,N_27281);
xor U27824 (N_27824,N_26698,N_26939);
and U27825 (N_27825,N_27118,N_26520);
nand U27826 (N_27826,N_26641,N_26467);
and U27827 (N_27827,N_27126,N_26986);
xor U27828 (N_27828,N_27374,N_26712);
nand U27829 (N_27829,N_27384,N_26956);
xnor U27830 (N_27830,N_27593,N_27420);
nand U27831 (N_27831,N_27447,N_27342);
xor U27832 (N_27832,N_27065,N_27210);
or U27833 (N_27833,N_27364,N_27415);
nand U27834 (N_27834,N_26442,N_27579);
and U27835 (N_27835,N_26844,N_26589);
or U27836 (N_27836,N_26559,N_27345);
xor U27837 (N_27837,N_27499,N_26626);
nand U27838 (N_27838,N_27032,N_26691);
nand U27839 (N_27839,N_26404,N_27217);
nor U27840 (N_27840,N_26989,N_26721);
and U27841 (N_27841,N_27296,N_27307);
nor U27842 (N_27842,N_26596,N_26517);
nand U27843 (N_27843,N_27332,N_26632);
xnor U27844 (N_27844,N_27208,N_26791);
nor U27845 (N_27845,N_26718,N_27026);
nand U27846 (N_27846,N_27255,N_27316);
xnor U27847 (N_27847,N_26484,N_26529);
nor U27848 (N_27848,N_27211,N_27292);
nor U27849 (N_27849,N_27030,N_27235);
or U27850 (N_27850,N_27586,N_26971);
or U27851 (N_27851,N_27466,N_26776);
and U27852 (N_27852,N_26542,N_27441);
or U27853 (N_27853,N_27019,N_26456);
nor U27854 (N_27854,N_27360,N_27005);
nor U27855 (N_27855,N_27112,N_26753);
nand U27856 (N_27856,N_27362,N_26628);
nor U27857 (N_27857,N_26463,N_26482);
nand U27858 (N_27858,N_26627,N_27438);
xnor U27859 (N_27859,N_27294,N_27594);
xor U27860 (N_27860,N_27058,N_26655);
and U27861 (N_27861,N_26838,N_27403);
nand U27862 (N_27862,N_27423,N_27046);
xor U27863 (N_27863,N_26851,N_26657);
nor U27864 (N_27864,N_26601,N_27176);
xor U27865 (N_27865,N_26468,N_27505);
and U27866 (N_27866,N_26690,N_27550);
and U27867 (N_27867,N_27012,N_26689);
nor U27868 (N_27868,N_26931,N_26669);
nand U27869 (N_27869,N_27109,N_27003);
nand U27870 (N_27870,N_27445,N_26620);
and U27871 (N_27871,N_27422,N_26666);
xnor U27872 (N_27872,N_26895,N_26555);
nand U27873 (N_27873,N_26894,N_27236);
nand U27874 (N_27874,N_27271,N_27389);
xnor U27875 (N_27875,N_26896,N_27312);
or U27876 (N_27876,N_27431,N_26574);
nand U27877 (N_27877,N_27346,N_26605);
xor U27878 (N_27878,N_27163,N_26551);
or U27879 (N_27879,N_27518,N_27355);
nand U27880 (N_27880,N_26471,N_26600);
xnor U27881 (N_27881,N_26564,N_27371);
or U27882 (N_27882,N_26590,N_27330);
xnor U27883 (N_27883,N_27279,N_26845);
xor U27884 (N_27884,N_27303,N_26634);
nor U27885 (N_27885,N_26816,N_27212);
nand U27886 (N_27886,N_26942,N_27076);
and U27887 (N_27887,N_27033,N_26489);
or U27888 (N_27888,N_27110,N_27157);
xor U27889 (N_27889,N_27549,N_27177);
nor U27890 (N_27890,N_26585,N_26553);
and U27891 (N_27891,N_26850,N_26964);
nand U27892 (N_27892,N_27090,N_27216);
nor U27893 (N_27893,N_27206,N_26566);
and U27894 (N_27894,N_27553,N_27276);
xnor U27895 (N_27895,N_27194,N_27493);
nor U27896 (N_27896,N_26420,N_27474);
nand U27897 (N_27897,N_27455,N_26959);
nor U27898 (N_27898,N_27514,N_26648);
xnor U27899 (N_27899,N_27185,N_26824);
nor U27900 (N_27900,N_26827,N_26519);
or U27901 (N_27901,N_26617,N_26419);
xor U27902 (N_27902,N_27315,N_26938);
nand U27903 (N_27903,N_27571,N_26444);
xor U27904 (N_27904,N_27024,N_27010);
xor U27905 (N_27905,N_27042,N_27082);
xor U27906 (N_27906,N_27363,N_26763);
xor U27907 (N_27907,N_26852,N_27370);
or U27908 (N_27908,N_27555,N_27546);
xor U27909 (N_27909,N_26481,N_27497);
nor U27910 (N_27910,N_26831,N_27552);
nand U27911 (N_27911,N_26701,N_26903);
and U27912 (N_27912,N_27201,N_26418);
and U27913 (N_27913,N_26515,N_27449);
xnor U27914 (N_27914,N_27548,N_26760);
xnor U27915 (N_27915,N_27335,N_27129);
nand U27916 (N_27916,N_26613,N_26433);
nor U27917 (N_27917,N_26727,N_27463);
and U27918 (N_27918,N_26803,N_26633);
nor U27919 (N_27919,N_26997,N_27139);
and U27920 (N_27920,N_27368,N_26606);
nor U27921 (N_27921,N_27037,N_27084);
and U27922 (N_27922,N_26609,N_26493);
or U27923 (N_27923,N_26474,N_27137);
or U27924 (N_27924,N_26967,N_27248);
or U27925 (N_27925,N_26548,N_27595);
nand U27926 (N_27926,N_26988,N_27343);
xnor U27927 (N_27927,N_26561,N_27386);
nand U27928 (N_27928,N_26714,N_27436);
and U27929 (N_27929,N_26663,N_26503);
nand U27930 (N_27930,N_26809,N_26910);
nand U27931 (N_27931,N_27230,N_27094);
nand U27932 (N_27932,N_27433,N_26949);
nand U27933 (N_27933,N_26854,N_27086);
and U27934 (N_27934,N_26952,N_26946);
xor U27935 (N_27935,N_27070,N_26726);
and U27936 (N_27936,N_27427,N_26970);
or U27937 (N_27937,N_26652,N_26587);
and U27938 (N_27938,N_26682,N_27117);
xnor U27939 (N_27939,N_27116,N_26597);
xor U27940 (N_27940,N_26878,N_26747);
or U27941 (N_27941,N_26756,N_26735);
nand U27942 (N_27942,N_27349,N_26651);
and U27943 (N_27943,N_27029,N_27528);
nor U27944 (N_27944,N_26793,N_27517);
or U27945 (N_27945,N_26432,N_26991);
xnor U27946 (N_27946,N_26577,N_26999);
or U27947 (N_27947,N_26996,N_26582);
nand U27948 (N_27948,N_27203,N_27301);
and U27949 (N_27949,N_27492,N_26840);
nand U27950 (N_27950,N_27242,N_26608);
nor U27951 (N_27951,N_26774,N_27050);
or U27952 (N_27952,N_26671,N_26604);
and U27953 (N_27953,N_26925,N_26599);
or U27954 (N_27954,N_27366,N_27170);
nand U27955 (N_27955,N_27502,N_26995);
nor U27956 (N_27956,N_27450,N_26722);
xnor U27957 (N_27957,N_26431,N_26823);
nor U27958 (N_27958,N_27559,N_26621);
or U27959 (N_27959,N_26943,N_26457);
nand U27960 (N_27960,N_27348,N_26528);
nand U27961 (N_27961,N_27532,N_26639);
nor U27962 (N_27962,N_27456,N_26842);
nand U27963 (N_27963,N_26766,N_27049);
and U27964 (N_27964,N_27377,N_26794);
nor U27965 (N_27965,N_27409,N_26447);
and U27966 (N_27966,N_27006,N_27071);
nand U27967 (N_27967,N_27096,N_27536);
nand U27968 (N_27968,N_26451,N_26498);
nand U27969 (N_27969,N_27140,N_26629);
xor U27970 (N_27970,N_26460,N_26638);
nand U27971 (N_27971,N_26804,N_27051);
xnor U27972 (N_27972,N_26713,N_27270);
nor U27973 (N_27973,N_26905,N_26562);
or U27974 (N_27974,N_27166,N_26654);
nand U27975 (N_27975,N_26411,N_26736);
xor U27976 (N_27976,N_26825,N_27034);
and U27977 (N_27977,N_27523,N_27576);
nand U27978 (N_27978,N_27200,N_27289);
or U27979 (N_27979,N_27568,N_26757);
xor U27980 (N_27980,N_27406,N_27079);
nand U27981 (N_27981,N_27411,N_27437);
and U27982 (N_27982,N_26700,N_26427);
or U27983 (N_27983,N_26511,N_26876);
and U27984 (N_27984,N_26647,N_27115);
nand U27985 (N_27985,N_26771,N_27237);
and U27986 (N_27986,N_27207,N_26572);
xnor U27987 (N_27987,N_26507,N_27057);
xor U27988 (N_27988,N_27418,N_26832);
and U27989 (N_27989,N_27205,N_27526);
and U27990 (N_27990,N_26914,N_26412);
nand U27991 (N_27991,N_27153,N_27286);
nor U27992 (N_27992,N_27314,N_27043);
or U27993 (N_27993,N_27496,N_27476);
xnor U27994 (N_27994,N_27577,N_26401);
nor U27995 (N_27995,N_27184,N_26472);
or U27996 (N_27996,N_27175,N_26998);
and U27997 (N_27997,N_27396,N_26775);
xor U27998 (N_27998,N_27429,N_26416);
nor U27999 (N_27999,N_27221,N_26645);
nand U28000 (N_28000,N_27092,N_26819);
xor U28001 (N_28001,N_27062,N_26821);
xor U28002 (N_28002,N_26537,N_27387);
and U28003 (N_28003,N_27365,N_27339);
and U28004 (N_28004,N_27244,N_27522);
xor U28005 (N_28005,N_26900,N_27125);
xnor U28006 (N_28006,N_26734,N_27080);
nand U28007 (N_28007,N_27421,N_27243);
or U28008 (N_28008,N_27402,N_26524);
xor U28009 (N_28009,N_26514,N_27104);
and U28010 (N_28010,N_27398,N_26464);
nand U28011 (N_28011,N_26926,N_26705);
or U28012 (N_28012,N_27407,N_26928);
nand U28013 (N_28013,N_26918,N_26478);
or U28014 (N_28014,N_27304,N_26919);
nor U28015 (N_28015,N_27087,N_26867);
xor U28016 (N_28016,N_27477,N_27459);
xnor U28017 (N_28017,N_27596,N_26624);
or U28018 (N_28018,N_27324,N_27491);
or U28019 (N_28019,N_26680,N_26890);
xnor U28020 (N_28020,N_26755,N_27556);
nand U28021 (N_28021,N_26494,N_26687);
and U28022 (N_28022,N_27192,N_27482);
xnor U28023 (N_28023,N_27587,N_26591);
xor U28024 (N_28024,N_27111,N_26787);
and U28025 (N_28025,N_26434,N_27124);
or U28026 (N_28026,N_27143,N_27404);
nand U28027 (N_28027,N_26450,N_26659);
nand U28028 (N_28028,N_27151,N_27527);
nand U28029 (N_28029,N_26686,N_27004);
xor U28030 (N_28030,N_26742,N_26779);
nand U28031 (N_28031,N_27494,N_26440);
and U28032 (N_28032,N_27228,N_26571);
or U28033 (N_28033,N_27578,N_27291);
nor U28034 (N_28034,N_27159,N_27325);
nor U28035 (N_28035,N_27439,N_26947);
nand U28036 (N_28036,N_27074,N_26452);
nand U28037 (N_28037,N_26565,N_26594);
nor U28038 (N_28038,N_26477,N_27485);
xor U28039 (N_28039,N_26541,N_26469);
or U28040 (N_28040,N_27138,N_26861);
nor U28041 (N_28041,N_27178,N_26812);
nand U28042 (N_28042,N_27425,N_26672);
or U28043 (N_28043,N_27495,N_26778);
nor U28044 (N_28044,N_26977,N_27537);
xnor U28045 (N_28045,N_27543,N_26513);
nand U28046 (N_28046,N_26711,N_26549);
nand U28047 (N_28047,N_27512,N_27145);
or U28048 (N_28048,N_26879,N_26491);
nand U28049 (N_28049,N_26909,N_27142);
and U28050 (N_28050,N_27430,N_27179);
nor U28051 (N_28051,N_27023,N_26922);
xnor U28052 (N_28052,N_26955,N_26806);
xnor U28053 (N_28053,N_27551,N_27259);
and U28054 (N_28054,N_26754,N_27232);
xor U28055 (N_28055,N_27458,N_27039);
or U28056 (N_28056,N_27319,N_26780);
nor U28057 (N_28057,N_27225,N_26994);
and U28058 (N_28058,N_26673,N_26693);
or U28059 (N_28059,N_26546,N_27260);
nand U28060 (N_28060,N_26920,N_26975);
or U28061 (N_28061,N_27529,N_26865);
or U28062 (N_28062,N_27516,N_26504);
nor U28063 (N_28063,N_27100,N_26820);
xnor U28064 (N_28064,N_27044,N_26635);
xnor U28065 (N_28065,N_26579,N_26888);
or U28066 (N_28066,N_27464,N_26846);
nand U28067 (N_28067,N_27017,N_27015);
or U28068 (N_28068,N_26984,N_26911);
and U28069 (N_28069,N_26677,N_27239);
nand U28070 (N_28070,N_26667,N_26855);
nor U28071 (N_28071,N_26719,N_27021);
nor U28072 (N_28072,N_27465,N_27434);
nand U28073 (N_28073,N_26786,N_26871);
and U28074 (N_28074,N_27561,N_27160);
or U28075 (N_28075,N_27198,N_26732);
xnor U28076 (N_28076,N_26422,N_27320);
or U28077 (N_28077,N_26930,N_26857);
nand U28078 (N_28078,N_26429,N_27490);
xnor U28079 (N_28079,N_26841,N_26731);
and U28080 (N_28080,N_27164,N_26576);
and U28081 (N_28081,N_26642,N_26512);
and U28082 (N_28082,N_27167,N_26487);
nor U28083 (N_28083,N_26948,N_27081);
nand U28084 (N_28084,N_26448,N_27257);
nor U28085 (N_28085,N_26940,N_26762);
and U28086 (N_28086,N_27148,N_27108);
and U28087 (N_28087,N_26882,N_27123);
nor U28088 (N_28088,N_27099,N_26408);
xor U28089 (N_28089,N_26625,N_26773);
or U28090 (N_28090,N_27563,N_26981);
or U28091 (N_28091,N_26445,N_27083);
and U28092 (N_28092,N_26539,N_26873);
xnor U28093 (N_28093,N_27264,N_27379);
and U28094 (N_28094,N_27238,N_26699);
xor U28095 (N_28095,N_26834,N_26568);
and U28096 (N_28096,N_26707,N_26423);
nand U28097 (N_28097,N_27038,N_27507);
nand U28098 (N_28098,N_26649,N_26744);
and U28099 (N_28099,N_26833,N_27273);
xor U28100 (N_28100,N_27448,N_26455);
xnor U28101 (N_28101,N_26650,N_27290);
or U28102 (N_28102,N_27052,N_27020);
or U28103 (N_28103,N_27564,N_27134);
or U28104 (N_28104,N_27509,N_27282);
or U28105 (N_28105,N_27392,N_27432);
xor U28106 (N_28106,N_26765,N_26588);
nand U28107 (N_28107,N_27367,N_26622);
nand U28108 (N_28108,N_27306,N_27462);
nand U28109 (N_28109,N_26441,N_26750);
and U28110 (N_28110,N_26752,N_26887);
or U28111 (N_28111,N_26643,N_26982);
nand U28112 (N_28112,N_26957,N_26595);
nor U28113 (N_28113,N_26815,N_27018);
nor U28114 (N_28114,N_27182,N_26458);
or U28115 (N_28115,N_27481,N_26923);
or U28116 (N_28116,N_27584,N_27498);
nor U28117 (N_28117,N_27161,N_26738);
and U28118 (N_28118,N_26898,N_27454);
nor U28119 (N_28119,N_26413,N_27318);
and U28120 (N_28120,N_27222,N_26817);
and U28121 (N_28121,N_26795,N_26612);
xor U28122 (N_28122,N_26904,N_26563);
nor U28123 (N_28123,N_26557,N_26929);
nand U28124 (N_28124,N_26935,N_26960);
nor U28125 (N_28125,N_27435,N_27269);
nor U28126 (N_28126,N_27395,N_26751);
nor U28127 (N_28127,N_26798,N_26670);
and U28128 (N_28128,N_26534,N_27209);
nand U28129 (N_28129,N_26603,N_27249);
and U28130 (N_28130,N_27531,N_27428);
nand U28131 (N_28131,N_27589,N_27442);
or U28132 (N_28132,N_26917,N_26640);
and U28133 (N_28133,N_26802,N_27189);
nor U28134 (N_28134,N_26614,N_27103);
or U28135 (N_28135,N_26630,N_27261);
or U28136 (N_28136,N_27501,N_27263);
and U28137 (N_28137,N_27385,N_26758);
nand U28138 (N_28138,N_27574,N_26535);
nor U28139 (N_28139,N_26710,N_27149);
nand U28140 (N_28140,N_27378,N_27417);
nor U28141 (N_28141,N_26709,N_26958);
and U28142 (N_28142,N_27582,N_26592);
nand U28143 (N_28143,N_26578,N_27469);
or U28144 (N_28144,N_27506,N_26811);
xnor U28145 (N_28145,N_27283,N_26860);
or U28146 (N_28146,N_27144,N_27583);
nand U28147 (N_28147,N_26428,N_26937);
nor U28148 (N_28148,N_26884,N_27508);
nand U28149 (N_28149,N_27174,N_26545);
and U28150 (N_28150,N_27488,N_26439);
nand U28151 (N_28151,N_27219,N_26808);
or U28152 (N_28152,N_27567,N_27515);
and U28153 (N_28153,N_27256,N_26792);
nor U28154 (N_28154,N_27340,N_26593);
nand U28155 (N_28155,N_26465,N_26473);
nand U28156 (N_28156,N_27119,N_26406);
xor U28157 (N_28157,N_26584,N_27388);
or U28158 (N_28158,N_27489,N_26872);
or U28159 (N_28159,N_26889,N_26637);
nor U28160 (N_28160,N_26583,N_26490);
nor U28161 (N_28161,N_27191,N_26950);
nor U28162 (N_28162,N_27246,N_26913);
xnor U28163 (N_28163,N_26866,N_27310);
and U28164 (N_28164,N_26915,N_27223);
and U28165 (N_28165,N_26674,N_27121);
nand U28166 (N_28166,N_27350,N_27202);
nor U28167 (N_28167,N_27479,N_26506);
or U28168 (N_28168,N_27560,N_26547);
nand U28169 (N_28169,N_26532,N_26859);
nor U28170 (N_28170,N_27101,N_27027);
and U28171 (N_28171,N_26575,N_26486);
or U28172 (N_28172,N_26716,N_26676);
and U28173 (N_28173,N_26932,N_27323);
and U28174 (N_28174,N_27452,N_27136);
nor U28175 (N_28175,N_26968,N_27040);
or U28176 (N_28176,N_27060,N_26965);
nor U28177 (N_28177,N_26405,N_26839);
nor U28178 (N_28178,N_26936,N_26826);
or U28179 (N_28179,N_26954,N_26573);
and U28180 (N_28180,N_26410,N_26864);
and U28181 (N_28181,N_27132,N_26602);
or U28182 (N_28182,N_27334,N_27562);
and U28183 (N_28183,N_26615,N_27539);
xnor U28184 (N_28184,N_26912,N_26927);
nand U28185 (N_28185,N_27359,N_26618);
nand U28186 (N_28186,N_27180,N_27565);
nor U28187 (N_28187,N_27183,N_27329);
xnor U28188 (N_28188,N_27091,N_26527);
nor U28189 (N_28189,N_26805,N_27268);
xnor U28190 (N_28190,N_27262,N_26720);
nor U28191 (N_28191,N_27147,N_27214);
nand U28192 (N_28192,N_27426,N_27408);
xnor U28193 (N_28193,N_26694,N_26767);
or U28194 (N_28194,N_26552,N_27400);
xnor U28195 (N_28195,N_27468,N_26739);
nand U28196 (N_28196,N_27036,N_26993);
nand U28197 (N_28197,N_27302,N_26543);
or U28198 (N_28198,N_27267,N_27570);
nand U28199 (N_28199,N_27120,N_27533);
nor U28200 (N_28200,N_26994,N_27376);
nor U28201 (N_28201,N_26895,N_27093);
nand U28202 (N_28202,N_26517,N_27112);
and U28203 (N_28203,N_26764,N_27073);
nor U28204 (N_28204,N_26702,N_27177);
or U28205 (N_28205,N_27431,N_27085);
nor U28206 (N_28206,N_26911,N_27365);
nor U28207 (N_28207,N_26589,N_27028);
or U28208 (N_28208,N_27409,N_27515);
nand U28209 (N_28209,N_26847,N_27340);
and U28210 (N_28210,N_27128,N_27480);
or U28211 (N_28211,N_26767,N_26649);
nand U28212 (N_28212,N_26569,N_26568);
and U28213 (N_28213,N_27199,N_26676);
and U28214 (N_28214,N_27456,N_26451);
nor U28215 (N_28215,N_27010,N_27412);
nor U28216 (N_28216,N_26532,N_27101);
and U28217 (N_28217,N_26963,N_26710);
nand U28218 (N_28218,N_26772,N_26898);
nor U28219 (N_28219,N_27489,N_26536);
xor U28220 (N_28220,N_27559,N_27455);
xnor U28221 (N_28221,N_26674,N_26809);
or U28222 (N_28222,N_27115,N_27203);
nor U28223 (N_28223,N_26626,N_26480);
and U28224 (N_28224,N_27167,N_26407);
xnor U28225 (N_28225,N_26976,N_26974);
or U28226 (N_28226,N_27358,N_26991);
nor U28227 (N_28227,N_26775,N_26979);
nand U28228 (N_28228,N_26638,N_26828);
or U28229 (N_28229,N_27065,N_26744);
nand U28230 (N_28230,N_26996,N_27354);
and U28231 (N_28231,N_26718,N_27515);
and U28232 (N_28232,N_26942,N_26508);
nor U28233 (N_28233,N_27151,N_26808);
or U28234 (N_28234,N_27237,N_26585);
or U28235 (N_28235,N_26633,N_27312);
xnor U28236 (N_28236,N_26962,N_26487);
nand U28237 (N_28237,N_27443,N_27256);
xor U28238 (N_28238,N_27380,N_27017);
nand U28239 (N_28239,N_27401,N_26505);
nand U28240 (N_28240,N_26555,N_26889);
nor U28241 (N_28241,N_26972,N_26731);
nor U28242 (N_28242,N_27156,N_26808);
or U28243 (N_28243,N_26905,N_26946);
and U28244 (N_28244,N_27450,N_27134);
xnor U28245 (N_28245,N_26779,N_27459);
nand U28246 (N_28246,N_27231,N_27210);
and U28247 (N_28247,N_27248,N_27186);
nor U28248 (N_28248,N_27113,N_27088);
or U28249 (N_28249,N_26651,N_26700);
and U28250 (N_28250,N_27592,N_26980);
nor U28251 (N_28251,N_27479,N_27558);
or U28252 (N_28252,N_27255,N_26493);
and U28253 (N_28253,N_27006,N_27131);
and U28254 (N_28254,N_26831,N_26830);
nand U28255 (N_28255,N_26784,N_26422);
nand U28256 (N_28256,N_27363,N_27003);
or U28257 (N_28257,N_26971,N_27014);
nor U28258 (N_28258,N_27498,N_26962);
nor U28259 (N_28259,N_27022,N_26994);
nand U28260 (N_28260,N_27146,N_27195);
or U28261 (N_28261,N_26404,N_26522);
and U28262 (N_28262,N_26703,N_26433);
nand U28263 (N_28263,N_27147,N_27278);
and U28264 (N_28264,N_26914,N_27496);
nand U28265 (N_28265,N_27566,N_26954);
and U28266 (N_28266,N_27012,N_26930);
or U28267 (N_28267,N_27519,N_27580);
and U28268 (N_28268,N_27007,N_26420);
xnor U28269 (N_28269,N_26859,N_27013);
and U28270 (N_28270,N_27151,N_26900);
nand U28271 (N_28271,N_27479,N_26890);
xor U28272 (N_28272,N_26545,N_27592);
and U28273 (N_28273,N_26562,N_27443);
or U28274 (N_28274,N_26760,N_26775);
xor U28275 (N_28275,N_27528,N_26859);
and U28276 (N_28276,N_26885,N_26554);
xor U28277 (N_28277,N_27580,N_26575);
nand U28278 (N_28278,N_26821,N_26953);
nand U28279 (N_28279,N_26799,N_26651);
xor U28280 (N_28280,N_27403,N_26706);
and U28281 (N_28281,N_27332,N_27238);
xnor U28282 (N_28282,N_26742,N_27147);
or U28283 (N_28283,N_26545,N_26985);
or U28284 (N_28284,N_27469,N_27528);
or U28285 (N_28285,N_26797,N_27538);
and U28286 (N_28286,N_26869,N_27318);
nand U28287 (N_28287,N_27520,N_26589);
nor U28288 (N_28288,N_27034,N_27318);
or U28289 (N_28289,N_27018,N_26449);
nand U28290 (N_28290,N_27040,N_26996);
nand U28291 (N_28291,N_27336,N_27206);
and U28292 (N_28292,N_27435,N_27168);
nor U28293 (N_28293,N_26750,N_26595);
nand U28294 (N_28294,N_27053,N_27054);
and U28295 (N_28295,N_26579,N_26871);
or U28296 (N_28296,N_26425,N_26897);
nor U28297 (N_28297,N_26405,N_26935);
and U28298 (N_28298,N_27532,N_27373);
or U28299 (N_28299,N_27207,N_26950);
or U28300 (N_28300,N_26998,N_26883);
and U28301 (N_28301,N_26907,N_27082);
or U28302 (N_28302,N_26841,N_26801);
and U28303 (N_28303,N_27180,N_26695);
and U28304 (N_28304,N_27084,N_27255);
and U28305 (N_28305,N_26585,N_26557);
nor U28306 (N_28306,N_27183,N_27244);
xnor U28307 (N_28307,N_27274,N_26580);
nand U28308 (N_28308,N_27536,N_26952);
or U28309 (N_28309,N_26831,N_27517);
xnor U28310 (N_28310,N_27237,N_26553);
xnor U28311 (N_28311,N_27397,N_26901);
nor U28312 (N_28312,N_27145,N_27247);
or U28313 (N_28313,N_27381,N_27436);
and U28314 (N_28314,N_27243,N_26648);
or U28315 (N_28315,N_26495,N_26910);
xor U28316 (N_28316,N_27306,N_26440);
nor U28317 (N_28317,N_27052,N_26970);
xnor U28318 (N_28318,N_26693,N_26886);
xnor U28319 (N_28319,N_27045,N_26788);
xor U28320 (N_28320,N_26729,N_27000);
nor U28321 (N_28321,N_26420,N_26733);
and U28322 (N_28322,N_26602,N_26844);
and U28323 (N_28323,N_26636,N_27455);
and U28324 (N_28324,N_26418,N_26523);
nor U28325 (N_28325,N_27241,N_27162);
or U28326 (N_28326,N_27199,N_27509);
nor U28327 (N_28327,N_27307,N_27457);
nor U28328 (N_28328,N_27114,N_26950);
nand U28329 (N_28329,N_26430,N_26916);
nor U28330 (N_28330,N_26703,N_27370);
and U28331 (N_28331,N_27591,N_26828);
and U28332 (N_28332,N_27098,N_26474);
and U28333 (N_28333,N_26756,N_26507);
xor U28334 (N_28334,N_27311,N_27520);
or U28335 (N_28335,N_27523,N_26562);
and U28336 (N_28336,N_26431,N_27179);
nand U28337 (N_28337,N_26653,N_26609);
xor U28338 (N_28338,N_26994,N_26516);
and U28339 (N_28339,N_27107,N_26973);
nand U28340 (N_28340,N_27294,N_27579);
nor U28341 (N_28341,N_27230,N_26720);
and U28342 (N_28342,N_26816,N_27576);
nor U28343 (N_28343,N_26506,N_27257);
xnor U28344 (N_28344,N_26605,N_27032);
or U28345 (N_28345,N_27165,N_27474);
nand U28346 (N_28346,N_26414,N_26743);
or U28347 (N_28347,N_26691,N_27207);
nor U28348 (N_28348,N_26461,N_27471);
or U28349 (N_28349,N_26734,N_27136);
nand U28350 (N_28350,N_27248,N_26643);
nand U28351 (N_28351,N_27017,N_26516);
and U28352 (N_28352,N_27464,N_26869);
or U28353 (N_28353,N_27008,N_27349);
xor U28354 (N_28354,N_27575,N_26891);
nand U28355 (N_28355,N_27014,N_26863);
xnor U28356 (N_28356,N_27209,N_27039);
xnor U28357 (N_28357,N_27519,N_27420);
nand U28358 (N_28358,N_26584,N_26412);
xor U28359 (N_28359,N_27378,N_26930);
or U28360 (N_28360,N_26592,N_26929);
or U28361 (N_28361,N_27346,N_27147);
or U28362 (N_28362,N_26667,N_27064);
xor U28363 (N_28363,N_27243,N_27496);
nand U28364 (N_28364,N_26799,N_26897);
xor U28365 (N_28365,N_27330,N_26499);
nor U28366 (N_28366,N_27239,N_26957);
or U28367 (N_28367,N_26793,N_26469);
nand U28368 (N_28368,N_27231,N_27225);
or U28369 (N_28369,N_27419,N_26767);
nor U28370 (N_28370,N_27206,N_27455);
nor U28371 (N_28371,N_27432,N_26544);
xor U28372 (N_28372,N_26947,N_26550);
or U28373 (N_28373,N_27546,N_26628);
or U28374 (N_28374,N_26726,N_26658);
xor U28375 (N_28375,N_26902,N_27529);
nand U28376 (N_28376,N_26690,N_27322);
xnor U28377 (N_28377,N_26454,N_26962);
and U28378 (N_28378,N_27450,N_26521);
and U28379 (N_28379,N_26583,N_26611);
and U28380 (N_28380,N_26664,N_27477);
nor U28381 (N_28381,N_26528,N_27497);
nor U28382 (N_28382,N_26777,N_27318);
or U28383 (N_28383,N_27502,N_27001);
xnor U28384 (N_28384,N_26404,N_27471);
xor U28385 (N_28385,N_26933,N_27087);
and U28386 (N_28386,N_26595,N_26940);
or U28387 (N_28387,N_26908,N_26806);
nand U28388 (N_28388,N_26800,N_27313);
or U28389 (N_28389,N_26579,N_26825);
and U28390 (N_28390,N_26980,N_26896);
or U28391 (N_28391,N_27553,N_26634);
or U28392 (N_28392,N_26709,N_27296);
and U28393 (N_28393,N_27381,N_26726);
and U28394 (N_28394,N_26411,N_26464);
and U28395 (N_28395,N_26550,N_26512);
nand U28396 (N_28396,N_27523,N_26441);
xnor U28397 (N_28397,N_27573,N_26873);
or U28398 (N_28398,N_26785,N_27587);
nor U28399 (N_28399,N_26558,N_27574);
and U28400 (N_28400,N_27365,N_27400);
nand U28401 (N_28401,N_26494,N_27346);
nor U28402 (N_28402,N_27024,N_27393);
nor U28403 (N_28403,N_27203,N_26726);
xnor U28404 (N_28404,N_26754,N_26880);
nor U28405 (N_28405,N_27224,N_27529);
nor U28406 (N_28406,N_27451,N_27294);
xor U28407 (N_28407,N_26780,N_26961);
and U28408 (N_28408,N_27167,N_26673);
and U28409 (N_28409,N_26948,N_27431);
and U28410 (N_28410,N_27559,N_26469);
nand U28411 (N_28411,N_27061,N_26625);
and U28412 (N_28412,N_26807,N_26447);
or U28413 (N_28413,N_26652,N_26576);
and U28414 (N_28414,N_27166,N_26865);
or U28415 (N_28415,N_26955,N_27108);
and U28416 (N_28416,N_27131,N_27214);
nand U28417 (N_28417,N_26547,N_26897);
nor U28418 (N_28418,N_27594,N_26606);
nand U28419 (N_28419,N_27346,N_27094);
nor U28420 (N_28420,N_26814,N_26595);
or U28421 (N_28421,N_27130,N_26460);
or U28422 (N_28422,N_27127,N_26406);
nor U28423 (N_28423,N_27331,N_26976);
xor U28424 (N_28424,N_27531,N_27097);
nor U28425 (N_28425,N_26947,N_26501);
xor U28426 (N_28426,N_26452,N_26652);
xnor U28427 (N_28427,N_26540,N_26816);
and U28428 (N_28428,N_27368,N_27292);
nor U28429 (N_28429,N_26671,N_27281);
xor U28430 (N_28430,N_26921,N_27386);
nor U28431 (N_28431,N_26546,N_27164);
nand U28432 (N_28432,N_26984,N_26706);
xor U28433 (N_28433,N_27064,N_27256);
xor U28434 (N_28434,N_27290,N_27118);
nor U28435 (N_28435,N_26893,N_26980);
or U28436 (N_28436,N_26512,N_27088);
xor U28437 (N_28437,N_27248,N_26585);
and U28438 (N_28438,N_27320,N_27501);
xor U28439 (N_28439,N_27115,N_27067);
xnor U28440 (N_28440,N_26440,N_27146);
xnor U28441 (N_28441,N_26764,N_27428);
nor U28442 (N_28442,N_27212,N_27366);
nand U28443 (N_28443,N_27306,N_27189);
or U28444 (N_28444,N_27542,N_26617);
or U28445 (N_28445,N_26484,N_27310);
and U28446 (N_28446,N_26775,N_26541);
nand U28447 (N_28447,N_27235,N_27047);
and U28448 (N_28448,N_26704,N_27057);
nand U28449 (N_28449,N_27399,N_27011);
or U28450 (N_28450,N_27406,N_27481);
or U28451 (N_28451,N_27565,N_26810);
and U28452 (N_28452,N_27029,N_26635);
or U28453 (N_28453,N_26672,N_27204);
and U28454 (N_28454,N_26561,N_27336);
nand U28455 (N_28455,N_26813,N_27432);
xnor U28456 (N_28456,N_26892,N_26558);
nand U28457 (N_28457,N_27079,N_27525);
nor U28458 (N_28458,N_27400,N_26453);
or U28459 (N_28459,N_27527,N_26849);
or U28460 (N_28460,N_26666,N_26772);
and U28461 (N_28461,N_26571,N_27578);
and U28462 (N_28462,N_27458,N_26942);
nor U28463 (N_28463,N_26937,N_27023);
nor U28464 (N_28464,N_27530,N_26445);
nand U28465 (N_28465,N_27322,N_26944);
nor U28466 (N_28466,N_27058,N_27021);
nor U28467 (N_28467,N_27541,N_27496);
nor U28468 (N_28468,N_26781,N_27122);
nand U28469 (N_28469,N_26902,N_27156);
xnor U28470 (N_28470,N_27406,N_26850);
xor U28471 (N_28471,N_26627,N_27318);
xor U28472 (N_28472,N_27354,N_27326);
xnor U28473 (N_28473,N_27376,N_26859);
xor U28474 (N_28474,N_26886,N_27147);
xor U28475 (N_28475,N_27421,N_27098);
xnor U28476 (N_28476,N_26743,N_27460);
and U28477 (N_28477,N_26564,N_27260);
or U28478 (N_28478,N_27328,N_27462);
nor U28479 (N_28479,N_27366,N_27336);
and U28480 (N_28480,N_26751,N_26827);
nor U28481 (N_28481,N_27007,N_27190);
nor U28482 (N_28482,N_26862,N_27482);
and U28483 (N_28483,N_26985,N_26847);
and U28484 (N_28484,N_27301,N_26617);
xnor U28485 (N_28485,N_26570,N_26738);
or U28486 (N_28486,N_26454,N_27277);
xor U28487 (N_28487,N_26632,N_27463);
nand U28488 (N_28488,N_26649,N_26412);
nor U28489 (N_28489,N_26671,N_26695);
xor U28490 (N_28490,N_27168,N_27129);
xnor U28491 (N_28491,N_26626,N_26520);
nor U28492 (N_28492,N_26598,N_27132);
xor U28493 (N_28493,N_27407,N_26811);
nor U28494 (N_28494,N_27440,N_27252);
nand U28495 (N_28495,N_27466,N_27555);
or U28496 (N_28496,N_27249,N_26599);
xor U28497 (N_28497,N_27388,N_26678);
nor U28498 (N_28498,N_26846,N_26969);
nor U28499 (N_28499,N_27058,N_26802);
nand U28500 (N_28500,N_26809,N_27011);
nand U28501 (N_28501,N_26675,N_27508);
nand U28502 (N_28502,N_27045,N_26553);
xor U28503 (N_28503,N_26971,N_27583);
xnor U28504 (N_28504,N_27229,N_27038);
nand U28505 (N_28505,N_27095,N_27519);
or U28506 (N_28506,N_27208,N_27241);
and U28507 (N_28507,N_26871,N_26683);
or U28508 (N_28508,N_27142,N_26867);
nor U28509 (N_28509,N_26569,N_26953);
or U28510 (N_28510,N_26426,N_27106);
nand U28511 (N_28511,N_26507,N_27463);
nor U28512 (N_28512,N_27371,N_26915);
or U28513 (N_28513,N_26935,N_27076);
nand U28514 (N_28514,N_26755,N_27113);
and U28515 (N_28515,N_26575,N_26436);
and U28516 (N_28516,N_26568,N_26800);
or U28517 (N_28517,N_26687,N_26523);
nand U28518 (N_28518,N_27059,N_26826);
nor U28519 (N_28519,N_27182,N_26629);
nor U28520 (N_28520,N_26532,N_27131);
and U28521 (N_28521,N_27353,N_27209);
nand U28522 (N_28522,N_27153,N_27579);
nand U28523 (N_28523,N_27148,N_27236);
xnor U28524 (N_28524,N_27231,N_27589);
and U28525 (N_28525,N_26401,N_27401);
xnor U28526 (N_28526,N_27181,N_27519);
xnor U28527 (N_28527,N_27343,N_27491);
xnor U28528 (N_28528,N_26403,N_26618);
or U28529 (N_28529,N_26686,N_26709);
and U28530 (N_28530,N_27542,N_26417);
or U28531 (N_28531,N_27093,N_26509);
nand U28532 (N_28532,N_26912,N_26673);
xnor U28533 (N_28533,N_27464,N_27567);
nand U28534 (N_28534,N_27444,N_27131);
xnor U28535 (N_28535,N_26476,N_26765);
nand U28536 (N_28536,N_27236,N_26673);
or U28537 (N_28537,N_26559,N_26599);
nand U28538 (N_28538,N_27392,N_27195);
or U28539 (N_28539,N_26558,N_27401);
or U28540 (N_28540,N_26484,N_26482);
or U28541 (N_28541,N_26975,N_26604);
or U28542 (N_28542,N_27585,N_27231);
nand U28543 (N_28543,N_26492,N_26609);
nand U28544 (N_28544,N_26645,N_27537);
nor U28545 (N_28545,N_26570,N_27040);
xor U28546 (N_28546,N_26572,N_26784);
xor U28547 (N_28547,N_26882,N_26742);
nand U28548 (N_28548,N_27081,N_27584);
nand U28549 (N_28549,N_27545,N_26409);
and U28550 (N_28550,N_27375,N_26529);
nand U28551 (N_28551,N_26879,N_26906);
xor U28552 (N_28552,N_27173,N_27587);
nor U28553 (N_28553,N_26835,N_26847);
xnor U28554 (N_28554,N_26831,N_26839);
nand U28555 (N_28555,N_27142,N_27074);
and U28556 (N_28556,N_27257,N_26970);
nor U28557 (N_28557,N_26744,N_26477);
and U28558 (N_28558,N_26676,N_26798);
and U28559 (N_28559,N_26766,N_26653);
nand U28560 (N_28560,N_27205,N_26479);
xnor U28561 (N_28561,N_27209,N_26594);
or U28562 (N_28562,N_26455,N_27246);
xnor U28563 (N_28563,N_26533,N_26812);
nor U28564 (N_28564,N_26673,N_27047);
and U28565 (N_28565,N_26763,N_27271);
xor U28566 (N_28566,N_27537,N_26867);
and U28567 (N_28567,N_26867,N_27424);
and U28568 (N_28568,N_27190,N_26730);
nor U28569 (N_28569,N_26798,N_27337);
nand U28570 (N_28570,N_26630,N_27295);
xnor U28571 (N_28571,N_27074,N_26460);
or U28572 (N_28572,N_26529,N_26550);
xor U28573 (N_28573,N_27002,N_27572);
xnor U28574 (N_28574,N_27568,N_26642);
xor U28575 (N_28575,N_27020,N_27193);
nand U28576 (N_28576,N_27075,N_26717);
nand U28577 (N_28577,N_26816,N_26780);
xor U28578 (N_28578,N_27249,N_27101);
nor U28579 (N_28579,N_27328,N_27550);
nor U28580 (N_28580,N_27193,N_27578);
xor U28581 (N_28581,N_27593,N_27074);
xnor U28582 (N_28582,N_27549,N_27310);
xnor U28583 (N_28583,N_27153,N_26747);
or U28584 (N_28584,N_26948,N_27234);
nor U28585 (N_28585,N_26550,N_26511);
and U28586 (N_28586,N_26648,N_27322);
or U28587 (N_28587,N_26930,N_27526);
nand U28588 (N_28588,N_27229,N_26849);
nor U28589 (N_28589,N_26688,N_26525);
xor U28590 (N_28590,N_26467,N_27058);
and U28591 (N_28591,N_26442,N_27357);
and U28592 (N_28592,N_27033,N_27066);
or U28593 (N_28593,N_27268,N_26753);
and U28594 (N_28594,N_27365,N_27371);
nand U28595 (N_28595,N_26450,N_26864);
or U28596 (N_28596,N_26678,N_27484);
and U28597 (N_28597,N_27195,N_27236);
nand U28598 (N_28598,N_26553,N_26790);
xor U28599 (N_28599,N_27587,N_26602);
or U28600 (N_28600,N_27489,N_26473);
xor U28601 (N_28601,N_27071,N_27349);
nor U28602 (N_28602,N_27505,N_26929);
nand U28603 (N_28603,N_26750,N_26927);
nor U28604 (N_28604,N_27250,N_26927);
nor U28605 (N_28605,N_27345,N_27351);
nand U28606 (N_28606,N_26892,N_26433);
xnor U28607 (N_28607,N_27049,N_27089);
and U28608 (N_28608,N_27425,N_26935);
nor U28609 (N_28609,N_26876,N_27069);
or U28610 (N_28610,N_27310,N_27357);
nor U28611 (N_28611,N_26659,N_27083);
nand U28612 (N_28612,N_27279,N_27208);
nand U28613 (N_28613,N_26427,N_27048);
xor U28614 (N_28614,N_27197,N_27397);
xor U28615 (N_28615,N_27040,N_26970);
nand U28616 (N_28616,N_27261,N_27585);
or U28617 (N_28617,N_26962,N_27439);
or U28618 (N_28618,N_27236,N_26834);
nand U28619 (N_28619,N_27267,N_27280);
nor U28620 (N_28620,N_26417,N_27386);
xor U28621 (N_28621,N_26990,N_27106);
nand U28622 (N_28622,N_27373,N_26763);
xor U28623 (N_28623,N_26889,N_26422);
xnor U28624 (N_28624,N_27534,N_26622);
nor U28625 (N_28625,N_27274,N_27445);
xnor U28626 (N_28626,N_26934,N_27408);
nand U28627 (N_28627,N_26631,N_27288);
nand U28628 (N_28628,N_26596,N_27504);
or U28629 (N_28629,N_27219,N_26673);
nand U28630 (N_28630,N_27561,N_26923);
and U28631 (N_28631,N_26995,N_26934);
and U28632 (N_28632,N_27237,N_26668);
or U28633 (N_28633,N_26705,N_27221);
xor U28634 (N_28634,N_27321,N_26867);
nor U28635 (N_28635,N_26619,N_27538);
or U28636 (N_28636,N_26475,N_27304);
nand U28637 (N_28637,N_27455,N_27010);
and U28638 (N_28638,N_27010,N_27315);
and U28639 (N_28639,N_26450,N_26492);
or U28640 (N_28640,N_27087,N_26450);
and U28641 (N_28641,N_27005,N_26978);
nor U28642 (N_28642,N_27088,N_27322);
and U28643 (N_28643,N_26818,N_27136);
nand U28644 (N_28644,N_26856,N_26968);
nand U28645 (N_28645,N_26429,N_27590);
nand U28646 (N_28646,N_27208,N_26920);
nand U28647 (N_28647,N_27116,N_27259);
xor U28648 (N_28648,N_27438,N_27416);
nand U28649 (N_28649,N_27455,N_26750);
nor U28650 (N_28650,N_27549,N_26750);
or U28651 (N_28651,N_26818,N_26694);
and U28652 (N_28652,N_26744,N_26967);
and U28653 (N_28653,N_27271,N_26833);
nor U28654 (N_28654,N_27179,N_27071);
and U28655 (N_28655,N_27597,N_27421);
or U28656 (N_28656,N_26880,N_27460);
nand U28657 (N_28657,N_27031,N_26596);
nand U28658 (N_28658,N_27598,N_26730);
and U28659 (N_28659,N_26592,N_26703);
nand U28660 (N_28660,N_26758,N_27223);
xnor U28661 (N_28661,N_27314,N_27029);
nand U28662 (N_28662,N_27051,N_26987);
nor U28663 (N_28663,N_26896,N_26478);
nor U28664 (N_28664,N_26431,N_27541);
and U28665 (N_28665,N_26996,N_27063);
nor U28666 (N_28666,N_26630,N_26938);
nand U28667 (N_28667,N_26835,N_26561);
nor U28668 (N_28668,N_26777,N_27511);
or U28669 (N_28669,N_26624,N_26522);
nor U28670 (N_28670,N_27080,N_27488);
xor U28671 (N_28671,N_27052,N_27185);
xor U28672 (N_28672,N_27040,N_26855);
xor U28673 (N_28673,N_26728,N_26892);
nand U28674 (N_28674,N_27040,N_26994);
nor U28675 (N_28675,N_26672,N_27330);
xor U28676 (N_28676,N_27024,N_26965);
nor U28677 (N_28677,N_27152,N_27035);
nor U28678 (N_28678,N_26901,N_27566);
and U28679 (N_28679,N_26603,N_26639);
nand U28680 (N_28680,N_26879,N_26887);
nand U28681 (N_28681,N_26993,N_27252);
xor U28682 (N_28682,N_26824,N_26400);
nor U28683 (N_28683,N_26776,N_26940);
or U28684 (N_28684,N_26887,N_27439);
xnor U28685 (N_28685,N_27140,N_27380);
or U28686 (N_28686,N_26880,N_27378);
nand U28687 (N_28687,N_26598,N_27344);
nor U28688 (N_28688,N_26442,N_27084);
nor U28689 (N_28689,N_27121,N_26518);
xor U28690 (N_28690,N_26458,N_27031);
or U28691 (N_28691,N_26588,N_26787);
and U28692 (N_28692,N_27239,N_27486);
and U28693 (N_28693,N_26701,N_27163);
nand U28694 (N_28694,N_26488,N_27304);
or U28695 (N_28695,N_26409,N_27328);
and U28696 (N_28696,N_27544,N_27498);
and U28697 (N_28697,N_27560,N_26723);
nor U28698 (N_28698,N_27156,N_27580);
nor U28699 (N_28699,N_27572,N_26543);
nor U28700 (N_28700,N_27030,N_26577);
or U28701 (N_28701,N_26733,N_27444);
and U28702 (N_28702,N_27337,N_27011);
nand U28703 (N_28703,N_27142,N_27299);
and U28704 (N_28704,N_27562,N_27524);
nand U28705 (N_28705,N_26824,N_27120);
xnor U28706 (N_28706,N_26565,N_27204);
and U28707 (N_28707,N_27335,N_27542);
and U28708 (N_28708,N_26947,N_26801);
xnor U28709 (N_28709,N_27575,N_27520);
xor U28710 (N_28710,N_26542,N_27091);
and U28711 (N_28711,N_27514,N_27111);
xnor U28712 (N_28712,N_27505,N_26951);
nand U28713 (N_28713,N_26946,N_26942);
nor U28714 (N_28714,N_27329,N_26426);
nand U28715 (N_28715,N_26457,N_26487);
nor U28716 (N_28716,N_26955,N_26603);
and U28717 (N_28717,N_27384,N_27098);
nor U28718 (N_28718,N_27337,N_26963);
or U28719 (N_28719,N_27251,N_27045);
xor U28720 (N_28720,N_27447,N_26448);
and U28721 (N_28721,N_27082,N_27004);
nand U28722 (N_28722,N_26583,N_26941);
nand U28723 (N_28723,N_26723,N_26975);
xor U28724 (N_28724,N_27368,N_27555);
and U28725 (N_28725,N_27203,N_27592);
nor U28726 (N_28726,N_26817,N_27325);
and U28727 (N_28727,N_26617,N_26753);
xor U28728 (N_28728,N_27196,N_27041);
nand U28729 (N_28729,N_27201,N_27020);
and U28730 (N_28730,N_26630,N_26494);
or U28731 (N_28731,N_27577,N_27343);
nand U28732 (N_28732,N_26904,N_27085);
xor U28733 (N_28733,N_26575,N_26576);
and U28734 (N_28734,N_27202,N_27136);
nor U28735 (N_28735,N_26463,N_26444);
nand U28736 (N_28736,N_26957,N_27287);
and U28737 (N_28737,N_27106,N_27543);
and U28738 (N_28738,N_27486,N_27475);
nand U28739 (N_28739,N_26970,N_27007);
nand U28740 (N_28740,N_26833,N_27073);
nand U28741 (N_28741,N_27222,N_27589);
and U28742 (N_28742,N_27553,N_26974);
and U28743 (N_28743,N_27354,N_26788);
or U28744 (N_28744,N_27416,N_27258);
xnor U28745 (N_28745,N_26813,N_26624);
or U28746 (N_28746,N_26424,N_27162);
nor U28747 (N_28747,N_26809,N_26426);
nor U28748 (N_28748,N_27375,N_27511);
nand U28749 (N_28749,N_27284,N_26807);
nand U28750 (N_28750,N_26772,N_26763);
nor U28751 (N_28751,N_26891,N_26678);
xor U28752 (N_28752,N_26674,N_26823);
or U28753 (N_28753,N_27039,N_27098);
and U28754 (N_28754,N_26675,N_26507);
or U28755 (N_28755,N_27057,N_27368);
or U28756 (N_28756,N_26743,N_27447);
or U28757 (N_28757,N_26961,N_26939);
and U28758 (N_28758,N_27206,N_27304);
or U28759 (N_28759,N_27170,N_26682);
nor U28760 (N_28760,N_26752,N_26450);
or U28761 (N_28761,N_27548,N_27107);
nor U28762 (N_28762,N_27571,N_26677);
xor U28763 (N_28763,N_27593,N_26806);
or U28764 (N_28764,N_27244,N_27138);
or U28765 (N_28765,N_26884,N_27483);
xor U28766 (N_28766,N_27337,N_27080);
or U28767 (N_28767,N_27139,N_27414);
nor U28768 (N_28768,N_26682,N_26514);
nand U28769 (N_28769,N_26519,N_27361);
and U28770 (N_28770,N_27437,N_26953);
nand U28771 (N_28771,N_26762,N_26718);
or U28772 (N_28772,N_27558,N_27085);
or U28773 (N_28773,N_26707,N_27019);
xor U28774 (N_28774,N_26522,N_26658);
xor U28775 (N_28775,N_26521,N_26436);
and U28776 (N_28776,N_27071,N_26444);
nand U28777 (N_28777,N_26584,N_26430);
nor U28778 (N_28778,N_26654,N_26957);
nand U28779 (N_28779,N_27209,N_26458);
and U28780 (N_28780,N_27348,N_27129);
nand U28781 (N_28781,N_26815,N_27542);
and U28782 (N_28782,N_26763,N_26410);
nand U28783 (N_28783,N_27332,N_27322);
or U28784 (N_28784,N_26652,N_27293);
and U28785 (N_28785,N_26505,N_26744);
nor U28786 (N_28786,N_26804,N_26723);
or U28787 (N_28787,N_26517,N_27577);
xor U28788 (N_28788,N_26747,N_26463);
xnor U28789 (N_28789,N_27420,N_27074);
or U28790 (N_28790,N_26626,N_26599);
nor U28791 (N_28791,N_26941,N_27591);
nand U28792 (N_28792,N_27396,N_27356);
or U28793 (N_28793,N_26949,N_27241);
nor U28794 (N_28794,N_26526,N_27392);
nand U28795 (N_28795,N_27414,N_26463);
nor U28796 (N_28796,N_27050,N_27015);
nand U28797 (N_28797,N_27112,N_26447);
or U28798 (N_28798,N_26572,N_26897);
xnor U28799 (N_28799,N_27118,N_26592);
and U28800 (N_28800,N_28251,N_27616);
xor U28801 (N_28801,N_27658,N_27716);
xor U28802 (N_28802,N_27931,N_28486);
or U28803 (N_28803,N_27882,N_27902);
xor U28804 (N_28804,N_28795,N_28367);
nor U28805 (N_28805,N_28422,N_27768);
xor U28806 (N_28806,N_27707,N_28062);
or U28807 (N_28807,N_28199,N_28359);
nand U28808 (N_28808,N_27974,N_27936);
nand U28809 (N_28809,N_28615,N_28789);
nor U28810 (N_28810,N_27606,N_28077);
or U28811 (N_28811,N_28449,N_28556);
and U28812 (N_28812,N_27761,N_27911);
xor U28813 (N_28813,N_27816,N_28351);
nand U28814 (N_28814,N_28553,N_27825);
xor U28815 (N_28815,N_27631,N_28190);
nor U28816 (N_28816,N_28492,N_28480);
and U28817 (N_28817,N_28316,N_28638);
nand U28818 (N_28818,N_28013,N_28511);
nor U28819 (N_28819,N_28014,N_28308);
and U28820 (N_28820,N_28252,N_27954);
xor U28821 (N_28821,N_28424,N_28103);
xnor U28822 (N_28822,N_28576,N_28734);
nor U28823 (N_28823,N_27907,N_28792);
or U28824 (N_28824,N_28610,N_28702);
nand U28825 (N_28825,N_28713,N_28546);
and U28826 (N_28826,N_27939,N_28330);
or U28827 (N_28827,N_28237,N_28264);
nand U28828 (N_28828,N_28698,N_27655);
xor U28829 (N_28829,N_28504,N_27983);
nand U28830 (N_28830,N_28398,N_27672);
or U28831 (N_28831,N_28570,N_27851);
nor U28832 (N_28832,N_27776,N_28481);
or U28833 (N_28833,N_28025,N_27806);
or U28834 (N_28834,N_28463,N_27702);
nor U28835 (N_28835,N_28297,N_28289);
and U28836 (N_28836,N_27796,N_28609);
nand U28837 (N_28837,N_28461,N_27856);
xor U28838 (N_28838,N_27626,N_27839);
and U28839 (N_28839,N_27727,N_28516);
or U28840 (N_28840,N_28366,N_28457);
nor U28841 (N_28841,N_28260,N_28709);
nor U28842 (N_28842,N_28361,N_28784);
and U28843 (N_28843,N_28519,N_28197);
or U28844 (N_28844,N_28592,N_28417);
nand U28845 (N_28845,N_27909,N_28079);
nor U28846 (N_28846,N_28106,N_28643);
xor U28847 (N_28847,N_27649,N_28121);
and U28848 (N_28848,N_28139,N_28224);
or U28849 (N_28849,N_28035,N_28547);
nand U28850 (N_28850,N_27892,N_28049);
and U28851 (N_28851,N_27987,N_27782);
or U28852 (N_28852,N_28098,N_28444);
nand U28853 (N_28853,N_28266,N_28329);
nor U28854 (N_28854,N_28600,N_28323);
xor U28855 (N_28855,N_28740,N_28384);
nor U28856 (N_28856,N_27959,N_28313);
or U28857 (N_28857,N_27832,N_27819);
nand U28858 (N_28858,N_27746,N_28798);
nand U28859 (N_28859,N_28350,N_28168);
xnor U28860 (N_28860,N_28467,N_28605);
or U28861 (N_28861,N_28766,N_28785);
nand U28862 (N_28862,N_28722,N_28127);
and U28863 (N_28863,N_28217,N_27656);
nor U28864 (N_28864,N_28451,N_27890);
nor U28865 (N_28865,N_28627,N_28128);
xnor U28866 (N_28866,N_28231,N_28660);
or U28867 (N_28867,N_28269,N_28063);
or U28868 (N_28868,N_28387,N_28626);
nor U28869 (N_28869,N_27664,N_28603);
or U28870 (N_28870,N_27717,N_28471);
or U28871 (N_28871,N_28774,N_28012);
and U28872 (N_28872,N_27641,N_28580);
nor U28873 (N_28873,N_27928,N_27878);
or U28874 (N_28874,N_27753,N_27917);
nor U28875 (N_28875,N_27901,N_28637);
nor U28876 (N_28876,N_28651,N_28542);
or U28877 (N_28877,N_27773,N_27805);
and U28878 (N_28878,N_28497,N_27934);
xnor U28879 (N_28879,N_28086,N_27704);
nand U28880 (N_28880,N_28137,N_27813);
xnor U28881 (N_28881,N_28443,N_28229);
xor U28882 (N_28882,N_28144,N_27925);
nor U28883 (N_28883,N_28697,N_27946);
xnor U28884 (N_28884,N_28657,N_27814);
and U28885 (N_28885,N_28665,N_27653);
xor U28886 (N_28886,N_28477,N_27845);
or U28887 (N_28887,N_28663,N_28623);
nor U28888 (N_28888,N_27705,N_28548);
xor U28889 (N_28889,N_27718,N_28036);
or U28890 (N_28890,N_28042,N_28183);
and U28891 (N_28891,N_28310,N_27644);
nor U28892 (N_28892,N_28270,N_28619);
nor U28893 (N_28893,N_27879,N_27975);
nor U28894 (N_28894,N_28379,N_28303);
nand U28895 (N_28895,N_27740,N_28239);
nor U28896 (N_28896,N_27899,N_27998);
nor U28897 (N_28897,N_28648,N_27972);
nand U28898 (N_28898,N_28423,N_27894);
nor U28899 (N_28899,N_28472,N_27857);
nand U28900 (N_28900,N_28671,N_28093);
or U28901 (N_28901,N_27682,N_28717);
and U28902 (N_28902,N_28724,N_28732);
nand U28903 (N_28903,N_28053,N_28514);
or U28904 (N_28904,N_28061,N_28584);
or U28905 (N_28905,N_28120,N_28321);
and U28906 (N_28906,N_27984,N_27777);
and U28907 (N_28907,N_28498,N_28325);
nand U28908 (N_28908,N_27745,N_27797);
nor U28909 (N_28909,N_28765,N_28757);
nand U28910 (N_28910,N_28135,N_27950);
xnor U28911 (N_28911,N_28097,N_27897);
nand U28912 (N_28912,N_28733,N_28527);
nor U28913 (N_28913,N_28221,N_28406);
xor U28914 (N_28914,N_28282,N_28394);
or U28915 (N_28915,N_27698,N_28117);
nor U28916 (N_28916,N_27802,N_27652);
nand U28917 (N_28917,N_28376,N_27895);
and U28918 (N_28918,N_28416,N_27600);
or U28919 (N_28919,N_27772,N_28725);
xor U28920 (N_28920,N_28711,N_28189);
nor U28921 (N_28921,N_27996,N_27948);
xor U28922 (N_28922,N_28009,N_28307);
or U28923 (N_28923,N_28150,N_28469);
xnor U28924 (N_28924,N_27980,N_27725);
xnor U28925 (N_28925,N_28390,N_28503);
nand U28926 (N_28926,N_28344,N_28293);
nand U28927 (N_28927,N_27968,N_28572);
nand U28928 (N_28928,N_27662,N_28425);
and U28929 (N_28929,N_28004,N_28292);
or U28930 (N_28930,N_28099,N_28726);
or U28931 (N_28931,N_28640,N_28142);
xnor U28932 (N_28932,N_28105,N_27699);
or U28933 (N_28933,N_28427,N_28368);
xnor U28934 (N_28934,N_28537,N_28218);
nor U28935 (N_28935,N_28540,N_27783);
nand U28936 (N_28936,N_28595,N_28616);
nand U28937 (N_28937,N_28696,N_28565);
nand U28938 (N_28938,N_28085,N_27951);
and U28939 (N_28939,N_28024,N_28283);
or U28940 (N_28940,N_28385,N_28747);
xor U28941 (N_28941,N_28440,N_28203);
xor U28942 (N_28942,N_28331,N_27860);
or U28943 (N_28943,N_28601,N_27926);
or U28944 (N_28944,N_28228,N_28631);
or U28945 (N_28945,N_28030,N_28618);
nor U28946 (N_28946,N_27774,N_28046);
and U28947 (N_28947,N_28000,N_27763);
or U28948 (N_28948,N_28092,N_28608);
xnor U28949 (N_28949,N_27927,N_27713);
and U28950 (N_28950,N_27651,N_27612);
or U28951 (N_28951,N_28163,N_27875);
xnor U28952 (N_28952,N_28191,N_28559);
or U28953 (N_28953,N_28058,N_27867);
and U28954 (N_28954,N_28372,N_28324);
or U28955 (N_28955,N_28112,N_27670);
nand U28956 (N_28956,N_27896,N_27888);
and U28957 (N_28957,N_28666,N_28412);
nor U28958 (N_28958,N_28573,N_28769);
nand U28959 (N_28959,N_27690,N_28018);
and U28960 (N_28960,N_28304,N_28352);
or U28961 (N_28961,N_28484,N_27685);
and U28962 (N_28962,N_27843,N_28295);
and U28963 (N_28963,N_27720,N_27712);
and U28964 (N_28964,N_27838,N_28005);
or U28965 (N_28965,N_27971,N_28544);
and U28966 (N_28966,N_28633,N_28291);
xnor U28967 (N_28967,N_28045,N_28781);
nor U28968 (N_28968,N_28154,N_27676);
or U28969 (N_28969,N_27886,N_27735);
xnor U28970 (N_28970,N_28082,N_28249);
or U28971 (N_28971,N_28288,N_27919);
nand U28972 (N_28972,N_28347,N_28256);
nor U28973 (N_28973,N_28760,N_28536);
and U28974 (N_28974,N_28534,N_28392);
and U28975 (N_28975,N_27637,N_28153);
nand U28976 (N_28976,N_27696,N_27826);
nand U28977 (N_28977,N_27615,N_28299);
nor U28978 (N_28978,N_28431,N_27823);
xor U28979 (N_28979,N_28555,N_27906);
nand U28980 (N_28980,N_28031,N_28284);
and U28981 (N_28981,N_28782,N_28509);
nor U28982 (N_28982,N_28539,N_28653);
xor U28983 (N_28983,N_28654,N_28635);
nand U28984 (N_28984,N_28743,N_27688);
nand U28985 (N_28985,N_28162,N_27608);
nand U28986 (N_28986,N_27765,N_27749);
nor U28987 (N_28987,N_28369,N_28131);
or U28988 (N_28988,N_28586,N_28797);
nand U28989 (N_28989,N_28083,N_27864);
or U28990 (N_28990,N_28628,N_28446);
or U28991 (N_28991,N_28320,N_28622);
nor U28992 (N_28992,N_27885,N_28250);
and U28993 (N_28993,N_28235,N_27962);
xor U28994 (N_28994,N_27957,N_27908);
nand U28995 (N_28995,N_27799,N_27821);
and U28996 (N_28996,N_28756,N_28023);
nor U28997 (N_28997,N_28317,N_27961);
xor U28998 (N_28998,N_28793,N_27918);
nor U28999 (N_28999,N_27611,N_27966);
nand U29000 (N_29000,N_28271,N_27710);
or U29001 (N_29001,N_28614,N_28181);
xnor U29002 (N_29002,N_27840,N_28575);
or U29003 (N_29003,N_27638,N_28505);
or U29004 (N_29004,N_28065,N_28302);
or U29005 (N_29005,N_27829,N_27764);
xnor U29006 (N_29006,N_28286,N_27937);
nor U29007 (N_29007,N_28479,N_27793);
nand U29008 (N_29008,N_28521,N_28647);
nor U29009 (N_29009,N_27981,N_27730);
xor U29010 (N_29010,N_27833,N_27876);
and U29011 (N_29011,N_27863,N_28335);
and U29012 (N_29012,N_27687,N_27929);
xnor U29013 (N_29013,N_27633,N_27800);
xnor U29014 (N_29014,N_28248,N_28763);
nor U29015 (N_29015,N_28211,N_28436);
or U29016 (N_29016,N_27995,N_28564);
nor U29017 (N_29017,N_28043,N_28612);
nand U29018 (N_29018,N_28124,N_28413);
and U29019 (N_29019,N_28166,N_28669);
or U29020 (N_29020,N_28448,N_28273);
nor U29021 (N_29021,N_27965,N_28102);
nor U29022 (N_29022,N_28363,N_28116);
or U29023 (N_29023,N_28475,N_27989);
nand U29024 (N_29024,N_28290,N_28185);
nor U29025 (N_29025,N_28175,N_28593);
nand U29026 (N_29026,N_28585,N_27920);
nand U29027 (N_29027,N_28187,N_27824);
or U29028 (N_29028,N_28489,N_27837);
nor U29029 (N_29029,N_27732,N_28141);
or U29030 (N_29030,N_28332,N_28501);
and U29031 (N_29031,N_28770,N_28474);
and U29032 (N_29032,N_28710,N_28753);
and U29033 (N_29033,N_28507,N_27643);
xnor U29034 (N_29034,N_28220,N_28315);
nand U29035 (N_29035,N_27757,N_27605);
nand U29036 (N_29036,N_28305,N_28579);
xor U29037 (N_29037,N_27775,N_28028);
nand U29038 (N_29038,N_28574,N_28500);
or U29039 (N_29039,N_28581,N_27744);
nor U29040 (N_29040,N_28535,N_28714);
or U29041 (N_29041,N_28690,N_28054);
nor U29042 (N_29042,N_28230,N_27870);
and U29043 (N_29043,N_27990,N_28021);
and U29044 (N_29044,N_27728,N_27669);
nand U29045 (N_29045,N_28037,N_28044);
xnor U29046 (N_29046,N_27741,N_28198);
nand U29047 (N_29047,N_28680,N_28122);
nand U29048 (N_29048,N_27750,N_28727);
nor U29049 (N_29049,N_28115,N_28208);
nand U29050 (N_29050,N_28263,N_28589);
nor U29051 (N_29051,N_28681,N_28353);
nand U29052 (N_29052,N_28206,N_27645);
or U29053 (N_29053,N_27809,N_27779);
nand U29054 (N_29054,N_27841,N_28438);
or U29055 (N_29055,N_28613,N_27747);
and U29056 (N_29056,N_28672,N_28225);
nand U29057 (N_29057,N_27635,N_27969);
or U29058 (N_29058,N_28050,N_28577);
xor U29059 (N_29059,N_27778,N_27963);
and U29060 (N_29060,N_28241,N_27780);
nand U29061 (N_29061,N_27988,N_28401);
nor U29062 (N_29062,N_27803,N_27976);
and U29063 (N_29063,N_27827,N_28405);
nor U29064 (N_29064,N_27915,N_27748);
and U29065 (N_29065,N_27881,N_28383);
or U29066 (N_29066,N_27810,N_28371);
nand U29067 (N_29067,N_28215,N_28739);
xor U29068 (N_29068,N_27785,N_27828);
nor U29069 (N_29069,N_28568,N_28728);
xor U29070 (N_29070,N_28502,N_28532);
nor U29071 (N_29071,N_28567,N_28531);
or U29072 (N_29072,N_28089,N_28704);
nand U29073 (N_29073,N_27850,N_28136);
xnor U29074 (N_29074,N_28196,N_27891);
nor U29075 (N_29075,N_28742,N_27629);
or U29076 (N_29076,N_27620,N_28255);
nor U29077 (N_29077,N_28238,N_27684);
nand U29078 (N_29078,N_28010,N_27752);
and U29079 (N_29079,N_28402,N_27887);
nand U29080 (N_29080,N_28530,N_27999);
nand U29081 (N_29081,N_28020,N_27743);
and U29082 (N_29082,N_28557,N_28148);
nor U29083 (N_29083,N_27848,N_27627);
nor U29084 (N_29084,N_28693,N_28634);
xor U29085 (N_29085,N_28694,N_27859);
nand U29086 (N_29086,N_28267,N_28219);
nor U29087 (N_29087,N_28339,N_28583);
or U29088 (N_29088,N_28072,N_28645);
and U29089 (N_29089,N_28470,N_28234);
xor U29090 (N_29090,N_27835,N_28257);
nor U29091 (N_29091,N_28718,N_28389);
xor U29092 (N_29092,N_27640,N_28377);
nor U29093 (N_29093,N_27898,N_28312);
nor U29094 (N_29094,N_28246,N_28378);
nor U29095 (N_29095,N_28151,N_28426);
xnor U29096 (N_29096,N_27683,N_27880);
nor U29097 (N_29097,N_28226,N_28674);
nor U29098 (N_29098,N_28172,N_28060);
and U29099 (N_29099,N_28015,N_28435);
and U29100 (N_29100,N_28716,N_28685);
or U29101 (N_29101,N_28354,N_28107);
nor U29102 (N_29102,N_28253,N_27942);
nand U29103 (N_29103,N_28796,N_28662);
nor U29104 (N_29104,N_28236,N_27923);
and U29105 (N_29105,N_28073,N_28155);
xnor U29106 (N_29106,N_28165,N_28675);
xnor U29107 (N_29107,N_28420,N_28032);
nor U29108 (N_29108,N_27769,N_28214);
xnor U29109 (N_29109,N_28644,N_27952);
nand U29110 (N_29110,N_28129,N_28499);
nor U29111 (N_29111,N_27602,N_28040);
nor U29112 (N_29112,N_27940,N_28356);
nand U29113 (N_29113,N_27729,N_28526);
and U29114 (N_29114,N_27650,N_28132);
or U29115 (N_29115,N_27634,N_28311);
and U29116 (N_29116,N_28160,N_28541);
xnor U29117 (N_29117,N_28750,N_27623);
xor U29118 (N_29118,N_28678,N_27862);
nor U29119 (N_29119,N_27830,N_28057);
or U29120 (N_29120,N_28775,N_28664);
nor U29121 (N_29121,N_28767,N_28466);
xnor U29122 (N_29122,N_28520,N_28545);
nor U29123 (N_29123,N_28207,N_28432);
nor U29124 (N_29124,N_28705,N_27758);
nor U29125 (N_29125,N_27603,N_28624);
nand U29126 (N_29126,N_28562,N_28382);
nand U29127 (N_29127,N_27930,N_28227);
nor U29128 (N_29128,N_28510,N_28611);
and U29129 (N_29129,N_27994,N_28161);
and U29130 (N_29130,N_28178,N_28091);
nor U29131 (N_29131,N_27665,N_27868);
xnor U29132 (N_29132,N_28066,N_28453);
xor U29133 (N_29133,N_28459,N_28393);
or U29134 (N_29134,N_27628,N_28524);
or U29135 (N_29135,N_28773,N_28429);
xnor U29136 (N_29136,N_28549,N_27977);
xor U29137 (N_29137,N_27861,N_28395);
xor U29138 (N_29138,N_28741,N_27834);
and U29139 (N_29139,N_28523,N_28374);
nor U29140 (N_29140,N_28319,N_28689);
or U29141 (N_29141,N_27795,N_28415);
nor U29142 (N_29142,N_28561,N_27893);
or U29143 (N_29143,N_27889,N_28649);
xor U29144 (N_29144,N_27791,N_28222);
nor U29145 (N_29145,N_28617,N_28341);
xnor U29146 (N_29146,N_28167,N_28587);
and U29147 (N_29147,N_27817,N_27706);
nor U29148 (N_29148,N_27808,N_27700);
or U29149 (N_29149,N_28688,N_28118);
xnor U29150 (N_29150,N_28076,N_28650);
nor U29151 (N_29151,N_28513,N_27770);
and U29152 (N_29152,N_28607,N_27723);
xnor U29153 (N_29153,N_28447,N_27953);
nor U29154 (N_29154,N_28414,N_28193);
nand U29155 (N_29155,N_28125,N_28794);
or U29156 (N_29156,N_27788,N_28119);
nand U29157 (N_29157,N_28296,N_28569);
nand U29158 (N_29158,N_28059,N_28488);
or U29159 (N_29159,N_28465,N_28095);
xnor U29160 (N_29160,N_28528,N_28701);
and U29161 (N_29161,N_28075,N_28194);
nor U29162 (N_29162,N_27865,N_28328);
nand U29163 (N_29163,N_28006,N_27836);
nor U29164 (N_29164,N_28008,N_28033);
or U29165 (N_29165,N_27666,N_27905);
xnor U29166 (N_29166,N_27947,N_28034);
or U29167 (N_29167,N_28146,N_28655);
xnor U29168 (N_29168,N_27792,N_28464);
or U29169 (N_29169,N_28179,N_28364);
and U29170 (N_29170,N_28630,N_28719);
nor U29171 (N_29171,N_28074,N_28778);
nor U29172 (N_29172,N_27842,N_28026);
nand U29173 (N_29173,N_28071,N_28776);
and U29174 (N_29174,N_28003,N_27914);
xor U29175 (N_29175,N_28301,N_27755);
and U29176 (N_29176,N_28764,N_27771);
xor U29177 (N_29177,N_27866,N_27703);
and U29178 (N_29178,N_27846,N_28067);
nor U29179 (N_29179,N_28388,N_28130);
xor U29180 (N_29180,N_27601,N_28563);
or U29181 (N_29181,N_28744,N_28606);
nand U29182 (N_29182,N_27804,N_27941);
or U29183 (N_29183,N_28708,N_27820);
nand U29184 (N_29184,N_28380,N_28355);
and U29185 (N_29185,N_28676,N_27609);
nor U29186 (N_29186,N_28596,N_28597);
or U29187 (N_29187,N_27991,N_27680);
nand U29188 (N_29188,N_28731,N_28349);
and U29189 (N_29189,N_28533,N_28108);
and U29190 (N_29190,N_28223,N_28751);
xnor U29191 (N_29191,N_28104,N_28748);
or U29192 (N_29192,N_27610,N_27913);
or U29193 (N_29193,N_28205,N_28204);
and U29194 (N_29194,N_28262,N_27943);
nand U29195 (N_29195,N_27648,N_28761);
or U29196 (N_29196,N_28343,N_27781);
or U29197 (N_29197,N_27877,N_27789);
nor U29198 (N_29198,N_27979,N_28096);
and U29199 (N_29199,N_27709,N_27715);
xnor U29200 (N_29200,N_28336,N_28683);
nand U29201 (N_29201,N_28621,N_28281);
nor U29202 (N_29202,N_28602,N_28670);
nand U29203 (N_29203,N_27967,N_28454);
nor U29204 (N_29204,N_28397,N_28703);
nor U29205 (N_29205,N_27674,N_28712);
and U29206 (N_29206,N_28791,N_28011);
nor U29207 (N_29207,N_28590,N_28538);
xor U29208 (N_29208,N_28242,N_28174);
xor U29209 (N_29209,N_27849,N_27912);
xor U29210 (N_29210,N_28213,N_28787);
and U29211 (N_29211,N_27964,N_28345);
nor U29212 (N_29212,N_28342,N_27617);
nand U29213 (N_29213,N_27986,N_28578);
nand U29214 (N_29214,N_28749,N_28069);
or U29215 (N_29215,N_28551,N_28306);
nor U29216 (N_29216,N_28090,N_27760);
and U29217 (N_29217,N_27997,N_28768);
xnor U29218 (N_29218,N_28314,N_27711);
xnor U29219 (N_29219,N_28491,N_27671);
nor U29220 (N_29220,N_28441,N_28133);
xnor U29221 (N_29221,N_28625,N_27973);
xnor U29222 (N_29222,N_28686,N_27738);
nor U29223 (N_29223,N_28110,N_27956);
or U29224 (N_29224,N_28200,N_27978);
and U29225 (N_29225,N_28051,N_28188);
nand U29226 (N_29226,N_28055,N_28038);
xor U29227 (N_29227,N_28494,N_28659);
or U29228 (N_29228,N_27807,N_28777);
nand U29229 (N_29229,N_28210,N_27724);
or U29230 (N_29230,N_27853,N_28706);
and U29231 (N_29231,N_28362,N_28375);
nor U29232 (N_29232,N_28735,N_27679);
nor U29233 (N_29233,N_27844,N_28430);
and U29234 (N_29234,N_28201,N_28745);
xor U29235 (N_29235,N_27960,N_28285);
xnor U29236 (N_29236,N_27636,N_28652);
nor U29237 (N_29237,N_28442,N_27639);
or U29238 (N_29238,N_27722,N_27767);
or U29239 (N_29239,N_27742,N_28598);
nor U29240 (N_29240,N_28668,N_27625);
nor U29241 (N_29241,N_28632,N_28604);
xnor U29242 (N_29242,N_28493,N_28468);
nand U29243 (N_29243,N_28259,N_27916);
nor U29244 (N_29244,N_28629,N_27714);
nand U29245 (N_29245,N_28278,N_28720);
and U29246 (N_29246,N_28280,N_27654);
xor U29247 (N_29247,N_28022,N_28746);
or U29248 (N_29248,N_28594,N_28048);
and U29249 (N_29249,N_28386,N_27701);
nand U29250 (N_29250,N_28340,N_27921);
nor U29251 (N_29251,N_28410,N_27621);
nor U29252 (N_29252,N_27855,N_28729);
nand U29253 (N_29253,N_28184,N_27619);
and U29254 (N_29254,N_28691,N_28418);
xnor U29255 (N_29255,N_27993,N_27736);
nor U29256 (N_29256,N_28111,N_28396);
xnor U29257 (N_29257,N_28552,N_28177);
or U29258 (N_29258,N_28245,N_28658);
nor U29259 (N_29259,N_28084,N_27647);
xor U29260 (N_29260,N_27910,N_28772);
nor U29261 (N_29261,N_27949,N_28599);
nand U29262 (N_29262,N_27903,N_27733);
nand U29263 (N_29263,N_28529,N_28571);
nand U29264 (N_29264,N_28243,N_28736);
and U29265 (N_29265,N_27992,N_28409);
and U29266 (N_29266,N_28326,N_28232);
nor U29267 (N_29267,N_28109,N_28790);
and U29268 (N_29268,N_28268,N_28554);
xor U29269 (N_29269,N_28164,N_28639);
nand U29270 (N_29270,N_27731,N_28483);
nor U29271 (N_29271,N_28149,N_28138);
or U29272 (N_29272,N_28202,N_27985);
nand U29273 (N_29273,N_28240,N_28287);
nand U29274 (N_29274,N_28695,N_27660);
and U29275 (N_29275,N_28348,N_28279);
nand U29276 (N_29276,N_28176,N_28508);
and U29277 (N_29277,N_27970,N_28300);
nand U29278 (N_29278,N_28407,N_28399);
nor U29279 (N_29279,N_28247,N_28512);
and U29280 (N_29280,N_28322,N_27958);
xnor U29281 (N_29281,N_28460,N_28799);
and U29282 (N_29282,N_27858,N_27604);
nand U29283 (N_29283,N_28017,N_27622);
or U29284 (N_29284,N_28558,N_28007);
or U29285 (N_29285,N_28357,N_27787);
nor U29286 (N_29286,N_28337,N_28327);
and U29287 (N_29287,N_28411,N_28758);
nor U29288 (N_29288,N_28365,N_28358);
nand U29289 (N_29289,N_28275,N_28707);
nand U29290 (N_29290,N_27697,N_28159);
xor U29291 (N_29291,N_27874,N_28759);
or U29292 (N_29292,N_27719,N_27614);
nor U29293 (N_29293,N_28591,N_28381);
nand U29294 (N_29294,N_27759,N_27873);
xnor U29295 (N_29295,N_27693,N_27872);
and U29296 (N_29296,N_28419,N_28433);
and U29297 (N_29297,N_28677,N_28244);
and U29298 (N_29298,N_28039,N_27618);
and U29299 (N_29299,N_27642,N_28455);
nor U29300 (N_29300,N_27694,N_27944);
xnor U29301 (N_29301,N_28274,N_27726);
and U29302 (N_29302,N_27852,N_28094);
xnor U29303 (N_29303,N_27756,N_28346);
nand U29304 (N_29304,N_28550,N_28019);
or U29305 (N_29305,N_27883,N_28518);
nor U29306 (N_29306,N_28487,N_28123);
nor U29307 (N_29307,N_28762,N_28370);
and U29308 (N_29308,N_28452,N_28113);
and U29309 (N_29309,N_28400,N_28730);
nor U29310 (N_29310,N_28458,N_28334);
nor U29311 (N_29311,N_28522,N_28360);
and U29312 (N_29312,N_28667,N_28041);
or U29313 (N_29313,N_28027,N_28180);
nor U29314 (N_29314,N_27798,N_27790);
and U29315 (N_29315,N_27607,N_28087);
and U29316 (N_29316,N_28140,N_28209);
or U29317 (N_29317,N_27721,N_28506);
nand U29318 (N_29318,N_28788,N_27668);
or U29319 (N_29319,N_28403,N_28212);
and U29320 (N_29320,N_27739,N_27737);
nand U29321 (N_29321,N_28421,N_28134);
or U29322 (N_29322,N_27678,N_27801);
nand U29323 (N_29323,N_28786,N_28081);
nand U29324 (N_29324,N_28029,N_28173);
nor U29325 (N_29325,N_28738,N_28642);
nor U29326 (N_29326,N_28318,N_27632);
and U29327 (N_29327,N_27762,N_27854);
nand U29328 (N_29328,N_28233,N_27847);
xor U29329 (N_29329,N_27935,N_28476);
and U29330 (N_29330,N_28182,N_27955);
and U29331 (N_29331,N_28408,N_28156);
xnor U29332 (N_29332,N_27818,N_28525);
or U29333 (N_29333,N_28152,N_28088);
nand U29334 (N_29334,N_28636,N_27754);
nand U29335 (N_29335,N_28170,N_28261);
nand U29336 (N_29336,N_27884,N_27871);
xnor U29337 (N_29337,N_27667,N_28752);
or U29338 (N_29338,N_28068,N_28294);
or U29339 (N_29339,N_28780,N_28439);
xor U29340 (N_29340,N_27624,N_27938);
and U29341 (N_29341,N_28272,N_28437);
or U29342 (N_29342,N_27630,N_28478);
or U29343 (N_29343,N_28656,N_28754);
or U29344 (N_29344,N_28404,N_28473);
nor U29345 (N_29345,N_28517,N_28047);
nor U29346 (N_29346,N_28582,N_28016);
nor U29347 (N_29347,N_28298,N_27812);
and U29348 (N_29348,N_27689,N_27708);
or U29349 (N_29349,N_28641,N_27924);
or U29350 (N_29350,N_28687,N_27686);
or U29351 (N_29351,N_27982,N_27811);
or U29352 (N_29352,N_28495,N_28078);
nand U29353 (N_29353,N_27692,N_27681);
xnor U29354 (N_29354,N_27822,N_28391);
nand U29355 (N_29355,N_28277,N_28682);
nor U29356 (N_29356,N_28482,N_27786);
and U29357 (N_29357,N_27922,N_28646);
xnor U29358 (N_29358,N_28700,N_28783);
nor U29359 (N_29359,N_27734,N_28001);
xnor U29360 (N_29360,N_28496,N_28333);
or U29361 (N_29361,N_27945,N_28715);
and U29362 (N_29362,N_27831,N_28002);
or U29363 (N_29363,N_28195,N_28064);
nand U29364 (N_29364,N_27659,N_28560);
and U29365 (N_29365,N_28157,N_28186);
and U29366 (N_29366,N_28070,N_28100);
xor U29367 (N_29367,N_28737,N_28169);
and U29368 (N_29368,N_28620,N_27661);
and U29369 (N_29369,N_27613,N_28254);
or U29370 (N_29370,N_27691,N_28434);
and U29371 (N_29371,N_28265,N_28588);
nand U29372 (N_29372,N_28080,N_27675);
and U29373 (N_29373,N_28258,N_28145);
or U29374 (N_29374,N_28126,N_28143);
nand U29375 (N_29375,N_27904,N_28276);
xnor U29376 (N_29376,N_27900,N_27751);
and U29377 (N_29377,N_27815,N_28101);
xnor U29378 (N_29378,N_28309,N_28462);
or U29379 (N_29379,N_28779,N_28692);
nor U29380 (N_29380,N_27933,N_28515);
nor U29381 (N_29381,N_27673,N_28428);
xor U29382 (N_29382,N_28566,N_28673);
nand U29383 (N_29383,N_27657,N_27784);
xnor U29384 (N_29384,N_28771,N_28158);
and U29385 (N_29385,N_27932,N_27663);
or U29386 (N_29386,N_28485,N_28490);
xor U29387 (N_29387,N_27646,N_28338);
or U29388 (N_29388,N_28723,N_28543);
xor U29389 (N_29389,N_27794,N_28373);
xnor U29390 (N_29390,N_28450,N_27677);
or U29391 (N_29391,N_28721,N_28147);
nand U29392 (N_29392,N_27869,N_28679);
nand U29393 (N_29393,N_28684,N_28216);
nor U29394 (N_29394,N_28052,N_27695);
nand U29395 (N_29395,N_28192,N_28445);
nand U29396 (N_29396,N_28171,N_28661);
nand U29397 (N_29397,N_28755,N_28699);
xnor U29398 (N_29398,N_28114,N_27766);
and U29399 (N_29399,N_28456,N_28056);
nor U29400 (N_29400,N_27726,N_27718);
nand U29401 (N_29401,N_28327,N_28499);
and U29402 (N_29402,N_28318,N_28038);
nand U29403 (N_29403,N_27852,N_28027);
nor U29404 (N_29404,N_28459,N_28602);
or U29405 (N_29405,N_28400,N_27994);
or U29406 (N_29406,N_28000,N_28621);
xnor U29407 (N_29407,N_27691,N_28066);
xnor U29408 (N_29408,N_28110,N_28421);
nand U29409 (N_29409,N_28334,N_27984);
or U29410 (N_29410,N_28439,N_28315);
and U29411 (N_29411,N_27839,N_28370);
nor U29412 (N_29412,N_28460,N_28697);
and U29413 (N_29413,N_28185,N_28059);
nor U29414 (N_29414,N_28135,N_28482);
and U29415 (N_29415,N_27971,N_28421);
and U29416 (N_29416,N_28566,N_28773);
nand U29417 (N_29417,N_28084,N_27744);
or U29418 (N_29418,N_28003,N_28583);
nand U29419 (N_29419,N_28760,N_27731);
and U29420 (N_29420,N_28182,N_28305);
or U29421 (N_29421,N_28370,N_28167);
or U29422 (N_29422,N_28358,N_28621);
xnor U29423 (N_29423,N_28239,N_27639);
xnor U29424 (N_29424,N_27681,N_28058);
and U29425 (N_29425,N_28423,N_28009);
nand U29426 (N_29426,N_28546,N_27804);
nor U29427 (N_29427,N_28768,N_28270);
nor U29428 (N_29428,N_28078,N_27614);
nand U29429 (N_29429,N_28767,N_27600);
nor U29430 (N_29430,N_27712,N_28228);
nand U29431 (N_29431,N_28400,N_27692);
nand U29432 (N_29432,N_28454,N_28349);
and U29433 (N_29433,N_27628,N_28332);
xnor U29434 (N_29434,N_27994,N_28640);
or U29435 (N_29435,N_28363,N_28287);
and U29436 (N_29436,N_28794,N_28307);
nand U29437 (N_29437,N_27889,N_27773);
nor U29438 (N_29438,N_28303,N_28456);
and U29439 (N_29439,N_28453,N_28624);
xor U29440 (N_29440,N_27904,N_28176);
nand U29441 (N_29441,N_27824,N_28265);
or U29442 (N_29442,N_27675,N_27620);
xor U29443 (N_29443,N_28370,N_27908);
nor U29444 (N_29444,N_27887,N_28620);
xor U29445 (N_29445,N_28751,N_27686);
or U29446 (N_29446,N_27892,N_27958);
xor U29447 (N_29447,N_28779,N_28708);
and U29448 (N_29448,N_28319,N_27873);
or U29449 (N_29449,N_27914,N_28518);
nor U29450 (N_29450,N_27715,N_27971);
or U29451 (N_29451,N_28746,N_28651);
nand U29452 (N_29452,N_28653,N_27856);
nand U29453 (N_29453,N_27763,N_28273);
or U29454 (N_29454,N_28195,N_28735);
nor U29455 (N_29455,N_28225,N_28053);
or U29456 (N_29456,N_28346,N_28483);
nand U29457 (N_29457,N_27804,N_27817);
or U29458 (N_29458,N_28740,N_28708);
nor U29459 (N_29459,N_28356,N_28293);
nor U29460 (N_29460,N_28071,N_27867);
nand U29461 (N_29461,N_27695,N_28367);
nand U29462 (N_29462,N_28211,N_27844);
nor U29463 (N_29463,N_28070,N_28660);
and U29464 (N_29464,N_27859,N_27708);
or U29465 (N_29465,N_28110,N_27900);
and U29466 (N_29466,N_27998,N_28774);
nor U29467 (N_29467,N_28791,N_27744);
nor U29468 (N_29468,N_28508,N_28516);
or U29469 (N_29469,N_28112,N_28050);
nand U29470 (N_29470,N_28360,N_28144);
nor U29471 (N_29471,N_27987,N_27774);
or U29472 (N_29472,N_28062,N_28291);
nor U29473 (N_29473,N_28135,N_27909);
nand U29474 (N_29474,N_27685,N_28442);
nand U29475 (N_29475,N_28606,N_28680);
or U29476 (N_29476,N_28473,N_28133);
and U29477 (N_29477,N_28484,N_28568);
xnor U29478 (N_29478,N_28385,N_27607);
or U29479 (N_29479,N_28726,N_28346);
or U29480 (N_29480,N_28234,N_28795);
nand U29481 (N_29481,N_28364,N_27725);
nor U29482 (N_29482,N_28712,N_27604);
xnor U29483 (N_29483,N_28288,N_28555);
and U29484 (N_29484,N_28113,N_28011);
nand U29485 (N_29485,N_28665,N_27698);
or U29486 (N_29486,N_28518,N_27793);
nand U29487 (N_29487,N_27603,N_28289);
and U29488 (N_29488,N_27915,N_28470);
nand U29489 (N_29489,N_28116,N_28481);
and U29490 (N_29490,N_28370,N_28200);
nor U29491 (N_29491,N_28794,N_28596);
xnor U29492 (N_29492,N_28176,N_27672);
xor U29493 (N_29493,N_28139,N_28205);
and U29494 (N_29494,N_28580,N_28647);
nor U29495 (N_29495,N_27985,N_27646);
and U29496 (N_29496,N_27903,N_27805);
and U29497 (N_29497,N_27600,N_27698);
nand U29498 (N_29498,N_28039,N_27746);
nor U29499 (N_29499,N_27995,N_27789);
or U29500 (N_29500,N_27664,N_27990);
nand U29501 (N_29501,N_27776,N_27809);
nor U29502 (N_29502,N_28784,N_28136);
nand U29503 (N_29503,N_27788,N_27611);
xnor U29504 (N_29504,N_27954,N_27660);
and U29505 (N_29505,N_28203,N_28105);
xor U29506 (N_29506,N_27996,N_28790);
or U29507 (N_29507,N_28173,N_28128);
xnor U29508 (N_29508,N_28666,N_27793);
xnor U29509 (N_29509,N_27793,N_28195);
or U29510 (N_29510,N_28401,N_28431);
and U29511 (N_29511,N_27785,N_28775);
xor U29512 (N_29512,N_27900,N_27734);
xnor U29513 (N_29513,N_27799,N_27926);
xor U29514 (N_29514,N_28301,N_27646);
and U29515 (N_29515,N_28308,N_28222);
xor U29516 (N_29516,N_27817,N_28157);
xnor U29517 (N_29517,N_28662,N_27985);
and U29518 (N_29518,N_28168,N_28279);
and U29519 (N_29519,N_27897,N_28176);
xor U29520 (N_29520,N_27955,N_27622);
nand U29521 (N_29521,N_28682,N_27923);
nand U29522 (N_29522,N_28730,N_27710);
and U29523 (N_29523,N_28378,N_28417);
nand U29524 (N_29524,N_28161,N_28095);
or U29525 (N_29525,N_27940,N_27976);
nand U29526 (N_29526,N_27899,N_27943);
and U29527 (N_29527,N_27715,N_28016);
nor U29528 (N_29528,N_28204,N_28153);
xor U29529 (N_29529,N_28694,N_27813);
and U29530 (N_29530,N_28503,N_28782);
or U29531 (N_29531,N_27977,N_28590);
or U29532 (N_29532,N_28202,N_28565);
and U29533 (N_29533,N_28683,N_28516);
nor U29534 (N_29534,N_28062,N_27929);
xor U29535 (N_29535,N_28420,N_28105);
xnor U29536 (N_29536,N_28089,N_27784);
nand U29537 (N_29537,N_28321,N_28590);
nor U29538 (N_29538,N_28598,N_28126);
xor U29539 (N_29539,N_28677,N_28404);
and U29540 (N_29540,N_27992,N_28468);
nand U29541 (N_29541,N_28725,N_28171);
nor U29542 (N_29542,N_27728,N_28563);
nor U29543 (N_29543,N_28601,N_27788);
and U29544 (N_29544,N_28008,N_28577);
or U29545 (N_29545,N_27930,N_28371);
and U29546 (N_29546,N_28319,N_28001);
nand U29547 (N_29547,N_28546,N_28342);
nand U29548 (N_29548,N_27981,N_27896);
or U29549 (N_29549,N_27876,N_28619);
and U29550 (N_29550,N_27940,N_28301);
or U29551 (N_29551,N_28125,N_27796);
and U29552 (N_29552,N_27683,N_28277);
nand U29553 (N_29553,N_28200,N_27936);
or U29554 (N_29554,N_28518,N_27723);
nor U29555 (N_29555,N_27647,N_28520);
nand U29556 (N_29556,N_28738,N_27878);
or U29557 (N_29557,N_28004,N_28400);
xnor U29558 (N_29558,N_27761,N_28087);
nand U29559 (N_29559,N_28617,N_28464);
and U29560 (N_29560,N_28512,N_28364);
nand U29561 (N_29561,N_28312,N_28158);
and U29562 (N_29562,N_28577,N_27856);
xnor U29563 (N_29563,N_27739,N_27889);
nor U29564 (N_29564,N_28258,N_28674);
nand U29565 (N_29565,N_27610,N_28787);
xnor U29566 (N_29566,N_28575,N_27891);
nand U29567 (N_29567,N_28741,N_28204);
and U29568 (N_29568,N_28329,N_28633);
xor U29569 (N_29569,N_28098,N_28262);
and U29570 (N_29570,N_28133,N_28276);
nand U29571 (N_29571,N_28768,N_28682);
and U29572 (N_29572,N_28476,N_28505);
nand U29573 (N_29573,N_27929,N_28474);
and U29574 (N_29574,N_28596,N_28208);
or U29575 (N_29575,N_28226,N_27724);
nor U29576 (N_29576,N_28139,N_28622);
nor U29577 (N_29577,N_28181,N_28791);
nand U29578 (N_29578,N_27625,N_27954);
nor U29579 (N_29579,N_27912,N_27937);
nand U29580 (N_29580,N_28536,N_28507);
nand U29581 (N_29581,N_28744,N_28713);
xnor U29582 (N_29582,N_28217,N_27662);
or U29583 (N_29583,N_27794,N_28030);
or U29584 (N_29584,N_28524,N_28365);
or U29585 (N_29585,N_28655,N_27986);
nand U29586 (N_29586,N_27814,N_28605);
and U29587 (N_29587,N_27665,N_27802);
nor U29588 (N_29588,N_28132,N_28193);
nand U29589 (N_29589,N_28247,N_28140);
or U29590 (N_29590,N_27629,N_28276);
nor U29591 (N_29591,N_27995,N_28111);
nor U29592 (N_29592,N_28282,N_27948);
nand U29593 (N_29593,N_28502,N_27670);
or U29594 (N_29594,N_28300,N_27860);
and U29595 (N_29595,N_27667,N_28030);
or U29596 (N_29596,N_28714,N_27951);
nor U29597 (N_29597,N_27695,N_27700);
and U29598 (N_29598,N_27893,N_28410);
and U29599 (N_29599,N_27972,N_28501);
nor U29600 (N_29600,N_28606,N_27884);
nor U29601 (N_29601,N_28448,N_27808);
xnor U29602 (N_29602,N_27839,N_27617);
nor U29603 (N_29603,N_27838,N_28199);
and U29604 (N_29604,N_27925,N_28448);
xor U29605 (N_29605,N_28417,N_27828);
nor U29606 (N_29606,N_28248,N_27654);
and U29607 (N_29607,N_28319,N_28764);
or U29608 (N_29608,N_28169,N_27621);
nor U29609 (N_29609,N_28467,N_28096);
xor U29610 (N_29610,N_28508,N_27944);
xnor U29611 (N_29611,N_28339,N_28490);
nor U29612 (N_29612,N_27903,N_28470);
nor U29613 (N_29613,N_28128,N_28617);
or U29614 (N_29614,N_28574,N_28296);
nand U29615 (N_29615,N_28083,N_28414);
or U29616 (N_29616,N_28689,N_27885);
or U29617 (N_29617,N_28286,N_27603);
xnor U29618 (N_29618,N_27860,N_28427);
nand U29619 (N_29619,N_28044,N_28627);
nand U29620 (N_29620,N_28558,N_28349);
or U29621 (N_29621,N_27834,N_27737);
nor U29622 (N_29622,N_28083,N_28019);
and U29623 (N_29623,N_28162,N_27694);
nand U29624 (N_29624,N_28776,N_28577);
nor U29625 (N_29625,N_28021,N_27928);
nor U29626 (N_29626,N_28115,N_27602);
nor U29627 (N_29627,N_28054,N_27768);
xor U29628 (N_29628,N_28724,N_28047);
xnor U29629 (N_29629,N_28130,N_28338);
xor U29630 (N_29630,N_28096,N_28114);
xnor U29631 (N_29631,N_28409,N_28262);
xnor U29632 (N_29632,N_27937,N_28204);
xor U29633 (N_29633,N_28246,N_28567);
and U29634 (N_29634,N_27881,N_27893);
nand U29635 (N_29635,N_28440,N_28763);
and U29636 (N_29636,N_28003,N_27834);
or U29637 (N_29637,N_28463,N_28339);
nor U29638 (N_29638,N_28564,N_28126);
nand U29639 (N_29639,N_28319,N_28307);
xor U29640 (N_29640,N_28192,N_28475);
nand U29641 (N_29641,N_28468,N_28719);
nor U29642 (N_29642,N_27975,N_27829);
and U29643 (N_29643,N_28544,N_27784);
nand U29644 (N_29644,N_28785,N_28695);
and U29645 (N_29645,N_28604,N_27838);
xnor U29646 (N_29646,N_28797,N_28491);
xnor U29647 (N_29647,N_28420,N_28331);
nor U29648 (N_29648,N_28441,N_28099);
nand U29649 (N_29649,N_28717,N_28034);
nor U29650 (N_29650,N_28159,N_27776);
or U29651 (N_29651,N_28407,N_27786);
nand U29652 (N_29652,N_28156,N_28100);
nand U29653 (N_29653,N_28693,N_28102);
nor U29654 (N_29654,N_28726,N_28160);
nor U29655 (N_29655,N_28634,N_28113);
and U29656 (N_29656,N_27969,N_28551);
xor U29657 (N_29657,N_28125,N_28048);
and U29658 (N_29658,N_27768,N_27723);
nand U29659 (N_29659,N_28155,N_28676);
nor U29660 (N_29660,N_28769,N_28175);
nor U29661 (N_29661,N_28356,N_28486);
nor U29662 (N_29662,N_28312,N_28186);
nor U29663 (N_29663,N_28034,N_28771);
nor U29664 (N_29664,N_28550,N_27903);
nand U29665 (N_29665,N_28715,N_27721);
nand U29666 (N_29666,N_27966,N_28429);
nand U29667 (N_29667,N_27998,N_28608);
nor U29668 (N_29668,N_28378,N_27963);
or U29669 (N_29669,N_28129,N_27970);
nor U29670 (N_29670,N_28707,N_28622);
and U29671 (N_29671,N_28738,N_28743);
and U29672 (N_29672,N_27673,N_27686);
xor U29673 (N_29673,N_27865,N_28321);
nor U29674 (N_29674,N_28287,N_28096);
xor U29675 (N_29675,N_28118,N_27760);
or U29676 (N_29676,N_28255,N_27948);
nor U29677 (N_29677,N_27724,N_28388);
and U29678 (N_29678,N_28282,N_28717);
or U29679 (N_29679,N_28570,N_28546);
nand U29680 (N_29680,N_28475,N_28703);
or U29681 (N_29681,N_28658,N_27786);
nand U29682 (N_29682,N_27933,N_27690);
nand U29683 (N_29683,N_28367,N_28146);
nor U29684 (N_29684,N_28648,N_27752);
and U29685 (N_29685,N_28270,N_27771);
nand U29686 (N_29686,N_27962,N_27733);
nand U29687 (N_29687,N_28146,N_28533);
and U29688 (N_29688,N_28430,N_28451);
nand U29689 (N_29689,N_27897,N_28129);
nand U29690 (N_29690,N_28531,N_27606);
nor U29691 (N_29691,N_28161,N_28218);
xnor U29692 (N_29692,N_28671,N_28348);
or U29693 (N_29693,N_28718,N_28385);
xor U29694 (N_29694,N_28296,N_28519);
and U29695 (N_29695,N_28337,N_28740);
or U29696 (N_29696,N_27836,N_28482);
xor U29697 (N_29697,N_28215,N_27862);
and U29698 (N_29698,N_27828,N_27645);
xnor U29699 (N_29699,N_27792,N_28738);
or U29700 (N_29700,N_28596,N_28268);
xnor U29701 (N_29701,N_28383,N_27636);
and U29702 (N_29702,N_28534,N_28518);
nor U29703 (N_29703,N_28603,N_28297);
or U29704 (N_29704,N_27787,N_28558);
nor U29705 (N_29705,N_27813,N_28722);
or U29706 (N_29706,N_28152,N_28629);
nand U29707 (N_29707,N_27946,N_28235);
nand U29708 (N_29708,N_28504,N_28229);
nor U29709 (N_29709,N_28678,N_28380);
xor U29710 (N_29710,N_27949,N_28668);
nand U29711 (N_29711,N_28405,N_27633);
and U29712 (N_29712,N_28706,N_28230);
nor U29713 (N_29713,N_27719,N_28217);
or U29714 (N_29714,N_28787,N_27804);
and U29715 (N_29715,N_28419,N_28765);
or U29716 (N_29716,N_28777,N_28775);
nand U29717 (N_29717,N_28332,N_28428);
and U29718 (N_29718,N_28466,N_27676);
and U29719 (N_29719,N_28127,N_28208);
nand U29720 (N_29720,N_28299,N_27891);
or U29721 (N_29721,N_28669,N_27635);
xnor U29722 (N_29722,N_28681,N_27674);
and U29723 (N_29723,N_28344,N_28657);
nand U29724 (N_29724,N_28686,N_28431);
or U29725 (N_29725,N_28636,N_28469);
nor U29726 (N_29726,N_28455,N_28767);
nor U29727 (N_29727,N_28449,N_28115);
nor U29728 (N_29728,N_27733,N_28335);
or U29729 (N_29729,N_28151,N_28456);
xor U29730 (N_29730,N_28086,N_28167);
nor U29731 (N_29731,N_28313,N_28429);
nor U29732 (N_29732,N_28588,N_27970);
or U29733 (N_29733,N_27776,N_28728);
nor U29734 (N_29734,N_27669,N_28663);
xnor U29735 (N_29735,N_27738,N_27932);
or U29736 (N_29736,N_28388,N_28568);
or U29737 (N_29737,N_28756,N_27700);
nor U29738 (N_29738,N_28107,N_28510);
nor U29739 (N_29739,N_27955,N_28540);
and U29740 (N_29740,N_27868,N_28493);
nor U29741 (N_29741,N_27754,N_28768);
nand U29742 (N_29742,N_27671,N_27956);
nor U29743 (N_29743,N_28798,N_28077);
or U29744 (N_29744,N_27961,N_28475);
and U29745 (N_29745,N_28093,N_28497);
and U29746 (N_29746,N_28622,N_28697);
xnor U29747 (N_29747,N_27829,N_27916);
nand U29748 (N_29748,N_28518,N_27615);
xor U29749 (N_29749,N_28758,N_28398);
and U29750 (N_29750,N_27778,N_28438);
or U29751 (N_29751,N_28665,N_28240);
or U29752 (N_29752,N_28577,N_28292);
nor U29753 (N_29753,N_28732,N_27670);
or U29754 (N_29754,N_27845,N_27921);
nor U29755 (N_29755,N_28295,N_28160);
nor U29756 (N_29756,N_28564,N_28570);
nor U29757 (N_29757,N_28406,N_27727);
xnor U29758 (N_29758,N_28118,N_28712);
xor U29759 (N_29759,N_28164,N_27656);
nor U29760 (N_29760,N_28605,N_27898);
xnor U29761 (N_29761,N_28775,N_28660);
xnor U29762 (N_29762,N_28002,N_28598);
and U29763 (N_29763,N_28562,N_28663);
nor U29764 (N_29764,N_27692,N_28099);
nor U29765 (N_29765,N_28490,N_28404);
nand U29766 (N_29766,N_27902,N_28426);
nand U29767 (N_29767,N_27784,N_28456);
nand U29768 (N_29768,N_28258,N_27658);
nor U29769 (N_29769,N_28166,N_28740);
nand U29770 (N_29770,N_28602,N_27874);
nand U29771 (N_29771,N_28787,N_28233);
xor U29772 (N_29772,N_28197,N_28697);
and U29773 (N_29773,N_28213,N_28027);
or U29774 (N_29774,N_27944,N_28011);
or U29775 (N_29775,N_28204,N_28260);
nand U29776 (N_29776,N_28798,N_28734);
or U29777 (N_29777,N_27876,N_28715);
and U29778 (N_29778,N_28300,N_28019);
xor U29779 (N_29779,N_28611,N_28451);
nor U29780 (N_29780,N_27896,N_28395);
and U29781 (N_29781,N_28090,N_28180);
xnor U29782 (N_29782,N_28710,N_28369);
nand U29783 (N_29783,N_28748,N_28543);
xor U29784 (N_29784,N_28625,N_28432);
nand U29785 (N_29785,N_27978,N_28196);
nand U29786 (N_29786,N_28060,N_27768);
nor U29787 (N_29787,N_28199,N_27670);
and U29788 (N_29788,N_28598,N_28658);
or U29789 (N_29789,N_28613,N_28603);
nand U29790 (N_29790,N_28245,N_27974);
nor U29791 (N_29791,N_28681,N_27626);
nor U29792 (N_29792,N_28497,N_27776);
nand U29793 (N_29793,N_28538,N_27671);
xor U29794 (N_29794,N_28747,N_28270);
xnor U29795 (N_29795,N_28285,N_27860);
or U29796 (N_29796,N_28554,N_28575);
nor U29797 (N_29797,N_28697,N_28519);
nand U29798 (N_29798,N_28233,N_27728);
and U29799 (N_29799,N_27988,N_28708);
xnor U29800 (N_29800,N_28675,N_28164);
or U29801 (N_29801,N_28549,N_27894);
xor U29802 (N_29802,N_27813,N_28619);
nand U29803 (N_29803,N_28457,N_28645);
nand U29804 (N_29804,N_27612,N_28671);
or U29805 (N_29805,N_27944,N_28177);
or U29806 (N_29806,N_27780,N_28438);
or U29807 (N_29807,N_28662,N_27869);
nand U29808 (N_29808,N_27645,N_28393);
and U29809 (N_29809,N_28525,N_27796);
xor U29810 (N_29810,N_28472,N_28195);
nor U29811 (N_29811,N_28758,N_28748);
xor U29812 (N_29812,N_28215,N_28119);
or U29813 (N_29813,N_28200,N_28204);
xnor U29814 (N_29814,N_28321,N_28479);
and U29815 (N_29815,N_28668,N_28630);
or U29816 (N_29816,N_28101,N_28544);
or U29817 (N_29817,N_28730,N_27981);
and U29818 (N_29818,N_28199,N_28219);
and U29819 (N_29819,N_28662,N_28558);
nor U29820 (N_29820,N_27681,N_28070);
xor U29821 (N_29821,N_28526,N_28120);
nor U29822 (N_29822,N_28592,N_27892);
nor U29823 (N_29823,N_28128,N_28461);
and U29824 (N_29824,N_28741,N_27664);
and U29825 (N_29825,N_28213,N_27882);
xor U29826 (N_29826,N_28568,N_28264);
and U29827 (N_29827,N_28132,N_27979);
nand U29828 (N_29828,N_28764,N_28468);
and U29829 (N_29829,N_28556,N_28231);
nor U29830 (N_29830,N_28656,N_28529);
or U29831 (N_29831,N_28575,N_28259);
and U29832 (N_29832,N_27721,N_28422);
and U29833 (N_29833,N_27974,N_27810);
nor U29834 (N_29834,N_28491,N_28645);
and U29835 (N_29835,N_27648,N_27864);
xnor U29836 (N_29836,N_27644,N_28772);
and U29837 (N_29837,N_28183,N_27877);
nand U29838 (N_29838,N_28618,N_27980);
nor U29839 (N_29839,N_28004,N_28032);
nor U29840 (N_29840,N_27785,N_28002);
nor U29841 (N_29841,N_27783,N_27817);
nand U29842 (N_29842,N_28222,N_27661);
or U29843 (N_29843,N_27678,N_27881);
and U29844 (N_29844,N_27855,N_28195);
and U29845 (N_29845,N_28126,N_27630);
and U29846 (N_29846,N_27874,N_28666);
xor U29847 (N_29847,N_27704,N_28088);
xor U29848 (N_29848,N_27724,N_28697);
or U29849 (N_29849,N_28159,N_27669);
and U29850 (N_29850,N_27618,N_28517);
nand U29851 (N_29851,N_28145,N_27692);
nor U29852 (N_29852,N_28536,N_27739);
nand U29853 (N_29853,N_27644,N_28301);
nor U29854 (N_29854,N_28447,N_28493);
nand U29855 (N_29855,N_27946,N_28685);
and U29856 (N_29856,N_27692,N_28123);
and U29857 (N_29857,N_27804,N_28644);
or U29858 (N_29858,N_28238,N_27998);
nand U29859 (N_29859,N_28118,N_28000);
xor U29860 (N_29860,N_27817,N_28025);
nor U29861 (N_29861,N_28676,N_27807);
xnor U29862 (N_29862,N_28748,N_27769);
and U29863 (N_29863,N_27697,N_28470);
or U29864 (N_29864,N_27748,N_28077);
or U29865 (N_29865,N_28749,N_27831);
nand U29866 (N_29866,N_27806,N_28409);
xor U29867 (N_29867,N_28237,N_27936);
nand U29868 (N_29868,N_28407,N_27735);
or U29869 (N_29869,N_28308,N_28413);
nand U29870 (N_29870,N_28533,N_28475);
nand U29871 (N_29871,N_28153,N_27732);
xnor U29872 (N_29872,N_27815,N_28099);
and U29873 (N_29873,N_27894,N_27736);
xnor U29874 (N_29874,N_28401,N_28376);
nor U29875 (N_29875,N_28440,N_27842);
and U29876 (N_29876,N_28423,N_27882);
or U29877 (N_29877,N_28237,N_28054);
or U29878 (N_29878,N_28309,N_27644);
nor U29879 (N_29879,N_28064,N_27667);
or U29880 (N_29880,N_28303,N_27796);
xnor U29881 (N_29881,N_27791,N_28379);
or U29882 (N_29882,N_28170,N_27864);
and U29883 (N_29883,N_28121,N_28617);
and U29884 (N_29884,N_28085,N_27760);
xor U29885 (N_29885,N_27717,N_28171);
xnor U29886 (N_29886,N_27821,N_28502);
or U29887 (N_29887,N_27853,N_28327);
or U29888 (N_29888,N_28123,N_28470);
or U29889 (N_29889,N_28051,N_28116);
xor U29890 (N_29890,N_27999,N_27770);
nor U29891 (N_29891,N_28620,N_28409);
nor U29892 (N_29892,N_27967,N_27812);
nand U29893 (N_29893,N_28098,N_27879);
xnor U29894 (N_29894,N_27669,N_28100);
nor U29895 (N_29895,N_28442,N_28712);
and U29896 (N_29896,N_28517,N_28229);
or U29897 (N_29897,N_27760,N_28596);
nand U29898 (N_29898,N_28420,N_28346);
xor U29899 (N_29899,N_28459,N_28660);
xor U29900 (N_29900,N_28512,N_27938);
and U29901 (N_29901,N_28044,N_28753);
nor U29902 (N_29902,N_27612,N_28068);
nand U29903 (N_29903,N_27852,N_27828);
xnor U29904 (N_29904,N_28158,N_28114);
and U29905 (N_29905,N_27633,N_27873);
nand U29906 (N_29906,N_28204,N_28330);
nand U29907 (N_29907,N_28662,N_28108);
and U29908 (N_29908,N_28110,N_28508);
nand U29909 (N_29909,N_28396,N_27944);
nor U29910 (N_29910,N_27847,N_28452);
xor U29911 (N_29911,N_28606,N_27912);
nand U29912 (N_29912,N_27638,N_28607);
nand U29913 (N_29913,N_28204,N_28593);
and U29914 (N_29914,N_28474,N_28317);
nor U29915 (N_29915,N_28794,N_28259);
nor U29916 (N_29916,N_28156,N_28753);
nand U29917 (N_29917,N_27613,N_28067);
xor U29918 (N_29918,N_27606,N_28775);
or U29919 (N_29919,N_28774,N_28729);
nand U29920 (N_29920,N_28751,N_28798);
nand U29921 (N_29921,N_27876,N_28664);
nand U29922 (N_29922,N_27641,N_28382);
or U29923 (N_29923,N_28529,N_28472);
nand U29924 (N_29924,N_27811,N_28234);
xnor U29925 (N_29925,N_28518,N_28377);
or U29926 (N_29926,N_28129,N_28784);
or U29927 (N_29927,N_28355,N_27993);
nor U29928 (N_29928,N_27710,N_27685);
nor U29929 (N_29929,N_27622,N_28655);
nand U29930 (N_29930,N_27727,N_28736);
or U29931 (N_29931,N_28761,N_27723);
or U29932 (N_29932,N_27713,N_28650);
nand U29933 (N_29933,N_27745,N_27899);
xor U29934 (N_29934,N_27856,N_28374);
and U29935 (N_29935,N_27650,N_27984);
and U29936 (N_29936,N_27925,N_28325);
nor U29937 (N_29937,N_28130,N_27947);
or U29938 (N_29938,N_28303,N_27705);
nor U29939 (N_29939,N_28241,N_28317);
or U29940 (N_29940,N_27928,N_28782);
nand U29941 (N_29941,N_28736,N_27625);
and U29942 (N_29942,N_28600,N_28328);
and U29943 (N_29943,N_28670,N_28767);
nand U29944 (N_29944,N_28760,N_27819);
nand U29945 (N_29945,N_27752,N_28392);
xnor U29946 (N_29946,N_27990,N_27834);
and U29947 (N_29947,N_28130,N_28786);
xnor U29948 (N_29948,N_27760,N_28082);
nor U29949 (N_29949,N_28237,N_28019);
xor U29950 (N_29950,N_28364,N_27966);
or U29951 (N_29951,N_27957,N_28069);
nor U29952 (N_29952,N_28667,N_28682);
and U29953 (N_29953,N_28168,N_28568);
nand U29954 (N_29954,N_28562,N_28284);
nor U29955 (N_29955,N_28275,N_27819);
xnor U29956 (N_29956,N_28387,N_27604);
nand U29957 (N_29957,N_28364,N_28125);
nand U29958 (N_29958,N_28265,N_27806);
xnor U29959 (N_29959,N_27667,N_27771);
xnor U29960 (N_29960,N_27991,N_28122);
or U29961 (N_29961,N_28313,N_27875);
nor U29962 (N_29962,N_27939,N_28561);
nand U29963 (N_29963,N_28102,N_28118);
or U29964 (N_29964,N_28154,N_28070);
or U29965 (N_29965,N_28532,N_27823);
xor U29966 (N_29966,N_28746,N_28048);
nor U29967 (N_29967,N_27903,N_28729);
nor U29968 (N_29968,N_28649,N_27765);
and U29969 (N_29969,N_28419,N_27729);
or U29970 (N_29970,N_28479,N_27791);
and U29971 (N_29971,N_27957,N_27941);
and U29972 (N_29972,N_27642,N_28619);
or U29973 (N_29973,N_28407,N_28460);
nand U29974 (N_29974,N_27752,N_28084);
and U29975 (N_29975,N_28177,N_28095);
and U29976 (N_29976,N_28202,N_28396);
nor U29977 (N_29977,N_28120,N_28206);
nor U29978 (N_29978,N_27771,N_28279);
and U29979 (N_29979,N_28302,N_28640);
and U29980 (N_29980,N_27628,N_28562);
nand U29981 (N_29981,N_27712,N_28695);
and U29982 (N_29982,N_27926,N_27603);
and U29983 (N_29983,N_27983,N_28586);
xor U29984 (N_29984,N_28389,N_28634);
nand U29985 (N_29985,N_28661,N_28561);
or U29986 (N_29986,N_27601,N_28638);
nor U29987 (N_29987,N_28397,N_28008);
and U29988 (N_29988,N_28303,N_27973);
nand U29989 (N_29989,N_27740,N_28713);
or U29990 (N_29990,N_28467,N_28639);
nor U29991 (N_29991,N_28503,N_28707);
xor U29992 (N_29992,N_27682,N_28798);
xor U29993 (N_29993,N_28228,N_27894);
nor U29994 (N_29994,N_28617,N_28729);
and U29995 (N_29995,N_28410,N_27811);
nor U29996 (N_29996,N_27798,N_27831);
xor U29997 (N_29997,N_27957,N_27912);
or U29998 (N_29998,N_28331,N_27783);
or U29999 (N_29999,N_27813,N_28112);
nand UO_0 (O_0,N_29076,N_28810);
nand UO_1 (O_1,N_29821,N_29865);
or UO_2 (O_2,N_28980,N_29189);
or UO_3 (O_3,N_28885,N_29128);
and UO_4 (O_4,N_29462,N_29774);
nand UO_5 (O_5,N_29481,N_29695);
or UO_6 (O_6,N_29374,N_29950);
xnor UO_7 (O_7,N_29122,N_29700);
nand UO_8 (O_8,N_28979,N_29438);
and UO_9 (O_9,N_29726,N_29044);
nor UO_10 (O_10,N_29061,N_29217);
nor UO_11 (O_11,N_29332,N_29977);
or UO_12 (O_12,N_29570,N_29553);
and UO_13 (O_13,N_28946,N_29706);
or UO_14 (O_14,N_29088,N_29798);
nor UO_15 (O_15,N_29324,N_29132);
and UO_16 (O_16,N_28812,N_29072);
or UO_17 (O_17,N_29897,N_29877);
xor UO_18 (O_18,N_29485,N_28884);
nand UO_19 (O_19,N_29247,N_29255);
xor UO_20 (O_20,N_29589,N_28813);
xnor UO_21 (O_21,N_29926,N_29796);
or UO_22 (O_22,N_29475,N_29530);
xnor UO_23 (O_23,N_28840,N_29022);
nand UO_24 (O_24,N_29509,N_28918);
or UO_25 (O_25,N_29141,N_29474);
xnor UO_26 (O_26,N_29371,N_29041);
or UO_27 (O_27,N_28814,N_29351);
or UO_28 (O_28,N_29758,N_29146);
or UO_29 (O_29,N_29498,N_29185);
or UO_30 (O_30,N_29435,N_29571);
and UO_31 (O_31,N_29263,N_29943);
or UO_32 (O_32,N_29080,N_29355);
nor UO_33 (O_33,N_29387,N_29499);
xor UO_34 (O_34,N_29607,N_29478);
or UO_35 (O_35,N_29031,N_29598);
and UO_36 (O_36,N_29736,N_29245);
nor UO_37 (O_37,N_29363,N_29461);
xnor UO_38 (O_38,N_29442,N_28953);
xnor UO_39 (O_39,N_29690,N_29439);
nor UO_40 (O_40,N_28988,N_29963);
xor UO_41 (O_41,N_29527,N_29696);
xnor UO_42 (O_42,N_29623,N_29864);
nand UO_43 (O_43,N_29221,N_29920);
and UO_44 (O_44,N_29555,N_29233);
or UO_45 (O_45,N_29754,N_29738);
nand UO_46 (O_46,N_29939,N_29325);
xnor UO_47 (O_47,N_29347,N_29767);
or UO_48 (O_48,N_29396,N_29647);
or UO_49 (O_49,N_29394,N_28905);
nor UO_50 (O_50,N_29138,N_29525);
or UO_51 (O_51,N_29861,N_29951);
xnor UO_52 (O_52,N_28952,N_29275);
nand UO_53 (O_53,N_29515,N_29884);
xor UO_54 (O_54,N_28955,N_29546);
or UO_55 (O_55,N_29984,N_29538);
xor UO_56 (O_56,N_29424,N_29914);
or UO_57 (O_57,N_29787,N_29673);
nand UO_58 (O_58,N_29399,N_29280);
or UO_59 (O_59,N_29075,N_29104);
nor UO_60 (O_60,N_29228,N_29933);
nand UO_61 (O_61,N_29824,N_29826);
xnor UO_62 (O_62,N_29569,N_29202);
xnor UO_63 (O_63,N_29123,N_29517);
and UO_64 (O_64,N_29505,N_29057);
xor UO_65 (O_65,N_28856,N_28935);
xor UO_66 (O_66,N_29974,N_29602);
or UO_67 (O_67,N_29265,N_29992);
or UO_68 (O_68,N_29340,N_29383);
nor UO_69 (O_69,N_29611,N_29831);
and UO_70 (O_70,N_29887,N_29526);
xor UO_71 (O_71,N_29356,N_29440);
xor UO_72 (O_72,N_29043,N_29973);
nor UO_73 (O_73,N_29628,N_29448);
nand UO_74 (O_74,N_29453,N_29846);
xnor UO_75 (O_75,N_29924,N_29411);
or UO_76 (O_76,N_28809,N_28919);
and UO_77 (O_77,N_29292,N_29875);
or UO_78 (O_78,N_29544,N_29282);
nor UO_79 (O_79,N_29425,N_29686);
nand UO_80 (O_80,N_29085,N_28879);
or UO_81 (O_81,N_29760,N_29307);
nand UO_82 (O_82,N_29070,N_29295);
xor UO_83 (O_83,N_29130,N_29004);
xor UO_84 (O_84,N_29249,N_29718);
nor UO_85 (O_85,N_29005,N_29502);
nor UO_86 (O_86,N_28848,N_29671);
and UO_87 (O_87,N_29523,N_29595);
nand UO_88 (O_88,N_29330,N_29014);
and UO_89 (O_89,N_29580,N_29936);
and UO_90 (O_90,N_29616,N_29894);
nand UO_91 (O_91,N_29501,N_29173);
or UO_92 (O_92,N_28976,N_29834);
xnor UO_93 (O_93,N_29844,N_29311);
or UO_94 (O_94,N_28831,N_29494);
or UO_95 (O_95,N_29968,N_29006);
or UO_96 (O_96,N_29388,N_29635);
and UO_97 (O_97,N_29522,N_29540);
xnor UO_98 (O_98,N_29337,N_29464);
or UO_99 (O_99,N_28862,N_29480);
and UO_100 (O_100,N_29379,N_29037);
and UO_101 (O_101,N_29719,N_28854);
nor UO_102 (O_102,N_29083,N_29048);
nor UO_103 (O_103,N_29631,N_29641);
nor UO_104 (O_104,N_28934,N_29373);
or UO_105 (O_105,N_29214,N_29863);
nand UO_106 (O_106,N_29880,N_29378);
and UO_107 (O_107,N_29640,N_28967);
and UO_108 (O_108,N_29513,N_29932);
nand UO_109 (O_109,N_29304,N_29678);
and UO_110 (O_110,N_28911,N_29841);
xor UO_111 (O_111,N_29294,N_29303);
and UO_112 (O_112,N_29215,N_29627);
nand UO_113 (O_113,N_29133,N_29857);
nor UO_114 (O_114,N_29717,N_29113);
nand UO_115 (O_115,N_29843,N_29915);
and UO_116 (O_116,N_29056,N_29261);
nand UO_117 (O_117,N_29913,N_29534);
nand UO_118 (O_118,N_28957,N_29446);
nand UO_119 (O_119,N_29300,N_29029);
nand UO_120 (O_120,N_29354,N_29590);
or UO_121 (O_121,N_28997,N_29588);
nand UO_122 (O_122,N_29472,N_29360);
nand UO_123 (O_123,N_29539,N_29893);
nor UO_124 (O_124,N_29966,N_29507);
nor UO_125 (O_125,N_29147,N_29630);
nand UO_126 (O_126,N_29591,N_29422);
nand UO_127 (O_127,N_29218,N_28815);
nor UO_128 (O_128,N_29953,N_29621);
or UO_129 (O_129,N_29151,N_29314);
nor UO_130 (O_130,N_28883,N_28846);
or UO_131 (O_131,N_28949,N_29871);
and UO_132 (O_132,N_29238,N_29322);
or UO_133 (O_133,N_29947,N_29782);
xor UO_134 (O_134,N_29962,N_29222);
nand UO_135 (O_135,N_28972,N_29203);
or UO_136 (O_136,N_29922,N_29904);
nand UO_137 (O_137,N_29883,N_29389);
nand UO_138 (O_138,N_29262,N_29847);
and UO_139 (O_139,N_29119,N_29366);
nor UO_140 (O_140,N_29154,N_29045);
xnor UO_141 (O_141,N_29308,N_28886);
nand UO_142 (O_142,N_28930,N_29870);
xor UO_143 (O_143,N_29035,N_29510);
xor UO_144 (O_144,N_28995,N_29753);
and UO_145 (O_145,N_29748,N_29701);
xor UO_146 (O_146,N_29476,N_28857);
nor UO_147 (O_147,N_28956,N_29949);
nor UO_148 (O_148,N_29972,N_29775);
or UO_149 (O_149,N_29855,N_29692);
nor UO_150 (O_150,N_28961,N_29998);
or UO_151 (O_151,N_29693,N_28820);
or UO_152 (O_152,N_28863,N_29771);
nor UO_153 (O_153,N_29646,N_28873);
xor UO_154 (O_154,N_29423,N_29090);
xor UO_155 (O_155,N_29801,N_29063);
or UO_156 (O_156,N_29162,N_29983);
nor UO_157 (O_157,N_29651,N_29670);
nor UO_158 (O_158,N_29250,N_28960);
nand UO_159 (O_159,N_29109,N_29482);
and UO_160 (O_160,N_29626,N_29930);
or UO_161 (O_161,N_29179,N_28917);
nor UO_162 (O_162,N_29667,N_29650);
nand UO_163 (O_163,N_29575,N_29227);
and UO_164 (O_164,N_29634,N_29059);
xor UO_165 (O_165,N_29199,N_29741);
or UO_166 (O_166,N_29068,N_29652);
xnor UO_167 (O_167,N_28920,N_29251);
nor UO_168 (O_168,N_29060,N_29783);
xnor UO_169 (O_169,N_29988,N_29769);
nand UO_170 (O_170,N_29687,N_29891);
nand UO_171 (O_171,N_29207,N_28944);
nand UO_172 (O_172,N_29323,N_29999);
or UO_173 (O_173,N_28966,N_29126);
xnor UO_174 (O_174,N_29042,N_29731);
nor UO_175 (O_175,N_29654,N_29994);
xor UO_176 (O_176,N_29709,N_29025);
nor UO_177 (O_177,N_28948,N_29003);
and UO_178 (O_178,N_29664,N_29566);
nand UO_179 (O_179,N_29483,N_29929);
nand UO_180 (O_180,N_29622,N_28978);
nor UO_181 (O_181,N_29459,N_29256);
nand UO_182 (O_182,N_29541,N_29506);
xor UO_183 (O_183,N_29702,N_29487);
nor UO_184 (O_184,N_29365,N_28903);
xor UO_185 (O_185,N_28924,N_29368);
nand UO_186 (O_186,N_28900,N_29028);
nor UO_187 (O_187,N_29143,N_29633);
or UO_188 (O_188,N_29528,N_29660);
nor UO_189 (O_189,N_29768,N_29034);
xnor UO_190 (O_190,N_29594,N_29500);
nand UO_191 (O_191,N_28914,N_29648);
or UO_192 (O_192,N_29645,N_29053);
nor UO_193 (O_193,N_29490,N_29859);
or UO_194 (O_194,N_29471,N_29152);
nor UO_195 (O_195,N_29762,N_29273);
xor UO_196 (O_196,N_29743,N_28823);
nand UO_197 (O_197,N_29370,N_29817);
nand UO_198 (O_198,N_29577,N_29554);
or UO_199 (O_199,N_28913,N_29927);
nand UO_200 (O_200,N_29981,N_29776);
nand UO_201 (O_201,N_29456,N_28906);
nand UO_202 (O_202,N_29401,N_28875);
nand UO_203 (O_203,N_29514,N_29069);
nor UO_204 (O_204,N_29101,N_29808);
or UO_205 (O_205,N_29892,N_29784);
and UO_206 (O_206,N_29071,N_29666);
nand UO_207 (O_207,N_29288,N_29866);
or UO_208 (O_208,N_29264,N_29313);
nor UO_209 (O_209,N_29198,N_29735);
nor UO_210 (O_210,N_29213,N_29867);
xor UO_211 (O_211,N_28929,N_29560);
and UO_212 (O_212,N_28825,N_28826);
and UO_213 (O_213,N_29803,N_29267);
and UO_214 (O_214,N_28842,N_29656);
xnor UO_215 (O_215,N_29606,N_29536);
xnor UO_216 (O_216,N_29610,N_29074);
nand UO_217 (O_217,N_29954,N_28975);
nor UO_218 (O_218,N_29862,N_29142);
or UO_219 (O_219,N_29643,N_29825);
or UO_220 (O_220,N_29087,N_29237);
and UO_221 (O_221,N_29420,N_29840);
nand UO_222 (O_222,N_29677,N_28888);
xnor UO_223 (O_223,N_28859,N_29699);
xor UO_224 (O_224,N_29961,N_29297);
xnor UO_225 (O_225,N_29730,N_29747);
or UO_226 (O_226,N_29441,N_29770);
xor UO_227 (O_227,N_29723,N_29653);
nor UO_228 (O_228,N_29912,N_29830);
nand UO_229 (O_229,N_29737,N_29597);
xnor UO_230 (O_230,N_28853,N_29728);
and UO_231 (O_231,N_29703,N_29377);
nor UO_232 (O_232,N_29270,N_29617);
nand UO_233 (O_233,N_28876,N_29176);
nand UO_234 (O_234,N_28971,N_28839);
or UO_235 (O_235,N_28894,N_29558);
nor UO_236 (O_236,N_29127,N_29727);
nor UO_237 (O_237,N_29694,N_29413);
and UO_238 (O_238,N_29751,N_28950);
nor UO_239 (O_239,N_28860,N_29935);
nor UO_240 (O_240,N_29081,N_29312);
and UO_241 (O_241,N_29008,N_28910);
or UO_242 (O_242,N_29605,N_29404);
or UO_243 (O_243,N_29624,N_29168);
xnor UO_244 (O_244,N_28984,N_29845);
and UO_245 (O_245,N_29204,N_29103);
or UO_246 (O_246,N_29985,N_29161);
xor UO_247 (O_247,N_29246,N_29367);
and UO_248 (O_248,N_29326,N_29752);
or UO_249 (O_249,N_28982,N_28824);
nand UO_250 (O_250,N_29814,N_28889);
nand UO_251 (O_251,N_29235,N_29910);
nand UO_252 (O_252,N_29970,N_29089);
xnor UO_253 (O_253,N_28925,N_29468);
nor UO_254 (O_254,N_29155,N_29272);
and UO_255 (O_255,N_29697,N_28945);
nand UO_256 (O_256,N_29452,N_28827);
or UO_257 (O_257,N_28915,N_28974);
and UO_258 (O_258,N_29339,N_29309);
or UO_259 (O_259,N_29305,N_29491);
and UO_260 (O_260,N_29036,N_29603);
or UO_261 (O_261,N_28908,N_29679);
nor UO_262 (O_262,N_29592,N_29524);
nand UO_263 (O_263,N_29187,N_29415);
xnor UO_264 (O_264,N_29231,N_29868);
and UO_265 (O_265,N_28927,N_28867);
and UO_266 (O_266,N_28865,N_29805);
nor UO_267 (O_267,N_28983,N_28850);
xor UO_268 (O_268,N_29269,N_29007);
or UO_269 (O_269,N_29188,N_28806);
and UO_270 (O_270,N_28987,N_29780);
and UO_271 (O_271,N_29649,N_29121);
or UO_272 (O_272,N_29921,N_28834);
or UO_273 (O_273,N_29144,N_29629);
nor UO_274 (O_274,N_29725,N_29010);
and UO_275 (O_275,N_29260,N_29742);
or UO_276 (O_276,N_29960,N_29020);
nor UO_277 (O_277,N_29918,N_29779);
xor UO_278 (O_278,N_29470,N_29663);
and UO_279 (O_279,N_29946,N_29084);
nor UO_280 (O_280,N_29548,N_29193);
nand UO_281 (O_281,N_29518,N_29574);
and UO_282 (O_282,N_29166,N_29094);
xnor UO_283 (O_283,N_29766,N_29615);
and UO_284 (O_284,N_29106,N_28866);
or UO_285 (O_285,N_29710,N_29682);
or UO_286 (O_286,N_29327,N_29637);
xnor UO_287 (O_287,N_29657,N_29903);
nor UO_288 (O_288,N_29165,N_29240);
xor UO_289 (O_289,N_29521,N_29079);
or UO_290 (O_290,N_29052,N_29197);
nor UO_291 (O_291,N_29876,N_29561);
nand UO_292 (O_292,N_29484,N_29015);
and UO_293 (O_293,N_29258,N_28954);
nor UO_294 (O_294,N_29225,N_29925);
or UO_295 (O_295,N_29901,N_29444);
xnor UO_296 (O_296,N_29271,N_29027);
xor UO_297 (O_297,N_29848,N_29975);
or UO_298 (O_298,N_29744,N_29206);
or UO_299 (O_299,N_28833,N_28985);
xor UO_300 (O_300,N_29689,N_29685);
and UO_301 (O_301,N_29713,N_29393);
nor UO_302 (O_302,N_29018,N_29431);
nor UO_303 (O_303,N_29669,N_29890);
xor UO_304 (O_304,N_28845,N_28921);
nand UO_305 (O_305,N_29287,N_28965);
nor UO_306 (O_306,N_29414,N_29334);
nand UO_307 (O_307,N_29819,N_29581);
or UO_308 (O_308,N_29795,N_29982);
nor UO_309 (O_309,N_29012,N_28990);
and UO_310 (O_310,N_29520,N_28818);
nand UO_311 (O_311,N_29996,N_29937);
and UO_312 (O_312,N_29436,N_28832);
xor UO_313 (O_313,N_29885,N_29364);
nor UO_314 (O_314,N_28882,N_29931);
nor UO_315 (O_315,N_29447,N_29145);
nor UO_316 (O_316,N_29124,N_29612);
and UO_317 (O_317,N_29811,N_29196);
or UO_318 (O_318,N_29065,N_29705);
nor UO_319 (O_319,N_29062,N_29078);
and UO_320 (O_320,N_29839,N_29781);
xnor UO_321 (O_321,N_29457,N_28821);
and UO_322 (O_322,N_29244,N_29907);
nor UO_323 (O_323,N_29150,N_29802);
xor UO_324 (O_324,N_29157,N_29220);
xnor UO_325 (O_325,N_29895,N_29310);
nor UO_326 (O_326,N_29114,N_29450);
nand UO_327 (O_327,N_29822,N_29095);
xor UO_328 (O_328,N_28933,N_29733);
or UO_329 (O_329,N_28928,N_29797);
nor UO_330 (O_330,N_29318,N_29965);
nand UO_331 (O_331,N_29572,N_28841);
or UO_332 (O_332,N_29407,N_29869);
nand UO_333 (O_333,N_28904,N_29158);
nor UO_334 (O_334,N_29403,N_28808);
or UO_335 (O_335,N_29136,N_29619);
nand UO_336 (O_336,N_29658,N_28964);
and UO_337 (O_337,N_29625,N_29684);
xnor UO_338 (O_338,N_29794,N_29416);
and UO_339 (O_339,N_29537,N_29849);
nand UO_340 (O_340,N_28916,N_29384);
or UO_341 (O_341,N_29900,N_29745);
xnor UO_342 (O_342,N_29519,N_29642);
nand UO_343 (O_343,N_28836,N_29291);
or UO_344 (O_344,N_29608,N_29286);
xor UO_345 (O_345,N_29545,N_29836);
and UO_346 (O_346,N_29241,N_29429);
or UO_347 (O_347,N_29372,N_29578);
xor UO_348 (O_348,N_29964,N_29969);
and UO_349 (O_349,N_29879,N_29746);
xor UO_350 (O_350,N_28970,N_29120);
nand UO_351 (O_351,N_29362,N_29788);
and UO_352 (O_352,N_28872,N_29655);
nand UO_353 (O_353,N_29274,N_29896);
xnor UO_354 (O_354,N_29812,N_29353);
or UO_355 (O_355,N_29091,N_29013);
and UO_356 (O_356,N_29940,N_29164);
xnor UO_357 (O_357,N_28878,N_29016);
nand UO_358 (O_358,N_28893,N_29881);
xnor UO_359 (O_359,N_29458,N_29281);
or UO_360 (O_360,N_29445,N_29317);
and UO_361 (O_361,N_29257,N_29711);
or UO_362 (O_362,N_28881,N_29175);
nor UO_363 (O_363,N_28998,N_29219);
xor UO_364 (O_364,N_29055,N_29804);
nand UO_365 (O_365,N_29898,N_28896);
nand UO_366 (O_366,N_28811,N_29564);
or UO_367 (O_367,N_28937,N_28963);
and UO_368 (O_368,N_29417,N_29156);
nor UO_369 (O_369,N_29466,N_29266);
nand UO_370 (O_370,N_28991,N_29243);
nor UO_371 (O_371,N_29391,N_28887);
xor UO_372 (O_372,N_29023,N_28828);
and UO_373 (O_373,N_29321,N_28968);
nand UO_374 (O_374,N_29201,N_29021);
or UO_375 (O_375,N_29467,N_29167);
xnor UO_376 (O_376,N_29613,N_29465);
nand UO_377 (O_377,N_28822,N_29997);
nor UO_378 (O_378,N_29899,N_29210);
nand UO_379 (O_379,N_29054,N_29110);
nor UO_380 (O_380,N_28871,N_29348);
nand UO_381 (O_381,N_29938,N_29421);
xor UO_382 (O_382,N_29708,N_29073);
xnor UO_383 (O_383,N_29516,N_29338);
xor UO_384 (O_384,N_29306,N_29889);
xnor UO_385 (O_385,N_29551,N_29665);
xnor UO_386 (O_386,N_29761,N_29967);
nor UO_387 (O_387,N_29698,N_29341);
nor UO_388 (O_388,N_29100,N_29749);
nand UO_389 (O_389,N_29092,N_28838);
xor UO_390 (O_390,N_29568,N_29017);
or UO_391 (O_391,N_29397,N_29837);
nor UO_392 (O_392,N_29587,N_29593);
xor UO_393 (O_393,N_29181,N_29350);
nor UO_394 (O_394,N_29638,N_29987);
nor UO_395 (O_395,N_29148,N_29511);
nor UO_396 (O_396,N_29632,N_29496);
or UO_397 (O_397,N_29923,N_29979);
or UO_398 (O_398,N_29343,N_29807);
and UO_399 (O_399,N_29820,N_28844);
nor UO_400 (O_400,N_29672,N_29386);
and UO_401 (O_401,N_28936,N_29342);
or UO_402 (O_402,N_29096,N_29721);
nand UO_403 (O_403,N_29177,N_29842);
or UO_404 (O_404,N_29361,N_29759);
nand UO_405 (O_405,N_28898,N_29550);
nor UO_406 (O_406,N_29239,N_29358);
nand UO_407 (O_407,N_29533,N_29504);
xnor UO_408 (O_408,N_29557,N_28800);
xor UO_409 (O_409,N_28977,N_29614);
nand UO_410 (O_410,N_29159,N_29732);
nand UO_411 (O_411,N_29543,N_29002);
nor UO_412 (O_412,N_29477,N_29601);
and UO_413 (O_413,N_29691,N_29194);
nor UO_414 (O_414,N_29046,N_29432);
nor UO_415 (O_415,N_29086,N_29434);
nand UO_416 (O_416,N_28926,N_29740);
nor UO_417 (O_417,N_29212,N_29582);
nor UO_418 (O_418,N_29191,N_29346);
nand UO_419 (O_419,N_28932,N_29077);
or UO_420 (O_420,N_28958,N_29229);
nor UO_421 (O_421,N_29427,N_29333);
and UO_422 (O_422,N_28892,N_29451);
nand UO_423 (O_423,N_29552,N_29359);
and UO_424 (O_424,N_29712,N_29433);
xnor UO_425 (O_425,N_28877,N_29385);
xnor UO_426 (O_426,N_29828,N_29223);
nor UO_427 (O_427,N_29596,N_29463);
xnor UO_428 (O_428,N_29800,N_29618);
and UO_429 (O_429,N_29944,N_29276);
xnor UO_430 (O_430,N_29116,N_28880);
or UO_431 (O_431,N_28981,N_29644);
nand UO_432 (O_432,N_29872,N_29289);
or UO_433 (O_433,N_29410,N_28943);
nand UO_434 (O_434,N_29688,N_29493);
nor UO_435 (O_435,N_29195,N_29492);
and UO_436 (O_436,N_28902,N_29716);
nand UO_437 (O_437,N_29756,N_29854);
nand UO_438 (O_438,N_28847,N_29928);
nand UO_439 (O_439,N_28923,N_29230);
nor UO_440 (O_440,N_29547,N_29856);
or UO_441 (O_441,N_29835,N_29958);
nor UO_442 (O_442,N_29402,N_29284);
nand UO_443 (O_443,N_29000,N_29454);
and UO_444 (O_444,N_29584,N_29298);
xor UO_445 (O_445,N_29290,N_29236);
nand UO_446 (O_446,N_29039,N_29714);
nor UO_447 (O_447,N_29254,N_29942);
nand UO_448 (O_448,N_29382,N_29163);
or UO_449 (O_449,N_29576,N_29182);
nor UO_450 (O_450,N_29171,N_28807);
xor UO_451 (O_451,N_28922,N_29409);
nand UO_452 (O_452,N_29040,N_29860);
and UO_453 (O_453,N_29636,N_29609);
or UO_454 (O_454,N_29178,N_28973);
and UO_455 (O_455,N_28897,N_29067);
xnor UO_456 (O_456,N_29785,N_29777);
nor UO_457 (O_457,N_29990,N_29345);
xnor UO_458 (O_458,N_29112,N_29604);
and UO_459 (O_459,N_29991,N_29882);
nor UO_460 (O_460,N_29512,N_29681);
nor UO_461 (O_461,N_29786,N_28843);
nand UO_462 (O_462,N_28849,N_29902);
or UO_463 (O_463,N_29833,N_29586);
xor UO_464 (O_464,N_28939,N_28993);
xor UO_465 (O_465,N_29380,N_29395);
xnor UO_466 (O_466,N_29174,N_29790);
and UO_467 (O_467,N_29832,N_29184);
nand UO_468 (O_468,N_29850,N_29226);
xnor UO_469 (O_469,N_29823,N_29851);
xnor UO_470 (O_470,N_28855,N_29945);
or UO_471 (O_471,N_29948,N_28940);
nand UO_472 (O_472,N_29418,N_29765);
nand UO_473 (O_473,N_29559,N_29392);
nor UO_474 (O_474,N_29799,N_28909);
and UO_475 (O_475,N_29909,N_29874);
nand UO_476 (O_476,N_29172,N_29556);
and UO_477 (O_477,N_29030,N_29328);
and UO_478 (O_478,N_29097,N_29426);
xor UO_479 (O_479,N_29993,N_29789);
nand UO_480 (O_480,N_28891,N_29763);
nor UO_481 (O_481,N_29792,N_29293);
xor UO_482 (O_482,N_29296,N_29278);
xnor UO_483 (O_483,N_28941,N_29405);
nand UO_484 (O_484,N_28801,N_29980);
xnor UO_485 (O_485,N_28931,N_29959);
or UO_486 (O_486,N_28959,N_29224);
and UO_487 (O_487,N_28858,N_29755);
and UO_488 (O_488,N_28864,N_29192);
nor UO_489 (O_489,N_29316,N_29058);
and UO_490 (O_490,N_29183,N_29209);
nor UO_491 (O_491,N_29573,N_29739);
and UO_492 (O_492,N_29376,N_29858);
and UO_493 (O_493,N_29398,N_28938);
or UO_494 (O_494,N_29724,N_29908);
xor UO_495 (O_495,N_29428,N_28852);
nor UO_496 (O_496,N_28890,N_29115);
xnor UO_497 (O_497,N_28819,N_29773);
and UO_498 (O_498,N_29208,N_29406);
or UO_499 (O_499,N_28907,N_29134);
nand UO_500 (O_500,N_29675,N_28895);
xor UO_501 (O_501,N_29234,N_29639);
nor UO_502 (O_502,N_29473,N_29888);
nand UO_503 (O_503,N_29390,N_29853);
nor UO_504 (O_504,N_29838,N_29715);
and UO_505 (O_505,N_28986,N_29659);
nand UO_506 (O_506,N_28874,N_29599);
nand UO_507 (O_507,N_29816,N_29449);
nor UO_508 (O_508,N_29720,N_28805);
xnor UO_509 (O_509,N_28861,N_29253);
nand UO_510 (O_510,N_29033,N_29049);
nor UO_511 (O_511,N_29336,N_29419);
xor UO_512 (O_512,N_28901,N_29118);
or UO_513 (O_513,N_29205,N_29169);
and UO_514 (O_514,N_29535,N_29186);
nor UO_515 (O_515,N_28851,N_29320);
xnor UO_516 (O_516,N_29302,N_29469);
xor UO_517 (O_517,N_29680,N_28912);
nand UO_518 (O_518,N_29455,N_29489);
or UO_519 (O_519,N_29986,N_29430);
nand UO_520 (O_520,N_28829,N_29562);
nand UO_521 (O_521,N_29140,N_29344);
xnor UO_522 (O_522,N_29565,N_29381);
nand UO_523 (O_523,N_29878,N_29301);
nand UO_524 (O_524,N_29757,N_29911);
xor UO_525 (O_525,N_29906,N_29919);
and UO_526 (O_526,N_28942,N_29722);
and UO_527 (O_527,N_28869,N_29661);
or UO_528 (O_528,N_28803,N_29674);
and UO_529 (O_529,N_29764,N_29460);
xor UO_530 (O_530,N_29093,N_29662);
or UO_531 (O_531,N_29956,N_29412);
nand UO_532 (O_532,N_29873,N_29408);
nand UO_533 (O_533,N_29995,N_29818);
or UO_534 (O_534,N_29211,N_29704);
and UO_535 (O_535,N_29252,N_29886);
nor UO_536 (O_536,N_29810,N_29529);
xnor UO_537 (O_537,N_29729,N_29813);
or UO_538 (O_538,N_29352,N_29242);
xnor UO_539 (O_539,N_29180,N_29809);
nor UO_540 (O_540,N_29051,N_28817);
nor UO_541 (O_541,N_29349,N_28989);
nand UO_542 (O_542,N_29917,N_29009);
nor UO_543 (O_543,N_29989,N_29683);
or UO_544 (O_544,N_29479,N_29542);
nand UO_545 (O_545,N_29375,N_28868);
and UO_546 (O_546,N_29299,N_29050);
and UO_547 (O_547,N_29852,N_29829);
nand UO_548 (O_548,N_29024,N_29105);
nor UO_549 (O_549,N_29026,N_29620);
nand UO_550 (O_550,N_29549,N_29315);
nand UO_551 (O_551,N_29563,N_29135);
xnor UO_552 (O_552,N_29283,N_29129);
and UO_553 (O_553,N_28999,N_29102);
xnor UO_554 (O_554,N_29139,N_28830);
or UO_555 (O_555,N_29583,N_29806);
and UO_556 (O_556,N_29131,N_29268);
or UO_557 (O_557,N_28947,N_29488);
nor UO_558 (O_558,N_29190,N_29495);
xnor UO_559 (O_559,N_29279,N_29064);
nand UO_560 (O_560,N_28969,N_28994);
or UO_561 (O_561,N_29750,N_29038);
nand UO_562 (O_562,N_29971,N_29707);
and UO_563 (O_563,N_29778,N_29319);
or UO_564 (O_564,N_29952,N_29827);
xor UO_565 (O_565,N_29137,N_29011);
xnor UO_566 (O_566,N_28835,N_28802);
or UO_567 (O_567,N_29125,N_29905);
xor UO_568 (O_568,N_29793,N_29585);
xor UO_569 (O_569,N_29600,N_29082);
xor UO_570 (O_570,N_29676,N_28870);
or UO_571 (O_571,N_29001,N_28837);
nor UO_572 (O_572,N_28816,N_28899);
nand UO_573 (O_573,N_29934,N_29248);
and UO_574 (O_574,N_29531,N_29200);
nand UO_575 (O_575,N_29032,N_29277);
or UO_576 (O_576,N_29329,N_29107);
xor UO_577 (O_577,N_29443,N_29170);
xor UO_578 (O_578,N_29369,N_29978);
nor UO_579 (O_579,N_29532,N_28951);
nor UO_580 (O_580,N_29579,N_29098);
or UO_581 (O_581,N_28996,N_29335);
nor UO_582 (O_582,N_29772,N_29285);
nor UO_583 (O_583,N_29099,N_29791);
xor UO_584 (O_584,N_29149,N_29216);
and UO_585 (O_585,N_29508,N_29117);
or UO_586 (O_586,N_29108,N_29668);
and UO_587 (O_587,N_29941,N_29497);
or UO_588 (O_588,N_29047,N_29567);
xor UO_589 (O_589,N_29232,N_29400);
nand UO_590 (O_590,N_29357,N_28962);
or UO_591 (O_591,N_28804,N_29916);
nor UO_592 (O_592,N_29734,N_29153);
and UO_593 (O_593,N_29815,N_29503);
nor UO_594 (O_594,N_29486,N_28992);
nand UO_595 (O_595,N_29160,N_29111);
or UO_596 (O_596,N_29957,N_29955);
or UO_597 (O_597,N_29259,N_29976);
xnor UO_598 (O_598,N_29019,N_29437);
nor UO_599 (O_599,N_29066,N_29331);
and UO_600 (O_600,N_29678,N_29402);
or UO_601 (O_601,N_28831,N_29601);
or UO_602 (O_602,N_29714,N_29230);
xor UO_603 (O_603,N_28935,N_29019);
and UO_604 (O_604,N_29481,N_29170);
nor UO_605 (O_605,N_29622,N_29926);
nand UO_606 (O_606,N_29007,N_29262);
nor UO_607 (O_607,N_29947,N_29788);
nand UO_608 (O_608,N_28898,N_29045);
or UO_609 (O_609,N_29024,N_29081);
or UO_610 (O_610,N_29603,N_29763);
nor UO_611 (O_611,N_29170,N_29404);
nand UO_612 (O_612,N_29793,N_29747);
xnor UO_613 (O_613,N_29061,N_29081);
and UO_614 (O_614,N_29853,N_29464);
nand UO_615 (O_615,N_29103,N_29793);
and UO_616 (O_616,N_29357,N_29523);
and UO_617 (O_617,N_29634,N_29450);
and UO_618 (O_618,N_29203,N_28995);
or UO_619 (O_619,N_29533,N_29363);
xor UO_620 (O_620,N_29286,N_29491);
nand UO_621 (O_621,N_28848,N_29658);
nor UO_622 (O_622,N_29869,N_29953);
and UO_623 (O_623,N_29435,N_29216);
or UO_624 (O_624,N_29502,N_28893);
nand UO_625 (O_625,N_29472,N_29206);
or UO_626 (O_626,N_29787,N_29438);
and UO_627 (O_627,N_28916,N_29997);
and UO_628 (O_628,N_29915,N_29819);
or UO_629 (O_629,N_29584,N_29956);
or UO_630 (O_630,N_29101,N_29542);
nand UO_631 (O_631,N_29796,N_28880);
nand UO_632 (O_632,N_29429,N_29861);
nand UO_633 (O_633,N_28979,N_29640);
xnor UO_634 (O_634,N_29048,N_29091);
xor UO_635 (O_635,N_29890,N_28912);
or UO_636 (O_636,N_29507,N_29249);
xor UO_637 (O_637,N_28985,N_29039);
nor UO_638 (O_638,N_29435,N_28966);
or UO_639 (O_639,N_29708,N_29282);
xnor UO_640 (O_640,N_29774,N_29179);
xnor UO_641 (O_641,N_28868,N_29879);
xnor UO_642 (O_642,N_28813,N_29995);
xor UO_643 (O_643,N_29508,N_29665);
xor UO_644 (O_644,N_29816,N_29849);
or UO_645 (O_645,N_28814,N_29697);
or UO_646 (O_646,N_29576,N_29296);
and UO_647 (O_647,N_29668,N_28865);
nand UO_648 (O_648,N_29390,N_29668);
and UO_649 (O_649,N_29962,N_29506);
or UO_650 (O_650,N_29383,N_29006);
nor UO_651 (O_651,N_29532,N_29525);
and UO_652 (O_652,N_29154,N_29532);
nor UO_653 (O_653,N_29184,N_29739);
nor UO_654 (O_654,N_29999,N_29683);
xor UO_655 (O_655,N_29412,N_29416);
nor UO_656 (O_656,N_29905,N_29418);
and UO_657 (O_657,N_29416,N_28984);
or UO_658 (O_658,N_29164,N_29072);
nor UO_659 (O_659,N_29951,N_29063);
or UO_660 (O_660,N_29541,N_29793);
nand UO_661 (O_661,N_28920,N_29134);
or UO_662 (O_662,N_29997,N_28875);
nand UO_663 (O_663,N_29167,N_29655);
nor UO_664 (O_664,N_28805,N_29410);
or UO_665 (O_665,N_29139,N_29400);
or UO_666 (O_666,N_29639,N_28977);
nor UO_667 (O_667,N_29773,N_29163);
and UO_668 (O_668,N_29230,N_29823);
xor UO_669 (O_669,N_28923,N_29304);
nor UO_670 (O_670,N_29082,N_29478);
nor UO_671 (O_671,N_29673,N_29108);
or UO_672 (O_672,N_29162,N_28821);
or UO_673 (O_673,N_29848,N_29427);
or UO_674 (O_674,N_29672,N_29721);
nor UO_675 (O_675,N_29646,N_28874);
nand UO_676 (O_676,N_29739,N_28856);
xor UO_677 (O_677,N_29436,N_29071);
or UO_678 (O_678,N_29121,N_29465);
nand UO_679 (O_679,N_29205,N_29974);
nand UO_680 (O_680,N_29666,N_29434);
nor UO_681 (O_681,N_29652,N_29512);
and UO_682 (O_682,N_29159,N_29070);
nand UO_683 (O_683,N_29923,N_29763);
xnor UO_684 (O_684,N_29018,N_29707);
or UO_685 (O_685,N_29374,N_29920);
nor UO_686 (O_686,N_28814,N_29404);
and UO_687 (O_687,N_29837,N_29847);
and UO_688 (O_688,N_29214,N_29742);
nand UO_689 (O_689,N_28888,N_29493);
or UO_690 (O_690,N_29962,N_29567);
nand UO_691 (O_691,N_29170,N_28912);
and UO_692 (O_692,N_29909,N_29370);
or UO_693 (O_693,N_29741,N_29641);
nand UO_694 (O_694,N_29725,N_29470);
nor UO_695 (O_695,N_29997,N_29856);
nand UO_696 (O_696,N_29818,N_29381);
and UO_697 (O_697,N_29494,N_29086);
nor UO_698 (O_698,N_29554,N_29042);
nand UO_699 (O_699,N_29381,N_29017);
xnor UO_700 (O_700,N_29011,N_28820);
nor UO_701 (O_701,N_28817,N_29151);
or UO_702 (O_702,N_29127,N_28934);
or UO_703 (O_703,N_28955,N_29944);
nor UO_704 (O_704,N_29670,N_29068);
nor UO_705 (O_705,N_29481,N_28823);
nor UO_706 (O_706,N_28847,N_29492);
xor UO_707 (O_707,N_29137,N_29532);
xnor UO_708 (O_708,N_29294,N_29879);
xnor UO_709 (O_709,N_29555,N_29708);
xor UO_710 (O_710,N_29688,N_29976);
or UO_711 (O_711,N_29308,N_29120);
nor UO_712 (O_712,N_29189,N_29643);
or UO_713 (O_713,N_29626,N_29622);
and UO_714 (O_714,N_29462,N_28801);
and UO_715 (O_715,N_29853,N_29167);
and UO_716 (O_716,N_29277,N_29772);
nor UO_717 (O_717,N_29442,N_29634);
nor UO_718 (O_718,N_29390,N_29340);
nand UO_719 (O_719,N_29558,N_29568);
or UO_720 (O_720,N_29584,N_29087);
nor UO_721 (O_721,N_28874,N_28993);
xnor UO_722 (O_722,N_29410,N_29169);
nor UO_723 (O_723,N_28970,N_28940);
and UO_724 (O_724,N_28931,N_29444);
nor UO_725 (O_725,N_29054,N_29265);
nor UO_726 (O_726,N_29697,N_29067);
or UO_727 (O_727,N_28851,N_29816);
and UO_728 (O_728,N_29663,N_29158);
and UO_729 (O_729,N_29921,N_28963);
and UO_730 (O_730,N_29169,N_29886);
nand UO_731 (O_731,N_29778,N_29422);
and UO_732 (O_732,N_29826,N_29383);
nand UO_733 (O_733,N_29871,N_29550);
or UO_734 (O_734,N_29013,N_28920);
and UO_735 (O_735,N_29057,N_29857);
nor UO_736 (O_736,N_29636,N_29893);
nand UO_737 (O_737,N_29528,N_29591);
nand UO_738 (O_738,N_29867,N_28940);
xor UO_739 (O_739,N_29820,N_29215);
or UO_740 (O_740,N_29095,N_29759);
nor UO_741 (O_741,N_28919,N_29751);
nand UO_742 (O_742,N_29462,N_29829);
and UO_743 (O_743,N_28876,N_29433);
nand UO_744 (O_744,N_28960,N_29466);
and UO_745 (O_745,N_29089,N_29603);
xor UO_746 (O_746,N_29845,N_28977);
or UO_747 (O_747,N_29667,N_29145);
and UO_748 (O_748,N_29461,N_29403);
nor UO_749 (O_749,N_29222,N_29139);
xor UO_750 (O_750,N_28855,N_28862);
and UO_751 (O_751,N_29575,N_29491);
or UO_752 (O_752,N_29512,N_29466);
xnor UO_753 (O_753,N_29572,N_29501);
or UO_754 (O_754,N_29311,N_29119);
xnor UO_755 (O_755,N_29264,N_29635);
xor UO_756 (O_756,N_29006,N_28976);
and UO_757 (O_757,N_29645,N_29123);
nand UO_758 (O_758,N_29783,N_29725);
nand UO_759 (O_759,N_28959,N_29574);
and UO_760 (O_760,N_29642,N_29236);
nand UO_761 (O_761,N_29466,N_29569);
nor UO_762 (O_762,N_29445,N_29001);
or UO_763 (O_763,N_29874,N_29351);
nor UO_764 (O_764,N_29154,N_29706);
xor UO_765 (O_765,N_28927,N_29436);
nand UO_766 (O_766,N_29674,N_29554);
nor UO_767 (O_767,N_29020,N_29901);
nand UO_768 (O_768,N_28974,N_29734);
nor UO_769 (O_769,N_29545,N_29770);
nor UO_770 (O_770,N_29518,N_29930);
and UO_771 (O_771,N_29678,N_29948);
nor UO_772 (O_772,N_29639,N_29771);
and UO_773 (O_773,N_29729,N_29091);
nand UO_774 (O_774,N_28868,N_29789);
and UO_775 (O_775,N_29064,N_29114);
or UO_776 (O_776,N_29185,N_29567);
nor UO_777 (O_777,N_29048,N_29442);
nand UO_778 (O_778,N_29107,N_29168);
nor UO_779 (O_779,N_29590,N_29607);
nand UO_780 (O_780,N_29477,N_29415);
xnor UO_781 (O_781,N_29873,N_28916);
xor UO_782 (O_782,N_28967,N_29753);
xor UO_783 (O_783,N_29551,N_29870);
and UO_784 (O_784,N_29945,N_28956);
or UO_785 (O_785,N_28918,N_29650);
or UO_786 (O_786,N_29526,N_29755);
or UO_787 (O_787,N_29058,N_29190);
nor UO_788 (O_788,N_29118,N_29199);
nor UO_789 (O_789,N_29923,N_28873);
xnor UO_790 (O_790,N_29478,N_29722);
nand UO_791 (O_791,N_29241,N_29575);
nand UO_792 (O_792,N_29356,N_29462);
xor UO_793 (O_793,N_29709,N_29882);
nor UO_794 (O_794,N_29804,N_29405);
nor UO_795 (O_795,N_29456,N_29415);
xor UO_796 (O_796,N_29506,N_29871);
or UO_797 (O_797,N_29546,N_29305);
or UO_798 (O_798,N_29556,N_28825);
or UO_799 (O_799,N_29673,N_29903);
nand UO_800 (O_800,N_29107,N_29843);
nor UO_801 (O_801,N_28967,N_28929);
and UO_802 (O_802,N_29410,N_28948);
or UO_803 (O_803,N_29102,N_29861);
xnor UO_804 (O_804,N_29462,N_29353);
and UO_805 (O_805,N_28825,N_29872);
or UO_806 (O_806,N_29813,N_28861);
nand UO_807 (O_807,N_29811,N_29734);
or UO_808 (O_808,N_29320,N_29768);
nand UO_809 (O_809,N_29940,N_29199);
or UO_810 (O_810,N_29975,N_29774);
and UO_811 (O_811,N_28874,N_29847);
or UO_812 (O_812,N_29501,N_28833);
xnor UO_813 (O_813,N_29503,N_29792);
and UO_814 (O_814,N_29515,N_29473);
nand UO_815 (O_815,N_29629,N_29764);
or UO_816 (O_816,N_29460,N_29090);
and UO_817 (O_817,N_29560,N_29658);
and UO_818 (O_818,N_28809,N_29857);
xor UO_819 (O_819,N_29046,N_29851);
nand UO_820 (O_820,N_29597,N_28901);
nand UO_821 (O_821,N_29095,N_28912);
nor UO_822 (O_822,N_29541,N_29519);
nor UO_823 (O_823,N_29264,N_29380);
xnor UO_824 (O_824,N_29072,N_29278);
nand UO_825 (O_825,N_29184,N_29510);
nand UO_826 (O_826,N_29271,N_29227);
or UO_827 (O_827,N_29364,N_29571);
or UO_828 (O_828,N_29350,N_29492);
or UO_829 (O_829,N_29699,N_29533);
or UO_830 (O_830,N_29020,N_29377);
nand UO_831 (O_831,N_28961,N_28931);
nand UO_832 (O_832,N_29814,N_28891);
xor UO_833 (O_833,N_29837,N_29975);
nor UO_834 (O_834,N_29413,N_29296);
nand UO_835 (O_835,N_29472,N_29645);
nand UO_836 (O_836,N_29171,N_28840);
nand UO_837 (O_837,N_29590,N_28871);
or UO_838 (O_838,N_28876,N_29901);
nand UO_839 (O_839,N_29855,N_29471);
nor UO_840 (O_840,N_29464,N_29096);
nand UO_841 (O_841,N_29220,N_29691);
and UO_842 (O_842,N_29819,N_29811);
xor UO_843 (O_843,N_29444,N_29517);
nor UO_844 (O_844,N_29981,N_29511);
or UO_845 (O_845,N_29471,N_28856);
nor UO_846 (O_846,N_29058,N_29586);
xnor UO_847 (O_847,N_29456,N_29327);
nor UO_848 (O_848,N_29047,N_29934);
xor UO_849 (O_849,N_29894,N_29775);
nand UO_850 (O_850,N_28800,N_29266);
nand UO_851 (O_851,N_29261,N_29810);
and UO_852 (O_852,N_29919,N_29578);
and UO_853 (O_853,N_29566,N_28942);
and UO_854 (O_854,N_29776,N_29019);
xnor UO_855 (O_855,N_29466,N_29247);
or UO_856 (O_856,N_29289,N_29033);
or UO_857 (O_857,N_29864,N_29577);
or UO_858 (O_858,N_29385,N_29738);
nand UO_859 (O_859,N_29712,N_29856);
xnor UO_860 (O_860,N_29607,N_28851);
or UO_861 (O_861,N_29302,N_29188);
or UO_862 (O_862,N_29553,N_29704);
nor UO_863 (O_863,N_29099,N_29862);
xnor UO_864 (O_864,N_29603,N_29839);
or UO_865 (O_865,N_29533,N_28897);
nor UO_866 (O_866,N_29157,N_29563);
nor UO_867 (O_867,N_29048,N_29049);
xor UO_868 (O_868,N_29720,N_29282);
and UO_869 (O_869,N_29804,N_29215);
xnor UO_870 (O_870,N_29866,N_29952);
nor UO_871 (O_871,N_29557,N_29711);
xnor UO_872 (O_872,N_29363,N_29707);
xnor UO_873 (O_873,N_29193,N_29784);
xor UO_874 (O_874,N_29121,N_29127);
or UO_875 (O_875,N_28941,N_29873);
xor UO_876 (O_876,N_29892,N_29840);
and UO_877 (O_877,N_28915,N_29370);
nand UO_878 (O_878,N_29203,N_29405);
or UO_879 (O_879,N_29286,N_29021);
nand UO_880 (O_880,N_29763,N_29683);
or UO_881 (O_881,N_28965,N_29777);
nor UO_882 (O_882,N_29936,N_29964);
xor UO_883 (O_883,N_29290,N_29705);
nor UO_884 (O_884,N_29418,N_29435);
or UO_885 (O_885,N_29754,N_29178);
nand UO_886 (O_886,N_29935,N_29230);
and UO_887 (O_887,N_29001,N_29284);
or UO_888 (O_888,N_28863,N_29036);
or UO_889 (O_889,N_29120,N_29367);
nor UO_890 (O_890,N_29204,N_29616);
xnor UO_891 (O_891,N_29830,N_28872);
and UO_892 (O_892,N_29470,N_29539);
xnor UO_893 (O_893,N_29683,N_29411);
and UO_894 (O_894,N_29477,N_29713);
nor UO_895 (O_895,N_29068,N_28850);
nand UO_896 (O_896,N_29869,N_29810);
xor UO_897 (O_897,N_29429,N_28810);
and UO_898 (O_898,N_28908,N_29965);
nor UO_899 (O_899,N_28890,N_29499);
xnor UO_900 (O_900,N_28946,N_28943);
or UO_901 (O_901,N_29441,N_28805);
xor UO_902 (O_902,N_29101,N_29574);
or UO_903 (O_903,N_29272,N_29556);
nand UO_904 (O_904,N_29002,N_29006);
and UO_905 (O_905,N_29181,N_29020);
and UO_906 (O_906,N_29938,N_29435);
xnor UO_907 (O_907,N_29567,N_29190);
and UO_908 (O_908,N_28903,N_29681);
xor UO_909 (O_909,N_29250,N_29943);
and UO_910 (O_910,N_29753,N_28866);
and UO_911 (O_911,N_29061,N_29264);
xnor UO_912 (O_912,N_29925,N_29200);
or UO_913 (O_913,N_29343,N_29371);
and UO_914 (O_914,N_29866,N_29026);
and UO_915 (O_915,N_28851,N_29688);
or UO_916 (O_916,N_29014,N_29845);
nand UO_917 (O_917,N_29123,N_29302);
or UO_918 (O_918,N_29365,N_29355);
and UO_919 (O_919,N_29163,N_29979);
nor UO_920 (O_920,N_29378,N_29495);
xor UO_921 (O_921,N_29575,N_29006);
nor UO_922 (O_922,N_29376,N_29184);
xor UO_923 (O_923,N_28834,N_29141);
and UO_924 (O_924,N_29662,N_29153);
nand UO_925 (O_925,N_29455,N_29647);
and UO_926 (O_926,N_28828,N_29268);
or UO_927 (O_927,N_29332,N_28812);
nor UO_928 (O_928,N_29918,N_29756);
nand UO_929 (O_929,N_29827,N_29683);
xnor UO_930 (O_930,N_29056,N_29475);
or UO_931 (O_931,N_29534,N_29519);
or UO_932 (O_932,N_29251,N_29254);
or UO_933 (O_933,N_28910,N_29487);
nand UO_934 (O_934,N_29339,N_29874);
or UO_935 (O_935,N_29262,N_29958);
and UO_936 (O_936,N_29034,N_29321);
nand UO_937 (O_937,N_29768,N_29727);
nand UO_938 (O_938,N_29638,N_29682);
xnor UO_939 (O_939,N_29313,N_29057);
xor UO_940 (O_940,N_29953,N_28820);
and UO_941 (O_941,N_29713,N_29418);
xnor UO_942 (O_942,N_29021,N_29797);
nor UO_943 (O_943,N_29592,N_29466);
nor UO_944 (O_944,N_28913,N_29175);
xnor UO_945 (O_945,N_29148,N_29960);
xor UO_946 (O_946,N_29587,N_28877);
and UO_947 (O_947,N_29058,N_28939);
nor UO_948 (O_948,N_29089,N_28921);
or UO_949 (O_949,N_29806,N_29606);
xnor UO_950 (O_950,N_29375,N_28930);
xnor UO_951 (O_951,N_29428,N_29992);
nor UO_952 (O_952,N_29290,N_29394);
xnor UO_953 (O_953,N_29898,N_29514);
xor UO_954 (O_954,N_29287,N_28891);
xor UO_955 (O_955,N_29765,N_29557);
and UO_956 (O_956,N_29173,N_29067);
nor UO_957 (O_957,N_29068,N_29691);
nand UO_958 (O_958,N_29878,N_29885);
and UO_959 (O_959,N_29125,N_29950);
nor UO_960 (O_960,N_28850,N_29842);
nor UO_961 (O_961,N_29813,N_29104);
or UO_962 (O_962,N_29819,N_29111);
or UO_963 (O_963,N_29090,N_29625);
and UO_964 (O_964,N_28924,N_29428);
nor UO_965 (O_965,N_28989,N_29343);
nand UO_966 (O_966,N_29821,N_29207);
or UO_967 (O_967,N_29544,N_28950);
or UO_968 (O_968,N_29751,N_29395);
nand UO_969 (O_969,N_29931,N_29928);
and UO_970 (O_970,N_29923,N_28954);
or UO_971 (O_971,N_29997,N_29843);
and UO_972 (O_972,N_29720,N_29717);
nand UO_973 (O_973,N_28925,N_29255);
nand UO_974 (O_974,N_28874,N_29760);
nor UO_975 (O_975,N_28964,N_29876);
nand UO_976 (O_976,N_29690,N_29753);
and UO_977 (O_977,N_29296,N_29213);
and UO_978 (O_978,N_29841,N_29679);
xor UO_979 (O_979,N_29387,N_29507);
nor UO_980 (O_980,N_29628,N_29900);
xnor UO_981 (O_981,N_29970,N_28954);
nand UO_982 (O_982,N_29194,N_29401);
nand UO_983 (O_983,N_29561,N_29394);
and UO_984 (O_984,N_28808,N_29793);
nor UO_985 (O_985,N_29772,N_29036);
nand UO_986 (O_986,N_29341,N_29448);
nor UO_987 (O_987,N_29002,N_29284);
and UO_988 (O_988,N_29689,N_29747);
xor UO_989 (O_989,N_29325,N_29332);
nor UO_990 (O_990,N_29054,N_29891);
nor UO_991 (O_991,N_29767,N_29684);
or UO_992 (O_992,N_29331,N_29342);
and UO_993 (O_993,N_29595,N_29918);
or UO_994 (O_994,N_29755,N_29125);
nor UO_995 (O_995,N_29281,N_28913);
nor UO_996 (O_996,N_29735,N_29563);
and UO_997 (O_997,N_28962,N_29424);
xor UO_998 (O_998,N_28967,N_29212);
nand UO_999 (O_999,N_29019,N_29137);
nor UO_1000 (O_1000,N_29201,N_28984);
nand UO_1001 (O_1001,N_29005,N_29221);
nor UO_1002 (O_1002,N_29016,N_29152);
nand UO_1003 (O_1003,N_29998,N_29446);
and UO_1004 (O_1004,N_28937,N_29148);
or UO_1005 (O_1005,N_29681,N_28986);
xnor UO_1006 (O_1006,N_29873,N_28991);
nand UO_1007 (O_1007,N_29256,N_29263);
nor UO_1008 (O_1008,N_29361,N_29726);
and UO_1009 (O_1009,N_29008,N_29926);
xnor UO_1010 (O_1010,N_29464,N_29014);
nor UO_1011 (O_1011,N_29177,N_29828);
nand UO_1012 (O_1012,N_29363,N_29675);
or UO_1013 (O_1013,N_29966,N_29984);
nand UO_1014 (O_1014,N_29087,N_28840);
xor UO_1015 (O_1015,N_29020,N_28933);
or UO_1016 (O_1016,N_29144,N_29557);
nor UO_1017 (O_1017,N_29750,N_29136);
nand UO_1018 (O_1018,N_29513,N_29003);
nand UO_1019 (O_1019,N_29195,N_29385);
nand UO_1020 (O_1020,N_29939,N_29559);
nand UO_1021 (O_1021,N_29618,N_29481);
nand UO_1022 (O_1022,N_29764,N_29065);
nand UO_1023 (O_1023,N_29443,N_29362);
xor UO_1024 (O_1024,N_29203,N_29438);
nand UO_1025 (O_1025,N_29132,N_29597);
nand UO_1026 (O_1026,N_29125,N_29035);
and UO_1027 (O_1027,N_29812,N_29583);
xor UO_1028 (O_1028,N_28965,N_29097);
or UO_1029 (O_1029,N_29131,N_29725);
and UO_1030 (O_1030,N_29924,N_29920);
or UO_1031 (O_1031,N_29362,N_29185);
and UO_1032 (O_1032,N_29345,N_29580);
and UO_1033 (O_1033,N_29671,N_29304);
nand UO_1034 (O_1034,N_29290,N_29141);
nor UO_1035 (O_1035,N_28846,N_29298);
nor UO_1036 (O_1036,N_29598,N_29837);
xnor UO_1037 (O_1037,N_29580,N_29955);
or UO_1038 (O_1038,N_29428,N_29606);
and UO_1039 (O_1039,N_29230,N_29315);
xor UO_1040 (O_1040,N_28937,N_28839);
nor UO_1041 (O_1041,N_29854,N_29438);
and UO_1042 (O_1042,N_28944,N_29263);
nand UO_1043 (O_1043,N_28971,N_29188);
or UO_1044 (O_1044,N_29918,N_29816);
nor UO_1045 (O_1045,N_29612,N_29043);
nand UO_1046 (O_1046,N_29155,N_29646);
nand UO_1047 (O_1047,N_29396,N_29266);
xnor UO_1048 (O_1048,N_29934,N_29577);
xor UO_1049 (O_1049,N_29098,N_28985);
xor UO_1050 (O_1050,N_28823,N_29349);
nor UO_1051 (O_1051,N_29160,N_29821);
and UO_1052 (O_1052,N_29844,N_29445);
or UO_1053 (O_1053,N_29056,N_29064);
or UO_1054 (O_1054,N_29773,N_28945);
xnor UO_1055 (O_1055,N_29143,N_28807);
and UO_1056 (O_1056,N_29839,N_29042);
or UO_1057 (O_1057,N_29455,N_29306);
and UO_1058 (O_1058,N_29087,N_29259);
or UO_1059 (O_1059,N_29441,N_29458);
and UO_1060 (O_1060,N_29188,N_29415);
or UO_1061 (O_1061,N_28885,N_28982);
or UO_1062 (O_1062,N_28833,N_29578);
xnor UO_1063 (O_1063,N_29845,N_29556);
nor UO_1064 (O_1064,N_29770,N_29453);
nor UO_1065 (O_1065,N_29009,N_29269);
nor UO_1066 (O_1066,N_29248,N_29207);
or UO_1067 (O_1067,N_29033,N_28813);
nand UO_1068 (O_1068,N_29347,N_29505);
nand UO_1069 (O_1069,N_29240,N_29022);
or UO_1070 (O_1070,N_29973,N_29617);
and UO_1071 (O_1071,N_29957,N_29485);
nor UO_1072 (O_1072,N_29586,N_29977);
and UO_1073 (O_1073,N_29954,N_29461);
xor UO_1074 (O_1074,N_29661,N_29621);
xor UO_1075 (O_1075,N_29185,N_29522);
or UO_1076 (O_1076,N_29824,N_29281);
or UO_1077 (O_1077,N_29670,N_29837);
xor UO_1078 (O_1078,N_29331,N_29426);
nor UO_1079 (O_1079,N_28995,N_29426);
and UO_1080 (O_1080,N_29631,N_29283);
and UO_1081 (O_1081,N_29397,N_29322);
or UO_1082 (O_1082,N_29945,N_29764);
nor UO_1083 (O_1083,N_28913,N_29738);
nand UO_1084 (O_1084,N_29481,N_29544);
and UO_1085 (O_1085,N_29327,N_29189);
or UO_1086 (O_1086,N_28833,N_29197);
or UO_1087 (O_1087,N_29123,N_29847);
nor UO_1088 (O_1088,N_29041,N_29266);
nor UO_1089 (O_1089,N_29340,N_29290);
nor UO_1090 (O_1090,N_29228,N_29844);
nand UO_1091 (O_1091,N_29470,N_29241);
and UO_1092 (O_1092,N_28988,N_28802);
xor UO_1093 (O_1093,N_29523,N_29469);
xor UO_1094 (O_1094,N_29140,N_29784);
xor UO_1095 (O_1095,N_29350,N_29020);
nor UO_1096 (O_1096,N_29428,N_29391);
xnor UO_1097 (O_1097,N_29100,N_29340);
nand UO_1098 (O_1098,N_29742,N_29747);
and UO_1099 (O_1099,N_29773,N_29798);
nand UO_1100 (O_1100,N_29207,N_29611);
xor UO_1101 (O_1101,N_28937,N_29882);
nand UO_1102 (O_1102,N_29745,N_28858);
and UO_1103 (O_1103,N_29003,N_29933);
or UO_1104 (O_1104,N_29817,N_29518);
or UO_1105 (O_1105,N_29623,N_29291);
xor UO_1106 (O_1106,N_28801,N_29588);
nor UO_1107 (O_1107,N_29745,N_29295);
and UO_1108 (O_1108,N_29318,N_29787);
nor UO_1109 (O_1109,N_29515,N_28899);
and UO_1110 (O_1110,N_28903,N_29836);
or UO_1111 (O_1111,N_28909,N_28841);
nor UO_1112 (O_1112,N_29343,N_29287);
or UO_1113 (O_1113,N_29883,N_28803);
xor UO_1114 (O_1114,N_29077,N_29791);
and UO_1115 (O_1115,N_29294,N_29998);
and UO_1116 (O_1116,N_29796,N_29978);
nor UO_1117 (O_1117,N_28920,N_29717);
xnor UO_1118 (O_1118,N_29235,N_29341);
nor UO_1119 (O_1119,N_29167,N_29934);
or UO_1120 (O_1120,N_28800,N_29576);
or UO_1121 (O_1121,N_29654,N_29237);
nor UO_1122 (O_1122,N_29950,N_29165);
nand UO_1123 (O_1123,N_29012,N_29408);
nor UO_1124 (O_1124,N_28958,N_28854);
nand UO_1125 (O_1125,N_29244,N_29430);
nor UO_1126 (O_1126,N_29671,N_29463);
nor UO_1127 (O_1127,N_29993,N_28806);
nand UO_1128 (O_1128,N_29793,N_29947);
nand UO_1129 (O_1129,N_29434,N_29949);
or UO_1130 (O_1130,N_29988,N_29784);
and UO_1131 (O_1131,N_29307,N_29973);
xnor UO_1132 (O_1132,N_29765,N_29960);
nand UO_1133 (O_1133,N_29221,N_29044);
or UO_1134 (O_1134,N_29547,N_28936);
or UO_1135 (O_1135,N_29574,N_29375);
nand UO_1136 (O_1136,N_29718,N_29302);
nand UO_1137 (O_1137,N_29979,N_29378);
or UO_1138 (O_1138,N_28925,N_29487);
xor UO_1139 (O_1139,N_29754,N_28963);
xnor UO_1140 (O_1140,N_28920,N_29834);
xor UO_1141 (O_1141,N_29981,N_29854);
nor UO_1142 (O_1142,N_29643,N_29671);
nand UO_1143 (O_1143,N_29687,N_29020);
nand UO_1144 (O_1144,N_29540,N_29597);
nor UO_1145 (O_1145,N_29833,N_29981);
and UO_1146 (O_1146,N_28924,N_29274);
and UO_1147 (O_1147,N_29916,N_29621);
nor UO_1148 (O_1148,N_29023,N_29431);
nand UO_1149 (O_1149,N_29897,N_29640);
or UO_1150 (O_1150,N_28942,N_29420);
nand UO_1151 (O_1151,N_29932,N_29528);
nor UO_1152 (O_1152,N_29207,N_29182);
nor UO_1153 (O_1153,N_29739,N_29443);
nor UO_1154 (O_1154,N_29926,N_29532);
or UO_1155 (O_1155,N_29819,N_29397);
nor UO_1156 (O_1156,N_29765,N_28829);
or UO_1157 (O_1157,N_29740,N_28805);
and UO_1158 (O_1158,N_29275,N_29905);
xnor UO_1159 (O_1159,N_28823,N_29107);
nand UO_1160 (O_1160,N_29907,N_29571);
xnor UO_1161 (O_1161,N_28873,N_29645);
nor UO_1162 (O_1162,N_29108,N_29772);
and UO_1163 (O_1163,N_29674,N_29579);
nand UO_1164 (O_1164,N_29297,N_29764);
xor UO_1165 (O_1165,N_29673,N_29490);
or UO_1166 (O_1166,N_29551,N_29118);
nor UO_1167 (O_1167,N_29210,N_28836);
nand UO_1168 (O_1168,N_29143,N_29351);
nand UO_1169 (O_1169,N_28900,N_29226);
nor UO_1170 (O_1170,N_28906,N_29854);
and UO_1171 (O_1171,N_29652,N_29516);
xnor UO_1172 (O_1172,N_28966,N_29659);
or UO_1173 (O_1173,N_29773,N_29607);
xnor UO_1174 (O_1174,N_29531,N_28850);
and UO_1175 (O_1175,N_29588,N_29065);
nor UO_1176 (O_1176,N_29853,N_29460);
nor UO_1177 (O_1177,N_29701,N_28869);
or UO_1178 (O_1178,N_29527,N_29873);
xnor UO_1179 (O_1179,N_29292,N_29175);
xnor UO_1180 (O_1180,N_29290,N_29329);
and UO_1181 (O_1181,N_29648,N_29500);
xnor UO_1182 (O_1182,N_29869,N_29764);
nand UO_1183 (O_1183,N_29666,N_29898);
xnor UO_1184 (O_1184,N_29362,N_28913);
and UO_1185 (O_1185,N_28956,N_29845);
xor UO_1186 (O_1186,N_29971,N_28835);
nor UO_1187 (O_1187,N_28955,N_29456);
xor UO_1188 (O_1188,N_29986,N_29502);
nand UO_1189 (O_1189,N_29005,N_29782);
nand UO_1190 (O_1190,N_29104,N_29456);
and UO_1191 (O_1191,N_29466,N_29733);
and UO_1192 (O_1192,N_29119,N_29369);
and UO_1193 (O_1193,N_29738,N_29521);
or UO_1194 (O_1194,N_29472,N_29156);
nor UO_1195 (O_1195,N_29819,N_29453);
nor UO_1196 (O_1196,N_29025,N_29695);
nor UO_1197 (O_1197,N_29504,N_29661);
or UO_1198 (O_1198,N_29932,N_29450);
and UO_1199 (O_1199,N_29257,N_29160);
or UO_1200 (O_1200,N_29998,N_29438);
nor UO_1201 (O_1201,N_29494,N_28969);
xnor UO_1202 (O_1202,N_28877,N_28924);
xor UO_1203 (O_1203,N_29339,N_29391);
or UO_1204 (O_1204,N_29324,N_28904);
xor UO_1205 (O_1205,N_29380,N_29154);
and UO_1206 (O_1206,N_28992,N_29904);
and UO_1207 (O_1207,N_29674,N_29854);
xnor UO_1208 (O_1208,N_29569,N_29071);
and UO_1209 (O_1209,N_29894,N_28954);
nor UO_1210 (O_1210,N_29072,N_29202);
nand UO_1211 (O_1211,N_28920,N_29119);
nand UO_1212 (O_1212,N_29622,N_29382);
xor UO_1213 (O_1213,N_28861,N_29987);
or UO_1214 (O_1214,N_28807,N_29483);
xnor UO_1215 (O_1215,N_29508,N_29299);
nor UO_1216 (O_1216,N_29482,N_29930);
or UO_1217 (O_1217,N_29517,N_29955);
and UO_1218 (O_1218,N_29086,N_28867);
and UO_1219 (O_1219,N_28899,N_29928);
xnor UO_1220 (O_1220,N_29406,N_29716);
or UO_1221 (O_1221,N_29384,N_29314);
and UO_1222 (O_1222,N_29838,N_29566);
xnor UO_1223 (O_1223,N_28800,N_29797);
xor UO_1224 (O_1224,N_29445,N_29622);
nand UO_1225 (O_1225,N_29411,N_29649);
xnor UO_1226 (O_1226,N_29314,N_28849);
or UO_1227 (O_1227,N_29741,N_28833);
and UO_1228 (O_1228,N_28910,N_29221);
nor UO_1229 (O_1229,N_29417,N_28976);
nand UO_1230 (O_1230,N_29501,N_29688);
or UO_1231 (O_1231,N_29038,N_29356);
nand UO_1232 (O_1232,N_29380,N_29862);
nor UO_1233 (O_1233,N_28831,N_29162);
or UO_1234 (O_1234,N_29472,N_29675);
nand UO_1235 (O_1235,N_29659,N_29752);
and UO_1236 (O_1236,N_29631,N_29652);
xor UO_1237 (O_1237,N_29103,N_29659);
nor UO_1238 (O_1238,N_29993,N_29787);
nand UO_1239 (O_1239,N_29223,N_28881);
xor UO_1240 (O_1240,N_29571,N_28979);
nor UO_1241 (O_1241,N_29627,N_29799);
nor UO_1242 (O_1242,N_29969,N_29101);
or UO_1243 (O_1243,N_29069,N_28983);
nand UO_1244 (O_1244,N_29846,N_29099);
nor UO_1245 (O_1245,N_29699,N_29165);
nand UO_1246 (O_1246,N_29599,N_28891);
or UO_1247 (O_1247,N_29036,N_29307);
nor UO_1248 (O_1248,N_29143,N_29509);
or UO_1249 (O_1249,N_29876,N_28968);
and UO_1250 (O_1250,N_29151,N_29264);
xnor UO_1251 (O_1251,N_29357,N_29711);
and UO_1252 (O_1252,N_29391,N_29245);
xor UO_1253 (O_1253,N_29172,N_29215);
and UO_1254 (O_1254,N_29672,N_29269);
xor UO_1255 (O_1255,N_29203,N_29818);
xnor UO_1256 (O_1256,N_29066,N_29541);
nand UO_1257 (O_1257,N_29740,N_29868);
or UO_1258 (O_1258,N_29964,N_29026);
or UO_1259 (O_1259,N_28812,N_29451);
xnor UO_1260 (O_1260,N_28917,N_29950);
and UO_1261 (O_1261,N_29579,N_29328);
xor UO_1262 (O_1262,N_29124,N_29091);
xnor UO_1263 (O_1263,N_29734,N_29755);
nand UO_1264 (O_1264,N_29766,N_29360);
nor UO_1265 (O_1265,N_29927,N_29888);
nand UO_1266 (O_1266,N_28930,N_29820);
xnor UO_1267 (O_1267,N_29518,N_28882);
xor UO_1268 (O_1268,N_29472,N_29319);
and UO_1269 (O_1269,N_29516,N_28919);
nor UO_1270 (O_1270,N_29469,N_29384);
xor UO_1271 (O_1271,N_29858,N_29560);
or UO_1272 (O_1272,N_29158,N_29576);
nor UO_1273 (O_1273,N_29245,N_29095);
and UO_1274 (O_1274,N_29981,N_29130);
nand UO_1275 (O_1275,N_29564,N_29248);
nand UO_1276 (O_1276,N_28826,N_29814);
xor UO_1277 (O_1277,N_29428,N_29064);
xnor UO_1278 (O_1278,N_29465,N_29790);
nand UO_1279 (O_1279,N_29208,N_29772);
nor UO_1280 (O_1280,N_29855,N_29637);
xor UO_1281 (O_1281,N_29360,N_29111);
nor UO_1282 (O_1282,N_29523,N_29151);
or UO_1283 (O_1283,N_28998,N_29105);
nor UO_1284 (O_1284,N_29232,N_29370);
and UO_1285 (O_1285,N_28878,N_28954);
nor UO_1286 (O_1286,N_29400,N_29248);
xnor UO_1287 (O_1287,N_28833,N_29690);
and UO_1288 (O_1288,N_29055,N_29512);
and UO_1289 (O_1289,N_29438,N_29879);
nor UO_1290 (O_1290,N_29851,N_29838);
nor UO_1291 (O_1291,N_29878,N_28914);
nor UO_1292 (O_1292,N_29275,N_29882);
or UO_1293 (O_1293,N_28874,N_28823);
nand UO_1294 (O_1294,N_29530,N_29610);
xor UO_1295 (O_1295,N_29646,N_29745);
and UO_1296 (O_1296,N_29607,N_29629);
nor UO_1297 (O_1297,N_29627,N_29466);
and UO_1298 (O_1298,N_29851,N_29234);
xnor UO_1299 (O_1299,N_29004,N_28818);
nor UO_1300 (O_1300,N_29879,N_29395);
or UO_1301 (O_1301,N_29054,N_29021);
nand UO_1302 (O_1302,N_29058,N_29906);
or UO_1303 (O_1303,N_29064,N_29304);
or UO_1304 (O_1304,N_29215,N_29388);
and UO_1305 (O_1305,N_29717,N_28821);
nor UO_1306 (O_1306,N_28823,N_29335);
or UO_1307 (O_1307,N_29568,N_28985);
and UO_1308 (O_1308,N_29089,N_29285);
xor UO_1309 (O_1309,N_29780,N_29821);
or UO_1310 (O_1310,N_28920,N_28880);
nand UO_1311 (O_1311,N_29997,N_29274);
and UO_1312 (O_1312,N_29824,N_28949);
xor UO_1313 (O_1313,N_28888,N_29838);
nor UO_1314 (O_1314,N_29771,N_28977);
or UO_1315 (O_1315,N_28968,N_29994);
and UO_1316 (O_1316,N_29404,N_29950);
nor UO_1317 (O_1317,N_29696,N_29255);
or UO_1318 (O_1318,N_28996,N_29873);
and UO_1319 (O_1319,N_29602,N_29021);
xnor UO_1320 (O_1320,N_29449,N_29720);
nor UO_1321 (O_1321,N_29405,N_29799);
xor UO_1322 (O_1322,N_29962,N_29885);
nand UO_1323 (O_1323,N_29705,N_29181);
xnor UO_1324 (O_1324,N_28977,N_29360);
xnor UO_1325 (O_1325,N_29326,N_28873);
nor UO_1326 (O_1326,N_28831,N_29821);
and UO_1327 (O_1327,N_29618,N_29993);
and UO_1328 (O_1328,N_29808,N_29759);
or UO_1329 (O_1329,N_29873,N_29860);
xor UO_1330 (O_1330,N_29552,N_29655);
nand UO_1331 (O_1331,N_29571,N_28826);
nor UO_1332 (O_1332,N_28888,N_29256);
nand UO_1333 (O_1333,N_29658,N_29994);
nor UO_1334 (O_1334,N_28893,N_28988);
or UO_1335 (O_1335,N_29708,N_29601);
nand UO_1336 (O_1336,N_29777,N_29136);
nor UO_1337 (O_1337,N_29313,N_28812);
xnor UO_1338 (O_1338,N_29908,N_29382);
or UO_1339 (O_1339,N_29438,N_29790);
nand UO_1340 (O_1340,N_29422,N_29305);
xor UO_1341 (O_1341,N_29479,N_29535);
nor UO_1342 (O_1342,N_29828,N_28879);
nand UO_1343 (O_1343,N_29306,N_29435);
nand UO_1344 (O_1344,N_29575,N_29320);
nor UO_1345 (O_1345,N_29150,N_28885);
or UO_1346 (O_1346,N_29882,N_29322);
nand UO_1347 (O_1347,N_29942,N_29085);
or UO_1348 (O_1348,N_29243,N_29993);
xnor UO_1349 (O_1349,N_29039,N_29227);
and UO_1350 (O_1350,N_29603,N_29508);
nand UO_1351 (O_1351,N_29622,N_29922);
and UO_1352 (O_1352,N_28998,N_28851);
nor UO_1353 (O_1353,N_28844,N_29004);
nand UO_1354 (O_1354,N_28942,N_29235);
and UO_1355 (O_1355,N_29995,N_28915);
or UO_1356 (O_1356,N_29614,N_29210);
xnor UO_1357 (O_1357,N_29529,N_29941);
xnor UO_1358 (O_1358,N_29417,N_29511);
nor UO_1359 (O_1359,N_29296,N_28910);
or UO_1360 (O_1360,N_29475,N_29915);
nand UO_1361 (O_1361,N_29448,N_29307);
xor UO_1362 (O_1362,N_29688,N_29928);
or UO_1363 (O_1363,N_29825,N_28872);
or UO_1364 (O_1364,N_29775,N_29481);
xor UO_1365 (O_1365,N_29908,N_29498);
nor UO_1366 (O_1366,N_29185,N_28940);
nand UO_1367 (O_1367,N_29664,N_29545);
or UO_1368 (O_1368,N_28824,N_29816);
or UO_1369 (O_1369,N_29262,N_29127);
xnor UO_1370 (O_1370,N_29157,N_28968);
xnor UO_1371 (O_1371,N_29433,N_29568);
and UO_1372 (O_1372,N_29054,N_29731);
xnor UO_1373 (O_1373,N_28998,N_29220);
and UO_1374 (O_1374,N_29519,N_29416);
xor UO_1375 (O_1375,N_29964,N_28922);
nand UO_1376 (O_1376,N_29532,N_29625);
xor UO_1377 (O_1377,N_29499,N_29474);
nor UO_1378 (O_1378,N_29929,N_29891);
or UO_1379 (O_1379,N_28977,N_28860);
and UO_1380 (O_1380,N_28970,N_29616);
nor UO_1381 (O_1381,N_28926,N_28917);
and UO_1382 (O_1382,N_28935,N_29703);
nor UO_1383 (O_1383,N_29986,N_29289);
or UO_1384 (O_1384,N_29828,N_29594);
nor UO_1385 (O_1385,N_29297,N_29958);
nor UO_1386 (O_1386,N_29798,N_29239);
nor UO_1387 (O_1387,N_29971,N_29836);
or UO_1388 (O_1388,N_29418,N_28918);
xnor UO_1389 (O_1389,N_29100,N_29245);
and UO_1390 (O_1390,N_28893,N_28887);
xnor UO_1391 (O_1391,N_29415,N_29876);
xnor UO_1392 (O_1392,N_29850,N_29884);
or UO_1393 (O_1393,N_29903,N_29443);
or UO_1394 (O_1394,N_29151,N_29193);
or UO_1395 (O_1395,N_28971,N_28913);
or UO_1396 (O_1396,N_28958,N_29581);
xnor UO_1397 (O_1397,N_29375,N_29225);
or UO_1398 (O_1398,N_29497,N_28915);
nand UO_1399 (O_1399,N_29478,N_29791);
or UO_1400 (O_1400,N_28940,N_29145);
xor UO_1401 (O_1401,N_29854,N_29848);
and UO_1402 (O_1402,N_29063,N_29451);
nor UO_1403 (O_1403,N_29628,N_29481);
and UO_1404 (O_1404,N_29431,N_29637);
xnor UO_1405 (O_1405,N_29683,N_29724);
and UO_1406 (O_1406,N_29484,N_29194);
nand UO_1407 (O_1407,N_29868,N_29755);
nor UO_1408 (O_1408,N_29568,N_29136);
or UO_1409 (O_1409,N_29016,N_29056);
or UO_1410 (O_1410,N_29578,N_29856);
or UO_1411 (O_1411,N_29262,N_29729);
xnor UO_1412 (O_1412,N_29224,N_29547);
or UO_1413 (O_1413,N_29619,N_29092);
nand UO_1414 (O_1414,N_29644,N_28972);
or UO_1415 (O_1415,N_28964,N_29086);
nor UO_1416 (O_1416,N_29973,N_29750);
nor UO_1417 (O_1417,N_29029,N_28829);
or UO_1418 (O_1418,N_28834,N_29132);
and UO_1419 (O_1419,N_29765,N_29469);
xnor UO_1420 (O_1420,N_29230,N_29090);
or UO_1421 (O_1421,N_29656,N_29345);
or UO_1422 (O_1422,N_29524,N_29059);
nand UO_1423 (O_1423,N_29151,N_28865);
xor UO_1424 (O_1424,N_28862,N_29609);
nand UO_1425 (O_1425,N_28828,N_28831);
and UO_1426 (O_1426,N_28881,N_29920);
nand UO_1427 (O_1427,N_28852,N_29584);
or UO_1428 (O_1428,N_29757,N_29244);
xnor UO_1429 (O_1429,N_29413,N_29589);
nor UO_1430 (O_1430,N_29037,N_29806);
and UO_1431 (O_1431,N_29118,N_29780);
xnor UO_1432 (O_1432,N_29359,N_29269);
nand UO_1433 (O_1433,N_29222,N_29775);
and UO_1434 (O_1434,N_29978,N_29622);
nor UO_1435 (O_1435,N_29208,N_29719);
nor UO_1436 (O_1436,N_29095,N_29295);
xnor UO_1437 (O_1437,N_29260,N_29017);
nor UO_1438 (O_1438,N_28880,N_29203);
and UO_1439 (O_1439,N_29245,N_28994);
or UO_1440 (O_1440,N_29876,N_29493);
and UO_1441 (O_1441,N_29278,N_29653);
nand UO_1442 (O_1442,N_29149,N_29212);
xnor UO_1443 (O_1443,N_29732,N_29181);
and UO_1444 (O_1444,N_29867,N_29073);
nor UO_1445 (O_1445,N_29703,N_29697);
or UO_1446 (O_1446,N_29715,N_28893);
or UO_1447 (O_1447,N_28910,N_29717);
xor UO_1448 (O_1448,N_29934,N_29816);
and UO_1449 (O_1449,N_29595,N_29803);
or UO_1450 (O_1450,N_29427,N_29423);
and UO_1451 (O_1451,N_29804,N_29680);
nor UO_1452 (O_1452,N_28901,N_29795);
and UO_1453 (O_1453,N_29586,N_28929);
nand UO_1454 (O_1454,N_29175,N_29770);
nand UO_1455 (O_1455,N_28894,N_29544);
xnor UO_1456 (O_1456,N_29853,N_29958);
and UO_1457 (O_1457,N_28972,N_29928);
xnor UO_1458 (O_1458,N_29292,N_29177);
xor UO_1459 (O_1459,N_28894,N_29870);
or UO_1460 (O_1460,N_29889,N_29853);
or UO_1461 (O_1461,N_29932,N_29888);
nand UO_1462 (O_1462,N_29225,N_29280);
and UO_1463 (O_1463,N_29206,N_29131);
nor UO_1464 (O_1464,N_29598,N_29239);
nand UO_1465 (O_1465,N_29061,N_29082);
or UO_1466 (O_1466,N_29990,N_29882);
xor UO_1467 (O_1467,N_29239,N_28907);
and UO_1468 (O_1468,N_29474,N_28928);
and UO_1469 (O_1469,N_29858,N_29969);
xnor UO_1470 (O_1470,N_29002,N_29550);
and UO_1471 (O_1471,N_29948,N_28961);
or UO_1472 (O_1472,N_29871,N_29296);
and UO_1473 (O_1473,N_29552,N_28827);
or UO_1474 (O_1474,N_29349,N_29379);
nand UO_1475 (O_1475,N_28973,N_28960);
nand UO_1476 (O_1476,N_29469,N_29329);
or UO_1477 (O_1477,N_29492,N_29728);
xor UO_1478 (O_1478,N_29305,N_29728);
nor UO_1479 (O_1479,N_29961,N_29724);
xnor UO_1480 (O_1480,N_28803,N_29614);
nor UO_1481 (O_1481,N_29654,N_29260);
nor UO_1482 (O_1482,N_29493,N_29084);
and UO_1483 (O_1483,N_29328,N_29776);
nand UO_1484 (O_1484,N_29308,N_29665);
and UO_1485 (O_1485,N_29027,N_29736);
or UO_1486 (O_1486,N_29529,N_29775);
or UO_1487 (O_1487,N_29826,N_29866);
and UO_1488 (O_1488,N_29825,N_28825);
xor UO_1489 (O_1489,N_29510,N_29480);
nand UO_1490 (O_1490,N_29150,N_29014);
nand UO_1491 (O_1491,N_28841,N_29575);
nor UO_1492 (O_1492,N_29791,N_28855);
nor UO_1493 (O_1493,N_29712,N_29918);
or UO_1494 (O_1494,N_28868,N_29641);
nor UO_1495 (O_1495,N_29625,N_29798);
or UO_1496 (O_1496,N_29089,N_29236);
nand UO_1497 (O_1497,N_29905,N_29074);
xor UO_1498 (O_1498,N_29153,N_29981);
nand UO_1499 (O_1499,N_29111,N_29785);
or UO_1500 (O_1500,N_29339,N_29557);
nor UO_1501 (O_1501,N_29843,N_28844);
xor UO_1502 (O_1502,N_28984,N_29542);
and UO_1503 (O_1503,N_29084,N_29220);
or UO_1504 (O_1504,N_28955,N_29033);
or UO_1505 (O_1505,N_29695,N_28853);
xnor UO_1506 (O_1506,N_29846,N_29148);
nor UO_1507 (O_1507,N_29210,N_29803);
xnor UO_1508 (O_1508,N_29926,N_29327);
nand UO_1509 (O_1509,N_29847,N_29412);
nand UO_1510 (O_1510,N_29688,N_29942);
or UO_1511 (O_1511,N_29414,N_29276);
nor UO_1512 (O_1512,N_29669,N_29371);
or UO_1513 (O_1513,N_29769,N_29941);
and UO_1514 (O_1514,N_29581,N_29207);
xor UO_1515 (O_1515,N_29213,N_29433);
and UO_1516 (O_1516,N_29831,N_29714);
xor UO_1517 (O_1517,N_29596,N_29516);
or UO_1518 (O_1518,N_29621,N_29247);
nand UO_1519 (O_1519,N_29739,N_29614);
xor UO_1520 (O_1520,N_29865,N_29152);
xor UO_1521 (O_1521,N_29408,N_28850);
xnor UO_1522 (O_1522,N_29684,N_29385);
nor UO_1523 (O_1523,N_29411,N_29163);
nor UO_1524 (O_1524,N_28858,N_29132);
or UO_1525 (O_1525,N_29351,N_28919);
nand UO_1526 (O_1526,N_29211,N_29095);
nand UO_1527 (O_1527,N_29690,N_29416);
xnor UO_1528 (O_1528,N_29437,N_29395);
nor UO_1529 (O_1529,N_29824,N_29788);
xor UO_1530 (O_1530,N_29238,N_29084);
nor UO_1531 (O_1531,N_28998,N_29584);
xnor UO_1532 (O_1532,N_29803,N_29750);
and UO_1533 (O_1533,N_28943,N_28977);
and UO_1534 (O_1534,N_29799,N_29265);
and UO_1535 (O_1535,N_29928,N_29721);
or UO_1536 (O_1536,N_29701,N_29002);
and UO_1537 (O_1537,N_28802,N_28842);
nand UO_1538 (O_1538,N_29089,N_29780);
nand UO_1539 (O_1539,N_28875,N_29922);
nor UO_1540 (O_1540,N_29073,N_29327);
and UO_1541 (O_1541,N_29860,N_29134);
xnor UO_1542 (O_1542,N_29562,N_29986);
or UO_1543 (O_1543,N_29558,N_29837);
and UO_1544 (O_1544,N_28959,N_29264);
xnor UO_1545 (O_1545,N_29203,N_29878);
or UO_1546 (O_1546,N_29795,N_29396);
xor UO_1547 (O_1547,N_29746,N_29179);
xnor UO_1548 (O_1548,N_29005,N_29634);
nand UO_1549 (O_1549,N_29335,N_29479);
nand UO_1550 (O_1550,N_29585,N_29940);
or UO_1551 (O_1551,N_29045,N_29473);
and UO_1552 (O_1552,N_29936,N_28895);
xnor UO_1553 (O_1553,N_29260,N_29490);
and UO_1554 (O_1554,N_29346,N_28939);
and UO_1555 (O_1555,N_29164,N_29956);
xor UO_1556 (O_1556,N_29605,N_29033);
xor UO_1557 (O_1557,N_29328,N_29415);
nand UO_1558 (O_1558,N_29249,N_28944);
xnor UO_1559 (O_1559,N_29758,N_28900);
nand UO_1560 (O_1560,N_29501,N_29228);
nor UO_1561 (O_1561,N_29411,N_29675);
nand UO_1562 (O_1562,N_29956,N_29511);
xnor UO_1563 (O_1563,N_29119,N_29267);
nor UO_1564 (O_1564,N_29347,N_29880);
xor UO_1565 (O_1565,N_29108,N_29245);
xnor UO_1566 (O_1566,N_28924,N_28838);
xor UO_1567 (O_1567,N_29986,N_29824);
nand UO_1568 (O_1568,N_29857,N_28985);
or UO_1569 (O_1569,N_29900,N_28824);
nand UO_1570 (O_1570,N_29861,N_29976);
or UO_1571 (O_1571,N_29830,N_28998);
nor UO_1572 (O_1572,N_29862,N_29005);
and UO_1573 (O_1573,N_29727,N_28830);
and UO_1574 (O_1574,N_28802,N_29136);
nor UO_1575 (O_1575,N_28969,N_29233);
xor UO_1576 (O_1576,N_29929,N_28932);
and UO_1577 (O_1577,N_29549,N_29711);
and UO_1578 (O_1578,N_29430,N_29556);
or UO_1579 (O_1579,N_29050,N_28981);
nor UO_1580 (O_1580,N_29113,N_29590);
nand UO_1581 (O_1581,N_29753,N_29417);
nor UO_1582 (O_1582,N_29612,N_29466);
or UO_1583 (O_1583,N_29935,N_29310);
xor UO_1584 (O_1584,N_29462,N_29589);
nand UO_1585 (O_1585,N_29459,N_29417);
nand UO_1586 (O_1586,N_28965,N_29650);
xnor UO_1587 (O_1587,N_29762,N_29374);
nand UO_1588 (O_1588,N_29917,N_29515);
nand UO_1589 (O_1589,N_28912,N_29855);
nor UO_1590 (O_1590,N_29023,N_29269);
nor UO_1591 (O_1591,N_29756,N_29704);
xnor UO_1592 (O_1592,N_29488,N_29762);
and UO_1593 (O_1593,N_29838,N_29574);
xnor UO_1594 (O_1594,N_29810,N_29666);
xnor UO_1595 (O_1595,N_29607,N_29654);
xor UO_1596 (O_1596,N_29321,N_29643);
or UO_1597 (O_1597,N_29439,N_29872);
nor UO_1598 (O_1598,N_29914,N_29481);
nand UO_1599 (O_1599,N_29817,N_29561);
nand UO_1600 (O_1600,N_29222,N_29067);
xor UO_1601 (O_1601,N_29149,N_29236);
and UO_1602 (O_1602,N_29014,N_29740);
or UO_1603 (O_1603,N_28807,N_29318);
nand UO_1604 (O_1604,N_29622,N_29665);
or UO_1605 (O_1605,N_29217,N_29890);
or UO_1606 (O_1606,N_29884,N_29961);
nor UO_1607 (O_1607,N_29616,N_29231);
and UO_1608 (O_1608,N_29224,N_29516);
or UO_1609 (O_1609,N_29167,N_29794);
and UO_1610 (O_1610,N_29565,N_29855);
nand UO_1611 (O_1611,N_29736,N_29851);
nor UO_1612 (O_1612,N_29669,N_28901);
and UO_1613 (O_1613,N_28946,N_29014);
and UO_1614 (O_1614,N_29385,N_29254);
nor UO_1615 (O_1615,N_29194,N_29705);
or UO_1616 (O_1616,N_29509,N_29250);
or UO_1617 (O_1617,N_28825,N_29580);
or UO_1618 (O_1618,N_29152,N_29921);
and UO_1619 (O_1619,N_29266,N_29620);
and UO_1620 (O_1620,N_29976,N_28932);
or UO_1621 (O_1621,N_29532,N_29471);
nand UO_1622 (O_1622,N_29762,N_29904);
nor UO_1623 (O_1623,N_29052,N_29442);
or UO_1624 (O_1624,N_28989,N_29637);
nor UO_1625 (O_1625,N_29305,N_28860);
xor UO_1626 (O_1626,N_29901,N_29255);
xor UO_1627 (O_1627,N_29388,N_29342);
and UO_1628 (O_1628,N_29678,N_29769);
and UO_1629 (O_1629,N_29179,N_29576);
or UO_1630 (O_1630,N_29657,N_29217);
xor UO_1631 (O_1631,N_29584,N_29226);
nor UO_1632 (O_1632,N_29179,N_29551);
nand UO_1633 (O_1633,N_28938,N_28805);
and UO_1634 (O_1634,N_29597,N_29301);
xnor UO_1635 (O_1635,N_28842,N_29782);
nor UO_1636 (O_1636,N_29955,N_29345);
or UO_1637 (O_1637,N_29457,N_29422);
or UO_1638 (O_1638,N_29787,N_29164);
nor UO_1639 (O_1639,N_29603,N_29293);
or UO_1640 (O_1640,N_29200,N_29077);
and UO_1641 (O_1641,N_29854,N_29425);
nor UO_1642 (O_1642,N_29625,N_29998);
or UO_1643 (O_1643,N_29902,N_28858);
and UO_1644 (O_1644,N_29949,N_28983);
nand UO_1645 (O_1645,N_29225,N_29996);
nor UO_1646 (O_1646,N_29034,N_29455);
nand UO_1647 (O_1647,N_29852,N_29029);
nand UO_1648 (O_1648,N_29252,N_29707);
nor UO_1649 (O_1649,N_29232,N_29008);
or UO_1650 (O_1650,N_29072,N_29635);
xnor UO_1651 (O_1651,N_29940,N_29516);
nor UO_1652 (O_1652,N_29395,N_29726);
or UO_1653 (O_1653,N_29323,N_29513);
and UO_1654 (O_1654,N_29806,N_29809);
xor UO_1655 (O_1655,N_29850,N_29231);
nor UO_1656 (O_1656,N_29473,N_29934);
nor UO_1657 (O_1657,N_29612,N_28951);
nor UO_1658 (O_1658,N_29391,N_28982);
or UO_1659 (O_1659,N_29243,N_29570);
or UO_1660 (O_1660,N_29855,N_29729);
nand UO_1661 (O_1661,N_28888,N_28839);
and UO_1662 (O_1662,N_29991,N_29849);
nor UO_1663 (O_1663,N_29979,N_29698);
nor UO_1664 (O_1664,N_29763,N_29496);
or UO_1665 (O_1665,N_29309,N_29342);
nor UO_1666 (O_1666,N_29288,N_29439);
and UO_1667 (O_1667,N_28846,N_29763);
xnor UO_1668 (O_1668,N_29475,N_28975);
xor UO_1669 (O_1669,N_28839,N_29347);
nand UO_1670 (O_1670,N_29073,N_29341);
nand UO_1671 (O_1671,N_29737,N_29122);
or UO_1672 (O_1672,N_28984,N_29238);
and UO_1673 (O_1673,N_28899,N_28804);
nor UO_1674 (O_1674,N_28827,N_28802);
nor UO_1675 (O_1675,N_29637,N_29875);
and UO_1676 (O_1676,N_29641,N_29445);
nand UO_1677 (O_1677,N_29851,N_28999);
xor UO_1678 (O_1678,N_29293,N_29996);
nor UO_1679 (O_1679,N_29339,N_29802);
xnor UO_1680 (O_1680,N_29764,N_29970);
nand UO_1681 (O_1681,N_29439,N_29529);
xor UO_1682 (O_1682,N_29578,N_29115);
nand UO_1683 (O_1683,N_28926,N_28825);
and UO_1684 (O_1684,N_29461,N_29282);
or UO_1685 (O_1685,N_28860,N_29301);
nand UO_1686 (O_1686,N_29963,N_29472);
and UO_1687 (O_1687,N_29875,N_29888);
xnor UO_1688 (O_1688,N_28994,N_29752);
xnor UO_1689 (O_1689,N_29228,N_28947);
or UO_1690 (O_1690,N_29564,N_29053);
nor UO_1691 (O_1691,N_29933,N_29235);
xnor UO_1692 (O_1692,N_29036,N_29113);
and UO_1693 (O_1693,N_29747,N_28978);
nand UO_1694 (O_1694,N_28813,N_29881);
xnor UO_1695 (O_1695,N_29712,N_29150);
nor UO_1696 (O_1696,N_29512,N_29317);
and UO_1697 (O_1697,N_29692,N_29099);
and UO_1698 (O_1698,N_29152,N_29496);
xnor UO_1699 (O_1699,N_29394,N_29989);
nand UO_1700 (O_1700,N_29607,N_29168);
or UO_1701 (O_1701,N_29296,N_29075);
or UO_1702 (O_1702,N_29368,N_29738);
xnor UO_1703 (O_1703,N_29576,N_29793);
and UO_1704 (O_1704,N_28994,N_29264);
or UO_1705 (O_1705,N_29230,N_29300);
nand UO_1706 (O_1706,N_29783,N_29178);
nor UO_1707 (O_1707,N_29027,N_29863);
or UO_1708 (O_1708,N_29267,N_29494);
nand UO_1709 (O_1709,N_29302,N_29994);
nor UO_1710 (O_1710,N_29351,N_29391);
or UO_1711 (O_1711,N_28831,N_29132);
xor UO_1712 (O_1712,N_29220,N_29496);
nor UO_1713 (O_1713,N_29619,N_29952);
and UO_1714 (O_1714,N_29831,N_29780);
or UO_1715 (O_1715,N_29419,N_29019);
nand UO_1716 (O_1716,N_29301,N_29313);
or UO_1717 (O_1717,N_29099,N_29977);
nand UO_1718 (O_1718,N_29524,N_29746);
nor UO_1719 (O_1719,N_28836,N_29613);
nor UO_1720 (O_1720,N_29235,N_28935);
nand UO_1721 (O_1721,N_29977,N_28838);
xnor UO_1722 (O_1722,N_29778,N_28965);
nor UO_1723 (O_1723,N_29612,N_29267);
nand UO_1724 (O_1724,N_29212,N_29322);
nand UO_1725 (O_1725,N_29742,N_29098);
and UO_1726 (O_1726,N_29452,N_29105);
and UO_1727 (O_1727,N_29376,N_29460);
and UO_1728 (O_1728,N_29839,N_29892);
or UO_1729 (O_1729,N_29950,N_29674);
and UO_1730 (O_1730,N_29861,N_29073);
or UO_1731 (O_1731,N_28997,N_29029);
xnor UO_1732 (O_1732,N_29592,N_29640);
nand UO_1733 (O_1733,N_29491,N_28920);
xor UO_1734 (O_1734,N_29606,N_29009);
nand UO_1735 (O_1735,N_29348,N_28842);
and UO_1736 (O_1736,N_28857,N_28874);
xor UO_1737 (O_1737,N_29443,N_29411);
and UO_1738 (O_1738,N_28882,N_29352);
and UO_1739 (O_1739,N_29653,N_29440);
or UO_1740 (O_1740,N_28880,N_29212);
xor UO_1741 (O_1741,N_28869,N_29144);
xnor UO_1742 (O_1742,N_28868,N_29445);
nor UO_1743 (O_1743,N_29547,N_29238);
and UO_1744 (O_1744,N_29246,N_28817);
nor UO_1745 (O_1745,N_29890,N_29071);
and UO_1746 (O_1746,N_29051,N_29425);
nand UO_1747 (O_1747,N_29115,N_29297);
and UO_1748 (O_1748,N_29806,N_28888);
xor UO_1749 (O_1749,N_29106,N_29867);
or UO_1750 (O_1750,N_29777,N_29551);
and UO_1751 (O_1751,N_29356,N_29233);
nor UO_1752 (O_1752,N_29642,N_29399);
xor UO_1753 (O_1753,N_29235,N_29557);
xor UO_1754 (O_1754,N_28839,N_29404);
nand UO_1755 (O_1755,N_29985,N_28980);
and UO_1756 (O_1756,N_28941,N_29278);
nor UO_1757 (O_1757,N_29910,N_29990);
xor UO_1758 (O_1758,N_29725,N_29776);
or UO_1759 (O_1759,N_29484,N_28833);
or UO_1760 (O_1760,N_29918,N_29857);
xor UO_1761 (O_1761,N_28815,N_29739);
and UO_1762 (O_1762,N_29276,N_29055);
or UO_1763 (O_1763,N_29606,N_29268);
and UO_1764 (O_1764,N_29585,N_29802);
and UO_1765 (O_1765,N_29130,N_29787);
nand UO_1766 (O_1766,N_29593,N_29080);
nor UO_1767 (O_1767,N_29193,N_28978);
xor UO_1768 (O_1768,N_29947,N_29875);
or UO_1769 (O_1769,N_28994,N_29569);
and UO_1770 (O_1770,N_29880,N_28930);
nand UO_1771 (O_1771,N_29890,N_28892);
and UO_1772 (O_1772,N_29919,N_29046);
nand UO_1773 (O_1773,N_29724,N_29575);
nor UO_1774 (O_1774,N_29217,N_29460);
or UO_1775 (O_1775,N_29858,N_29740);
nand UO_1776 (O_1776,N_29223,N_29929);
nand UO_1777 (O_1777,N_29916,N_29813);
and UO_1778 (O_1778,N_29946,N_28980);
nor UO_1779 (O_1779,N_29180,N_29166);
nand UO_1780 (O_1780,N_29062,N_29958);
or UO_1781 (O_1781,N_29336,N_29414);
and UO_1782 (O_1782,N_28885,N_29692);
or UO_1783 (O_1783,N_29304,N_29446);
xnor UO_1784 (O_1784,N_29317,N_28937);
nor UO_1785 (O_1785,N_29563,N_29041);
xnor UO_1786 (O_1786,N_29572,N_29095);
or UO_1787 (O_1787,N_29618,N_28856);
nand UO_1788 (O_1788,N_29137,N_29319);
and UO_1789 (O_1789,N_29781,N_29261);
and UO_1790 (O_1790,N_29494,N_28852);
xor UO_1791 (O_1791,N_29476,N_29640);
nand UO_1792 (O_1792,N_28809,N_28901);
nand UO_1793 (O_1793,N_29610,N_29123);
or UO_1794 (O_1794,N_29040,N_29205);
and UO_1795 (O_1795,N_29520,N_29500);
xnor UO_1796 (O_1796,N_29283,N_29189);
xor UO_1797 (O_1797,N_29996,N_28916);
nand UO_1798 (O_1798,N_29382,N_29320);
nor UO_1799 (O_1799,N_29668,N_29296);
and UO_1800 (O_1800,N_28931,N_29336);
xor UO_1801 (O_1801,N_29203,N_29471);
xnor UO_1802 (O_1802,N_29758,N_28860);
nor UO_1803 (O_1803,N_29432,N_28981);
xnor UO_1804 (O_1804,N_29802,N_29988);
or UO_1805 (O_1805,N_29533,N_29277);
or UO_1806 (O_1806,N_29766,N_28810);
nand UO_1807 (O_1807,N_29458,N_29929);
and UO_1808 (O_1808,N_29933,N_29742);
nand UO_1809 (O_1809,N_29603,N_29114);
or UO_1810 (O_1810,N_29855,N_29719);
nor UO_1811 (O_1811,N_28998,N_28907);
or UO_1812 (O_1812,N_29005,N_28830);
nand UO_1813 (O_1813,N_29314,N_29834);
or UO_1814 (O_1814,N_29857,N_29268);
xnor UO_1815 (O_1815,N_28874,N_29108);
nand UO_1816 (O_1816,N_29951,N_29059);
and UO_1817 (O_1817,N_28904,N_29423);
xor UO_1818 (O_1818,N_29724,N_29285);
nand UO_1819 (O_1819,N_29830,N_29913);
or UO_1820 (O_1820,N_29441,N_29152);
nor UO_1821 (O_1821,N_29541,N_28943);
nor UO_1822 (O_1822,N_29612,N_29831);
xor UO_1823 (O_1823,N_29651,N_29450);
xnor UO_1824 (O_1824,N_29769,N_28932);
nand UO_1825 (O_1825,N_29401,N_29964);
or UO_1826 (O_1826,N_28943,N_29136);
nand UO_1827 (O_1827,N_28982,N_29248);
nand UO_1828 (O_1828,N_29676,N_29548);
and UO_1829 (O_1829,N_29366,N_29033);
xor UO_1830 (O_1830,N_28858,N_29339);
nand UO_1831 (O_1831,N_28970,N_29587);
nor UO_1832 (O_1832,N_29120,N_28917);
or UO_1833 (O_1833,N_29736,N_29467);
nand UO_1834 (O_1834,N_28970,N_29079);
nand UO_1835 (O_1835,N_29251,N_29515);
nand UO_1836 (O_1836,N_29114,N_29334);
and UO_1837 (O_1837,N_29771,N_28807);
or UO_1838 (O_1838,N_29908,N_28876);
or UO_1839 (O_1839,N_29083,N_29125);
xnor UO_1840 (O_1840,N_29181,N_29358);
nand UO_1841 (O_1841,N_29875,N_28820);
or UO_1842 (O_1842,N_28814,N_29146);
xnor UO_1843 (O_1843,N_29725,N_29658);
and UO_1844 (O_1844,N_29299,N_28907);
nor UO_1845 (O_1845,N_29035,N_29461);
nor UO_1846 (O_1846,N_29547,N_29061);
nor UO_1847 (O_1847,N_29593,N_29097);
xnor UO_1848 (O_1848,N_28974,N_29121);
or UO_1849 (O_1849,N_29352,N_29323);
nor UO_1850 (O_1850,N_29019,N_29014);
xor UO_1851 (O_1851,N_29018,N_28874);
xor UO_1852 (O_1852,N_29533,N_29874);
nand UO_1853 (O_1853,N_29078,N_29583);
nand UO_1854 (O_1854,N_29400,N_29949);
nor UO_1855 (O_1855,N_29941,N_29924);
nand UO_1856 (O_1856,N_29615,N_29143);
or UO_1857 (O_1857,N_29710,N_29650);
and UO_1858 (O_1858,N_29083,N_28911);
xor UO_1859 (O_1859,N_29836,N_29228);
xor UO_1860 (O_1860,N_29986,N_29095);
xnor UO_1861 (O_1861,N_29715,N_29298);
xor UO_1862 (O_1862,N_29746,N_29506);
or UO_1863 (O_1863,N_29692,N_28991);
nor UO_1864 (O_1864,N_29249,N_29243);
nor UO_1865 (O_1865,N_29898,N_29897);
and UO_1866 (O_1866,N_29522,N_29376);
nand UO_1867 (O_1867,N_29941,N_29456);
and UO_1868 (O_1868,N_28922,N_28883);
nor UO_1869 (O_1869,N_29577,N_28818);
nor UO_1870 (O_1870,N_28870,N_29789);
or UO_1871 (O_1871,N_29636,N_29958);
xor UO_1872 (O_1872,N_29086,N_29089);
xor UO_1873 (O_1873,N_29100,N_29627);
xor UO_1874 (O_1874,N_29734,N_29698);
nor UO_1875 (O_1875,N_29240,N_29678);
and UO_1876 (O_1876,N_28819,N_28999);
nand UO_1877 (O_1877,N_28894,N_29205);
and UO_1878 (O_1878,N_29731,N_29946);
or UO_1879 (O_1879,N_29162,N_29248);
nor UO_1880 (O_1880,N_28847,N_28930);
nand UO_1881 (O_1881,N_29715,N_29897);
nor UO_1882 (O_1882,N_29907,N_29286);
or UO_1883 (O_1883,N_29665,N_29601);
nand UO_1884 (O_1884,N_29214,N_29130);
and UO_1885 (O_1885,N_29988,N_29375);
nor UO_1886 (O_1886,N_28918,N_29366);
xnor UO_1887 (O_1887,N_29566,N_29356);
nand UO_1888 (O_1888,N_29934,N_29911);
nor UO_1889 (O_1889,N_29020,N_28871);
nor UO_1890 (O_1890,N_29043,N_29574);
xor UO_1891 (O_1891,N_29016,N_29285);
or UO_1892 (O_1892,N_29960,N_29214);
and UO_1893 (O_1893,N_29859,N_29090);
xor UO_1894 (O_1894,N_28864,N_29565);
and UO_1895 (O_1895,N_29534,N_29184);
or UO_1896 (O_1896,N_29820,N_29971);
and UO_1897 (O_1897,N_29503,N_29918);
nor UO_1898 (O_1898,N_29825,N_29621);
nand UO_1899 (O_1899,N_29868,N_29790);
nor UO_1900 (O_1900,N_29159,N_29797);
or UO_1901 (O_1901,N_29078,N_29594);
nor UO_1902 (O_1902,N_29845,N_29910);
nand UO_1903 (O_1903,N_29435,N_29309);
and UO_1904 (O_1904,N_29652,N_29976);
and UO_1905 (O_1905,N_29057,N_29286);
nor UO_1906 (O_1906,N_29835,N_29853);
and UO_1907 (O_1907,N_29775,N_29740);
nand UO_1908 (O_1908,N_29113,N_29389);
or UO_1909 (O_1909,N_29248,N_29461);
or UO_1910 (O_1910,N_29990,N_29760);
or UO_1911 (O_1911,N_29705,N_29840);
or UO_1912 (O_1912,N_29138,N_29148);
or UO_1913 (O_1913,N_28948,N_29271);
nand UO_1914 (O_1914,N_29566,N_29447);
or UO_1915 (O_1915,N_29508,N_28891);
or UO_1916 (O_1916,N_29836,N_29573);
and UO_1917 (O_1917,N_29047,N_28970);
or UO_1918 (O_1918,N_29357,N_28876);
and UO_1919 (O_1919,N_29423,N_29131);
xor UO_1920 (O_1920,N_29268,N_29985);
or UO_1921 (O_1921,N_29641,N_28911);
nor UO_1922 (O_1922,N_28962,N_29020);
nor UO_1923 (O_1923,N_28827,N_28896);
xnor UO_1924 (O_1924,N_29530,N_29796);
and UO_1925 (O_1925,N_29156,N_29746);
nand UO_1926 (O_1926,N_29872,N_29071);
or UO_1927 (O_1927,N_29139,N_29156);
or UO_1928 (O_1928,N_29695,N_29799);
and UO_1929 (O_1929,N_29538,N_29898);
nand UO_1930 (O_1930,N_29464,N_29947);
nand UO_1931 (O_1931,N_29663,N_29656);
and UO_1932 (O_1932,N_29112,N_29583);
xnor UO_1933 (O_1933,N_29214,N_29391);
nand UO_1934 (O_1934,N_29470,N_29347);
xnor UO_1935 (O_1935,N_29942,N_29859);
nand UO_1936 (O_1936,N_28900,N_29651);
and UO_1937 (O_1937,N_29326,N_29845);
or UO_1938 (O_1938,N_29809,N_29377);
xnor UO_1939 (O_1939,N_28832,N_28941);
nor UO_1940 (O_1940,N_29746,N_29388);
nor UO_1941 (O_1941,N_29412,N_29536);
and UO_1942 (O_1942,N_29041,N_29191);
nor UO_1943 (O_1943,N_29798,N_29772);
nand UO_1944 (O_1944,N_28975,N_29935);
nor UO_1945 (O_1945,N_29463,N_29863);
nand UO_1946 (O_1946,N_29736,N_29438);
nand UO_1947 (O_1947,N_29498,N_29785);
xnor UO_1948 (O_1948,N_29783,N_29078);
or UO_1949 (O_1949,N_28843,N_29733);
or UO_1950 (O_1950,N_29282,N_29307);
or UO_1951 (O_1951,N_28881,N_29566);
nor UO_1952 (O_1952,N_29373,N_29667);
xnor UO_1953 (O_1953,N_29803,N_29476);
or UO_1954 (O_1954,N_29526,N_29580);
or UO_1955 (O_1955,N_29021,N_29343);
xor UO_1956 (O_1956,N_28805,N_29502);
or UO_1957 (O_1957,N_29622,N_28815);
xnor UO_1958 (O_1958,N_29420,N_29734);
xor UO_1959 (O_1959,N_29409,N_29477);
and UO_1960 (O_1960,N_29788,N_29829);
nand UO_1961 (O_1961,N_29279,N_28911);
or UO_1962 (O_1962,N_29366,N_29628);
or UO_1963 (O_1963,N_29850,N_28974);
and UO_1964 (O_1964,N_29991,N_29629);
nand UO_1965 (O_1965,N_29347,N_29320);
xnor UO_1966 (O_1966,N_29063,N_29895);
nor UO_1967 (O_1967,N_29663,N_29685);
nor UO_1968 (O_1968,N_29595,N_29291);
xnor UO_1969 (O_1969,N_29372,N_29399);
xnor UO_1970 (O_1970,N_29435,N_29089);
or UO_1971 (O_1971,N_29514,N_29300);
nor UO_1972 (O_1972,N_29768,N_29883);
nand UO_1973 (O_1973,N_29078,N_29533);
or UO_1974 (O_1974,N_29838,N_29335);
xor UO_1975 (O_1975,N_29768,N_28981);
xnor UO_1976 (O_1976,N_29312,N_28909);
xnor UO_1977 (O_1977,N_29188,N_29149);
xor UO_1978 (O_1978,N_29479,N_29379);
nor UO_1979 (O_1979,N_29955,N_29405);
nor UO_1980 (O_1980,N_29688,N_29002);
or UO_1981 (O_1981,N_28805,N_29958);
nor UO_1982 (O_1982,N_29999,N_29365);
nor UO_1983 (O_1983,N_29327,N_29979);
xor UO_1984 (O_1984,N_29457,N_29444);
xor UO_1985 (O_1985,N_29745,N_29497);
xor UO_1986 (O_1986,N_29801,N_28973);
xor UO_1987 (O_1987,N_28917,N_29190);
nand UO_1988 (O_1988,N_29001,N_29536);
or UO_1989 (O_1989,N_28898,N_29995);
or UO_1990 (O_1990,N_29714,N_29627);
xnor UO_1991 (O_1991,N_29609,N_29019);
nor UO_1992 (O_1992,N_29252,N_29675);
xnor UO_1993 (O_1993,N_29346,N_29986);
xor UO_1994 (O_1994,N_29329,N_29066);
nand UO_1995 (O_1995,N_29998,N_29424);
xnor UO_1996 (O_1996,N_29686,N_29079);
xor UO_1997 (O_1997,N_29652,N_29558);
nor UO_1998 (O_1998,N_29191,N_29941);
and UO_1999 (O_1999,N_29924,N_29289);
nand UO_2000 (O_2000,N_28870,N_29688);
and UO_2001 (O_2001,N_28813,N_29354);
xnor UO_2002 (O_2002,N_29886,N_28921);
or UO_2003 (O_2003,N_29122,N_29596);
xor UO_2004 (O_2004,N_28929,N_29574);
nand UO_2005 (O_2005,N_28908,N_29520);
or UO_2006 (O_2006,N_28800,N_29832);
or UO_2007 (O_2007,N_28898,N_29452);
nand UO_2008 (O_2008,N_29262,N_28965);
nand UO_2009 (O_2009,N_29531,N_29291);
and UO_2010 (O_2010,N_28965,N_29571);
xor UO_2011 (O_2011,N_28988,N_29069);
nor UO_2012 (O_2012,N_29767,N_29034);
nand UO_2013 (O_2013,N_29748,N_28898);
nand UO_2014 (O_2014,N_29380,N_29690);
nor UO_2015 (O_2015,N_29773,N_29262);
or UO_2016 (O_2016,N_29541,N_29788);
or UO_2017 (O_2017,N_29799,N_29748);
xor UO_2018 (O_2018,N_29577,N_29530);
nand UO_2019 (O_2019,N_29176,N_28982);
and UO_2020 (O_2020,N_28834,N_29597);
nand UO_2021 (O_2021,N_29976,N_29082);
nand UO_2022 (O_2022,N_29798,N_29694);
xor UO_2023 (O_2023,N_29809,N_29378);
and UO_2024 (O_2024,N_29422,N_28998);
nand UO_2025 (O_2025,N_28970,N_29023);
nand UO_2026 (O_2026,N_29003,N_29223);
nand UO_2027 (O_2027,N_29450,N_29284);
nor UO_2028 (O_2028,N_28922,N_29057);
and UO_2029 (O_2029,N_29325,N_28999);
and UO_2030 (O_2030,N_29596,N_28940);
and UO_2031 (O_2031,N_29756,N_28912);
or UO_2032 (O_2032,N_29092,N_29924);
nor UO_2033 (O_2033,N_29488,N_29862);
or UO_2034 (O_2034,N_29143,N_28804);
nor UO_2035 (O_2035,N_28932,N_29628);
nand UO_2036 (O_2036,N_29559,N_29159);
nand UO_2037 (O_2037,N_28957,N_29190);
nand UO_2038 (O_2038,N_29869,N_29239);
and UO_2039 (O_2039,N_29109,N_29076);
or UO_2040 (O_2040,N_29128,N_29197);
or UO_2041 (O_2041,N_29752,N_29968);
and UO_2042 (O_2042,N_28885,N_29814);
nor UO_2043 (O_2043,N_29214,N_29360);
nor UO_2044 (O_2044,N_28915,N_29115);
xor UO_2045 (O_2045,N_29442,N_29330);
nand UO_2046 (O_2046,N_29849,N_29240);
or UO_2047 (O_2047,N_29541,N_29487);
nand UO_2048 (O_2048,N_29443,N_28841);
xnor UO_2049 (O_2049,N_29254,N_29709);
or UO_2050 (O_2050,N_29130,N_29866);
xnor UO_2051 (O_2051,N_29189,N_29756);
or UO_2052 (O_2052,N_29266,N_29941);
or UO_2053 (O_2053,N_29472,N_29986);
nor UO_2054 (O_2054,N_29008,N_29695);
and UO_2055 (O_2055,N_28858,N_28808);
or UO_2056 (O_2056,N_28935,N_29952);
nor UO_2057 (O_2057,N_29352,N_29505);
nand UO_2058 (O_2058,N_28935,N_28855);
xor UO_2059 (O_2059,N_28900,N_29833);
nand UO_2060 (O_2060,N_29793,N_29526);
xor UO_2061 (O_2061,N_29938,N_29849);
and UO_2062 (O_2062,N_29915,N_29821);
xor UO_2063 (O_2063,N_29739,N_29178);
and UO_2064 (O_2064,N_29332,N_29209);
xnor UO_2065 (O_2065,N_28930,N_29291);
nor UO_2066 (O_2066,N_29273,N_29103);
and UO_2067 (O_2067,N_29139,N_29513);
xor UO_2068 (O_2068,N_29558,N_29189);
and UO_2069 (O_2069,N_29399,N_29910);
nor UO_2070 (O_2070,N_29411,N_29850);
nand UO_2071 (O_2071,N_29764,N_29447);
nand UO_2072 (O_2072,N_28863,N_29545);
xor UO_2073 (O_2073,N_29895,N_29812);
and UO_2074 (O_2074,N_29870,N_28851);
or UO_2075 (O_2075,N_29395,N_29878);
xor UO_2076 (O_2076,N_29246,N_29404);
and UO_2077 (O_2077,N_29427,N_29707);
or UO_2078 (O_2078,N_29897,N_29163);
and UO_2079 (O_2079,N_29280,N_29425);
nor UO_2080 (O_2080,N_29705,N_29592);
and UO_2081 (O_2081,N_28907,N_29709);
and UO_2082 (O_2082,N_28827,N_29239);
nand UO_2083 (O_2083,N_29511,N_29048);
and UO_2084 (O_2084,N_28855,N_28822);
nand UO_2085 (O_2085,N_29195,N_29174);
or UO_2086 (O_2086,N_29702,N_29474);
nor UO_2087 (O_2087,N_29879,N_29702);
or UO_2088 (O_2088,N_29028,N_29228);
nor UO_2089 (O_2089,N_29837,N_29775);
nor UO_2090 (O_2090,N_29092,N_29492);
and UO_2091 (O_2091,N_28855,N_28818);
nand UO_2092 (O_2092,N_29318,N_29037);
and UO_2093 (O_2093,N_29924,N_28867);
nand UO_2094 (O_2094,N_29968,N_28935);
xor UO_2095 (O_2095,N_29234,N_29617);
or UO_2096 (O_2096,N_29323,N_29739);
or UO_2097 (O_2097,N_29094,N_29637);
nand UO_2098 (O_2098,N_29672,N_29068);
nand UO_2099 (O_2099,N_29359,N_29036);
or UO_2100 (O_2100,N_28901,N_29890);
nor UO_2101 (O_2101,N_29846,N_29644);
and UO_2102 (O_2102,N_29187,N_28999);
nand UO_2103 (O_2103,N_29410,N_29729);
xnor UO_2104 (O_2104,N_29336,N_28888);
xnor UO_2105 (O_2105,N_29012,N_29126);
or UO_2106 (O_2106,N_29672,N_29982);
nor UO_2107 (O_2107,N_29149,N_29688);
nor UO_2108 (O_2108,N_29840,N_28890);
nor UO_2109 (O_2109,N_29207,N_29803);
or UO_2110 (O_2110,N_29741,N_29298);
and UO_2111 (O_2111,N_29011,N_29659);
nor UO_2112 (O_2112,N_29571,N_28858);
and UO_2113 (O_2113,N_29804,N_29910);
and UO_2114 (O_2114,N_29985,N_29024);
xor UO_2115 (O_2115,N_29822,N_29121);
nor UO_2116 (O_2116,N_29676,N_29099);
or UO_2117 (O_2117,N_29971,N_29287);
and UO_2118 (O_2118,N_29880,N_29594);
or UO_2119 (O_2119,N_29002,N_29447);
and UO_2120 (O_2120,N_29975,N_29841);
nand UO_2121 (O_2121,N_28906,N_29955);
xnor UO_2122 (O_2122,N_29180,N_28996);
or UO_2123 (O_2123,N_29674,N_29063);
nor UO_2124 (O_2124,N_29001,N_29105);
or UO_2125 (O_2125,N_28892,N_28916);
and UO_2126 (O_2126,N_29844,N_29889);
nand UO_2127 (O_2127,N_29957,N_29150);
xor UO_2128 (O_2128,N_29893,N_29273);
and UO_2129 (O_2129,N_29511,N_29615);
or UO_2130 (O_2130,N_29501,N_29261);
or UO_2131 (O_2131,N_29382,N_29055);
and UO_2132 (O_2132,N_29986,N_29905);
nor UO_2133 (O_2133,N_29975,N_29015);
nor UO_2134 (O_2134,N_29115,N_29059);
nor UO_2135 (O_2135,N_29104,N_29587);
nor UO_2136 (O_2136,N_29245,N_29586);
nand UO_2137 (O_2137,N_29172,N_29260);
nand UO_2138 (O_2138,N_29856,N_29086);
xnor UO_2139 (O_2139,N_28972,N_29850);
xnor UO_2140 (O_2140,N_29931,N_29476);
xnor UO_2141 (O_2141,N_29428,N_29690);
and UO_2142 (O_2142,N_29377,N_29175);
nand UO_2143 (O_2143,N_29401,N_29702);
xnor UO_2144 (O_2144,N_28802,N_29816);
nor UO_2145 (O_2145,N_28893,N_29696);
nor UO_2146 (O_2146,N_29441,N_29071);
and UO_2147 (O_2147,N_29338,N_29895);
nand UO_2148 (O_2148,N_29052,N_29279);
and UO_2149 (O_2149,N_29941,N_28806);
nand UO_2150 (O_2150,N_29708,N_29227);
xor UO_2151 (O_2151,N_29810,N_29575);
nor UO_2152 (O_2152,N_28857,N_29262);
and UO_2153 (O_2153,N_29037,N_29516);
nor UO_2154 (O_2154,N_29847,N_28966);
nor UO_2155 (O_2155,N_29948,N_29430);
nor UO_2156 (O_2156,N_29148,N_29850);
nor UO_2157 (O_2157,N_29820,N_29888);
nand UO_2158 (O_2158,N_29404,N_29055);
or UO_2159 (O_2159,N_29308,N_29738);
nor UO_2160 (O_2160,N_29753,N_29908);
nor UO_2161 (O_2161,N_28964,N_29719);
xnor UO_2162 (O_2162,N_29351,N_29385);
nand UO_2163 (O_2163,N_29143,N_29582);
nor UO_2164 (O_2164,N_29447,N_28901);
nand UO_2165 (O_2165,N_29081,N_29675);
nand UO_2166 (O_2166,N_29898,N_29427);
xnor UO_2167 (O_2167,N_29230,N_28824);
nor UO_2168 (O_2168,N_28954,N_29132);
nand UO_2169 (O_2169,N_28922,N_29385);
or UO_2170 (O_2170,N_29161,N_29330);
or UO_2171 (O_2171,N_28891,N_29140);
nand UO_2172 (O_2172,N_29251,N_29168);
nor UO_2173 (O_2173,N_29581,N_29373);
xor UO_2174 (O_2174,N_29864,N_29832);
or UO_2175 (O_2175,N_29511,N_28821);
nand UO_2176 (O_2176,N_28929,N_29810);
xor UO_2177 (O_2177,N_28993,N_29808);
xnor UO_2178 (O_2178,N_29742,N_29623);
and UO_2179 (O_2179,N_29409,N_29615);
xnor UO_2180 (O_2180,N_29726,N_29097);
and UO_2181 (O_2181,N_29815,N_29733);
and UO_2182 (O_2182,N_29544,N_29119);
and UO_2183 (O_2183,N_29302,N_29165);
nor UO_2184 (O_2184,N_29738,N_29293);
nor UO_2185 (O_2185,N_29590,N_29069);
nand UO_2186 (O_2186,N_29866,N_29255);
xnor UO_2187 (O_2187,N_29567,N_29769);
or UO_2188 (O_2188,N_29627,N_29360);
or UO_2189 (O_2189,N_29792,N_29658);
or UO_2190 (O_2190,N_29804,N_29701);
xor UO_2191 (O_2191,N_29180,N_29230);
and UO_2192 (O_2192,N_29254,N_29836);
and UO_2193 (O_2193,N_29739,N_29772);
nor UO_2194 (O_2194,N_29397,N_29525);
and UO_2195 (O_2195,N_29921,N_29550);
nor UO_2196 (O_2196,N_29188,N_29642);
nor UO_2197 (O_2197,N_29100,N_29382);
and UO_2198 (O_2198,N_29025,N_29061);
and UO_2199 (O_2199,N_29769,N_29880);
and UO_2200 (O_2200,N_29865,N_28928);
or UO_2201 (O_2201,N_29391,N_29475);
xor UO_2202 (O_2202,N_29937,N_29089);
or UO_2203 (O_2203,N_29341,N_29434);
or UO_2204 (O_2204,N_29248,N_28834);
nor UO_2205 (O_2205,N_29224,N_29257);
and UO_2206 (O_2206,N_29869,N_29891);
and UO_2207 (O_2207,N_29183,N_29447);
xor UO_2208 (O_2208,N_29142,N_29699);
or UO_2209 (O_2209,N_29212,N_28839);
and UO_2210 (O_2210,N_29974,N_29210);
nand UO_2211 (O_2211,N_29095,N_29032);
nand UO_2212 (O_2212,N_29710,N_29721);
and UO_2213 (O_2213,N_29484,N_29027);
nand UO_2214 (O_2214,N_29917,N_29812);
nand UO_2215 (O_2215,N_29823,N_29309);
nor UO_2216 (O_2216,N_28982,N_29657);
xnor UO_2217 (O_2217,N_29685,N_28966);
or UO_2218 (O_2218,N_29651,N_29181);
or UO_2219 (O_2219,N_29692,N_29661);
and UO_2220 (O_2220,N_29332,N_29662);
xor UO_2221 (O_2221,N_29193,N_29888);
and UO_2222 (O_2222,N_29726,N_29226);
or UO_2223 (O_2223,N_28869,N_29069);
xor UO_2224 (O_2224,N_29473,N_28861);
xor UO_2225 (O_2225,N_29672,N_29338);
nand UO_2226 (O_2226,N_29504,N_29236);
nand UO_2227 (O_2227,N_28963,N_29690);
nand UO_2228 (O_2228,N_29125,N_29116);
or UO_2229 (O_2229,N_29643,N_28959);
or UO_2230 (O_2230,N_29815,N_29240);
and UO_2231 (O_2231,N_29149,N_28954);
nand UO_2232 (O_2232,N_29323,N_29054);
nor UO_2233 (O_2233,N_29174,N_28872);
and UO_2234 (O_2234,N_29945,N_28990);
xnor UO_2235 (O_2235,N_29791,N_29759);
and UO_2236 (O_2236,N_29681,N_29916);
or UO_2237 (O_2237,N_28923,N_29801);
nand UO_2238 (O_2238,N_29481,N_28818);
or UO_2239 (O_2239,N_29891,N_29048);
or UO_2240 (O_2240,N_29753,N_29377);
and UO_2241 (O_2241,N_29168,N_29327);
xor UO_2242 (O_2242,N_29035,N_29979);
or UO_2243 (O_2243,N_29223,N_29143);
xnor UO_2244 (O_2244,N_29183,N_29346);
or UO_2245 (O_2245,N_29306,N_29493);
or UO_2246 (O_2246,N_29483,N_29204);
nor UO_2247 (O_2247,N_29916,N_29410);
xor UO_2248 (O_2248,N_29715,N_29424);
xor UO_2249 (O_2249,N_29537,N_29012);
or UO_2250 (O_2250,N_29304,N_29334);
and UO_2251 (O_2251,N_29202,N_29329);
xnor UO_2252 (O_2252,N_29372,N_29788);
xor UO_2253 (O_2253,N_28853,N_29684);
xnor UO_2254 (O_2254,N_29236,N_29818);
nor UO_2255 (O_2255,N_29776,N_29702);
or UO_2256 (O_2256,N_28864,N_29522);
and UO_2257 (O_2257,N_29558,N_28933);
nand UO_2258 (O_2258,N_29751,N_29565);
or UO_2259 (O_2259,N_29468,N_29920);
or UO_2260 (O_2260,N_29665,N_29140);
nor UO_2261 (O_2261,N_29548,N_29152);
nand UO_2262 (O_2262,N_29543,N_29720);
xor UO_2263 (O_2263,N_29619,N_29953);
nor UO_2264 (O_2264,N_29419,N_29135);
nor UO_2265 (O_2265,N_29290,N_28921);
or UO_2266 (O_2266,N_28837,N_29301);
or UO_2267 (O_2267,N_29428,N_29455);
nor UO_2268 (O_2268,N_29800,N_29828);
or UO_2269 (O_2269,N_29017,N_29225);
and UO_2270 (O_2270,N_29807,N_28825);
xnor UO_2271 (O_2271,N_29007,N_29191);
xor UO_2272 (O_2272,N_28841,N_28878);
or UO_2273 (O_2273,N_29943,N_29537);
or UO_2274 (O_2274,N_29329,N_29415);
or UO_2275 (O_2275,N_28819,N_29106);
xnor UO_2276 (O_2276,N_29568,N_29929);
and UO_2277 (O_2277,N_29486,N_29451);
nand UO_2278 (O_2278,N_28902,N_28823);
and UO_2279 (O_2279,N_29962,N_29141);
nand UO_2280 (O_2280,N_28934,N_29228);
nor UO_2281 (O_2281,N_29334,N_29644);
nor UO_2282 (O_2282,N_29887,N_29757);
nor UO_2283 (O_2283,N_29747,N_29004);
and UO_2284 (O_2284,N_29016,N_29822);
nand UO_2285 (O_2285,N_29406,N_28913);
xor UO_2286 (O_2286,N_29835,N_29709);
and UO_2287 (O_2287,N_29277,N_29319);
nand UO_2288 (O_2288,N_29108,N_29200);
and UO_2289 (O_2289,N_29408,N_29552);
nand UO_2290 (O_2290,N_29261,N_28846);
nand UO_2291 (O_2291,N_29656,N_29995);
or UO_2292 (O_2292,N_29189,N_29399);
nor UO_2293 (O_2293,N_29154,N_28989);
xor UO_2294 (O_2294,N_29056,N_29163);
and UO_2295 (O_2295,N_29195,N_29864);
nor UO_2296 (O_2296,N_29087,N_29384);
and UO_2297 (O_2297,N_28917,N_29258);
nor UO_2298 (O_2298,N_29290,N_29604);
nand UO_2299 (O_2299,N_29731,N_29156);
or UO_2300 (O_2300,N_29260,N_29068);
nand UO_2301 (O_2301,N_29753,N_29200);
nand UO_2302 (O_2302,N_29119,N_29553);
xnor UO_2303 (O_2303,N_29087,N_28899);
and UO_2304 (O_2304,N_28865,N_29230);
and UO_2305 (O_2305,N_29533,N_29965);
or UO_2306 (O_2306,N_29446,N_29252);
nor UO_2307 (O_2307,N_29632,N_28854);
nor UO_2308 (O_2308,N_29071,N_29488);
nand UO_2309 (O_2309,N_29041,N_29619);
or UO_2310 (O_2310,N_29543,N_29753);
nand UO_2311 (O_2311,N_29219,N_29170);
or UO_2312 (O_2312,N_29046,N_29985);
xor UO_2313 (O_2313,N_29610,N_29288);
nor UO_2314 (O_2314,N_29816,N_29852);
nor UO_2315 (O_2315,N_29794,N_29424);
nand UO_2316 (O_2316,N_29046,N_29884);
and UO_2317 (O_2317,N_29418,N_29720);
nand UO_2318 (O_2318,N_29704,N_28817);
or UO_2319 (O_2319,N_29089,N_29784);
or UO_2320 (O_2320,N_29318,N_29067);
xor UO_2321 (O_2321,N_29790,N_29906);
or UO_2322 (O_2322,N_29987,N_29145);
xnor UO_2323 (O_2323,N_29390,N_29851);
xor UO_2324 (O_2324,N_29548,N_29175);
and UO_2325 (O_2325,N_29659,N_29499);
nand UO_2326 (O_2326,N_29690,N_29631);
nand UO_2327 (O_2327,N_29018,N_29744);
and UO_2328 (O_2328,N_29410,N_29828);
nand UO_2329 (O_2329,N_29324,N_29867);
nor UO_2330 (O_2330,N_29414,N_29268);
nor UO_2331 (O_2331,N_28833,N_29437);
or UO_2332 (O_2332,N_29941,N_29507);
nand UO_2333 (O_2333,N_29355,N_29944);
xnor UO_2334 (O_2334,N_28944,N_29988);
and UO_2335 (O_2335,N_29279,N_29587);
nand UO_2336 (O_2336,N_29769,N_29785);
nor UO_2337 (O_2337,N_29328,N_29939);
nor UO_2338 (O_2338,N_29572,N_29923);
xor UO_2339 (O_2339,N_29483,N_29655);
nand UO_2340 (O_2340,N_29741,N_29780);
nand UO_2341 (O_2341,N_29059,N_29453);
or UO_2342 (O_2342,N_29807,N_29806);
or UO_2343 (O_2343,N_29176,N_29590);
or UO_2344 (O_2344,N_29597,N_29211);
and UO_2345 (O_2345,N_29163,N_29099);
and UO_2346 (O_2346,N_29331,N_29720);
nand UO_2347 (O_2347,N_29334,N_29467);
and UO_2348 (O_2348,N_29331,N_29141);
or UO_2349 (O_2349,N_29291,N_29179);
nand UO_2350 (O_2350,N_29838,N_29332);
and UO_2351 (O_2351,N_29486,N_29864);
or UO_2352 (O_2352,N_29707,N_29287);
nor UO_2353 (O_2353,N_29299,N_29594);
nand UO_2354 (O_2354,N_28823,N_29478);
nor UO_2355 (O_2355,N_29740,N_29627);
and UO_2356 (O_2356,N_28873,N_29291);
nand UO_2357 (O_2357,N_29934,N_29054);
and UO_2358 (O_2358,N_29864,N_29330);
nor UO_2359 (O_2359,N_29855,N_29106);
or UO_2360 (O_2360,N_29781,N_29652);
and UO_2361 (O_2361,N_29906,N_28941);
or UO_2362 (O_2362,N_28820,N_29621);
nor UO_2363 (O_2363,N_28961,N_29463);
or UO_2364 (O_2364,N_29287,N_28817);
or UO_2365 (O_2365,N_29338,N_29211);
or UO_2366 (O_2366,N_29339,N_29394);
nand UO_2367 (O_2367,N_29473,N_29144);
and UO_2368 (O_2368,N_29171,N_28817);
nor UO_2369 (O_2369,N_29851,N_29932);
and UO_2370 (O_2370,N_29451,N_29591);
nand UO_2371 (O_2371,N_29504,N_29834);
nand UO_2372 (O_2372,N_29443,N_28903);
or UO_2373 (O_2373,N_29882,N_29482);
nor UO_2374 (O_2374,N_29496,N_29386);
nor UO_2375 (O_2375,N_28905,N_29432);
xor UO_2376 (O_2376,N_29267,N_29438);
and UO_2377 (O_2377,N_29825,N_29608);
and UO_2378 (O_2378,N_29509,N_29040);
nor UO_2379 (O_2379,N_28836,N_29376);
or UO_2380 (O_2380,N_29116,N_28961);
and UO_2381 (O_2381,N_29019,N_29338);
nor UO_2382 (O_2382,N_29657,N_28856);
xnor UO_2383 (O_2383,N_29499,N_29892);
xor UO_2384 (O_2384,N_29435,N_28834);
nor UO_2385 (O_2385,N_29196,N_29567);
or UO_2386 (O_2386,N_29765,N_29028);
xnor UO_2387 (O_2387,N_29999,N_28900);
nor UO_2388 (O_2388,N_29661,N_29131);
xor UO_2389 (O_2389,N_28804,N_29407);
and UO_2390 (O_2390,N_29528,N_29153);
nand UO_2391 (O_2391,N_28855,N_29449);
and UO_2392 (O_2392,N_29433,N_29175);
nor UO_2393 (O_2393,N_28897,N_29239);
nand UO_2394 (O_2394,N_29791,N_29747);
xor UO_2395 (O_2395,N_29880,N_29331);
nor UO_2396 (O_2396,N_28810,N_29393);
xnor UO_2397 (O_2397,N_29580,N_29642);
or UO_2398 (O_2398,N_29692,N_29058);
xor UO_2399 (O_2399,N_29347,N_29264);
or UO_2400 (O_2400,N_29059,N_29077);
xor UO_2401 (O_2401,N_29714,N_28807);
or UO_2402 (O_2402,N_28874,N_29442);
or UO_2403 (O_2403,N_29423,N_29243);
or UO_2404 (O_2404,N_28845,N_29387);
nor UO_2405 (O_2405,N_28894,N_28991);
or UO_2406 (O_2406,N_29803,N_29740);
and UO_2407 (O_2407,N_29356,N_28968);
or UO_2408 (O_2408,N_29173,N_29119);
nand UO_2409 (O_2409,N_29942,N_29634);
nor UO_2410 (O_2410,N_28875,N_29072);
xnor UO_2411 (O_2411,N_29117,N_29965);
or UO_2412 (O_2412,N_28934,N_29018);
nand UO_2413 (O_2413,N_28844,N_28969);
nand UO_2414 (O_2414,N_29803,N_29273);
xnor UO_2415 (O_2415,N_29864,N_29796);
and UO_2416 (O_2416,N_28913,N_29191);
xnor UO_2417 (O_2417,N_29416,N_29870);
xor UO_2418 (O_2418,N_28839,N_29293);
and UO_2419 (O_2419,N_29619,N_29606);
xor UO_2420 (O_2420,N_29797,N_29552);
nor UO_2421 (O_2421,N_28885,N_29965);
or UO_2422 (O_2422,N_29195,N_29300);
xor UO_2423 (O_2423,N_29277,N_29665);
nor UO_2424 (O_2424,N_29306,N_29482);
nand UO_2425 (O_2425,N_29248,N_28804);
xnor UO_2426 (O_2426,N_29809,N_29465);
xor UO_2427 (O_2427,N_29833,N_29007);
xor UO_2428 (O_2428,N_29283,N_29217);
and UO_2429 (O_2429,N_29005,N_29241);
nand UO_2430 (O_2430,N_29408,N_29132);
and UO_2431 (O_2431,N_29146,N_29036);
or UO_2432 (O_2432,N_29018,N_29554);
and UO_2433 (O_2433,N_29030,N_28987);
nor UO_2434 (O_2434,N_29672,N_29992);
nand UO_2435 (O_2435,N_28983,N_29858);
nor UO_2436 (O_2436,N_29670,N_29654);
xnor UO_2437 (O_2437,N_29752,N_29001);
or UO_2438 (O_2438,N_29288,N_29471);
or UO_2439 (O_2439,N_29332,N_29907);
nor UO_2440 (O_2440,N_29916,N_29780);
nand UO_2441 (O_2441,N_29873,N_29717);
nor UO_2442 (O_2442,N_29682,N_29093);
xor UO_2443 (O_2443,N_29084,N_29349);
nor UO_2444 (O_2444,N_29854,N_28902);
nand UO_2445 (O_2445,N_29893,N_29834);
or UO_2446 (O_2446,N_29291,N_29120);
nor UO_2447 (O_2447,N_29147,N_29023);
and UO_2448 (O_2448,N_28931,N_29355);
xnor UO_2449 (O_2449,N_28898,N_29707);
or UO_2450 (O_2450,N_29379,N_29949);
nor UO_2451 (O_2451,N_29355,N_29629);
nor UO_2452 (O_2452,N_29748,N_29766);
nand UO_2453 (O_2453,N_29305,N_29958);
or UO_2454 (O_2454,N_28824,N_29010);
nand UO_2455 (O_2455,N_29591,N_29037);
or UO_2456 (O_2456,N_29505,N_28966);
or UO_2457 (O_2457,N_28896,N_29160);
or UO_2458 (O_2458,N_29840,N_29283);
xnor UO_2459 (O_2459,N_29803,N_29589);
nand UO_2460 (O_2460,N_29440,N_29070);
nor UO_2461 (O_2461,N_29777,N_29743);
nor UO_2462 (O_2462,N_29791,N_29704);
nand UO_2463 (O_2463,N_29602,N_29397);
and UO_2464 (O_2464,N_29776,N_29647);
nand UO_2465 (O_2465,N_29256,N_29028);
xnor UO_2466 (O_2466,N_29954,N_28904);
nand UO_2467 (O_2467,N_28802,N_29043);
nand UO_2468 (O_2468,N_29415,N_29973);
and UO_2469 (O_2469,N_29181,N_29459);
xor UO_2470 (O_2470,N_29483,N_29722);
nor UO_2471 (O_2471,N_29231,N_29304);
xnor UO_2472 (O_2472,N_29633,N_28808);
xor UO_2473 (O_2473,N_29441,N_29299);
nand UO_2474 (O_2474,N_29623,N_29833);
xor UO_2475 (O_2475,N_28811,N_29052);
nor UO_2476 (O_2476,N_29148,N_29090);
nor UO_2477 (O_2477,N_29351,N_29133);
and UO_2478 (O_2478,N_29033,N_29675);
nor UO_2479 (O_2479,N_29499,N_29963);
and UO_2480 (O_2480,N_29631,N_29299);
xor UO_2481 (O_2481,N_29373,N_28951);
or UO_2482 (O_2482,N_29986,N_29945);
or UO_2483 (O_2483,N_29159,N_29380);
xnor UO_2484 (O_2484,N_29898,N_29076);
and UO_2485 (O_2485,N_29490,N_29489);
and UO_2486 (O_2486,N_29880,N_28966);
or UO_2487 (O_2487,N_29874,N_29215);
and UO_2488 (O_2488,N_29281,N_29771);
and UO_2489 (O_2489,N_29326,N_29964);
nor UO_2490 (O_2490,N_29222,N_28908);
xor UO_2491 (O_2491,N_29552,N_29777);
xnor UO_2492 (O_2492,N_29538,N_29372);
nor UO_2493 (O_2493,N_28819,N_29227);
or UO_2494 (O_2494,N_29608,N_29236);
nand UO_2495 (O_2495,N_29405,N_29473);
nand UO_2496 (O_2496,N_29402,N_29798);
and UO_2497 (O_2497,N_29701,N_28818);
nor UO_2498 (O_2498,N_28939,N_28944);
nor UO_2499 (O_2499,N_29581,N_29068);
or UO_2500 (O_2500,N_29892,N_29125);
nor UO_2501 (O_2501,N_29257,N_29204);
nor UO_2502 (O_2502,N_29190,N_29625);
xnor UO_2503 (O_2503,N_29157,N_29345);
xnor UO_2504 (O_2504,N_29702,N_29996);
or UO_2505 (O_2505,N_29180,N_29878);
nor UO_2506 (O_2506,N_29783,N_29147);
or UO_2507 (O_2507,N_29256,N_29616);
or UO_2508 (O_2508,N_29318,N_29308);
nand UO_2509 (O_2509,N_29525,N_29120);
and UO_2510 (O_2510,N_29693,N_28843);
or UO_2511 (O_2511,N_29622,N_29616);
nand UO_2512 (O_2512,N_28932,N_29664);
xnor UO_2513 (O_2513,N_29939,N_29384);
or UO_2514 (O_2514,N_29327,N_29005);
nand UO_2515 (O_2515,N_29429,N_28996);
or UO_2516 (O_2516,N_28880,N_29315);
nand UO_2517 (O_2517,N_29671,N_29826);
and UO_2518 (O_2518,N_29228,N_29575);
xor UO_2519 (O_2519,N_29861,N_29238);
and UO_2520 (O_2520,N_29158,N_29806);
nand UO_2521 (O_2521,N_29566,N_29799);
xor UO_2522 (O_2522,N_29447,N_29379);
and UO_2523 (O_2523,N_29337,N_28922);
and UO_2524 (O_2524,N_29992,N_29432);
or UO_2525 (O_2525,N_29950,N_29070);
nand UO_2526 (O_2526,N_29006,N_29182);
xnor UO_2527 (O_2527,N_29382,N_29314);
nand UO_2528 (O_2528,N_29701,N_29435);
or UO_2529 (O_2529,N_29311,N_28834);
and UO_2530 (O_2530,N_29398,N_29925);
and UO_2531 (O_2531,N_29760,N_29245);
nand UO_2532 (O_2532,N_29984,N_29693);
nor UO_2533 (O_2533,N_29052,N_29111);
and UO_2534 (O_2534,N_29455,N_29495);
nand UO_2535 (O_2535,N_29164,N_28884);
or UO_2536 (O_2536,N_29979,N_29804);
xor UO_2537 (O_2537,N_29747,N_29456);
nand UO_2538 (O_2538,N_28928,N_29846);
xnor UO_2539 (O_2539,N_29775,N_29557);
nor UO_2540 (O_2540,N_29829,N_29790);
or UO_2541 (O_2541,N_28843,N_29388);
nand UO_2542 (O_2542,N_29588,N_29818);
nand UO_2543 (O_2543,N_29751,N_29875);
nand UO_2544 (O_2544,N_29479,N_29994);
nor UO_2545 (O_2545,N_29238,N_28985);
nand UO_2546 (O_2546,N_29240,N_29185);
and UO_2547 (O_2547,N_29390,N_29138);
and UO_2548 (O_2548,N_29338,N_29566);
nor UO_2549 (O_2549,N_29526,N_28821);
xor UO_2550 (O_2550,N_29391,N_29702);
xor UO_2551 (O_2551,N_28935,N_29657);
nor UO_2552 (O_2552,N_28900,N_28925);
and UO_2553 (O_2553,N_29046,N_28810);
xnor UO_2554 (O_2554,N_29814,N_29654);
or UO_2555 (O_2555,N_29309,N_29991);
xnor UO_2556 (O_2556,N_29534,N_29673);
or UO_2557 (O_2557,N_29642,N_28996);
and UO_2558 (O_2558,N_29762,N_29630);
or UO_2559 (O_2559,N_29619,N_29989);
and UO_2560 (O_2560,N_28874,N_29121);
and UO_2561 (O_2561,N_29908,N_29204);
nor UO_2562 (O_2562,N_29661,N_29867);
nor UO_2563 (O_2563,N_28870,N_28959);
and UO_2564 (O_2564,N_29169,N_29301);
nor UO_2565 (O_2565,N_29636,N_29403);
or UO_2566 (O_2566,N_29941,N_29206);
or UO_2567 (O_2567,N_29055,N_29075);
nand UO_2568 (O_2568,N_29350,N_29746);
and UO_2569 (O_2569,N_29910,N_29926);
xnor UO_2570 (O_2570,N_28886,N_29882);
nor UO_2571 (O_2571,N_29076,N_29399);
and UO_2572 (O_2572,N_29979,N_29903);
nand UO_2573 (O_2573,N_29880,N_29996);
nand UO_2574 (O_2574,N_28933,N_29365);
nor UO_2575 (O_2575,N_29597,N_29136);
xnor UO_2576 (O_2576,N_28818,N_29733);
or UO_2577 (O_2577,N_29576,N_29428);
nand UO_2578 (O_2578,N_29599,N_29307);
nor UO_2579 (O_2579,N_29577,N_29056);
or UO_2580 (O_2580,N_29880,N_29073);
nand UO_2581 (O_2581,N_29879,N_29942);
nand UO_2582 (O_2582,N_28806,N_29332);
or UO_2583 (O_2583,N_29039,N_29407);
nand UO_2584 (O_2584,N_29247,N_29926);
and UO_2585 (O_2585,N_29480,N_29770);
and UO_2586 (O_2586,N_29558,N_28946);
or UO_2587 (O_2587,N_29773,N_29847);
or UO_2588 (O_2588,N_29320,N_29262);
nand UO_2589 (O_2589,N_29900,N_29891);
or UO_2590 (O_2590,N_28939,N_28911);
and UO_2591 (O_2591,N_28824,N_29087);
and UO_2592 (O_2592,N_29482,N_29957);
nor UO_2593 (O_2593,N_29166,N_29484);
xnor UO_2594 (O_2594,N_29413,N_29880);
nand UO_2595 (O_2595,N_29325,N_29344);
and UO_2596 (O_2596,N_29535,N_29232);
nor UO_2597 (O_2597,N_28903,N_29029);
or UO_2598 (O_2598,N_29151,N_29029);
nor UO_2599 (O_2599,N_29120,N_29077);
or UO_2600 (O_2600,N_29890,N_29746);
and UO_2601 (O_2601,N_29768,N_29559);
nand UO_2602 (O_2602,N_29643,N_28893);
nand UO_2603 (O_2603,N_29975,N_29939);
xor UO_2604 (O_2604,N_29416,N_28909);
nand UO_2605 (O_2605,N_29308,N_29268);
and UO_2606 (O_2606,N_29427,N_29597);
nand UO_2607 (O_2607,N_28945,N_29644);
xor UO_2608 (O_2608,N_29584,N_29599);
or UO_2609 (O_2609,N_29414,N_29662);
xnor UO_2610 (O_2610,N_29780,N_29181);
nand UO_2611 (O_2611,N_29857,N_28960);
nand UO_2612 (O_2612,N_29837,N_28939);
and UO_2613 (O_2613,N_29691,N_29569);
and UO_2614 (O_2614,N_29127,N_29448);
and UO_2615 (O_2615,N_29268,N_29249);
nor UO_2616 (O_2616,N_29024,N_29964);
and UO_2617 (O_2617,N_29890,N_29836);
and UO_2618 (O_2618,N_29650,N_29154);
and UO_2619 (O_2619,N_29804,N_29316);
nand UO_2620 (O_2620,N_29774,N_28912);
nor UO_2621 (O_2621,N_29518,N_28837);
or UO_2622 (O_2622,N_28856,N_28977);
and UO_2623 (O_2623,N_29900,N_29117);
nor UO_2624 (O_2624,N_29632,N_29752);
or UO_2625 (O_2625,N_28977,N_29109);
nor UO_2626 (O_2626,N_29001,N_29568);
xor UO_2627 (O_2627,N_29079,N_29560);
xnor UO_2628 (O_2628,N_29015,N_29786);
and UO_2629 (O_2629,N_29888,N_29953);
and UO_2630 (O_2630,N_29624,N_28871);
or UO_2631 (O_2631,N_29549,N_29433);
xor UO_2632 (O_2632,N_29713,N_29937);
nand UO_2633 (O_2633,N_29478,N_29837);
and UO_2634 (O_2634,N_28968,N_29461);
nand UO_2635 (O_2635,N_28862,N_29623);
nor UO_2636 (O_2636,N_29248,N_29735);
nand UO_2637 (O_2637,N_29668,N_29600);
or UO_2638 (O_2638,N_29061,N_28961);
nand UO_2639 (O_2639,N_29282,N_29592);
or UO_2640 (O_2640,N_29618,N_29829);
nor UO_2641 (O_2641,N_29115,N_28923);
nor UO_2642 (O_2642,N_29898,N_29428);
or UO_2643 (O_2643,N_29073,N_29429);
and UO_2644 (O_2644,N_28930,N_29393);
or UO_2645 (O_2645,N_29900,N_29582);
xnor UO_2646 (O_2646,N_29252,N_29984);
or UO_2647 (O_2647,N_29461,N_29399);
nand UO_2648 (O_2648,N_29114,N_29130);
or UO_2649 (O_2649,N_29628,N_29454);
or UO_2650 (O_2650,N_29740,N_29598);
xor UO_2651 (O_2651,N_29620,N_29272);
and UO_2652 (O_2652,N_29811,N_29151);
or UO_2653 (O_2653,N_29253,N_29010);
and UO_2654 (O_2654,N_29162,N_29191);
nor UO_2655 (O_2655,N_29075,N_29382);
nor UO_2656 (O_2656,N_29471,N_29464);
nand UO_2657 (O_2657,N_29531,N_28886);
nand UO_2658 (O_2658,N_29452,N_29609);
nor UO_2659 (O_2659,N_29590,N_29071);
nand UO_2660 (O_2660,N_29411,N_29225);
nand UO_2661 (O_2661,N_28866,N_29032);
and UO_2662 (O_2662,N_29668,N_29697);
and UO_2663 (O_2663,N_28935,N_29123);
nor UO_2664 (O_2664,N_29700,N_29977);
or UO_2665 (O_2665,N_29811,N_29488);
xnor UO_2666 (O_2666,N_29578,N_29390);
and UO_2667 (O_2667,N_29857,N_29184);
and UO_2668 (O_2668,N_29734,N_29672);
nand UO_2669 (O_2669,N_29681,N_29061);
and UO_2670 (O_2670,N_29228,N_29003);
xor UO_2671 (O_2671,N_29142,N_29550);
xor UO_2672 (O_2672,N_29125,N_29334);
or UO_2673 (O_2673,N_29968,N_29678);
nand UO_2674 (O_2674,N_29942,N_28808);
and UO_2675 (O_2675,N_29938,N_28878);
nor UO_2676 (O_2676,N_29102,N_29615);
nand UO_2677 (O_2677,N_29326,N_29130);
or UO_2678 (O_2678,N_28945,N_29277);
nor UO_2679 (O_2679,N_29552,N_28844);
or UO_2680 (O_2680,N_28892,N_29063);
nand UO_2681 (O_2681,N_29106,N_29254);
xnor UO_2682 (O_2682,N_28889,N_29456);
nor UO_2683 (O_2683,N_28871,N_29232);
nand UO_2684 (O_2684,N_29332,N_29570);
nor UO_2685 (O_2685,N_29078,N_28999);
or UO_2686 (O_2686,N_29323,N_29840);
nor UO_2687 (O_2687,N_29465,N_29348);
and UO_2688 (O_2688,N_29126,N_29914);
nor UO_2689 (O_2689,N_29309,N_29700);
and UO_2690 (O_2690,N_29658,N_29237);
or UO_2691 (O_2691,N_28870,N_29928);
and UO_2692 (O_2692,N_29969,N_29436);
or UO_2693 (O_2693,N_29275,N_29735);
and UO_2694 (O_2694,N_29591,N_28800);
or UO_2695 (O_2695,N_28972,N_28968);
xor UO_2696 (O_2696,N_29255,N_29150);
and UO_2697 (O_2697,N_28845,N_28958);
nor UO_2698 (O_2698,N_28862,N_29059);
nand UO_2699 (O_2699,N_29081,N_29554);
nor UO_2700 (O_2700,N_29327,N_29512);
or UO_2701 (O_2701,N_29012,N_29918);
nor UO_2702 (O_2702,N_28906,N_29461);
nor UO_2703 (O_2703,N_28852,N_29665);
nor UO_2704 (O_2704,N_28805,N_29058);
nand UO_2705 (O_2705,N_29160,N_29386);
xor UO_2706 (O_2706,N_29191,N_29193);
and UO_2707 (O_2707,N_29634,N_29722);
nand UO_2708 (O_2708,N_29628,N_28924);
nor UO_2709 (O_2709,N_28972,N_29376);
and UO_2710 (O_2710,N_29545,N_29148);
and UO_2711 (O_2711,N_29163,N_29190);
xor UO_2712 (O_2712,N_29677,N_29751);
and UO_2713 (O_2713,N_29352,N_29733);
xor UO_2714 (O_2714,N_29291,N_29294);
nor UO_2715 (O_2715,N_29049,N_29295);
nand UO_2716 (O_2716,N_29418,N_29637);
xor UO_2717 (O_2717,N_29125,N_28901);
xnor UO_2718 (O_2718,N_28996,N_29147);
nor UO_2719 (O_2719,N_29321,N_29863);
or UO_2720 (O_2720,N_29403,N_29071);
xor UO_2721 (O_2721,N_29090,N_29972);
or UO_2722 (O_2722,N_29911,N_29809);
xor UO_2723 (O_2723,N_29812,N_29182);
xnor UO_2724 (O_2724,N_29460,N_29511);
and UO_2725 (O_2725,N_28808,N_29401);
nor UO_2726 (O_2726,N_28877,N_29584);
and UO_2727 (O_2727,N_29724,N_29642);
and UO_2728 (O_2728,N_29557,N_28916);
xor UO_2729 (O_2729,N_29542,N_29523);
and UO_2730 (O_2730,N_29743,N_29345);
nand UO_2731 (O_2731,N_28907,N_29098);
xnor UO_2732 (O_2732,N_29625,N_29545);
nand UO_2733 (O_2733,N_29358,N_29832);
or UO_2734 (O_2734,N_29901,N_29944);
xnor UO_2735 (O_2735,N_29730,N_29311);
nand UO_2736 (O_2736,N_29307,N_29220);
xor UO_2737 (O_2737,N_29773,N_29430);
and UO_2738 (O_2738,N_29994,N_29417);
xor UO_2739 (O_2739,N_28990,N_29761);
xor UO_2740 (O_2740,N_29229,N_29142);
or UO_2741 (O_2741,N_29907,N_28806);
nor UO_2742 (O_2742,N_29797,N_29874);
nor UO_2743 (O_2743,N_29033,N_29749);
nand UO_2744 (O_2744,N_29386,N_29460);
and UO_2745 (O_2745,N_29938,N_28950);
xnor UO_2746 (O_2746,N_28986,N_29889);
and UO_2747 (O_2747,N_29957,N_29147);
and UO_2748 (O_2748,N_29667,N_29754);
or UO_2749 (O_2749,N_28961,N_29706);
nor UO_2750 (O_2750,N_29318,N_29880);
nand UO_2751 (O_2751,N_29711,N_29144);
or UO_2752 (O_2752,N_29738,N_29829);
or UO_2753 (O_2753,N_29730,N_29624);
or UO_2754 (O_2754,N_29695,N_29915);
xnor UO_2755 (O_2755,N_29606,N_29969);
xor UO_2756 (O_2756,N_29840,N_29122);
nand UO_2757 (O_2757,N_29545,N_29598);
or UO_2758 (O_2758,N_29063,N_29085);
nor UO_2759 (O_2759,N_29186,N_29229);
or UO_2760 (O_2760,N_29210,N_29825);
or UO_2761 (O_2761,N_29836,N_29280);
nor UO_2762 (O_2762,N_29513,N_29752);
or UO_2763 (O_2763,N_28993,N_29478);
nand UO_2764 (O_2764,N_29597,N_29011);
nand UO_2765 (O_2765,N_29026,N_29599);
xnor UO_2766 (O_2766,N_29952,N_29236);
and UO_2767 (O_2767,N_29492,N_29523);
and UO_2768 (O_2768,N_29598,N_29208);
or UO_2769 (O_2769,N_29888,N_29495);
xor UO_2770 (O_2770,N_29226,N_28852);
nand UO_2771 (O_2771,N_29032,N_28995);
and UO_2772 (O_2772,N_29703,N_29173);
or UO_2773 (O_2773,N_29307,N_29005);
xnor UO_2774 (O_2774,N_29186,N_28984);
nor UO_2775 (O_2775,N_29322,N_29584);
nand UO_2776 (O_2776,N_29838,N_29010);
and UO_2777 (O_2777,N_29035,N_29522);
xor UO_2778 (O_2778,N_29498,N_29351);
xnor UO_2779 (O_2779,N_29538,N_28805);
nand UO_2780 (O_2780,N_29363,N_29101);
or UO_2781 (O_2781,N_29785,N_29351);
and UO_2782 (O_2782,N_29369,N_29359);
nor UO_2783 (O_2783,N_29369,N_29751);
and UO_2784 (O_2784,N_29797,N_29377);
xor UO_2785 (O_2785,N_29812,N_29599);
nand UO_2786 (O_2786,N_29659,N_29440);
and UO_2787 (O_2787,N_29956,N_29284);
and UO_2788 (O_2788,N_29337,N_29548);
and UO_2789 (O_2789,N_29491,N_29176);
nor UO_2790 (O_2790,N_29227,N_29262);
xnor UO_2791 (O_2791,N_29191,N_29636);
xor UO_2792 (O_2792,N_28987,N_29643);
or UO_2793 (O_2793,N_28839,N_29445);
nor UO_2794 (O_2794,N_29965,N_29244);
or UO_2795 (O_2795,N_28979,N_29782);
and UO_2796 (O_2796,N_28872,N_28825);
nand UO_2797 (O_2797,N_29820,N_29184);
or UO_2798 (O_2798,N_29646,N_29290);
nand UO_2799 (O_2799,N_29620,N_29128);
nor UO_2800 (O_2800,N_29357,N_29771);
or UO_2801 (O_2801,N_29595,N_29666);
and UO_2802 (O_2802,N_28997,N_29090);
nand UO_2803 (O_2803,N_29712,N_29571);
nand UO_2804 (O_2804,N_29655,N_29490);
or UO_2805 (O_2805,N_29560,N_29347);
nand UO_2806 (O_2806,N_28891,N_29039);
and UO_2807 (O_2807,N_29187,N_29044);
xor UO_2808 (O_2808,N_29425,N_29341);
nor UO_2809 (O_2809,N_29921,N_29355);
xor UO_2810 (O_2810,N_29787,N_29191);
nand UO_2811 (O_2811,N_29656,N_29831);
nand UO_2812 (O_2812,N_29276,N_29338);
xor UO_2813 (O_2813,N_29085,N_29024);
xor UO_2814 (O_2814,N_29877,N_29538);
nand UO_2815 (O_2815,N_28920,N_29520);
or UO_2816 (O_2816,N_29662,N_28909);
xnor UO_2817 (O_2817,N_29533,N_29297);
nand UO_2818 (O_2818,N_29324,N_28970);
xnor UO_2819 (O_2819,N_29473,N_28823);
nor UO_2820 (O_2820,N_29159,N_29743);
nand UO_2821 (O_2821,N_29676,N_29520);
and UO_2822 (O_2822,N_29726,N_28884);
nand UO_2823 (O_2823,N_29939,N_29738);
nor UO_2824 (O_2824,N_29929,N_29808);
xnor UO_2825 (O_2825,N_29876,N_29314);
and UO_2826 (O_2826,N_29998,N_29752);
nor UO_2827 (O_2827,N_29707,N_29682);
nor UO_2828 (O_2828,N_29454,N_29248);
or UO_2829 (O_2829,N_29049,N_28863);
and UO_2830 (O_2830,N_29088,N_29108);
xnor UO_2831 (O_2831,N_29277,N_28835);
xnor UO_2832 (O_2832,N_29945,N_29211);
xor UO_2833 (O_2833,N_28822,N_29199);
and UO_2834 (O_2834,N_28960,N_29943);
nand UO_2835 (O_2835,N_29402,N_29914);
nor UO_2836 (O_2836,N_29586,N_29708);
or UO_2837 (O_2837,N_29906,N_29396);
or UO_2838 (O_2838,N_29759,N_29472);
nor UO_2839 (O_2839,N_29552,N_29004);
or UO_2840 (O_2840,N_28888,N_29002);
xnor UO_2841 (O_2841,N_29306,N_29365);
xnor UO_2842 (O_2842,N_29715,N_29605);
nand UO_2843 (O_2843,N_28853,N_29979);
or UO_2844 (O_2844,N_28959,N_29735);
and UO_2845 (O_2845,N_29322,N_29739);
and UO_2846 (O_2846,N_29043,N_29818);
and UO_2847 (O_2847,N_29070,N_28955);
and UO_2848 (O_2848,N_29572,N_28973);
and UO_2849 (O_2849,N_29680,N_28943);
xor UO_2850 (O_2850,N_29680,N_29476);
nand UO_2851 (O_2851,N_29696,N_28995);
and UO_2852 (O_2852,N_29664,N_29265);
nor UO_2853 (O_2853,N_29740,N_29907);
or UO_2854 (O_2854,N_29663,N_29001);
or UO_2855 (O_2855,N_29863,N_29656);
nor UO_2856 (O_2856,N_29486,N_29354);
or UO_2857 (O_2857,N_28824,N_29418);
nand UO_2858 (O_2858,N_29901,N_29614);
nand UO_2859 (O_2859,N_29672,N_28924);
and UO_2860 (O_2860,N_29388,N_29325);
xnor UO_2861 (O_2861,N_29658,N_29890);
nand UO_2862 (O_2862,N_29926,N_28801);
and UO_2863 (O_2863,N_29100,N_29693);
nor UO_2864 (O_2864,N_29960,N_29008);
nand UO_2865 (O_2865,N_29957,N_29350);
or UO_2866 (O_2866,N_28983,N_29880);
nor UO_2867 (O_2867,N_29807,N_29686);
and UO_2868 (O_2868,N_29921,N_29532);
xor UO_2869 (O_2869,N_28821,N_29888);
nand UO_2870 (O_2870,N_29781,N_29122);
and UO_2871 (O_2871,N_29907,N_29405);
xor UO_2872 (O_2872,N_28844,N_29434);
nor UO_2873 (O_2873,N_29794,N_29934);
and UO_2874 (O_2874,N_29969,N_29320);
and UO_2875 (O_2875,N_28981,N_29107);
and UO_2876 (O_2876,N_29658,N_29720);
and UO_2877 (O_2877,N_29571,N_29240);
or UO_2878 (O_2878,N_29595,N_29039);
and UO_2879 (O_2879,N_28948,N_29061);
nand UO_2880 (O_2880,N_29073,N_29368);
and UO_2881 (O_2881,N_29185,N_29679);
and UO_2882 (O_2882,N_28834,N_28929);
nand UO_2883 (O_2883,N_29185,N_28827);
xnor UO_2884 (O_2884,N_29675,N_29355);
xor UO_2885 (O_2885,N_29902,N_29851);
nand UO_2886 (O_2886,N_29455,N_28880);
nor UO_2887 (O_2887,N_29451,N_29013);
xor UO_2888 (O_2888,N_28816,N_28944);
nand UO_2889 (O_2889,N_29279,N_29019);
or UO_2890 (O_2890,N_29313,N_28997);
nand UO_2891 (O_2891,N_29580,N_29194);
or UO_2892 (O_2892,N_28835,N_29756);
and UO_2893 (O_2893,N_29340,N_28817);
nor UO_2894 (O_2894,N_28942,N_29990);
or UO_2895 (O_2895,N_29729,N_29508);
nand UO_2896 (O_2896,N_29717,N_29524);
nand UO_2897 (O_2897,N_29339,N_28849);
xor UO_2898 (O_2898,N_28979,N_28877);
nor UO_2899 (O_2899,N_29716,N_29530);
nand UO_2900 (O_2900,N_29617,N_29968);
or UO_2901 (O_2901,N_29112,N_29779);
xor UO_2902 (O_2902,N_28999,N_28838);
nor UO_2903 (O_2903,N_29168,N_29733);
and UO_2904 (O_2904,N_28855,N_29762);
xor UO_2905 (O_2905,N_29604,N_29227);
and UO_2906 (O_2906,N_29605,N_29839);
nor UO_2907 (O_2907,N_29103,N_29458);
nand UO_2908 (O_2908,N_29508,N_29142);
xor UO_2909 (O_2909,N_29644,N_29642);
or UO_2910 (O_2910,N_28828,N_29776);
or UO_2911 (O_2911,N_29032,N_29475);
xnor UO_2912 (O_2912,N_29243,N_29740);
nand UO_2913 (O_2913,N_29021,N_29366);
or UO_2914 (O_2914,N_29729,N_29453);
or UO_2915 (O_2915,N_29987,N_29690);
nor UO_2916 (O_2916,N_29024,N_29038);
or UO_2917 (O_2917,N_29847,N_28860);
xor UO_2918 (O_2918,N_29800,N_29297);
xor UO_2919 (O_2919,N_29208,N_29905);
xor UO_2920 (O_2920,N_29531,N_29290);
nand UO_2921 (O_2921,N_29196,N_29663);
and UO_2922 (O_2922,N_29427,N_29526);
or UO_2923 (O_2923,N_29967,N_28817);
xor UO_2924 (O_2924,N_29823,N_29787);
xnor UO_2925 (O_2925,N_29263,N_29161);
nand UO_2926 (O_2926,N_29445,N_29591);
nor UO_2927 (O_2927,N_29371,N_28973);
and UO_2928 (O_2928,N_29134,N_29785);
xnor UO_2929 (O_2929,N_29456,N_29297);
nand UO_2930 (O_2930,N_29919,N_29339);
nor UO_2931 (O_2931,N_29169,N_29411);
xnor UO_2932 (O_2932,N_28993,N_28867);
nor UO_2933 (O_2933,N_29807,N_29529);
xnor UO_2934 (O_2934,N_29155,N_29897);
nand UO_2935 (O_2935,N_28926,N_28874);
nand UO_2936 (O_2936,N_29877,N_29267);
nand UO_2937 (O_2937,N_28893,N_29745);
and UO_2938 (O_2938,N_29463,N_29010);
or UO_2939 (O_2939,N_28826,N_28845);
and UO_2940 (O_2940,N_29674,N_28904);
or UO_2941 (O_2941,N_29832,N_29171);
nand UO_2942 (O_2942,N_29909,N_29416);
and UO_2943 (O_2943,N_29200,N_28875);
nor UO_2944 (O_2944,N_29046,N_29234);
and UO_2945 (O_2945,N_28840,N_29311);
and UO_2946 (O_2946,N_29455,N_28857);
xor UO_2947 (O_2947,N_29936,N_28847);
xor UO_2948 (O_2948,N_29921,N_29432);
nand UO_2949 (O_2949,N_29657,N_28881);
or UO_2950 (O_2950,N_28928,N_29422);
or UO_2951 (O_2951,N_28975,N_29167);
nor UO_2952 (O_2952,N_28975,N_29842);
nand UO_2953 (O_2953,N_29365,N_29824);
nand UO_2954 (O_2954,N_29322,N_29978);
or UO_2955 (O_2955,N_29842,N_29111);
and UO_2956 (O_2956,N_29390,N_29072);
xnor UO_2957 (O_2957,N_28853,N_29047);
or UO_2958 (O_2958,N_29002,N_29481);
nand UO_2959 (O_2959,N_29367,N_29085);
or UO_2960 (O_2960,N_29452,N_28932);
xnor UO_2961 (O_2961,N_29418,N_29910);
nand UO_2962 (O_2962,N_28966,N_29865);
xor UO_2963 (O_2963,N_29378,N_29533);
nor UO_2964 (O_2964,N_28918,N_29592);
or UO_2965 (O_2965,N_28949,N_29544);
and UO_2966 (O_2966,N_29732,N_29150);
or UO_2967 (O_2967,N_29167,N_29832);
nor UO_2968 (O_2968,N_28806,N_29168);
or UO_2969 (O_2969,N_29021,N_29786);
xor UO_2970 (O_2970,N_29778,N_29939);
or UO_2971 (O_2971,N_29490,N_29377);
nor UO_2972 (O_2972,N_29612,N_29972);
and UO_2973 (O_2973,N_28817,N_29667);
nor UO_2974 (O_2974,N_29297,N_29438);
xnor UO_2975 (O_2975,N_29417,N_29463);
xor UO_2976 (O_2976,N_29529,N_29343);
or UO_2977 (O_2977,N_29400,N_29978);
and UO_2978 (O_2978,N_29029,N_29098);
and UO_2979 (O_2979,N_28879,N_29681);
and UO_2980 (O_2980,N_29597,N_29494);
nor UO_2981 (O_2981,N_29949,N_28852);
xor UO_2982 (O_2982,N_29741,N_29911);
nor UO_2983 (O_2983,N_29963,N_28925);
or UO_2984 (O_2984,N_29220,N_29364);
or UO_2985 (O_2985,N_28996,N_29032);
xnor UO_2986 (O_2986,N_28913,N_29772);
and UO_2987 (O_2987,N_28861,N_29264);
nand UO_2988 (O_2988,N_29815,N_29001);
nor UO_2989 (O_2989,N_28902,N_29803);
or UO_2990 (O_2990,N_28962,N_29967);
xnor UO_2991 (O_2991,N_29300,N_29643);
xor UO_2992 (O_2992,N_29842,N_29582);
and UO_2993 (O_2993,N_29726,N_29799);
nor UO_2994 (O_2994,N_29405,N_29094);
nand UO_2995 (O_2995,N_28811,N_28888);
and UO_2996 (O_2996,N_29616,N_29497);
nor UO_2997 (O_2997,N_29347,N_29554);
xor UO_2998 (O_2998,N_29297,N_28964);
and UO_2999 (O_2999,N_29837,N_29291);
and UO_3000 (O_3000,N_29528,N_28834);
nor UO_3001 (O_3001,N_29963,N_29189);
and UO_3002 (O_3002,N_29982,N_28849);
nand UO_3003 (O_3003,N_29155,N_29455);
nand UO_3004 (O_3004,N_28823,N_29491);
nor UO_3005 (O_3005,N_29010,N_28909);
and UO_3006 (O_3006,N_28974,N_29872);
nor UO_3007 (O_3007,N_29583,N_29059);
and UO_3008 (O_3008,N_29834,N_28840);
nor UO_3009 (O_3009,N_29759,N_29063);
or UO_3010 (O_3010,N_28853,N_29693);
or UO_3011 (O_3011,N_29462,N_29211);
nand UO_3012 (O_3012,N_28835,N_29217);
nand UO_3013 (O_3013,N_29235,N_29240);
or UO_3014 (O_3014,N_29926,N_29447);
xnor UO_3015 (O_3015,N_29119,N_28949);
nor UO_3016 (O_3016,N_29793,N_29744);
and UO_3017 (O_3017,N_29897,N_29926);
or UO_3018 (O_3018,N_29120,N_29246);
xor UO_3019 (O_3019,N_29455,N_29260);
nand UO_3020 (O_3020,N_29573,N_28916);
xnor UO_3021 (O_3021,N_29140,N_29407);
nor UO_3022 (O_3022,N_28888,N_29502);
and UO_3023 (O_3023,N_29246,N_29060);
xnor UO_3024 (O_3024,N_29905,N_28912);
nor UO_3025 (O_3025,N_29413,N_29435);
xnor UO_3026 (O_3026,N_29073,N_29145);
or UO_3027 (O_3027,N_29488,N_29191);
xnor UO_3028 (O_3028,N_29554,N_28974);
nand UO_3029 (O_3029,N_29552,N_29418);
nor UO_3030 (O_3030,N_29749,N_29819);
nor UO_3031 (O_3031,N_29863,N_28893);
xor UO_3032 (O_3032,N_29203,N_29841);
or UO_3033 (O_3033,N_29778,N_29667);
nor UO_3034 (O_3034,N_28925,N_28801);
nand UO_3035 (O_3035,N_29953,N_28899);
nor UO_3036 (O_3036,N_29318,N_28990);
or UO_3037 (O_3037,N_29682,N_29595);
or UO_3038 (O_3038,N_29502,N_29098);
nand UO_3039 (O_3039,N_29491,N_29220);
or UO_3040 (O_3040,N_29550,N_29912);
or UO_3041 (O_3041,N_29411,N_29983);
nor UO_3042 (O_3042,N_29376,N_29037);
xor UO_3043 (O_3043,N_29466,N_29739);
nor UO_3044 (O_3044,N_29369,N_29420);
nor UO_3045 (O_3045,N_29750,N_28959);
or UO_3046 (O_3046,N_29673,N_29973);
nor UO_3047 (O_3047,N_29266,N_29341);
nor UO_3048 (O_3048,N_29856,N_29109);
and UO_3049 (O_3049,N_29946,N_28970);
xor UO_3050 (O_3050,N_29392,N_29964);
nand UO_3051 (O_3051,N_29923,N_29404);
or UO_3052 (O_3052,N_28974,N_29107);
or UO_3053 (O_3053,N_29486,N_29106);
or UO_3054 (O_3054,N_29294,N_29385);
or UO_3055 (O_3055,N_29175,N_29964);
xor UO_3056 (O_3056,N_28825,N_29474);
and UO_3057 (O_3057,N_29064,N_29619);
xnor UO_3058 (O_3058,N_29779,N_29768);
nor UO_3059 (O_3059,N_29921,N_29894);
xor UO_3060 (O_3060,N_29316,N_29077);
and UO_3061 (O_3061,N_29086,N_29841);
or UO_3062 (O_3062,N_29038,N_29749);
nand UO_3063 (O_3063,N_28982,N_29520);
xnor UO_3064 (O_3064,N_29495,N_29513);
nor UO_3065 (O_3065,N_28866,N_29807);
nor UO_3066 (O_3066,N_29181,N_29021);
and UO_3067 (O_3067,N_29649,N_29725);
xnor UO_3068 (O_3068,N_28973,N_29002);
nand UO_3069 (O_3069,N_29053,N_29302);
and UO_3070 (O_3070,N_28831,N_29479);
xnor UO_3071 (O_3071,N_28962,N_29835);
or UO_3072 (O_3072,N_29178,N_29830);
and UO_3073 (O_3073,N_28824,N_29634);
xor UO_3074 (O_3074,N_29170,N_29629);
nand UO_3075 (O_3075,N_29936,N_29784);
nand UO_3076 (O_3076,N_28888,N_29599);
and UO_3077 (O_3077,N_29534,N_29181);
or UO_3078 (O_3078,N_28946,N_29029);
xor UO_3079 (O_3079,N_29300,N_29887);
nor UO_3080 (O_3080,N_29243,N_29749);
nor UO_3081 (O_3081,N_29661,N_29917);
xnor UO_3082 (O_3082,N_29357,N_29890);
nand UO_3083 (O_3083,N_29985,N_29350);
and UO_3084 (O_3084,N_29192,N_29590);
xor UO_3085 (O_3085,N_29221,N_29715);
nand UO_3086 (O_3086,N_29344,N_29314);
nand UO_3087 (O_3087,N_29736,N_29076);
or UO_3088 (O_3088,N_29615,N_29735);
and UO_3089 (O_3089,N_29259,N_29935);
or UO_3090 (O_3090,N_29122,N_29769);
nor UO_3091 (O_3091,N_29151,N_29962);
or UO_3092 (O_3092,N_29298,N_29242);
nor UO_3093 (O_3093,N_29880,N_29327);
nor UO_3094 (O_3094,N_29884,N_29037);
or UO_3095 (O_3095,N_29684,N_29053);
and UO_3096 (O_3096,N_29426,N_29834);
or UO_3097 (O_3097,N_29245,N_29324);
nand UO_3098 (O_3098,N_29140,N_29673);
nor UO_3099 (O_3099,N_29893,N_29207);
or UO_3100 (O_3100,N_28981,N_29689);
and UO_3101 (O_3101,N_29408,N_29007);
or UO_3102 (O_3102,N_29291,N_29299);
and UO_3103 (O_3103,N_29833,N_29876);
or UO_3104 (O_3104,N_29621,N_29453);
xor UO_3105 (O_3105,N_29928,N_29670);
xor UO_3106 (O_3106,N_29892,N_29015);
or UO_3107 (O_3107,N_29749,N_29710);
and UO_3108 (O_3108,N_29504,N_29155);
xor UO_3109 (O_3109,N_29367,N_28891);
nand UO_3110 (O_3110,N_29914,N_29482);
nor UO_3111 (O_3111,N_29988,N_29487);
xnor UO_3112 (O_3112,N_29347,N_29053);
nor UO_3113 (O_3113,N_29552,N_29369);
xor UO_3114 (O_3114,N_29156,N_29879);
nor UO_3115 (O_3115,N_29939,N_29492);
nor UO_3116 (O_3116,N_29164,N_29861);
xor UO_3117 (O_3117,N_29726,N_29640);
nor UO_3118 (O_3118,N_29103,N_29932);
nand UO_3119 (O_3119,N_29616,N_28917);
and UO_3120 (O_3120,N_28851,N_29461);
and UO_3121 (O_3121,N_29924,N_29463);
and UO_3122 (O_3122,N_29325,N_29508);
nor UO_3123 (O_3123,N_29878,N_29873);
nor UO_3124 (O_3124,N_29137,N_29242);
nand UO_3125 (O_3125,N_29585,N_29883);
xor UO_3126 (O_3126,N_29794,N_29974);
and UO_3127 (O_3127,N_28850,N_29551);
nand UO_3128 (O_3128,N_28938,N_29764);
and UO_3129 (O_3129,N_29385,N_29500);
nor UO_3130 (O_3130,N_29360,N_28877);
nor UO_3131 (O_3131,N_29105,N_29765);
and UO_3132 (O_3132,N_29772,N_28916);
or UO_3133 (O_3133,N_28928,N_29656);
nand UO_3134 (O_3134,N_29515,N_29301);
nor UO_3135 (O_3135,N_29480,N_29695);
nand UO_3136 (O_3136,N_29740,N_28894);
xnor UO_3137 (O_3137,N_29873,N_29958);
and UO_3138 (O_3138,N_29560,N_29624);
xor UO_3139 (O_3139,N_29194,N_29339);
and UO_3140 (O_3140,N_28913,N_29798);
nor UO_3141 (O_3141,N_29645,N_29616);
or UO_3142 (O_3142,N_29849,N_28876);
or UO_3143 (O_3143,N_28970,N_29473);
and UO_3144 (O_3144,N_29690,N_29344);
xnor UO_3145 (O_3145,N_29713,N_29346);
and UO_3146 (O_3146,N_29351,N_29327);
or UO_3147 (O_3147,N_29979,N_29421);
or UO_3148 (O_3148,N_28999,N_29830);
xor UO_3149 (O_3149,N_29289,N_29887);
xor UO_3150 (O_3150,N_29502,N_29439);
nor UO_3151 (O_3151,N_29262,N_29937);
nor UO_3152 (O_3152,N_28944,N_28839);
nand UO_3153 (O_3153,N_29362,N_29198);
or UO_3154 (O_3154,N_29883,N_29522);
nor UO_3155 (O_3155,N_29178,N_29177);
or UO_3156 (O_3156,N_29310,N_29574);
nor UO_3157 (O_3157,N_28801,N_28940);
nand UO_3158 (O_3158,N_29234,N_29164);
xnor UO_3159 (O_3159,N_29250,N_29633);
and UO_3160 (O_3160,N_29910,N_29985);
nor UO_3161 (O_3161,N_29786,N_29566);
nor UO_3162 (O_3162,N_29172,N_29822);
or UO_3163 (O_3163,N_29940,N_29174);
nor UO_3164 (O_3164,N_29452,N_28888);
nand UO_3165 (O_3165,N_29257,N_29027);
or UO_3166 (O_3166,N_29696,N_28926);
nor UO_3167 (O_3167,N_28866,N_29541);
xnor UO_3168 (O_3168,N_29370,N_29886);
xnor UO_3169 (O_3169,N_29311,N_29623);
nor UO_3170 (O_3170,N_29094,N_29067);
nand UO_3171 (O_3171,N_29814,N_29966);
and UO_3172 (O_3172,N_29316,N_29164);
nor UO_3173 (O_3173,N_29410,N_29903);
nand UO_3174 (O_3174,N_29304,N_29900);
nor UO_3175 (O_3175,N_29769,N_29694);
xnor UO_3176 (O_3176,N_29557,N_29070);
xor UO_3177 (O_3177,N_29997,N_29048);
or UO_3178 (O_3178,N_29393,N_29085);
nand UO_3179 (O_3179,N_29181,N_29757);
nor UO_3180 (O_3180,N_29579,N_29950);
nor UO_3181 (O_3181,N_28855,N_29021);
and UO_3182 (O_3182,N_28936,N_29925);
or UO_3183 (O_3183,N_29547,N_29923);
xor UO_3184 (O_3184,N_29817,N_29953);
nor UO_3185 (O_3185,N_29068,N_29033);
xor UO_3186 (O_3186,N_28818,N_28973);
nand UO_3187 (O_3187,N_29647,N_28910);
or UO_3188 (O_3188,N_29828,N_29806);
and UO_3189 (O_3189,N_29573,N_29204);
xnor UO_3190 (O_3190,N_29821,N_29348);
and UO_3191 (O_3191,N_29937,N_29916);
xnor UO_3192 (O_3192,N_29213,N_28865);
xor UO_3193 (O_3193,N_29764,N_29793);
and UO_3194 (O_3194,N_29848,N_29317);
and UO_3195 (O_3195,N_29296,N_29193);
and UO_3196 (O_3196,N_29652,N_29055);
and UO_3197 (O_3197,N_28999,N_29866);
nor UO_3198 (O_3198,N_29724,N_28967);
nor UO_3199 (O_3199,N_28820,N_29194);
or UO_3200 (O_3200,N_29817,N_29492);
nand UO_3201 (O_3201,N_29989,N_29056);
and UO_3202 (O_3202,N_29557,N_29424);
or UO_3203 (O_3203,N_29766,N_29227);
nand UO_3204 (O_3204,N_29470,N_29515);
xnor UO_3205 (O_3205,N_29957,N_29205);
and UO_3206 (O_3206,N_29802,N_29034);
nor UO_3207 (O_3207,N_28948,N_29209);
nor UO_3208 (O_3208,N_29799,N_29508);
nor UO_3209 (O_3209,N_29706,N_29910);
nor UO_3210 (O_3210,N_28944,N_29769);
xnor UO_3211 (O_3211,N_28998,N_29242);
xor UO_3212 (O_3212,N_28863,N_29517);
or UO_3213 (O_3213,N_29348,N_29540);
or UO_3214 (O_3214,N_29924,N_29701);
nand UO_3215 (O_3215,N_28825,N_29839);
and UO_3216 (O_3216,N_28959,N_29325);
or UO_3217 (O_3217,N_29906,N_29177);
nor UO_3218 (O_3218,N_29705,N_29271);
nor UO_3219 (O_3219,N_29937,N_29025);
nor UO_3220 (O_3220,N_29200,N_29451);
nor UO_3221 (O_3221,N_28922,N_29144);
or UO_3222 (O_3222,N_29337,N_29557);
nor UO_3223 (O_3223,N_29539,N_29813);
nand UO_3224 (O_3224,N_28951,N_29546);
nor UO_3225 (O_3225,N_29091,N_29400);
nand UO_3226 (O_3226,N_28980,N_29916);
and UO_3227 (O_3227,N_29218,N_29052);
and UO_3228 (O_3228,N_29868,N_28944);
nand UO_3229 (O_3229,N_29608,N_29009);
xor UO_3230 (O_3230,N_29575,N_29369);
and UO_3231 (O_3231,N_29473,N_29925);
nand UO_3232 (O_3232,N_29713,N_28823);
nor UO_3233 (O_3233,N_29149,N_29829);
nand UO_3234 (O_3234,N_29875,N_29738);
xor UO_3235 (O_3235,N_29829,N_29837);
nand UO_3236 (O_3236,N_29924,N_29708);
or UO_3237 (O_3237,N_29148,N_29373);
nor UO_3238 (O_3238,N_29178,N_29114);
nor UO_3239 (O_3239,N_29811,N_29442);
nand UO_3240 (O_3240,N_28955,N_29085);
nand UO_3241 (O_3241,N_29489,N_28888);
nor UO_3242 (O_3242,N_29415,N_29933);
xnor UO_3243 (O_3243,N_29340,N_29676);
nor UO_3244 (O_3244,N_28872,N_29539);
xor UO_3245 (O_3245,N_29032,N_29143);
and UO_3246 (O_3246,N_29333,N_29650);
nand UO_3247 (O_3247,N_29109,N_29168);
nand UO_3248 (O_3248,N_29688,N_29535);
nor UO_3249 (O_3249,N_29050,N_29738);
xor UO_3250 (O_3250,N_28842,N_29256);
nor UO_3251 (O_3251,N_29762,N_29393);
and UO_3252 (O_3252,N_29338,N_29667);
nand UO_3253 (O_3253,N_28933,N_29314);
xnor UO_3254 (O_3254,N_29949,N_29441);
or UO_3255 (O_3255,N_29324,N_29890);
or UO_3256 (O_3256,N_29295,N_29595);
xnor UO_3257 (O_3257,N_29658,N_29615);
nand UO_3258 (O_3258,N_29068,N_29955);
nand UO_3259 (O_3259,N_29932,N_28808);
xor UO_3260 (O_3260,N_29122,N_29399);
nor UO_3261 (O_3261,N_28965,N_29211);
and UO_3262 (O_3262,N_29130,N_29863);
xor UO_3263 (O_3263,N_29859,N_28861);
xnor UO_3264 (O_3264,N_28982,N_29768);
nor UO_3265 (O_3265,N_29186,N_28883);
or UO_3266 (O_3266,N_29487,N_29435);
nand UO_3267 (O_3267,N_29205,N_29396);
nand UO_3268 (O_3268,N_29616,N_29184);
nand UO_3269 (O_3269,N_29780,N_29670);
nand UO_3270 (O_3270,N_29419,N_29205);
nor UO_3271 (O_3271,N_29647,N_29465);
xor UO_3272 (O_3272,N_29580,N_29622);
and UO_3273 (O_3273,N_29004,N_29818);
or UO_3274 (O_3274,N_29983,N_29558);
nor UO_3275 (O_3275,N_29275,N_29488);
or UO_3276 (O_3276,N_29012,N_29050);
and UO_3277 (O_3277,N_28815,N_29101);
and UO_3278 (O_3278,N_28893,N_29638);
and UO_3279 (O_3279,N_29387,N_29076);
xnor UO_3280 (O_3280,N_29736,N_28949);
and UO_3281 (O_3281,N_29965,N_29257);
nor UO_3282 (O_3282,N_29327,N_29223);
nand UO_3283 (O_3283,N_29232,N_29273);
nand UO_3284 (O_3284,N_29039,N_29826);
and UO_3285 (O_3285,N_29548,N_29974);
or UO_3286 (O_3286,N_29997,N_29283);
xor UO_3287 (O_3287,N_29266,N_29537);
xor UO_3288 (O_3288,N_29932,N_29797);
xor UO_3289 (O_3289,N_29989,N_29539);
nor UO_3290 (O_3290,N_29356,N_29960);
nor UO_3291 (O_3291,N_29237,N_28824);
and UO_3292 (O_3292,N_29940,N_29265);
xnor UO_3293 (O_3293,N_28964,N_28866);
nand UO_3294 (O_3294,N_29067,N_29954);
or UO_3295 (O_3295,N_28901,N_28849);
xnor UO_3296 (O_3296,N_29876,N_29650);
or UO_3297 (O_3297,N_29810,N_29654);
nand UO_3298 (O_3298,N_29663,N_29877);
and UO_3299 (O_3299,N_29665,N_29293);
or UO_3300 (O_3300,N_28952,N_29109);
nor UO_3301 (O_3301,N_29242,N_29526);
or UO_3302 (O_3302,N_28817,N_29597);
xor UO_3303 (O_3303,N_29033,N_28874);
and UO_3304 (O_3304,N_29985,N_29679);
nor UO_3305 (O_3305,N_29260,N_29457);
nor UO_3306 (O_3306,N_28904,N_29337);
and UO_3307 (O_3307,N_29860,N_29051);
and UO_3308 (O_3308,N_29640,N_29009);
and UO_3309 (O_3309,N_29951,N_29926);
or UO_3310 (O_3310,N_29681,N_29112);
xor UO_3311 (O_3311,N_28924,N_28911);
nand UO_3312 (O_3312,N_29146,N_29988);
and UO_3313 (O_3313,N_29852,N_29286);
and UO_3314 (O_3314,N_29639,N_29985);
nand UO_3315 (O_3315,N_29062,N_29891);
nor UO_3316 (O_3316,N_29064,N_29613);
nand UO_3317 (O_3317,N_28869,N_29148);
nor UO_3318 (O_3318,N_29173,N_29861);
or UO_3319 (O_3319,N_28925,N_29514);
nor UO_3320 (O_3320,N_29608,N_29356);
or UO_3321 (O_3321,N_29681,N_29212);
xor UO_3322 (O_3322,N_29011,N_29434);
xnor UO_3323 (O_3323,N_29464,N_28915);
xnor UO_3324 (O_3324,N_29788,N_29759);
or UO_3325 (O_3325,N_29915,N_29080);
xnor UO_3326 (O_3326,N_29773,N_29247);
xnor UO_3327 (O_3327,N_29093,N_29271);
nor UO_3328 (O_3328,N_29986,N_29411);
nor UO_3329 (O_3329,N_29207,N_29894);
and UO_3330 (O_3330,N_29868,N_29469);
or UO_3331 (O_3331,N_29318,N_29801);
nand UO_3332 (O_3332,N_28898,N_28941);
or UO_3333 (O_3333,N_29359,N_29984);
xor UO_3334 (O_3334,N_29733,N_29042);
nand UO_3335 (O_3335,N_28888,N_29758);
and UO_3336 (O_3336,N_29786,N_28975);
or UO_3337 (O_3337,N_29381,N_29957);
or UO_3338 (O_3338,N_29737,N_29138);
nor UO_3339 (O_3339,N_29831,N_29712);
nor UO_3340 (O_3340,N_29100,N_29262);
and UO_3341 (O_3341,N_29308,N_29635);
or UO_3342 (O_3342,N_29422,N_29595);
or UO_3343 (O_3343,N_29036,N_28810);
nor UO_3344 (O_3344,N_29183,N_29882);
or UO_3345 (O_3345,N_29536,N_29521);
nor UO_3346 (O_3346,N_29125,N_29478);
or UO_3347 (O_3347,N_29510,N_29141);
and UO_3348 (O_3348,N_28983,N_29638);
and UO_3349 (O_3349,N_29882,N_28980);
nor UO_3350 (O_3350,N_29123,N_29636);
nor UO_3351 (O_3351,N_29078,N_29877);
nand UO_3352 (O_3352,N_29089,N_29051);
and UO_3353 (O_3353,N_29338,N_29809);
xnor UO_3354 (O_3354,N_29074,N_29109);
or UO_3355 (O_3355,N_29096,N_29997);
nor UO_3356 (O_3356,N_29069,N_29025);
xor UO_3357 (O_3357,N_29445,N_29465);
nand UO_3358 (O_3358,N_29918,N_28877);
nand UO_3359 (O_3359,N_29062,N_29291);
or UO_3360 (O_3360,N_29659,N_29917);
nor UO_3361 (O_3361,N_29298,N_29051);
nand UO_3362 (O_3362,N_28849,N_29074);
nor UO_3363 (O_3363,N_29198,N_29749);
xor UO_3364 (O_3364,N_29384,N_28945);
nor UO_3365 (O_3365,N_29354,N_29831);
nor UO_3366 (O_3366,N_29773,N_28840);
and UO_3367 (O_3367,N_29356,N_29346);
nor UO_3368 (O_3368,N_29163,N_29681);
or UO_3369 (O_3369,N_29815,N_28920);
nand UO_3370 (O_3370,N_29135,N_29430);
nor UO_3371 (O_3371,N_28843,N_29833);
or UO_3372 (O_3372,N_29487,N_28874);
nor UO_3373 (O_3373,N_29534,N_29476);
nor UO_3374 (O_3374,N_29934,N_29603);
or UO_3375 (O_3375,N_28866,N_29698);
or UO_3376 (O_3376,N_28868,N_29177);
nand UO_3377 (O_3377,N_29034,N_29863);
and UO_3378 (O_3378,N_29688,N_29997);
and UO_3379 (O_3379,N_28828,N_29732);
or UO_3380 (O_3380,N_29375,N_28923);
xnor UO_3381 (O_3381,N_29759,N_28881);
or UO_3382 (O_3382,N_29478,N_29584);
xnor UO_3383 (O_3383,N_29603,N_29586);
nand UO_3384 (O_3384,N_29632,N_29887);
nor UO_3385 (O_3385,N_29314,N_29154);
xor UO_3386 (O_3386,N_28845,N_29350);
or UO_3387 (O_3387,N_29362,N_29587);
xor UO_3388 (O_3388,N_29289,N_29873);
nor UO_3389 (O_3389,N_29103,N_29120);
or UO_3390 (O_3390,N_29126,N_29407);
nor UO_3391 (O_3391,N_29346,N_29797);
nor UO_3392 (O_3392,N_29048,N_29765);
or UO_3393 (O_3393,N_29263,N_29913);
nand UO_3394 (O_3394,N_28904,N_29602);
nor UO_3395 (O_3395,N_28850,N_29980);
and UO_3396 (O_3396,N_29907,N_29920);
xnor UO_3397 (O_3397,N_29821,N_29944);
xnor UO_3398 (O_3398,N_29392,N_29880);
nor UO_3399 (O_3399,N_29270,N_29667);
and UO_3400 (O_3400,N_29736,N_29978);
and UO_3401 (O_3401,N_29930,N_29048);
and UO_3402 (O_3402,N_29275,N_29976);
xor UO_3403 (O_3403,N_29438,N_29147);
and UO_3404 (O_3404,N_29966,N_28931);
nand UO_3405 (O_3405,N_29159,N_29520);
nand UO_3406 (O_3406,N_29961,N_28988);
nand UO_3407 (O_3407,N_28973,N_29491);
or UO_3408 (O_3408,N_29787,N_29499);
nand UO_3409 (O_3409,N_29479,N_29468);
and UO_3410 (O_3410,N_29064,N_28995);
xor UO_3411 (O_3411,N_29484,N_29635);
nor UO_3412 (O_3412,N_29936,N_29788);
nor UO_3413 (O_3413,N_29759,N_29433);
and UO_3414 (O_3414,N_28841,N_29008);
or UO_3415 (O_3415,N_29760,N_29569);
xnor UO_3416 (O_3416,N_29801,N_29655);
or UO_3417 (O_3417,N_29152,N_29384);
or UO_3418 (O_3418,N_29226,N_29141);
nor UO_3419 (O_3419,N_29197,N_29383);
nand UO_3420 (O_3420,N_29238,N_29403);
or UO_3421 (O_3421,N_28892,N_29576);
xor UO_3422 (O_3422,N_29768,N_28930);
and UO_3423 (O_3423,N_29478,N_28819);
xor UO_3424 (O_3424,N_28891,N_29828);
nor UO_3425 (O_3425,N_29711,N_29941);
or UO_3426 (O_3426,N_29751,N_29418);
xnor UO_3427 (O_3427,N_29994,N_29378);
or UO_3428 (O_3428,N_29812,N_29103);
and UO_3429 (O_3429,N_29893,N_29838);
nand UO_3430 (O_3430,N_29150,N_29587);
nor UO_3431 (O_3431,N_29643,N_29873);
nor UO_3432 (O_3432,N_29417,N_29793);
or UO_3433 (O_3433,N_29354,N_28810);
or UO_3434 (O_3434,N_28813,N_29831);
xor UO_3435 (O_3435,N_29626,N_29639);
nor UO_3436 (O_3436,N_29600,N_29415);
xnor UO_3437 (O_3437,N_28899,N_29415);
and UO_3438 (O_3438,N_29083,N_28949);
and UO_3439 (O_3439,N_29928,N_28821);
xor UO_3440 (O_3440,N_28924,N_29979);
and UO_3441 (O_3441,N_29924,N_28948);
or UO_3442 (O_3442,N_29506,N_29113);
and UO_3443 (O_3443,N_29687,N_29654);
xnor UO_3444 (O_3444,N_29523,N_29149);
nand UO_3445 (O_3445,N_29364,N_28867);
xor UO_3446 (O_3446,N_28807,N_29679);
or UO_3447 (O_3447,N_29904,N_29178);
xnor UO_3448 (O_3448,N_29797,N_28975);
or UO_3449 (O_3449,N_29597,N_29920);
or UO_3450 (O_3450,N_29912,N_29356);
and UO_3451 (O_3451,N_28903,N_29791);
xor UO_3452 (O_3452,N_29080,N_29481);
nor UO_3453 (O_3453,N_29819,N_29557);
nand UO_3454 (O_3454,N_29274,N_28897);
nor UO_3455 (O_3455,N_29702,N_29503);
nand UO_3456 (O_3456,N_29382,N_29946);
and UO_3457 (O_3457,N_29040,N_29471);
or UO_3458 (O_3458,N_29335,N_29960);
or UO_3459 (O_3459,N_29349,N_29512);
or UO_3460 (O_3460,N_29029,N_29275);
and UO_3461 (O_3461,N_28944,N_29274);
and UO_3462 (O_3462,N_28876,N_29140);
nor UO_3463 (O_3463,N_29979,N_29085);
or UO_3464 (O_3464,N_29482,N_29332);
xnor UO_3465 (O_3465,N_29944,N_28808);
xnor UO_3466 (O_3466,N_29947,N_29158);
or UO_3467 (O_3467,N_28924,N_29768);
or UO_3468 (O_3468,N_29320,N_29762);
nor UO_3469 (O_3469,N_29686,N_29018);
or UO_3470 (O_3470,N_29708,N_29971);
nand UO_3471 (O_3471,N_29967,N_28890);
and UO_3472 (O_3472,N_29941,N_29789);
or UO_3473 (O_3473,N_29597,N_29174);
or UO_3474 (O_3474,N_29897,N_29993);
nor UO_3475 (O_3475,N_29808,N_29715);
and UO_3476 (O_3476,N_29600,N_29564);
xor UO_3477 (O_3477,N_29649,N_29385);
nor UO_3478 (O_3478,N_29596,N_29923);
xnor UO_3479 (O_3479,N_29823,N_29588);
nand UO_3480 (O_3480,N_29435,N_29767);
or UO_3481 (O_3481,N_29205,N_29760);
or UO_3482 (O_3482,N_28899,N_28946);
xnor UO_3483 (O_3483,N_29120,N_29104);
or UO_3484 (O_3484,N_29279,N_29835);
nor UO_3485 (O_3485,N_29421,N_29127);
or UO_3486 (O_3486,N_29566,N_29217);
xnor UO_3487 (O_3487,N_29938,N_29796);
or UO_3488 (O_3488,N_29669,N_29521);
or UO_3489 (O_3489,N_29806,N_28963);
nor UO_3490 (O_3490,N_28920,N_29610);
nor UO_3491 (O_3491,N_29224,N_29730);
nor UO_3492 (O_3492,N_29077,N_29243);
and UO_3493 (O_3493,N_29756,N_29695);
xnor UO_3494 (O_3494,N_29490,N_29007);
nand UO_3495 (O_3495,N_28931,N_29329);
and UO_3496 (O_3496,N_29596,N_29087);
nand UO_3497 (O_3497,N_29397,N_29474);
nor UO_3498 (O_3498,N_29668,N_28958);
nand UO_3499 (O_3499,N_29320,N_29123);
endmodule